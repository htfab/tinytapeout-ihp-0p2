module tt_um_vc32_cpu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire clknet_leaf_0_clk;
 wire \cpu.addr[10] ;
 wire \cpu.addr[11] ;
 wire \cpu.addr[12] ;
 wire \cpu.addr[13] ;
 wire \cpu.addr[14] ;
 wire \cpu.addr[15] ;
 wire \cpu.addr[1] ;
 wire \cpu.addr[2] ;
 wire \cpu.addr[3] ;
 wire \cpu.addr[4] ;
 wire \cpu.addr[5] ;
 wire \cpu.addr[6] ;
 wire \cpu.addr[7] ;
 wire \cpu.addr[8] ;
 wire \cpu.addr[9] ;
 wire \cpu.br ;
 wire \cpu.cond[0] ;
 wire \cpu.cond[1] ;
 wire \cpu.cond[2] ;
 wire \cpu.d_flush_all ;
 wire \cpu.d_rstrobe_d ;
 wire \cpu.d_wstrobe_d ;
 wire \cpu.dcache.flush_write ;
 wire \cpu.dcache.r_data[0][0] ;
 wire \cpu.dcache.r_data[0][10] ;
 wire \cpu.dcache.r_data[0][11] ;
 wire \cpu.dcache.r_data[0][12] ;
 wire \cpu.dcache.r_data[0][13] ;
 wire \cpu.dcache.r_data[0][14] ;
 wire \cpu.dcache.r_data[0][15] ;
 wire \cpu.dcache.r_data[0][16] ;
 wire \cpu.dcache.r_data[0][17] ;
 wire \cpu.dcache.r_data[0][18] ;
 wire \cpu.dcache.r_data[0][19] ;
 wire \cpu.dcache.r_data[0][1] ;
 wire \cpu.dcache.r_data[0][20] ;
 wire \cpu.dcache.r_data[0][21] ;
 wire \cpu.dcache.r_data[0][22] ;
 wire \cpu.dcache.r_data[0][23] ;
 wire \cpu.dcache.r_data[0][24] ;
 wire \cpu.dcache.r_data[0][25] ;
 wire \cpu.dcache.r_data[0][26] ;
 wire \cpu.dcache.r_data[0][27] ;
 wire \cpu.dcache.r_data[0][28] ;
 wire \cpu.dcache.r_data[0][29] ;
 wire \cpu.dcache.r_data[0][2] ;
 wire \cpu.dcache.r_data[0][30] ;
 wire \cpu.dcache.r_data[0][31] ;
 wire \cpu.dcache.r_data[0][3] ;
 wire \cpu.dcache.r_data[0][4] ;
 wire \cpu.dcache.r_data[0][5] ;
 wire \cpu.dcache.r_data[0][6] ;
 wire \cpu.dcache.r_data[0][7] ;
 wire \cpu.dcache.r_data[0][8] ;
 wire \cpu.dcache.r_data[0][9] ;
 wire \cpu.dcache.r_data[1][0] ;
 wire \cpu.dcache.r_data[1][10] ;
 wire \cpu.dcache.r_data[1][11] ;
 wire \cpu.dcache.r_data[1][12] ;
 wire \cpu.dcache.r_data[1][13] ;
 wire \cpu.dcache.r_data[1][14] ;
 wire \cpu.dcache.r_data[1][15] ;
 wire \cpu.dcache.r_data[1][16] ;
 wire \cpu.dcache.r_data[1][17] ;
 wire \cpu.dcache.r_data[1][18] ;
 wire \cpu.dcache.r_data[1][19] ;
 wire \cpu.dcache.r_data[1][1] ;
 wire \cpu.dcache.r_data[1][20] ;
 wire \cpu.dcache.r_data[1][21] ;
 wire \cpu.dcache.r_data[1][22] ;
 wire \cpu.dcache.r_data[1][23] ;
 wire \cpu.dcache.r_data[1][24] ;
 wire \cpu.dcache.r_data[1][25] ;
 wire \cpu.dcache.r_data[1][26] ;
 wire \cpu.dcache.r_data[1][27] ;
 wire \cpu.dcache.r_data[1][28] ;
 wire \cpu.dcache.r_data[1][29] ;
 wire \cpu.dcache.r_data[1][2] ;
 wire \cpu.dcache.r_data[1][30] ;
 wire \cpu.dcache.r_data[1][31] ;
 wire \cpu.dcache.r_data[1][3] ;
 wire \cpu.dcache.r_data[1][4] ;
 wire \cpu.dcache.r_data[1][5] ;
 wire \cpu.dcache.r_data[1][6] ;
 wire \cpu.dcache.r_data[1][7] ;
 wire \cpu.dcache.r_data[1][8] ;
 wire \cpu.dcache.r_data[1][9] ;
 wire \cpu.dcache.r_data[2][0] ;
 wire \cpu.dcache.r_data[2][10] ;
 wire \cpu.dcache.r_data[2][11] ;
 wire \cpu.dcache.r_data[2][12] ;
 wire \cpu.dcache.r_data[2][13] ;
 wire \cpu.dcache.r_data[2][14] ;
 wire \cpu.dcache.r_data[2][15] ;
 wire \cpu.dcache.r_data[2][16] ;
 wire \cpu.dcache.r_data[2][17] ;
 wire \cpu.dcache.r_data[2][18] ;
 wire \cpu.dcache.r_data[2][19] ;
 wire \cpu.dcache.r_data[2][1] ;
 wire \cpu.dcache.r_data[2][20] ;
 wire \cpu.dcache.r_data[2][21] ;
 wire \cpu.dcache.r_data[2][22] ;
 wire \cpu.dcache.r_data[2][23] ;
 wire \cpu.dcache.r_data[2][24] ;
 wire \cpu.dcache.r_data[2][25] ;
 wire \cpu.dcache.r_data[2][26] ;
 wire \cpu.dcache.r_data[2][27] ;
 wire \cpu.dcache.r_data[2][28] ;
 wire \cpu.dcache.r_data[2][29] ;
 wire \cpu.dcache.r_data[2][2] ;
 wire \cpu.dcache.r_data[2][30] ;
 wire \cpu.dcache.r_data[2][31] ;
 wire \cpu.dcache.r_data[2][3] ;
 wire \cpu.dcache.r_data[2][4] ;
 wire \cpu.dcache.r_data[2][5] ;
 wire \cpu.dcache.r_data[2][6] ;
 wire \cpu.dcache.r_data[2][7] ;
 wire \cpu.dcache.r_data[2][8] ;
 wire \cpu.dcache.r_data[2][9] ;
 wire \cpu.dcache.r_data[3][0] ;
 wire \cpu.dcache.r_data[3][10] ;
 wire \cpu.dcache.r_data[3][11] ;
 wire \cpu.dcache.r_data[3][12] ;
 wire \cpu.dcache.r_data[3][13] ;
 wire \cpu.dcache.r_data[3][14] ;
 wire \cpu.dcache.r_data[3][15] ;
 wire \cpu.dcache.r_data[3][16] ;
 wire \cpu.dcache.r_data[3][17] ;
 wire \cpu.dcache.r_data[3][18] ;
 wire \cpu.dcache.r_data[3][19] ;
 wire \cpu.dcache.r_data[3][1] ;
 wire \cpu.dcache.r_data[3][20] ;
 wire \cpu.dcache.r_data[3][21] ;
 wire \cpu.dcache.r_data[3][22] ;
 wire \cpu.dcache.r_data[3][23] ;
 wire \cpu.dcache.r_data[3][24] ;
 wire \cpu.dcache.r_data[3][25] ;
 wire \cpu.dcache.r_data[3][26] ;
 wire \cpu.dcache.r_data[3][27] ;
 wire \cpu.dcache.r_data[3][28] ;
 wire \cpu.dcache.r_data[3][29] ;
 wire \cpu.dcache.r_data[3][2] ;
 wire \cpu.dcache.r_data[3][30] ;
 wire \cpu.dcache.r_data[3][31] ;
 wire \cpu.dcache.r_data[3][3] ;
 wire \cpu.dcache.r_data[3][4] ;
 wire \cpu.dcache.r_data[3][5] ;
 wire \cpu.dcache.r_data[3][6] ;
 wire \cpu.dcache.r_data[3][7] ;
 wire \cpu.dcache.r_data[3][8] ;
 wire \cpu.dcache.r_data[3][9] ;
 wire \cpu.dcache.r_data[4][0] ;
 wire \cpu.dcache.r_data[4][10] ;
 wire \cpu.dcache.r_data[4][11] ;
 wire \cpu.dcache.r_data[4][12] ;
 wire \cpu.dcache.r_data[4][13] ;
 wire \cpu.dcache.r_data[4][14] ;
 wire \cpu.dcache.r_data[4][15] ;
 wire \cpu.dcache.r_data[4][16] ;
 wire \cpu.dcache.r_data[4][17] ;
 wire \cpu.dcache.r_data[4][18] ;
 wire \cpu.dcache.r_data[4][19] ;
 wire \cpu.dcache.r_data[4][1] ;
 wire \cpu.dcache.r_data[4][20] ;
 wire \cpu.dcache.r_data[4][21] ;
 wire \cpu.dcache.r_data[4][22] ;
 wire \cpu.dcache.r_data[4][23] ;
 wire \cpu.dcache.r_data[4][24] ;
 wire \cpu.dcache.r_data[4][25] ;
 wire \cpu.dcache.r_data[4][26] ;
 wire \cpu.dcache.r_data[4][27] ;
 wire \cpu.dcache.r_data[4][28] ;
 wire \cpu.dcache.r_data[4][29] ;
 wire \cpu.dcache.r_data[4][2] ;
 wire \cpu.dcache.r_data[4][30] ;
 wire \cpu.dcache.r_data[4][31] ;
 wire \cpu.dcache.r_data[4][3] ;
 wire \cpu.dcache.r_data[4][4] ;
 wire \cpu.dcache.r_data[4][5] ;
 wire \cpu.dcache.r_data[4][6] ;
 wire \cpu.dcache.r_data[4][7] ;
 wire \cpu.dcache.r_data[4][8] ;
 wire \cpu.dcache.r_data[4][9] ;
 wire \cpu.dcache.r_data[5][0] ;
 wire \cpu.dcache.r_data[5][10] ;
 wire \cpu.dcache.r_data[5][11] ;
 wire \cpu.dcache.r_data[5][12] ;
 wire \cpu.dcache.r_data[5][13] ;
 wire \cpu.dcache.r_data[5][14] ;
 wire \cpu.dcache.r_data[5][15] ;
 wire \cpu.dcache.r_data[5][16] ;
 wire \cpu.dcache.r_data[5][17] ;
 wire \cpu.dcache.r_data[5][18] ;
 wire \cpu.dcache.r_data[5][19] ;
 wire \cpu.dcache.r_data[5][1] ;
 wire \cpu.dcache.r_data[5][20] ;
 wire \cpu.dcache.r_data[5][21] ;
 wire \cpu.dcache.r_data[5][22] ;
 wire \cpu.dcache.r_data[5][23] ;
 wire \cpu.dcache.r_data[5][24] ;
 wire \cpu.dcache.r_data[5][25] ;
 wire \cpu.dcache.r_data[5][26] ;
 wire \cpu.dcache.r_data[5][27] ;
 wire \cpu.dcache.r_data[5][28] ;
 wire \cpu.dcache.r_data[5][29] ;
 wire \cpu.dcache.r_data[5][2] ;
 wire \cpu.dcache.r_data[5][30] ;
 wire \cpu.dcache.r_data[5][31] ;
 wire \cpu.dcache.r_data[5][3] ;
 wire \cpu.dcache.r_data[5][4] ;
 wire \cpu.dcache.r_data[5][5] ;
 wire \cpu.dcache.r_data[5][6] ;
 wire \cpu.dcache.r_data[5][7] ;
 wire \cpu.dcache.r_data[5][8] ;
 wire \cpu.dcache.r_data[5][9] ;
 wire \cpu.dcache.r_data[6][0] ;
 wire \cpu.dcache.r_data[6][10] ;
 wire \cpu.dcache.r_data[6][11] ;
 wire \cpu.dcache.r_data[6][12] ;
 wire \cpu.dcache.r_data[6][13] ;
 wire \cpu.dcache.r_data[6][14] ;
 wire \cpu.dcache.r_data[6][15] ;
 wire \cpu.dcache.r_data[6][16] ;
 wire \cpu.dcache.r_data[6][17] ;
 wire \cpu.dcache.r_data[6][18] ;
 wire \cpu.dcache.r_data[6][19] ;
 wire \cpu.dcache.r_data[6][1] ;
 wire \cpu.dcache.r_data[6][20] ;
 wire \cpu.dcache.r_data[6][21] ;
 wire \cpu.dcache.r_data[6][22] ;
 wire \cpu.dcache.r_data[6][23] ;
 wire \cpu.dcache.r_data[6][24] ;
 wire \cpu.dcache.r_data[6][25] ;
 wire \cpu.dcache.r_data[6][26] ;
 wire \cpu.dcache.r_data[6][27] ;
 wire \cpu.dcache.r_data[6][28] ;
 wire \cpu.dcache.r_data[6][29] ;
 wire \cpu.dcache.r_data[6][2] ;
 wire \cpu.dcache.r_data[6][30] ;
 wire \cpu.dcache.r_data[6][31] ;
 wire \cpu.dcache.r_data[6][3] ;
 wire \cpu.dcache.r_data[6][4] ;
 wire \cpu.dcache.r_data[6][5] ;
 wire \cpu.dcache.r_data[6][6] ;
 wire \cpu.dcache.r_data[6][7] ;
 wire \cpu.dcache.r_data[6][8] ;
 wire \cpu.dcache.r_data[6][9] ;
 wire \cpu.dcache.r_data[7][0] ;
 wire \cpu.dcache.r_data[7][10] ;
 wire \cpu.dcache.r_data[7][11] ;
 wire \cpu.dcache.r_data[7][12] ;
 wire \cpu.dcache.r_data[7][13] ;
 wire \cpu.dcache.r_data[7][14] ;
 wire \cpu.dcache.r_data[7][15] ;
 wire \cpu.dcache.r_data[7][16] ;
 wire \cpu.dcache.r_data[7][17] ;
 wire \cpu.dcache.r_data[7][18] ;
 wire \cpu.dcache.r_data[7][19] ;
 wire \cpu.dcache.r_data[7][1] ;
 wire \cpu.dcache.r_data[7][20] ;
 wire \cpu.dcache.r_data[7][21] ;
 wire \cpu.dcache.r_data[7][22] ;
 wire \cpu.dcache.r_data[7][23] ;
 wire \cpu.dcache.r_data[7][24] ;
 wire \cpu.dcache.r_data[7][25] ;
 wire \cpu.dcache.r_data[7][26] ;
 wire \cpu.dcache.r_data[7][27] ;
 wire \cpu.dcache.r_data[7][28] ;
 wire \cpu.dcache.r_data[7][29] ;
 wire \cpu.dcache.r_data[7][2] ;
 wire \cpu.dcache.r_data[7][30] ;
 wire \cpu.dcache.r_data[7][31] ;
 wire \cpu.dcache.r_data[7][3] ;
 wire \cpu.dcache.r_data[7][4] ;
 wire \cpu.dcache.r_data[7][5] ;
 wire \cpu.dcache.r_data[7][6] ;
 wire \cpu.dcache.r_data[7][7] ;
 wire \cpu.dcache.r_data[7][8] ;
 wire \cpu.dcache.r_data[7][9] ;
 wire \cpu.dcache.r_dirty[0] ;
 wire \cpu.dcache.r_dirty[1] ;
 wire \cpu.dcache.r_dirty[2] ;
 wire \cpu.dcache.r_dirty[3] ;
 wire \cpu.dcache.r_dirty[4] ;
 wire \cpu.dcache.r_dirty[5] ;
 wire \cpu.dcache.r_dirty[6] ;
 wire \cpu.dcache.r_dirty[7] ;
 wire \cpu.dcache.r_offset[0] ;
 wire \cpu.dcache.r_offset[1] ;
 wire \cpu.dcache.r_offset[2] ;
 wire \cpu.dcache.r_tag[0][10] ;
 wire \cpu.dcache.r_tag[0][11] ;
 wire \cpu.dcache.r_tag[0][12] ;
 wire \cpu.dcache.r_tag[0][13] ;
 wire \cpu.dcache.r_tag[0][14] ;
 wire \cpu.dcache.r_tag[0][15] ;
 wire \cpu.dcache.r_tag[0][16] ;
 wire \cpu.dcache.r_tag[0][17] ;
 wire \cpu.dcache.r_tag[0][18] ;
 wire \cpu.dcache.r_tag[0][19] ;
 wire \cpu.dcache.r_tag[0][20] ;
 wire \cpu.dcache.r_tag[0][21] ;
 wire \cpu.dcache.r_tag[0][22] ;
 wire \cpu.dcache.r_tag[0][23] ;
 wire \cpu.dcache.r_tag[0][5] ;
 wire \cpu.dcache.r_tag[0][6] ;
 wire \cpu.dcache.r_tag[0][7] ;
 wire \cpu.dcache.r_tag[0][8] ;
 wire \cpu.dcache.r_tag[0][9] ;
 wire \cpu.dcache.r_tag[1][10] ;
 wire \cpu.dcache.r_tag[1][11] ;
 wire \cpu.dcache.r_tag[1][12] ;
 wire \cpu.dcache.r_tag[1][13] ;
 wire \cpu.dcache.r_tag[1][14] ;
 wire \cpu.dcache.r_tag[1][15] ;
 wire \cpu.dcache.r_tag[1][16] ;
 wire \cpu.dcache.r_tag[1][17] ;
 wire \cpu.dcache.r_tag[1][18] ;
 wire \cpu.dcache.r_tag[1][19] ;
 wire \cpu.dcache.r_tag[1][20] ;
 wire \cpu.dcache.r_tag[1][21] ;
 wire \cpu.dcache.r_tag[1][22] ;
 wire \cpu.dcache.r_tag[1][23] ;
 wire \cpu.dcache.r_tag[1][5] ;
 wire \cpu.dcache.r_tag[1][6] ;
 wire \cpu.dcache.r_tag[1][7] ;
 wire \cpu.dcache.r_tag[1][8] ;
 wire \cpu.dcache.r_tag[1][9] ;
 wire \cpu.dcache.r_tag[2][10] ;
 wire \cpu.dcache.r_tag[2][11] ;
 wire \cpu.dcache.r_tag[2][12] ;
 wire \cpu.dcache.r_tag[2][13] ;
 wire \cpu.dcache.r_tag[2][14] ;
 wire \cpu.dcache.r_tag[2][15] ;
 wire \cpu.dcache.r_tag[2][16] ;
 wire \cpu.dcache.r_tag[2][17] ;
 wire \cpu.dcache.r_tag[2][18] ;
 wire \cpu.dcache.r_tag[2][19] ;
 wire \cpu.dcache.r_tag[2][20] ;
 wire \cpu.dcache.r_tag[2][21] ;
 wire \cpu.dcache.r_tag[2][22] ;
 wire \cpu.dcache.r_tag[2][23] ;
 wire \cpu.dcache.r_tag[2][5] ;
 wire \cpu.dcache.r_tag[2][6] ;
 wire \cpu.dcache.r_tag[2][7] ;
 wire \cpu.dcache.r_tag[2][8] ;
 wire \cpu.dcache.r_tag[2][9] ;
 wire \cpu.dcache.r_tag[3][10] ;
 wire \cpu.dcache.r_tag[3][11] ;
 wire \cpu.dcache.r_tag[3][12] ;
 wire \cpu.dcache.r_tag[3][13] ;
 wire \cpu.dcache.r_tag[3][14] ;
 wire \cpu.dcache.r_tag[3][15] ;
 wire \cpu.dcache.r_tag[3][16] ;
 wire \cpu.dcache.r_tag[3][17] ;
 wire \cpu.dcache.r_tag[3][18] ;
 wire \cpu.dcache.r_tag[3][19] ;
 wire \cpu.dcache.r_tag[3][20] ;
 wire \cpu.dcache.r_tag[3][21] ;
 wire \cpu.dcache.r_tag[3][22] ;
 wire \cpu.dcache.r_tag[3][23] ;
 wire \cpu.dcache.r_tag[3][5] ;
 wire \cpu.dcache.r_tag[3][6] ;
 wire \cpu.dcache.r_tag[3][7] ;
 wire \cpu.dcache.r_tag[3][8] ;
 wire \cpu.dcache.r_tag[3][9] ;
 wire \cpu.dcache.r_tag[4][10] ;
 wire \cpu.dcache.r_tag[4][11] ;
 wire \cpu.dcache.r_tag[4][12] ;
 wire \cpu.dcache.r_tag[4][13] ;
 wire \cpu.dcache.r_tag[4][14] ;
 wire \cpu.dcache.r_tag[4][15] ;
 wire \cpu.dcache.r_tag[4][16] ;
 wire \cpu.dcache.r_tag[4][17] ;
 wire \cpu.dcache.r_tag[4][18] ;
 wire \cpu.dcache.r_tag[4][19] ;
 wire \cpu.dcache.r_tag[4][20] ;
 wire \cpu.dcache.r_tag[4][21] ;
 wire \cpu.dcache.r_tag[4][22] ;
 wire \cpu.dcache.r_tag[4][23] ;
 wire \cpu.dcache.r_tag[4][5] ;
 wire \cpu.dcache.r_tag[4][6] ;
 wire \cpu.dcache.r_tag[4][7] ;
 wire \cpu.dcache.r_tag[4][8] ;
 wire \cpu.dcache.r_tag[4][9] ;
 wire \cpu.dcache.r_tag[5][10] ;
 wire \cpu.dcache.r_tag[5][11] ;
 wire \cpu.dcache.r_tag[5][12] ;
 wire \cpu.dcache.r_tag[5][13] ;
 wire \cpu.dcache.r_tag[5][14] ;
 wire \cpu.dcache.r_tag[5][15] ;
 wire \cpu.dcache.r_tag[5][16] ;
 wire \cpu.dcache.r_tag[5][17] ;
 wire \cpu.dcache.r_tag[5][18] ;
 wire \cpu.dcache.r_tag[5][19] ;
 wire \cpu.dcache.r_tag[5][20] ;
 wire \cpu.dcache.r_tag[5][21] ;
 wire \cpu.dcache.r_tag[5][22] ;
 wire \cpu.dcache.r_tag[5][23] ;
 wire \cpu.dcache.r_tag[5][5] ;
 wire \cpu.dcache.r_tag[5][6] ;
 wire \cpu.dcache.r_tag[5][7] ;
 wire \cpu.dcache.r_tag[5][8] ;
 wire \cpu.dcache.r_tag[5][9] ;
 wire \cpu.dcache.r_tag[6][10] ;
 wire \cpu.dcache.r_tag[6][11] ;
 wire \cpu.dcache.r_tag[6][12] ;
 wire \cpu.dcache.r_tag[6][13] ;
 wire \cpu.dcache.r_tag[6][14] ;
 wire \cpu.dcache.r_tag[6][15] ;
 wire \cpu.dcache.r_tag[6][16] ;
 wire \cpu.dcache.r_tag[6][17] ;
 wire \cpu.dcache.r_tag[6][18] ;
 wire \cpu.dcache.r_tag[6][19] ;
 wire \cpu.dcache.r_tag[6][20] ;
 wire \cpu.dcache.r_tag[6][21] ;
 wire \cpu.dcache.r_tag[6][22] ;
 wire \cpu.dcache.r_tag[6][23] ;
 wire \cpu.dcache.r_tag[6][5] ;
 wire \cpu.dcache.r_tag[6][6] ;
 wire \cpu.dcache.r_tag[6][7] ;
 wire \cpu.dcache.r_tag[6][8] ;
 wire \cpu.dcache.r_tag[6][9] ;
 wire \cpu.dcache.r_tag[7][10] ;
 wire \cpu.dcache.r_tag[7][11] ;
 wire \cpu.dcache.r_tag[7][12] ;
 wire \cpu.dcache.r_tag[7][13] ;
 wire \cpu.dcache.r_tag[7][14] ;
 wire \cpu.dcache.r_tag[7][15] ;
 wire \cpu.dcache.r_tag[7][16] ;
 wire \cpu.dcache.r_tag[7][17] ;
 wire \cpu.dcache.r_tag[7][18] ;
 wire \cpu.dcache.r_tag[7][19] ;
 wire \cpu.dcache.r_tag[7][20] ;
 wire \cpu.dcache.r_tag[7][21] ;
 wire \cpu.dcache.r_tag[7][22] ;
 wire \cpu.dcache.r_tag[7][23] ;
 wire \cpu.dcache.r_tag[7][5] ;
 wire \cpu.dcache.r_tag[7][6] ;
 wire \cpu.dcache.r_tag[7][7] ;
 wire \cpu.dcache.r_tag[7][8] ;
 wire \cpu.dcache.r_tag[7][9] ;
 wire \cpu.dcache.r_valid[0] ;
 wire \cpu.dcache.r_valid[1] ;
 wire \cpu.dcache.r_valid[2] ;
 wire \cpu.dcache.r_valid[3] ;
 wire \cpu.dcache.r_valid[4] ;
 wire \cpu.dcache.r_valid[5] ;
 wire \cpu.dcache.r_valid[6] ;
 wire \cpu.dcache.r_valid[7] ;
 wire \cpu.dcache.wdata[0] ;
 wire \cpu.dcache.wdata[10] ;
 wire \cpu.dcache.wdata[11] ;
 wire \cpu.dcache.wdata[12] ;
 wire \cpu.dcache.wdata[13] ;
 wire \cpu.dcache.wdata[14] ;
 wire \cpu.dcache.wdata[15] ;
 wire \cpu.dcache.wdata[1] ;
 wire \cpu.dcache.wdata[2] ;
 wire \cpu.dcache.wdata[3] ;
 wire \cpu.dcache.wdata[4] ;
 wire \cpu.dcache.wdata[5] ;
 wire \cpu.dcache.wdata[6] ;
 wire \cpu.dcache.wdata[7] ;
 wire \cpu.dcache.wdata[8] ;
 wire \cpu.dcache.wdata[9] ;
 wire \cpu.dec.div ;
 wire \cpu.dec.do_flush_all ;
 wire \cpu.dec.do_flush_write ;
 wire \cpu.dec.do_inv_mmu ;
 wire \cpu.dec.imm[0] ;
 wire \cpu.dec.imm[10] ;
 wire \cpu.dec.imm[11] ;
 wire \cpu.dec.imm[12] ;
 wire \cpu.dec.imm[13] ;
 wire \cpu.dec.imm[14] ;
 wire \cpu.dec.imm[15] ;
 wire \cpu.dec.imm[1] ;
 wire \cpu.dec.imm[2] ;
 wire \cpu.dec.imm[3] ;
 wire \cpu.dec.imm[4] ;
 wire \cpu.dec.imm[5] ;
 wire \cpu.dec.imm[6] ;
 wire \cpu.dec.imm[7] ;
 wire \cpu.dec.imm[8] ;
 wire \cpu.dec.imm[9] ;
 wire \cpu.dec.io ;
 wire \cpu.dec.iready ;
 wire \cpu.dec.jmp ;
 wire \cpu.dec.load ;
 wire \cpu.dec.mult ;
 wire \cpu.dec.needs_rs2 ;
 wire \cpu.dec.r_op[10] ;
 wire \cpu.dec.r_op[1] ;
 wire \cpu.dec.r_op[2] ;
 wire \cpu.dec.r_op[3] ;
 wire \cpu.dec.r_op[4] ;
 wire \cpu.dec.r_op[5] ;
 wire \cpu.dec.r_op[6] ;
 wire \cpu.dec.r_op[7] ;
 wire \cpu.dec.r_op[8] ;
 wire \cpu.dec.r_op[9] ;
 wire \cpu.dec.r_rd[0] ;
 wire \cpu.dec.r_rd[1] ;
 wire \cpu.dec.r_rd[2] ;
 wire \cpu.dec.r_rd[3] ;
 wire \cpu.dec.r_rs1[0] ;
 wire \cpu.dec.r_rs1[1] ;
 wire \cpu.dec.r_rs1[2] ;
 wire \cpu.dec.r_rs1[3] ;
 wire \cpu.dec.r_rs2[0] ;
 wire \cpu.dec.r_rs2[1] ;
 wire \cpu.dec.r_rs2[2] ;
 wire \cpu.dec.r_rs2[3] ;
 wire \cpu.dec.r_rs2_inv ;
 wire \cpu.dec.r_rs2_pc ;
 wire \cpu.dec.r_set_cc ;
 wire \cpu.dec.r_store ;
 wire \cpu.dec.r_swapsp ;
 wire \cpu.dec.r_sys_call ;
 wire \cpu.dec.r_trap ;
 wire \cpu.dec.supmode ;
 wire \cpu.dec.user_io ;
 wire \cpu.ex.c_div_running ;
 wire \cpu.ex.c_mult[0] ;
 wire \cpu.ex.c_mult[10] ;
 wire \cpu.ex.c_mult[11] ;
 wire \cpu.ex.c_mult[12] ;
 wire \cpu.ex.c_mult[13] ;
 wire \cpu.ex.c_mult[14] ;
 wire \cpu.ex.c_mult[15] ;
 wire \cpu.ex.c_mult[1] ;
 wire \cpu.ex.c_mult[2] ;
 wire \cpu.ex.c_mult[3] ;
 wire \cpu.ex.c_mult[4] ;
 wire \cpu.ex.c_mult[5] ;
 wire \cpu.ex.c_mult[6] ;
 wire \cpu.ex.c_mult[7] ;
 wire \cpu.ex.c_mult[8] ;
 wire \cpu.ex.c_mult[9] ;
 wire \cpu.ex.c_mult_off[0] ;
 wire \cpu.ex.c_mult_off[1] ;
 wire \cpu.ex.c_mult_off[2] ;
 wire \cpu.ex.c_mult_off[3] ;
 wire \cpu.ex.c_mult_running ;
 wire \cpu.ex.genblk3.c_supmode ;
 wire \cpu.ex.genblk3.r_mmu_d_proxy ;
 wire \cpu.ex.genblk3.r_mmu_enable ;
 wire \cpu.ex.genblk3.r_prev_supmode ;
 wire \cpu.ex.i_flush_all ;
 wire \cpu.ex.ifetch ;
 wire \cpu.ex.io_access ;
 wire \cpu.ex.mmu_read[12] ;
 wire \cpu.ex.mmu_read[13] ;
 wire \cpu.ex.mmu_read[14] ;
 wire \cpu.ex.mmu_read[15] ;
 wire \cpu.ex.mmu_read[1] ;
 wire \cpu.ex.mmu_read[2] ;
 wire \cpu.ex.mmu_read[3] ;
 wire \cpu.ex.mmu_reg_data[0] ;
 wire \cpu.ex.pc[10] ;
 wire \cpu.ex.pc[11] ;
 wire \cpu.ex.pc[12] ;
 wire \cpu.ex.pc[13] ;
 wire \cpu.ex.pc[14] ;
 wire \cpu.ex.pc[15] ;
 wire \cpu.ex.pc[1] ;
 wire \cpu.ex.pc[2] ;
 wire \cpu.ex.pc[3] ;
 wire \cpu.ex.pc[4] ;
 wire \cpu.ex.pc[5] ;
 wire \cpu.ex.pc[6] ;
 wire \cpu.ex.pc[7] ;
 wire \cpu.ex.pc[8] ;
 wire \cpu.ex.pc[9] ;
 wire \cpu.ex.r_10[0] ;
 wire \cpu.ex.r_10[10] ;
 wire \cpu.ex.r_10[11] ;
 wire \cpu.ex.r_10[12] ;
 wire \cpu.ex.r_10[13] ;
 wire \cpu.ex.r_10[14] ;
 wire \cpu.ex.r_10[15] ;
 wire \cpu.ex.r_10[1] ;
 wire \cpu.ex.r_10[2] ;
 wire \cpu.ex.r_10[3] ;
 wire \cpu.ex.r_10[4] ;
 wire \cpu.ex.r_10[5] ;
 wire \cpu.ex.r_10[6] ;
 wire \cpu.ex.r_10[7] ;
 wire \cpu.ex.r_10[8] ;
 wire \cpu.ex.r_10[9] ;
 wire \cpu.ex.r_11[0] ;
 wire \cpu.ex.r_11[10] ;
 wire \cpu.ex.r_11[11] ;
 wire \cpu.ex.r_11[12] ;
 wire \cpu.ex.r_11[13] ;
 wire \cpu.ex.r_11[14] ;
 wire \cpu.ex.r_11[15] ;
 wire \cpu.ex.r_11[1] ;
 wire \cpu.ex.r_11[2] ;
 wire \cpu.ex.r_11[3] ;
 wire \cpu.ex.r_11[4] ;
 wire \cpu.ex.r_11[5] ;
 wire \cpu.ex.r_11[6] ;
 wire \cpu.ex.r_11[7] ;
 wire \cpu.ex.r_11[8] ;
 wire \cpu.ex.r_11[9] ;
 wire \cpu.ex.r_12[0] ;
 wire \cpu.ex.r_12[10] ;
 wire \cpu.ex.r_12[11] ;
 wire \cpu.ex.r_12[12] ;
 wire \cpu.ex.r_12[13] ;
 wire \cpu.ex.r_12[14] ;
 wire \cpu.ex.r_12[15] ;
 wire \cpu.ex.r_12[1] ;
 wire \cpu.ex.r_12[2] ;
 wire \cpu.ex.r_12[3] ;
 wire \cpu.ex.r_12[4] ;
 wire \cpu.ex.r_12[5] ;
 wire \cpu.ex.r_12[6] ;
 wire \cpu.ex.r_12[7] ;
 wire \cpu.ex.r_12[8] ;
 wire \cpu.ex.r_12[9] ;
 wire \cpu.ex.r_13[0] ;
 wire \cpu.ex.r_13[10] ;
 wire \cpu.ex.r_13[11] ;
 wire \cpu.ex.r_13[12] ;
 wire \cpu.ex.r_13[13] ;
 wire \cpu.ex.r_13[14] ;
 wire \cpu.ex.r_13[15] ;
 wire \cpu.ex.r_13[1] ;
 wire \cpu.ex.r_13[2] ;
 wire \cpu.ex.r_13[3] ;
 wire \cpu.ex.r_13[4] ;
 wire \cpu.ex.r_13[5] ;
 wire \cpu.ex.r_13[6] ;
 wire \cpu.ex.r_13[7] ;
 wire \cpu.ex.r_13[8] ;
 wire \cpu.ex.r_13[9] ;
 wire \cpu.ex.r_14[0] ;
 wire \cpu.ex.r_14[10] ;
 wire \cpu.ex.r_14[11] ;
 wire \cpu.ex.r_14[12] ;
 wire \cpu.ex.r_14[13] ;
 wire \cpu.ex.r_14[14] ;
 wire \cpu.ex.r_14[15] ;
 wire \cpu.ex.r_14[1] ;
 wire \cpu.ex.r_14[2] ;
 wire \cpu.ex.r_14[3] ;
 wire \cpu.ex.r_14[4] ;
 wire \cpu.ex.r_14[5] ;
 wire \cpu.ex.r_14[6] ;
 wire \cpu.ex.r_14[7] ;
 wire \cpu.ex.r_14[8] ;
 wire \cpu.ex.r_14[9] ;
 wire \cpu.ex.r_15[0] ;
 wire \cpu.ex.r_15[10] ;
 wire \cpu.ex.r_15[11] ;
 wire \cpu.ex.r_15[12] ;
 wire \cpu.ex.r_15[13] ;
 wire \cpu.ex.r_15[14] ;
 wire \cpu.ex.r_15[15] ;
 wire \cpu.ex.r_15[1] ;
 wire \cpu.ex.r_15[2] ;
 wire \cpu.ex.r_15[3] ;
 wire \cpu.ex.r_15[4] ;
 wire \cpu.ex.r_15[5] ;
 wire \cpu.ex.r_15[6] ;
 wire \cpu.ex.r_15[7] ;
 wire \cpu.ex.r_15[8] ;
 wire \cpu.ex.r_15[9] ;
 wire \cpu.ex.r_8[0] ;
 wire \cpu.ex.r_8[10] ;
 wire \cpu.ex.r_8[11] ;
 wire \cpu.ex.r_8[12] ;
 wire \cpu.ex.r_8[13] ;
 wire \cpu.ex.r_8[14] ;
 wire \cpu.ex.r_8[15] ;
 wire \cpu.ex.r_8[1] ;
 wire \cpu.ex.r_8[2] ;
 wire \cpu.ex.r_8[3] ;
 wire \cpu.ex.r_8[4] ;
 wire \cpu.ex.r_8[5] ;
 wire \cpu.ex.r_8[6] ;
 wire \cpu.ex.r_8[7] ;
 wire \cpu.ex.r_8[8] ;
 wire \cpu.ex.r_8[9] ;
 wire \cpu.ex.r_9[0] ;
 wire \cpu.ex.r_9[10] ;
 wire \cpu.ex.r_9[11] ;
 wire \cpu.ex.r_9[12] ;
 wire \cpu.ex.r_9[13] ;
 wire \cpu.ex.r_9[14] ;
 wire \cpu.ex.r_9[15] ;
 wire \cpu.ex.r_9[1] ;
 wire \cpu.ex.r_9[2] ;
 wire \cpu.ex.r_9[3] ;
 wire \cpu.ex.r_9[4] ;
 wire \cpu.ex.r_9[5] ;
 wire \cpu.ex.r_9[6] ;
 wire \cpu.ex.r_9[7] ;
 wire \cpu.ex.r_9[8] ;
 wire \cpu.ex.r_9[9] ;
 wire \cpu.ex.r_branch_stall ;
 wire \cpu.ex.r_cc ;
 wire \cpu.ex.r_div_running ;
 wire \cpu.ex.r_epc[10] ;
 wire \cpu.ex.r_epc[11] ;
 wire \cpu.ex.r_epc[12] ;
 wire \cpu.ex.r_epc[13] ;
 wire \cpu.ex.r_epc[14] ;
 wire \cpu.ex.r_epc[15] ;
 wire \cpu.ex.r_epc[1] ;
 wire \cpu.ex.r_epc[2] ;
 wire \cpu.ex.r_epc[3] ;
 wire \cpu.ex.r_epc[4] ;
 wire \cpu.ex.r_epc[5] ;
 wire \cpu.ex.r_epc[6] ;
 wire \cpu.ex.r_epc[7] ;
 wire \cpu.ex.r_epc[8] ;
 wire \cpu.ex.r_epc[9] ;
 wire \cpu.ex.r_ie ;
 wire \cpu.ex.r_lr[10] ;
 wire \cpu.ex.r_lr[11] ;
 wire \cpu.ex.r_lr[12] ;
 wire \cpu.ex.r_lr[13] ;
 wire \cpu.ex.r_lr[14] ;
 wire \cpu.ex.r_lr[15] ;
 wire \cpu.ex.r_lr[1] ;
 wire \cpu.ex.r_lr[2] ;
 wire \cpu.ex.r_lr[3] ;
 wire \cpu.ex.r_lr[4] ;
 wire \cpu.ex.r_lr[5] ;
 wire \cpu.ex.r_lr[6] ;
 wire \cpu.ex.r_lr[7] ;
 wire \cpu.ex.r_lr[8] ;
 wire \cpu.ex.r_lr[9] ;
 wire \cpu.ex.r_mult[0] ;
 wire \cpu.ex.r_mult[10] ;
 wire \cpu.ex.r_mult[11] ;
 wire \cpu.ex.r_mult[12] ;
 wire \cpu.ex.r_mult[13] ;
 wire \cpu.ex.r_mult[14] ;
 wire \cpu.ex.r_mult[15] ;
 wire \cpu.ex.r_mult[16] ;
 wire \cpu.ex.r_mult[17] ;
 wire \cpu.ex.r_mult[18] ;
 wire \cpu.ex.r_mult[19] ;
 wire \cpu.ex.r_mult[1] ;
 wire \cpu.ex.r_mult[20] ;
 wire \cpu.ex.r_mult[21] ;
 wire \cpu.ex.r_mult[22] ;
 wire \cpu.ex.r_mult[23] ;
 wire \cpu.ex.r_mult[24] ;
 wire \cpu.ex.r_mult[25] ;
 wire \cpu.ex.r_mult[26] ;
 wire \cpu.ex.r_mult[27] ;
 wire \cpu.ex.r_mult[28] ;
 wire \cpu.ex.r_mult[29] ;
 wire \cpu.ex.r_mult[2] ;
 wire \cpu.ex.r_mult[30] ;
 wire \cpu.ex.r_mult[31] ;
 wire \cpu.ex.r_mult[3] ;
 wire \cpu.ex.r_mult[4] ;
 wire \cpu.ex.r_mult[5] ;
 wire \cpu.ex.r_mult[6] ;
 wire \cpu.ex.r_mult[7] ;
 wire \cpu.ex.r_mult[8] ;
 wire \cpu.ex.r_mult[9] ;
 wire \cpu.ex.r_mult_off[0] ;
 wire \cpu.ex.r_mult_off[1] ;
 wire \cpu.ex.r_mult_off[2] ;
 wire \cpu.ex.r_mult_off[3] ;
 wire \cpu.ex.r_mult_running ;
 wire \cpu.ex.r_prev_ie ;
 wire \cpu.ex.r_read_stall ;
 wire \cpu.ex.r_set_cc ;
 wire \cpu.ex.r_sp[10] ;
 wire \cpu.ex.r_sp[11] ;
 wire \cpu.ex.r_sp[12] ;
 wire \cpu.ex.r_sp[13] ;
 wire \cpu.ex.r_sp[14] ;
 wire \cpu.ex.r_sp[15] ;
 wire \cpu.ex.r_sp[1] ;
 wire \cpu.ex.r_sp[2] ;
 wire \cpu.ex.r_sp[3] ;
 wire \cpu.ex.r_sp[4] ;
 wire \cpu.ex.r_sp[5] ;
 wire \cpu.ex.r_sp[6] ;
 wire \cpu.ex.r_sp[7] ;
 wire \cpu.ex.r_sp[8] ;
 wire \cpu.ex.r_sp[9] ;
 wire \cpu.ex.r_stmp[0] ;
 wire \cpu.ex.r_stmp[10] ;
 wire \cpu.ex.r_stmp[11] ;
 wire \cpu.ex.r_stmp[12] ;
 wire \cpu.ex.r_stmp[13] ;
 wire \cpu.ex.r_stmp[14] ;
 wire \cpu.ex.r_stmp[15] ;
 wire \cpu.ex.r_stmp[1] ;
 wire \cpu.ex.r_stmp[2] ;
 wire \cpu.ex.r_stmp[3] ;
 wire \cpu.ex.r_stmp[4] ;
 wire \cpu.ex.r_stmp[5] ;
 wire \cpu.ex.r_stmp[6] ;
 wire \cpu.ex.r_stmp[7] ;
 wire \cpu.ex.r_stmp[8] ;
 wire \cpu.ex.r_stmp[9] ;
 wire \cpu.ex.r_wb_addr[0] ;
 wire \cpu.ex.r_wb_addr[1] ;
 wire \cpu.ex.r_wb_addr[2] ;
 wire \cpu.ex.r_wb_addr[3] ;
 wire \cpu.ex.r_wb_swapsp ;
 wire \cpu.ex.r_wb_valid ;
 wire \cpu.ex.r_wmask[0] ;
 wire \cpu.ex.r_wmask[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[0] ;
 wire \cpu.genblk1.mmu.r_valid_d[10] ;
 wire \cpu.genblk1.mmu.r_valid_d[11] ;
 wire \cpu.genblk1.mmu.r_valid_d[12] ;
 wire \cpu.genblk1.mmu.r_valid_d[13] ;
 wire \cpu.genblk1.mmu.r_valid_d[14] ;
 wire \cpu.genblk1.mmu.r_valid_d[15] ;
 wire \cpu.genblk1.mmu.r_valid_d[16] ;
 wire \cpu.genblk1.mmu.r_valid_d[17] ;
 wire \cpu.genblk1.mmu.r_valid_d[18] ;
 wire \cpu.genblk1.mmu.r_valid_d[19] ;
 wire \cpu.genblk1.mmu.r_valid_d[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[20] ;
 wire \cpu.genblk1.mmu.r_valid_d[21] ;
 wire \cpu.genblk1.mmu.r_valid_d[22] ;
 wire \cpu.genblk1.mmu.r_valid_d[23] ;
 wire \cpu.genblk1.mmu.r_valid_d[24] ;
 wire \cpu.genblk1.mmu.r_valid_d[25] ;
 wire \cpu.genblk1.mmu.r_valid_d[26] ;
 wire \cpu.genblk1.mmu.r_valid_d[27] ;
 wire \cpu.genblk1.mmu.r_valid_d[28] ;
 wire \cpu.genblk1.mmu.r_valid_d[29] ;
 wire \cpu.genblk1.mmu.r_valid_d[2] ;
 wire \cpu.genblk1.mmu.r_valid_d[30] ;
 wire \cpu.genblk1.mmu.r_valid_d[31] ;
 wire \cpu.genblk1.mmu.r_valid_d[3] ;
 wire \cpu.genblk1.mmu.r_valid_d[4] ;
 wire \cpu.genblk1.mmu.r_valid_d[5] ;
 wire \cpu.genblk1.mmu.r_valid_d[6] ;
 wire \cpu.genblk1.mmu.r_valid_d[7] ;
 wire \cpu.genblk1.mmu.r_valid_d[8] ;
 wire \cpu.genblk1.mmu.r_valid_d[9] ;
 wire \cpu.genblk1.mmu.r_valid_i[0] ;
 wire \cpu.genblk1.mmu.r_valid_i[10] ;
 wire \cpu.genblk1.mmu.r_valid_i[11] ;
 wire \cpu.genblk1.mmu.r_valid_i[12] ;
 wire \cpu.genblk1.mmu.r_valid_i[13] ;
 wire \cpu.genblk1.mmu.r_valid_i[14] ;
 wire \cpu.genblk1.mmu.r_valid_i[15] ;
 wire \cpu.genblk1.mmu.r_valid_i[16] ;
 wire \cpu.genblk1.mmu.r_valid_i[17] ;
 wire \cpu.genblk1.mmu.r_valid_i[18] ;
 wire \cpu.genblk1.mmu.r_valid_i[19] ;
 wire \cpu.genblk1.mmu.r_valid_i[1] ;
 wire \cpu.genblk1.mmu.r_valid_i[20] ;
 wire \cpu.genblk1.mmu.r_valid_i[21] ;
 wire \cpu.genblk1.mmu.r_valid_i[22] ;
 wire \cpu.genblk1.mmu.r_valid_i[23] ;
 wire \cpu.genblk1.mmu.r_valid_i[24] ;
 wire \cpu.genblk1.mmu.r_valid_i[25] ;
 wire \cpu.genblk1.mmu.r_valid_i[26] ;
 wire \cpu.genblk1.mmu.r_valid_i[27] ;
 wire \cpu.genblk1.mmu.r_valid_i[28] ;
 wire \cpu.genblk1.mmu.r_valid_i[29] ;
 wire \cpu.genblk1.mmu.r_valid_i[2] ;
 wire \cpu.genblk1.mmu.r_valid_i[30] ;
 wire \cpu.genblk1.mmu.r_valid_i[31] ;
 wire \cpu.genblk1.mmu.r_valid_i[3] ;
 wire \cpu.genblk1.mmu.r_valid_i[4] ;
 wire \cpu.genblk1.mmu.r_valid_i[5] ;
 wire \cpu.genblk1.mmu.r_valid_i[6] ;
 wire \cpu.genblk1.mmu.r_valid_i[7] ;
 wire \cpu.genblk1.mmu.r_valid_i[8] ;
 wire \cpu.genblk1.mmu.r_valid_i[9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][9] ;
 wire \cpu.genblk1.mmu.r_writeable_d[0] ;
 wire \cpu.genblk1.mmu.r_writeable_d[10] ;
 wire \cpu.genblk1.mmu.r_writeable_d[11] ;
 wire \cpu.genblk1.mmu.r_writeable_d[12] ;
 wire \cpu.genblk1.mmu.r_writeable_d[13] ;
 wire \cpu.genblk1.mmu.r_writeable_d[14] ;
 wire \cpu.genblk1.mmu.r_writeable_d[15] ;
 wire \cpu.genblk1.mmu.r_writeable_d[16] ;
 wire \cpu.genblk1.mmu.r_writeable_d[17] ;
 wire \cpu.genblk1.mmu.r_writeable_d[18] ;
 wire \cpu.genblk1.mmu.r_writeable_d[19] ;
 wire \cpu.genblk1.mmu.r_writeable_d[1] ;
 wire \cpu.genblk1.mmu.r_writeable_d[20] ;
 wire \cpu.genblk1.mmu.r_writeable_d[21] ;
 wire \cpu.genblk1.mmu.r_writeable_d[22] ;
 wire \cpu.genblk1.mmu.r_writeable_d[23] ;
 wire \cpu.genblk1.mmu.r_writeable_d[24] ;
 wire \cpu.genblk1.mmu.r_writeable_d[25] ;
 wire \cpu.genblk1.mmu.r_writeable_d[26] ;
 wire \cpu.genblk1.mmu.r_writeable_d[27] ;
 wire \cpu.genblk1.mmu.r_writeable_d[28] ;
 wire \cpu.genblk1.mmu.r_writeable_d[29] ;
 wire \cpu.genblk1.mmu.r_writeable_d[2] ;
 wire \cpu.genblk1.mmu.r_writeable_d[30] ;
 wire \cpu.genblk1.mmu.r_writeable_d[31] ;
 wire \cpu.genblk1.mmu.r_writeable_d[3] ;
 wire \cpu.genblk1.mmu.r_writeable_d[4] ;
 wire \cpu.genblk1.mmu.r_writeable_d[5] ;
 wire \cpu.genblk1.mmu.r_writeable_d[6] ;
 wire \cpu.genblk1.mmu.r_writeable_d[7] ;
 wire \cpu.genblk1.mmu.r_writeable_d[8] ;
 wire \cpu.genblk1.mmu.r_writeable_d[9] ;
 wire \cpu.gpio.genblk1[3].srcs_o[0] ;
 wire \cpu.gpio.genblk1[3].srcs_o[11] ;
 wire \cpu.gpio.genblk1[3].srcs_o[1] ;
 wire \cpu.gpio.genblk1[3].srcs_o[2] ;
 wire \cpu.gpio.genblk1[3].srcs_o[3] ;
 wire \cpu.gpio.genblk1[3].srcs_o[4] ;
 wire \cpu.gpio.genblk1[3].srcs_o[5] ;
 wire \cpu.gpio.genblk1[3].srcs_o[6] ;
 wire \cpu.gpio.genblk1[3].srcs_o[7] ;
 wire \cpu.gpio.genblk1[3].srcs_o[8] ;
 wire \cpu.gpio.genblk1[4].srcs_o[0] ;
 wire \cpu.gpio.genblk1[5].srcs_o[0] ;
 wire \cpu.gpio.genblk1[6].srcs_o[0] ;
 wire \cpu.gpio.genblk1[7].srcs_o[0] ;
 wire \cpu.gpio.genblk2[4].srcs_io[0] ;
 wire \cpu.gpio.genblk2[5].srcs_io[0] ;
 wire \cpu.gpio.genblk2[6].srcs_io[0] ;
 wire \cpu.gpio.genblk2[7].srcs_io[0] ;
 wire \cpu.gpio.r_enable_in[0] ;
 wire \cpu.gpio.r_enable_in[1] ;
 wire \cpu.gpio.r_enable_in[2] ;
 wire \cpu.gpio.r_enable_in[3] ;
 wire \cpu.gpio.r_enable_in[4] ;
 wire \cpu.gpio.r_enable_in[5] ;
 wire \cpu.gpio.r_enable_in[6] ;
 wire \cpu.gpio.r_enable_in[7] ;
 wire \cpu.gpio.r_enable_io[4] ;
 wire \cpu.gpio.r_enable_io[5] ;
 wire \cpu.gpio.r_enable_io[6] ;
 wire \cpu.gpio.r_enable_io[7] ;
 wire \cpu.gpio.r_spi_miso_src[0][0] ;
 wire \cpu.gpio.r_spi_miso_src[0][1] ;
 wire \cpu.gpio.r_spi_miso_src[0][2] ;
 wire \cpu.gpio.r_spi_miso_src[0][3] ;
 wire \cpu.gpio.r_spi_miso_src[1][0] ;
 wire \cpu.gpio.r_spi_miso_src[1][1] ;
 wire \cpu.gpio.r_spi_miso_src[1][2] ;
 wire \cpu.gpio.r_spi_miso_src[1][3] ;
 wire \cpu.gpio.r_src_io[4][0] ;
 wire \cpu.gpio.r_src_io[4][1] ;
 wire \cpu.gpio.r_src_io[4][2] ;
 wire \cpu.gpio.r_src_io[4][3] ;
 wire \cpu.gpio.r_src_io[5][0] ;
 wire \cpu.gpio.r_src_io[5][1] ;
 wire \cpu.gpio.r_src_io[5][2] ;
 wire \cpu.gpio.r_src_io[5][3] ;
 wire \cpu.gpio.r_src_io[6][0] ;
 wire \cpu.gpio.r_src_io[6][1] ;
 wire \cpu.gpio.r_src_io[6][2] ;
 wire \cpu.gpio.r_src_io[6][3] ;
 wire \cpu.gpio.r_src_io[7][0] ;
 wire \cpu.gpio.r_src_io[7][1] ;
 wire \cpu.gpio.r_src_io[7][2] ;
 wire \cpu.gpio.r_src_io[7][3] ;
 wire \cpu.gpio.r_src_o[3][0] ;
 wire \cpu.gpio.r_src_o[3][1] ;
 wire \cpu.gpio.r_src_o[3][2] ;
 wire \cpu.gpio.r_src_o[3][3] ;
 wire \cpu.gpio.r_src_o[4][0] ;
 wire \cpu.gpio.r_src_o[4][1] ;
 wire \cpu.gpio.r_src_o[4][2] ;
 wire \cpu.gpio.r_src_o[4][3] ;
 wire \cpu.gpio.r_src_o[5][0] ;
 wire \cpu.gpio.r_src_o[5][1] ;
 wire \cpu.gpio.r_src_o[5][2] ;
 wire \cpu.gpio.r_src_o[5][3] ;
 wire \cpu.gpio.r_src_o[6][0] ;
 wire \cpu.gpio.r_src_o[6][1] ;
 wire \cpu.gpio.r_src_o[6][2] ;
 wire \cpu.gpio.r_src_o[6][3] ;
 wire \cpu.gpio.r_src_o[7][0] ;
 wire \cpu.gpio.r_src_o[7][1] ;
 wire \cpu.gpio.r_src_o[7][2] ;
 wire \cpu.gpio.r_src_o[7][3] ;
 wire \cpu.gpio.r_uart_rx_src[0] ;
 wire \cpu.gpio.r_uart_rx_src[1] ;
 wire \cpu.gpio.r_uart_rx_src[2] ;
 wire \cpu.gpio.uart_rx ;
 wire \cpu.i_wstrobe_d ;
 wire \cpu.icache.r_data[0][0] ;
 wire \cpu.icache.r_data[0][10] ;
 wire \cpu.icache.r_data[0][11] ;
 wire \cpu.icache.r_data[0][12] ;
 wire \cpu.icache.r_data[0][13] ;
 wire \cpu.icache.r_data[0][14] ;
 wire \cpu.icache.r_data[0][15] ;
 wire \cpu.icache.r_data[0][16] ;
 wire \cpu.icache.r_data[0][17] ;
 wire \cpu.icache.r_data[0][18] ;
 wire \cpu.icache.r_data[0][19] ;
 wire \cpu.icache.r_data[0][1] ;
 wire \cpu.icache.r_data[0][20] ;
 wire \cpu.icache.r_data[0][21] ;
 wire \cpu.icache.r_data[0][22] ;
 wire \cpu.icache.r_data[0][23] ;
 wire \cpu.icache.r_data[0][24] ;
 wire \cpu.icache.r_data[0][25] ;
 wire \cpu.icache.r_data[0][26] ;
 wire \cpu.icache.r_data[0][27] ;
 wire \cpu.icache.r_data[0][28] ;
 wire \cpu.icache.r_data[0][29] ;
 wire \cpu.icache.r_data[0][2] ;
 wire \cpu.icache.r_data[0][30] ;
 wire \cpu.icache.r_data[0][31] ;
 wire \cpu.icache.r_data[0][3] ;
 wire \cpu.icache.r_data[0][4] ;
 wire \cpu.icache.r_data[0][5] ;
 wire \cpu.icache.r_data[0][6] ;
 wire \cpu.icache.r_data[0][7] ;
 wire \cpu.icache.r_data[0][8] ;
 wire \cpu.icache.r_data[0][9] ;
 wire \cpu.icache.r_data[1][0] ;
 wire \cpu.icache.r_data[1][10] ;
 wire \cpu.icache.r_data[1][11] ;
 wire \cpu.icache.r_data[1][12] ;
 wire \cpu.icache.r_data[1][13] ;
 wire \cpu.icache.r_data[1][14] ;
 wire \cpu.icache.r_data[1][15] ;
 wire \cpu.icache.r_data[1][16] ;
 wire \cpu.icache.r_data[1][17] ;
 wire \cpu.icache.r_data[1][18] ;
 wire \cpu.icache.r_data[1][19] ;
 wire \cpu.icache.r_data[1][1] ;
 wire \cpu.icache.r_data[1][20] ;
 wire \cpu.icache.r_data[1][21] ;
 wire \cpu.icache.r_data[1][22] ;
 wire \cpu.icache.r_data[1][23] ;
 wire \cpu.icache.r_data[1][24] ;
 wire \cpu.icache.r_data[1][25] ;
 wire \cpu.icache.r_data[1][26] ;
 wire \cpu.icache.r_data[1][27] ;
 wire \cpu.icache.r_data[1][28] ;
 wire \cpu.icache.r_data[1][29] ;
 wire \cpu.icache.r_data[1][2] ;
 wire \cpu.icache.r_data[1][30] ;
 wire \cpu.icache.r_data[1][31] ;
 wire \cpu.icache.r_data[1][3] ;
 wire \cpu.icache.r_data[1][4] ;
 wire \cpu.icache.r_data[1][5] ;
 wire \cpu.icache.r_data[1][6] ;
 wire \cpu.icache.r_data[1][7] ;
 wire \cpu.icache.r_data[1][8] ;
 wire \cpu.icache.r_data[1][9] ;
 wire \cpu.icache.r_data[2][0] ;
 wire \cpu.icache.r_data[2][10] ;
 wire \cpu.icache.r_data[2][11] ;
 wire \cpu.icache.r_data[2][12] ;
 wire \cpu.icache.r_data[2][13] ;
 wire \cpu.icache.r_data[2][14] ;
 wire \cpu.icache.r_data[2][15] ;
 wire \cpu.icache.r_data[2][16] ;
 wire \cpu.icache.r_data[2][17] ;
 wire \cpu.icache.r_data[2][18] ;
 wire \cpu.icache.r_data[2][19] ;
 wire \cpu.icache.r_data[2][1] ;
 wire \cpu.icache.r_data[2][20] ;
 wire \cpu.icache.r_data[2][21] ;
 wire \cpu.icache.r_data[2][22] ;
 wire \cpu.icache.r_data[2][23] ;
 wire \cpu.icache.r_data[2][24] ;
 wire \cpu.icache.r_data[2][25] ;
 wire \cpu.icache.r_data[2][26] ;
 wire \cpu.icache.r_data[2][27] ;
 wire \cpu.icache.r_data[2][28] ;
 wire \cpu.icache.r_data[2][29] ;
 wire \cpu.icache.r_data[2][2] ;
 wire \cpu.icache.r_data[2][30] ;
 wire \cpu.icache.r_data[2][31] ;
 wire \cpu.icache.r_data[2][3] ;
 wire \cpu.icache.r_data[2][4] ;
 wire \cpu.icache.r_data[2][5] ;
 wire \cpu.icache.r_data[2][6] ;
 wire \cpu.icache.r_data[2][7] ;
 wire \cpu.icache.r_data[2][8] ;
 wire \cpu.icache.r_data[2][9] ;
 wire \cpu.icache.r_data[3][0] ;
 wire \cpu.icache.r_data[3][10] ;
 wire \cpu.icache.r_data[3][11] ;
 wire \cpu.icache.r_data[3][12] ;
 wire \cpu.icache.r_data[3][13] ;
 wire \cpu.icache.r_data[3][14] ;
 wire \cpu.icache.r_data[3][15] ;
 wire \cpu.icache.r_data[3][16] ;
 wire \cpu.icache.r_data[3][17] ;
 wire \cpu.icache.r_data[3][18] ;
 wire \cpu.icache.r_data[3][19] ;
 wire \cpu.icache.r_data[3][1] ;
 wire \cpu.icache.r_data[3][20] ;
 wire \cpu.icache.r_data[3][21] ;
 wire \cpu.icache.r_data[3][22] ;
 wire \cpu.icache.r_data[3][23] ;
 wire \cpu.icache.r_data[3][24] ;
 wire \cpu.icache.r_data[3][25] ;
 wire \cpu.icache.r_data[3][26] ;
 wire \cpu.icache.r_data[3][27] ;
 wire \cpu.icache.r_data[3][28] ;
 wire \cpu.icache.r_data[3][29] ;
 wire \cpu.icache.r_data[3][2] ;
 wire \cpu.icache.r_data[3][30] ;
 wire \cpu.icache.r_data[3][31] ;
 wire \cpu.icache.r_data[3][3] ;
 wire \cpu.icache.r_data[3][4] ;
 wire \cpu.icache.r_data[3][5] ;
 wire \cpu.icache.r_data[3][6] ;
 wire \cpu.icache.r_data[3][7] ;
 wire \cpu.icache.r_data[3][8] ;
 wire \cpu.icache.r_data[3][9] ;
 wire \cpu.icache.r_data[4][0] ;
 wire \cpu.icache.r_data[4][10] ;
 wire \cpu.icache.r_data[4][11] ;
 wire \cpu.icache.r_data[4][12] ;
 wire \cpu.icache.r_data[4][13] ;
 wire \cpu.icache.r_data[4][14] ;
 wire \cpu.icache.r_data[4][15] ;
 wire \cpu.icache.r_data[4][16] ;
 wire \cpu.icache.r_data[4][17] ;
 wire \cpu.icache.r_data[4][18] ;
 wire \cpu.icache.r_data[4][19] ;
 wire \cpu.icache.r_data[4][1] ;
 wire \cpu.icache.r_data[4][20] ;
 wire \cpu.icache.r_data[4][21] ;
 wire \cpu.icache.r_data[4][22] ;
 wire \cpu.icache.r_data[4][23] ;
 wire \cpu.icache.r_data[4][24] ;
 wire \cpu.icache.r_data[4][25] ;
 wire \cpu.icache.r_data[4][26] ;
 wire \cpu.icache.r_data[4][27] ;
 wire \cpu.icache.r_data[4][28] ;
 wire \cpu.icache.r_data[4][29] ;
 wire \cpu.icache.r_data[4][2] ;
 wire \cpu.icache.r_data[4][30] ;
 wire \cpu.icache.r_data[4][31] ;
 wire \cpu.icache.r_data[4][3] ;
 wire \cpu.icache.r_data[4][4] ;
 wire \cpu.icache.r_data[4][5] ;
 wire \cpu.icache.r_data[4][6] ;
 wire \cpu.icache.r_data[4][7] ;
 wire \cpu.icache.r_data[4][8] ;
 wire \cpu.icache.r_data[4][9] ;
 wire \cpu.icache.r_data[5][0] ;
 wire \cpu.icache.r_data[5][10] ;
 wire \cpu.icache.r_data[5][11] ;
 wire \cpu.icache.r_data[5][12] ;
 wire \cpu.icache.r_data[5][13] ;
 wire \cpu.icache.r_data[5][14] ;
 wire \cpu.icache.r_data[5][15] ;
 wire \cpu.icache.r_data[5][16] ;
 wire \cpu.icache.r_data[5][17] ;
 wire \cpu.icache.r_data[5][18] ;
 wire \cpu.icache.r_data[5][19] ;
 wire \cpu.icache.r_data[5][1] ;
 wire \cpu.icache.r_data[5][20] ;
 wire \cpu.icache.r_data[5][21] ;
 wire \cpu.icache.r_data[5][22] ;
 wire \cpu.icache.r_data[5][23] ;
 wire \cpu.icache.r_data[5][24] ;
 wire \cpu.icache.r_data[5][25] ;
 wire \cpu.icache.r_data[5][26] ;
 wire \cpu.icache.r_data[5][27] ;
 wire \cpu.icache.r_data[5][28] ;
 wire \cpu.icache.r_data[5][29] ;
 wire \cpu.icache.r_data[5][2] ;
 wire \cpu.icache.r_data[5][30] ;
 wire \cpu.icache.r_data[5][31] ;
 wire \cpu.icache.r_data[5][3] ;
 wire \cpu.icache.r_data[5][4] ;
 wire \cpu.icache.r_data[5][5] ;
 wire \cpu.icache.r_data[5][6] ;
 wire \cpu.icache.r_data[5][7] ;
 wire \cpu.icache.r_data[5][8] ;
 wire \cpu.icache.r_data[5][9] ;
 wire \cpu.icache.r_data[6][0] ;
 wire \cpu.icache.r_data[6][10] ;
 wire \cpu.icache.r_data[6][11] ;
 wire \cpu.icache.r_data[6][12] ;
 wire \cpu.icache.r_data[6][13] ;
 wire \cpu.icache.r_data[6][14] ;
 wire \cpu.icache.r_data[6][15] ;
 wire \cpu.icache.r_data[6][16] ;
 wire \cpu.icache.r_data[6][17] ;
 wire \cpu.icache.r_data[6][18] ;
 wire \cpu.icache.r_data[6][19] ;
 wire \cpu.icache.r_data[6][1] ;
 wire \cpu.icache.r_data[6][20] ;
 wire \cpu.icache.r_data[6][21] ;
 wire \cpu.icache.r_data[6][22] ;
 wire \cpu.icache.r_data[6][23] ;
 wire \cpu.icache.r_data[6][24] ;
 wire \cpu.icache.r_data[6][25] ;
 wire \cpu.icache.r_data[6][26] ;
 wire \cpu.icache.r_data[6][27] ;
 wire \cpu.icache.r_data[6][28] ;
 wire \cpu.icache.r_data[6][29] ;
 wire \cpu.icache.r_data[6][2] ;
 wire \cpu.icache.r_data[6][30] ;
 wire \cpu.icache.r_data[6][31] ;
 wire \cpu.icache.r_data[6][3] ;
 wire \cpu.icache.r_data[6][4] ;
 wire \cpu.icache.r_data[6][5] ;
 wire \cpu.icache.r_data[6][6] ;
 wire \cpu.icache.r_data[6][7] ;
 wire \cpu.icache.r_data[6][8] ;
 wire \cpu.icache.r_data[6][9] ;
 wire \cpu.icache.r_data[7][0] ;
 wire \cpu.icache.r_data[7][10] ;
 wire \cpu.icache.r_data[7][11] ;
 wire \cpu.icache.r_data[7][12] ;
 wire \cpu.icache.r_data[7][13] ;
 wire \cpu.icache.r_data[7][14] ;
 wire \cpu.icache.r_data[7][15] ;
 wire \cpu.icache.r_data[7][16] ;
 wire \cpu.icache.r_data[7][17] ;
 wire \cpu.icache.r_data[7][18] ;
 wire \cpu.icache.r_data[7][19] ;
 wire \cpu.icache.r_data[7][1] ;
 wire \cpu.icache.r_data[7][20] ;
 wire \cpu.icache.r_data[7][21] ;
 wire \cpu.icache.r_data[7][22] ;
 wire \cpu.icache.r_data[7][23] ;
 wire \cpu.icache.r_data[7][24] ;
 wire \cpu.icache.r_data[7][25] ;
 wire \cpu.icache.r_data[7][26] ;
 wire \cpu.icache.r_data[7][27] ;
 wire \cpu.icache.r_data[7][28] ;
 wire \cpu.icache.r_data[7][29] ;
 wire \cpu.icache.r_data[7][2] ;
 wire \cpu.icache.r_data[7][30] ;
 wire \cpu.icache.r_data[7][31] ;
 wire \cpu.icache.r_data[7][3] ;
 wire \cpu.icache.r_data[7][4] ;
 wire \cpu.icache.r_data[7][5] ;
 wire \cpu.icache.r_data[7][6] ;
 wire \cpu.icache.r_data[7][7] ;
 wire \cpu.icache.r_data[7][8] ;
 wire \cpu.icache.r_data[7][9] ;
 wire \cpu.icache.r_offset[0] ;
 wire \cpu.icache.r_offset[1] ;
 wire \cpu.icache.r_offset[2] ;
 wire \cpu.icache.r_tag[0][10] ;
 wire \cpu.icache.r_tag[0][11] ;
 wire \cpu.icache.r_tag[0][12] ;
 wire \cpu.icache.r_tag[0][13] ;
 wire \cpu.icache.r_tag[0][14] ;
 wire \cpu.icache.r_tag[0][15] ;
 wire \cpu.icache.r_tag[0][16] ;
 wire \cpu.icache.r_tag[0][17] ;
 wire \cpu.icache.r_tag[0][18] ;
 wire \cpu.icache.r_tag[0][19] ;
 wire \cpu.icache.r_tag[0][20] ;
 wire \cpu.icache.r_tag[0][21] ;
 wire \cpu.icache.r_tag[0][22] ;
 wire \cpu.icache.r_tag[0][23] ;
 wire \cpu.icache.r_tag[0][5] ;
 wire \cpu.icache.r_tag[0][6] ;
 wire \cpu.icache.r_tag[0][7] ;
 wire \cpu.icache.r_tag[0][8] ;
 wire \cpu.icache.r_tag[0][9] ;
 wire \cpu.icache.r_tag[1][10] ;
 wire \cpu.icache.r_tag[1][11] ;
 wire \cpu.icache.r_tag[1][12] ;
 wire \cpu.icache.r_tag[1][13] ;
 wire \cpu.icache.r_tag[1][14] ;
 wire \cpu.icache.r_tag[1][15] ;
 wire \cpu.icache.r_tag[1][16] ;
 wire \cpu.icache.r_tag[1][17] ;
 wire \cpu.icache.r_tag[1][18] ;
 wire \cpu.icache.r_tag[1][19] ;
 wire \cpu.icache.r_tag[1][20] ;
 wire \cpu.icache.r_tag[1][21] ;
 wire \cpu.icache.r_tag[1][22] ;
 wire \cpu.icache.r_tag[1][23] ;
 wire \cpu.icache.r_tag[1][5] ;
 wire \cpu.icache.r_tag[1][6] ;
 wire \cpu.icache.r_tag[1][7] ;
 wire \cpu.icache.r_tag[1][8] ;
 wire \cpu.icache.r_tag[1][9] ;
 wire \cpu.icache.r_tag[2][10] ;
 wire \cpu.icache.r_tag[2][11] ;
 wire \cpu.icache.r_tag[2][12] ;
 wire \cpu.icache.r_tag[2][13] ;
 wire \cpu.icache.r_tag[2][14] ;
 wire \cpu.icache.r_tag[2][15] ;
 wire \cpu.icache.r_tag[2][16] ;
 wire \cpu.icache.r_tag[2][17] ;
 wire \cpu.icache.r_tag[2][18] ;
 wire \cpu.icache.r_tag[2][19] ;
 wire \cpu.icache.r_tag[2][20] ;
 wire \cpu.icache.r_tag[2][21] ;
 wire \cpu.icache.r_tag[2][22] ;
 wire \cpu.icache.r_tag[2][23] ;
 wire \cpu.icache.r_tag[2][5] ;
 wire \cpu.icache.r_tag[2][6] ;
 wire \cpu.icache.r_tag[2][7] ;
 wire \cpu.icache.r_tag[2][8] ;
 wire \cpu.icache.r_tag[2][9] ;
 wire \cpu.icache.r_tag[3][10] ;
 wire \cpu.icache.r_tag[3][11] ;
 wire \cpu.icache.r_tag[3][12] ;
 wire \cpu.icache.r_tag[3][13] ;
 wire \cpu.icache.r_tag[3][14] ;
 wire \cpu.icache.r_tag[3][15] ;
 wire \cpu.icache.r_tag[3][16] ;
 wire \cpu.icache.r_tag[3][17] ;
 wire \cpu.icache.r_tag[3][18] ;
 wire \cpu.icache.r_tag[3][19] ;
 wire \cpu.icache.r_tag[3][20] ;
 wire \cpu.icache.r_tag[3][21] ;
 wire \cpu.icache.r_tag[3][22] ;
 wire \cpu.icache.r_tag[3][23] ;
 wire \cpu.icache.r_tag[3][5] ;
 wire \cpu.icache.r_tag[3][6] ;
 wire \cpu.icache.r_tag[3][7] ;
 wire \cpu.icache.r_tag[3][8] ;
 wire \cpu.icache.r_tag[3][9] ;
 wire \cpu.icache.r_tag[4][10] ;
 wire \cpu.icache.r_tag[4][11] ;
 wire \cpu.icache.r_tag[4][12] ;
 wire \cpu.icache.r_tag[4][13] ;
 wire \cpu.icache.r_tag[4][14] ;
 wire \cpu.icache.r_tag[4][15] ;
 wire \cpu.icache.r_tag[4][16] ;
 wire \cpu.icache.r_tag[4][17] ;
 wire \cpu.icache.r_tag[4][18] ;
 wire \cpu.icache.r_tag[4][19] ;
 wire \cpu.icache.r_tag[4][20] ;
 wire \cpu.icache.r_tag[4][21] ;
 wire \cpu.icache.r_tag[4][22] ;
 wire \cpu.icache.r_tag[4][23] ;
 wire \cpu.icache.r_tag[4][5] ;
 wire \cpu.icache.r_tag[4][6] ;
 wire \cpu.icache.r_tag[4][7] ;
 wire \cpu.icache.r_tag[4][8] ;
 wire \cpu.icache.r_tag[4][9] ;
 wire \cpu.icache.r_tag[5][10] ;
 wire \cpu.icache.r_tag[5][11] ;
 wire \cpu.icache.r_tag[5][12] ;
 wire \cpu.icache.r_tag[5][13] ;
 wire \cpu.icache.r_tag[5][14] ;
 wire \cpu.icache.r_tag[5][15] ;
 wire \cpu.icache.r_tag[5][16] ;
 wire \cpu.icache.r_tag[5][17] ;
 wire \cpu.icache.r_tag[5][18] ;
 wire \cpu.icache.r_tag[5][19] ;
 wire \cpu.icache.r_tag[5][20] ;
 wire \cpu.icache.r_tag[5][21] ;
 wire \cpu.icache.r_tag[5][22] ;
 wire \cpu.icache.r_tag[5][23] ;
 wire \cpu.icache.r_tag[5][5] ;
 wire \cpu.icache.r_tag[5][6] ;
 wire \cpu.icache.r_tag[5][7] ;
 wire \cpu.icache.r_tag[5][8] ;
 wire \cpu.icache.r_tag[5][9] ;
 wire \cpu.icache.r_tag[6][10] ;
 wire \cpu.icache.r_tag[6][11] ;
 wire \cpu.icache.r_tag[6][12] ;
 wire \cpu.icache.r_tag[6][13] ;
 wire \cpu.icache.r_tag[6][14] ;
 wire \cpu.icache.r_tag[6][15] ;
 wire \cpu.icache.r_tag[6][16] ;
 wire \cpu.icache.r_tag[6][17] ;
 wire \cpu.icache.r_tag[6][18] ;
 wire \cpu.icache.r_tag[6][19] ;
 wire \cpu.icache.r_tag[6][20] ;
 wire \cpu.icache.r_tag[6][21] ;
 wire \cpu.icache.r_tag[6][22] ;
 wire \cpu.icache.r_tag[6][23] ;
 wire \cpu.icache.r_tag[6][5] ;
 wire \cpu.icache.r_tag[6][6] ;
 wire \cpu.icache.r_tag[6][7] ;
 wire \cpu.icache.r_tag[6][8] ;
 wire \cpu.icache.r_tag[6][9] ;
 wire \cpu.icache.r_tag[7][10] ;
 wire \cpu.icache.r_tag[7][11] ;
 wire \cpu.icache.r_tag[7][12] ;
 wire \cpu.icache.r_tag[7][13] ;
 wire \cpu.icache.r_tag[7][14] ;
 wire \cpu.icache.r_tag[7][15] ;
 wire \cpu.icache.r_tag[7][16] ;
 wire \cpu.icache.r_tag[7][17] ;
 wire \cpu.icache.r_tag[7][18] ;
 wire \cpu.icache.r_tag[7][19] ;
 wire \cpu.icache.r_tag[7][20] ;
 wire \cpu.icache.r_tag[7][21] ;
 wire \cpu.icache.r_tag[7][22] ;
 wire \cpu.icache.r_tag[7][23] ;
 wire \cpu.icache.r_tag[7][5] ;
 wire \cpu.icache.r_tag[7][6] ;
 wire \cpu.icache.r_tag[7][7] ;
 wire \cpu.icache.r_tag[7][8] ;
 wire \cpu.icache.r_tag[7][9] ;
 wire \cpu.icache.r_valid[0] ;
 wire \cpu.icache.r_valid[1] ;
 wire \cpu.icache.r_valid[2] ;
 wire \cpu.icache.r_valid[3] ;
 wire \cpu.icache.r_valid[4] ;
 wire \cpu.icache.r_valid[5] ;
 wire \cpu.icache.r_valid[6] ;
 wire \cpu.icache.r_valid[7] ;
 wire \cpu.intr.r_clock ;
 wire \cpu.intr.r_clock_cmp[0] ;
 wire \cpu.intr.r_clock_cmp[10] ;
 wire \cpu.intr.r_clock_cmp[11] ;
 wire \cpu.intr.r_clock_cmp[12] ;
 wire \cpu.intr.r_clock_cmp[13] ;
 wire \cpu.intr.r_clock_cmp[14] ;
 wire \cpu.intr.r_clock_cmp[15] ;
 wire \cpu.intr.r_clock_cmp[16] ;
 wire \cpu.intr.r_clock_cmp[17] ;
 wire \cpu.intr.r_clock_cmp[18] ;
 wire \cpu.intr.r_clock_cmp[19] ;
 wire \cpu.intr.r_clock_cmp[1] ;
 wire \cpu.intr.r_clock_cmp[20] ;
 wire \cpu.intr.r_clock_cmp[21] ;
 wire \cpu.intr.r_clock_cmp[22] ;
 wire \cpu.intr.r_clock_cmp[23] ;
 wire \cpu.intr.r_clock_cmp[24] ;
 wire \cpu.intr.r_clock_cmp[25] ;
 wire \cpu.intr.r_clock_cmp[26] ;
 wire \cpu.intr.r_clock_cmp[27] ;
 wire \cpu.intr.r_clock_cmp[28] ;
 wire \cpu.intr.r_clock_cmp[29] ;
 wire \cpu.intr.r_clock_cmp[2] ;
 wire \cpu.intr.r_clock_cmp[30] ;
 wire \cpu.intr.r_clock_cmp[31] ;
 wire \cpu.intr.r_clock_cmp[3] ;
 wire \cpu.intr.r_clock_cmp[4] ;
 wire \cpu.intr.r_clock_cmp[5] ;
 wire \cpu.intr.r_clock_cmp[6] ;
 wire \cpu.intr.r_clock_cmp[7] ;
 wire \cpu.intr.r_clock_cmp[8] ;
 wire \cpu.intr.r_clock_cmp[9] ;
 wire \cpu.intr.r_clock_count[0] ;
 wire \cpu.intr.r_clock_count[10] ;
 wire \cpu.intr.r_clock_count[11] ;
 wire \cpu.intr.r_clock_count[12] ;
 wire \cpu.intr.r_clock_count[13] ;
 wire \cpu.intr.r_clock_count[14] ;
 wire \cpu.intr.r_clock_count[15] ;
 wire \cpu.intr.r_clock_count[16] ;
 wire \cpu.intr.r_clock_count[17] ;
 wire \cpu.intr.r_clock_count[18] ;
 wire \cpu.intr.r_clock_count[19] ;
 wire \cpu.intr.r_clock_count[1] ;
 wire \cpu.intr.r_clock_count[20] ;
 wire \cpu.intr.r_clock_count[21] ;
 wire \cpu.intr.r_clock_count[22] ;
 wire \cpu.intr.r_clock_count[23] ;
 wire \cpu.intr.r_clock_count[24] ;
 wire \cpu.intr.r_clock_count[25] ;
 wire \cpu.intr.r_clock_count[26] ;
 wire \cpu.intr.r_clock_count[27] ;
 wire \cpu.intr.r_clock_count[28] ;
 wire \cpu.intr.r_clock_count[29] ;
 wire \cpu.intr.r_clock_count[2] ;
 wire \cpu.intr.r_clock_count[30] ;
 wire \cpu.intr.r_clock_count[31] ;
 wire \cpu.intr.r_clock_count[3] ;
 wire \cpu.intr.r_clock_count[4] ;
 wire \cpu.intr.r_clock_count[5] ;
 wire \cpu.intr.r_clock_count[6] ;
 wire \cpu.intr.r_clock_count[7] ;
 wire \cpu.intr.r_clock_count[8] ;
 wire \cpu.intr.r_clock_count[9] ;
 wire \cpu.intr.r_enable[0] ;
 wire \cpu.intr.r_enable[1] ;
 wire \cpu.intr.r_enable[2] ;
 wire \cpu.intr.r_enable[3] ;
 wire \cpu.intr.r_enable[4] ;
 wire \cpu.intr.r_enable[5] ;
 wire \cpu.intr.r_swi ;
 wire \cpu.intr.r_timer ;
 wire \cpu.intr.r_timer_count[0] ;
 wire \cpu.intr.r_timer_count[10] ;
 wire \cpu.intr.r_timer_count[11] ;
 wire \cpu.intr.r_timer_count[12] ;
 wire \cpu.intr.r_timer_count[13] ;
 wire \cpu.intr.r_timer_count[14] ;
 wire \cpu.intr.r_timer_count[15] ;
 wire \cpu.intr.r_timer_count[16] ;
 wire \cpu.intr.r_timer_count[17] ;
 wire \cpu.intr.r_timer_count[18] ;
 wire \cpu.intr.r_timer_count[19] ;
 wire \cpu.intr.r_timer_count[1] ;
 wire \cpu.intr.r_timer_count[20] ;
 wire \cpu.intr.r_timer_count[21] ;
 wire \cpu.intr.r_timer_count[22] ;
 wire \cpu.intr.r_timer_count[23] ;
 wire \cpu.intr.r_timer_count[2] ;
 wire \cpu.intr.r_timer_count[3] ;
 wire \cpu.intr.r_timer_count[4] ;
 wire \cpu.intr.r_timer_count[5] ;
 wire \cpu.intr.r_timer_count[6] ;
 wire \cpu.intr.r_timer_count[7] ;
 wire \cpu.intr.r_timer_count[8] ;
 wire \cpu.intr.r_timer_count[9] ;
 wire \cpu.intr.r_timer_reload[0] ;
 wire \cpu.intr.r_timer_reload[10] ;
 wire \cpu.intr.r_timer_reload[11] ;
 wire \cpu.intr.r_timer_reload[12] ;
 wire \cpu.intr.r_timer_reload[13] ;
 wire \cpu.intr.r_timer_reload[14] ;
 wire \cpu.intr.r_timer_reload[15] ;
 wire \cpu.intr.r_timer_reload[16] ;
 wire \cpu.intr.r_timer_reload[17] ;
 wire \cpu.intr.r_timer_reload[18] ;
 wire \cpu.intr.r_timer_reload[19] ;
 wire \cpu.intr.r_timer_reload[1] ;
 wire \cpu.intr.r_timer_reload[20] ;
 wire \cpu.intr.r_timer_reload[21] ;
 wire \cpu.intr.r_timer_reload[22] ;
 wire \cpu.intr.r_timer_reload[23] ;
 wire \cpu.intr.r_timer_reload[2] ;
 wire \cpu.intr.r_timer_reload[3] ;
 wire \cpu.intr.r_timer_reload[4] ;
 wire \cpu.intr.r_timer_reload[5] ;
 wire \cpu.intr.r_timer_reload[6] ;
 wire \cpu.intr.r_timer_reload[7] ;
 wire \cpu.intr.r_timer_reload[8] ;
 wire \cpu.intr.r_timer_reload[9] ;
 wire \cpu.intr.spi_intr ;
 wire \cpu.qspi.c_rstrobe_d ;
 wire \cpu.qspi.c_wstrobe_d ;
 wire \cpu.qspi.c_wstrobe_i ;
 wire \cpu.qspi.r_count[0] ;
 wire \cpu.qspi.r_count[1] ;
 wire \cpu.qspi.r_count[2] ;
 wire \cpu.qspi.r_count[3] ;
 wire \cpu.qspi.r_count[4] ;
 wire \cpu.qspi.r_ind ;
 wire \cpu.qspi.r_mask[0] ;
 wire \cpu.qspi.r_mask[1] ;
 wire \cpu.qspi.r_mask[2] ;
 wire \cpu.qspi.r_quad[0] ;
 wire \cpu.qspi.r_quad[1] ;
 wire \cpu.qspi.r_quad[2] ;
 wire \cpu.qspi.r_read_delay[0][0] ;
 wire \cpu.qspi.r_read_delay[0][1] ;
 wire \cpu.qspi.r_read_delay[0][2] ;
 wire \cpu.qspi.r_read_delay[0][3] ;
 wire \cpu.qspi.r_read_delay[1][0] ;
 wire \cpu.qspi.r_read_delay[1][1] ;
 wire \cpu.qspi.r_read_delay[1][2] ;
 wire \cpu.qspi.r_read_delay[1][3] ;
 wire \cpu.qspi.r_read_delay[2][0] ;
 wire \cpu.qspi.r_read_delay[2][1] ;
 wire \cpu.qspi.r_read_delay[2][2] ;
 wire \cpu.qspi.r_read_delay[2][3] ;
 wire \cpu.qspi.r_rom_mode[0] ;
 wire \cpu.qspi.r_rom_mode[1] ;
 wire \cpu.qspi.r_state[0] ;
 wire \cpu.qspi.r_state[10] ;
 wire \cpu.qspi.r_state[11] ;
 wire \cpu.qspi.r_state[12] ;
 wire \cpu.qspi.r_state[13] ;
 wire \cpu.qspi.r_state[14] ;
 wire \cpu.qspi.r_state[15] ;
 wire \cpu.qspi.r_state[16] ;
 wire \cpu.qspi.r_state[17] ;
 wire \cpu.qspi.r_state[1] ;
 wire \cpu.qspi.r_state[2] ;
 wire \cpu.qspi.r_state[3] ;
 wire \cpu.qspi.r_state[4] ;
 wire \cpu.qspi.r_state[5] ;
 wire \cpu.qspi.r_state[6] ;
 wire \cpu.qspi.r_state[7] ;
 wire \cpu.qspi.r_state[8] ;
 wire \cpu.qspi.r_state[9] ;
 wire \cpu.r_clk_invert ;
 wire \cpu.spi.r_bits[0] ;
 wire \cpu.spi.r_bits[1] ;
 wire \cpu.spi.r_bits[2] ;
 wire \cpu.spi.r_clk_count[0][0] ;
 wire \cpu.spi.r_clk_count[0][1] ;
 wire \cpu.spi.r_clk_count[0][2] ;
 wire \cpu.spi.r_clk_count[0][3] ;
 wire \cpu.spi.r_clk_count[0][4] ;
 wire \cpu.spi.r_clk_count[0][5] ;
 wire \cpu.spi.r_clk_count[0][6] ;
 wire \cpu.spi.r_clk_count[0][7] ;
 wire \cpu.spi.r_clk_count[1][0] ;
 wire \cpu.spi.r_clk_count[1][1] ;
 wire \cpu.spi.r_clk_count[1][2] ;
 wire \cpu.spi.r_clk_count[1][3] ;
 wire \cpu.spi.r_clk_count[1][4] ;
 wire \cpu.spi.r_clk_count[1][5] ;
 wire \cpu.spi.r_clk_count[1][6] ;
 wire \cpu.spi.r_clk_count[1][7] ;
 wire \cpu.spi.r_clk_count[2][0] ;
 wire \cpu.spi.r_clk_count[2][1] ;
 wire \cpu.spi.r_clk_count[2][2] ;
 wire \cpu.spi.r_clk_count[2][3] ;
 wire \cpu.spi.r_clk_count[2][4] ;
 wire \cpu.spi.r_clk_count[2][5] ;
 wire \cpu.spi.r_clk_count[2][6] ;
 wire \cpu.spi.r_clk_count[2][7] ;
 wire \cpu.spi.r_count[0] ;
 wire \cpu.spi.r_count[1] ;
 wire \cpu.spi.r_count[2] ;
 wire \cpu.spi.r_count[3] ;
 wire \cpu.spi.r_count[4] ;
 wire \cpu.spi.r_count[5] ;
 wire \cpu.spi.r_count[6] ;
 wire \cpu.spi.r_count[7] ;
 wire \cpu.spi.r_in[0] ;
 wire \cpu.spi.r_in[1] ;
 wire \cpu.spi.r_in[2] ;
 wire \cpu.spi.r_in[3] ;
 wire \cpu.spi.r_in[4] ;
 wire \cpu.spi.r_in[5] ;
 wire \cpu.spi.r_in[6] ;
 wire \cpu.spi.r_in[7] ;
 wire \cpu.spi.r_mode[0][0] ;
 wire \cpu.spi.r_mode[0][1] ;
 wire \cpu.spi.r_mode[1][0] ;
 wire \cpu.spi.r_mode[1][1] ;
 wire \cpu.spi.r_mode[2][0] ;
 wire \cpu.spi.r_mode[2][1] ;
 wire \cpu.spi.r_out[0] ;
 wire \cpu.spi.r_out[1] ;
 wire \cpu.spi.r_out[2] ;
 wire \cpu.spi.r_out[3] ;
 wire \cpu.spi.r_out[4] ;
 wire \cpu.spi.r_out[5] ;
 wire \cpu.spi.r_out[6] ;
 wire \cpu.spi.r_out[7] ;
 wire \cpu.spi.r_ready ;
 wire \cpu.spi.r_searching ;
 wire \cpu.spi.r_sel[0] ;
 wire \cpu.spi.r_sel[1] ;
 wire \cpu.spi.r_src[0] ;
 wire \cpu.spi.r_src[1] ;
 wire \cpu.spi.r_src[2] ;
 wire \cpu.spi.r_state[0] ;
 wire \cpu.spi.r_state[1] ;
 wire \cpu.spi.r_state[2] ;
 wire \cpu.spi.r_state[3] ;
 wire \cpu.spi.r_state[4] ;
 wire \cpu.spi.r_state[5] ;
 wire \cpu.spi.r_state[6] ;
 wire \cpu.spi.r_timeout[0] ;
 wire \cpu.spi.r_timeout[1] ;
 wire \cpu.spi.r_timeout[2] ;
 wire \cpu.spi.r_timeout[3] ;
 wire \cpu.spi.r_timeout[4] ;
 wire \cpu.spi.r_timeout[5] ;
 wire \cpu.spi.r_timeout[6] ;
 wire \cpu.spi.r_timeout[7] ;
 wire \cpu.spi.r_timeout_count[0] ;
 wire \cpu.spi.r_timeout_count[1] ;
 wire \cpu.spi.r_timeout_count[2] ;
 wire \cpu.spi.r_timeout_count[3] ;
 wire \cpu.spi.r_timeout_count[4] ;
 wire \cpu.spi.r_timeout_count[5] ;
 wire \cpu.spi.r_timeout_count[6] ;
 wire \cpu.spi.r_timeout_count[7] ;
 wire \cpu.uart.r_div[0] ;
 wire \cpu.uart.r_div[10] ;
 wire \cpu.uart.r_div[11] ;
 wire \cpu.uart.r_div[1] ;
 wire \cpu.uart.r_div[2] ;
 wire \cpu.uart.r_div[3] ;
 wire \cpu.uart.r_div[4] ;
 wire \cpu.uart.r_div[5] ;
 wire \cpu.uart.r_div[6] ;
 wire \cpu.uart.r_div[7] ;
 wire \cpu.uart.r_div[8] ;
 wire \cpu.uart.r_div[9] ;
 wire \cpu.uart.r_div_value[0] ;
 wire \cpu.uart.r_div_value[10] ;
 wire \cpu.uart.r_div_value[11] ;
 wire \cpu.uart.r_div_value[1] ;
 wire \cpu.uart.r_div_value[2] ;
 wire \cpu.uart.r_div_value[3] ;
 wire \cpu.uart.r_div_value[4] ;
 wire \cpu.uart.r_div_value[5] ;
 wire \cpu.uart.r_div_value[6] ;
 wire \cpu.uart.r_div_value[7] ;
 wire \cpu.uart.r_div_value[8] ;
 wire \cpu.uart.r_div_value[9] ;
 wire \cpu.uart.r_ib[0] ;
 wire \cpu.uart.r_ib[1] ;
 wire \cpu.uart.r_ib[2] ;
 wire \cpu.uart.r_ib[3] ;
 wire \cpu.uart.r_ib[4] ;
 wire \cpu.uart.r_ib[5] ;
 wire \cpu.uart.r_ib[6] ;
 wire \cpu.uart.r_in[0] ;
 wire \cpu.uart.r_in[1] ;
 wire \cpu.uart.r_in[2] ;
 wire \cpu.uart.r_in[3] ;
 wire \cpu.uart.r_in[4] ;
 wire \cpu.uart.r_in[5] ;
 wire \cpu.uart.r_in[6] ;
 wire \cpu.uart.r_in[7] ;
 wire \cpu.uart.r_out[0] ;
 wire \cpu.uart.r_out[1] ;
 wire \cpu.uart.r_out[2] ;
 wire \cpu.uart.r_out[3] ;
 wire \cpu.uart.r_out[4] ;
 wire \cpu.uart.r_out[5] ;
 wire \cpu.uart.r_out[6] ;
 wire \cpu.uart.r_out[7] ;
 wire \cpu.uart.r_r ;
 wire \cpu.uart.r_r_int ;
 wire \cpu.uart.r_r_invert ;
 wire \cpu.uart.r_rcnt[0] ;
 wire \cpu.uart.r_rcnt[1] ;
 wire \cpu.uart.r_rstate[0] ;
 wire \cpu.uart.r_rstate[1] ;
 wire \cpu.uart.r_rstate[2] ;
 wire \cpu.uart.r_rstate[3] ;
 wire \cpu.uart.r_x_int ;
 wire \cpu.uart.r_x_invert ;
 wire \cpu.uart.r_xcnt[0] ;
 wire \cpu.uart.r_xcnt[1] ;
 wire \cpu.uart.r_xstate[0] ;
 wire \cpu.uart.r_xstate[1] ;
 wire \cpu.uart.r_xstate[2] ;
 wire \cpu.uart.r_xstate[3] ;
 wire r_reset;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;

 sg13g2_buf_1 _14994_ (.A(\cpu.dec.r_op[5] ),
    .X(_08255_));
 sg13g2_buf_1 _14995_ (.A(_08255_),
    .X(_08256_));
 sg13g2_buf_1 _14996_ (.A(\cpu.ex.pc[1] ),
    .X(_08257_));
 sg13g2_buf_1 _14997_ (.A(_08257_),
    .X(_08258_));
 sg13g2_inv_1 _14998_ (.Y(_08259_),
    .A(_00204_));
 sg13g2_buf_2 _14999_ (.A(_00190_),
    .X(_08260_));
 sg13g2_buf_1 _15000_ (.A(net1130),
    .X(_08261_));
 sg13g2_buf_1 _15001_ (.A(\cpu.ex.pc[2] ),
    .X(_08262_));
 sg13g2_buf_1 _15002_ (.A(_08262_),
    .X(_08263_));
 sg13g2_buf_2 _15003_ (.A(\cpu.ex.pc[4] ),
    .X(_08264_));
 sg13g2_buf_1 _15004_ (.A(\cpu.ex.pc[3] ),
    .X(_08265_));
 sg13g2_nor2b_1 _15005_ (.A(_08264_),
    .B_N(_08265_),
    .Y(_08266_));
 sg13g2_buf_1 _15006_ (.A(_08265_),
    .X(_08267_));
 sg13g2_nand2b_1 _15007_ (.Y(_08268_),
    .B(_08264_),
    .A_N(net1069));
 sg13g2_o21ai_1 _15008_ (.B1(_08268_),
    .Y(_08269_),
    .A1(net1070),
    .A2(_08266_));
 sg13g2_and2_1 _15009_ (.A(net1071),
    .B(_08269_),
    .X(_08270_));
 sg13g2_buf_2 _15010_ (.A(_08270_),
    .X(_08271_));
 sg13g2_nor2_1 _15011_ (.A(_08263_),
    .B(net1130),
    .Y(_08272_));
 sg13g2_mux2_1 _15012_ (.A0(\cpu.icache.r_data[7][26] ),
    .A1(\cpu.icache.r_data[3][26] ),
    .S(net1130),
    .X(_08273_));
 sg13g2_a22oi_1 _15013_ (.Y(_08274_),
    .B1(_08273_),
    .B2(net1070),
    .A2(_08272_),
    .A1(\cpu.icache.r_data[6][26] ));
 sg13g2_buf_1 _15014_ (.A(_08267_),
    .X(_08275_));
 sg13g2_buf_2 _15015_ (.A(net931),
    .X(_08276_));
 sg13g2_nand2b_1 _15016_ (.Y(_08277_),
    .B(net797),
    .A_N(_08274_));
 sg13g2_inv_1 _15017_ (.Y(_08278_),
    .A(_08262_));
 sg13g2_buf_2 _15018_ (.A(_08278_),
    .X(_08279_));
 sg13g2_and2_1 _15019_ (.A(net930),
    .B(_08266_),
    .X(_08280_));
 sg13g2_buf_1 _15020_ (.A(_08280_),
    .X(_08281_));
 sg13g2_nor2_1 _15021_ (.A(_08265_),
    .B(net1130),
    .Y(_08282_));
 sg13g2_buf_1 _15022_ (.A(_08282_),
    .X(_08283_));
 sg13g2_and2_1 _15023_ (.A(net1070),
    .B(net929),
    .X(_08284_));
 sg13g2_buf_2 _15024_ (.A(_08284_),
    .X(_08285_));
 sg13g2_a22oi_1 _15025_ (.Y(_08286_),
    .B1(_08285_),
    .B2(\cpu.icache.r_data[5][26] ),
    .A2(_08281_),
    .A1(\cpu.icache.r_data[2][26] ));
 sg13g2_nor3_1 _15026_ (.A(_08278_),
    .B(net1069),
    .C(_08264_),
    .Y(_08287_));
 sg13g2_buf_2 _15027_ (.A(_08287_),
    .X(_08288_));
 sg13g2_nor3_1 _15028_ (.A(net1070),
    .B(net1069),
    .C(net1130),
    .Y(_08289_));
 sg13g2_buf_1 _15029_ (.A(_08289_),
    .X(_08290_));
 sg13g2_a22oi_1 _15030_ (.Y(_08291_),
    .B1(net796),
    .B2(\cpu.icache.r_data[4][26] ),
    .A2(_08288_),
    .A1(\cpu.icache.r_data[1][26] ));
 sg13g2_nand3_1 _15031_ (.B(_08286_),
    .C(_08291_),
    .A(_08277_),
    .Y(_08292_));
 sg13g2_a21oi_1 _15032_ (.A1(_08259_),
    .A2(_08271_),
    .Y(_08293_),
    .B1(_08292_));
 sg13g2_nand2_1 _15033_ (.Y(_08294_),
    .A(_00203_),
    .B(_08271_));
 sg13g2_nand2_1 _15034_ (.Y(_08295_),
    .A(net1071),
    .B(_08269_));
 sg13g2_and2_1 _15035_ (.A(net1070),
    .B(_08265_),
    .X(_08296_));
 sg13g2_buf_2 _15036_ (.A(_08296_),
    .X(_08297_));
 sg13g2_and2_1 _15037_ (.A(_08260_),
    .B(_08297_),
    .X(_08298_));
 sg13g2_buf_1 _15038_ (.A(_08298_),
    .X(_08299_));
 sg13g2_buf_1 _15039_ (.A(_08272_),
    .X(_08300_));
 sg13g2_mux2_1 _15040_ (.A0(\cpu.icache.r_data[4][10] ),
    .A1(\cpu.icache.r_data[6][10] ),
    .S(net1069),
    .X(_08301_));
 sg13g2_a22oi_1 _15041_ (.Y(_08302_),
    .B1(net795),
    .B2(_08301_),
    .A2(_08299_),
    .A1(\cpu.icache.r_data[3][10] ));
 sg13g2_a22oi_1 _15042_ (.Y(_08303_),
    .B1(_08281_),
    .B2(\cpu.icache.r_data[2][10] ),
    .A2(_08288_),
    .A1(\cpu.icache.r_data[1][10] ));
 sg13g2_nor2b_1 _15043_ (.A(_08260_),
    .B_N(_08297_),
    .Y(_08304_));
 sg13g2_buf_2 _15044_ (.A(_08304_),
    .X(_08305_));
 sg13g2_a22oi_1 _15045_ (.Y(_08306_),
    .B1(_08285_),
    .B2(\cpu.icache.r_data[5][10] ),
    .A2(_08305_),
    .A1(\cpu.icache.r_data[7][10] ));
 sg13g2_nand4_1 _15046_ (.B(_08302_),
    .C(_08303_),
    .A(_08295_),
    .Y(_08307_),
    .D(_08306_));
 sg13g2_a21oi_1 _15047_ (.A1(_08294_),
    .A2(_08307_),
    .Y(_08308_),
    .B1(net1072));
 sg13g2_a21oi_1 _15048_ (.A1(net1072),
    .A2(_08293_),
    .Y(_08309_),
    .B1(_08308_));
 sg13g2_buf_1 _15049_ (.A(_08309_),
    .X(_08310_));
 sg13g2_inv_2 _15050_ (.Y(_08311_),
    .A(_08310_));
 sg13g2_buf_1 _15051_ (.A(_08258_),
    .X(_08312_));
 sg13g2_buf_1 _15052_ (.A(_08312_),
    .X(_08313_));
 sg13g2_buf_1 _15053_ (.A(net796),
    .X(_08314_));
 sg13g2_buf_1 _15054_ (.A(_08297_),
    .X(_08315_));
 sg13g2_buf_1 _15055_ (.A(net1130),
    .X(_08316_));
 sg13g2_buf_1 _15056_ (.A(net1068),
    .X(_08317_));
 sg13g2_mux2_1 _15057_ (.A0(\cpu.icache.r_data[7][0] ),
    .A1(\cpu.icache.r_data[3][0] ),
    .S(net927),
    .X(_08318_));
 sg13g2_a22oi_1 _15058_ (.Y(_08319_),
    .B1(net704),
    .B2(_08318_),
    .A2(net705),
    .A1(\cpu.icache.r_data[4][0] ));
 sg13g2_buf_1 _15059_ (.A(_08288_),
    .X(_08320_));
 sg13g2_buf_1 _15060_ (.A(net703),
    .X(_08321_));
 sg13g2_buf_1 _15061_ (.A(_08281_),
    .X(_08322_));
 sg13g2_buf_1 _15062_ (.A(net640),
    .X(_08323_));
 sg13g2_a22oi_1 _15063_ (.Y(_08324_),
    .B1(net556),
    .B2(\cpu.icache.r_data[2][0] ),
    .A2(net641),
    .A1(\cpu.icache.r_data[1][0] ));
 sg13g2_and2_1 _15064_ (.A(net931),
    .B(_08272_),
    .X(_08325_));
 sg13g2_buf_2 _15065_ (.A(_08325_),
    .X(_08326_));
 sg13g2_buf_2 _15066_ (.A(_08326_),
    .X(_08327_));
 sg13g2_buf_1 _15067_ (.A(_08285_),
    .X(_08328_));
 sg13g2_buf_1 _15068_ (.A(net638),
    .X(_08329_));
 sg13g2_a22oi_1 _15069_ (.Y(_08330_),
    .B1(net555),
    .B2(\cpu.icache.r_data[5][0] ),
    .A2(net639),
    .A1(\cpu.icache.r_data[6][0] ));
 sg13g2_nand3_1 _15070_ (.B(_08324_),
    .C(_08330_),
    .A(_08319_),
    .Y(_08331_));
 sg13g2_buf_1 _15071_ (.A(_08295_),
    .X(_08332_));
 sg13g2_buf_1 _15072_ (.A(net637),
    .X(_08333_));
 sg13g2_mux2_1 _15073_ (.A0(\cpu.icache.r_data[0][0] ),
    .A1(_08331_),
    .S(net554),
    .X(_08334_));
 sg13g2_buf_1 _15074_ (.A(net1072),
    .X(_08335_));
 sg13g2_mux2_1 _15075_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(net927),
    .X(_08336_));
 sg13g2_buf_1 _15076_ (.A(net931),
    .X(_08337_));
 sg13g2_buf_1 _15077_ (.A(net793),
    .X(_08338_));
 sg13g2_a22oi_1 _15078_ (.Y(_08339_),
    .B1(_08336_),
    .B2(net702),
    .A2(net929),
    .A1(\cpu.icache.r_data[5][16] ));
 sg13g2_buf_1 _15079_ (.A(_08263_),
    .X(_08340_));
 sg13g2_buf_2 _15080_ (.A(net925),
    .X(_08341_));
 sg13g2_buf_1 _15081_ (.A(net792),
    .X(_08342_));
 sg13g2_nand2b_1 _15082_ (.Y(_08343_),
    .B(net701),
    .A_N(_08339_));
 sg13g2_buf_1 _15083_ (.A(_08271_),
    .X(_08344_));
 sg13g2_buf_1 _15084_ (.A(net553),
    .X(_08345_));
 sg13g2_a22oi_1 _15085_ (.Y(_08346_),
    .B1(net705),
    .B2(\cpu.icache.r_data[4][16] ),
    .A2(net641),
    .A1(\cpu.icache.r_data[1][16] ));
 sg13g2_buf_1 _15086_ (.A(_08281_),
    .X(_08347_));
 sg13g2_buf_1 _15087_ (.A(net636),
    .X(_08348_));
 sg13g2_a22oi_1 _15088_ (.Y(_08349_),
    .B1(net639),
    .B2(\cpu.icache.r_data[6][16] ),
    .A2(net552),
    .A1(\cpu.icache.r_data[2][16] ));
 sg13g2_nand2_1 _15089_ (.Y(_08350_),
    .A(_08346_),
    .B(_08349_));
 sg13g2_a21oi_1 _15090_ (.A1(\cpu.icache.r_data[0][16] ),
    .A2(net483),
    .Y(_08351_),
    .B1(_08350_));
 sg13g2_nand3_1 _15091_ (.B(_08343_),
    .C(_08351_),
    .A(net926),
    .Y(_08352_));
 sg13g2_o21ai_1 _15092_ (.B1(_08352_),
    .Y(_08353_),
    .A1(net794),
    .A2(_08334_));
 sg13g2_buf_2 _15093_ (.A(_08353_),
    .X(_08354_));
 sg13g2_buf_1 _15094_ (.A(_08288_),
    .X(_08355_));
 sg13g2_a22oi_1 _15095_ (.Y(_08356_),
    .B1(net640),
    .B2(\cpu.icache.r_data[2][1] ),
    .A2(net700),
    .A1(\cpu.icache.r_data[1][1] ));
 sg13g2_buf_2 _15096_ (.A(_08299_),
    .X(_08357_));
 sg13g2_a22oi_1 _15097_ (.Y(_08358_),
    .B1(_08326_),
    .B2(\cpu.icache.r_data[6][1] ),
    .A2(net551),
    .A1(\cpu.icache.r_data[3][1] ));
 sg13g2_nor2_1 _15098_ (.A(net1070),
    .B(net931),
    .Y(_08359_));
 sg13g2_mux2_1 _15099_ (.A0(\cpu.icache.r_data[5][1] ),
    .A1(\cpu.icache.r_data[7][1] ),
    .S(net1069),
    .X(_08360_));
 sg13g2_a22oi_1 _15100_ (.Y(_08361_),
    .B1(_08360_),
    .B2(net925),
    .A2(_08359_),
    .A1(\cpu.icache.r_data[4][1] ));
 sg13g2_or2_1 _15101_ (.X(_08362_),
    .B(_08361_),
    .A(net927));
 sg13g2_nand3_1 _15102_ (.B(_08358_),
    .C(_08362_),
    .A(_08356_),
    .Y(_08363_));
 sg13g2_buf_1 _15103_ (.A(_08332_),
    .X(_08364_));
 sg13g2_mux2_1 _15104_ (.A0(\cpu.icache.r_data[0][1] ),
    .A1(_08363_),
    .S(net550),
    .X(_08365_));
 sg13g2_buf_1 _15105_ (.A(net1071),
    .X(_08366_));
 sg13g2_mux2_1 _15106_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(net924),
    .X(_08367_));
 sg13g2_a22oi_1 _15107_ (.Y(_08368_),
    .B1(_08367_),
    .B2(net793),
    .A2(net929),
    .A1(\cpu.icache.r_data[5][17] ));
 sg13g2_nand2b_1 _15108_ (.Y(_08369_),
    .B(net701),
    .A_N(_08368_));
 sg13g2_buf_2 _15109_ (.A(net796),
    .X(_08370_));
 sg13g2_a22oi_1 _15110_ (.Y(_08371_),
    .B1(net699),
    .B2(\cpu.icache.r_data[4][17] ),
    .A2(net703),
    .A1(\cpu.icache.r_data[1][17] ));
 sg13g2_a22oi_1 _15111_ (.Y(_08372_),
    .B1(_08326_),
    .B2(\cpu.icache.r_data[6][17] ),
    .A2(net636),
    .A1(\cpu.icache.r_data[2][17] ));
 sg13g2_nand2_1 _15112_ (.Y(_08373_),
    .A(_08371_),
    .B(_08372_));
 sg13g2_a21oi_1 _15113_ (.A1(\cpu.icache.r_data[0][17] ),
    .A2(net553),
    .Y(_08374_),
    .B1(_08373_));
 sg13g2_nand3_1 _15114_ (.B(_08369_),
    .C(_08374_),
    .A(net1072),
    .Y(_08375_));
 sg13g2_o21ai_1 _15115_ (.B1(_08375_),
    .Y(_08376_),
    .A1(net928),
    .A2(_08365_));
 sg13g2_buf_2 _15116_ (.A(_08376_),
    .X(_08377_));
 sg13g2_inv_1 _15117_ (.Y(_08378_),
    .A(_08377_));
 sg13g2_buf_1 _15118_ (.A(_08378_),
    .X(_08379_));
 sg13g2_nor2_1 _15119_ (.A(_08354_),
    .B(net223),
    .Y(_08380_));
 sg13g2_buf_1 _15120_ (.A(_08380_),
    .X(_08381_));
 sg13g2_buf_1 _15121_ (.A(_08355_),
    .X(_08382_));
 sg13g2_a22oi_1 _15122_ (.Y(_08383_),
    .B1(net556),
    .B2(\cpu.icache.r_data[2][31] ),
    .A2(net635),
    .A1(\cpu.icache.r_data[1][31] ));
 sg13g2_mux2_1 _15123_ (.A0(\cpu.icache.r_data[7][31] ),
    .A1(\cpu.icache.r_data[3][31] ),
    .S(_08317_),
    .X(_08384_));
 sg13g2_a22oi_1 _15124_ (.Y(_08385_),
    .B1(net704),
    .B2(_08384_),
    .A2(_08314_),
    .A1(\cpu.icache.r_data[4][31] ));
 sg13g2_a22oi_1 _15125_ (.Y(_08386_),
    .B1(_08329_),
    .B2(\cpu.icache.r_data[5][31] ),
    .A2(net639),
    .A1(\cpu.icache.r_data[6][31] ));
 sg13g2_nand2b_1 _15126_ (.Y(_08387_),
    .B(net553),
    .A_N(_00202_));
 sg13g2_nand4_1 _15127_ (.B(_08385_),
    .C(_08386_),
    .A(_08383_),
    .Y(_08388_),
    .D(_08387_));
 sg13g2_inv_1 _15128_ (.Y(_08389_),
    .A(_08257_));
 sg13g2_buf_1 _15129_ (.A(_08389_),
    .X(_08390_));
 sg13g2_nand2_1 _15130_ (.Y(_08391_),
    .A(_00201_),
    .B(net553));
 sg13g2_buf_1 _15131_ (.A(net637),
    .X(_08392_));
 sg13g2_buf_1 _15132_ (.A(_08285_),
    .X(_08393_));
 sg13g2_a22oi_1 _15133_ (.Y(_08394_),
    .B1(net634),
    .B2(\cpu.icache.r_data[5][15] ),
    .A2(net705),
    .A1(\cpu.icache.r_data[4][15] ));
 sg13g2_a22oi_1 _15134_ (.Y(_08395_),
    .B1(net552),
    .B2(\cpu.icache.r_data[2][15] ),
    .A2(_08321_),
    .A1(\cpu.icache.r_data[1][15] ));
 sg13g2_mux2_1 _15135_ (.A0(\cpu.icache.r_data[7][15] ),
    .A1(\cpu.icache.r_data[3][15] ),
    .S(net1068),
    .X(_08396_));
 sg13g2_buf_1 _15136_ (.A(net925),
    .X(_08397_));
 sg13g2_a22oi_1 _15137_ (.Y(_08398_),
    .B1(_08396_),
    .B2(net791),
    .A2(net795),
    .A1(\cpu.icache.r_data[6][15] ));
 sg13g2_buf_1 _15138_ (.A(net797),
    .X(_08399_));
 sg13g2_nand2b_1 _15139_ (.Y(_08400_),
    .B(net698),
    .A_N(_08398_));
 sg13g2_nand4_1 _15140_ (.B(_08394_),
    .C(_08395_),
    .A(net549),
    .Y(_08401_),
    .D(_08400_));
 sg13g2_and3_1 _15141_ (.X(_08402_),
    .A(net923),
    .B(_08391_),
    .C(_08401_));
 sg13g2_a21oi_1 _15142_ (.A1(net926),
    .A2(_08388_),
    .Y(_08403_),
    .B1(_08402_));
 sg13g2_buf_1 _15143_ (.A(_08403_),
    .X(_08404_));
 sg13g2_nand2_1 _15144_ (.Y(_08405_),
    .A(\cpu.icache.r_data[0][14] ),
    .B(_08271_));
 sg13g2_mux4_1 _15145_ (.S0(net925),
    .A0(\cpu.icache.r_data[4][14] ),
    .A1(\cpu.icache.r_data[5][14] ),
    .A2(\cpu.icache.r_data[6][14] ),
    .A3(\cpu.icache.r_data[7][14] ),
    .S1(net797),
    .X(_08406_));
 sg13g2_nand2b_1 _15146_ (.Y(_08407_),
    .B(_08406_),
    .A_N(net927));
 sg13g2_nand2_1 _15147_ (.Y(_08408_),
    .A(\cpu.icache.r_data[2][14] ),
    .B(net552));
 sg13g2_a22oi_1 _15148_ (.Y(_08409_),
    .B1(net551),
    .B2(\cpu.icache.r_data[3][14] ),
    .A2(net700),
    .A1(\cpu.icache.r_data[1][14] ));
 sg13g2_nand4_1 _15149_ (.B(_08407_),
    .C(_08408_),
    .A(_08405_),
    .Y(_08410_),
    .D(_08409_));
 sg13g2_nand2_1 _15150_ (.Y(_08411_),
    .A(\cpu.icache.r_data[0][30] ),
    .B(_08271_));
 sg13g2_mux2_1 _15151_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(net1071),
    .X(_08412_));
 sg13g2_a22oi_1 _15152_ (.Y(_08413_),
    .B1(_08412_),
    .B2(_08340_),
    .A2(_08300_),
    .A1(\cpu.icache.r_data[6][30] ));
 sg13g2_nand2b_1 _15153_ (.Y(_08414_),
    .B(net793),
    .A_N(_08413_));
 sg13g2_a22oi_1 _15154_ (.Y(_08415_),
    .B1(net796),
    .B2(\cpu.icache.r_data[4][30] ),
    .A2(net703),
    .A1(\cpu.icache.r_data[1][30] ));
 sg13g2_a22oi_1 _15155_ (.Y(_08416_),
    .B1(net638),
    .B2(\cpu.icache.r_data[5][30] ),
    .A2(net636),
    .A1(\cpu.icache.r_data[2][30] ));
 sg13g2_nand4_1 _15156_ (.B(_08414_),
    .C(_08415_),
    .A(_08411_),
    .Y(_08417_),
    .D(_08416_));
 sg13g2_or2_1 _15157_ (.X(_08418_),
    .B(_08417_),
    .A(_08389_));
 sg13g2_o21ai_1 _15158_ (.B1(_08418_),
    .Y(_08419_),
    .A1(net928),
    .A2(_08410_));
 sg13g2_buf_1 _15159_ (.A(_08419_),
    .X(_08420_));
 sg13g2_mux2_1 _15160_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(net1068),
    .X(_08421_));
 sg13g2_a22oi_1 _15161_ (.Y(_08422_),
    .B1(_08421_),
    .B2(net791),
    .A2(net795),
    .A1(\cpu.icache.r_data[6][29] ));
 sg13g2_nand2b_1 _15162_ (.Y(_08423_),
    .B(net698),
    .A_N(_08422_));
 sg13g2_a22oi_1 _15163_ (.Y(_08424_),
    .B1(net640),
    .B2(\cpu.icache.r_data[2][29] ),
    .A2(net699),
    .A1(\cpu.icache.r_data[4][29] ));
 sg13g2_a22oi_1 _15164_ (.Y(_08425_),
    .B1(net638),
    .B2(\cpu.icache.r_data[5][29] ),
    .A2(net700),
    .A1(\cpu.icache.r_data[1][29] ));
 sg13g2_nand3_1 _15165_ (.B(_08424_),
    .C(_08425_),
    .A(_08423_),
    .Y(_08426_));
 sg13g2_a21oi_1 _15166_ (.A1(\cpu.icache.r_data[0][29] ),
    .A2(net483),
    .Y(_08427_),
    .B1(_08426_));
 sg13g2_nand2b_1 _15167_ (.Y(_08428_),
    .B(net553),
    .A_N(\cpu.icache.r_data[0][13] ));
 sg13g2_a22oi_1 _15168_ (.Y(_08429_),
    .B1(net638),
    .B2(\cpu.icache.r_data[5][13] ),
    .A2(net700),
    .A1(\cpu.icache.r_data[1][13] ));
 sg13g2_a22oi_1 _15169_ (.Y(_08430_),
    .B1(net551),
    .B2(\cpu.icache.r_data[3][13] ),
    .A2(net640),
    .A1(\cpu.icache.r_data[2][13] ));
 sg13g2_mux2_1 _15170_ (.A0(\cpu.icache.r_data[4][13] ),
    .A1(\cpu.icache.r_data[6][13] ),
    .S(net931),
    .X(_08431_));
 sg13g2_a22oi_1 _15171_ (.Y(_08432_),
    .B1(_08431_),
    .B2(net930),
    .A2(_08297_),
    .A1(\cpu.icache.r_data[7][13] ));
 sg13g2_or2_1 _15172_ (.X(_08433_),
    .B(_08432_),
    .A(net927));
 sg13g2_nand4_1 _15173_ (.B(_08429_),
    .C(_08430_),
    .A(net550),
    .Y(_08434_),
    .D(_08433_));
 sg13g2_a21oi_1 _15174_ (.A1(_08428_),
    .A2(_08434_),
    .Y(_08435_),
    .B1(net1072));
 sg13g2_a21o_1 _15175_ (.A2(_08427_),
    .A1(net926),
    .B1(_08435_),
    .X(_08436_));
 sg13g2_buf_1 _15176_ (.A(_08436_),
    .X(_08437_));
 sg13g2_nand2_1 _15177_ (.Y(_08438_),
    .A(_08420_),
    .B(_08437_));
 sg13g2_nor2_1 _15178_ (.A(_08404_),
    .B(_08438_),
    .Y(_08439_));
 sg13g2_buf_2 _15179_ (.A(_08439_),
    .X(_08440_));
 sg13g2_nand2_1 _15180_ (.Y(_08441_),
    .A(net172),
    .B(_08440_));
 sg13g2_inv_1 _15181_ (.Y(_08442_),
    .A(_00206_));
 sg13g2_mux2_1 _15182_ (.A0(\cpu.icache.r_data[7][27] ),
    .A1(\cpu.icache.r_data[3][27] ),
    .S(net1071),
    .X(_08443_));
 sg13g2_a22oi_1 _15183_ (.Y(_08444_),
    .B1(_08443_),
    .B2(net925),
    .A2(_08300_),
    .A1(\cpu.icache.r_data[6][27] ));
 sg13g2_nand2b_1 _15184_ (.Y(_08445_),
    .B(net793),
    .A_N(_08444_));
 sg13g2_a22oi_1 _15185_ (.Y(_08446_),
    .B1(_08370_),
    .B2(\cpu.icache.r_data[4][27] ),
    .A2(net703),
    .A1(\cpu.icache.r_data[1][27] ));
 sg13g2_a22oi_1 _15186_ (.Y(_08447_),
    .B1(net638),
    .B2(\cpu.icache.r_data[5][27] ),
    .A2(net636),
    .A1(\cpu.icache.r_data[2][27] ));
 sg13g2_nand3_1 _15187_ (.B(_08446_),
    .C(_08447_),
    .A(_08445_),
    .Y(_08448_));
 sg13g2_a21oi_1 _15188_ (.A1(_08442_),
    .A2(net553),
    .Y(_08449_),
    .B1(_08448_));
 sg13g2_nand2_1 _15189_ (.Y(_08450_),
    .A(_00205_),
    .B(_08271_));
 sg13g2_a22oi_1 _15190_ (.Y(_08451_),
    .B1(net638),
    .B2(\cpu.icache.r_data[5][11] ),
    .A2(net796),
    .A1(\cpu.icache.r_data[4][11] ));
 sg13g2_a22oi_1 _15191_ (.Y(_08452_),
    .B1(net636),
    .B2(\cpu.icache.r_data[2][11] ),
    .A2(net703),
    .A1(\cpu.icache.r_data[1][11] ));
 sg13g2_mux2_1 _15192_ (.A0(\cpu.icache.r_data[7][11] ),
    .A1(\cpu.icache.r_data[3][11] ),
    .S(net1071),
    .X(_08453_));
 sg13g2_a22oi_1 _15193_ (.Y(_08454_),
    .B1(_08453_),
    .B2(net925),
    .A2(net795),
    .A1(\cpu.icache.r_data[6][11] ));
 sg13g2_nand2b_1 _15194_ (.Y(_08455_),
    .B(net793),
    .A_N(_08454_));
 sg13g2_nand4_1 _15195_ (.B(_08451_),
    .C(_08452_),
    .A(net637),
    .Y(_08456_),
    .D(_08455_));
 sg13g2_a21oi_1 _15196_ (.A1(_08450_),
    .A2(_08456_),
    .Y(_08457_),
    .B1(net1072));
 sg13g2_a21oi_1 _15197_ (.A1(net928),
    .A2(_08449_),
    .Y(_08458_),
    .B1(_08457_));
 sg13g2_buf_1 _15198_ (.A(_08458_),
    .X(_08459_));
 sg13g2_buf_1 _15199_ (.A(net336),
    .X(_08460_));
 sg13g2_nor3_1 _15200_ (.A(_08311_),
    .B(_08441_),
    .C(net295),
    .Y(_08461_));
 sg13g2_buf_2 _15201_ (.A(_00189_),
    .X(_08462_));
 sg13g2_buf_1 _15202_ (.A(\cpu.ex.genblk3.r_mmu_enable ),
    .X(_08463_));
 sg13g2_inv_2 _15203_ (.Y(_08464_),
    .A(net1129));
 sg13g2_buf_1 _15204_ (.A(\cpu.ex.io_access ),
    .X(_08465_));
 sg13g2_buf_2 _15205_ (.A(\cpu.ex.r_wmask[1] ),
    .X(_08466_));
 sg13g2_nor2_1 _15206_ (.A(_08466_),
    .B(\cpu.ex.r_wmask[0] ),
    .Y(_08467_));
 sg13g2_buf_2 _15207_ (.A(_08467_),
    .X(_08468_));
 sg13g2_nor3_1 _15208_ (.A(_08464_),
    .B(_08465_),
    .C(_08468_),
    .Y(_08469_));
 sg13g2_buf_1 _15209_ (.A(\cpu.addr[15] ),
    .X(_08470_));
 sg13g2_inv_1 _15210_ (.Y(_08471_),
    .A(_08470_));
 sg13g2_buf_2 _15211_ (.A(_08471_),
    .X(_08472_));
 sg13g2_buf_8 _15212_ (.A(\cpu.ex.ifetch ),
    .X(_08473_));
 sg13g2_inv_2 _15213_ (.Y(_08474_),
    .A(net1128));
 sg13g2_buf_1 _15214_ (.A(\cpu.ex.genblk3.r_mmu_d_proxy ),
    .X(_08475_));
 sg13g2_buf_2 _15215_ (.A(_00193_),
    .X(_08476_));
 sg13g2_a21oi_1 _15216_ (.A1(_08474_),
    .A2(_08475_),
    .Y(_08477_),
    .B1(_08476_));
 sg13g2_buf_1 _15217_ (.A(_08477_),
    .X(_08478_));
 sg13g2_buf_2 _15218_ (.A(\cpu.addr[13] ),
    .X(_08479_));
 sg13g2_buf_8 _15219_ (.A(\cpu.addr[12] ),
    .X(_08480_));
 sg13g2_buf_8 _15220_ (.A(_08480_),
    .X(_08481_));
 sg13g2_nand2b_1 _15221_ (.Y(_08482_),
    .B(net1067),
    .A_N(_08479_));
 sg13g2_buf_1 _15222_ (.A(_08482_),
    .X(_08483_));
 sg13g2_buf_8 _15223_ (.A(\cpu.addr[14] ),
    .X(_08484_));
 sg13g2_buf_8 _15224_ (.A(_08484_),
    .X(_08485_));
 sg13g2_mux2_1 _15225_ (.A0(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .S(net1066),
    .X(_08486_));
 sg13g2_nor2_1 _15226_ (.A(_08483_),
    .B(_08486_),
    .Y(_08487_));
 sg13g2_nor3_1 _15227_ (.A(_08472_),
    .B(_08478_),
    .C(_08487_),
    .Y(_08488_));
 sg13g2_inv_1 _15228_ (.Y(_08489_),
    .A(_08479_));
 sg13g2_nor2_1 _15229_ (.A(net1067),
    .B(_08489_),
    .Y(_08490_));
 sg13g2_buf_1 _15230_ (.A(_08484_),
    .X(_08491_));
 sg13g2_buf_1 _15231_ (.A(_08484_),
    .X(_08492_));
 sg13g2_nand2b_1 _15232_ (.Y(_08493_),
    .B(net1064),
    .A_N(\cpu.genblk1.mmu.r_writeable_d[14] ));
 sg13g2_o21ai_1 _15233_ (.B1(_08493_),
    .Y(_08494_),
    .A1(net1065),
    .A2(\cpu.genblk1.mmu.r_writeable_d[10] ));
 sg13g2_buf_8 _15234_ (.A(_08479_),
    .X(_08495_));
 sg13g2_nor2_1 _15235_ (.A(net1067),
    .B(_08495_),
    .Y(_08496_));
 sg13g2_nand2b_1 _15236_ (.Y(_08497_),
    .B(net1064),
    .A_N(\cpu.genblk1.mmu.r_writeable_d[12] ));
 sg13g2_o21ai_1 _15237_ (.B1(_08497_),
    .Y(_08498_),
    .A1(net1065),
    .A2(\cpu.genblk1.mmu.r_writeable_d[8] ));
 sg13g2_nand2_1 _15238_ (.Y(_08499_),
    .A(net1067),
    .B(net1063));
 sg13g2_mux2_1 _15239_ (.A0(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .S(net1066),
    .X(_08500_));
 sg13g2_nor2_1 _15240_ (.A(_08499_),
    .B(_08500_),
    .Y(_08501_));
 sg13g2_a221oi_1 _15241_ (.B2(_08498_),
    .C1(_08501_),
    .B1(_08496_),
    .A1(_08490_),
    .Y(_08502_),
    .A2(_08494_));
 sg13g2_a21o_1 _15242_ (.A2(_08475_),
    .A1(_08474_),
    .B1(_08476_),
    .X(_08503_));
 sg13g2_buf_4 _15243_ (.X(_08504_),
    .A(_08503_));
 sg13g2_mux2_1 _15244_ (.A0(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .S(net1064),
    .X(_08505_));
 sg13g2_nor2_1 _15245_ (.A(_08499_),
    .B(_08505_),
    .Y(_08506_));
 sg13g2_nor3_1 _15246_ (.A(_08472_),
    .B(_08504_),
    .C(_08506_),
    .Y(_08507_));
 sg13g2_nand2b_1 _15247_ (.Y(_08508_),
    .B(net1064),
    .A_N(\cpu.genblk1.mmu.r_writeable_d[28] ));
 sg13g2_o21ai_1 _15248_ (.B1(_08508_),
    .Y(_08509_),
    .A1(net1065),
    .A2(\cpu.genblk1.mmu.r_writeable_d[24] ));
 sg13g2_nand2b_1 _15249_ (.Y(_08510_),
    .B(net1065),
    .A_N(\cpu.genblk1.mmu.r_writeable_d[30] ));
 sg13g2_o21ai_1 _15250_ (.B1(_08510_),
    .Y(_08511_),
    .A1(net1065),
    .A2(\cpu.genblk1.mmu.r_writeable_d[26] ));
 sg13g2_mux2_1 _15251_ (.A0(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .S(net1066),
    .X(_08512_));
 sg13g2_nor2_1 _15252_ (.A(_08483_),
    .B(_08512_),
    .Y(_08513_));
 sg13g2_a221oi_1 _15253_ (.B2(_08490_),
    .C1(_08513_),
    .B1(_08511_),
    .A1(_08496_),
    .Y(_08514_),
    .A2(_08509_));
 sg13g2_a22oi_1 _15254_ (.Y(_08515_),
    .B1(_08507_),
    .B2(_08514_),
    .A2(_08502_),
    .A1(_08488_));
 sg13g2_mux2_1 _15255_ (.A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .S(net1064),
    .X(_08516_));
 sg13g2_or2_1 _15256_ (.X(_08517_),
    .B(_08516_),
    .A(_08483_));
 sg13g2_nand2b_1 _15257_ (.Y(_08518_),
    .B(net1066),
    .A_N(\cpu.genblk1.mmu.r_writeable_d[6] ));
 sg13g2_o21ai_1 _15258_ (.B1(_08518_),
    .Y(_08519_),
    .A1(net1065),
    .A2(\cpu.genblk1.mmu.r_writeable_d[2] ));
 sg13g2_nand2b_1 _15259_ (.Y(_08520_),
    .B(net1064),
    .A_N(\cpu.genblk1.mmu.r_writeable_d[4] ));
 sg13g2_o21ai_1 _15260_ (.B1(_08520_),
    .Y(_08521_),
    .A1(_08491_),
    .A2(\cpu.genblk1.mmu.r_writeable_d[0] ));
 sg13g2_mux2_1 _15261_ (.A0(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .S(net1066),
    .X(_08522_));
 sg13g2_nor2_1 _15262_ (.A(_08499_),
    .B(_08522_),
    .Y(_08523_));
 sg13g2_a221oi_1 _15263_ (.B2(_08496_),
    .C1(_08523_),
    .B1(_08521_),
    .A1(_08490_),
    .Y(_08524_),
    .A2(_08519_));
 sg13g2_nand4_1 _15264_ (.B(_08504_),
    .C(_08517_),
    .A(_08472_),
    .Y(_08525_),
    .D(_08524_));
 sg13g2_mux2_1 _15265_ (.A0(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .S(net1064),
    .X(_08526_));
 sg13g2_or2_1 _15266_ (.X(_08527_),
    .B(_08526_),
    .A(_08499_));
 sg13g2_nand2b_1 _15267_ (.Y(_08528_),
    .B(_08485_),
    .A_N(\cpu.genblk1.mmu.r_writeable_d[20] ));
 sg13g2_o21ai_1 _15268_ (.B1(_08528_),
    .Y(_08529_),
    .A1(net1065),
    .A2(\cpu.genblk1.mmu.r_writeable_d[16] ));
 sg13g2_nand2b_1 _15269_ (.Y(_08530_),
    .B(net1064),
    .A_N(\cpu.genblk1.mmu.r_writeable_d[22] ));
 sg13g2_o21ai_1 _15270_ (.B1(_08530_),
    .Y(_08531_),
    .A1(net1065),
    .A2(\cpu.genblk1.mmu.r_writeable_d[18] ));
 sg13g2_mux2_1 _15271_ (.A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .S(_08485_),
    .X(_08532_));
 sg13g2_nor2_1 _15272_ (.A(_08483_),
    .B(_08532_),
    .Y(_08533_));
 sg13g2_a221oi_1 _15273_ (.B2(_08490_),
    .C1(_08533_),
    .B1(_08531_),
    .A1(_08496_),
    .Y(_08534_),
    .A2(_08529_));
 sg13g2_nand4_1 _15274_ (.B(_08478_),
    .C(_08527_),
    .A(_08472_),
    .Y(_08535_),
    .D(_08534_));
 sg13g2_nand4_1 _15275_ (.B(_08515_),
    .C(_08525_),
    .A(_08469_),
    .Y(_08536_),
    .D(_08535_));
 sg13g2_buf_2 _15276_ (.A(_08536_),
    .X(_08537_));
 sg13g2_buf_4 _15277_ (.X(_08538_),
    .A(\cpu.ex.pc[15] ));
 sg13g2_buf_8 _15278_ (.A(\cpu.ex.pc[14] ),
    .X(_08539_));
 sg13g2_buf_8 _15279_ (.A(_08539_),
    .X(_08540_));
 sg13g2_mux2_1 _15280_ (.A0(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[20] ),
    .S(net1062),
    .X(_08541_));
 sg13g2_mux2_1 _15281_ (.A0(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[22] ),
    .S(_08540_),
    .X(_08542_));
 sg13g2_mux2_1 _15282_ (.A0(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[21] ),
    .S(net1062),
    .X(_08543_));
 sg13g2_mux2_1 _15283_ (.A0(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[23] ),
    .S(_08540_),
    .X(_08544_));
 sg13g2_buf_4 _15284_ (.X(_08545_),
    .A(\cpu.ex.pc[13] ));
 sg13g2_buf_2 _15285_ (.A(\cpu.ex.pc[12] ),
    .X(_08546_));
 sg13g2_buf_2 _15286_ (.A(_08546_),
    .X(_08547_));
 sg13g2_mux4_1 _15287_ (.S0(_08545_),
    .A0(_08541_),
    .A1(_08542_),
    .A2(_08543_),
    .A3(_08544_),
    .S1(_08547_),
    .X(_08548_));
 sg13g2_buf_1 _15288_ (.A(\cpu.dec.supmode ),
    .X(_08549_));
 sg13g2_nand3_1 _15289_ (.B(net1129),
    .C(_08473_),
    .A(net1127),
    .Y(_08550_));
 sg13g2_or3_1 _15290_ (.A(_08538_),
    .B(_08548_),
    .C(_08550_),
    .X(_08551_));
 sg13g2_nand2_1 _15291_ (.Y(_08552_),
    .A(\cpu.ex.genblk3.r_mmu_enable ),
    .B(net1128));
 sg13g2_mux2_1 _15292_ (.A0(\cpu.genblk1.mmu.r_valid_i[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[4] ),
    .S(_08539_),
    .X(_08553_));
 sg13g2_mux2_1 _15293_ (.A0(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[6] ),
    .S(_08539_),
    .X(_08554_));
 sg13g2_mux2_1 _15294_ (.A0(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[5] ),
    .S(_08539_),
    .X(_08555_));
 sg13g2_mux2_1 _15295_ (.A0(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[7] ),
    .S(_08539_),
    .X(_08556_));
 sg13g2_mux4_1 _15296_ (.S0(_08545_),
    .A0(_08553_),
    .A1(_08554_),
    .A2(_08555_),
    .A3(_08556_),
    .S1(_08546_),
    .X(_08557_));
 sg13g2_or4_1 _15297_ (.A(_08538_),
    .B(net1127),
    .C(_08552_),
    .D(_08557_),
    .X(_08558_));
 sg13g2_inv_2 _15298_ (.Y(_08559_),
    .A(_08538_));
 sg13g2_buf_8 _15299_ (.A(_08539_),
    .X(_08560_));
 sg13g2_mux2_1 _15300_ (.A0(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[28] ),
    .S(_08560_),
    .X(_08561_));
 sg13g2_mux2_1 _15301_ (.A0(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[29] ),
    .S(_08560_),
    .X(_08562_));
 sg13g2_mux2_1 _15302_ (.A0(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[30] ),
    .S(net1062),
    .X(_08563_));
 sg13g2_mux2_1 _15303_ (.A0(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[31] ),
    .S(net1062),
    .X(_08564_));
 sg13g2_mux4_1 _15304_ (.S0(_08546_),
    .A0(_08561_),
    .A1(_08562_),
    .A2(_08563_),
    .A3(_08564_),
    .S1(_08545_),
    .X(_08565_));
 sg13g2_or3_1 _15305_ (.A(_08559_),
    .B(_08550_),
    .C(_08565_),
    .X(_08566_));
 sg13g2_mux2_1 _15306_ (.A0(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[12] ),
    .S(net1062),
    .X(_08567_));
 sg13g2_mux2_1 _15307_ (.A0(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[13] ),
    .S(net1062),
    .X(_08568_));
 sg13g2_mux2_1 _15308_ (.A0(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[14] ),
    .S(net1062),
    .X(_08569_));
 sg13g2_mux2_1 _15309_ (.A0(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[15] ),
    .S(net1062),
    .X(_08570_));
 sg13g2_mux4_1 _15310_ (.S0(_08546_),
    .A0(_08567_),
    .A1(_08568_),
    .A2(_08569_),
    .A3(_08570_),
    .S1(_08545_),
    .X(_08571_));
 sg13g2_or4_1 _15311_ (.A(_08559_),
    .B(net1127),
    .C(_08552_),
    .D(_08571_),
    .X(_08572_));
 sg13g2_nand4_1 _15312_ (.B(_08558_),
    .C(_08566_),
    .A(_08551_),
    .Y(_08573_),
    .D(_08572_));
 sg13g2_buf_2 _15313_ (.A(_08573_),
    .X(_08574_));
 sg13g2_buf_1 _15314_ (.A(\cpu.ex.r_read_stall ),
    .X(_08575_));
 sg13g2_inv_2 _15315_ (.Y(_08576_),
    .A(_08575_));
 sg13g2_nand3_1 _15316_ (.B(_08576_),
    .C(_08468_),
    .A(_08462_),
    .Y(_08577_));
 sg13g2_inv_1 _15317_ (.Y(_08578_),
    .A(_08462_));
 sg13g2_buf_1 _15318_ (.A(_08575_),
    .X(_08579_));
 sg13g2_buf_8 _15319_ (.A(_00198_),
    .X(_08580_));
 sg13g2_a21o_1 _15320_ (.A2(\cpu.cond[0] ),
    .A1(\cpu.ex.mmu_reg_data[0] ),
    .B1(_08580_),
    .X(_08581_));
 sg13g2_buf_1 _15321_ (.A(\cpu.ex.mmu_reg_data[0] ),
    .X(_08582_));
 sg13g2_buf_1 _15322_ (.A(\cpu.cond[0] ),
    .X(_08583_));
 sg13g2_nor2b_1 _15323_ (.A(net1126),
    .B_N(net1125),
    .Y(_08584_));
 sg13g2_nand2_1 _15324_ (.Y(_08585_),
    .A(net1129),
    .B(_00197_));
 sg13g2_a221oi_1 _15325_ (.B2(_08580_),
    .C1(_08585_),
    .B1(_08584_),
    .A1(_08576_),
    .Y(_08586_),
    .A2(_08581_));
 sg13g2_o21ai_1 _15326_ (.B1(_08586_),
    .Y(_08587_),
    .A1(_08578_),
    .A2(net1060));
 sg13g2_buf_1 _15327_ (.A(_08470_),
    .X(_08588_));
 sg13g2_mux4_1 _15328_ (.S0(net1067),
    .A0(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[31] ),
    .S1(net1066),
    .X(_08589_));
 sg13g2_nand3_1 _15329_ (.B(net1059),
    .C(_08589_),
    .A(net1063),
    .Y(_08590_));
 sg13g2_mux4_1 _15330_ (.S0(net1067),
    .A0(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[23] ),
    .S1(_08484_),
    .X(_08591_));
 sg13g2_nand3_1 _15331_ (.B(_08472_),
    .C(_08591_),
    .A(net1063),
    .Y(_08592_));
 sg13g2_mux4_1 _15332_ (.S0(_08480_),
    .A0(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[29] ),
    .S1(_08484_),
    .X(_08593_));
 sg13g2_nor2b_1 _15333_ (.A(net1063),
    .B_N(_08470_),
    .Y(_08594_));
 sg13g2_mux4_1 _15334_ (.S0(net1067),
    .A0(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[21] ),
    .S1(net1066),
    .X(_08595_));
 sg13g2_nor2_1 _15335_ (.A(net1063),
    .B(net1059),
    .Y(_08596_));
 sg13g2_a22oi_1 _15336_ (.Y(_08597_),
    .B1(_08595_),
    .B2(_08596_),
    .A2(_08594_),
    .A1(_08593_));
 sg13g2_nand4_1 _15337_ (.B(_08590_),
    .C(_08592_),
    .A(_08478_),
    .Y(_08598_),
    .D(_08597_));
 sg13g2_buf_1 _15338_ (.A(net1066),
    .X(_08599_));
 sg13g2_mux4_1 _15339_ (.S0(net1067),
    .A0(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[15] ),
    .S1(net1063),
    .X(_08600_));
 sg13g2_nand3_1 _15340_ (.B(net1059),
    .C(_08600_),
    .A(net922),
    .Y(_08601_));
 sg13g2_mux4_1 _15341_ (.S0(_08480_),
    .A0(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[7] ),
    .S1(net1063),
    .X(_08602_));
 sg13g2_nand3_1 _15342_ (.B(_08472_),
    .C(_08602_),
    .A(_08491_),
    .Y(_08603_));
 sg13g2_mux4_1 _15343_ (.S0(_08480_),
    .A0(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[11] ),
    .S1(_08479_),
    .X(_08604_));
 sg13g2_nor2b_1 _15344_ (.A(_08492_),
    .B_N(_08470_),
    .Y(_08605_));
 sg13g2_mux4_1 _15345_ (.S0(_08480_),
    .A0(\cpu.genblk1.mmu.r_valid_d[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[2] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[3] ),
    .S1(net1063),
    .X(_08606_));
 sg13g2_nor2_1 _15346_ (.A(_08492_),
    .B(net1059),
    .Y(_08607_));
 sg13g2_a22oi_1 _15347_ (.Y(_08608_),
    .B1(_08606_),
    .B2(_08607_),
    .A2(_08605_),
    .A1(_08604_));
 sg13g2_nand4_1 _15348_ (.B(_08601_),
    .C(_08603_),
    .A(_08504_),
    .Y(_08609_),
    .D(_08608_));
 sg13g2_inv_1 _15349_ (.Y(_08610_),
    .A(_08465_));
 sg13g2_a21oi_1 _15350_ (.A1(net1129),
    .A2(net1058),
    .Y(_08611_),
    .B1(_08586_));
 sg13g2_a221oi_1 _15351_ (.B2(_08609_),
    .C1(_08611_),
    .B1(_08598_),
    .A1(_08468_),
    .Y(_08612_),
    .A2(_08587_));
 sg13g2_a21oi_2 _15352_ (.B1(_08612_),
    .Y(_08613_),
    .A2(_08577_),
    .A1(_08574_));
 sg13g2_nand2_1 _15353_ (.Y(_08614_),
    .A(_08537_),
    .B(_08613_));
 sg13g2_buf_1 _15354_ (.A(_08614_),
    .X(_08615_));
 sg13g2_buf_1 _15355_ (.A(_08615_),
    .X(_08616_));
 sg13g2_buf_2 _15356_ (.A(_08547_),
    .X(_08617_));
 sg13g2_buf_1 _15357_ (.A(net921),
    .X(_08618_));
 sg13g2_buf_1 _15358_ (.A(net1129),
    .X(_08619_));
 sg13g2_buf_1 _15359_ (.A(net1127),
    .X(_08620_));
 sg13g2_buf_1 _15360_ (.A(net1056),
    .X(_08621_));
 sg13g2_buf_2 _15361_ (.A(_08547_),
    .X(_08622_));
 sg13g2_buf_2 _15362_ (.A(net919),
    .X(_08623_));
 sg13g2_buf_1 _15363_ (.A(_08545_),
    .X(_08624_));
 sg13g2_buf_1 _15364_ (.A(net1055),
    .X(_08625_));
 sg13g2_mux4_1 _15365_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .S1(net918),
    .X(_08626_));
 sg13g2_mux4_1 _15366_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .S1(net918),
    .X(_08627_));
 sg13g2_buf_2 _15367_ (.A(net919),
    .X(_08628_));
 sg13g2_buf_1 _15368_ (.A(_08545_),
    .X(_08629_));
 sg13g2_buf_1 _15369_ (.A(net1054),
    .X(_08630_));
 sg13g2_mux4_1 _15370_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .S1(net917),
    .X(_08631_));
 sg13g2_mux4_1 _15371_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .S1(net917),
    .X(_08632_));
 sg13g2_buf_2 _15372_ (.A(_08559_),
    .X(_08633_));
 sg13g2_buf_1 _15373_ (.A(net1061),
    .X(_08634_));
 sg13g2_mux4_1 _15374_ (.S0(net916),
    .A0(_08626_),
    .A1(_08627_),
    .A2(_08631_),
    .A3(_08632_),
    .S1(net915),
    .X(_08635_));
 sg13g2_nand2_1 _15375_ (.Y(_08636_),
    .A(net920),
    .B(_08635_));
 sg13g2_mux4_1 _15376_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .S1(net918),
    .X(_08637_));
 sg13g2_mux4_1 _15377_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .S1(net918),
    .X(_08638_));
 sg13g2_buf_2 _15378_ (.A(net919),
    .X(_08639_));
 sg13g2_buf_1 _15379_ (.A(net1054),
    .X(_08640_));
 sg13g2_mux4_1 _15380_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .S1(_08640_),
    .X(_08641_));
 sg13g2_mux4_1 _15381_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .S1(net914),
    .X(_08642_));
 sg13g2_buf_1 _15382_ (.A(net1061),
    .X(_08643_));
 sg13g2_mux4_1 _15383_ (.S0(net916),
    .A0(_08637_),
    .A1(_08638_),
    .A2(_08641_),
    .A3(_08642_),
    .S1(net913),
    .X(_08644_));
 sg13g2_nand2b_1 _15384_ (.Y(_08645_),
    .B(_08644_),
    .A_N(_08620_));
 sg13g2_nand3_1 _15385_ (.B(_08636_),
    .C(_08645_),
    .A(net1057),
    .Y(_08646_));
 sg13g2_o21ai_1 _15386_ (.B1(_08646_),
    .Y(_08647_),
    .A1(net790),
    .A2(net1057));
 sg13g2_buf_2 _15387_ (.A(_08647_),
    .X(_08648_));
 sg13g2_buf_1 _15388_ (.A(net554),
    .X(_08649_));
 sg13g2_buf_1 _15389_ (.A(_08321_),
    .X(_08650_));
 sg13g2_buf_1 _15390_ (.A(net699),
    .X(_08651_));
 sg13g2_a22oi_1 _15391_ (.Y(_08652_),
    .B1(net633),
    .B2(\cpu.icache.r_tag[4][12] ),
    .A2(net548),
    .A1(\cpu.icache.r_tag[1][12] ));
 sg13g2_buf_1 _15392_ (.A(net640),
    .X(_08653_));
 sg13g2_buf_2 _15393_ (.A(net551),
    .X(_08654_));
 sg13g2_buf_1 _15394_ (.A(net481),
    .X(_08655_));
 sg13g2_a22oi_1 _15395_ (.Y(_08656_),
    .B1(net425),
    .B2(\cpu.icache.r_tag[3][12] ),
    .A2(net547),
    .A1(\cpu.icache.r_tag[2][12] ));
 sg13g2_buf_1 _15396_ (.A(net927),
    .X(_08657_));
 sg13g2_mux2_1 _15397_ (.A0(\cpu.icache.r_tag[5][12] ),
    .A1(\cpu.icache.r_tag[7][12] ),
    .S(net793),
    .X(_08658_));
 sg13g2_nor2b_1 _15398_ (.A(net1070),
    .B_N(net1069),
    .Y(_08659_));
 sg13g2_buf_2 _15399_ (.A(_08659_),
    .X(_08660_));
 sg13g2_a22oi_1 _15400_ (.Y(_08661_),
    .B1(_08660_),
    .B2(\cpu.icache.r_tag[6][12] ),
    .A2(_08658_),
    .A1(net792));
 sg13g2_or2_1 _15401_ (.X(_08662_),
    .B(_08661_),
    .A(net786));
 sg13g2_nand4_1 _15402_ (.B(_08652_),
    .C(_08656_),
    .A(net482),
    .Y(_08663_),
    .D(_08662_));
 sg13g2_o21ai_1 _15403_ (.B1(_08663_),
    .Y(_08664_),
    .A1(\cpu.icache.r_tag[0][12] ),
    .A2(net482));
 sg13g2_xor2_1 _15404_ (.B(_08664_),
    .A(net384),
    .X(_08665_));
 sg13g2_buf_1 _15405_ (.A(net1055),
    .X(_08666_));
 sg13g2_mux4_1 _15406_ (.S0(_08623_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .S1(_08625_),
    .X(_08667_));
 sg13g2_mux4_1 _15407_ (.S0(_08623_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .S1(_08625_),
    .X(_08668_));
 sg13g2_mux4_1 _15408_ (.S0(_08628_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .S1(_08630_),
    .X(_08669_));
 sg13g2_mux4_1 _15409_ (.S0(_08628_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .S1(_08630_),
    .X(_08670_));
 sg13g2_mux4_1 _15410_ (.S0(net916),
    .A0(_08667_),
    .A1(_08668_),
    .A2(_08669_),
    .A3(_08670_),
    .S1(net915),
    .X(_08671_));
 sg13g2_nand2_1 _15411_ (.Y(_08672_),
    .A(net920),
    .B(_08671_));
 sg13g2_mux4_1 _15412_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .S1(net918),
    .X(_08673_));
 sg13g2_mux4_1 _15413_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .S1(net918),
    .X(_08674_));
 sg13g2_mux4_1 _15414_ (.S0(_08639_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .S1(_08640_),
    .X(_08675_));
 sg13g2_mux4_1 _15415_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .S1(net917),
    .X(_08676_));
 sg13g2_mux4_1 _15416_ (.S0(net916),
    .A0(_08673_),
    .A1(_08674_),
    .A2(_08675_),
    .A3(_08676_),
    .S1(net915),
    .X(_08677_));
 sg13g2_nand2b_1 _15417_ (.Y(_08678_),
    .B(_08677_),
    .A_N(net920));
 sg13g2_nand3_1 _15418_ (.B(_08672_),
    .C(_08678_),
    .A(net1057),
    .Y(_08679_));
 sg13g2_o21ai_1 _15419_ (.B1(_08679_),
    .Y(_08680_),
    .A1(net912),
    .A2(net1057));
 sg13g2_buf_2 _15420_ (.A(_08680_),
    .X(_08681_));
 sg13g2_buf_1 _15421_ (.A(net635),
    .X(_08682_));
 sg13g2_buf_2 _15422_ (.A(net633),
    .X(_08683_));
 sg13g2_a22oi_1 _15423_ (.Y(_08684_),
    .B1(_08683_),
    .B2(\cpu.icache.r_tag[4][13] ),
    .A2(_08682_),
    .A1(\cpu.icache.r_tag[1][13] ));
 sg13g2_buf_1 _15424_ (.A(net556),
    .X(_08685_));
 sg13g2_a22oi_1 _15425_ (.Y(_08686_),
    .B1(_08655_),
    .B2(\cpu.icache.r_tag[3][13] ),
    .A2(_08685_),
    .A1(\cpu.icache.r_tag[2][13] ));
 sg13g2_mux2_1 _15426_ (.A0(\cpu.icache.r_tag[5][13] ),
    .A1(\cpu.icache.r_tag[7][13] ),
    .S(_08337_),
    .X(_08687_));
 sg13g2_a22oi_1 _15427_ (.Y(_08688_),
    .B1(_08687_),
    .B2(net701),
    .A2(_08660_),
    .A1(\cpu.icache.r_tag[6][13] ));
 sg13g2_or2_1 _15428_ (.X(_08689_),
    .B(_08688_),
    .A(net786));
 sg13g2_nand4_1 _15429_ (.B(_08684_),
    .C(_08686_),
    .A(net482),
    .Y(_08690_),
    .D(_08689_));
 sg13g2_o21ai_1 _15430_ (.B1(_08690_),
    .Y(_08691_),
    .A1(\cpu.icache.r_tag[0][13] ),
    .A2(net482));
 sg13g2_xor2_1 _15431_ (.B(_08691_),
    .A(net383),
    .X(_08692_));
 sg13g2_nor2_1 _15432_ (.A(_08665_),
    .B(_08692_),
    .Y(_08693_));
 sg13g2_buf_2 _15433_ (.A(_00192_),
    .X(_08694_));
 sg13g2_buf_1 _15434_ (.A(_08694_),
    .X(_08695_));
 sg13g2_buf_2 _15435_ (.A(_08547_),
    .X(_08696_));
 sg13g2_buf_1 _15436_ (.A(net1054),
    .X(_08697_));
 sg13g2_mux4_1 _15437_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S1(net910),
    .X(_08698_));
 sg13g2_mux4_1 _15438_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S1(net910),
    .X(_08699_));
 sg13g2_buf_2 _15439_ (.A(_08547_),
    .X(_08700_));
 sg13g2_mux4_1 _15440_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S1(net910),
    .X(_08701_));
 sg13g2_mux4_1 _15441_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S1(net910),
    .X(_08702_));
 sg13g2_buf_2 _15442_ (.A(_08559_),
    .X(_08703_));
 sg13g2_mux4_1 _15443_ (.S0(net908),
    .A0(_08698_),
    .A1(_08699_),
    .A2(_08701_),
    .A3(_08702_),
    .S1(_08643_),
    .X(_08704_));
 sg13g2_mux4_1 _15444_ (.S0(_08696_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S1(_08697_),
    .X(_08705_));
 sg13g2_mux4_1 _15445_ (.S0(_08696_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S1(_08697_),
    .X(_08706_));
 sg13g2_buf_1 _15446_ (.A(_08545_),
    .X(_08707_));
 sg13g2_mux4_1 _15447_ (.S0(_08700_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S1(net1052),
    .X(_08708_));
 sg13g2_mux4_1 _15448_ (.S0(_08700_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S1(_08707_),
    .X(_08709_));
 sg13g2_mux4_1 _15449_ (.S0(_08703_),
    .A0(_08705_),
    .A1(_08706_),
    .A2(_08708_),
    .A3(_08709_),
    .S1(_08643_),
    .X(_08710_));
 sg13g2_mux2_1 _15450_ (.A0(_08704_),
    .A1(_08710_),
    .S(net1056),
    .X(_08711_));
 sg13g2_nand2b_1 _15451_ (.Y(_08712_),
    .B(_08711_),
    .A_N(net1053));
 sg13g2_buf_1 _15452_ (.A(_08712_),
    .X(_08713_));
 sg13g2_mux4_1 _15453_ (.S0(net791),
    .A0(\cpu.icache.r_tag[4][20] ),
    .A1(\cpu.icache.r_tag[5][20] ),
    .A2(\cpu.icache.r_tag[6][20] ),
    .A3(\cpu.icache.r_tag[7][20] ),
    .S1(_08337_),
    .X(_08714_));
 sg13g2_nand2b_1 _15454_ (.Y(_08715_),
    .B(_08714_),
    .A_N(_08657_));
 sg13g2_nand2_1 _15455_ (.Y(_08716_),
    .A(\cpu.icache.r_tag[1][20] ),
    .B(net548));
 sg13g2_a22oi_1 _15456_ (.Y(_08717_),
    .B1(net481),
    .B2(\cpu.icache.r_tag[3][20] ),
    .A2(net556),
    .A1(\cpu.icache.r_tag[2][20] ));
 sg13g2_nand4_1 _15457_ (.B(_08715_),
    .C(_08716_),
    .A(net554),
    .Y(_08718_),
    .D(_08717_));
 sg13g2_o21ai_1 _15458_ (.B1(_08718_),
    .Y(_08719_),
    .A1(\cpu.icache.r_tag[0][20] ),
    .A2(net482));
 sg13g2_xnor2_1 _15459_ (.Y(_08720_),
    .A(net479),
    .B(_08719_));
 sg13g2_buf_2 _15460_ (.A(net921),
    .X(_08721_));
 sg13g2_buf_1 _15461_ (.A(net1055),
    .X(_08722_));
 sg13g2_mux4_1 _15462_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S1(net907),
    .X(_08723_));
 sg13g2_mux4_1 _15463_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S1(net907),
    .X(_08724_));
 sg13g2_mux4_1 _15464_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S1(net907),
    .X(_08725_));
 sg13g2_mux4_1 _15465_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S1(net907),
    .X(_08726_));
 sg13g2_mux4_1 _15466_ (.S0(net916),
    .A0(_08723_),
    .A1(_08724_),
    .A2(_08725_),
    .A3(_08726_),
    .S1(net915),
    .X(_08727_));
 sg13g2_mux4_1 _15467_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S1(net907),
    .X(_08728_));
 sg13g2_mux4_1 _15468_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S1(net907),
    .X(_08729_));
 sg13g2_mux4_1 _15469_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S1(net918),
    .X(_08730_));
 sg13g2_mux4_1 _15470_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S1(net918),
    .X(_08731_));
 sg13g2_mux4_1 _15471_ (.S0(net916),
    .A0(_08728_),
    .A1(_08729_),
    .A2(_08730_),
    .A3(_08731_),
    .S1(net915),
    .X(_08732_));
 sg13g2_mux2_1 _15472_ (.A0(_08727_),
    .A1(_08732_),
    .S(net920),
    .X(_08733_));
 sg13g2_nand2b_1 _15473_ (.Y(_08734_),
    .B(_08733_),
    .A_N(net1053));
 sg13g2_buf_2 _15474_ (.A(_08734_),
    .X(_08735_));
 sg13g2_buf_1 _15475_ (.A(net549),
    .X(_08736_));
 sg13g2_a22oi_1 _15476_ (.Y(_08737_),
    .B1(net633),
    .B2(\cpu.icache.r_tag[4][19] ),
    .A2(net548),
    .A1(\cpu.icache.r_tag[1][19] ));
 sg13g2_a22oi_1 _15477_ (.Y(_08738_),
    .B1(net481),
    .B2(\cpu.icache.r_tag[3][19] ),
    .A2(net547),
    .A1(\cpu.icache.r_tag[2][19] ));
 sg13g2_mux2_1 _15478_ (.A0(\cpu.icache.r_tag[5][19] ),
    .A1(\cpu.icache.r_tag[7][19] ),
    .S(net797),
    .X(_08739_));
 sg13g2_a22oi_1 _15479_ (.Y(_08740_),
    .B1(_08739_),
    .B2(net792),
    .A2(_08660_),
    .A1(\cpu.icache.r_tag[6][19] ));
 sg13g2_or2_1 _15480_ (.X(_08741_),
    .B(_08740_),
    .A(net786));
 sg13g2_nand4_1 _15481_ (.B(_08737_),
    .C(_08738_),
    .A(net478),
    .Y(_08742_),
    .D(_08741_));
 sg13g2_o21ai_1 _15482_ (.B1(_08742_),
    .Y(_08743_),
    .A1(\cpu.icache.r_tag[0][19] ),
    .A2(_08649_));
 sg13g2_xor2_1 _15483_ (.B(_08743_),
    .A(net424),
    .X(_08744_));
 sg13g2_inv_1 _15484_ (.Y(_08745_),
    .A(_08744_));
 sg13g2_mux4_1 _15485_ (.S0(net921),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .S1(net1055),
    .X(_08746_));
 sg13g2_mux4_1 _15486_ (.S0(_08617_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .S1(_08624_),
    .X(_08747_));
 sg13g2_mux4_1 _15487_ (.S0(net919),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .S1(net1054),
    .X(_08748_));
 sg13g2_mux4_1 _15488_ (.S0(net919),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .S1(net1054),
    .X(_08749_));
 sg13g2_mux4_1 _15489_ (.S0(_08559_),
    .A0(_08746_),
    .A1(_08747_),
    .A2(_08748_),
    .A3(_08749_),
    .S1(net1061),
    .X(_08750_));
 sg13g2_mux4_1 _15490_ (.S0(net919),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .S1(net1054),
    .X(_08751_));
 sg13g2_mux4_1 _15491_ (.S0(net919),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .S1(_08624_),
    .X(_08752_));
 sg13g2_mux4_1 _15492_ (.S0(net919),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .S1(net1054),
    .X(_08753_));
 sg13g2_mux4_1 _15493_ (.S0(_08622_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .S1(_08629_),
    .X(_08754_));
 sg13g2_mux4_1 _15494_ (.S0(_08559_),
    .A0(_08751_),
    .A1(_08752_),
    .A2(_08753_),
    .A3(_08754_),
    .S1(net1061),
    .X(_08755_));
 sg13g2_mux2_1 _15495_ (.A0(_08750_),
    .A1(_08755_),
    .S(net1056),
    .X(_08756_));
 sg13g2_nand2b_1 _15496_ (.Y(_08757_),
    .B(_08756_),
    .A_N(net1053));
 sg13g2_buf_2 _15497_ (.A(_08757_),
    .X(_08758_));
 sg13g2_nand2_1 _15498_ (.Y(_08759_),
    .A(\cpu.icache.r_tag[1][23] ),
    .B(net548));
 sg13g2_a22oi_1 _15499_ (.Y(_08760_),
    .B1(net639),
    .B2(\cpu.icache.r_tag[6][23] ),
    .A2(net633),
    .A1(\cpu.icache.r_tag[4][23] ));
 sg13g2_and2_1 _15500_ (.A(net931),
    .B(net1068),
    .X(_08761_));
 sg13g2_a22oi_1 _15501_ (.Y(_08762_),
    .B1(_08761_),
    .B2(\cpu.icache.r_tag[3][23] ),
    .A2(net929),
    .A1(\cpu.icache.r_tag[5][23] ));
 sg13g2_nor2_1 _15502_ (.A(net930),
    .B(_08762_),
    .Y(_08763_));
 sg13g2_a221oi_1 _15503_ (.B2(\cpu.icache.r_tag[7][23] ),
    .C1(_08763_),
    .B1(_08305_),
    .A1(\cpu.icache.r_tag[2][23] ),
    .Y(_08764_),
    .A2(net556));
 sg13g2_nand4_1 _15504_ (.B(_08759_),
    .C(_08760_),
    .A(net478),
    .Y(_08765_),
    .D(_08764_));
 sg13g2_o21ai_1 _15505_ (.B1(_08765_),
    .Y(_08766_),
    .A1(\cpu.icache.r_tag[0][23] ),
    .A2(_08649_));
 sg13g2_xor2_1 _15506_ (.B(_08766_),
    .A(net477),
    .X(_08767_));
 sg13g2_inv_1 _15507_ (.Y(_08768_),
    .A(\cpu.ex.pc[11] ));
 sg13g2_buf_1 _15508_ (.A(_08768_),
    .X(_08769_));
 sg13g2_a22oi_1 _15509_ (.Y(_08770_),
    .B1(net638),
    .B2(\cpu.icache.r_tag[5][11] ),
    .A2(_08326_),
    .A1(\cpu.icache.r_tag[6][11] ));
 sg13g2_mux2_1 _15510_ (.A0(\cpu.icache.r_tag[7][11] ),
    .A1(\cpu.icache.r_tag[3][11] ),
    .S(net1068),
    .X(_08771_));
 sg13g2_a22oi_1 _15511_ (.Y(_08772_),
    .B1(_08297_),
    .B2(_08771_),
    .A2(net796),
    .A1(\cpu.icache.r_tag[4][11] ));
 sg13g2_a22oi_1 _15512_ (.Y(_08773_),
    .B1(_08322_),
    .B2(\cpu.icache.r_tag[2][11] ),
    .A2(net700),
    .A1(\cpu.icache.r_tag[1][11] ));
 sg13g2_nand4_1 _15513_ (.B(_08770_),
    .C(_08772_),
    .A(_08364_),
    .Y(_08774_),
    .D(_08773_));
 sg13g2_o21ai_1 _15514_ (.B1(_08774_),
    .Y(_08775_),
    .A1(\cpu.icache.r_tag[0][11] ),
    .A2(net549));
 sg13g2_xnor2_1 _15515_ (.Y(_08776_),
    .A(net1051),
    .B(_08775_));
 sg13g2_buf_2 _15516_ (.A(\cpu.ex.pc[6] ),
    .X(_08777_));
 sg13g2_a22oi_1 _15517_ (.Y(_08778_),
    .B1(_08328_),
    .B2(\cpu.icache.r_tag[5][6] ),
    .A2(net551),
    .A1(\cpu.icache.r_tag[3][6] ));
 sg13g2_a22oi_1 _15518_ (.Y(_08779_),
    .B1(_08305_),
    .B2(\cpu.icache.r_tag[7][6] ),
    .A2(net636),
    .A1(\cpu.icache.r_tag[2][6] ));
 sg13g2_buf_1 _15519_ (.A(net795),
    .X(_08780_));
 sg13g2_mux2_1 _15520_ (.A0(\cpu.icache.r_tag[4][6] ),
    .A1(\cpu.icache.r_tag[6][6] ),
    .S(_08275_),
    .X(_08781_));
 sg13g2_a22oi_1 _15521_ (.Y(_08782_),
    .B1(net697),
    .B2(_08781_),
    .A2(net703),
    .A1(\cpu.icache.r_tag[1][6] ));
 sg13g2_nand4_1 _15522_ (.B(_08778_),
    .C(_08779_),
    .A(net637),
    .Y(_08783_),
    .D(_08782_));
 sg13g2_o21ai_1 _15523_ (.B1(_08783_),
    .Y(_08784_),
    .A1(\cpu.icache.r_tag[0][6] ),
    .A2(net549));
 sg13g2_xor2_1 _15524_ (.B(_08784_),
    .A(_08777_),
    .X(_08785_));
 sg13g2_buf_2 _15525_ (.A(\cpu.ex.pc[9] ),
    .X(_08786_));
 sg13g2_inv_1 _15526_ (.Y(_08787_),
    .A(_08786_));
 sg13g2_buf_1 _15527_ (.A(_08787_),
    .X(_08788_));
 sg13g2_a22oi_1 _15528_ (.Y(_08789_),
    .B1(_08326_),
    .B2(\cpu.icache.r_tag[6][9] ),
    .A2(_08322_),
    .A1(\cpu.icache.r_tag[2][9] ));
 sg13g2_a22oi_1 _15529_ (.Y(_08790_),
    .B1(_08370_),
    .B2(\cpu.icache.r_tag[4][9] ),
    .A2(_08355_),
    .A1(\cpu.icache.r_tag[1][9] ));
 sg13g2_mux2_1 _15530_ (.A0(\cpu.icache.r_tag[7][9] ),
    .A1(\cpu.icache.r_tag[3][9] ),
    .S(_08261_),
    .X(_08791_));
 sg13g2_a22oi_1 _15531_ (.Y(_08792_),
    .B1(_08791_),
    .B2(net797),
    .A2(net929),
    .A1(\cpu.icache.r_tag[5][9] ));
 sg13g2_nand2b_1 _15532_ (.Y(_08793_),
    .B(net791),
    .A_N(_08792_));
 sg13g2_nand4_1 _15533_ (.B(_08789_),
    .C(_08790_),
    .A(_08364_),
    .Y(_08794_),
    .D(_08793_));
 sg13g2_o21ai_1 _15534_ (.B1(_08794_),
    .Y(_08795_),
    .A1(\cpu.icache.r_tag[0][9] ),
    .A2(net549));
 sg13g2_xnor2_1 _15535_ (.Y(_08796_),
    .A(net906),
    .B(_08795_));
 sg13g2_buf_1 _15536_ (.A(\cpu.ex.pc[7] ),
    .X(_08797_));
 sg13g2_a22oi_1 _15537_ (.Y(_08798_),
    .B1(net699),
    .B2(\cpu.icache.r_tag[4][7] ),
    .A2(net703),
    .A1(\cpu.icache.r_tag[1][7] ));
 sg13g2_a22oi_1 _15538_ (.Y(_08799_),
    .B1(net551),
    .B2(\cpu.icache.r_tag[3][7] ),
    .A2(net636),
    .A1(\cpu.icache.r_tag[2][7] ));
 sg13g2_mux2_1 _15539_ (.A0(\cpu.icache.r_tag[5][7] ),
    .A1(\cpu.icache.r_tag[7][7] ),
    .S(net1069),
    .X(_08800_));
 sg13g2_a22oi_1 _15540_ (.Y(_08801_),
    .B1(_08800_),
    .B2(net925),
    .A2(_08660_),
    .A1(\cpu.icache.r_tag[6][7] ));
 sg13g2_or2_1 _15541_ (.X(_08802_),
    .B(_08801_),
    .A(net924));
 sg13g2_nand4_1 _15542_ (.B(_08798_),
    .C(_08799_),
    .A(net637),
    .Y(_08803_),
    .D(_08802_));
 sg13g2_o21ai_1 _15543_ (.B1(_08803_),
    .Y(_08804_),
    .A1(\cpu.icache.r_tag[0][7] ),
    .A2(_08392_));
 sg13g2_xor2_1 _15544_ (.B(_08804_),
    .A(_08797_),
    .X(_08805_));
 sg13g2_nand4_1 _15545_ (.B(_08785_),
    .C(_08796_),
    .A(_08776_),
    .Y(_08806_),
    .D(_08805_));
 sg13g2_buf_1 _15546_ (.A(\cpu.ex.pc[10] ),
    .X(_08807_));
 sg13g2_a22oi_1 _15547_ (.Y(_08808_),
    .B1(_08305_),
    .B2(\cpu.icache.r_tag[7][10] ),
    .A2(_08326_),
    .A1(\cpu.icache.r_tag[6][10] ));
 sg13g2_and2_1 _15548_ (.A(\cpu.icache.r_tag[4][10] ),
    .B(_08290_),
    .X(_08809_));
 sg13g2_a221oi_1 _15549_ (.B2(\cpu.icache.r_tag[5][10] ),
    .C1(_08809_),
    .B1(_08285_),
    .A1(\cpu.icache.r_tag[2][10] ),
    .Y(_08810_),
    .A2(net636));
 sg13g2_a22oi_1 _15550_ (.Y(_08811_),
    .B1(_08357_),
    .B2(\cpu.icache.r_tag[3][10] ),
    .A2(net703),
    .A1(\cpu.icache.r_tag[1][10] ));
 sg13g2_nand4_1 _15551_ (.B(_08808_),
    .C(_08810_),
    .A(net637),
    .Y(_08812_),
    .D(_08811_));
 sg13g2_o21ai_1 _15552_ (.B1(_08812_),
    .Y(_08813_),
    .A1(\cpu.icache.r_tag[0][10] ),
    .A2(_08392_));
 sg13g2_xor2_1 _15553_ (.B(_08813_),
    .A(_08807_),
    .X(_08814_));
 sg13g2_mux4_1 _15554_ (.S0(net792),
    .A0(\cpu.icache.r_valid[4] ),
    .A1(\cpu.icache.r_valid[5] ),
    .A2(\cpu.icache.r_valid[6] ),
    .A3(\cpu.icache.r_valid[7] ),
    .S1(net702),
    .X(_08815_));
 sg13g2_mux4_1 _15555_ (.S0(net792),
    .A0(\cpu.icache.r_valid[0] ),
    .A1(\cpu.icache.r_valid[1] ),
    .A2(\cpu.icache.r_valid[2] ),
    .A3(\cpu.icache.r_valid[3] ),
    .S1(net698),
    .X(_08816_));
 sg13g2_inv_2 _15556_ (.Y(_08817_),
    .A(_08264_));
 sg13g2_mux2_1 _15557_ (.A0(_08815_),
    .A1(_08816_),
    .S(_08817_),
    .X(_08818_));
 sg13g2_inv_1 _15558_ (.Y(_08819_),
    .A(\cpu.ex.pc[8] ));
 sg13g2_buf_1 _15559_ (.A(_08819_),
    .X(_08820_));
 sg13g2_a22oi_1 _15560_ (.Y(_08821_),
    .B1(_08326_),
    .B2(\cpu.icache.r_tag[6][8] ),
    .A2(_08347_),
    .A1(\cpu.icache.r_tag[2][8] ));
 sg13g2_a22oi_1 _15561_ (.Y(_08822_),
    .B1(_08290_),
    .B2(\cpu.icache.r_tag[4][8] ),
    .A2(_08320_),
    .A1(\cpu.icache.r_tag[1][8] ));
 sg13g2_mux2_1 _15562_ (.A0(\cpu.icache.r_tag[7][8] ),
    .A1(\cpu.icache.r_tag[3][8] ),
    .S(_08261_),
    .X(_08823_));
 sg13g2_a22oi_1 _15563_ (.Y(_08824_),
    .B1(_08823_),
    .B2(_08275_),
    .A2(net929),
    .A1(\cpu.icache.r_tag[5][8] ));
 sg13g2_nand2b_1 _15564_ (.Y(_08825_),
    .B(net791),
    .A_N(_08824_));
 sg13g2_nand4_1 _15565_ (.B(_08821_),
    .C(_08822_),
    .A(_08332_),
    .Y(_08826_),
    .D(_08825_));
 sg13g2_o21ai_1 _15566_ (.B1(_08826_),
    .Y(_08827_),
    .A1(\cpu.icache.r_tag[0][8] ),
    .A2(net550));
 sg13g2_xnor2_1 _15567_ (.Y(_08828_),
    .A(net1050),
    .B(_08827_));
 sg13g2_buf_2 _15568_ (.A(\cpu.ex.pc[5] ),
    .X(_08829_));
 sg13g2_a22oi_1 _15569_ (.Y(_08830_),
    .B1(_08328_),
    .B2(\cpu.icache.r_tag[5][5] ),
    .A2(_08320_),
    .A1(\cpu.icache.r_tag[1][5] ));
 sg13g2_a22oi_1 _15570_ (.Y(_08831_),
    .B1(_08357_),
    .B2(\cpu.icache.r_tag[3][5] ),
    .A2(_08347_),
    .A1(\cpu.icache.r_tag[2][5] ));
 sg13g2_mux2_1 _15571_ (.A0(\cpu.icache.r_tag[4][5] ),
    .A1(\cpu.icache.r_tag[6][5] ),
    .S(_08267_),
    .X(_08832_));
 sg13g2_a22oi_1 _15572_ (.Y(_08833_),
    .B1(_08832_),
    .B2(net930),
    .A2(_08297_),
    .A1(\cpu.icache.r_tag[7][5] ));
 sg13g2_or2_1 _15573_ (.X(_08834_),
    .B(_08833_),
    .A(net924));
 sg13g2_nand4_1 _15574_ (.B(_08830_),
    .C(_08831_),
    .A(net637),
    .Y(_08835_),
    .D(_08834_));
 sg13g2_o21ai_1 _15575_ (.B1(_08835_),
    .Y(_08836_),
    .A1(\cpu.icache.r_tag[0][5] ),
    .A2(net550));
 sg13g2_xor2_1 _15576_ (.B(_08836_),
    .A(_08829_),
    .X(_08837_));
 sg13g2_nand4_1 _15577_ (.B(_08818_),
    .C(_08828_),
    .A(_08814_),
    .Y(_08838_),
    .D(_08837_));
 sg13g2_nor3_1 _15578_ (.A(_08767_),
    .B(_08806_),
    .C(_08838_),
    .Y(_08839_));
 sg13g2_nand4_1 _15579_ (.B(_08720_),
    .C(_08745_),
    .A(_08693_),
    .Y(_08840_),
    .D(_08839_));
 sg13g2_mux4_1 _15580_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S1(net917),
    .X(_08841_));
 sg13g2_mux4_1 _15581_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S1(net917),
    .X(_08842_));
 sg13g2_buf_2 _15582_ (.A(_08547_),
    .X(_08843_));
 sg13g2_buf_1 _15583_ (.A(net1054),
    .X(_08844_));
 sg13g2_mux4_1 _15584_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S1(net904),
    .X(_08845_));
 sg13g2_mux4_1 _15585_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S1(net914),
    .X(_08846_));
 sg13g2_mux4_1 _15586_ (.S0(net916),
    .A0(_08841_),
    .A1(_08842_),
    .A2(_08845_),
    .A3(_08846_),
    .S1(net913),
    .X(_08847_));
 sg13g2_mux4_1 _15587_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S1(net914),
    .X(_08848_));
 sg13g2_mux4_1 _15588_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S1(net917),
    .X(_08849_));
 sg13g2_mux4_1 _15589_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S1(net904),
    .X(_08850_));
 sg13g2_mux4_1 _15590_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S1(net904),
    .X(_08851_));
 sg13g2_mux4_1 _15591_ (.S0(net908),
    .A0(_08848_),
    .A1(_08849_),
    .A2(_08850_),
    .A3(_08851_),
    .S1(net913),
    .X(_08852_));
 sg13g2_mux2_1 _15592_ (.A0(_08847_),
    .A1(_08852_),
    .S(net1056),
    .X(_08853_));
 sg13g2_nand2b_1 _15593_ (.Y(_08854_),
    .B(_08853_),
    .A_N(net1053));
 sg13g2_buf_2 _15594_ (.A(_08854_),
    .X(_08855_));
 sg13g2_mux2_1 _15595_ (.A0(\cpu.icache.r_tag[7][18] ),
    .A1(\cpu.icache.r_tag[3][18] ),
    .S(_08317_),
    .X(_08856_));
 sg13g2_a22oi_1 _15596_ (.Y(_08857_),
    .B1(net704),
    .B2(_08856_),
    .A2(net633),
    .A1(\cpu.icache.r_tag[4][18] ));
 sg13g2_a22oi_1 _15597_ (.Y(_08858_),
    .B1(net555),
    .B2(\cpu.icache.r_tag[5][18] ),
    .A2(net548),
    .A1(\cpu.icache.r_tag[1][18] ));
 sg13g2_a22oi_1 _15598_ (.Y(_08859_),
    .B1(net639),
    .B2(\cpu.icache.r_tag[6][18] ),
    .A2(net547),
    .A1(\cpu.icache.r_tag[2][18] ));
 sg13g2_nand3_1 _15599_ (.B(_08858_),
    .C(_08859_),
    .A(_08857_),
    .Y(_08860_));
 sg13g2_mux2_1 _15600_ (.A0(\cpu.icache.r_tag[0][18] ),
    .A1(_08860_),
    .S(net478),
    .X(_08861_));
 sg13g2_xor2_1 _15601_ (.B(_08861_),
    .A(_08855_),
    .X(_08862_));
 sg13g2_mux4_1 _15602_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S1(net1052),
    .X(_08863_));
 sg13g2_mux4_1 _15603_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S1(net1052),
    .X(_08864_));
 sg13g2_buf_2 _15604_ (.A(_08547_),
    .X(_08865_));
 sg13g2_buf_1 _15605_ (.A(_08545_),
    .X(_08866_));
 sg13g2_mux4_1 _15606_ (.S0(net903),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S1(net1049),
    .X(_08867_));
 sg13g2_mux4_1 _15607_ (.S0(net903),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S1(net1049),
    .X(_08868_));
 sg13g2_mux4_1 _15608_ (.S0(_08538_),
    .A0(_08863_),
    .A1(_08864_),
    .A2(_08867_),
    .A3(_08868_),
    .S1(net1127),
    .X(_08869_));
 sg13g2_a21oi_1 _15609_ (.A1(net1057),
    .A2(_08869_),
    .Y(_08870_),
    .B1(net915));
 sg13g2_inv_1 _15610_ (.Y(_08871_),
    .A(net1061));
 sg13g2_mux4_1 _15611_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S1(net910),
    .X(_08872_));
 sg13g2_mux4_1 _15612_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S1(net910),
    .X(_08873_));
 sg13g2_mux4_1 _15613_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S1(net1052),
    .X(_08874_));
 sg13g2_mux4_1 _15614_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S1(net1052),
    .X(_08875_));
 sg13g2_mux4_1 _15615_ (.S0(_08538_),
    .A0(_08872_),
    .A1(_08873_),
    .A2(_08874_),
    .A3(_08875_),
    .S1(net1056),
    .X(_08876_));
 sg13g2_nor3_1 _15616_ (.A(_08871_),
    .B(_08464_),
    .C(_08876_),
    .Y(_08877_));
 sg13g2_or2_1 _15617_ (.X(_08878_),
    .B(_08877_),
    .A(_08870_));
 sg13g2_buf_2 _15618_ (.A(_08878_),
    .X(_08879_));
 sg13g2_a22oi_1 _15619_ (.Y(_08880_),
    .B1(net555),
    .B2(\cpu.icache.r_tag[5][14] ),
    .A2(net705),
    .A1(\cpu.icache.r_tag[4][14] ));
 sg13g2_a22oi_1 _15620_ (.Y(_08881_),
    .B1(_08323_),
    .B2(\cpu.icache.r_tag[2][14] ),
    .A2(net635),
    .A1(\cpu.icache.r_tag[1][14] ));
 sg13g2_mux2_1 _15621_ (.A0(\cpu.icache.r_tag[7][14] ),
    .A1(\cpu.icache.r_tag[3][14] ),
    .S(net924),
    .X(_08882_));
 sg13g2_a22oi_1 _15622_ (.Y(_08883_),
    .B1(_08882_),
    .B2(net792),
    .A2(_08780_),
    .A1(\cpu.icache.r_tag[6][14] ));
 sg13g2_nand2b_1 _15623_ (.Y(_08884_),
    .B(net702),
    .A_N(_08883_));
 sg13g2_nand4_1 _15624_ (.B(_08880_),
    .C(_08881_),
    .A(net554),
    .Y(_08885_),
    .D(_08884_));
 sg13g2_o21ai_1 _15625_ (.B1(_08885_),
    .Y(_08886_),
    .A1(\cpu.icache.r_tag[0][14] ),
    .A2(net478));
 sg13g2_xnor2_1 _15626_ (.Y(_08887_),
    .A(net476),
    .B(_08886_));
 sg13g2_mux4_1 _15627_ (.S0(net903),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S1(net1049),
    .X(_08888_));
 sg13g2_mux4_1 _15628_ (.S0(net903),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S1(net1049),
    .X(_08889_));
 sg13g2_mux4_1 _15629_ (.S0(net921),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S1(net1055),
    .X(_08890_));
 sg13g2_mux4_1 _15630_ (.S0(net921),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S1(net1055),
    .X(_08891_));
 sg13g2_mux4_1 _15631_ (.S0(net908),
    .A0(_08888_),
    .A1(_08889_),
    .A2(_08890_),
    .A3(_08891_),
    .S1(net913),
    .X(_08892_));
 sg13g2_mux4_1 _15632_ (.S0(net903),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S1(net1049),
    .X(_08893_));
 sg13g2_mux4_1 _15633_ (.S0(net903),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S1(net1049),
    .X(_08894_));
 sg13g2_mux4_1 _15634_ (.S0(net921),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S1(net1055),
    .X(_08895_));
 sg13g2_mux4_1 _15635_ (.S0(net921),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S1(net1055),
    .X(_08896_));
 sg13g2_mux4_1 _15636_ (.S0(net908),
    .A0(_08893_),
    .A1(_08894_),
    .A2(_08895_),
    .A3(_08896_),
    .S1(net1061),
    .X(_08897_));
 sg13g2_mux2_1 _15637_ (.A0(_08892_),
    .A1(_08897_),
    .S(net1056),
    .X(_08898_));
 sg13g2_nand2b_1 _15638_ (.Y(_08899_),
    .B(_08898_),
    .A_N(net1053));
 sg13g2_buf_2 _15639_ (.A(_08899_),
    .X(_08900_));
 sg13g2_and2_1 _15640_ (.A(\cpu.icache.r_tag[4][17] ),
    .B(net699),
    .X(_08901_));
 sg13g2_a221oi_1 _15641_ (.B2(\cpu.icache.r_tag[5][17] ),
    .C1(_08901_),
    .B1(_08393_),
    .A1(\cpu.icache.r_tag[7][17] ),
    .Y(_08902_),
    .A2(_08305_));
 sg13g2_a22oi_1 _15642_ (.Y(_08903_),
    .B1(net639),
    .B2(\cpu.icache.r_tag[6][17] ),
    .A2(_08654_),
    .A1(\cpu.icache.r_tag[3][17] ));
 sg13g2_a22oi_1 _15643_ (.Y(_08904_),
    .B1(_08323_),
    .B2(\cpu.icache.r_tag[2][17] ),
    .A2(net635),
    .A1(\cpu.icache.r_tag[1][17] ));
 sg13g2_nand4_1 _15644_ (.B(_08902_),
    .C(_08903_),
    .A(net554),
    .Y(_08905_),
    .D(_08904_));
 sg13g2_o21ai_1 _15645_ (.B1(_08905_),
    .Y(_08906_),
    .A1(\cpu.icache.r_tag[0][17] ),
    .A2(_08736_));
 sg13g2_xnor2_1 _15646_ (.Y(_08907_),
    .A(_08900_),
    .B(_08906_));
 sg13g2_mux4_1 _15647_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S1(net912),
    .X(_08908_));
 sg13g2_mux4_1 _15648_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S1(net912),
    .X(_08909_));
 sg13g2_mux4_1 _15649_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S1(net907),
    .X(_08910_));
 sg13g2_mux4_1 _15650_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S1(net907),
    .X(_08911_));
 sg13g2_mux4_1 _15651_ (.S0(_08633_),
    .A0(_08908_),
    .A1(_08909_),
    .A2(_08910_),
    .A3(_08911_),
    .S1(_08634_),
    .X(_08912_));
 sg13g2_mux4_1 _15652_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S1(net912),
    .X(_08913_));
 sg13g2_mux4_1 _15653_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S1(net912),
    .X(_08914_));
 sg13g2_mux4_1 _15654_ (.S0(_08721_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S1(_08722_),
    .X(_08915_));
 sg13g2_mux4_1 _15655_ (.S0(_08721_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S1(_08722_),
    .X(_08916_));
 sg13g2_mux4_1 _15656_ (.S0(_08633_),
    .A0(_08913_),
    .A1(_08914_),
    .A2(_08915_),
    .A3(_08916_),
    .S1(_08634_),
    .X(_08917_));
 sg13g2_mux2_1 _15657_ (.A0(_08912_),
    .A1(_08917_),
    .S(_08621_),
    .X(_08918_));
 sg13g2_nand2b_1 _15658_ (.Y(_08919_),
    .B(_08918_),
    .A_N(net1053));
 sg13g2_buf_1 _15659_ (.A(_08919_),
    .X(_08920_));
 sg13g2_a22oi_1 _15660_ (.Y(_08921_),
    .B1(_08654_),
    .B2(\cpu.icache.r_tag[3][21] ),
    .A2(net547),
    .A1(\cpu.icache.r_tag[2][21] ));
 sg13g2_buf_1 _15661_ (.A(net639),
    .X(_08922_));
 sg13g2_a22oi_1 _15662_ (.Y(_08923_),
    .B1(net544),
    .B2(\cpu.icache.r_tag[6][21] ),
    .A2(_08650_),
    .A1(\cpu.icache.r_tag[1][21] ));
 sg13g2_mux2_1 _15663_ (.A0(\cpu.icache.r_tag[5][21] ),
    .A1(\cpu.icache.r_tag[7][21] ),
    .S(_08276_),
    .X(_08924_));
 sg13g2_a22oi_1 _15664_ (.Y(_08925_),
    .B1(_08924_),
    .B2(net792),
    .A2(_08359_),
    .A1(\cpu.icache.r_tag[4][21] ));
 sg13g2_or2_1 _15665_ (.X(_08926_),
    .B(_08925_),
    .A(_08657_));
 sg13g2_nand4_1 _15666_ (.B(_08921_),
    .C(_08923_),
    .A(net478),
    .Y(_08927_),
    .D(_08926_));
 sg13g2_o21ai_1 _15667_ (.B1(_08927_),
    .Y(_08928_),
    .A1(\cpu.icache.r_tag[0][21] ),
    .A2(net482));
 sg13g2_xor2_1 _15668_ (.B(_08928_),
    .A(net422),
    .X(_08929_));
 sg13g2_inv_1 _15669_ (.Y(_08930_),
    .A(_08929_));
 sg13g2_and4_1 _15670_ (.A(_08862_),
    .B(_08887_),
    .C(_08907_),
    .D(_08930_),
    .X(_08931_));
 sg13g2_mux4_1 _15671_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S1(net914),
    .X(_08932_));
 sg13g2_mux4_1 _15672_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S1(net914),
    .X(_08933_));
 sg13g2_mux4_1 _15673_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S1(net904),
    .X(_08934_));
 sg13g2_mux4_1 _15674_ (.S0(_08843_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S1(_08844_),
    .X(_08935_));
 sg13g2_mux4_1 _15675_ (.S0(net908),
    .A0(_08932_),
    .A1(_08933_),
    .A2(_08934_),
    .A3(_08935_),
    .S1(net913),
    .X(_08936_));
 sg13g2_mux4_1 _15676_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S1(net904),
    .X(_08937_));
 sg13g2_mux4_1 _15677_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S1(net914),
    .X(_08938_));
 sg13g2_mux4_1 _15678_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S1(net910),
    .X(_08939_));
 sg13g2_mux4_1 _15679_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S1(net910),
    .X(_08940_));
 sg13g2_mux4_1 _15680_ (.S0(net908),
    .A0(_08937_),
    .A1(_08938_),
    .A2(_08939_),
    .A3(_08940_),
    .S1(net913),
    .X(_08941_));
 sg13g2_mux2_1 _15681_ (.A0(_08936_),
    .A1(_08941_),
    .S(net1056),
    .X(_08942_));
 sg13g2_nand2b_1 _15682_ (.Y(_08943_),
    .B(_08942_),
    .A_N(net1053));
 sg13g2_buf_2 _15683_ (.A(_08943_),
    .X(_08944_));
 sg13g2_nand2_1 _15684_ (.Y(_08945_),
    .A(\cpu.icache.r_tag[4][16] ),
    .B(_08651_));
 sg13g2_a22oi_1 _15685_ (.Y(_08946_),
    .B1(_08327_),
    .B2(\cpu.icache.r_tag[6][16] ),
    .A2(_08653_),
    .A1(\cpu.icache.r_tag[2][16] ));
 sg13g2_buf_1 _15686_ (.A(_08305_),
    .X(_08947_));
 sg13g2_a22oi_1 _15687_ (.Y(_08948_),
    .B1(_08761_),
    .B2(\cpu.icache.r_tag[3][16] ),
    .A2(net929),
    .A1(\cpu.icache.r_tag[5][16] ));
 sg13g2_nor2_1 _15688_ (.A(_08279_),
    .B(_08948_),
    .Y(_08949_));
 sg13g2_a221oi_1 _15689_ (.B2(\cpu.icache.r_tag[7][16] ),
    .C1(_08949_),
    .B1(_08947_),
    .A1(\cpu.icache.r_tag[1][16] ),
    .Y(_08950_),
    .A2(_08382_));
 sg13g2_nand4_1 _15690_ (.B(_08945_),
    .C(_08946_),
    .A(net478),
    .Y(_08951_),
    .D(_08950_));
 sg13g2_o21ai_1 _15691_ (.B1(_08951_),
    .Y(_08952_),
    .A1(\cpu.icache.r_tag[0][16] ),
    .A2(net482));
 sg13g2_xnor2_1 _15692_ (.Y(_08953_),
    .A(net421),
    .B(_08952_));
 sg13g2_mux4_1 _15693_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S1(net917),
    .X(_08954_));
 sg13g2_mux4_1 _15694_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S1(net917),
    .X(_08955_));
 sg13g2_mux4_1 _15695_ (.S0(_08843_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S1(_08844_),
    .X(_08956_));
 sg13g2_mux4_1 _15696_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S1(net904),
    .X(_08957_));
 sg13g2_mux4_1 _15697_ (.S0(net908),
    .A0(_08954_),
    .A1(_08955_),
    .A2(_08956_),
    .A3(_08957_),
    .S1(net913),
    .X(_08958_));
 sg13g2_mux4_1 _15698_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S1(net914),
    .X(_08959_));
 sg13g2_mux4_1 _15699_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S1(net914),
    .X(_08960_));
 sg13g2_mux4_1 _15700_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S1(net904),
    .X(_08961_));
 sg13g2_mux4_1 _15701_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S1(net904),
    .X(_08962_));
 sg13g2_mux4_1 _15702_ (.S0(net908),
    .A0(_08959_),
    .A1(_08960_),
    .A2(_08961_),
    .A3(_08962_),
    .S1(net913),
    .X(_08963_));
 sg13g2_mux2_1 _15703_ (.A0(_08958_),
    .A1(_08963_),
    .S(net1056),
    .X(_08964_));
 sg13g2_nand2b_1 _15704_ (.Y(_08965_),
    .B(_08964_),
    .A_N(_08695_));
 sg13g2_buf_1 _15705_ (.A(_08965_),
    .X(_08966_));
 sg13g2_a22oi_1 _15706_ (.Y(_08967_),
    .B1(_08653_),
    .B2(\cpu.icache.r_tag[2][22] ),
    .A2(_08650_),
    .A1(\cpu.icache.r_tag[1][22] ));
 sg13g2_a22oi_1 _15707_ (.Y(_08968_),
    .B1(_08327_),
    .B2(\cpu.icache.r_tag[6][22] ),
    .A2(_08651_),
    .A1(\cpu.icache.r_tag[4][22] ));
 sg13g2_mux2_1 _15708_ (.A0(\cpu.icache.r_tag[7][22] ),
    .A1(\cpu.icache.r_tag[3][22] ),
    .S(net924),
    .X(_08969_));
 sg13g2_a22oi_1 _15709_ (.Y(_08970_),
    .B1(_08969_),
    .B2(net698),
    .A2(_08283_),
    .A1(\cpu.icache.r_tag[5][22] ));
 sg13g2_nand2b_1 _15710_ (.Y(_08971_),
    .B(_08342_),
    .A_N(_08970_));
 sg13g2_nand3_1 _15711_ (.B(_08968_),
    .C(_08971_),
    .A(_08967_),
    .Y(_08972_));
 sg13g2_mux2_1 _15712_ (.A0(\cpu.icache.r_tag[0][22] ),
    .A1(_08972_),
    .S(net478),
    .X(_08973_));
 sg13g2_xor2_1 _15713_ (.B(_08973_),
    .A(net420),
    .X(_08974_));
 sg13g2_mux4_1 _15714_ (.S0(_08865_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S1(_08866_),
    .X(_08975_));
 sg13g2_mux4_1 _15715_ (.S0(net903),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S1(net1049),
    .X(_08976_));
 sg13g2_mux4_1 _15716_ (.S0(net921),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S1(_08866_),
    .X(_08977_));
 sg13g2_mux4_1 _15717_ (.S0(_08865_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S1(net1049),
    .X(_08978_));
 sg13g2_mux4_1 _15718_ (.S0(net1061),
    .A0(_08975_),
    .A1(_08976_),
    .A2(_08977_),
    .A3(_08978_),
    .S1(_08549_),
    .X(_08979_));
 sg13g2_a21oi_1 _15719_ (.A1(net1057),
    .A2(_08979_),
    .Y(_08980_),
    .B1(_08538_));
 sg13g2_mux4_1 _15720_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S1(_08707_),
    .X(_08981_));
 sg13g2_mux4_1 _15721_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S1(net1052),
    .X(_08982_));
 sg13g2_mux4_1 _15722_ (.S0(net903),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S1(net1052),
    .X(_08983_));
 sg13g2_mux4_1 _15723_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S1(net1052),
    .X(_08984_));
 sg13g2_mux4_1 _15724_ (.S0(net1061),
    .A0(_08981_),
    .A1(_08982_),
    .A2(_08983_),
    .A3(_08984_),
    .S1(_08620_),
    .X(_08985_));
 sg13g2_nor3_1 _15725_ (.A(net916),
    .B(_08464_),
    .C(_08985_),
    .Y(_08986_));
 sg13g2_or2_1 _15726_ (.X(_08987_),
    .B(_08986_),
    .A(_08980_));
 sg13g2_buf_2 _15727_ (.A(_08987_),
    .X(_08988_));
 sg13g2_a22oi_1 _15728_ (.Y(_08989_),
    .B1(net705),
    .B2(\cpu.icache.r_tag[4][15] ),
    .A2(_08382_),
    .A1(\cpu.icache.r_tag[1][15] ));
 sg13g2_a22oi_1 _15729_ (.Y(_08990_),
    .B1(_08329_),
    .B2(\cpu.icache.r_tag[5][15] ),
    .A2(_08348_),
    .A1(\cpu.icache.r_tag[2][15] ));
 sg13g2_mux2_1 _15730_ (.A0(\cpu.icache.r_tag[7][15] ),
    .A1(\cpu.icache.r_tag[3][15] ),
    .S(net924),
    .X(_08991_));
 sg13g2_a22oi_1 _15731_ (.Y(_08992_),
    .B1(_08991_),
    .B2(_08341_),
    .A2(_08780_),
    .A1(\cpu.icache.r_tag[6][15] ));
 sg13g2_nand2b_1 _15732_ (.Y(_08993_),
    .B(net702),
    .A_N(_08992_));
 sg13g2_nand4_1 _15733_ (.B(_08989_),
    .C(_08990_),
    .A(_08333_),
    .Y(_08994_),
    .D(_08993_));
 sg13g2_o21ai_1 _15734_ (.B1(_08994_),
    .Y(_08995_),
    .A1(\cpu.icache.r_tag[0][15] ),
    .A2(net478));
 sg13g2_xnor2_1 _15735_ (.Y(_08996_),
    .A(net474),
    .B(_08995_));
 sg13g2_nand4_1 _15736_ (.B(_08953_),
    .C(_08974_),
    .A(_08931_),
    .Y(_08997_),
    .D(_08996_));
 sg13g2_nor4_1 _15737_ (.A(_08462_),
    .B(_08616_),
    .C(_08840_),
    .D(_08997_),
    .Y(_08998_));
 sg13g2_buf_1 _15738_ (.A(_08998_),
    .X(_08999_));
 sg13g2_buf_1 _15739_ (.A(_08999_),
    .X(_09000_));
 sg13g2_mux2_1 _15740_ (.A0(net1073),
    .A1(_08461_),
    .S(net119),
    .X(_00016_));
 sg13g2_buf_2 _15741_ (.A(\cpu.dec.r_op[4] ),
    .X(_09001_));
 sg13g2_buf_1 _15742_ (.A(_09001_),
    .X(_09002_));
 sg13g2_nand2_1 _15743_ (.Y(_09003_),
    .A(_08862_),
    .B(_08953_));
 sg13g2_nand2b_1 _15744_ (.Y(_09004_),
    .B(_08974_),
    .A_N(_08767_));
 sg13g2_nor2_1 _15745_ (.A(_09003_),
    .B(_09004_),
    .Y(_09005_));
 sg13g2_nand3_1 _15746_ (.B(_08907_),
    .C(_08996_),
    .A(_08887_),
    .Y(_09006_));
 sg13g2_nand4_1 _15747_ (.B(_08814_),
    .C(_08818_),
    .A(_08796_),
    .Y(_09007_),
    .D(_08828_));
 sg13g2_nand4_1 _15748_ (.B(_08785_),
    .C(_08805_),
    .A(_08776_),
    .Y(_09008_),
    .D(_08837_));
 sg13g2_nor2_1 _15749_ (.A(_09007_),
    .B(_09008_),
    .Y(_09009_));
 sg13g2_nand2_1 _15750_ (.Y(_09010_),
    .A(_08720_),
    .B(_09009_));
 sg13g2_nor4_1 _15751_ (.A(_08744_),
    .B(_08929_),
    .C(_09006_),
    .D(_09010_),
    .Y(_09011_));
 sg13g2_nand3_1 _15752_ (.B(_09005_),
    .C(_09011_),
    .A(_08693_),
    .Y(_09012_));
 sg13g2_nor3_1 _15753_ (.A(_08462_),
    .B(net294),
    .C(_09012_),
    .Y(_09013_));
 sg13g2_buf_2 _15754_ (.A(_09013_),
    .X(_09014_));
 sg13g2_inv_1 _15755_ (.Y(_09015_),
    .A(_09014_));
 sg13g2_buf_1 _15756_ (.A(_09015_),
    .X(_09016_));
 sg13g2_buf_1 _15757_ (.A(net89),
    .X(_09017_));
 sg13g2_inv_1 _15758_ (.Y(_09018_),
    .A(_00212_));
 sg13g2_mux2_1 _15759_ (.A0(\cpu.icache.r_data[7][28] ),
    .A1(\cpu.icache.r_data[3][28] ),
    .S(net1071),
    .X(_09019_));
 sg13g2_a22oi_1 _15760_ (.Y(_09020_),
    .B1(_09019_),
    .B2(net925),
    .A2(net795),
    .A1(\cpu.icache.r_data[6][28] ));
 sg13g2_nand2b_1 _15761_ (.Y(_09021_),
    .B(_08276_),
    .A_N(_09020_));
 sg13g2_a22oi_1 _15762_ (.Y(_09022_),
    .B1(net796),
    .B2(\cpu.icache.r_data[4][28] ),
    .A2(_08288_),
    .A1(\cpu.icache.r_data[1][28] ));
 sg13g2_a22oi_1 _15763_ (.Y(_09023_),
    .B1(_08285_),
    .B2(\cpu.icache.r_data[5][28] ),
    .A2(_08281_),
    .A1(\cpu.icache.r_data[2][28] ));
 sg13g2_nand3_1 _15764_ (.B(_09022_),
    .C(_09023_),
    .A(_09021_),
    .Y(_09024_));
 sg13g2_a21oi_1 _15765_ (.A1(_09018_),
    .A2(net553),
    .Y(_09025_),
    .B1(_09024_));
 sg13g2_nand2_1 _15766_ (.Y(_09026_),
    .A(_00211_),
    .B(_08271_));
 sg13g2_a22oi_1 _15767_ (.Y(_09027_),
    .B1(net796),
    .B2(\cpu.icache.r_data[4][12] ),
    .A2(_08288_),
    .A1(\cpu.icache.r_data[1][12] ));
 sg13g2_a22oi_1 _15768_ (.Y(_09028_),
    .B1(_08299_),
    .B2(\cpu.icache.r_data[3][12] ),
    .A2(_08281_),
    .A1(\cpu.icache.r_data[2][12] ));
 sg13g2_mux2_1 _15769_ (.A0(\cpu.icache.r_data[5][12] ),
    .A1(\cpu.icache.r_data[7][12] ),
    .S(net1069),
    .X(_09029_));
 sg13g2_a22oi_1 _15770_ (.Y(_09030_),
    .B1(_09029_),
    .B2(net1070),
    .A2(_08660_),
    .A1(\cpu.icache.r_data[6][12] ));
 sg13g2_or2_1 _15771_ (.X(_09031_),
    .B(_09030_),
    .A(net924));
 sg13g2_nand4_1 _15772_ (.B(_09027_),
    .C(_09028_),
    .A(net637),
    .Y(_09032_),
    .D(_09031_));
 sg13g2_a21oi_1 _15773_ (.A1(_09026_),
    .A2(_09032_),
    .Y(_09033_),
    .B1(_08258_));
 sg13g2_a21o_1 _15774_ (.A2(_09025_),
    .A1(net928),
    .B1(_09033_),
    .X(_09034_));
 sg13g2_buf_2 _15775_ (.A(_09034_),
    .X(_09035_));
 sg13g2_buf_1 _15776_ (.A(_09035_),
    .X(_09036_));
 sg13g2_and2_1 _15777_ (.A(_08310_),
    .B(_08458_),
    .X(_09037_));
 sg13g2_buf_1 _15778_ (.A(_09037_),
    .X(_09038_));
 sg13g2_a21o_1 _15779_ (.A2(_08388_),
    .A1(net926),
    .B1(_08402_),
    .X(_09039_));
 sg13g2_buf_1 _15780_ (.A(_09039_),
    .X(_09040_));
 sg13g2_mux2_1 _15781_ (.A0(_08417_),
    .A1(_08410_),
    .S(net923),
    .X(_09041_));
 sg13g2_buf_1 _15782_ (.A(_09041_),
    .X(_09042_));
 sg13g2_a21oi_1 _15783_ (.A1(_08335_),
    .A2(_08427_),
    .Y(_09043_),
    .B1(_08435_));
 sg13g2_buf_1 _15784_ (.A(_09043_),
    .X(_09044_));
 sg13g2_nor2_1 _15785_ (.A(_09042_),
    .B(_09044_),
    .Y(_09045_));
 sg13g2_buf_2 _15786_ (.A(_09045_),
    .X(_09046_));
 sg13g2_nand2_1 _15787_ (.Y(_09047_),
    .A(net292),
    .B(_09046_));
 sg13g2_buf_2 _15788_ (.A(_09047_),
    .X(_09048_));
 sg13g2_inv_1 _15789_ (.Y(_09049_),
    .A(_08354_));
 sg13g2_nand2_1 _15790_ (.Y(_09050_),
    .A(_09049_),
    .B(net223));
 sg13g2_buf_1 _15791_ (.A(_09050_),
    .X(_09051_));
 sg13g2_nor2_2 _15792_ (.A(_09048_),
    .B(_09051_),
    .Y(_09052_));
 sg13g2_nand2_1 _15793_ (.Y(_09053_),
    .A(_09038_),
    .B(_09052_));
 sg13g2_nor2_1 _15794_ (.A(_00210_),
    .B(net550),
    .Y(_09054_));
 sg13g2_mux2_1 _15795_ (.A0(\cpu.icache.r_data[4][22] ),
    .A1(\cpu.icache.r_data[6][22] ),
    .S(net797),
    .X(_09055_));
 sg13g2_a22oi_1 _15796_ (.Y(_09056_),
    .B1(_09055_),
    .B2(net930),
    .A2(net704),
    .A1(\cpu.icache.r_data[7][22] ));
 sg13g2_nor2_1 _15797_ (.A(net786),
    .B(_09056_),
    .Y(_09057_));
 sg13g2_a22oi_1 _15798_ (.Y(_09058_),
    .B1(net552),
    .B2(\cpu.icache.r_data[2][22] ),
    .A2(net641),
    .A1(\cpu.icache.r_data[1][22] ));
 sg13g2_a22oi_1 _15799_ (.Y(_09059_),
    .B1(net634),
    .B2(\cpu.icache.r_data[5][22] ),
    .A2(net551),
    .A1(\cpu.icache.r_data[3][22] ));
 sg13g2_nand2_1 _15800_ (.Y(_09060_),
    .A(_09058_),
    .B(_09059_));
 sg13g2_nor3_1 _15801_ (.A(_09054_),
    .B(_09057_),
    .C(_09060_),
    .Y(_09061_));
 sg13g2_nand2_1 _15802_ (.Y(_09062_),
    .A(_00209_),
    .B(net553));
 sg13g2_a22oi_1 _15803_ (.Y(_09063_),
    .B1(net699),
    .B2(\cpu.icache.r_data[4][6] ),
    .A2(net700),
    .A1(\cpu.icache.r_data[1][6] ));
 sg13g2_a22oi_1 _15804_ (.Y(_09064_),
    .B1(net551),
    .B2(\cpu.icache.r_data[3][6] ),
    .A2(net640),
    .A1(\cpu.icache.r_data[2][6] ));
 sg13g2_mux2_1 _15805_ (.A0(\cpu.icache.r_data[5][6] ),
    .A1(\cpu.icache.r_data[7][6] ),
    .S(net931),
    .X(_09065_));
 sg13g2_a22oi_1 _15806_ (.Y(_09066_),
    .B1(_09065_),
    .B2(_08340_),
    .A2(_08660_),
    .A1(\cpu.icache.r_data[6][6] ));
 sg13g2_or2_1 _15807_ (.X(_09067_),
    .B(_09066_),
    .A(net927));
 sg13g2_nand4_1 _15808_ (.B(_09063_),
    .C(_09064_),
    .A(net550),
    .Y(_09068_),
    .D(_09067_));
 sg13g2_a21oi_1 _15809_ (.A1(_09062_),
    .A2(_09068_),
    .Y(_09069_),
    .B1(net928));
 sg13g2_a21oi_2 _15810_ (.B1(_09069_),
    .Y(_09070_),
    .A2(_09061_),
    .A1(_08335_));
 sg13g2_buf_1 _15811_ (.A(_09070_),
    .X(_09071_));
 sg13g2_inv_2 _15812_ (.Y(_09072_),
    .A(net290));
 sg13g2_inv_1 _15813_ (.Y(_09073_),
    .A(_00208_));
 sg13g2_mux2_1 _15814_ (.A0(\cpu.icache.r_data[7][21] ),
    .A1(\cpu.icache.r_data[3][21] ),
    .S(net927),
    .X(_09074_));
 sg13g2_a22oi_1 _15815_ (.Y(_09075_),
    .B1(_09074_),
    .B2(_08341_),
    .A2(net697),
    .A1(\cpu.icache.r_data[6][21] ));
 sg13g2_nand2b_1 _15816_ (.Y(_09076_),
    .B(_08338_),
    .A_N(_09075_));
 sg13g2_a22oi_1 _15817_ (.Y(_09077_),
    .B1(net633),
    .B2(\cpu.icache.r_data[4][21] ),
    .A2(net548),
    .A1(\cpu.icache.r_data[1][21] ));
 sg13g2_buf_1 _15818_ (.A(_08393_),
    .X(_09078_));
 sg13g2_a22oi_1 _15819_ (.Y(_09079_),
    .B1(net542),
    .B2(\cpu.icache.r_data[5][21] ),
    .A2(net547),
    .A1(\cpu.icache.r_data[2][21] ));
 sg13g2_nand3_1 _15820_ (.B(_09077_),
    .C(_09079_),
    .A(_09076_),
    .Y(_09080_));
 sg13g2_a21oi_1 _15821_ (.A1(_09073_),
    .A2(_08345_),
    .Y(_09081_),
    .B1(_09080_));
 sg13g2_nand2_1 _15822_ (.Y(_09082_),
    .A(_00207_),
    .B(net483));
 sg13g2_a22oi_1 _15823_ (.Y(_09083_),
    .B1(net633),
    .B2(\cpu.icache.r_data[4][5] ),
    .A2(net548),
    .A1(\cpu.icache.r_data[1][5] ));
 sg13g2_a22oi_1 _15824_ (.Y(_09084_),
    .B1(net639),
    .B2(\cpu.icache.r_data[6][5] ),
    .A2(net547),
    .A1(\cpu.icache.r_data[2][5] ));
 sg13g2_mux2_1 _15825_ (.A0(\cpu.icache.r_data[7][5] ),
    .A1(\cpu.icache.r_data[3][5] ),
    .S(_08366_),
    .X(_09085_));
 sg13g2_a22oi_1 _15826_ (.Y(_09086_),
    .B1(_09085_),
    .B2(_08399_),
    .A2(net929),
    .A1(\cpu.icache.r_data[5][5] ));
 sg13g2_nand2b_1 _15827_ (.Y(_09087_),
    .B(_08342_),
    .A_N(_09086_));
 sg13g2_nand4_1 _15828_ (.B(_09083_),
    .C(_09084_),
    .A(_08736_),
    .Y(_09088_),
    .D(_09087_));
 sg13g2_a21oi_1 _15829_ (.A1(_09082_),
    .A2(_09088_),
    .Y(_09089_),
    .B1(net926));
 sg13g2_a21oi_1 _15830_ (.A1(net794),
    .A2(_09081_),
    .Y(_09090_),
    .B1(_09089_));
 sg13g2_buf_1 _15831_ (.A(_09090_),
    .X(_09091_));
 sg13g2_inv_1 _15832_ (.Y(_09092_),
    .A(net289));
 sg13g2_buf_1 _15833_ (.A(_09092_),
    .X(_09093_));
 sg13g2_nand2_1 _15834_ (.Y(_09094_),
    .A(_09072_),
    .B(net222));
 sg13g2_nor4_1 _15835_ (.A(net89),
    .B(_09036_),
    .C(_09053_),
    .D(_09094_),
    .Y(_09095_));
 sg13g2_a21o_1 _15836_ (.A2(_09017_),
    .A1(net1048),
    .B1(_09095_),
    .X(_00015_));
 sg13g2_nand2_1 _15837_ (.Y(_09096_),
    .A(_09036_),
    .B(_09071_));
 sg13g2_buf_1 _15838_ (.A(_08310_),
    .X(_09097_));
 sg13g2_o21ai_1 _15839_ (.B1(net288),
    .Y(_09098_),
    .A1(net222),
    .A2(_09096_));
 sg13g2_nand4_1 _15840_ (.B(_08440_),
    .C(net295),
    .A(net172),
    .Y(_09099_),
    .D(_09098_));
 sg13g2_buf_1 _15841_ (.A(\cpu.dec.r_op[2] ),
    .X(_09100_));
 sg13g2_buf_1 _15842_ (.A(net1124),
    .X(_09101_));
 sg13g2_nand2_1 _15843_ (.Y(_09102_),
    .A(net1047),
    .B(net89));
 sg13g2_o21ai_1 _15844_ (.B1(_09102_),
    .Y(_00013_),
    .A1(net79),
    .A2(_09099_));
 sg13g2_buf_1 _15845_ (.A(_08999_),
    .X(_09103_));
 sg13g2_buf_1 _15846_ (.A(net118),
    .X(_09104_));
 sg13g2_nor2b_1 _15847_ (.A(_08441_),
    .B_N(_09038_),
    .Y(_09105_));
 sg13g2_nand2_1 _15848_ (.Y(_09106_),
    .A(_09035_),
    .B(_09072_));
 sg13g2_nor2_1 _15849_ (.A(net222),
    .B(_09106_),
    .Y(_09107_));
 sg13g2_nor2_1 _15850_ (.A(_09035_),
    .B(_09070_),
    .Y(_09108_));
 sg13g2_nand4_1 _15851_ (.B(_09052_),
    .C(net289),
    .A(_09038_),
    .Y(_09109_),
    .D(_09108_));
 sg13g2_inv_1 _15852_ (.Y(_09110_),
    .A(_00218_));
 sg13g2_mux2_1 _15853_ (.A0(\cpu.icache.r_data[4][20] ),
    .A1(\cpu.icache.r_data[6][20] ),
    .S(net793),
    .X(_09111_));
 sg13g2_a22oi_1 _15854_ (.Y(_09112_),
    .B1(net697),
    .B2(_09111_),
    .A2(net556),
    .A1(\cpu.icache.r_data[2][20] ));
 sg13g2_a22oi_1 _15855_ (.Y(_09113_),
    .B1(_08305_),
    .B2(\cpu.icache.r_data[7][20] ),
    .A2(net481),
    .A1(\cpu.icache.r_data[3][20] ));
 sg13g2_a22oi_1 _15856_ (.Y(_09114_),
    .B1(net555),
    .B2(\cpu.icache.r_data[5][20] ),
    .A2(net635),
    .A1(\cpu.icache.r_data[1][20] ));
 sg13g2_nand3_1 _15857_ (.B(_09113_),
    .C(_09114_),
    .A(_09112_),
    .Y(_09115_));
 sg13g2_a21oi_1 _15858_ (.A1(_09110_),
    .A2(net483),
    .Y(_09116_),
    .B1(_09115_));
 sg13g2_nand2_1 _15859_ (.Y(_09117_),
    .A(_00217_),
    .B(_08345_));
 sg13g2_a22oi_1 _15860_ (.Y(_09118_),
    .B1(net555),
    .B2(\cpu.icache.r_data[5][4] ),
    .A2(net705),
    .A1(\cpu.icache.r_data[4][4] ));
 sg13g2_a22oi_1 _15861_ (.Y(_09119_),
    .B1(net556),
    .B2(\cpu.icache.r_data[2][4] ),
    .A2(net635),
    .A1(\cpu.icache.r_data[1][4] ));
 sg13g2_mux2_1 _15862_ (.A0(\cpu.icache.r_data[7][4] ),
    .A1(\cpu.icache.r_data[3][4] ),
    .S(_08316_),
    .X(_09120_));
 sg13g2_a22oi_1 _15863_ (.Y(_09121_),
    .B1(_09120_),
    .B2(_08397_),
    .A2(net697),
    .A1(\cpu.icache.r_data[6][4] ));
 sg13g2_nand2b_1 _15864_ (.Y(_09122_),
    .B(_08399_),
    .A_N(_09121_));
 sg13g2_nand4_1 _15865_ (.B(_09118_),
    .C(_09119_),
    .A(net554),
    .Y(_09123_),
    .D(_09122_));
 sg13g2_a21oi_1 _15866_ (.A1(_09117_),
    .A2(_09123_),
    .Y(_09124_),
    .B1(net928));
 sg13g2_a21oi_1 _15867_ (.A1(net794),
    .A2(_09116_),
    .Y(_09125_),
    .B1(_09124_));
 sg13g2_buf_1 _15868_ (.A(_09125_),
    .X(_09126_));
 sg13g2_buf_1 _15869_ (.A(_09126_),
    .X(_09127_));
 sg13g2_a22oi_1 _15870_ (.Y(_09128_),
    .B1(net634),
    .B2(\cpu.icache.r_data[5][2] ),
    .A2(net699),
    .A1(\cpu.icache.r_data[4][2] ));
 sg13g2_a22oi_1 _15871_ (.Y(_09129_),
    .B1(net640),
    .B2(\cpu.icache.r_data[2][2] ),
    .A2(net700),
    .A1(\cpu.icache.r_data[1][2] ));
 sg13g2_mux2_1 _15872_ (.A0(\cpu.icache.r_data[7][2] ),
    .A1(\cpu.icache.r_data[3][2] ),
    .S(net1068),
    .X(_09130_));
 sg13g2_a22oi_1 _15873_ (.Y(_09131_),
    .B1(_09130_),
    .B2(net791),
    .A2(net795),
    .A1(\cpu.icache.r_data[6][2] ));
 sg13g2_nand2b_1 _15874_ (.Y(_09132_),
    .B(net698),
    .A_N(_09131_));
 sg13g2_and4_1 _15875_ (.A(net549),
    .B(_09128_),
    .C(_09129_),
    .D(_09132_),
    .X(_09133_));
 sg13g2_a21oi_1 _15876_ (.A1(_00213_),
    .A2(net483),
    .Y(_09134_),
    .B1(_09133_));
 sg13g2_nor2_1 _15877_ (.A(_00214_),
    .B(net554),
    .Y(_09135_));
 sg13g2_mux2_1 _15878_ (.A0(\cpu.icache.r_data[7][18] ),
    .A1(\cpu.icache.r_data[3][18] ),
    .S(net1068),
    .X(_09136_));
 sg13g2_a22oi_1 _15879_ (.Y(_09137_),
    .B1(_09136_),
    .B2(net791),
    .A2(net697),
    .A1(\cpu.icache.r_data[6][18] ));
 sg13g2_nand2b_1 _15880_ (.Y(_09138_),
    .B(net698),
    .A_N(_09137_));
 sg13g2_a22oi_1 _15881_ (.Y(_09139_),
    .B1(net705),
    .B2(\cpu.icache.r_data[4][18] ),
    .A2(net641),
    .A1(\cpu.icache.r_data[1][18] ));
 sg13g2_a22oi_1 _15882_ (.Y(_09140_),
    .B1(net634),
    .B2(\cpu.icache.r_data[5][18] ),
    .A2(net552),
    .A1(\cpu.icache.r_data[2][18] ));
 sg13g2_nand3_1 _15883_ (.B(_09139_),
    .C(_09140_),
    .A(_09138_),
    .Y(_09141_));
 sg13g2_or3_1 _15884_ (.A(net923),
    .B(_09135_),
    .C(_09141_),
    .X(_09142_));
 sg13g2_o21ai_1 _15885_ (.B1(_09142_),
    .Y(_09143_),
    .A1(net926),
    .A2(_09134_));
 sg13g2_buf_2 _15886_ (.A(_09143_),
    .X(_09144_));
 sg13g2_inv_2 _15887_ (.Y(_09145_),
    .A(_09144_));
 sg13g2_inv_1 _15888_ (.Y(_09146_),
    .A(_00216_));
 sg13g2_mux2_1 _15889_ (.A0(\cpu.icache.r_data[7][19] ),
    .A1(\cpu.icache.r_data[3][19] ),
    .S(net1068),
    .X(_09147_));
 sg13g2_a22oi_1 _15890_ (.Y(_09148_),
    .B1(_09147_),
    .B2(net791),
    .A2(net697),
    .A1(\cpu.icache.r_data[6][19] ));
 sg13g2_nand2b_1 _15891_ (.Y(_09149_),
    .B(net698),
    .A_N(_09148_));
 sg13g2_a22oi_1 _15892_ (.Y(_09150_),
    .B1(net705),
    .B2(\cpu.icache.r_data[4][19] ),
    .A2(net641),
    .A1(\cpu.icache.r_data[1][19] ));
 sg13g2_a22oi_1 _15893_ (.Y(_09151_),
    .B1(net634),
    .B2(\cpu.icache.r_data[5][19] ),
    .A2(net552),
    .A1(\cpu.icache.r_data[2][19] ));
 sg13g2_nand3_1 _15894_ (.B(_09150_),
    .C(_09151_),
    .A(_09149_),
    .Y(_09152_));
 sg13g2_a21oi_1 _15895_ (.A1(_09146_),
    .A2(net483),
    .Y(_09153_),
    .B1(_09152_));
 sg13g2_nand2_1 _15896_ (.Y(_09154_),
    .A(_00215_),
    .B(net483));
 sg13g2_mux2_1 _15897_ (.A0(\cpu.icache.r_data[4][3] ),
    .A1(\cpu.icache.r_data[6][3] ),
    .S(net797),
    .X(_09155_));
 sg13g2_a22oi_1 _15898_ (.Y(_09156_),
    .B1(net697),
    .B2(_09155_),
    .A2(net481),
    .A1(\cpu.icache.r_data[3][3] ));
 sg13g2_a22oi_1 _15899_ (.Y(_09157_),
    .B1(net552),
    .B2(\cpu.icache.r_data[2][3] ),
    .A2(net641),
    .A1(\cpu.icache.r_data[1][3] ));
 sg13g2_a22oi_1 _15900_ (.Y(_09158_),
    .B1(net634),
    .B2(\cpu.icache.r_data[5][3] ),
    .A2(_08305_),
    .A1(\cpu.icache.r_data[7][3] ));
 sg13g2_nand4_1 _15901_ (.B(_09156_),
    .C(_09157_),
    .A(net549),
    .Y(_09159_),
    .D(_09158_));
 sg13g2_a21oi_1 _15902_ (.A1(_09154_),
    .A2(_09159_),
    .Y(_09160_),
    .B1(net928));
 sg13g2_a21oi_1 _15903_ (.A1(net926),
    .A2(_09153_),
    .Y(_09161_),
    .B1(_09160_));
 sg13g2_buf_1 _15904_ (.A(_09161_),
    .X(_09162_));
 sg13g2_nand2_1 _15905_ (.Y(_09163_),
    .A(_09145_),
    .B(net246));
 sg13g2_nor3_1 _15906_ (.A(_09109_),
    .B(net221),
    .C(_09163_),
    .Y(_09164_));
 sg13g2_a21oi_1 _15907_ (.A1(_09105_),
    .A2(_09107_),
    .Y(_09165_),
    .B1(_09164_));
 sg13g2_buf_2 _15908_ (.A(\cpu.dec.r_op[3] ),
    .X(_09166_));
 sg13g2_buf_1 _15909_ (.A(_09166_),
    .X(_09167_));
 sg13g2_nor2_1 _15910_ (.A(net1046),
    .B(net119),
    .Y(_09168_));
 sg13g2_a21oi_1 _15911_ (.A1(net107),
    .A2(_09165_),
    .Y(_00014_),
    .B1(_09168_));
 sg13g2_nor2_2 _15912_ (.A(_09070_),
    .B(net289),
    .Y(_09169_));
 sg13g2_a21o_1 _15913_ (.A2(_09116_),
    .A1(_08313_),
    .B1(_09124_),
    .X(_09170_));
 sg13g2_buf_1 _15914_ (.A(_09170_),
    .X(_09171_));
 sg13g2_inv_1 _15915_ (.Y(_09172_),
    .A(_09161_));
 sg13g2_nand2_2 _15916_ (.Y(_09173_),
    .A(_09144_),
    .B(_09172_));
 sg13g2_nor2_2 _15917_ (.A(_09171_),
    .B(_09173_),
    .Y(_09174_));
 sg13g2_buf_1 _15918_ (.A(_09051_),
    .X(_09175_));
 sg13g2_nand3_1 _15919_ (.B(_09090_),
    .C(_09108_),
    .A(_09038_),
    .Y(_09176_));
 sg13g2_buf_2 _15920_ (.A(_09176_),
    .X(_09177_));
 sg13g2_nor3_2 _15921_ (.A(_09048_),
    .B(net144),
    .C(_09177_),
    .Y(_09178_));
 sg13g2_a22oi_1 _15922_ (.Y(_09179_),
    .B1(_09174_),
    .B2(_09178_),
    .A2(_09105_),
    .A1(_09169_));
 sg13g2_buf_2 _15923_ (.A(\cpu.dec.r_op[6] ),
    .X(_09180_));
 sg13g2_buf_1 _15924_ (.A(_09180_),
    .X(_09181_));
 sg13g2_nor2_1 _15925_ (.A(net1045),
    .B(net119),
    .Y(_09182_));
 sg13g2_a21oi_1 _15926_ (.A1(net107),
    .A2(_09179_),
    .Y(_00017_),
    .B1(_09182_));
 sg13g2_buf_1 _15927_ (.A(\cpu.spi.r_count[7] ),
    .X(_09183_));
 sg13g2_buf_1 _15928_ (.A(\cpu.spi.r_count[3] ),
    .X(_09184_));
 sg13g2_buf_1 _15929_ (.A(\cpu.spi.r_count[0] ),
    .X(_09185_));
 sg13g2_buf_1 _15930_ (.A(\cpu.spi.r_count[1] ),
    .X(_09186_));
 sg13g2_nor2_1 _15931_ (.A(_09185_),
    .B(_09186_),
    .Y(_09187_));
 sg13g2_nand2b_1 _15932_ (.Y(_09188_),
    .B(_09187_),
    .A_N(\cpu.spi.r_count[2] ));
 sg13g2_nor3_1 _15933_ (.A(_09184_),
    .B(\cpu.spi.r_count[4] ),
    .C(_09188_),
    .Y(_09189_));
 sg13g2_nor2b_1 _15934_ (.A(\cpu.spi.r_count[5] ),
    .B_N(_09189_),
    .Y(_09190_));
 sg13g2_nor2b_1 _15935_ (.A(\cpu.spi.r_count[6] ),
    .B_N(_09190_),
    .Y(_09191_));
 sg13g2_nand2b_1 _15936_ (.Y(_09192_),
    .B(_09191_),
    .A_N(_09183_));
 sg13g2_buf_1 _15937_ (.A(_09192_),
    .X(_09193_));
 sg13g2_buf_1 _15938_ (.A(_09193_),
    .X(_09194_));
 sg13g2_buf_1 _15939_ (.A(\cpu.spi.r_state[1] ),
    .X(_09195_));
 sg13g2_inv_2 _15940_ (.Y(_09196_),
    .A(_09195_));
 sg13g2_buf_1 _15941_ (.A(\cpu.addr[3] ),
    .X(_09197_));
 sg13g2_buf_1 _15942_ (.A(_09197_),
    .X(_09198_));
 sg13g2_buf_1 _15943_ (.A(net1044),
    .X(_09199_));
 sg13g2_buf_1 _15944_ (.A(net902),
    .X(_09200_));
 sg13g2_buf_1 _15945_ (.A(net784),
    .X(_09201_));
 sg13g2_buf_1 _15946_ (.A(\cpu.addr[8] ),
    .X(_09202_));
 sg13g2_buf_1 _15947_ (.A(_09202_),
    .X(_09203_));
 sg13g2_buf_1 _15948_ (.A(\cpu.addr[7] ),
    .X(_09204_));
 sg13g2_buf_1 _15949_ (.A(_09204_),
    .X(_09205_));
 sg13g2_buf_2 _15950_ (.A(\cpu.addr[6] ),
    .X(_09206_));
 sg13g2_nand3b_1 _15951_ (.B(net1042),
    .C(_09206_),
    .Y(_09207_),
    .A_N(net1043));
 sg13g2_buf_2 _15952_ (.A(_09207_),
    .X(_09208_));
 sg13g2_buf_1 _15953_ (.A(_08465_),
    .X(_09209_));
 sg13g2_buf_1 _15954_ (.A(\cpu.ex.r_wmask[0] ),
    .X(_09210_));
 sg13g2_or2_1 _15955_ (.X(_09211_),
    .B(net1123),
    .A(_08466_));
 sg13g2_buf_1 _15956_ (.A(\cpu.dec.r_trap ),
    .X(_09212_));
 sg13g2_nor2_2 _15957_ (.A(_09212_),
    .B(_08615_),
    .Y(_09213_));
 sg13g2_buf_1 _15958_ (.A(\cpu.intr.r_enable[4] ),
    .X(_09214_));
 sg13g2_buf_1 _15959_ (.A(ui_in[2]),
    .X(_09215_));
 sg13g2_nand2_1 _15960_ (.Y(_09216_),
    .A(\cpu.gpio.r_enable_in[2] ),
    .B(_09215_));
 sg13g2_buf_1 _15961_ (.A(ui_in[7]),
    .X(_09217_));
 sg13g2_nand2_1 _15962_ (.Y(_09218_),
    .A(\cpu.gpio.r_enable_in[7] ),
    .B(_09217_));
 sg13g2_buf_1 _15963_ (.A(\cpu.gpio.r_enable_in[0] ),
    .X(_09219_));
 sg13g2_buf_1 _15964_ (.A(ui_in[0]),
    .X(_09220_));
 sg13g2_buf_1 _15965_ (.A(\cpu.gpio.r_enable_in[6] ),
    .X(_09221_));
 sg13g2_buf_1 _15966_ (.A(ui_in[6]),
    .X(_09222_));
 sg13g2_a22oi_1 _15967_ (.Y(_09223_),
    .B1(_09221_),
    .B2(_09222_),
    .A2(_09220_),
    .A1(_09219_));
 sg13g2_and3_1 _15968_ (.X(_09224_),
    .A(_09216_),
    .B(_09218_),
    .C(_09223_));
 sg13g2_buf_1 _15969_ (.A(\cpu.gpio.r_enable_in[1] ),
    .X(_09225_));
 sg13g2_buf_1 _15970_ (.A(ui_in[1]),
    .X(_09226_));
 sg13g2_buf_1 _15971_ (.A(uio_in[7]),
    .X(_09227_));
 sg13g2_a22oi_1 _15972_ (.Y(_09228_),
    .B1(\cpu.gpio.r_enable_io[7] ),
    .B2(_09227_),
    .A2(_09226_),
    .A1(_09225_));
 sg13g2_buf_1 _15973_ (.A(\cpu.gpio.r_enable_in[3] ),
    .X(_09229_));
 sg13g2_buf_1 _15974_ (.A(ui_in[3]),
    .X(_09230_));
 sg13g2_buf_1 _15975_ (.A(uio_in[6]),
    .X(_09231_));
 sg13g2_a22oi_1 _15976_ (.Y(_09232_),
    .B1(\cpu.gpio.r_enable_io[6] ),
    .B2(_09231_),
    .A2(_09230_),
    .A1(_09229_));
 sg13g2_buf_1 _15977_ (.A(\cpu.gpio.r_enable_in[4] ),
    .X(_09233_));
 sg13g2_buf_1 _15978_ (.A(ui_in[4]),
    .X(_09234_));
 sg13g2_buf_1 _15979_ (.A(\cpu.gpio.r_enable_in[5] ),
    .X(_09235_));
 sg13g2_buf_1 _15980_ (.A(ui_in[5]),
    .X(_09236_));
 sg13g2_a22oi_1 _15981_ (.Y(_09237_),
    .B1(_09235_),
    .B2(_09236_),
    .A2(_09234_),
    .A1(_09233_));
 sg13g2_buf_1 _15982_ (.A(\cpu.gpio.r_enable_io[4] ),
    .X(_09238_));
 sg13g2_buf_1 _15983_ (.A(uio_in[4]),
    .X(_09239_));
 sg13g2_buf_1 _15984_ (.A(\cpu.gpio.r_enable_io[5] ),
    .X(_09240_));
 sg13g2_buf_1 _15985_ (.A(uio_in[5]),
    .X(_09241_));
 sg13g2_a22oi_1 _15986_ (.Y(_09242_),
    .B1(_09240_),
    .B2(_09241_),
    .A2(_09239_),
    .A1(_09238_));
 sg13g2_and4_1 _15987_ (.A(_09228_),
    .B(_09232_),
    .C(_09237_),
    .D(_09242_),
    .X(_09243_));
 sg13g2_nand2_1 _15988_ (.Y(_09244_),
    .A(_09224_),
    .B(_09243_));
 sg13g2_buf_1 _15989_ (.A(\cpu.intr.r_timer ),
    .X(_09245_));
 sg13g2_buf_1 _15990_ (.A(\cpu.intr.r_enable[3] ),
    .X(_09246_));
 sg13g2_a22oi_1 _15991_ (.Y(_09247_),
    .B1(_09246_),
    .B2(\cpu.intr.r_swi ),
    .A2(\cpu.intr.r_enable[2] ),
    .A1(_09245_));
 sg13g2_buf_1 _15992_ (.A(\cpu.uart.r_x_int ),
    .X(_09248_));
 sg13g2_buf_1 _15993_ (.A(\cpu.uart.r_r_int ),
    .X(_09249_));
 sg13g2_o21ai_1 _15994_ (.B1(\cpu.intr.r_enable[0] ),
    .Y(_09250_),
    .A1(_09248_),
    .A2(_09249_));
 sg13g2_buf_1 _15995_ (.A(\cpu.intr.r_enable[1] ),
    .X(_09251_));
 sg13g2_buf_1 _15996_ (.A(\cpu.intr.spi_intr ),
    .X(_09252_));
 sg13g2_buf_1 _15997_ (.A(\cpu.intr.r_enable[5] ),
    .X(_09253_));
 sg13g2_a22oi_1 _15998_ (.Y(_09254_),
    .B1(_09252_),
    .B2(_09253_),
    .A2(_09251_),
    .A1(\cpu.intr.r_clock ));
 sg13g2_nand3_1 _15999_ (.B(_09250_),
    .C(_09254_),
    .A(_09247_),
    .Y(_09255_));
 sg13g2_a21oi_1 _16000_ (.A1(_09214_),
    .A2(_09244_),
    .Y(_09256_),
    .B1(_09255_));
 sg13g2_buf_2 _16001_ (.A(\cpu.ex.r_ie ),
    .X(_09257_));
 sg13g2_nor2b_2 _16002_ (.A(_09256_),
    .B_N(_09257_),
    .Y(_09258_));
 sg13g2_nand2_1 _16003_ (.Y(_09259_),
    .A(net1127),
    .B(_09258_));
 sg13g2_nand4_1 _16004_ (.B(_09211_),
    .C(_09213_),
    .A(net1041),
    .Y(_09260_),
    .D(_09259_));
 sg13g2_buf_1 _16005_ (.A(_09260_),
    .X(_09261_));
 sg13g2_nor3_1 _16006_ (.A(net696),
    .B(_09208_),
    .C(_09261_),
    .Y(_09262_));
 sg13g2_buf_2 _16007_ (.A(_09262_),
    .X(_09263_));
 sg13g2_nor2_1 _16008_ (.A(_09196_),
    .B(_09263_),
    .Y(_09264_));
 sg13g2_buf_1 _16009_ (.A(_09264_),
    .X(_09265_));
 sg13g2_buf_2 _16010_ (.A(_09201_),
    .X(_09266_));
 sg13g2_buf_2 _16011_ (.A(\cpu.addr[2] ),
    .X(_09267_));
 sg13g2_buf_1 _16012_ (.A(_09267_),
    .X(_09268_));
 sg13g2_buf_1 _16013_ (.A(net1040),
    .X(_09269_));
 sg13g2_buf_1 _16014_ (.A(net901),
    .X(_09270_));
 sg13g2_buf_2 _16015_ (.A(\cpu.addr[1] ),
    .X(_09271_));
 sg13g2_buf_1 _16016_ (.A(_09271_),
    .X(_09272_));
 sg13g2_buf_1 _16017_ (.A(_09272_),
    .X(_09273_));
 sg13g2_nand2_1 _16018_ (.Y(_09274_),
    .A(_09213_),
    .B(_09259_));
 sg13g2_or4_1 _16019_ (.A(_00197_),
    .B(net783),
    .C(_09273_),
    .D(_09274_),
    .X(_09275_));
 sg13g2_inv_1 _16020_ (.Y(_09276_),
    .A(_08580_));
 sg13g2_nor2_1 _16021_ (.A(net1126),
    .B(_08580_),
    .Y(_09277_));
 sg13g2_a21oi_1 _16022_ (.A1(net1126),
    .A2(net1060),
    .Y(_09278_),
    .B1(_09277_));
 sg13g2_nand2_1 _16023_ (.Y(_09279_),
    .A(net1125),
    .B(_09278_));
 sg13g2_o21ai_1 _16024_ (.B1(_09279_),
    .Y(_09280_),
    .A1(_09276_),
    .A2(net1060));
 sg13g2_buf_1 _16025_ (.A(_09280_),
    .X(_09281_));
 sg13g2_nor4_2 _16026_ (.A(net632),
    .B(_09208_),
    .C(_09275_),
    .Y(_09282_),
    .D(_09281_));
 sg13g2_buf_1 _16027_ (.A(\cpu.spi.r_state[3] ),
    .X(_09283_));
 sg13g2_a21oi_1 _16028_ (.A1(_09265_),
    .A2(_09282_),
    .Y(_09284_),
    .B1(_09283_));
 sg13g2_buf_2 _16029_ (.A(\cpu.spi.r_state[0] ),
    .X(_09285_));
 sg13g2_buf_1 _16030_ (.A(net783),
    .X(_09286_));
 sg13g2_buf_1 _16031_ (.A(net900),
    .X(_09287_));
 sg13g2_nor2_1 _16032_ (.A(net695),
    .B(net782),
    .Y(_09288_));
 sg13g2_buf_2 _16033_ (.A(_09288_),
    .X(_09289_));
 sg13g2_nand2_1 _16034_ (.Y(_09290_),
    .A(_09263_),
    .B(_09289_));
 sg13g2_nand2b_1 _16035_ (.Y(_09291_),
    .B(net1),
    .A_N(r_reset));
 sg13g2_buf_2 _16036_ (.A(_09291_),
    .X(_09292_));
 sg13g2_buf_1 _16037_ (.A(_09292_),
    .X(_09293_));
 sg13g2_buf_2 _16038_ (.A(net899),
    .X(_09294_));
 sg13g2_a21oi_1 _16039_ (.A1(_09285_),
    .A2(_09290_),
    .Y(_09295_),
    .B1(net781));
 sg13g2_o21ai_1 _16040_ (.B1(_09295_),
    .Y(_00029_),
    .A1(_09194_),
    .A2(_09284_));
 sg13g2_buf_2 _16041_ (.A(net781),
    .X(_09296_));
 sg13g2_buf_1 _16042_ (.A(_09296_),
    .X(_09297_));
 sg13g2_inv_1 _16043_ (.Y(_09298_),
    .A(_09282_));
 sg13g2_buf_1 _16044_ (.A(\cpu.spi.r_bits[0] ),
    .X(_09299_));
 sg13g2_buf_1 _16045_ (.A(\cpu.spi.r_bits[1] ),
    .X(_09300_));
 sg13g2_nor3_1 _16046_ (.A(_09299_),
    .B(_09300_),
    .C(\cpu.spi.r_bits[2] ),
    .Y(_09301_));
 sg13g2_buf_1 _16047_ (.A(\cpu.spi.r_timeout_count[7] ),
    .X(_09302_));
 sg13g2_buf_1 _16048_ (.A(\cpu.spi.r_timeout_count[0] ),
    .X(_09303_));
 sg13g2_buf_1 _16049_ (.A(\cpu.spi.r_timeout_count[1] ),
    .X(_09304_));
 sg13g2_or3_1 _16050_ (.A(_09303_),
    .B(_09304_),
    .C(\cpu.spi.r_timeout_count[2] ),
    .X(_09305_));
 sg13g2_buf_1 _16051_ (.A(_09305_),
    .X(_09306_));
 sg13g2_or2_1 _16052_ (.X(_09307_),
    .B(_09306_),
    .A(\cpu.spi.r_timeout_count[3] ));
 sg13g2_buf_1 _16053_ (.A(_09307_),
    .X(_09308_));
 sg13g2_or2_1 _16054_ (.X(_09309_),
    .B(_09308_),
    .A(\cpu.spi.r_timeout_count[4] ));
 sg13g2_buf_1 _16055_ (.A(_09309_),
    .X(_09310_));
 sg13g2_or2_1 _16056_ (.X(_09311_),
    .B(_09310_),
    .A(\cpu.spi.r_timeout_count[5] ));
 sg13g2_buf_1 _16057_ (.A(_09311_),
    .X(_09312_));
 sg13g2_or2_1 _16058_ (.X(_09313_),
    .B(_09312_),
    .A(\cpu.spi.r_timeout_count[6] ));
 sg13g2_buf_1 _16059_ (.A(_09313_),
    .X(_09314_));
 sg13g2_o21ai_1 _16060_ (.B1(\cpu.spi.r_searching ),
    .Y(_09315_),
    .A1(_09302_),
    .A2(_09314_));
 sg13g2_nand2_1 _16061_ (.Y(_09316_),
    .A(_09301_),
    .B(_09315_));
 sg13g2_buf_1 _16062_ (.A(\cpu.spi.r_in[3] ),
    .X(_09317_));
 sg13g2_buf_1 _16063_ (.A(\cpu.spi.r_in[6] ),
    .X(_09318_));
 sg13g2_buf_1 _16064_ (.A(\cpu.spi.r_in[1] ),
    .X(_09319_));
 sg13g2_buf_1 _16065_ (.A(\cpu.spi.r_in[0] ),
    .X(_09320_));
 sg13g2_nand2_1 _16066_ (.Y(_09321_),
    .A(_09319_),
    .B(_09320_));
 sg13g2_nand3_1 _16067_ (.B(_09318_),
    .C(_09321_),
    .A(_09317_),
    .Y(_09322_));
 sg13g2_buf_1 _16068_ (.A(\cpu.spi.r_in[2] ),
    .X(_09323_));
 sg13g2_buf_1 _16069_ (.A(\cpu.spi.r_in[5] ),
    .X(_09324_));
 sg13g2_buf_1 _16070_ (.A(\cpu.spi.r_in[4] ),
    .X(_09325_));
 sg13g2_nand4_1 _16071_ (.B(_09324_),
    .C(_09325_),
    .A(_09323_),
    .Y(_09326_),
    .D(\cpu.spi.r_in[7] ));
 sg13g2_nor2_1 _16072_ (.A(_09322_),
    .B(_09326_),
    .Y(_09327_));
 sg13g2_o21ai_1 _16073_ (.B1(\cpu.spi.r_searching ),
    .Y(_09328_),
    .A1(_00220_),
    .A2(_09327_));
 sg13g2_buf_1 _16074_ (.A(_09328_),
    .X(_09329_));
 sg13g2_a21oi_1 _16075_ (.A1(_09316_),
    .A2(_09329_),
    .Y(_09330_),
    .B1(_09193_));
 sg13g2_buf_1 _16076_ (.A(\cpu.spi.r_state[6] ),
    .X(_09331_));
 sg13g2_buf_1 _16077_ (.A(_09331_),
    .X(_09332_));
 sg13g2_a22oi_1 _16078_ (.Y(_09333_),
    .B1(_09330_),
    .B2(net1038),
    .A2(_09298_),
    .A1(_09265_));
 sg13g2_nor2_1 _16079_ (.A(net631),
    .B(_09333_),
    .Y(_00030_));
 sg13g2_nor2b_1 _16080_ (.A(_09183_),
    .B_N(_09191_),
    .Y(_09334_));
 sg13g2_buf_1 _16081_ (.A(_09334_),
    .X(_09335_));
 sg13g2_buf_1 _16082_ (.A(net473),
    .X(_09336_));
 sg13g2_nand4_1 _16083_ (.B(net418),
    .C(_09316_),
    .A(net1038),
    .Y(_09337_),
    .D(_09329_));
 sg13g2_buf_1 _16084_ (.A(_09337_),
    .X(_09338_));
 sg13g2_buf_1 _16085_ (.A(\cpu.spi.r_state[2] ),
    .X(_09339_));
 sg13g2_buf_1 _16086_ (.A(_09196_),
    .X(_09340_));
 sg13g2_inv_2 _16087_ (.Y(_09341_),
    .A(net1044));
 sg13g2_buf_1 _16088_ (.A(_09341_),
    .X(_09342_));
 sg13g2_nor2_1 _16089_ (.A(_09208_),
    .B(_09261_),
    .Y(_09343_));
 sg13g2_buf_2 _16090_ (.A(_09343_),
    .X(_09344_));
 sg13g2_nand2_1 _16091_ (.Y(_09345_),
    .A(net780),
    .B(_09344_));
 sg13g2_buf_1 _16092_ (.A(_09345_),
    .X(_09346_));
 sg13g2_buf_1 _16093_ (.A(\cpu.spi.r_state[4] ),
    .X(_09347_));
 sg13g2_nor3_1 _16094_ (.A(\cpu.spi.r_state[5] ),
    .B(net1121),
    .C(net419),
    .Y(_09348_));
 sg13g2_o21ai_1 _16095_ (.B1(_09348_),
    .Y(_09349_),
    .A1(net898),
    .A2(net117));
 sg13g2_o21ai_1 _16096_ (.B1(_09349_),
    .Y(_09350_),
    .A1(net1122),
    .A2(_09336_));
 sg13g2_buf_2 _16097_ (.A(net781),
    .X(_09351_));
 sg13g2_buf_1 _16098_ (.A(_09351_),
    .X(_09352_));
 sg13g2_a21oi_1 _16099_ (.A1(_09338_),
    .A2(_09350_),
    .Y(_00031_),
    .B1(net630));
 sg13g2_buf_1 _16100_ (.A(_09351_),
    .X(_09353_));
 sg13g2_nor3_1 _16101_ (.A(_09353_),
    .B(_09336_),
    .C(_09284_),
    .Y(_00032_));
 sg13g2_buf_1 _16102_ (.A(_09263_),
    .X(_09354_));
 sg13g2_nand3_1 _16103_ (.B(net143),
    .C(_09289_),
    .A(_09285_),
    .Y(_09355_));
 sg13g2_nand2_1 _16104_ (.Y(_09356_),
    .A(net1121),
    .B(net419));
 sg13g2_a21oi_1 _16105_ (.A1(_09355_),
    .A2(_09356_),
    .Y(_00033_),
    .B1(net630));
 sg13g2_buf_1 _16106_ (.A(_09195_),
    .X(_09357_));
 sg13g2_buf_1 _16107_ (.A(net1037),
    .X(_09358_));
 sg13g2_a21oi_1 _16108_ (.A1(_09358_),
    .A2(net143),
    .Y(_09359_),
    .B1(\cpu.spi.r_state[5] ));
 sg13g2_nor3_1 _16109_ (.A(net629),
    .B(net418),
    .C(_09359_),
    .Y(_00034_));
 sg13g2_nand2_1 _16110_ (.Y(_09360_),
    .A(net1038),
    .B(net419));
 sg13g2_nand2_1 _16111_ (.Y(_09361_),
    .A(net1122),
    .B(net418));
 sg13g2_a21oi_1 _16112_ (.A1(_09360_),
    .A2(_09361_),
    .Y(_00035_),
    .B1(net630));
 sg13g2_buf_2 _16113_ (.A(\cpu.ex.r_mult_off[0] ),
    .X(_09362_));
 sg13g2_inv_1 _16114_ (.Y(_09363_),
    .A(\cpu.dec.mult ));
 sg13g2_nand3b_1 _16115_ (.B(\cpu.dec.iready ),
    .C(_00199_),
    .Y(_09364_),
    .A_N(\cpu.ex.r_branch_stall ));
 sg13g2_buf_1 _16116_ (.A(_09364_),
    .X(_09365_));
 sg13g2_nor3_1 _16117_ (.A(_09363_),
    .B(_09292_),
    .C(net1036),
    .Y(_09366_));
 sg13g2_buf_2 _16118_ (.A(_09366_),
    .X(_09367_));
 sg13g2_inv_1 _16119_ (.Y(_09368_),
    .A(\cpu.dec.div ));
 sg13g2_nor3_1 _16120_ (.A(_09368_),
    .B(_09292_),
    .C(net1036),
    .Y(_09369_));
 sg13g2_buf_2 _16121_ (.A(_09369_),
    .X(_09370_));
 sg13g2_nor2_2 _16122_ (.A(_09367_),
    .B(_09370_),
    .Y(_09371_));
 sg13g2_nand2_1 _16123_ (.Y(_09372_),
    .A(_09362_),
    .B(_09371_));
 sg13g2_buf_2 _16124_ (.A(_09372_),
    .X(\cpu.ex.c_mult_off[0] ));
 sg13g2_buf_1 _16125_ (.A(\cpu.ex.r_div_running ),
    .X(_09373_));
 sg13g2_buf_2 _16126_ (.A(\cpu.ex.r_mult_off[1] ),
    .X(_09374_));
 sg13g2_buf_2 _16127_ (.A(\cpu.ex.r_mult_off[2] ),
    .X(_09375_));
 sg13g2_buf_2 _16128_ (.A(\cpu.ex.r_mult_off[3] ),
    .X(_09376_));
 sg13g2_nor4_2 _16129_ (.A(_09374_),
    .B(_09375_),
    .C(_09376_),
    .Y(_09377_),
    .D(\cpu.ex.c_mult_off[0] ));
 sg13g2_buf_1 _16130_ (.A(_09370_),
    .X(_09378_));
 sg13g2_buf_1 _16131_ (.A(net694),
    .X(_09379_));
 sg13g2_nor2b_1 _16132_ (.A(r_reset),
    .B_N(net1),
    .Y(_09380_));
 sg13g2_buf_1 _16133_ (.A(_09380_),
    .X(_09381_));
 sg13g2_o21ai_1 _16134_ (.B1(_09381_),
    .Y(_09382_),
    .A1(_09373_),
    .A2(net628));
 sg13g2_a21oi_1 _16135_ (.A1(_09373_),
    .A2(_09377_),
    .Y(\cpu.ex.c_div_running ),
    .B1(_09382_));
 sg13g2_buf_1 _16136_ (.A(\cpu.ex.r_mult_running ),
    .X(_09383_));
 sg13g2_or3_1 _16137_ (.A(_09363_),
    .B(_09292_),
    .C(net1036),
    .X(_09384_));
 sg13g2_buf_1 _16138_ (.A(_09384_),
    .X(_09385_));
 sg13g2_buf_8 _16139_ (.A(_09385_),
    .X(_09386_));
 sg13g2_nand2b_1 _16140_ (.Y(_09387_),
    .B(net693),
    .A_N(net1120));
 sg13g2_buf_2 _16141_ (.A(_09387_),
    .X(_09388_));
 sg13g2_nand2_1 _16142_ (.Y(_09389_),
    .A(_09381_),
    .B(_09388_));
 sg13g2_a21oi_1 _16143_ (.A1(net1120),
    .A2(_09377_),
    .Y(\cpu.ex.c_mult_running ),
    .B1(_09389_));
 sg13g2_buf_1 _16144_ (.A(\cpu.qspi.r_state[17] ),
    .X(_09390_));
 sg13g2_buf_1 _16145_ (.A(\cpu.dcache.flush_write ),
    .X(_09391_));
 sg13g2_buf_2 _16146_ (.A(\cpu.addr[4] ),
    .X(_09392_));
 sg13g2_and2_1 _16147_ (.A(_09392_),
    .B(_09197_),
    .X(_09393_));
 sg13g2_buf_1 _16148_ (.A(_09393_),
    .X(_09394_));
 sg13g2_and2_1 _16149_ (.A(net1040),
    .B(_09394_),
    .X(_09395_));
 sg13g2_buf_1 _16150_ (.A(_09395_),
    .X(_09396_));
 sg13g2_buf_1 _16151_ (.A(_09396_),
    .X(_09397_));
 sg13g2_buf_1 _16152_ (.A(_00225_),
    .X(_09398_));
 sg13g2_nand2_1 _16153_ (.Y(_09399_),
    .A(_09267_),
    .B(net1119));
 sg13g2_nor2_1 _16154_ (.A(_09198_),
    .B(_09399_),
    .Y(_09400_));
 sg13g2_buf_1 _16155_ (.A(_09400_),
    .X(_09401_));
 sg13g2_buf_1 _16156_ (.A(_09401_),
    .X(_09402_));
 sg13g2_buf_1 _16157_ (.A(net692),
    .X(_09403_));
 sg13g2_a22oi_1 _16158_ (.Y(_09404_),
    .B1(net626),
    .B2(\cpu.dcache.r_tag[1][12] ),
    .A2(net627),
    .A1(\cpu.dcache.r_tag[7][12] ));
 sg13g2_nor2b_1 _16159_ (.A(_09267_),
    .B_N(_00225_),
    .Y(_09405_));
 sg13g2_and2_1 _16160_ (.A(net1044),
    .B(_09405_),
    .X(_09406_));
 sg13g2_buf_1 _16161_ (.A(_09406_),
    .X(_09407_));
 sg13g2_buf_1 _16162_ (.A(_09407_),
    .X(_09408_));
 sg13g2_buf_1 _16163_ (.A(net691),
    .X(_09409_));
 sg13g2_and3_1 _16164_ (.X(_09410_),
    .A(net1040),
    .B(net1044),
    .C(net1119));
 sg13g2_buf_1 _16165_ (.A(_09410_),
    .X(_09411_));
 sg13g2_buf_1 _16166_ (.A(_09411_),
    .X(_09412_));
 sg13g2_buf_1 _16167_ (.A(net690),
    .X(_09413_));
 sg13g2_a22oi_1 _16168_ (.Y(_09414_),
    .B1(net624),
    .B2(\cpu.dcache.r_tag[3][12] ),
    .A2(net625),
    .A1(\cpu.dcache.r_tag[2][12] ));
 sg13g2_nor2b_1 _16169_ (.A(_09267_),
    .B_N(_09392_),
    .Y(_09415_));
 sg13g2_buf_2 _16170_ (.A(_09415_),
    .X(_09416_));
 sg13g2_and2_1 _16171_ (.A(net1044),
    .B(_09416_),
    .X(_09417_));
 sg13g2_buf_2 _16172_ (.A(_09417_),
    .X(_09418_));
 sg13g2_buf_1 _16173_ (.A(net689),
    .X(_09419_));
 sg13g2_nor2b_1 _16174_ (.A(_09197_),
    .B_N(_09267_),
    .Y(_09420_));
 sg13g2_buf_2 _16175_ (.A(_09420_),
    .X(_09421_));
 sg13g2_and2_1 _16176_ (.A(_09392_),
    .B(_09421_),
    .X(_09422_));
 sg13g2_buf_1 _16177_ (.A(_09422_),
    .X(_09423_));
 sg13g2_buf_2 _16178_ (.A(_09423_),
    .X(_09424_));
 sg13g2_a22oi_1 _16179_ (.Y(_09425_),
    .B1(net622),
    .B2(\cpu.dcache.r_tag[5][12] ),
    .A2(net623),
    .A1(\cpu.dcache.r_tag[6][12] ));
 sg13g2_inv_1 _16180_ (.Y(_09426_),
    .A(_00241_));
 sg13g2_nor2_1 _16181_ (.A(_09392_),
    .B(_09197_),
    .Y(_09427_));
 sg13g2_and2_1 _16182_ (.A(_09399_),
    .B(_09427_),
    .X(_09428_));
 sg13g2_buf_2 _16183_ (.A(_09428_),
    .X(_09429_));
 sg13g2_buf_1 _16184_ (.A(_09429_),
    .X(_09430_));
 sg13g2_and2_1 _16185_ (.A(_09341_),
    .B(_09416_),
    .X(_09431_));
 sg13g2_buf_2 _16186_ (.A(_09431_),
    .X(_09432_));
 sg13g2_buf_1 _16187_ (.A(_09432_),
    .X(_09433_));
 sg13g2_a22oi_1 _16188_ (.Y(_09434_),
    .B1(net621),
    .B2(\cpu.dcache.r_tag[4][12] ),
    .A2(net688),
    .A1(_09426_));
 sg13g2_nand4_1 _16189_ (.B(_09414_),
    .C(_09425_),
    .A(_09404_),
    .Y(_09435_),
    .D(_09434_));
 sg13g2_buf_1 _16190_ (.A(_08504_),
    .X(_09436_));
 sg13g2_buf_4 _16191_ (.X(_09437_),
    .A(_08481_));
 sg13g2_buf_8 _16192_ (.A(_09437_),
    .X(_09438_));
 sg13g2_buf_8 _16193_ (.A(_08495_),
    .X(_09439_));
 sg13g2_buf_1 _16194_ (.A(_09439_),
    .X(_09440_));
 sg13g2_mux4_1 _16195_ (.S0(net779),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .S1(net778),
    .X(_09441_));
 sg13g2_buf_1 _16196_ (.A(_09439_),
    .X(_09442_));
 sg13g2_mux4_1 _16197_ (.S0(net779),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .S1(net777),
    .X(_09443_));
 sg13g2_mux4_1 _16198_ (.S0(_09438_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .S1(_09440_),
    .X(_09444_));
 sg13g2_mux4_1 _16199_ (.S0(net779),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .S1(net778),
    .X(_09445_));
 sg13g2_buf_2 _16200_ (.A(_08472_),
    .X(_09446_));
 sg13g2_buf_2 _16201_ (.A(net922),
    .X(_09447_));
 sg13g2_mux4_1 _16202_ (.S0(net776),
    .A0(_09441_),
    .A1(_09443_),
    .A2(_09444_),
    .A3(_09445_),
    .S1(net775),
    .X(_09448_));
 sg13g2_buf_1 _16203_ (.A(_08478_),
    .X(_09449_));
 sg13g2_buf_2 _16204_ (.A(_09439_),
    .X(_09450_));
 sg13g2_mux4_1 _16205_ (.S0(_09437_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .S1(net774),
    .X(_09451_));
 sg13g2_buf_2 _16206_ (.A(_08481_),
    .X(_09452_));
 sg13g2_mux4_1 _16207_ (.S0(net896),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .S1(net774),
    .X(_09453_));
 sg13g2_mux4_1 _16208_ (.S0(_09437_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .S1(_09439_),
    .X(_09454_));
 sg13g2_mux4_1 _16209_ (.S0(_09437_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .S1(net774),
    .X(_09455_));
 sg13g2_buf_2 _16210_ (.A(_08472_),
    .X(_09456_));
 sg13g2_mux4_1 _16211_ (.S0(net773),
    .A0(_09451_),
    .A1(_09453_),
    .A2(_09454_),
    .A3(_09455_),
    .S1(net922),
    .X(_09457_));
 sg13g2_and2_1 _16212_ (.A(net686),
    .B(_09457_),
    .X(_09458_));
 sg13g2_a21oi_1 _16213_ (.A1(net687),
    .A2(_09448_),
    .Y(_09459_),
    .B1(_09458_));
 sg13g2_buf_8 _16214_ (.A(net779),
    .X(_09460_));
 sg13g2_buf_1 _16215_ (.A(net685),
    .X(_09461_));
 sg13g2_nor2_1 _16216_ (.A(net1129),
    .B(_09461_),
    .Y(_09462_));
 sg13g2_a21oi_1 _16217_ (.A1(net1057),
    .A2(_09459_),
    .Y(_09463_),
    .B1(_09462_));
 sg13g2_buf_1 _16218_ (.A(_09463_),
    .X(_09464_));
 sg13g2_xor2_1 _16219_ (.B(net382),
    .A(_09435_),
    .X(_09465_));
 sg13g2_a22oi_1 _16220_ (.Y(_09466_),
    .B1(net623),
    .B2(\cpu.dcache.r_tag[6][13] ),
    .A2(net692),
    .A1(\cpu.dcache.r_tag[1][13] ));
 sg13g2_a22oi_1 _16221_ (.Y(_09467_),
    .B1(net624),
    .B2(\cpu.dcache.r_tag[3][13] ),
    .A2(net625),
    .A1(\cpu.dcache.r_tag[2][13] ));
 sg13g2_a22oi_1 _16222_ (.Y(_09468_),
    .B1(net622),
    .B2(\cpu.dcache.r_tag[5][13] ),
    .A2(net627),
    .A1(\cpu.dcache.r_tag[7][13] ));
 sg13g2_inv_1 _16223_ (.Y(_09469_),
    .A(_00242_));
 sg13g2_a22oi_1 _16224_ (.Y(_09470_),
    .B1(net621),
    .B2(\cpu.dcache.r_tag[4][13] ),
    .A2(net688),
    .A1(_09469_));
 sg13g2_nand4_1 _16225_ (.B(_09467_),
    .C(_09468_),
    .A(_09466_),
    .Y(_09471_),
    .D(_09470_));
 sg13g2_buf_8 _16226_ (.A(_09437_),
    .X(_09472_));
 sg13g2_buf_2 _16227_ (.A(_09439_),
    .X(_09473_));
 sg13g2_mux4_1 _16228_ (.S0(net772),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .S1(net771),
    .X(_09474_));
 sg13g2_mux4_1 _16229_ (.S0(net772),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .S1(net771),
    .X(_09475_));
 sg13g2_buf_2 _16230_ (.A(_09439_),
    .X(_09476_));
 sg13g2_mux4_1 _16231_ (.S0(net896),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .S1(net770),
    .X(_09477_));
 sg13g2_buf_8 _16232_ (.A(_09437_),
    .X(_09478_));
 sg13g2_mux4_1 _16233_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .S1(net770),
    .X(_09479_));
 sg13g2_mux4_1 _16234_ (.S0(net773),
    .A0(_09474_),
    .A1(_09475_),
    .A2(_09477_),
    .A3(_09479_),
    .S1(net922),
    .X(_09480_));
 sg13g2_mux4_1 _16235_ (.S0(_09478_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .S1(_09476_),
    .X(_09481_));
 sg13g2_mux4_1 _16236_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .S1(net770),
    .X(_09482_));
 sg13g2_mux4_1 _16237_ (.S0(net896),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .S1(net774),
    .X(_09483_));
 sg13g2_mux4_1 _16238_ (.S0(net896),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .S1(net774),
    .X(_09484_));
 sg13g2_mux4_1 _16239_ (.S0(net773),
    .A0(_09481_),
    .A1(_09482_),
    .A2(_09483_),
    .A3(_09484_),
    .S1(net922),
    .X(_09485_));
 sg13g2_mux2_1 _16240_ (.A0(_09480_),
    .A1(_09485_),
    .S(net687),
    .X(_09486_));
 sg13g2_nand2_1 _16241_ (.Y(_09487_),
    .A(_08463_),
    .B(_09486_));
 sg13g2_o21ai_1 _16242_ (.B1(_09487_),
    .Y(_09488_),
    .A1(_08619_),
    .A2(_08489_));
 sg13g2_buf_1 _16243_ (.A(_09488_),
    .X(_09489_));
 sg13g2_xor2_1 _16244_ (.B(net381),
    .A(_09471_),
    .X(_09490_));
 sg13g2_nor2_1 _16245_ (.A(_09465_),
    .B(_09490_),
    .Y(_09491_));
 sg13g2_inv_1 _16246_ (.Y(_09492_),
    .A(_09491_));
 sg13g2_buf_8 _16247_ (.A(net779),
    .X(_09493_));
 sg13g2_buf_2 _16248_ (.A(net778),
    .X(_09494_));
 sg13g2_mux4_1 _16249_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .S1(net683),
    .X(_09495_));
 sg13g2_buf_8 _16250_ (.A(net779),
    .X(_09496_));
 sg13g2_buf_2 _16251_ (.A(net778),
    .X(_09497_));
 sg13g2_mux4_1 _16252_ (.S0(net682),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .S1(net681),
    .X(_09498_));
 sg13g2_buf_8 _16253_ (.A(_09437_),
    .X(_09499_));
 sg13g2_buf_8 _16254_ (.A(net768),
    .X(_09500_));
 sg13g2_buf_2 _16255_ (.A(net778),
    .X(_09501_));
 sg13g2_mux4_1 _16256_ (.S0(net680),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .S1(net679),
    .X(_09502_));
 sg13g2_mux4_1 _16257_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .S1(net683),
    .X(_09503_));
 sg13g2_mux4_1 _16258_ (.S0(net776),
    .A0(_09495_),
    .A1(_09498_),
    .A2(_09502_),
    .A3(_09503_),
    .S1(net775),
    .X(_09504_));
 sg13g2_nand2_1 _16259_ (.Y(_09505_),
    .A(net686),
    .B(_09504_));
 sg13g2_mux4_1 _16260_ (.S0(_09493_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .S1(_09494_),
    .X(_09506_));
 sg13g2_mux4_1 _16261_ (.S0(_09493_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .S1(_09494_),
    .X(_09507_));
 sg13g2_mux4_1 _16262_ (.S0(net680),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .S1(net679),
    .X(_09508_));
 sg13g2_mux4_1 _16263_ (.S0(net680),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .S1(net679),
    .X(_09509_));
 sg13g2_mux4_1 _16264_ (.S0(net776),
    .A0(_09506_),
    .A1(_09507_),
    .A2(_09508_),
    .A3(_09509_),
    .S1(net775),
    .X(_09510_));
 sg13g2_nand2_1 _16265_ (.Y(_09511_),
    .A(net687),
    .B(_09510_));
 sg13g2_a21oi_1 _16266_ (.A1(_09505_),
    .A2(_09511_),
    .Y(_09512_),
    .B1(_08694_));
 sg13g2_buf_1 _16267_ (.A(_09512_),
    .X(_09513_));
 sg13g2_inv_1 _16268_ (.Y(_09514_),
    .A(_00246_));
 sg13g2_buf_1 _16269_ (.A(_09427_),
    .X(_09515_));
 sg13g2_nand2_1 _16270_ (.Y(_09516_),
    .A(_09399_),
    .B(net895));
 sg13g2_buf_2 _16271_ (.A(_09516_),
    .X(_09517_));
 sg13g2_a22oi_1 _16272_ (.Y(_09518_),
    .B1(net622),
    .B2(\cpu.dcache.r_tag[5][17] ),
    .A2(net692),
    .A1(\cpu.dcache.r_tag[1][17] ));
 sg13g2_a22oi_1 _16273_ (.Y(_09519_),
    .B1(net624),
    .B2(\cpu.dcache.r_tag[3][17] ),
    .A2(net625),
    .A1(\cpu.dcache.r_tag[2][17] ));
 sg13g2_and2_1 _16274_ (.A(net1040),
    .B(net1044),
    .X(_09520_));
 sg13g2_buf_2 _16275_ (.A(_09520_),
    .X(_09521_));
 sg13g2_mux2_1 _16276_ (.A0(\cpu.dcache.r_tag[4][17] ),
    .A1(\cpu.dcache.r_tag[6][17] ),
    .S(net902),
    .X(_09522_));
 sg13g2_inv_1 _16277_ (.Y(_09523_),
    .A(net1040));
 sg13g2_buf_1 _16278_ (.A(_09523_),
    .X(_09524_));
 sg13g2_a22oi_1 _16279_ (.Y(_09525_),
    .B1(_09522_),
    .B2(_09524_),
    .A2(_09521_),
    .A1(\cpu.dcache.r_tag[7][17] ));
 sg13g2_buf_1 _16280_ (.A(_09392_),
    .X(_09526_));
 sg13g2_nand2b_1 _16281_ (.Y(_09527_),
    .B(_09526_),
    .A_N(_09525_));
 sg13g2_nand4_1 _16282_ (.B(_09518_),
    .C(_09519_),
    .A(_09517_),
    .Y(_09528_),
    .D(_09527_));
 sg13g2_o21ai_1 _16283_ (.B1(_09528_),
    .Y(_09529_),
    .A1(_09514_),
    .A2(_09517_));
 sg13g2_xor2_1 _16284_ (.B(_09529_),
    .A(net380),
    .X(_09530_));
 sg13g2_a22oi_1 _16285_ (.Y(_09531_),
    .B1(net621),
    .B2(\cpu.dcache.r_tag[4][14] ),
    .A2(net626),
    .A1(\cpu.dcache.r_tag[1][14] ));
 sg13g2_a22oi_1 _16286_ (.Y(_09532_),
    .B1(net624),
    .B2(\cpu.dcache.r_tag[3][14] ),
    .A2(net625),
    .A1(\cpu.dcache.r_tag[2][14] ));
 sg13g2_buf_1 _16287_ (.A(net622),
    .X(_09533_));
 sg13g2_a22oi_1 _16288_ (.Y(_09534_),
    .B1(net541),
    .B2(\cpu.dcache.r_tag[5][14] ),
    .A2(net623),
    .A1(\cpu.dcache.r_tag[6][14] ));
 sg13g2_inv_1 _16289_ (.Y(_09535_),
    .A(_00243_));
 sg13g2_a22oi_1 _16290_ (.Y(_09536_),
    .B1(net688),
    .B2(_09535_),
    .A2(net627),
    .A1(\cpu.dcache.r_tag[7][14] ));
 sg13g2_nand4_1 _16291_ (.B(_09532_),
    .C(_09534_),
    .A(_09531_),
    .Y(_09537_),
    .D(_09536_));
 sg13g2_buf_2 _16292_ (.A(net775),
    .X(_09538_));
 sg13g2_buf_2 _16293_ (.A(_09437_),
    .X(_09539_));
 sg13g2_mux4_1 _16294_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .S1(net777),
    .X(_09540_));
 sg13g2_mux4_1 _16295_ (.S0(net680),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .S1(net679),
    .X(_09541_));
 sg13g2_mux4_1 _16296_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .S1(net777),
    .X(_09542_));
 sg13g2_mux4_1 _16297_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .S1(net777),
    .X(_09543_));
 sg13g2_mux4_1 _16298_ (.S0(_08504_),
    .A0(_09540_),
    .A1(_09541_),
    .A2(_09542_),
    .A3(_09543_),
    .S1(net1059),
    .X(_09544_));
 sg13g2_nand2_1 _16299_ (.Y(_09545_),
    .A(_08619_),
    .B(_09544_));
 sg13g2_mux4_1 _16300_ (.S0(net680),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .S1(net679),
    .X(_09546_));
 sg13g2_mux4_1 _16301_ (.S0(net680),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .S1(net679),
    .X(_09547_));
 sg13g2_mux4_1 _16302_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .S1(net777),
    .X(_09548_));
 sg13g2_mux4_1 _16303_ (.S0(_09539_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .S1(_09442_),
    .X(_09549_));
 sg13g2_mux4_1 _16304_ (.S0(_08504_),
    .A0(_09546_),
    .A1(_09547_),
    .A2(_09548_),
    .A3(_09549_),
    .S1(_08588_),
    .X(_09550_));
 sg13g2_o21ai_1 _16305_ (.B1(net678),
    .Y(_09551_),
    .A1(_08464_),
    .A2(_09550_));
 sg13g2_o21ai_1 _16306_ (.B1(_09551_),
    .Y(_09552_),
    .A1(net678),
    .A2(_09545_));
 sg13g2_buf_1 _16307_ (.A(_09552_),
    .X(_09553_));
 sg13g2_xnor2_1 _16308_ (.Y(_09554_),
    .A(_09537_),
    .B(net379));
 sg13g2_buf_1 _16309_ (.A(net1035),
    .X(_09555_));
 sg13g2_mux2_1 _16310_ (.A0(\cpu.dcache.r_tag[5][11] ),
    .A1(\cpu.dcache.r_tag[7][11] ),
    .S(net902),
    .X(_09556_));
 sg13g2_nor2_2 _16311_ (.A(net901),
    .B(net902),
    .Y(_09557_));
 sg13g2_a22oi_1 _16312_ (.Y(_09558_),
    .B1(_09557_),
    .B2(\cpu.dcache.r_tag[4][11] ),
    .A2(_09556_),
    .A1(net901));
 sg13g2_inv_1 _16313_ (.Y(_09559_),
    .A(_09558_));
 sg13g2_a22oi_1 _16314_ (.Y(_09560_),
    .B1(net690),
    .B2(\cpu.dcache.r_tag[3][11] ),
    .A2(net691),
    .A1(\cpu.dcache.r_tag[2][11] ));
 sg13g2_nand2_1 _16315_ (.Y(_09561_),
    .A(\cpu.dcache.r_tag[1][11] ),
    .B(_09401_));
 sg13g2_inv_1 _16316_ (.Y(_09562_),
    .A(_00240_));
 sg13g2_a22oi_1 _16317_ (.Y(_09563_),
    .B1(_09429_),
    .B2(_09562_),
    .A2(net689),
    .A1(\cpu.dcache.r_tag[6][11] ));
 sg13g2_nand3_1 _16318_ (.B(_09561_),
    .C(_09563_),
    .A(_09560_),
    .Y(_09564_));
 sg13g2_a21oi_1 _16319_ (.A1(net894),
    .A2(_09559_),
    .Y(_09565_),
    .B1(_09564_));
 sg13g2_xor2_1 _16320_ (.B(_09565_),
    .A(_00239_),
    .X(_09566_));
 sg13g2_buf_2 _16321_ (.A(_00227_),
    .X(_09567_));
 sg13g2_inv_1 _16322_ (.Y(_09568_),
    .A(_09567_));
 sg13g2_a22oi_1 _16323_ (.Y(_09569_),
    .B1(_09432_),
    .B2(\cpu.dcache.r_tag[4][5] ),
    .A2(net690),
    .A1(\cpu.dcache.r_tag[3][5] ));
 sg13g2_a22oi_1 _16324_ (.Y(_09570_),
    .B1(net691),
    .B2(\cpu.dcache.r_tag[2][5] ),
    .A2(net627),
    .A1(\cpu.dcache.r_tag[7][5] ));
 sg13g2_a22oi_1 _16325_ (.Y(_09571_),
    .B1(net622),
    .B2(\cpu.dcache.r_tag[5][5] ),
    .A2(_09401_),
    .A1(\cpu.dcache.r_tag[1][5] ));
 sg13g2_inv_1 _16326_ (.Y(_09572_),
    .A(_00228_));
 sg13g2_a22oi_1 _16327_ (.Y(_09573_),
    .B1(net688),
    .B2(_09572_),
    .A2(net689),
    .A1(\cpu.dcache.r_tag[6][5] ));
 sg13g2_and4_1 _16328_ (.A(_09569_),
    .B(_09570_),
    .C(_09571_),
    .D(_09573_),
    .X(_09574_));
 sg13g2_xnor2_1 _16329_ (.Y(_09575_),
    .A(net1034),
    .B(_09574_));
 sg13g2_inv_1 _16330_ (.Y(_09576_),
    .A(_00230_));
 sg13g2_a22oi_1 _16331_ (.Y(_09577_),
    .B1(net688),
    .B2(_09576_),
    .A2(net622),
    .A1(\cpu.dcache.r_tag[5][6] ));
 sg13g2_a22oi_1 _16332_ (.Y(_09578_),
    .B1(net689),
    .B2(\cpu.dcache.r_tag[6][6] ),
    .A2(net692),
    .A1(\cpu.dcache.r_tag[1][6] ));
 sg13g2_a22oi_1 _16333_ (.Y(_09579_),
    .B1(_09432_),
    .B2(\cpu.dcache.r_tag[4][6] ),
    .A2(net690),
    .A1(\cpu.dcache.r_tag[3][6] ));
 sg13g2_a22oi_1 _16334_ (.Y(_09580_),
    .B1(net691),
    .B2(\cpu.dcache.r_tag[2][6] ),
    .A2(net627),
    .A1(\cpu.dcache.r_tag[7][6] ));
 sg13g2_nand4_1 _16335_ (.B(_09578_),
    .C(_09579_),
    .A(_09577_),
    .Y(_09581_),
    .D(_09580_));
 sg13g2_xnor2_1 _16336_ (.Y(_09582_),
    .A(_00229_),
    .B(_09581_));
 sg13g2_nand2_1 _16337_ (.Y(_09583_),
    .A(net1035),
    .B(\cpu.dcache.r_tag[4][8] ));
 sg13g2_or2_1 _16338_ (.X(_09584_),
    .B(_00234_),
    .A(net1035));
 sg13g2_a21oi_1 _16339_ (.A1(_09583_),
    .A2(_09584_),
    .Y(_09585_),
    .B1(net901));
 sg13g2_or2_1 _16340_ (.X(_09586_),
    .B(net1119),
    .A(net1035));
 sg13g2_nor2_1 _16341_ (.A(_00234_),
    .B(_09586_),
    .Y(_09587_));
 sg13g2_o21ai_1 _16342_ (.B1(_09341_),
    .Y(_09588_),
    .A1(_09585_),
    .A2(_09587_));
 sg13g2_a22oi_1 _16343_ (.Y(_09589_),
    .B1(net689),
    .B2(\cpu.dcache.r_tag[6][8] ),
    .A2(_09401_),
    .A1(\cpu.dcache.r_tag[1][8] ));
 sg13g2_a22oi_1 _16344_ (.Y(_09590_),
    .B1(net690),
    .B2(\cpu.dcache.r_tag[3][8] ),
    .A2(_09407_),
    .A1(\cpu.dcache.r_tag[2][8] ));
 sg13g2_a22oi_1 _16345_ (.Y(_09591_),
    .B1(_09423_),
    .B2(\cpu.dcache.r_tag[5][8] ),
    .A2(_09396_),
    .A1(\cpu.dcache.r_tag[7][8] ));
 sg13g2_nand4_1 _16346_ (.B(_09589_),
    .C(_09590_),
    .A(_09588_),
    .Y(_09592_),
    .D(_09591_));
 sg13g2_xor2_1 _16347_ (.B(_09592_),
    .A(_00233_),
    .X(_09593_));
 sg13g2_inv_1 _16348_ (.Y(_09594_),
    .A(\cpu.dcache.r_tag[4][9] ));
 sg13g2_nor2b_1 _16349_ (.A(net1044),
    .B_N(_09392_),
    .Y(_09595_));
 sg13g2_nand2_1 _16350_ (.Y(_09596_),
    .A(net1119),
    .B(\cpu.dcache.r_tag[2][9] ));
 sg13g2_a221oi_1 _16351_ (.B2(net902),
    .C1(net1040),
    .B1(_09596_),
    .A1(_09594_),
    .Y(_09597_),
    .A2(_09595_));
 sg13g2_mux2_1 _16352_ (.A0(\cpu.dcache.r_tag[6][9] ),
    .A1(\cpu.dcache.r_tag[7][9] ),
    .S(net1040),
    .X(_09598_));
 sg13g2_a22oi_1 _16353_ (.Y(_09599_),
    .B1(_09598_),
    .B2(_09394_),
    .A2(_09411_),
    .A1(\cpu.dcache.r_tag[3][9] ));
 sg13g2_nand2b_1 _16354_ (.Y(_09600_),
    .B(_09599_),
    .A_N(_09597_));
 sg13g2_a22oi_1 _16355_ (.Y(_09601_),
    .B1(\cpu.dcache.r_tag[1][9] ),
    .B2(net1119),
    .A2(\cpu.dcache.r_tag[5][9] ),
    .A1(net1035));
 sg13g2_o21ai_1 _16356_ (.B1(_09586_),
    .Y(_09602_),
    .A1(_09523_),
    .A2(_09601_));
 sg13g2_and2_1 _16357_ (.A(_09341_),
    .B(_09602_),
    .X(_09603_));
 sg13g2_nand2_1 _16358_ (.Y(_09604_),
    .A(_00236_),
    .B(_09429_));
 sg13g2_o21ai_1 _16359_ (.B1(_09604_),
    .Y(_09605_),
    .A1(_09600_),
    .A2(_09603_));
 sg13g2_xnor2_1 _16360_ (.Y(_09606_),
    .A(_00235_),
    .B(_09605_));
 sg13g2_a22oi_1 _16361_ (.Y(_09607_),
    .B1(\cpu.dcache.r_tag[1][7] ),
    .B2(_09398_),
    .A2(\cpu.dcache.r_tag[5][7] ),
    .A1(net1035));
 sg13g2_nand3_1 _16362_ (.B(_09398_),
    .C(\cpu.dcache.r_tag[3][7] ),
    .A(_09199_),
    .Y(_09608_));
 sg13g2_o21ai_1 _16363_ (.B1(_09608_),
    .Y(_09609_),
    .A1(net902),
    .A2(_09607_));
 sg13g2_nand2_1 _16364_ (.Y(_09610_),
    .A(_09269_),
    .B(_09609_));
 sg13g2_mux2_1 _16365_ (.A0(\cpu.dcache.r_tag[4][7] ),
    .A1(\cpu.dcache.r_tag[6][7] ),
    .S(net1044),
    .X(_09611_));
 sg13g2_a22oi_1 _16366_ (.Y(_09612_),
    .B1(_09611_),
    .B2(_09523_),
    .A2(_09521_),
    .A1(\cpu.dcache.r_tag[7][7] ));
 sg13g2_nand2b_1 _16367_ (.Y(_09613_),
    .B(net1035),
    .A_N(_09612_));
 sg13g2_inv_1 _16368_ (.Y(_09614_),
    .A(_00232_));
 sg13g2_a22oi_1 _16369_ (.Y(_09615_),
    .B1(_09429_),
    .B2(_09614_),
    .A2(net691),
    .A1(\cpu.dcache.r_tag[2][7] ));
 sg13g2_nand3_1 _16370_ (.B(_09613_),
    .C(_09615_),
    .A(_09610_),
    .Y(_09616_));
 sg13g2_xor2_1 _16371_ (.B(_09616_),
    .A(_00231_),
    .X(_09617_));
 sg13g2_inv_1 _16372_ (.Y(_09618_),
    .A(_00238_));
 sg13g2_a22oi_1 _16373_ (.Y(_09619_),
    .B1(_09432_),
    .B2(\cpu.dcache.r_tag[4][10] ),
    .A2(_09429_),
    .A1(_09618_));
 sg13g2_a22oi_1 _16374_ (.Y(_09620_),
    .B1(net689),
    .B2(\cpu.dcache.r_tag[6][10] ),
    .A2(_09401_),
    .A1(\cpu.dcache.r_tag[1][10] ));
 sg13g2_a22oi_1 _16375_ (.Y(_09621_),
    .B1(_09411_),
    .B2(\cpu.dcache.r_tag[3][10] ),
    .A2(_09396_),
    .A1(\cpu.dcache.r_tag[7][10] ));
 sg13g2_a22oi_1 _16376_ (.Y(_09622_),
    .B1(_09423_),
    .B2(\cpu.dcache.r_tag[5][10] ),
    .A2(_09407_),
    .A1(\cpu.dcache.r_tag[2][10] ));
 sg13g2_nand4_1 _16377_ (.B(_09620_),
    .C(_09621_),
    .A(_09619_),
    .Y(_09623_),
    .D(_09622_));
 sg13g2_xor2_1 _16378_ (.B(_09623_),
    .A(_00237_),
    .X(_09624_));
 sg13g2_nand4_1 _16379_ (.B(_09606_),
    .C(_09617_),
    .A(_09593_),
    .Y(_09625_),
    .D(_09624_));
 sg13g2_nor4_1 _16380_ (.A(_09566_),
    .B(_09575_),
    .C(_09582_),
    .D(_09625_),
    .Y(_09626_));
 sg13g2_mux4_1 _16381_ (.S0(net680),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .S1(net679),
    .X(_09627_));
 sg13g2_mux4_1 _16382_ (.S0(net680),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .S1(net679),
    .X(_09628_));
 sg13g2_mux4_1 _16383_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .S1(net777),
    .X(_09629_));
 sg13g2_mux4_1 _16384_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .S1(net777),
    .X(_09630_));
 sg13g2_mux4_1 _16385_ (.S0(net776),
    .A0(_09627_),
    .A1(_09628_),
    .A2(_09629_),
    .A3(_09630_),
    .S1(net775),
    .X(_09631_));
 sg13g2_nand2_1 _16386_ (.Y(_09632_),
    .A(net686),
    .B(_09631_));
 sg13g2_mux4_1 _16387_ (.S0(_09500_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .S1(_09501_),
    .X(_09633_));
 sg13g2_mux4_1 _16388_ (.S0(_09500_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .S1(_09501_),
    .X(_09634_));
 sg13g2_mux4_1 _16389_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .S1(_09442_),
    .X(_09635_));
 sg13g2_mux4_1 _16390_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .S1(net777),
    .X(_09636_));
 sg13g2_mux4_1 _16391_ (.S0(_09446_),
    .A0(_09633_),
    .A1(_09634_),
    .A2(_09635_),
    .A3(_09636_),
    .S1(_09447_),
    .X(_09637_));
 sg13g2_nand2_1 _16392_ (.Y(_09638_),
    .A(net687),
    .B(_09637_));
 sg13g2_a21oi_1 _16393_ (.A1(_09632_),
    .A2(_09638_),
    .Y(_09639_),
    .B1(_08694_));
 sg13g2_buf_1 _16394_ (.A(_09639_),
    .X(_09640_));
 sg13g2_buf_1 _16395_ (.A(net688),
    .X(_09641_));
 sg13g2_a22oi_1 _16396_ (.Y(_09642_),
    .B1(net691),
    .B2(\cpu.dcache.r_tag[2][23] ),
    .A2(net692),
    .A1(\cpu.dcache.r_tag[1][23] ));
 sg13g2_a22oi_1 _16397_ (.Y(_09643_),
    .B1(_09412_),
    .B2(\cpu.dcache.r_tag[3][23] ),
    .A2(net627),
    .A1(\cpu.dcache.r_tag[7][23] ));
 sg13g2_mux2_1 _16398_ (.A0(\cpu.dcache.r_tag[4][23] ),
    .A1(\cpu.dcache.r_tag[6][23] ),
    .S(_09198_),
    .X(_09644_));
 sg13g2_a22oi_1 _16399_ (.Y(_09645_),
    .B1(_09644_),
    .B2(_09523_),
    .A2(_09421_),
    .A1(\cpu.dcache.r_tag[5][23] ));
 sg13g2_nand2b_1 _16400_ (.Y(_09646_),
    .B(net1035),
    .A_N(_09645_));
 sg13g2_and4_1 _16401_ (.A(_09517_),
    .B(_09642_),
    .C(_09643_),
    .D(_09646_),
    .X(_09647_));
 sg13g2_a21oi_1 _16402_ (.A1(_00249_),
    .A2(net619),
    .Y(_09648_),
    .B1(_09647_));
 sg13g2_xnor2_1 _16403_ (.Y(_09649_),
    .A(net378),
    .B(_09648_));
 sg13g2_nand4_1 _16404_ (.B(_09554_),
    .C(_09626_),
    .A(_09530_),
    .Y(_09650_),
    .D(_09649_));
 sg13g2_mux4_1 _16405_ (.S0(net779),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .S1(net778),
    .X(_09651_));
 sg13g2_mux4_1 _16406_ (.S0(net779),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .S1(_09440_),
    .X(_09652_));
 sg13g2_buf_2 _16407_ (.A(_09439_),
    .X(_09653_));
 sg13g2_mux4_1 _16408_ (.S0(net768),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .S1(net765),
    .X(_09654_));
 sg13g2_mux4_1 _16409_ (.S0(net768),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .S1(net765),
    .X(_09655_));
 sg13g2_mux4_1 _16410_ (.S0(net773),
    .A0(_09651_),
    .A1(_09652_),
    .A2(_09654_),
    .A3(_09655_),
    .S1(net775),
    .X(_09656_));
 sg13g2_nand2_1 _16411_ (.Y(_09657_),
    .A(net686),
    .B(_09656_));
 sg13g2_mux4_1 _16412_ (.S0(net768),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .S1(net765),
    .X(_09658_));
 sg13g2_mux4_1 _16413_ (.S0(_09499_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .S1(net778),
    .X(_09659_));
 sg13g2_mux4_1 _16414_ (.S0(_09472_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .S1(_09653_),
    .X(_09660_));
 sg13g2_mux4_1 _16415_ (.S0(net768),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .S1(net765),
    .X(_09661_));
 sg13g2_mux4_1 _16416_ (.S0(net773),
    .A0(_09658_),
    .A1(_09659_),
    .A2(_09660_),
    .A3(_09661_),
    .S1(net775),
    .X(_09662_));
 sg13g2_nand2_1 _16417_ (.Y(_09663_),
    .A(_09436_),
    .B(_09662_));
 sg13g2_a21oi_1 _16418_ (.A1(_09657_),
    .A2(_09663_),
    .Y(_09664_),
    .B1(_08694_));
 sg13g2_buf_1 _16419_ (.A(_09664_),
    .X(_09665_));
 sg13g2_a22oi_1 _16420_ (.Y(_09666_),
    .B1(net622),
    .B2(\cpu.dcache.r_tag[5][19] ),
    .A2(net689),
    .A1(\cpu.dcache.r_tag[6][19] ));
 sg13g2_a22oi_1 _16421_ (.Y(_09667_),
    .B1(net692),
    .B2(\cpu.dcache.r_tag[1][19] ),
    .A2(net627),
    .A1(\cpu.dcache.r_tag[7][19] ));
 sg13g2_inv_1 _16422_ (.Y(_09668_),
    .A(_00248_));
 sg13g2_a22oi_1 _16423_ (.Y(_09669_),
    .B1(_09432_),
    .B2(\cpu.dcache.r_tag[4][19] ),
    .A2(_09430_),
    .A1(_09668_));
 sg13g2_a22oi_1 _16424_ (.Y(_09670_),
    .B1(net690),
    .B2(\cpu.dcache.r_tag[3][19] ),
    .A2(_09408_),
    .A1(\cpu.dcache.r_tag[2][19] ));
 sg13g2_nand4_1 _16425_ (.B(_09667_),
    .C(_09669_),
    .A(_09666_),
    .Y(_09671_),
    .D(_09670_));
 sg13g2_xnor2_1 _16426_ (.Y(_09672_),
    .A(net417),
    .B(_09671_));
 sg13g2_mux4_1 _16427_ (.S0(net768),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .S1(net765),
    .X(_09673_));
 sg13g2_mux4_1 _16428_ (.S0(net768),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .S1(net765),
    .X(_09674_));
 sg13g2_mux4_1 _16429_ (.S0(net772),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .S1(net771),
    .X(_09675_));
 sg13g2_mux4_1 _16430_ (.S0(net772),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .S1(net771),
    .X(_09676_));
 sg13g2_mux4_1 _16431_ (.S0(net773),
    .A0(_09673_),
    .A1(_09674_),
    .A2(_09675_),
    .A3(_09676_),
    .S1(net775),
    .X(_09677_));
 sg13g2_nand2_1 _16432_ (.Y(_09678_),
    .A(net686),
    .B(_09677_));
 sg13g2_mux4_1 _16433_ (.S0(net768),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .S1(_09653_),
    .X(_09679_));
 sg13g2_mux4_1 _16434_ (.S0(_09499_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .S1(net765),
    .X(_09680_));
 sg13g2_mux4_1 _16435_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .S1(net771),
    .X(_09681_));
 sg13g2_mux4_1 _16436_ (.S0(_09478_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .S1(_09473_),
    .X(_09682_));
 sg13g2_mux4_1 _16437_ (.S0(_09456_),
    .A0(_09679_),
    .A1(_09680_),
    .A2(_09681_),
    .A3(_09682_),
    .S1(_09447_),
    .X(_09683_));
 sg13g2_nand2_1 _16438_ (.Y(_09684_),
    .A(_09436_),
    .B(_09683_));
 sg13g2_a21oi_1 _16439_ (.A1(_09678_),
    .A2(_09684_),
    .Y(_09685_),
    .B1(_08694_));
 sg13g2_buf_1 _16440_ (.A(_09685_),
    .X(_09686_));
 sg13g2_a22oi_1 _16441_ (.Y(_09687_),
    .B1(net622),
    .B2(\cpu.dcache.r_tag[5][16] ),
    .A2(_09397_),
    .A1(\cpu.dcache.r_tag[7][16] ));
 sg13g2_a22oi_1 _16442_ (.Y(_09688_),
    .B1(_09418_),
    .B2(\cpu.dcache.r_tag[6][16] ),
    .A2(_09402_),
    .A1(\cpu.dcache.r_tag[1][16] ));
 sg13g2_inv_1 _16443_ (.Y(_09689_),
    .A(_00245_));
 sg13g2_a22oi_1 _16444_ (.Y(_09690_),
    .B1(_09432_),
    .B2(\cpu.dcache.r_tag[4][16] ),
    .A2(_09429_),
    .A1(_09689_));
 sg13g2_a22oi_1 _16445_ (.Y(_09691_),
    .B1(net690),
    .B2(\cpu.dcache.r_tag[3][16] ),
    .A2(net691),
    .A1(\cpu.dcache.r_tag[2][16] ));
 sg13g2_nand4_1 _16446_ (.B(_09688_),
    .C(_09690_),
    .A(_09687_),
    .Y(_09692_),
    .D(_09691_));
 sg13g2_xnor2_1 _16447_ (.Y(_09693_),
    .A(net416),
    .B(_09692_));
 sg13g2_a22oi_1 _16448_ (.Y(_09694_),
    .B1(_09418_),
    .B2(\cpu.dcache.r_tag[6][15] ),
    .A2(net690),
    .A1(\cpu.dcache.r_tag[3][15] ));
 sg13g2_a22oi_1 _16449_ (.Y(_09695_),
    .B1(_09424_),
    .B2(\cpu.dcache.r_tag[5][15] ),
    .A2(_09402_),
    .A1(\cpu.dcache.r_tag[1][15] ));
 sg13g2_a22oi_1 _16450_ (.Y(_09696_),
    .B1(_09432_),
    .B2(\cpu.dcache.r_tag[4][15] ),
    .A2(net691),
    .A1(\cpu.dcache.r_tag[2][15] ));
 sg13g2_inv_1 _16451_ (.Y(_09697_),
    .A(_00244_));
 sg13g2_a22oi_1 _16452_ (.Y(_09698_),
    .B1(_09430_),
    .B2(_09697_),
    .A2(_09397_),
    .A1(\cpu.dcache.r_tag[7][15] ));
 sg13g2_nand4_1 _16453_ (.B(_09695_),
    .C(_09696_),
    .A(_09694_),
    .Y(_09699_),
    .D(_09698_));
 sg13g2_mux4_1 _16454_ (.S0(net896),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .S1(net774),
    .X(_09700_));
 sg13g2_mux4_1 _16455_ (.S0(net896),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .S1(_09476_),
    .X(_09701_));
 sg13g2_mux4_1 _16456_ (.S0(net896),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .S1(net774),
    .X(_09702_));
 sg13g2_mux4_1 _16457_ (.S0(_09452_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .S1(_09450_),
    .X(_09703_));
 sg13g2_mux4_1 _16458_ (.S0(_08504_),
    .A0(_09700_),
    .A1(_09701_),
    .A2(_09702_),
    .A3(_09703_),
    .S1(net922),
    .X(_09704_));
 sg13g2_nand2_1 _16459_ (.Y(_09705_),
    .A(_08463_),
    .B(_09704_));
 sg13g2_mux4_1 _16460_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .S1(net770),
    .X(_09706_));
 sg13g2_mux4_1 _16461_ (.S0(_09472_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .S1(_09473_),
    .X(_09707_));
 sg13g2_mux4_1 _16462_ (.S0(net896),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .S1(net774),
    .X(_09708_));
 sg13g2_mux4_1 _16463_ (.S0(_09452_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .S1(_09450_),
    .X(_09709_));
 sg13g2_mux4_1 _16464_ (.S0(_08504_),
    .A0(_09706_),
    .A1(_09707_),
    .A2(_09708_),
    .A3(_09709_),
    .S1(net922),
    .X(_09710_));
 sg13g2_o21ai_1 _16465_ (.B1(net1059),
    .Y(_09711_),
    .A1(_08464_),
    .A2(_09710_));
 sg13g2_o21ai_1 _16466_ (.B1(_09711_),
    .Y(_09712_),
    .A1(net1059),
    .A2(_09705_));
 sg13g2_buf_1 _16467_ (.A(_09712_),
    .X(_09713_));
 sg13g2_xnor2_1 _16468_ (.Y(_09714_),
    .A(_09699_),
    .B(net415));
 sg13g2_mux4_1 _16469_ (.S0(net772),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .S1(net771),
    .X(_09715_));
 sg13g2_mux4_1 _16470_ (.S0(net772),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .S1(net765),
    .X(_09716_));
 sg13g2_mux4_1 _16471_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .S1(net770),
    .X(_09717_));
 sg13g2_mux4_1 _16472_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .S1(net770),
    .X(_09718_));
 sg13g2_mux4_1 _16473_ (.S0(net773),
    .A0(_09715_),
    .A1(_09716_),
    .A2(_09717_),
    .A3(_09718_),
    .S1(_08599_),
    .X(_09719_));
 sg13g2_nand2_1 _16474_ (.Y(_09720_),
    .A(_09449_),
    .B(_09719_));
 sg13g2_mux4_1 _16475_ (.S0(net772),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .S1(net771),
    .X(_09721_));
 sg13g2_mux4_1 _16476_ (.S0(net772),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .S1(net771),
    .X(_09722_));
 sg13g2_mux4_1 _16477_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .S1(net770),
    .X(_09723_));
 sg13g2_mux4_1 _16478_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .S1(net770),
    .X(_09724_));
 sg13g2_mux4_1 _16479_ (.S0(net773),
    .A0(_09721_),
    .A1(_09722_),
    .A2(_09723_),
    .A3(_09724_),
    .S1(_08599_),
    .X(_09725_));
 sg13g2_nand2_1 _16480_ (.Y(_09726_),
    .A(net687),
    .B(_09725_));
 sg13g2_a21oi_2 _16481_ (.B1(_08694_),
    .Y(_09727_),
    .A2(_09726_),
    .A1(_09720_));
 sg13g2_buf_1 _16482_ (.A(_09727_),
    .X(_09728_));
 sg13g2_nand2_1 _16483_ (.Y(_09729_),
    .A(\cpu.dcache.r_tag[2][20] ),
    .B(net625));
 sg13g2_a22oi_1 _16484_ (.Y(_09730_),
    .B1(_09433_),
    .B2(\cpu.dcache.r_tag[4][20] ),
    .A2(net688),
    .A1(\cpu.dcache.r_tag[0][20] ));
 sg13g2_a22oi_1 _16485_ (.Y(_09731_),
    .B1(net624),
    .B2(\cpu.dcache.r_tag[3][20] ),
    .A2(net692),
    .A1(\cpu.dcache.r_tag[1][20] ));
 sg13g2_nor2_2 _16486_ (.A(net1040),
    .B(_09341_),
    .Y(_09732_));
 sg13g2_mux2_1 _16487_ (.A0(\cpu.dcache.r_tag[5][20] ),
    .A1(\cpu.dcache.r_tag[7][20] ),
    .S(net902),
    .X(_09733_));
 sg13g2_a22oi_1 _16488_ (.Y(_09734_),
    .B1(_09733_),
    .B2(net901),
    .A2(_09732_),
    .A1(\cpu.dcache.r_tag[6][20] ));
 sg13g2_nand2b_1 _16489_ (.Y(_09735_),
    .B(_09526_),
    .A_N(_09734_));
 sg13g2_nand4_1 _16490_ (.B(_09730_),
    .C(_09731_),
    .A(_09729_),
    .Y(_09736_),
    .D(_09735_));
 sg13g2_xnor2_1 _16491_ (.Y(_09737_),
    .A(net414),
    .B(_09736_));
 sg13g2_and4_1 _16492_ (.A(_09672_),
    .B(_09693_),
    .C(_09714_),
    .D(_09737_),
    .X(_09738_));
 sg13g2_buf_2 _16493_ (.A(net778),
    .X(_09739_));
 sg13g2_mux4_1 _16494_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .S1(_09739_),
    .X(_09740_));
 sg13g2_mux4_1 _16495_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .S1(net677),
    .X(_09741_));
 sg13g2_mux4_1 _16496_ (.S0(net682),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .S1(net681),
    .X(_09742_));
 sg13g2_mux4_1 _16497_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .S1(net677),
    .X(_09743_));
 sg13g2_buf_2 _16498_ (.A(_09446_),
    .X(_09744_));
 sg13g2_mux4_1 _16499_ (.S0(_09744_),
    .A0(_09740_),
    .A1(_09741_),
    .A2(_09742_),
    .A3(_09743_),
    .S1(net678),
    .X(_09745_));
 sg13g2_nand2_1 _16500_ (.Y(_09746_),
    .A(net686),
    .B(_09745_));
 sg13g2_mux4_1 _16501_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .S1(net677),
    .X(_09747_));
 sg13g2_mux4_1 _16502_ (.S0(_09460_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .S1(_09739_),
    .X(_09748_));
 sg13g2_mux4_1 _16503_ (.S0(_09496_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .S1(_09497_),
    .X(_09749_));
 sg13g2_mux4_1 _16504_ (.S0(_09496_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .S1(_09497_),
    .X(_09750_));
 sg13g2_mux4_1 _16505_ (.S0(net776),
    .A0(_09747_),
    .A1(_09748_),
    .A2(_09749_),
    .A3(_09750_),
    .S1(net678),
    .X(_09751_));
 sg13g2_nand2_1 _16506_ (.Y(_09752_),
    .A(net687),
    .B(_09751_));
 sg13g2_a21oi_2 _16507_ (.B1(net1053),
    .Y(_09753_),
    .A2(_09752_),
    .A1(_09746_));
 sg13g2_buf_1 _16508_ (.A(_09753_),
    .X(_09754_));
 sg13g2_a22oi_1 _16509_ (.Y(_09755_),
    .B1(_09419_),
    .B2(\cpu.dcache.r_tag[6][18] ),
    .A2(net626),
    .A1(\cpu.dcache.r_tag[1][18] ));
 sg13g2_a22oi_1 _16510_ (.Y(_09756_),
    .B1(_09413_),
    .B2(\cpu.dcache.r_tag[3][18] ),
    .A2(_09409_),
    .A1(\cpu.dcache.r_tag[2][18] ));
 sg13g2_buf_1 _16511_ (.A(net627),
    .X(_09757_));
 sg13g2_a22oi_1 _16512_ (.Y(_09758_),
    .B1(_09533_),
    .B2(\cpu.dcache.r_tag[5][18] ),
    .A2(_09757_),
    .A1(\cpu.dcache.r_tag[7][18] ));
 sg13g2_inv_1 _16513_ (.Y(_09759_),
    .A(_00247_));
 sg13g2_a22oi_1 _16514_ (.Y(_09760_),
    .B1(_09433_),
    .B2(\cpu.dcache.r_tag[4][18] ),
    .A2(net688),
    .A1(_09759_));
 sg13g2_nand4_1 _16515_ (.B(_09756_),
    .C(_09758_),
    .A(_09755_),
    .Y(_09761_),
    .D(_09760_));
 sg13g2_xnor2_1 _16516_ (.Y(_09762_),
    .A(net377),
    .B(_09761_));
 sg13g2_mux4_1 _16517_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .S1(net677),
    .X(_09763_));
 sg13g2_mux4_1 _16518_ (.S0(_09460_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .S1(net677),
    .X(_09764_));
 sg13g2_mux4_1 _16519_ (.S0(net682),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .S1(net681),
    .X(_09765_));
 sg13g2_mux4_1 _16520_ (.S0(net682),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .S1(net681),
    .X(_09766_));
 sg13g2_mux4_1 _16521_ (.S0(_09744_),
    .A0(_09763_),
    .A1(_09764_),
    .A2(_09765_),
    .A3(_09766_),
    .S1(net678),
    .X(_09767_));
 sg13g2_nand2_1 _16522_ (.Y(_09768_),
    .A(net686),
    .B(_09767_));
 sg13g2_mux4_1 _16523_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .S1(net677),
    .X(_09769_));
 sg13g2_mux4_1 _16524_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .S1(net677),
    .X(_09770_));
 sg13g2_mux4_1 _16525_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .S1(net683),
    .X(_09771_));
 sg13g2_mux4_1 _16526_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .S1(net683),
    .X(_09772_));
 sg13g2_mux4_1 _16527_ (.S0(net776),
    .A0(_09769_),
    .A1(_09770_),
    .A2(_09771_),
    .A3(_09772_),
    .S1(net678),
    .X(_09773_));
 sg13g2_nand2_1 _16528_ (.Y(_09774_),
    .A(net687),
    .B(_09773_));
 sg13g2_a21oi_2 _16529_ (.B1(_08695_),
    .Y(_09775_),
    .A2(_09774_),
    .A1(_09768_));
 sg13g2_buf_1 _16530_ (.A(_09775_),
    .X(_09776_));
 sg13g2_a22oi_1 _16531_ (.Y(_09777_),
    .B1(_09412_),
    .B2(\cpu.dcache.r_tag[3][22] ),
    .A2(_09408_),
    .A1(\cpu.dcache.r_tag[2][22] ));
 sg13g2_a22oi_1 _16532_ (.Y(_09778_),
    .B1(_09432_),
    .B2(\cpu.dcache.r_tag[4][22] ),
    .A2(_09396_),
    .A1(\cpu.dcache.r_tag[7][22] ));
 sg13g2_a22oi_1 _16533_ (.Y(_09779_),
    .B1(_09424_),
    .B2(\cpu.dcache.r_tag[5][22] ),
    .A2(net689),
    .A1(\cpu.dcache.r_tag[6][22] ));
 sg13g2_nand3_1 _16534_ (.B(_09778_),
    .C(_09779_),
    .A(_09777_),
    .Y(_09780_));
 sg13g2_nand2b_1 _16535_ (.Y(_09781_),
    .B(_09515_),
    .A_N(\cpu.dcache.r_tag[0][22] ));
 sg13g2_o21ai_1 _16536_ (.B1(_09781_),
    .Y(_09782_),
    .A1(_09515_),
    .A2(_09780_));
 sg13g2_o21ai_1 _16537_ (.B1(_09403_),
    .Y(_09783_),
    .A1(\cpu.dcache.r_tag[1][22] ),
    .A2(_09780_));
 sg13g2_o21ai_1 _16538_ (.B1(_09783_),
    .Y(_09784_),
    .A1(_09403_),
    .A2(_09782_));
 sg13g2_xnor2_1 _16539_ (.Y(_09785_),
    .A(net376),
    .B(_09784_));
 sg13g2_mux4_1 _16540_ (.S0(net682),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .S1(net681),
    .X(_09786_));
 sg13g2_mux4_1 _16541_ (.S0(net682),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .S1(net681),
    .X(_09787_));
 sg13g2_mux4_1 _16542_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .S1(net683),
    .X(_09788_));
 sg13g2_mux4_1 _16543_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .S1(net683),
    .X(_09789_));
 sg13g2_mux4_1 _16544_ (.S0(net776),
    .A0(_09786_),
    .A1(_09787_),
    .A2(_09788_),
    .A3(_09789_),
    .S1(_09538_),
    .X(_09790_));
 sg13g2_nand2_1 _16545_ (.Y(_09791_),
    .A(net686),
    .B(_09790_));
 sg13g2_mux4_1 _16546_ (.S0(net682),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .S1(net681),
    .X(_09792_));
 sg13g2_mux4_1 _16547_ (.S0(net682),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .S1(net681),
    .X(_09793_));
 sg13g2_mux4_1 _16548_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .S1(net683),
    .X(_09794_));
 sg13g2_mux4_1 _16549_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .S1(net683),
    .X(_09795_));
 sg13g2_mux4_1 _16550_ (.S0(net776),
    .A0(_09792_),
    .A1(_09793_),
    .A2(_09794_),
    .A3(_09795_),
    .S1(_09538_),
    .X(_09796_));
 sg13g2_nand2_1 _16551_ (.Y(_09797_),
    .A(net687),
    .B(_09796_));
 sg13g2_a21oi_1 _16552_ (.A1(_09791_),
    .A2(_09797_),
    .Y(_09798_),
    .B1(_08694_));
 sg13g2_buf_1 _16553_ (.A(_09798_),
    .X(_09799_));
 sg13g2_a22oi_1 _16554_ (.Y(_09800_),
    .B1(_09413_),
    .B2(\cpu.dcache.r_tag[3][21] ),
    .A2(_09409_),
    .A1(\cpu.dcache.r_tag[2][21] ));
 sg13g2_a22oi_1 _16555_ (.Y(_09801_),
    .B1(net623),
    .B2(\cpu.dcache.r_tag[6][21] ),
    .A2(net692),
    .A1(\cpu.dcache.r_tag[1][21] ));
 sg13g2_mux2_1 _16556_ (.A0(\cpu.dcache.r_tag[5][21] ),
    .A1(\cpu.dcache.r_tag[7][21] ),
    .S(net902),
    .X(_09802_));
 sg13g2_a22oi_1 _16557_ (.Y(_09803_),
    .B1(_09802_),
    .B2(_09269_),
    .A2(_09557_),
    .A1(\cpu.dcache.r_tag[4][21] ));
 sg13g2_nand2b_1 _16558_ (.Y(_09804_),
    .B(net894),
    .A_N(_09803_));
 sg13g2_nand4_1 _16559_ (.B(_09800_),
    .C(_09801_),
    .A(_09517_),
    .Y(_09805_),
    .D(_09804_));
 sg13g2_o21ai_1 _16560_ (.B1(_09805_),
    .Y(_09806_),
    .A1(\cpu.dcache.r_tag[0][21] ),
    .A2(_09517_));
 sg13g2_xor2_1 _16561_ (.B(_09806_),
    .A(net375),
    .X(_09807_));
 sg13g2_nand4_1 _16562_ (.B(_09762_),
    .C(_09785_),
    .A(_09738_),
    .Y(_09808_),
    .D(_09807_));
 sg13g2_nor4_1 _16563_ (.A(_09391_),
    .B(_09492_),
    .C(_09650_),
    .D(_09808_),
    .Y(_09809_));
 sg13g2_inv_1 _16564_ (.Y(_09810_),
    .A(_09392_));
 sg13g2_buf_1 _16565_ (.A(_09810_),
    .X(_09811_));
 sg13g2_mux4_1 _16566_ (.S0(_09270_),
    .A0(\cpu.dcache.r_valid[0] ),
    .A1(\cpu.dcache.r_valid[1] ),
    .A2(\cpu.dcache.r_valid[2] ),
    .A3(\cpu.dcache.r_valid[3] ),
    .S1(net784),
    .X(_09812_));
 sg13g2_mux4_1 _16567_ (.S0(net901),
    .A0(\cpu.dcache.r_valid[4] ),
    .A1(\cpu.dcache.r_valid[5] ),
    .A2(\cpu.dcache.r_valid[6] ),
    .A3(\cpu.dcache.r_valid[7] ),
    .S1(net784),
    .X(_09813_));
 sg13g2_and2_1 _16568_ (.A(_09555_),
    .B(_09813_),
    .X(_09814_));
 sg13g2_a21oi_2 _16569_ (.B1(_09814_),
    .Y(_09815_),
    .A2(_09812_),
    .A1(net893));
 sg13g2_mux4_1 _16570_ (.S0(net901),
    .A0(\cpu.dcache.r_dirty[4] ),
    .A1(\cpu.dcache.r_dirty[5] ),
    .A2(\cpu.dcache.r_dirty[6] ),
    .A3(\cpu.dcache.r_dirty[7] ),
    .S1(_09200_),
    .X(_09816_));
 sg13g2_mux4_1 _16571_ (.S0(net901),
    .A0(\cpu.dcache.r_dirty[0] ),
    .A1(\cpu.dcache.r_dirty[1] ),
    .A2(\cpu.dcache.r_dirty[2] ),
    .A3(\cpu.dcache.r_dirty[3] ),
    .S1(_09200_),
    .X(_09817_));
 sg13g2_mux2_1 _16572_ (.A0(_09816_),
    .A1(_09817_),
    .S(net893),
    .X(_09818_));
 sg13g2_nand3_1 _16573_ (.B(_09259_),
    .C(_09818_),
    .A(_09213_),
    .Y(_09819_));
 sg13g2_nor3_1 _16574_ (.A(_09809_),
    .B(_09815_),
    .C(_09819_),
    .Y(_09820_));
 sg13g2_inv_1 _16575_ (.Y(_09821_),
    .A(_09820_));
 sg13g2_or3_1 _16576_ (.A(_09492_),
    .B(_09650_),
    .C(_09808_),
    .X(_09822_));
 sg13g2_buf_1 _16577_ (.A(_09822_),
    .X(_09823_));
 sg13g2_inv_1 _16578_ (.Y(_09824_),
    .A(_09391_));
 sg13g2_o21ai_1 _16579_ (.B1(_09824_),
    .Y(_09825_),
    .A1(_09823_),
    .A2(_09815_));
 sg13g2_nand3_1 _16580_ (.B(_09213_),
    .C(_09259_),
    .A(net1058),
    .Y(_09826_));
 sg13g2_a21oi_1 _16581_ (.A1(_09821_),
    .A2(_09825_),
    .Y(_09827_),
    .B1(_09826_));
 sg13g2_nand2_1 _16582_ (.Y(_09828_),
    .A(_08468_),
    .B(_09281_));
 sg13g2_a22oi_1 _16583_ (.Y(_09829_),
    .B1(_09827_),
    .B2(_09828_),
    .A2(_09012_),
    .A1(net1128));
 sg13g2_buf_1 _16584_ (.A(_09829_),
    .X(_09830_));
 sg13g2_nand2_1 _16585_ (.Y(_09831_),
    .A(_09390_),
    .B(_09830_));
 sg13g2_buf_1 _16586_ (.A(\cpu.qspi.r_state[7] ),
    .X(_09832_));
 sg13g2_buf_1 _16587_ (.A(\cpu.qspi.r_ind ),
    .X(_09833_));
 sg13g2_buf_1 _16588_ (.A(_00250_),
    .X(_09834_));
 sg13g2_buf_1 _16589_ (.A(\cpu.qspi.r_count[0] ),
    .X(_09835_));
 sg13g2_buf_2 _16590_ (.A(\cpu.qspi.r_count[1] ),
    .X(_09836_));
 sg13g2_buf_1 _16591_ (.A(\cpu.qspi.r_count[2] ),
    .X(_09837_));
 sg13g2_nor3_1 _16592_ (.A(_09835_),
    .B(_09836_),
    .C(_09837_),
    .Y(_09838_));
 sg13g2_nor2b_1 _16593_ (.A(\cpu.qspi.r_count[3] ),
    .B_N(_09838_),
    .Y(_09839_));
 sg13g2_buf_1 _16594_ (.A(_09839_),
    .X(_09840_));
 sg13g2_and2_1 _16595_ (.A(_09834_),
    .B(_09840_),
    .X(_09841_));
 sg13g2_buf_1 _16596_ (.A(_09841_),
    .X(_09842_));
 sg13g2_buf_2 _16597_ (.A(\cpu.qspi.r_state[2] ),
    .X(_09843_));
 sg13g2_buf_1 _16598_ (.A(\cpu.qspi.r_state[1] ),
    .X(_09844_));
 sg13g2_a221oi_1 _16599_ (.B2(_09843_),
    .C1(_09844_),
    .B1(_09842_),
    .A1(_09832_),
    .Y(_09845_),
    .A2(_09833_));
 sg13g2_a21oi_1 _16600_ (.A1(_09831_),
    .A2(_09845_),
    .Y(_00026_),
    .B1(net630));
 sg13g2_buf_1 _16601_ (.A(\cpu.qspi.r_state[16] ),
    .X(_09846_));
 sg13g2_nand2_1 _16602_ (.Y(_09847_),
    .A(_09834_),
    .B(_09840_));
 sg13g2_buf_2 _16603_ (.A(_09847_),
    .X(_09848_));
 sg13g2_and2_1 _16604_ (.A(_08474_),
    .B(_09820_),
    .X(_09849_));
 sg13g2_buf_1 _16605_ (.A(_09849_),
    .X(_09850_));
 sg13g2_buf_2 _16606_ (.A(\cpu.qspi.r_state[8] ),
    .X(_09851_));
 sg13g2_a22oi_1 _16607_ (.Y(_09852_),
    .B1(net142),
    .B2(_09851_),
    .A2(_09848_),
    .A1(net1118));
 sg13g2_nor2_1 _16608_ (.A(net631),
    .B(_09852_),
    .Y(_00025_));
 sg13g2_buf_2 _16609_ (.A(\cpu.qspi.r_state[4] ),
    .X(_09853_));
 sg13g2_buf_1 _16610_ (.A(\cpu.qspi.r_state[9] ),
    .X(_09854_));
 sg13g2_a21oi_1 _16611_ (.A1(_09853_),
    .A2(_09842_),
    .Y(_09855_),
    .B1(_09854_));
 sg13g2_nor2_1 _16612_ (.A(net631),
    .B(_09855_),
    .Y(_00022_));
 sg13g2_buf_1 _16613_ (.A(_08474_),
    .X(_09856_));
 sg13g2_nor2_1 _16614_ (.A(_08474_),
    .B(_08757_),
    .Y(_09857_));
 sg13g2_a21oi_1 _16615_ (.A1(net892),
    .A2(net378),
    .Y(_09858_),
    .B1(_09857_));
 sg13g2_inv_1 _16616_ (.Y(_09859_),
    .A(\cpu.qspi.r_rom_mode[0] ));
 sg13g2_mux2_1 _16617_ (.A0(_09850_),
    .A1(_09858_),
    .S(_09859_),
    .X(_09860_));
 sg13g2_buf_1 _16618_ (.A(\cpu.qspi.r_rom_mode[1] ),
    .X(_09861_));
 sg13g2_nor2b_1 _16619_ (.A(_09860_),
    .B_N(_09861_),
    .Y(_09862_));
 sg13g2_buf_1 _16620_ (.A(_09862_),
    .X(_09863_));
 sg13g2_nor3_1 _16621_ (.A(\cpu.qspi.r_rom_mode[0] ),
    .B(_09861_),
    .C(_09858_),
    .Y(_09864_));
 sg13g2_buf_1 _16622_ (.A(_09864_),
    .X(_09865_));
 sg13g2_nor2_1 _16623_ (.A(net245),
    .B(net88),
    .Y(_09866_));
 sg13g2_and2_1 _16624_ (.A(\cpu.qspi.r_quad[2] ),
    .B(net245),
    .X(_09867_));
 sg13g2_a221oi_1 _16625_ (.B2(\cpu.qspi.r_quad[0] ),
    .C1(_09867_),
    .B1(_09866_),
    .A1(\cpu.qspi.r_quad[1] ),
    .Y(_09868_),
    .A2(net88));
 sg13g2_buf_2 _16626_ (.A(_09868_),
    .X(_09869_));
 sg13g2_inv_1 _16627_ (.Y(_09870_),
    .A(_09390_));
 sg13g2_nor2_1 _16628_ (.A(_09870_),
    .B(_09830_),
    .Y(_09871_));
 sg13g2_a22oi_1 _16629_ (.Y(_09872_),
    .B1(_09869_),
    .B2(_09871_),
    .A2(_09848_),
    .A1(_09853_));
 sg13g2_nor2_1 _16630_ (.A(net631),
    .B(_09872_),
    .Y(_00028_));
 sg13g2_nand2_1 _16631_ (.Y(_09873_),
    .A(_09843_),
    .B(_09848_));
 sg13g2_buf_1 _16632_ (.A(\cpu.qspi.r_state[14] ),
    .X(_09874_));
 sg13g2_nand2_1 _16633_ (.Y(_09875_),
    .A(net1117),
    .B(_09842_));
 sg13g2_a21oi_1 _16634_ (.A1(_09873_),
    .A2(_09875_),
    .Y(_00027_),
    .B1(net630));
 sg13g2_inv_1 _16635_ (.Y(_09876_),
    .A(_09832_));
 sg13g2_buf_1 _16636_ (.A(_09381_),
    .X(_09877_));
 sg13g2_buf_1 _16637_ (.A(net891),
    .X(_09878_));
 sg13g2_buf_1 _16638_ (.A(net764),
    .X(_09879_));
 sg13g2_o21ai_1 _16639_ (.B1(net675),
    .Y(_00021_),
    .A1(_09876_),
    .A2(_09833_));
 sg13g2_buf_1 _16640_ (.A(\cpu.dec.r_op[10] ),
    .X(_09880_));
 sg13g2_nor4_1 _16641_ (.A(_09015_),
    .B(net288),
    .C(_08441_),
    .D(net295),
    .Y(_09881_));
 sg13g2_a21o_1 _16642_ (.A2(_09017_),
    .A1(net1116),
    .B1(_09881_),
    .X(_00011_));
 sg13g2_buf_1 _16643_ (.A(net289),
    .X(_09882_));
 sg13g2_nor2_1 _16644_ (.A(net244),
    .B(_09096_),
    .Y(_09883_));
 sg13g2_nor2b_1 _16645_ (.A(net288),
    .B_N(net295),
    .Y(_09884_));
 sg13g2_a22oi_1 _16646_ (.Y(_09885_),
    .B1(_09884_),
    .B2(_09052_),
    .A2(_09883_),
    .A1(_09105_));
 sg13g2_buf_1 _16647_ (.A(\cpu.dec.r_op[9] ),
    .X(_09886_));
 sg13g2_buf_1 _16648_ (.A(net1115),
    .X(_09887_));
 sg13g2_nor2_1 _16649_ (.A(net1033),
    .B(net119),
    .Y(_09888_));
 sg13g2_a21oi_1 _16650_ (.A1(net107),
    .A2(_09885_),
    .Y(_00020_),
    .B1(_09888_));
 sg13g2_buf_2 _16651_ (.A(\cpu.dec.r_op[8] ),
    .X(_09889_));
 sg13g2_buf_1 _16652_ (.A(_09889_),
    .X(_09890_));
 sg13g2_inv_1 _16653_ (.Y(_09891_),
    .A(net1032));
 sg13g2_buf_1 _16654_ (.A(_09014_),
    .X(_09892_));
 sg13g2_buf_1 _16655_ (.A(_09049_),
    .X(_09893_));
 sg13g2_nor2_1 _16656_ (.A(net195),
    .B(_08377_),
    .Y(_09894_));
 sg13g2_buf_2 _16657_ (.A(_09894_),
    .X(_09895_));
 sg13g2_nor2_1 _16658_ (.A(_09040_),
    .B(_08438_),
    .Y(_09896_));
 sg13g2_buf_2 _16659_ (.A(_09896_),
    .X(_09897_));
 sg13g2_nand3_1 _16660_ (.B(_09895_),
    .C(_09897_),
    .A(_09103_),
    .Y(_09898_));
 sg13g2_o21ai_1 _16661_ (.B1(_09898_),
    .Y(_00019_),
    .A1(_09891_),
    .A2(_09892_));
 sg13g2_buf_1 _16662_ (.A(_00275_),
    .X(_09899_));
 sg13g2_buf_1 _16663_ (.A(\cpu.qspi.r_state[12] ),
    .X(_09900_));
 sg13g2_buf_1 _16664_ (.A(_09900_),
    .X(_09901_));
 sg13g2_nand2_1 _16665_ (.Y(_09902_),
    .A(net1031),
    .B(_09848_));
 sg13g2_a21oi_1 _16666_ (.A1(_09899_),
    .A2(_09902_),
    .Y(_00023_),
    .B1(net630));
 sg13g2_nor2b_1 _16667_ (.A(_09053_),
    .B_N(_09883_),
    .Y(_09903_));
 sg13g2_buf_1 _16668_ (.A(_09171_),
    .X(_09904_));
 sg13g2_nor2_1 _16669_ (.A(_09144_),
    .B(net246),
    .Y(_09905_));
 sg13g2_nand3_1 _16670_ (.B(net220),
    .C(_09905_),
    .A(_09178_),
    .Y(_09906_));
 sg13g2_nor2b_1 _16671_ (.A(_09903_),
    .B_N(_09906_),
    .Y(_09907_));
 sg13g2_buf_1 _16672_ (.A(\cpu.dec.r_op[1] ),
    .X(_09908_));
 sg13g2_nor2_1 _16673_ (.A(_09908_),
    .B(_09000_),
    .Y(_09909_));
 sg13g2_a21oi_1 _16674_ (.A1(_09104_),
    .A2(_09907_),
    .Y(_00012_),
    .B1(_09909_));
 sg13g2_buf_1 _16675_ (.A(\cpu.qspi.r_state[5] ),
    .X(_09910_));
 sg13g2_inv_1 _16676_ (.Y(_09911_),
    .A(net1114));
 sg13g2_nand2_1 _16677_ (.Y(_09912_),
    .A(net1117),
    .B(_09848_));
 sg13g2_a21oi_1 _16678_ (.A1(_09911_),
    .A2(_09912_),
    .Y(_00024_),
    .B1(_09352_));
 sg13g2_buf_1 _16679_ (.A(_09144_),
    .X(_09913_));
 sg13g2_buf_1 _16680_ (.A(net246),
    .X(_09914_));
 sg13g2_nand4_1 _16681_ (.B(_09913_),
    .C(net220),
    .A(_09108_),
    .Y(_09915_),
    .D(net219));
 sg13g2_nand3_1 _16682_ (.B(_09052_),
    .C(_09882_),
    .A(_09038_),
    .Y(_09916_));
 sg13g2_a21oi_1 _16683_ (.A1(_09096_),
    .A2(_09915_),
    .Y(_09917_),
    .B1(_09916_));
 sg13g2_buf_2 _16684_ (.A(_09014_),
    .X(_09918_));
 sg13g2_mux2_1 _16685_ (.A0(\cpu.dec.r_op[7] ),
    .A1(_09917_),
    .S(net105),
    .X(_00018_));
 sg13g2_buf_1 _16686_ (.A(\cpu.uart.r_div[11] ),
    .X(_09919_));
 sg13g2_nor3_1 _16687_ (.A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ),
    .C(\cpu.uart.r_div[2] ),
    .Y(_09920_));
 sg13g2_nor2b_1 _16688_ (.A(\cpu.uart.r_div[3] ),
    .B_N(_09920_),
    .Y(_09921_));
 sg13g2_nor2b_1 _16689_ (.A(\cpu.uart.r_div[4] ),
    .B_N(_09921_),
    .Y(_09922_));
 sg13g2_nor2b_1 _16690_ (.A(\cpu.uart.r_div[5] ),
    .B_N(_09922_),
    .Y(_09923_));
 sg13g2_nor2b_1 _16691_ (.A(\cpu.uart.r_div[6] ),
    .B_N(_09923_),
    .Y(_09924_));
 sg13g2_nand2b_1 _16692_ (.Y(_09925_),
    .B(_09924_),
    .A_N(\cpu.uart.r_div[7] ));
 sg13g2_nor2_1 _16693_ (.A(\cpu.uart.r_div[8] ),
    .B(_09925_),
    .Y(_09926_));
 sg13g2_nand2b_1 _16694_ (.Y(_09927_),
    .B(_09926_),
    .A_N(\cpu.uart.r_div[9] ));
 sg13g2_buf_1 _16695_ (.A(_09927_),
    .X(_09928_));
 sg13g2_nor3_1 _16696_ (.A(\cpu.uart.r_div[10] ),
    .B(_09919_),
    .C(_09928_),
    .Y(_09929_));
 sg13g2_buf_2 _16697_ (.A(_09929_),
    .X(_09930_));
 sg13g2_nor2_1 _16698_ (.A(net781),
    .B(_09930_),
    .Y(_09931_));
 sg13g2_buf_1 _16699_ (.A(_09931_),
    .X(_09932_));
 sg13g2_buf_1 _16700_ (.A(net242),
    .X(_09933_));
 sg13g2_mux2_1 _16701_ (.A0(\cpu.uart.r_div_value[0] ),
    .A1(_00277_),
    .S(net218),
    .X(_00079_));
 sg13g2_xnor2_1 _16702_ (.Y(_09934_),
    .A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ));
 sg13g2_mux2_1 _16703_ (.A0(\cpu.uart.r_div_value[1] ),
    .A1(_09934_),
    .S(net218),
    .X(_00082_));
 sg13g2_o21ai_1 _16704_ (.B1(\cpu.uart.r_div[2] ),
    .Y(_09935_),
    .A1(\cpu.uart.r_div[0] ),
    .A2(\cpu.uart.r_div[1] ));
 sg13g2_nor2b_1 _16705_ (.A(_09920_),
    .B_N(_09935_),
    .Y(_09936_));
 sg13g2_nor2_1 _16706_ (.A(\cpu.uart.r_div_value[2] ),
    .B(_09932_),
    .Y(_09937_));
 sg13g2_a21oi_1 _16707_ (.A1(net218),
    .A2(_09936_),
    .Y(_00083_),
    .B1(_09937_));
 sg13g2_xnor2_1 _16708_ (.Y(_09938_),
    .A(\cpu.uart.r_div[3] ),
    .B(_09920_));
 sg13g2_nor2_1 _16709_ (.A(\cpu.uart.r_div_value[3] ),
    .B(net242),
    .Y(_09939_));
 sg13g2_a21oi_1 _16710_ (.A1(net218),
    .A2(_09938_),
    .Y(_00084_),
    .B1(_09939_));
 sg13g2_xnor2_1 _16711_ (.Y(_09940_),
    .A(\cpu.uart.r_div[4] ),
    .B(_09921_));
 sg13g2_nor2_1 _16712_ (.A(\cpu.uart.r_div_value[4] ),
    .B(net242),
    .Y(_09941_));
 sg13g2_a21oi_1 _16713_ (.A1(net218),
    .A2(_09940_),
    .Y(_00085_),
    .B1(_09941_));
 sg13g2_xnor2_1 _16714_ (.Y(_09942_),
    .A(\cpu.uart.r_div[5] ),
    .B(_09922_));
 sg13g2_nor2_1 _16715_ (.A(\cpu.uart.r_div_value[5] ),
    .B(net242),
    .Y(_09943_));
 sg13g2_a21oi_1 _16716_ (.A1(net218),
    .A2(_09942_),
    .Y(_00086_),
    .B1(_09943_));
 sg13g2_xnor2_1 _16717_ (.Y(_09944_),
    .A(\cpu.uart.r_div[6] ),
    .B(_09923_));
 sg13g2_nor2_1 _16718_ (.A(\cpu.uart.r_div_value[6] ),
    .B(net242),
    .Y(_09945_));
 sg13g2_a21oi_1 _16719_ (.A1(net218),
    .A2(_09944_),
    .Y(_00087_),
    .B1(_09945_));
 sg13g2_xnor2_1 _16720_ (.Y(_09946_),
    .A(\cpu.uart.r_div[7] ),
    .B(_09924_));
 sg13g2_nor2_1 _16721_ (.A(\cpu.uart.r_div_value[7] ),
    .B(net242),
    .Y(_09947_));
 sg13g2_a21oi_1 _16722_ (.A1(_09933_),
    .A2(_09946_),
    .Y(_00088_),
    .B1(_09947_));
 sg13g2_xor2_1 _16723_ (.B(_09925_),
    .A(\cpu.uart.r_div[8] ),
    .X(_09948_));
 sg13g2_nor2_1 _16724_ (.A(\cpu.uart.r_div_value[8] ),
    .B(net242),
    .Y(_09949_));
 sg13g2_a21oi_1 _16725_ (.A1(net218),
    .A2(_09948_),
    .Y(_00089_),
    .B1(_09949_));
 sg13g2_xnor2_1 _16726_ (.Y(_09950_),
    .A(\cpu.uart.r_div[9] ),
    .B(_09926_));
 sg13g2_nor2_1 _16727_ (.A(\cpu.uart.r_div_value[9] ),
    .B(net242),
    .Y(_09951_));
 sg13g2_a21oi_1 _16728_ (.A1(_09933_),
    .A2(_09950_),
    .Y(_00090_),
    .B1(_09951_));
 sg13g2_buf_1 _16729_ (.A(\cpu.uart.r_div_value[10] ),
    .X(_09952_));
 sg13g2_inv_1 _16730_ (.Y(_09953_),
    .A(_09952_));
 sg13g2_buf_1 _16731_ (.A(_09351_),
    .X(_09954_));
 sg13g2_nand2_1 _16732_ (.Y(_09955_),
    .A(net891),
    .B(_09928_));
 sg13g2_o21ai_1 _16733_ (.B1(_09955_),
    .Y(_09956_),
    .A1(_09919_),
    .A2(_09952_));
 sg13g2_inv_1 _16734_ (.Y(_09957_),
    .A(\cpu.uart.r_div[10] ));
 sg13g2_nor3_1 _16735_ (.A(_09957_),
    .B(_09351_),
    .C(_09928_),
    .Y(_09958_));
 sg13g2_a221oi_1 _16736_ (.B2(_09957_),
    .C1(_09958_),
    .B1(_09956_),
    .A1(_09953_),
    .Y(_00080_),
    .A2(net618));
 sg13g2_nor2_1 _16737_ (.A(\cpu.uart.r_div[10] ),
    .B(_09928_),
    .Y(_09959_));
 sg13g2_nand2_1 _16738_ (.Y(_09960_),
    .A(_09919_),
    .B(net764));
 sg13g2_o21ai_1 _16739_ (.B1(\cpu.uart.r_div_value[11] ),
    .Y(_09961_),
    .A1(_09351_),
    .A2(_09930_));
 sg13g2_o21ai_1 _16740_ (.B1(_09961_),
    .Y(_00081_),
    .A1(_09959_),
    .A2(_09960_));
 sg13g2_buf_1 _16741_ (.A(\cpu.intr.r_timer_count[19] ),
    .X(_09962_));
 sg13g2_buf_1 _16742_ (.A(\cpu.intr.r_timer_count[18] ),
    .X(_09963_));
 sg13g2_buf_1 _16743_ (.A(\cpu.intr.r_timer_count[17] ),
    .X(_09964_));
 sg13g2_buf_1 _16744_ (.A(\cpu.intr.r_timer_count[16] ),
    .X(_09965_));
 sg13g2_buf_1 _16745_ (.A(\cpu.intr.r_timer_count[10] ),
    .X(_09966_));
 sg13g2_buf_1 _16746_ (.A(\cpu.intr.r_timer_count[7] ),
    .X(_09967_));
 sg13g2_buf_1 _16747_ (.A(\cpu.intr.r_timer_count[1] ),
    .X(_09968_));
 sg13g2_nor3_1 _16748_ (.A(_09968_),
    .B(\cpu.intr.r_timer_count[0] ),
    .C(\cpu.intr.r_timer_count[2] ),
    .Y(_09969_));
 sg13g2_nor2b_1 _16749_ (.A(\cpu.intr.r_timer_count[3] ),
    .B_N(_09969_),
    .Y(_09970_));
 sg13g2_nor2b_1 _16750_ (.A(\cpu.intr.r_timer_count[4] ),
    .B_N(_09970_),
    .Y(_09971_));
 sg13g2_nor2b_1 _16751_ (.A(\cpu.intr.r_timer_count[5] ),
    .B_N(_09971_),
    .Y(_09972_));
 sg13g2_nand2b_1 _16752_ (.Y(_09973_),
    .B(_09972_),
    .A_N(\cpu.intr.r_timer_count[6] ));
 sg13g2_nor3_1 _16753_ (.A(_09967_),
    .B(\cpu.intr.r_timer_count[8] ),
    .C(_09973_),
    .Y(_09974_));
 sg13g2_nand2b_1 _16754_ (.Y(_09975_),
    .B(_09974_),
    .A_N(\cpu.intr.r_timer_count[9] ));
 sg13g2_nor3_1 _16755_ (.A(\cpu.intr.r_timer_count[11] ),
    .B(_09966_),
    .C(_09975_),
    .Y(_09976_));
 sg13g2_nor2b_1 _16756_ (.A(\cpu.intr.r_timer_count[12] ),
    .B_N(_09976_),
    .Y(_09977_));
 sg13g2_nor2b_1 _16757_ (.A(\cpu.intr.r_timer_count[13] ),
    .B_N(_09977_),
    .Y(_09978_));
 sg13g2_nor2b_1 _16758_ (.A(\cpu.intr.r_timer_count[14] ),
    .B_N(_09978_),
    .Y(_09979_));
 sg13g2_nand2b_1 _16759_ (.Y(_09980_),
    .B(_09979_),
    .A_N(\cpu.intr.r_timer_count[15] ));
 sg13g2_nor3_1 _16760_ (.A(_09964_),
    .B(_09965_),
    .C(_09980_),
    .Y(_09981_));
 sg13g2_nor2b_1 _16761_ (.A(_09963_),
    .B_N(_09981_),
    .Y(_09982_));
 sg13g2_nand2b_1 _16762_ (.Y(_09983_),
    .B(_09982_),
    .A_N(_09962_));
 sg13g2_buf_1 _16763_ (.A(_09983_),
    .X(_09984_));
 sg13g2_buf_1 _16764_ (.A(\cpu.intr.r_timer_count[21] ),
    .X(_09985_));
 sg13g2_buf_2 _16765_ (.A(\cpu.intr.r_timer_count[20] ),
    .X(_09986_));
 sg13g2_buf_1 _16766_ (.A(\cpu.intr.r_timer_count[23] ),
    .X(_09987_));
 sg13g2_buf_1 _16767_ (.A(\cpu.intr.r_timer_count[22] ),
    .X(_09988_));
 sg13g2_nor4_2 _16768_ (.A(_09985_),
    .B(_09986_),
    .C(_09987_),
    .Y(_09989_),
    .D(_09988_));
 sg13g2_nand2b_1 _16769_ (.Y(_09990_),
    .B(_09989_),
    .A_N(_09984_));
 sg13g2_buf_2 _16770_ (.A(_09990_),
    .X(_09991_));
 sg13g2_buf_1 _16771_ (.A(net782),
    .X(_09992_));
 sg13g2_buf_1 _16772_ (.A(net674),
    .X(_09993_));
 sg13g2_buf_1 _16773_ (.A(net540),
    .X(_09994_));
 sg13g2_buf_1 _16774_ (.A(net472),
    .X(_09995_));
 sg13g2_buf_1 _16775_ (.A(net413),
    .X(_09996_));
 sg13g2_buf_1 _16776_ (.A(net374),
    .X(_09997_));
 sg13g2_buf_1 _16777_ (.A(\cpu.addr[5] ),
    .X(_09998_));
 sg13g2_buf_1 _16778_ (.A(_09998_),
    .X(_09999_));
 sg13g2_nor3_2 _16779_ (.A(net1030),
    .B(net1043),
    .C(net1042),
    .Y(_10000_));
 sg13g2_nand2_2 _16780_ (.Y(_10001_),
    .A(_09206_),
    .B(_10000_));
 sg13g2_nor2_1 _16781_ (.A(_09261_),
    .B(_10001_),
    .Y(_10002_));
 sg13g2_buf_1 _16782_ (.A(_10002_),
    .X(_10003_));
 sg13g2_nand3_1 _16783_ (.B(_09997_),
    .C(net171),
    .A(net617),
    .Y(_10004_));
 sg13g2_buf_1 _16784_ (.A(_10004_),
    .X(_10005_));
 sg13g2_nand2_1 _16785_ (.Y(_10006_),
    .A(_09991_),
    .B(_10005_));
 sg13g2_buf_2 _16786_ (.A(_10006_),
    .X(_10007_));
 sg13g2_buf_8 _16787_ (.A(_10007_),
    .X(_10008_));
 sg13g2_mux2_1 _16788_ (.A0(_00283_),
    .A1(\cpu.intr.r_timer_reload[0] ),
    .S(net70),
    .X(_00055_));
 sg13g2_buf_8 _16789_ (.A(_10007_),
    .X(_10009_));
 sg13g2_xor2_1 _16790_ (.B(\cpu.intr.r_timer_count[0] ),
    .A(_09968_),
    .X(_10010_));
 sg13g2_nand2_1 _16791_ (.Y(_10011_),
    .A(\cpu.intr.r_timer_reload[1] ),
    .B(net70));
 sg13g2_o21ai_1 _16792_ (.B1(_10011_),
    .Y(_00066_),
    .A1(net69),
    .A2(_10010_));
 sg13g2_o21ai_1 _16793_ (.B1(\cpu.intr.r_timer_count[2] ),
    .Y(_10012_),
    .A1(_09968_),
    .A2(\cpu.intr.r_timer_count[0] ));
 sg13g2_nor2b_1 _16794_ (.A(_09969_),
    .B_N(_10012_),
    .Y(_10013_));
 sg13g2_nand2_1 _16795_ (.Y(_10014_),
    .A(\cpu.intr.r_timer_reload[2] ),
    .B(net70));
 sg13g2_o21ai_1 _16796_ (.B1(_10014_),
    .Y(_00071_),
    .A1(net69),
    .A2(_10013_));
 sg13g2_xnor2_1 _16797_ (.Y(_10015_),
    .A(\cpu.intr.r_timer_count[3] ),
    .B(_09969_));
 sg13g2_nand2_1 _16798_ (.Y(_10016_),
    .A(\cpu.intr.r_timer_reload[3] ),
    .B(_10008_));
 sg13g2_o21ai_1 _16799_ (.B1(_10016_),
    .Y(_00072_),
    .A1(net69),
    .A2(_10015_));
 sg13g2_xnor2_1 _16800_ (.Y(_10017_),
    .A(\cpu.intr.r_timer_count[4] ),
    .B(_09970_));
 sg13g2_nand2_1 _16801_ (.Y(_10018_),
    .A(\cpu.intr.r_timer_reload[4] ),
    .B(_10008_));
 sg13g2_o21ai_1 _16802_ (.B1(_10018_),
    .Y(_00073_),
    .A1(net69),
    .A2(_10017_));
 sg13g2_xnor2_1 _16803_ (.Y(_10019_),
    .A(\cpu.intr.r_timer_count[5] ),
    .B(_09971_));
 sg13g2_buf_8 _16804_ (.A(_10007_),
    .X(_10020_));
 sg13g2_nand2_1 _16805_ (.Y(_10021_),
    .A(\cpu.intr.r_timer_reload[5] ),
    .B(net68));
 sg13g2_o21ai_1 _16806_ (.B1(_10021_),
    .Y(_00074_),
    .A1(_10009_),
    .A2(_10019_));
 sg13g2_xnor2_1 _16807_ (.Y(_10022_),
    .A(\cpu.intr.r_timer_count[6] ),
    .B(_09972_));
 sg13g2_nand2_1 _16808_ (.Y(_10023_),
    .A(\cpu.intr.r_timer_reload[6] ),
    .B(net68));
 sg13g2_o21ai_1 _16809_ (.B1(_10023_),
    .Y(_00075_),
    .A1(net69),
    .A2(_10022_));
 sg13g2_xor2_1 _16810_ (.B(_09973_),
    .A(_09967_),
    .X(_10024_));
 sg13g2_nand2_1 _16811_ (.Y(_10025_),
    .A(\cpu.intr.r_timer_reload[7] ),
    .B(_10020_));
 sg13g2_o21ai_1 _16812_ (.B1(_10025_),
    .Y(_00076_),
    .A1(net69),
    .A2(_10024_));
 sg13g2_nor2_1 _16813_ (.A(_09967_),
    .B(_09973_),
    .Y(_10026_));
 sg13g2_xnor2_1 _16814_ (.Y(_10027_),
    .A(\cpu.intr.r_timer_count[8] ),
    .B(_10026_));
 sg13g2_nand2_1 _16815_ (.Y(_10028_),
    .A(\cpu.intr.r_timer_reload[8] ),
    .B(_10020_));
 sg13g2_o21ai_1 _16816_ (.B1(_10028_),
    .Y(_00077_),
    .A1(_10009_),
    .A2(_10027_));
 sg13g2_xnor2_1 _16817_ (.Y(_10029_),
    .A(\cpu.intr.r_timer_count[9] ),
    .B(_09974_));
 sg13g2_nand2_1 _16818_ (.Y(_10030_),
    .A(\cpu.intr.r_timer_reload[9] ),
    .B(net68));
 sg13g2_o21ai_1 _16819_ (.B1(_10030_),
    .Y(_00078_),
    .A1(net69),
    .A2(_10029_));
 sg13g2_xor2_1 _16820_ (.B(_09975_),
    .A(_09966_),
    .X(_10031_));
 sg13g2_nand2_1 _16821_ (.Y(_10032_),
    .A(\cpu.intr.r_timer_reload[10] ),
    .B(net68));
 sg13g2_o21ai_1 _16822_ (.B1(_10032_),
    .Y(_00056_),
    .A1(net69),
    .A2(_10031_));
 sg13g2_o21ai_1 _16823_ (.B1(\cpu.intr.r_timer_count[11] ),
    .Y(_10033_),
    .A1(_09966_),
    .A2(_09975_));
 sg13g2_nor2b_1 _16824_ (.A(_09976_),
    .B_N(_10033_),
    .Y(_10034_));
 sg13g2_nand2_1 _16825_ (.Y(_10035_),
    .A(\cpu.intr.r_timer_reload[11] ),
    .B(net68));
 sg13g2_o21ai_1 _16826_ (.B1(_10035_),
    .Y(_00057_),
    .A1(net70),
    .A2(_10034_));
 sg13g2_xnor2_1 _16827_ (.Y(_10036_),
    .A(\cpu.intr.r_timer_count[12] ),
    .B(_09976_));
 sg13g2_nand2_1 _16828_ (.Y(_10037_),
    .A(\cpu.intr.r_timer_reload[12] ),
    .B(net68));
 sg13g2_o21ai_1 _16829_ (.B1(_10037_),
    .Y(_00058_),
    .A1(net70),
    .A2(_10036_));
 sg13g2_xnor2_1 _16830_ (.Y(_10038_),
    .A(\cpu.intr.r_timer_count[13] ),
    .B(_09977_));
 sg13g2_nand2_1 _16831_ (.Y(_10039_),
    .A(\cpu.intr.r_timer_reload[13] ),
    .B(net68));
 sg13g2_o21ai_1 _16832_ (.B1(_10039_),
    .Y(_00059_),
    .A1(net70),
    .A2(_10038_));
 sg13g2_xnor2_1 _16833_ (.Y(_10040_),
    .A(\cpu.intr.r_timer_count[14] ),
    .B(_09978_));
 sg13g2_nand2_1 _16834_ (.Y(_10041_),
    .A(\cpu.intr.r_timer_reload[14] ),
    .B(net68));
 sg13g2_o21ai_1 _16835_ (.B1(_10041_),
    .Y(_00060_),
    .A1(net70),
    .A2(_10040_));
 sg13g2_xnor2_1 _16836_ (.Y(_10042_),
    .A(\cpu.intr.r_timer_count[15] ),
    .B(_09979_));
 sg13g2_nand2_1 _16837_ (.Y(_10043_),
    .A(\cpu.intr.r_timer_reload[15] ),
    .B(_10007_));
 sg13g2_o21ai_1 _16838_ (.B1(_10043_),
    .Y(_00061_),
    .A1(net70),
    .A2(_10042_));
 sg13g2_nor4_1 _16839_ (.A(_09964_),
    .B(_09962_),
    .C(_09963_),
    .D(\cpu.intr.r_timer_reload[16] ),
    .Y(_10044_));
 sg13g2_a21oi_1 _16840_ (.A1(_09989_),
    .A2(_10044_),
    .Y(_10045_),
    .B1(_09965_));
 sg13g2_mux2_1 _16841_ (.A0(_10045_),
    .A1(_09965_),
    .S(_09980_),
    .X(_10046_));
 sg13g2_buf_1 _16842_ (.A(\cpu.dcache.wdata[0] ),
    .X(_10047_));
 sg13g2_buf_1 _16843_ (.A(_10047_),
    .X(_10048_));
 sg13g2_buf_1 _16844_ (.A(net1029),
    .X(_10049_));
 sg13g2_inv_2 _16845_ (.Y(_10050_),
    .A(_09271_));
 sg13g2_buf_1 _16846_ (.A(_10050_),
    .X(_10051_));
 sg13g2_buf_1 _16847_ (.A(net889),
    .X(_10052_));
 sg13g2_buf_1 _16848_ (.A(net763),
    .X(_10053_));
 sg13g2_buf_2 _16849_ (.A(net673),
    .X(_10054_));
 sg13g2_nand2_1 _16850_ (.Y(_10055_),
    .A(net695),
    .B(_09394_));
 sg13g2_buf_1 _16851_ (.A(_10055_),
    .X(_10056_));
 sg13g2_buf_2 _16852_ (.A(_09206_),
    .X(_10057_));
 sg13g2_and2_1 _16853_ (.A(net1028),
    .B(_10000_),
    .X(_10058_));
 sg13g2_buf_1 _16854_ (.A(_10058_),
    .X(_10059_));
 sg13g2_nand2b_1 _16855_ (.Y(_10060_),
    .B(_10059_),
    .A_N(_09261_));
 sg13g2_buf_1 _16856_ (.A(_10060_),
    .X(_10061_));
 sg13g2_nor3_1 _16857_ (.A(net616),
    .B(net539),
    .C(_10061_),
    .Y(_10062_));
 sg13g2_buf_2 _16858_ (.A(_10062_),
    .X(_10063_));
 sg13g2_buf_1 _16859_ (.A(_10063_),
    .X(_10064_));
 sg13g2_mux2_1 _16860_ (.A0(_10046_),
    .A1(_10049_),
    .S(net104),
    .X(_00062_));
 sg13g2_inv_1 _16861_ (.Y(_10065_),
    .A(_10005_));
 sg13g2_o21ai_1 _16862_ (.B1(_09964_),
    .Y(_10066_),
    .A1(_09965_),
    .A2(_09980_));
 sg13g2_nand2b_1 _16863_ (.Y(_10067_),
    .B(_10066_),
    .A_N(_09981_));
 sg13g2_o21ai_1 _16864_ (.B1(_10067_),
    .Y(_10068_),
    .A1(\cpu.intr.r_timer_reload[17] ),
    .A2(_09991_));
 sg13g2_buf_1 _16865_ (.A(\cpu.dcache.wdata[1] ),
    .X(_10069_));
 sg13g2_buf_1 _16866_ (.A(_10069_),
    .X(_10070_));
 sg13g2_nand2_1 _16867_ (.Y(_10071_),
    .A(net1027),
    .B(_10063_));
 sg13g2_o21ai_1 _16868_ (.B1(_10071_),
    .Y(_00063_),
    .A1(_10065_),
    .A2(_10068_));
 sg13g2_xor2_1 _16869_ (.B(_09981_),
    .A(_09963_),
    .X(_10072_));
 sg13g2_o21ai_1 _16870_ (.B1(_10072_),
    .Y(_10073_),
    .A1(\cpu.intr.r_timer_reload[18] ),
    .A2(_09991_));
 sg13g2_buf_1 _16871_ (.A(\cpu.dcache.wdata[2] ),
    .X(_10074_));
 sg13g2_buf_1 _16872_ (.A(_10074_),
    .X(_10075_));
 sg13g2_nand2_1 _16873_ (.Y(_10076_),
    .A(net1026),
    .B(_10063_));
 sg13g2_o21ai_1 _16874_ (.B1(_10076_),
    .Y(_00064_),
    .A1(_10065_),
    .A2(_10073_));
 sg13g2_xor2_1 _16875_ (.B(_09982_),
    .A(_09962_),
    .X(_10077_));
 sg13g2_o21ai_1 _16876_ (.B1(_10077_),
    .Y(_10078_),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .A2(_09991_));
 sg13g2_buf_1 _16877_ (.A(\cpu.dcache.wdata[3] ),
    .X(_10079_));
 sg13g2_buf_1 _16878_ (.A(net1113),
    .X(_10080_));
 sg13g2_nand2_1 _16879_ (.Y(_10081_),
    .A(_10080_),
    .B(_10063_));
 sg13g2_o21ai_1 _16880_ (.B1(_10081_),
    .Y(_00065_),
    .A1(net104),
    .A2(_10078_));
 sg13g2_nor2b_1 _16881_ (.A(\cpu.intr.r_timer_reload[20] ),
    .B_N(_09989_),
    .Y(_10082_));
 sg13g2_nor3_1 _16882_ (.A(_09986_),
    .B(_09984_),
    .C(_10082_),
    .Y(_10083_));
 sg13g2_a21oi_1 _16883_ (.A1(_09986_),
    .A2(_09984_),
    .Y(_10084_),
    .B1(_10083_));
 sg13g2_buf_2 _16884_ (.A(\cpu.dcache.wdata[4] ),
    .X(_10085_));
 sg13g2_buf_1 _16885_ (.A(_10085_),
    .X(_10086_));
 sg13g2_nor2_1 _16886_ (.A(net1024),
    .B(_10005_),
    .Y(_10087_));
 sg13g2_a21oi_1 _16887_ (.A1(_10005_),
    .A2(_10084_),
    .Y(_00067_),
    .B1(_10087_));
 sg13g2_nor2_1 _16888_ (.A(_09986_),
    .B(_09984_),
    .Y(_10088_));
 sg13g2_xor2_1 _16889_ (.B(_10088_),
    .A(_09985_),
    .X(_10089_));
 sg13g2_o21ai_1 _16890_ (.B1(_10089_),
    .Y(_10090_),
    .A1(\cpu.intr.r_timer_reload[21] ),
    .A2(_09991_));
 sg13g2_buf_2 _16891_ (.A(\cpu.dcache.wdata[5] ),
    .X(_10091_));
 sg13g2_buf_1 _16892_ (.A(_10091_),
    .X(_10092_));
 sg13g2_nand2_1 _16893_ (.Y(_10093_),
    .A(_10092_),
    .B(_10063_));
 sg13g2_o21ai_1 _16894_ (.B1(_10093_),
    .Y(_00068_),
    .A1(_10065_),
    .A2(_10090_));
 sg13g2_nor3_1 _16895_ (.A(_09985_),
    .B(_09986_),
    .C(_09984_),
    .Y(_10094_));
 sg13g2_xor2_1 _16896_ (.B(_10094_),
    .A(_09988_),
    .X(_10095_));
 sg13g2_o21ai_1 _16897_ (.B1(_10095_),
    .Y(_10096_),
    .A1(\cpu.intr.r_timer_reload[22] ),
    .A2(_09991_));
 sg13g2_buf_2 _16898_ (.A(\cpu.dcache.wdata[6] ),
    .X(_10097_));
 sg13g2_buf_1 _16899_ (.A(_10097_),
    .X(_10098_));
 sg13g2_nand2_1 _16900_ (.Y(_10099_),
    .A(net1022),
    .B(_10063_));
 sg13g2_o21ai_1 _16901_ (.B1(_10099_),
    .Y(_00069_),
    .A1(_10065_),
    .A2(_10096_));
 sg13g2_nor2b_1 _16902_ (.A(_09987_),
    .B_N(\cpu.intr.r_timer_reload[23] ),
    .Y(_10100_));
 sg13g2_nor2b_1 _16903_ (.A(_09988_),
    .B_N(_10094_),
    .Y(_10101_));
 sg13g2_mux2_1 _16904_ (.A0(_09987_),
    .A1(_10100_),
    .S(_10101_),
    .X(_10102_));
 sg13g2_buf_2 _16905_ (.A(\cpu.dcache.wdata[7] ),
    .X(_10103_));
 sg13g2_buf_1 _16906_ (.A(_10103_),
    .X(_10104_));
 sg13g2_buf_1 _16907_ (.A(net1021),
    .X(_10105_));
 sg13g2_mux2_1 _16908_ (.A0(_10102_),
    .A1(net888),
    .S(_10064_),
    .X(_00070_));
 sg13g2_buf_1 _16909_ (.A(net674),
    .X(_10106_));
 sg13g2_buf_1 _16910_ (.A(net615),
    .X(_10107_));
 sg13g2_nor2b_1 _16911_ (.A(net538),
    .B_N(net1029),
    .Y(_10108_));
 sg13g2_nand2_1 _16912_ (.Y(_10109_),
    .A(_09341_),
    .B(_09416_));
 sg13g2_buf_2 _16913_ (.A(_10109_),
    .X(_10110_));
 sg13g2_nor2_1 _16914_ (.A(_10110_),
    .B(_10061_),
    .Y(_10111_));
 sg13g2_buf_2 _16915_ (.A(_10111_),
    .X(_10112_));
 sg13g2_buf_1 _16916_ (.A(_10112_),
    .X(_10113_));
 sg13g2_mux2_1 _16917_ (.A0(_00284_),
    .A1(_10108_),
    .S(net103),
    .X(_00036_));
 sg13g2_inv_1 _16918_ (.Y(_10114_),
    .A(_10069_));
 sg13g2_buf_1 _16919_ (.A(_10114_),
    .X(_10115_));
 sg13g2_buf_1 _16920_ (.A(net887),
    .X(_10116_));
 sg13g2_nand2_1 _16921_ (.Y(_10117_),
    .A(net616),
    .B(_10112_));
 sg13g2_buf_1 _16922_ (.A(_10117_),
    .X(_10118_));
 sg13g2_nor2_1 _16923_ (.A(net783),
    .B(_10050_),
    .Y(_10119_));
 sg13g2_buf_2 _16924_ (.A(_10119_),
    .X(_10120_));
 sg13g2_and2_1 _16925_ (.A(_09595_),
    .B(_10120_),
    .X(_10121_));
 sg13g2_buf_1 _16926_ (.A(_10121_),
    .X(_10122_));
 sg13g2_buf_1 _16927_ (.A(_10122_),
    .X(_10123_));
 sg13g2_buf_1 _16928_ (.A(_10123_),
    .X(_10124_));
 sg13g2_nand2_1 _16929_ (.Y(_10125_),
    .A(net171),
    .B(net373));
 sg13g2_buf_1 _16930_ (.A(_10125_),
    .X(_10126_));
 sg13g2_buf_1 _16931_ (.A(_10126_),
    .X(_10127_));
 sg13g2_buf_2 _16932_ (.A(\cpu.intr.r_clock_count[0] ),
    .X(_10128_));
 sg13g2_buf_2 _16933_ (.A(\cpu.intr.r_clock_count[1] ),
    .X(_10129_));
 sg13g2_xor2_1 _16934_ (.B(_10129_),
    .A(_10128_),
    .X(_10130_));
 sg13g2_nand3_1 _16935_ (.B(net102),
    .C(_10130_),
    .A(_10118_),
    .Y(_10131_));
 sg13g2_o21ai_1 _16936_ (.B1(_10131_),
    .Y(_00043_),
    .A1(net762),
    .A2(_10118_));
 sg13g2_buf_1 _16937_ (.A(_10074_),
    .X(_10132_));
 sg13g2_buf_1 _16938_ (.A(net1020),
    .X(_10133_));
 sg13g2_buf_1 _16939_ (.A(_09993_),
    .X(_10134_));
 sg13g2_nor3_1 _16940_ (.A(net537),
    .B(_10110_),
    .C(_10061_),
    .Y(_10135_));
 sg13g2_buf_1 _16941_ (.A(_10135_),
    .X(_10136_));
 sg13g2_buf_1 _16942_ (.A(net116),
    .X(_10137_));
 sg13g2_and2_1 _16943_ (.A(net171),
    .B(net412),
    .X(_10138_));
 sg13g2_buf_1 _16944_ (.A(_10138_),
    .X(_10139_));
 sg13g2_buf_1 _16945_ (.A(_10139_),
    .X(_10140_));
 sg13g2_buf_1 _16946_ (.A(net100),
    .X(_10141_));
 sg13g2_buf_1 _16947_ (.A(\cpu.intr.r_clock_count[2] ),
    .X(_10142_));
 sg13g2_nand2_1 _16948_ (.Y(_10143_),
    .A(_10128_),
    .B(_10129_));
 sg13g2_xor2_1 _16949_ (.B(_10143_),
    .A(_10142_),
    .X(_10144_));
 sg13g2_nor3_1 _16950_ (.A(net101),
    .B(net86),
    .C(_10144_),
    .Y(_10145_));
 sg13g2_a21o_1 _16951_ (.A2(net101),
    .A1(net886),
    .B1(_10145_),
    .X(_00044_));
 sg13g2_buf_1 _16952_ (.A(net1025),
    .X(_10146_));
 sg13g2_buf_1 _16953_ (.A(\cpu.intr.r_clock_count[3] ),
    .X(_10147_));
 sg13g2_nand2_1 _16954_ (.Y(_10148_),
    .A(_10129_),
    .B(_10142_));
 sg13g2_nor2_1 _16955_ (.A(_00284_),
    .B(_10148_),
    .Y(_10149_));
 sg13g2_xnor2_1 _16956_ (.Y(_10150_),
    .A(_10147_),
    .B(_10149_));
 sg13g2_nor3_1 _16957_ (.A(net116),
    .B(net86),
    .C(_10150_),
    .Y(_10151_));
 sg13g2_a21o_1 _16958_ (.A2(net101),
    .A1(net885),
    .B1(_10151_),
    .X(_00045_));
 sg13g2_buf_1 _16959_ (.A(_10086_),
    .X(_10152_));
 sg13g2_buf_2 _16960_ (.A(\cpu.intr.r_clock_count[4] ),
    .X(_10153_));
 sg13g2_and4_1 _16961_ (.A(_10128_),
    .B(_10129_),
    .C(_10142_),
    .D(_10147_),
    .X(_10154_));
 sg13g2_buf_1 _16962_ (.A(_10154_),
    .X(_10155_));
 sg13g2_xnor2_1 _16963_ (.Y(_10156_),
    .A(_10153_),
    .B(_10155_));
 sg13g2_nor3_1 _16964_ (.A(net116),
    .B(net86),
    .C(_10156_),
    .Y(_10157_));
 sg13g2_a21o_1 _16965_ (.A2(net101),
    .A1(net884),
    .B1(_10157_),
    .X(_00046_));
 sg13g2_buf_1 _16966_ (.A(_10092_),
    .X(_10158_));
 sg13g2_buf_2 _16967_ (.A(\cpu.intr.r_clock_count[5] ),
    .X(_10159_));
 sg13g2_and3_1 _16968_ (.X(_10160_),
    .A(_10147_),
    .B(_10153_),
    .C(_10149_));
 sg13g2_buf_1 _16969_ (.A(_10160_),
    .X(_10161_));
 sg13g2_xnor2_1 _16970_ (.Y(_10162_),
    .A(_10159_),
    .B(_10161_));
 sg13g2_nor3_1 _16971_ (.A(_10136_),
    .B(_10140_),
    .C(_10162_),
    .Y(_10163_));
 sg13g2_a21o_1 _16972_ (.A2(_10137_),
    .A1(net883),
    .B1(_10163_),
    .X(_00047_));
 sg13g2_buf_1 _16973_ (.A(net1022),
    .X(_10164_));
 sg13g2_buf_2 _16974_ (.A(\cpu.intr.r_clock_count[6] ),
    .X(_10165_));
 sg13g2_and2_1 _16975_ (.A(_10153_),
    .B(_10155_),
    .X(_10166_));
 sg13g2_buf_1 _16976_ (.A(_10166_),
    .X(_10167_));
 sg13g2_nand2_1 _16977_ (.Y(_10168_),
    .A(_10159_),
    .B(_10167_));
 sg13g2_xor2_1 _16978_ (.B(_10168_),
    .A(_10165_),
    .X(_10169_));
 sg13g2_nor3_1 _16979_ (.A(net116),
    .B(net100),
    .C(_10169_),
    .Y(_10170_));
 sg13g2_a21o_1 _16980_ (.A2(_10137_),
    .A1(net882),
    .B1(_10170_),
    .X(_00048_));
 sg13g2_buf_1 _16981_ (.A(\cpu.intr.r_clock_count[7] ),
    .X(_10171_));
 sg13g2_nand3_1 _16982_ (.B(_10165_),
    .C(_10161_),
    .A(_10159_),
    .Y(_10172_));
 sg13g2_xor2_1 _16983_ (.B(_10172_),
    .A(_10171_),
    .X(_10173_));
 sg13g2_nor3_1 _16984_ (.A(net116),
    .B(net100),
    .C(_10173_),
    .Y(_10174_));
 sg13g2_a21o_1 _16985_ (.A2(net101),
    .A1(net888),
    .B1(_10174_),
    .X(_00049_));
 sg13g2_buf_2 _16986_ (.A(\cpu.intr.r_clock_count[8] ),
    .X(_10175_));
 sg13g2_nand2_1 _16987_ (.Y(_10176_),
    .A(_10153_),
    .B(_10155_));
 sg13g2_nand3_1 _16988_ (.B(_10165_),
    .C(_10171_),
    .A(_10159_),
    .Y(_10177_));
 sg13g2_nor2_1 _16989_ (.A(_10176_),
    .B(_10177_),
    .Y(_10178_));
 sg13g2_xnor2_1 _16990_ (.Y(_10179_),
    .A(_10175_),
    .B(_10178_));
 sg13g2_buf_1 _16991_ (.A(net616),
    .X(_10180_));
 sg13g2_buf_2 _16992_ (.A(\cpu.dcache.wdata[8] ),
    .X(_10181_));
 sg13g2_nand3_1 _16993_ (.B(_10181_),
    .C(_10113_),
    .A(net536),
    .Y(_10182_));
 sg13g2_o21ai_1 _16994_ (.B1(_10182_),
    .Y(_00050_),
    .A1(_10113_),
    .A2(_10179_));
 sg13g2_buf_2 _16995_ (.A(\cpu.intr.r_clock_count[9] ),
    .X(_10183_));
 sg13g2_nand2_1 _16996_ (.Y(_10184_),
    .A(_10175_),
    .B(_10178_));
 sg13g2_xor2_1 _16997_ (.B(_10184_),
    .A(_10183_),
    .X(_10185_));
 sg13g2_buf_2 _16998_ (.A(\cpu.dcache.wdata[9] ),
    .X(_10186_));
 sg13g2_nand3_1 _16999_ (.B(_10186_),
    .C(net103),
    .A(net536),
    .Y(_10187_));
 sg13g2_o21ai_1 _17000_ (.B1(_10187_),
    .Y(_00051_),
    .A1(net103),
    .A2(_10185_));
 sg13g2_buf_1 _17001_ (.A(\cpu.intr.r_clock_count[10] ),
    .X(_10188_));
 sg13g2_nand3_1 _17002_ (.B(_10183_),
    .C(_10178_),
    .A(_10175_),
    .Y(_10189_));
 sg13g2_xor2_1 _17003_ (.B(_10189_),
    .A(_10188_),
    .X(_10190_));
 sg13g2_buf_2 _17004_ (.A(\cpu.dcache.wdata[10] ),
    .X(_10191_));
 sg13g2_nand3_1 _17005_ (.B(_10191_),
    .C(_10112_),
    .A(net536),
    .Y(_10192_));
 sg13g2_o21ai_1 _17006_ (.B1(_10192_),
    .Y(_00037_),
    .A1(net103),
    .A2(_10190_));
 sg13g2_buf_2 _17007_ (.A(\cpu.intr.r_clock_count[11] ),
    .X(_10193_));
 sg13g2_nand3_1 _17008_ (.B(_10183_),
    .C(_10188_),
    .A(_10175_),
    .Y(_10194_));
 sg13g2_nor2_1 _17009_ (.A(_10177_),
    .B(_10194_),
    .Y(_10195_));
 sg13g2_and2_1 _17010_ (.A(_10161_),
    .B(_10195_),
    .X(_10196_));
 sg13g2_xnor2_1 _17011_ (.Y(_10197_),
    .A(_10193_),
    .B(_10196_));
 sg13g2_buf_2 _17012_ (.A(\cpu.dcache.wdata[11] ),
    .X(_10198_));
 sg13g2_nand3_1 _17013_ (.B(_10198_),
    .C(_10112_),
    .A(net536),
    .Y(_10199_));
 sg13g2_o21ai_1 _17014_ (.B1(_10199_),
    .Y(_00038_),
    .A1(net103),
    .A2(_10197_));
 sg13g2_buf_1 _17015_ (.A(\cpu.intr.r_clock_count[12] ),
    .X(_10200_));
 sg13g2_nand3_1 _17016_ (.B(_10167_),
    .C(_10195_),
    .A(_10193_),
    .Y(_10201_));
 sg13g2_xor2_1 _17017_ (.B(_10201_),
    .A(_10200_),
    .X(_10202_));
 sg13g2_buf_2 _17018_ (.A(\cpu.dcache.wdata[12] ),
    .X(_10203_));
 sg13g2_nand3_1 _17019_ (.B(_10203_),
    .C(_10112_),
    .A(net536),
    .Y(_10204_));
 sg13g2_o21ai_1 _17020_ (.B1(_10204_),
    .Y(_00039_),
    .A1(net103),
    .A2(_10202_));
 sg13g2_buf_2 _17021_ (.A(\cpu.dcache.wdata[13] ),
    .X(_10205_));
 sg13g2_buf_1 _17022_ (.A(\cpu.intr.r_clock_count[13] ),
    .X(_10206_));
 sg13g2_nand4_1 _17023_ (.B(_10200_),
    .C(_10161_),
    .A(_10193_),
    .Y(_10207_),
    .D(_10195_));
 sg13g2_xor2_1 _17024_ (.B(_10207_),
    .A(_10206_),
    .X(_10208_));
 sg13g2_nor3_1 _17025_ (.A(net116),
    .B(net100),
    .C(_10208_),
    .Y(_10209_));
 sg13g2_a21o_1 _17026_ (.A2(net101),
    .A1(_10205_),
    .B1(_10209_),
    .X(_00040_));
 sg13g2_buf_2 _17027_ (.A(\cpu.intr.r_clock_count[14] ),
    .X(_10210_));
 sg13g2_and4_1 _17028_ (.A(_10193_),
    .B(_10200_),
    .C(_10206_),
    .D(_10195_),
    .X(_10211_));
 sg13g2_buf_1 _17029_ (.A(_10211_),
    .X(_10212_));
 sg13g2_nand2_1 _17030_ (.Y(_10213_),
    .A(_10167_),
    .B(_10212_));
 sg13g2_xor2_1 _17031_ (.B(_10213_),
    .A(_10210_),
    .X(_10214_));
 sg13g2_buf_2 _17032_ (.A(\cpu.dcache.wdata[14] ),
    .X(_10215_));
 sg13g2_nand3_1 _17033_ (.B(_10215_),
    .C(_10112_),
    .A(net536),
    .Y(_10216_));
 sg13g2_o21ai_1 _17034_ (.B1(_10216_),
    .Y(_00041_),
    .A1(net103),
    .A2(_10214_));
 sg13g2_buf_2 _17035_ (.A(\cpu.intr.r_clock_count[15] ),
    .X(_10217_));
 sg13g2_nand3_1 _17036_ (.B(_10161_),
    .C(_10212_),
    .A(_10210_),
    .Y(_10218_));
 sg13g2_xor2_1 _17037_ (.B(_10218_),
    .A(_10217_),
    .X(_10219_));
 sg13g2_buf_2 _17038_ (.A(\cpu.dcache.wdata[15] ),
    .X(_10220_));
 sg13g2_nand3_1 _17039_ (.B(_10220_),
    .C(_10112_),
    .A(net536),
    .Y(_10221_));
 sg13g2_o21ai_1 _17040_ (.B1(_10221_),
    .Y(_00042_),
    .A1(net103),
    .A2(_10219_));
 sg13g2_buf_1 _17041_ (.A(\cpu.ex.r_wb_valid ),
    .X(_10222_));
 sg13g2_buf_1 _17042_ (.A(\cpu.ex.r_set_cc ),
    .X(_10223_));
 sg13g2_inv_1 _17043_ (.Y(_10224_),
    .A(net1112));
 sg13g2_buf_1 _17044_ (.A(\cpu.ex.r_wb_addr[3] ),
    .X(_10225_));
 sg13g2_inv_1 _17045_ (.Y(_10226_),
    .A(net1111));
 sg13g2_buf_1 _17046_ (.A(\cpu.ex.r_wb_addr[2] ),
    .X(_10227_));
 sg13g2_nand2_1 _17047_ (.Y(_10228_),
    .A(_10226_),
    .B(net1110));
 sg13g2_buf_2 _17048_ (.A(\cpu.ex.r_wb_addr[1] ),
    .X(_10229_));
 sg13g2_buf_8 _17049_ (.A(_10229_),
    .X(_10230_));
 sg13g2_buf_1 _17050_ (.A(\cpu.ex.r_wb_addr[0] ),
    .X(_10231_));
 sg13g2_buf_1 _17051_ (.A(_10231_),
    .X(_10232_));
 sg13g2_nand2_1 _17052_ (.Y(_10233_),
    .A(net1019),
    .B(net1018));
 sg13g2_nor3_1 _17053_ (.A(_10224_),
    .B(_10228_),
    .C(_10233_),
    .Y(_10234_));
 sg13g2_a21o_1 _17054_ (.A2(_10223_),
    .A1(net1112),
    .B1(_10234_),
    .X(_10235_));
 sg13g2_buf_2 _17055_ (.A(_10235_),
    .X(_10236_));
 sg13g2_buf_1 _17056_ (.A(_10236_),
    .X(_10237_));
 sg13g2_buf_1 _17057_ (.A(net677),
    .X(_10238_));
 sg13g2_nor4_1 _17058_ (.A(_10230_),
    .B(_10231_),
    .C(net1111),
    .D(net1110),
    .Y(_10239_));
 sg13g2_nand2b_1 _17059_ (.Y(_10240_),
    .B(net1112),
    .A_N(_10239_));
 sg13g2_buf_2 _17060_ (.A(\cpu.dec.r_rs2[2] ),
    .X(_10241_));
 sg13g2_xnor2_1 _17061_ (.Y(_10242_),
    .A(net1110),
    .B(_10241_));
 sg13g2_buf_2 _17062_ (.A(\cpu.dec.r_rs2[0] ),
    .X(_10243_));
 sg13g2_xnor2_1 _17063_ (.Y(_10244_),
    .A(_10231_),
    .B(_10243_));
 sg13g2_buf_2 _17064_ (.A(\cpu.dec.r_rs2[3] ),
    .X(_10245_));
 sg13g2_xnor2_1 _17065_ (.Y(_10246_),
    .A(net1111),
    .B(_10245_));
 sg13g2_buf_8 _17066_ (.A(\cpu.dec.r_rs2[1] ),
    .X(_10247_));
 sg13g2_xnor2_1 _17067_ (.Y(_10248_),
    .A(_10229_),
    .B(_10247_));
 sg13g2_nand4_1 _17068_ (.B(_10244_),
    .C(_10246_),
    .A(_10242_),
    .Y(_10249_),
    .D(_10248_));
 sg13g2_buf_1 _17069_ (.A(_10249_),
    .X(_10250_));
 sg13g2_nor2_1 _17070_ (.A(_10240_),
    .B(_10250_),
    .Y(_10251_));
 sg13g2_buf_8 _17071_ (.A(_10251_),
    .X(_10252_));
 sg13g2_buf_1 _17072_ (.A(net613),
    .X(_10253_));
 sg13g2_buf_8 _17073_ (.A(_10247_),
    .X(_10254_));
 sg13g2_buf_8 _17074_ (.A(net1017),
    .X(_10255_));
 sg13g2_buf_8 _17075_ (.A(net881),
    .X(_10256_));
 sg13g2_buf_8 _17076_ (.A(_10256_),
    .X(_10257_));
 sg13g2_buf_1 _17077_ (.A(net672),
    .X(_10258_));
 sg13g2_buf_8 _17078_ (.A(_10243_),
    .X(_10259_));
 sg13g2_inv_2 _17079_ (.Y(_10260_),
    .A(net1016));
 sg13g2_buf_1 _17080_ (.A(_10260_),
    .X(_10261_));
 sg13g2_buf_1 _17081_ (.A(net760),
    .X(_10262_));
 sg13g2_buf_8 _17082_ (.A(_10245_),
    .X(_10263_));
 sg13g2_nor2b_1 _17083_ (.A(_10241_),
    .B_N(net1015),
    .Y(_10264_));
 sg13g2_buf_1 _17084_ (.A(_10264_),
    .X(_10265_));
 sg13g2_buf_1 _17085_ (.A(_10265_),
    .X(_10266_));
 sg13g2_nor2b_1 _17086_ (.A(_10245_),
    .B_N(_10241_),
    .Y(_10267_));
 sg13g2_buf_1 _17087_ (.A(_10267_),
    .X(_10268_));
 sg13g2_buf_2 _17088_ (.A(\cpu.ex.r_mult[29] ),
    .X(_10269_));
 sg13g2_a22oi_1 _17089_ (.Y(_10270_),
    .B1(net880),
    .B2(_10269_),
    .A2(net670),
    .A1(\cpu.ex.r_11[13] ));
 sg13g2_nand3_1 _17090_ (.B(net671),
    .C(net880),
    .A(\cpu.ex.r_stmp[13] ),
    .Y(_10271_));
 sg13g2_o21ai_1 _17091_ (.B1(_10271_),
    .Y(_10272_),
    .A1(net671),
    .A2(_10270_));
 sg13g2_buf_8 _17092_ (.A(_10241_),
    .X(_10273_));
 sg13g2_nand3_1 _17093_ (.B(_10254_),
    .C(net1014),
    .A(_10243_),
    .Y(_10274_));
 sg13g2_buf_1 _17094_ (.A(_10274_),
    .X(_10275_));
 sg13g2_buf_2 _17095_ (.A(net1016),
    .X(_10276_));
 sg13g2_buf_8 _17096_ (.A(net879),
    .X(_10277_));
 sg13g2_buf_1 _17097_ (.A(net1014),
    .X(_10278_));
 sg13g2_buf_8 _17098_ (.A(net878),
    .X(_10279_));
 sg13g2_nor3_1 _17099_ (.A(net759),
    .B(net672),
    .C(net758),
    .Y(_10280_));
 sg13g2_nand2_1 _17100_ (.Y(_10281_),
    .A(\cpu.ex.r_8[13] ),
    .B(_10280_));
 sg13g2_o21ai_1 _17101_ (.B1(_10281_),
    .Y(_10282_),
    .A1(_00269_),
    .A2(_10275_));
 sg13g2_buf_8 _17102_ (.A(net1015),
    .X(_10283_));
 sg13g2_buf_8 _17103_ (.A(net877),
    .X(_10284_));
 sg13g2_buf_8 _17104_ (.A(net757),
    .X(_10285_));
 sg13g2_buf_1 _17105_ (.A(net669),
    .X(_10286_));
 sg13g2_buf_1 _17106_ (.A(_10278_),
    .X(_10287_));
 sg13g2_buf_1 _17107_ (.A(net756),
    .X(_10288_));
 sg13g2_nor2b_1 _17108_ (.A(_10243_),
    .B_N(_10247_),
    .Y(_10289_));
 sg13g2_buf_2 _17109_ (.A(_10289_),
    .X(_10290_));
 sg13g2_buf_1 _17110_ (.A(_10290_),
    .X(_10291_));
 sg13g2_mux2_1 _17111_ (.A0(\cpu.ex.r_sp[13] ),
    .A1(\cpu.ex.r_10[13] ),
    .S(net611),
    .X(_10292_));
 sg13g2_nor2_1 _17112_ (.A(_10247_),
    .B(_10245_),
    .Y(_10293_));
 sg13g2_buf_2 _17113_ (.A(_10293_),
    .X(_10294_));
 sg13g2_buf_1 _17114_ (.A(net759),
    .X(_10295_));
 sg13g2_buf_1 _17115_ (.A(net667),
    .X(_10296_));
 sg13g2_and2_1 _17116_ (.A(\cpu.ex.r_lr[13] ),
    .B(net610),
    .X(_10297_));
 sg13g2_a22oi_1 _17117_ (.Y(_10298_),
    .B1(_10294_),
    .B2(_10297_),
    .A2(_10292_),
    .A1(net755));
 sg13g2_nor2b_2 _17118_ (.A(net879),
    .B_N(net877),
    .Y(_10299_));
 sg13g2_mux2_1 _17119_ (.A0(\cpu.ex.r_12[13] ),
    .A1(\cpu.ex.r_14[13] ),
    .S(net612),
    .X(_10300_));
 sg13g2_nand3_1 _17120_ (.B(_10299_),
    .C(_10300_),
    .A(net668),
    .Y(_10301_));
 sg13g2_o21ai_1 _17121_ (.B1(_10301_),
    .Y(_10302_),
    .A1(net668),
    .A2(_10298_));
 sg13g2_a221oi_1 _17122_ (.B2(net611),
    .C1(_10302_),
    .B1(_10282_),
    .A1(net612),
    .Y(_10303_),
    .A2(_10272_));
 sg13g2_buf_1 _17123_ (.A(\cpu.ex.mmu_read[13] ),
    .X(_10304_));
 sg13g2_mux2_1 _17124_ (.A0(_10304_),
    .A1(\cpu.ex.r_13[13] ),
    .S(net611),
    .X(_10305_));
 sg13g2_a22oi_1 _17125_ (.Y(_10306_),
    .B1(_10305_),
    .B2(net668),
    .A2(net670),
    .A1(\cpu.ex.r_9[13] ));
 sg13g2_nor2_1 _17126_ (.A(_10263_),
    .B(net1014),
    .Y(_10307_));
 sg13g2_buf_2 _17127_ (.A(_10307_),
    .X(_10308_));
 sg13g2_nand3_1 _17128_ (.B(net612),
    .C(_10308_),
    .A(\cpu.ex.r_epc[13] ),
    .Y(_10309_));
 sg13g2_o21ai_1 _17129_ (.B1(_10309_),
    .Y(_10310_),
    .A1(net612),
    .A2(_10306_));
 sg13g2_nand2_1 _17130_ (.Y(_10311_),
    .A(net610),
    .B(_10310_));
 sg13g2_nor2_1 _17131_ (.A(net1016),
    .B(net1017),
    .Y(_10312_));
 sg13g2_nand2_1 _17132_ (.Y(_10313_),
    .A(_10308_),
    .B(_10312_));
 sg13g2_o21ai_1 _17133_ (.B1(_10313_),
    .Y(_10314_),
    .A1(_10240_),
    .A2(_10250_));
 sg13g2_buf_2 _17134_ (.A(_10314_),
    .X(_10315_));
 sg13g2_a21oi_1 _17135_ (.A1(_10303_),
    .A2(_10311_),
    .Y(_10316_),
    .B1(_10315_));
 sg13g2_a21o_1 _17136_ (.A2(net534),
    .A1(net614),
    .B1(_10316_),
    .X(_10317_));
 sg13g2_buf_1 _17137_ (.A(\cpu.dec.needs_rs2 ),
    .X(_10318_));
 sg13g2_buf_1 _17138_ (.A(_10318_),
    .X(_10319_));
 sg13g2_mux2_1 _17139_ (.A0(\cpu.dec.imm[13] ),
    .A1(_10317_),
    .S(net1013),
    .X(_10320_));
 sg13g2_buf_1 _17140_ (.A(\cpu.dec.r_rs2_pc ),
    .X(_10321_));
 sg13g2_buf_2 _17141_ (.A(\cpu.dec.r_rs2_inv ),
    .X(_10322_));
 sg13g2_or2_1 _17142_ (.X(_10323_),
    .B(_10322_),
    .A(_10321_));
 sg13g2_buf_1 _17143_ (.A(_10323_),
    .X(_10324_));
 sg13g2_buf_1 _17144_ (.A(_10321_),
    .X(_10325_));
 sg13g2_buf_1 _17145_ (.A(net1012),
    .X(_10326_));
 sg13g2_nand2b_1 _17146_ (.Y(_10327_),
    .B(net876),
    .A_N(net912));
 sg13g2_o21ai_1 _17147_ (.B1(_10327_),
    .Y(_10328_),
    .A1(_10320_),
    .A2(_10324_));
 sg13g2_buf_1 _17148_ (.A(_10328_),
    .X(_10329_));
 sg13g2_buf_1 _17149_ (.A(_10329_),
    .X(_10330_));
 sg13g2_buf_2 _17150_ (.A(_00298_),
    .X(_10331_));
 sg13g2_nor2_1 _17151_ (.A(_10224_),
    .B(_10239_),
    .Y(_10332_));
 sg13g2_and4_1 _17152_ (.A(_10242_),
    .B(_10244_),
    .C(_10246_),
    .D(_10248_),
    .X(_10333_));
 sg13g2_a22oi_1 _17153_ (.Y(_10334_),
    .B1(_10308_),
    .B2(_10312_),
    .A2(_10333_),
    .A1(_10332_));
 sg13g2_buf_2 _17154_ (.A(_10334_),
    .X(_10335_));
 sg13g2_buf_8 _17155_ (.A(_10335_),
    .X(_10336_));
 sg13g2_nand3b_1 _17156_ (.B(net669),
    .C(\cpu.ex.r_14[12] ),
    .Y(_10337_),
    .A_N(net667));
 sg13g2_buf_1 _17157_ (.A(\cpu.ex.r_mult[28] ),
    .X(_10338_));
 sg13g2_nand3b_1 _17158_ (.B(net667),
    .C(_10338_),
    .Y(_10339_),
    .A_N(net669));
 sg13g2_inv_1 _17159_ (.Y(_10340_),
    .A(_10254_));
 sg13g2_buf_1 _17160_ (.A(_10340_),
    .X(_10341_));
 sg13g2_a21o_1 _17161_ (.A2(_10339_),
    .A1(_10337_),
    .B1(net754),
    .X(_10342_));
 sg13g2_nor2b_1 _17162_ (.A(_10247_),
    .B_N(_10245_),
    .Y(_10343_));
 sg13g2_buf_2 _17163_ (.A(_10343_),
    .X(_10344_));
 sg13g2_buf_8 _17164_ (.A(_10344_),
    .X(_10345_));
 sg13g2_nand3_1 _17165_ (.B(net610),
    .C(net753),
    .A(\cpu.ex.r_13[12] ),
    .Y(_10346_));
 sg13g2_nor2b_1 _17166_ (.A(_10245_),
    .B_N(_10247_),
    .Y(_10347_));
 sg13g2_buf_1 _17167_ (.A(_10347_),
    .X(_10348_));
 sg13g2_nand3_1 _17168_ (.B(net671),
    .C(net875),
    .A(\cpu.ex.r_stmp[12] ),
    .Y(_10349_));
 sg13g2_and4_1 _17169_ (.A(net668),
    .B(_10342_),
    .C(_10346_),
    .D(_10349_),
    .X(_10350_));
 sg13g2_inv_1 _17170_ (.Y(_10351_),
    .A(net1014));
 sg13g2_buf_1 _17171_ (.A(_10351_),
    .X(_10352_));
 sg13g2_buf_1 _17172_ (.A(net752),
    .X(_10353_));
 sg13g2_nand3_1 _17173_ (.B(net671),
    .C(net753),
    .A(\cpu.ex.r_8[12] ),
    .Y(_10354_));
 sg13g2_inv_4 _17174_ (.A(_10263_),
    .Y(_10355_));
 sg13g2_and2_1 _17175_ (.A(_10243_),
    .B(net1017),
    .X(_10356_));
 sg13g2_buf_2 _17176_ (.A(_10356_),
    .X(_10357_));
 sg13g2_nand3_1 _17177_ (.B(_10355_),
    .C(_10357_),
    .A(\cpu.ex.r_epc[12] ),
    .Y(_10358_));
 sg13g2_nor2b_1 _17178_ (.A(net1017),
    .B_N(_10243_),
    .Y(_10359_));
 sg13g2_buf_1 _17179_ (.A(_10359_),
    .X(_10360_));
 sg13g2_mux2_1 _17180_ (.A0(\cpu.ex.r_lr[12] ),
    .A1(\cpu.ex.r_9[12] ),
    .S(net669),
    .X(_10361_));
 sg13g2_nand2_1 _17181_ (.Y(_10362_),
    .A(net751),
    .B(_10361_));
 sg13g2_and4_1 _17182_ (.A(net666),
    .B(_10354_),
    .C(_10358_),
    .D(_10362_),
    .X(_10363_));
 sg13g2_nor2b_1 _17183_ (.A(_00268_),
    .B_N(net668),
    .Y(_10364_));
 sg13g2_nor2b_1 _17184_ (.A(net668),
    .B_N(\cpu.ex.r_11[12] ),
    .Y(_10365_));
 sg13g2_o21ai_1 _17185_ (.B1(net612),
    .Y(_10366_),
    .A1(_10364_),
    .A2(_10365_));
 sg13g2_nor2b_1 _17186_ (.A(_10241_),
    .B_N(_10247_),
    .Y(_10367_));
 sg13g2_buf_1 _17187_ (.A(_10367_),
    .X(_10368_));
 sg13g2_nor2b_2 _17188_ (.A(net761),
    .B_N(net878),
    .Y(_10369_));
 sg13g2_a22oi_1 _17189_ (.Y(_10370_),
    .B1(_10369_),
    .B2(\cpu.ex.r_12[12] ),
    .A2(_10368_),
    .A1(\cpu.ex.r_10[12] ));
 sg13g2_buf_1 _17190_ (.A(\cpu.ex.mmu_read[12] ),
    .X(_10371_));
 sg13g2_nand2_1 _17191_ (.Y(_10372_),
    .A(net1108),
    .B(_10369_));
 sg13g2_buf_1 _17192_ (.A(\cpu.ex.r_sp[12] ),
    .X(_10373_));
 sg13g2_nand2_1 _17193_ (.Y(_10374_),
    .A(_10373_),
    .B(_10368_));
 sg13g2_mux4_1 _17194_ (.S0(net671),
    .A0(_10366_),
    .A1(_10370_),
    .A2(_10372_),
    .A3(_10374_),
    .S1(_10355_),
    .X(_10375_));
 sg13g2_o21ai_1 _17195_ (.B1(_10375_),
    .Y(_10376_),
    .A1(_10350_),
    .A2(_10363_));
 sg13g2_a22oi_1 _17196_ (.Y(_10377_),
    .B1(net533),
    .B2(_10376_),
    .A2(net534),
    .A1(net620));
 sg13g2_nor2_1 _17197_ (.A(net1013),
    .B(\cpu.dec.imm[12] ),
    .Y(_10378_));
 sg13g2_a21oi_1 _17198_ (.A1(net1013),
    .A2(_10377_),
    .Y(_10379_),
    .B1(_10378_));
 sg13g2_nand2b_1 _17199_ (.Y(_10380_),
    .B(net876),
    .A_N(_08639_));
 sg13g2_o21ai_1 _17200_ (.B1(_10380_),
    .Y(_10381_),
    .A1(_10324_),
    .A2(_10379_));
 sg13g2_buf_2 _17201_ (.A(_10381_),
    .X(_10382_));
 sg13g2_inv_1 _17202_ (.Y(_10383_),
    .A(_10382_));
 sg13g2_inv_1 _17203_ (.Y(_10384_),
    .A(_10331_));
 sg13g2_nand2_1 _17204_ (.Y(_10385_),
    .A(_08768_),
    .B(net876));
 sg13g2_buf_1 _17205_ (.A(\cpu.addr[11] ),
    .X(_10386_));
 sg13g2_and2_1 _17206_ (.A(net1015),
    .B(net1014),
    .X(_10387_));
 sg13g2_buf_1 _17207_ (.A(_10387_),
    .X(_10388_));
 sg13g2_and2_1 _17208_ (.A(_10388_),
    .B(net755),
    .X(_10389_));
 sg13g2_buf_1 _17209_ (.A(net1014),
    .X(_10390_));
 sg13g2_and2_1 _17210_ (.A(net874),
    .B(_10344_),
    .X(_10391_));
 sg13g2_buf_1 _17211_ (.A(_10391_),
    .X(_10392_));
 sg13g2_mux2_1 _17212_ (.A0(\cpu.ex.r_12[11] ),
    .A1(\cpu.ex.r_13[11] ),
    .S(_10295_),
    .X(_10393_));
 sg13g2_a22oi_1 _17213_ (.Y(_10394_),
    .B1(_10392_),
    .B2(_10393_),
    .A2(_10389_),
    .A1(\cpu.ex.r_14[11] ));
 sg13g2_buf_1 _17214_ (.A(\cpu.ex.r_sp[11] ),
    .X(_10395_));
 sg13g2_mux2_1 _17215_ (.A0(_10395_),
    .A1(\cpu.ex.r_stmp[11] ),
    .S(_10287_),
    .X(_10396_));
 sg13g2_a22oi_1 _17216_ (.Y(_10397_),
    .B1(_10396_),
    .B2(_10355_),
    .A2(_10266_),
    .A1(\cpu.ex.r_10[11] ));
 sg13g2_nand2b_1 _17217_ (.Y(_10398_),
    .B(_10291_),
    .A_N(_10397_));
 sg13g2_and2_1 _17218_ (.A(\cpu.ex.r_8[11] ),
    .B(_10280_),
    .X(_10399_));
 sg13g2_nor2_1 _17219_ (.A(_00267_),
    .B(_10275_),
    .Y(_10400_));
 sg13g2_o21ai_1 _17220_ (.B1(net611),
    .Y(_10401_),
    .A1(_10399_),
    .A2(_10400_));
 sg13g2_inv_1 _17221_ (.Y(_10402_),
    .A(\cpu.ex.r_mult[27] ));
 sg13g2_nor4_1 _17222_ (.A(_10402_),
    .B(net754),
    .C(net611),
    .D(_10353_),
    .Y(_10403_));
 sg13g2_mux4_1 _17223_ (.S0(net672),
    .A0(\cpu.ex.r_lr[11] ),
    .A1(\cpu.ex.r_epc[11] ),
    .A2(\cpu.ex.r_9[11] ),
    .A3(\cpu.ex.r_11[11] ),
    .S1(net757),
    .X(_10404_));
 sg13g2_and2_1 _17224_ (.A(net666),
    .B(_10404_),
    .X(_10405_));
 sg13g2_o21ai_1 _17225_ (.B1(_10296_),
    .Y(_10406_),
    .A1(_10403_),
    .A2(_10405_));
 sg13g2_nand4_1 _17226_ (.B(_10398_),
    .C(_10401_),
    .A(_10394_),
    .Y(_10407_),
    .D(_10406_));
 sg13g2_inv_1 _17227_ (.Y(_10408_),
    .A(net1109));
 sg13g2_buf_1 _17228_ (.A(_10408_),
    .X(_10409_));
 sg13g2_a221oi_1 _17229_ (.B2(_10407_),
    .C1(net873),
    .B1(net533),
    .A1(net1107),
    .Y(_10410_),
    .A2(net534));
 sg13g2_nor2_1 _17230_ (.A(_10319_),
    .B(\cpu.dec.imm[11] ),
    .Y(_10411_));
 sg13g2_nor2_1 _17231_ (.A(_10321_),
    .B(_10322_),
    .Y(_10412_));
 sg13g2_buf_1 _17232_ (.A(_10412_),
    .X(_10413_));
 sg13g2_buf_1 _17233_ (.A(_10413_),
    .X(_10414_));
 sg13g2_o21ai_1 _17234_ (.B1(net750),
    .Y(_10415_),
    .A1(_10410_),
    .A2(_10411_));
 sg13g2_nand2_1 _17235_ (.Y(_10416_),
    .A(_10385_),
    .B(_10415_));
 sg13g2_buf_1 _17236_ (.A(_10416_),
    .X(_10417_));
 sg13g2_buf_1 _17237_ (.A(\cpu.ex.r_mult[26] ),
    .X(_10418_));
 sg13g2_a22oi_1 _17238_ (.Y(_10419_),
    .B1(_10417_),
    .B2(net1106),
    .A2(_10382_),
    .A1(_10384_));
 sg13g2_a21o_1 _17239_ (.A2(_10383_),
    .A1(_10331_),
    .B1(_10419_),
    .X(_10420_));
 sg13g2_buf_1 _17240_ (.A(_10420_),
    .X(_10421_));
 sg13g2_inv_1 _17241_ (.Y(_10422_),
    .A(_10421_));
 sg13g2_and2_1 _17242_ (.A(net170),
    .B(_10422_),
    .X(_10423_));
 sg13g2_buf_1 _17243_ (.A(_10338_),
    .X(_10424_));
 sg13g2_nand2b_1 _17244_ (.Y(_10425_),
    .B(_10421_),
    .A_N(net170));
 sg13g2_and2_1 _17245_ (.A(net1011),
    .B(_10425_),
    .X(_10426_));
 sg13g2_or3_1 _17246_ (.A(_09368_),
    .B(_09292_),
    .C(net1036),
    .X(_10427_));
 sg13g2_buf_1 _17247_ (.A(_10427_),
    .X(_10428_));
 sg13g2_o21ai_1 _17248_ (.B1(net749),
    .Y(_10429_),
    .A1(_10423_),
    .A2(_10426_));
 sg13g2_buf_1 _17249_ (.A(_10429_),
    .X(_10430_));
 sg13g2_nor2_1 _17250_ (.A(_10408_),
    .B(_10324_),
    .Y(_10431_));
 sg13g2_or2_1 _17251_ (.X(_10432_),
    .B(net874),
    .A(net877));
 sg13g2_buf_1 _17252_ (.A(_10432_),
    .X(_10433_));
 sg13g2_nor2_1 _17253_ (.A(net754),
    .B(_10433_),
    .Y(_10434_));
 sg13g2_a22oi_1 _17254_ (.Y(_10435_),
    .B1(_10434_),
    .B2(\cpu.ex.r_epc[3] ),
    .A2(_10392_),
    .A1(\cpu.ex.r_13[3] ));
 sg13g2_buf_1 _17255_ (.A(\cpu.ex.r_sp[3] ),
    .X(_10436_));
 sg13g2_a221oi_1 _17256_ (.B2(_10436_),
    .C1(net667),
    .B1(_10434_),
    .A1(\cpu.ex.r_12[3] ),
    .Y(_10437_),
    .A2(_10392_));
 sg13g2_a21oi_1 _17257_ (.A1(net667),
    .A2(_10435_),
    .Y(_10438_),
    .B1(_10437_));
 sg13g2_mux2_1 _17258_ (.A0(\cpu.ex.r_8[3] ),
    .A1(\cpu.ex.r_10[3] ),
    .S(net881),
    .X(_10439_));
 sg13g2_mux2_1 _17259_ (.A0(\cpu.ex.r_lr[3] ),
    .A1(\cpu.ex.r_9[3] ),
    .S(net877),
    .X(_10440_));
 sg13g2_a22oi_1 _17260_ (.Y(_10441_),
    .B1(_10440_),
    .B2(net751),
    .A2(_10439_),
    .A1(_10299_));
 sg13g2_nor2_1 _17261_ (.A(net756),
    .B(_10441_),
    .Y(_10442_));
 sg13g2_nand3_1 _17262_ (.B(_10388_),
    .C(_10290_),
    .A(\cpu.ex.r_14[3] ),
    .Y(_10443_));
 sg13g2_buf_1 _17263_ (.A(\cpu.ex.mmu_read[3] ),
    .X(_10444_));
 sg13g2_mux2_1 _17264_ (.A0(net1129),
    .A1(_10444_),
    .S(net879),
    .X(_10445_));
 sg13g2_nand3_1 _17265_ (.B(_10294_),
    .C(_10445_),
    .A(net758),
    .Y(_10446_));
 sg13g2_nand2_1 _17266_ (.Y(_10447_),
    .A(_10443_),
    .B(_10446_));
 sg13g2_nand2_1 _17267_ (.Y(_10448_),
    .A(net879),
    .B(_10255_));
 sg13g2_a22oi_1 _17268_ (.Y(_10449_),
    .B1(net880),
    .B2(\cpu.ex.r_mult[19] ),
    .A2(net670),
    .A1(\cpu.ex.r_11[3] ));
 sg13g2_nor2_1 _17269_ (.A(_10448_),
    .B(_10449_),
    .Y(_10450_));
 sg13g2_nor2_1 _17270_ (.A(net1016),
    .B(net1015),
    .Y(_10451_));
 sg13g2_buf_2 _17271_ (.A(_10451_),
    .X(_10452_));
 sg13g2_and2_1 _17272_ (.A(net879),
    .B(net877),
    .X(_10453_));
 sg13g2_buf_2 _17273_ (.A(_10453_),
    .X(_10454_));
 sg13g2_inv_1 _17274_ (.Y(_10455_),
    .A(_00259_));
 sg13g2_a22oi_1 _17275_ (.Y(_10456_),
    .B1(_10454_),
    .B2(_10455_),
    .A2(_10452_),
    .A1(\cpu.ex.r_stmp[3] ));
 sg13g2_and2_1 _17276_ (.A(net1017),
    .B(_10241_),
    .X(_10457_));
 sg13g2_buf_1 _17277_ (.A(_10457_),
    .X(_10458_));
 sg13g2_nor2b_1 _17278_ (.A(_10456_),
    .B_N(_10458_),
    .Y(_10459_));
 sg13g2_or4_1 _17279_ (.A(_10442_),
    .B(_10447_),
    .C(_10450_),
    .D(_10459_),
    .X(_10460_));
 sg13g2_o21ai_1 _17280_ (.B1(_10336_),
    .Y(_10461_),
    .A1(_10438_),
    .A2(_10460_));
 sg13g2_nand2_1 _17281_ (.Y(_10462_),
    .A(_09199_),
    .B(net613));
 sg13g2_nand3_1 _17282_ (.B(_10461_),
    .C(_10462_),
    .A(_10431_),
    .Y(_10463_));
 sg13g2_buf_1 _17283_ (.A(_10463_),
    .X(_10464_));
 sg13g2_buf_1 _17284_ (.A(\cpu.dec.imm[3] ),
    .X(_10465_));
 sg13g2_nor2_1 _17285_ (.A(_10465_),
    .B(net1109),
    .Y(_10466_));
 sg13g2_inv_1 _17286_ (.Y(_10467_),
    .A(net1012));
 sg13g2_nor2_1 _17287_ (.A(_08265_),
    .B(_10467_),
    .Y(_10468_));
 sg13g2_a21oi_1 _17288_ (.A1(_10413_),
    .A2(_10466_),
    .Y(_10469_),
    .B1(_10468_));
 sg13g2_buf_1 _17289_ (.A(_10469_),
    .X(_10470_));
 sg13g2_nand2_1 _17290_ (.Y(_10471_),
    .A(net879),
    .B(net874));
 sg13g2_buf_1 _17291_ (.A(\cpu.ex.mmu_read[2] ),
    .X(_10472_));
 sg13g2_and2_1 _17292_ (.A(net881),
    .B(net1015),
    .X(_10473_));
 sg13g2_inv_1 _17293_ (.Y(_10474_),
    .A(_00258_));
 sg13g2_a22oi_1 _17294_ (.Y(_10475_),
    .B1(_10473_),
    .B2(_10474_),
    .A2(_10294_),
    .A1(_10472_));
 sg13g2_nor2_1 _17295_ (.A(_10471_),
    .B(_10475_),
    .Y(_10476_));
 sg13g2_nand2b_1 _17296_ (.Y(_10477_),
    .B(net1015),
    .A_N(_10273_));
 sg13g2_buf_2 _17297_ (.A(_10477_),
    .X(_10478_));
 sg13g2_a22oi_1 _17298_ (.Y(_10479_),
    .B1(_10357_),
    .B2(\cpu.ex.r_11[2] ),
    .A2(_10312_),
    .A1(\cpu.ex.r_8[2] ));
 sg13g2_nor2_1 _17299_ (.A(_10478_),
    .B(_10479_),
    .Y(_10480_));
 sg13g2_nand2_1 _17300_ (.Y(_10481_),
    .A(net881),
    .B(_10308_));
 sg13g2_buf_1 _17301_ (.A(\cpu.ex.r_sp[2] ),
    .X(_10482_));
 sg13g2_and2_1 _17302_ (.A(\cpu.ex.r_epc[2] ),
    .B(net1016),
    .X(_10483_));
 sg13g2_a21oi_1 _17303_ (.A1(_10482_),
    .A2(_10260_),
    .Y(_10484_),
    .B1(_10483_));
 sg13g2_nand3_1 _17304_ (.B(net880),
    .C(_10357_),
    .A(\cpu.ex.r_mult[18] ),
    .Y(_10485_));
 sg13g2_o21ai_1 _17305_ (.B1(_10485_),
    .Y(_10486_),
    .A1(_10481_),
    .A2(_10484_));
 sg13g2_mux2_1 _17306_ (.A0(\cpu.ex.r_10[2] ),
    .A1(\cpu.ex.r_14[2] ),
    .S(_10273_),
    .X(_10487_));
 sg13g2_nand3_1 _17307_ (.B(_10290_),
    .C(_10487_),
    .A(_10283_),
    .Y(_10488_));
 sg13g2_mux2_1 _17308_ (.A0(\cpu.ex.r_lr[2] ),
    .A1(\cpu.ex.r_9[2] ),
    .S(net1015),
    .X(_10489_));
 sg13g2_nand3_1 _17309_ (.B(net751),
    .C(_10489_),
    .A(net752),
    .Y(_10490_));
 sg13g2_mux2_1 _17310_ (.A0(net1127),
    .A1(\cpu.ex.r_stmp[2] ),
    .S(net1017),
    .X(_10491_));
 sg13g2_nand3_1 _17311_ (.B(_10452_),
    .C(_10491_),
    .A(net878),
    .Y(_10492_));
 sg13g2_mux2_1 _17312_ (.A0(\cpu.ex.r_12[2] ),
    .A1(\cpu.ex.r_13[2] ),
    .S(net1016),
    .X(_10493_));
 sg13g2_nand3_1 _17313_ (.B(net753),
    .C(_10493_),
    .A(net874),
    .Y(_10494_));
 sg13g2_nand4_1 _17314_ (.B(_10490_),
    .C(_10492_),
    .A(_10488_),
    .Y(_10495_),
    .D(_10494_));
 sg13g2_or4_1 _17315_ (.A(_10476_),
    .B(_10480_),
    .C(_10486_),
    .D(_10495_),
    .X(_10496_));
 sg13g2_nand2_1 _17316_ (.Y(_10497_),
    .A(net1109),
    .B(_10413_));
 sg13g2_a221oi_1 _17317_ (.B2(_10496_),
    .C1(_10497_),
    .B1(_10336_),
    .A1(_09268_),
    .Y(_10498_),
    .A2(net613));
 sg13g2_buf_1 _17318_ (.A(_10498_),
    .X(_10499_));
 sg13g2_buf_1 _17319_ (.A(\cpu.dec.imm[2] ),
    .X(_10500_));
 sg13g2_nor3_1 _17320_ (.A(_10500_),
    .B(net1109),
    .C(_10324_),
    .Y(_10501_));
 sg13g2_a21o_1 _17321_ (.A2(_10321_),
    .A1(_08278_),
    .B1(_10501_),
    .X(_10502_));
 sg13g2_buf_1 _17322_ (.A(_10502_),
    .X(_10503_));
 sg13g2_nor2_1 _17323_ (.A(_10499_),
    .B(_10503_),
    .Y(_10504_));
 sg13g2_buf_2 _17324_ (.A(_10504_),
    .X(_10505_));
 sg13g2_a21oi_1 _17325_ (.A1(_10464_),
    .A2(_10470_),
    .Y(_10506_),
    .B1(_10505_));
 sg13g2_buf_2 _17326_ (.A(_10506_),
    .X(_10507_));
 sg13g2_buf_1 _17327_ (.A(_00305_),
    .X(_10508_));
 sg13g2_and3_1 _17328_ (.X(_10509_),
    .A(_10431_),
    .B(_10461_),
    .C(_10462_));
 sg13g2_buf_2 _17329_ (.A(_10509_),
    .X(_10510_));
 sg13g2_a21o_1 _17330_ (.A2(_10466_),
    .A1(_10413_),
    .B1(_10468_),
    .X(_10511_));
 sg13g2_buf_2 _17331_ (.A(_10511_),
    .X(_10512_));
 sg13g2_nor2_2 _17332_ (.A(_10510_),
    .B(_10512_),
    .Y(_10513_));
 sg13g2_buf_1 _17333_ (.A(_00306_),
    .X(_10514_));
 sg13g2_a21oi_1 _17334_ (.A1(net1105),
    .A2(_10513_),
    .Y(_10515_),
    .B1(_10514_));
 sg13g2_nand2_1 _17335_ (.Y(_10516_),
    .A(net749),
    .B(_10515_));
 sg13g2_inv_1 _17336_ (.Y(_10517_),
    .A(_10516_));
 sg13g2_buf_1 _17337_ (.A(_00307_),
    .X(_10518_));
 sg13g2_nor2_1 _17338_ (.A(_10518_),
    .B(_09370_),
    .Y(_10519_));
 sg13g2_buf_1 _17339_ (.A(\cpu.dec.imm[1] ),
    .X(_10520_));
 sg13g2_inv_1 _17340_ (.Y(_10521_),
    .A(_10520_));
 sg13g2_nand2_1 _17341_ (.Y(_10522_),
    .A(_09271_),
    .B(net613));
 sg13g2_mux2_1 _17342_ (.A0(_10521_),
    .A1(_10522_),
    .S(net1109),
    .X(_10523_));
 sg13g2_inv_1 _17343_ (.Y(_10524_),
    .A(\cpu.ex.r_mult[17] ));
 sg13g2_mux2_1 _17344_ (.A0(_00257_),
    .A1(_10524_),
    .S(_10355_),
    .X(_10525_));
 sg13g2_buf_1 _17345_ (.A(\cpu.ex.r_prev_ie ),
    .X(_10526_));
 sg13g2_mux2_1 _17346_ (.A0(_10526_),
    .A1(\cpu.ex.mmu_read[1] ),
    .S(_10243_),
    .X(_10527_));
 sg13g2_nand3_1 _17347_ (.B(_10294_),
    .C(_10527_),
    .A(net874),
    .Y(_10528_));
 sg13g2_o21ai_1 _17348_ (.B1(_10528_),
    .Y(_10529_),
    .A1(_10275_),
    .A2(_10525_));
 sg13g2_and3_1 _17349_ (.X(_10530_),
    .A(\cpu.ex.r_11[1] ),
    .B(_10265_),
    .C(_10357_));
 sg13g2_nand2_1 _17350_ (.Y(_10531_),
    .A(net874),
    .B(_10344_));
 sg13g2_and2_1 _17351_ (.A(\cpu.ex.r_13[1] ),
    .B(_10243_),
    .X(_10532_));
 sg13g2_a21oi_1 _17352_ (.A1(\cpu.ex.r_12[1] ),
    .A2(_10260_),
    .Y(_10533_),
    .B1(_10532_));
 sg13g2_mux2_1 _17353_ (.A0(\cpu.ex.r_stmp[1] ),
    .A1(\cpu.ex.r_14[1] ),
    .S(net1015),
    .X(_10534_));
 sg13g2_nand3_1 _17354_ (.B(_10290_),
    .C(_10534_),
    .A(net874),
    .Y(_10535_));
 sg13g2_o21ai_1 _17355_ (.B1(_10535_),
    .Y(_10536_),
    .A1(_10531_),
    .A2(_10533_));
 sg13g2_nor3_1 _17356_ (.A(_10529_),
    .B(_10530_),
    .C(_10536_),
    .Y(_10537_));
 sg13g2_a22oi_1 _17357_ (.Y(_10538_),
    .B1(_10344_),
    .B2(\cpu.ex.r_9[1] ),
    .A2(_10348_),
    .A1(\cpu.ex.r_epc[1] ));
 sg13g2_buf_1 _17358_ (.A(\cpu.ex.r_sp[1] ),
    .X(_10539_));
 sg13g2_a221oi_1 _17359_ (.B2(\cpu.ex.r_8[1] ),
    .C1(net1016),
    .B1(_10344_),
    .A1(_10539_),
    .Y(_10540_),
    .A2(_10348_));
 sg13g2_a21oi_1 _17360_ (.A1(net879),
    .A2(_10538_),
    .Y(_10541_),
    .B1(_10540_));
 sg13g2_nand3_1 _17361_ (.B(net877),
    .C(_10290_),
    .A(\cpu.ex.r_10[1] ),
    .Y(_10542_));
 sg13g2_nand3_1 _17362_ (.B(net1016),
    .C(_10294_),
    .A(\cpu.ex.r_lr[1] ),
    .Y(_10543_));
 sg13g2_nand2_1 _17363_ (.Y(_10544_),
    .A(_10542_),
    .B(_10543_));
 sg13g2_o21ai_1 _17364_ (.B1(net752),
    .Y(_10545_),
    .A1(_10541_),
    .A2(_10544_));
 sg13g2_nand2_1 _17365_ (.Y(_10546_),
    .A(net1109),
    .B(_10335_));
 sg13g2_a21o_1 _17366_ (.A2(_10545_),
    .A1(_10537_),
    .B1(_10546_),
    .X(_10547_));
 sg13g2_nand3_1 _17367_ (.B(_10523_),
    .C(_10547_),
    .A(_10413_),
    .Y(_10548_));
 sg13g2_buf_1 _17368_ (.A(_10548_),
    .X(_10549_));
 sg13g2_nand2_1 _17369_ (.Y(_10550_),
    .A(_08389_),
    .B(_10321_));
 sg13g2_nand2_1 _17370_ (.Y(_10551_),
    .A(_10549_),
    .B(_10550_));
 sg13g2_buf_2 _17371_ (.A(_10551_),
    .X(_10552_));
 sg13g2_nor2_1 _17372_ (.A(_10519_),
    .B(_10552_),
    .Y(_10553_));
 sg13g2_xor2_1 _17373_ (.B(_09374_),
    .A(_09362_),
    .X(_10554_));
 sg13g2_and3_1 _17374_ (.X(_10555_),
    .A(net693),
    .B(net749),
    .C(_10554_));
 sg13g2_buf_8 _17375_ (.A(_10555_),
    .X(_10556_));
 sg13g2_buf_1 _17376_ (.A(_10556_),
    .X(_10557_));
 sg13g2_nor3_1 _17377_ (.A(_09362_),
    .B(_09374_),
    .C(_09375_),
    .Y(_10558_));
 sg13g2_xnor2_1 _17378_ (.Y(_10559_),
    .A(_09376_),
    .B(_10558_));
 sg13g2_and3_1 _17379_ (.X(_10560_),
    .A(_09385_),
    .B(net749),
    .C(_10559_));
 sg13g2_buf_1 _17380_ (.A(_10560_),
    .X(_10561_));
 sg13g2_inv_2 _17381_ (.Y(\cpu.ex.c_mult_off[3] ),
    .A(net609));
 sg13g2_buf_2 _17382_ (.A(\cpu.dec.r_rs1[3] ),
    .X(_10562_));
 sg13g2_buf_8 _17383_ (.A(\cpu.dec.r_rs1[2] ),
    .X(_10563_));
 sg13g2_nor2_1 _17384_ (.A(_10562_),
    .B(_10563_),
    .Y(_10564_));
 sg13g2_buf_1 _17385_ (.A(_10564_),
    .X(_10565_));
 sg13g2_buf_2 _17386_ (.A(\cpu.dec.r_rs1[0] ),
    .X(_10566_));
 sg13g2_buf_8 _17387_ (.A(\cpu.dec.r_rs1[1] ),
    .X(_10567_));
 sg13g2_nor2_1 _17388_ (.A(_10566_),
    .B(_10567_),
    .Y(_10568_));
 sg13g2_buf_2 _17389_ (.A(_10568_),
    .X(_10569_));
 sg13g2_a21oi_1 _17390_ (.A1(net872),
    .A2(_10569_),
    .Y(_10570_),
    .B1(_00271_));
 sg13g2_nand2_1 _17391_ (.Y(_10571_),
    .A(_09214_),
    .B(_09257_));
 sg13g2_a21o_1 _17392_ (.A2(_09243_),
    .A1(_09224_),
    .B1(_10571_),
    .X(_10572_));
 sg13g2_a21oi_1 _17393_ (.A1(_09257_),
    .A2(_09255_),
    .Y(_10573_),
    .B1(_09212_));
 sg13g2_nand3_1 _17394_ (.B(_10572_),
    .C(_10573_),
    .A(_10570_),
    .Y(_10574_));
 sg13g2_buf_1 _17395_ (.A(_10574_),
    .X(_10575_));
 sg13g2_nand3b_1 _17396_ (.B(_08537_),
    .C(_08613_),
    .Y(_10576_),
    .A_N(_10575_));
 sg13g2_buf_8 _17397_ (.A(_10576_),
    .X(_10577_));
 sg13g2_buf_1 _17398_ (.A(\cpu.br ),
    .X(_10578_));
 sg13g2_inv_2 _17399_ (.Y(_10579_),
    .A(_10578_));
 sg13g2_nor2_1 _17400_ (.A(_10579_),
    .B(_00295_),
    .Y(_10580_));
 sg13g2_and4_1 _17401_ (.A(_08469_),
    .B(_08515_),
    .C(_08525_),
    .D(_08535_),
    .X(_10581_));
 sg13g2_buf_2 _17402_ (.A(_10581_),
    .X(_10582_));
 sg13g2_buf_8 _17403_ (.A(_10566_),
    .X(_10583_));
 sg13g2_buf_8 _17404_ (.A(_10583_),
    .X(_10584_));
 sg13g2_buf_8 _17405_ (.A(net871),
    .X(_10585_));
 sg13g2_buf_1 _17406_ (.A(net748),
    .X(_10586_));
 sg13g2_buf_8 _17407_ (.A(_10562_),
    .X(_10587_));
 sg13g2_buf_8 _17408_ (.A(_10563_),
    .X(_10588_));
 sg13g2_nor2b_1 _17409_ (.A(net1009),
    .B_N(net1008),
    .Y(_10589_));
 sg13g2_buf_2 _17410_ (.A(_10589_),
    .X(_10590_));
 sg13g2_nor2b_1 _17411_ (.A(net1008),
    .B_N(_10562_),
    .Y(_10591_));
 sg13g2_buf_2 _17412_ (.A(_10591_),
    .X(_10592_));
 sg13g2_a22oi_1 _17413_ (.Y(_10593_),
    .B1(_10592_),
    .B2(\cpu.ex.r_10[2] ),
    .A2(_10590_),
    .A1(\cpu.ex.r_stmp[2] ));
 sg13g2_a22oi_1 _17414_ (.Y(_10594_),
    .B1(_10592_),
    .B2(\cpu.ex.r_8[2] ),
    .A2(_10590_),
    .A1(net1127));
 sg13g2_buf_8 _17415_ (.A(_10567_),
    .X(_10595_));
 sg13g2_inv_2 _17416_ (.Y(_10596_),
    .A(net1007));
 sg13g2_buf_1 _17417_ (.A(_10596_),
    .X(_10597_));
 sg13g2_mux2_1 _17418_ (.A0(_10593_),
    .A1(_10594_),
    .S(net747),
    .X(_10598_));
 sg13g2_nor2_1 _17419_ (.A(net665),
    .B(_10598_),
    .Y(_10599_));
 sg13g2_buf_1 _17420_ (.A(_10595_),
    .X(_10600_));
 sg13g2_buf_8 _17421_ (.A(net870),
    .X(_10601_));
 sg13g2_buf_8 _17422_ (.A(net1008),
    .X(_10602_));
 sg13g2_buf_1 _17423_ (.A(net869),
    .X(_10603_));
 sg13g2_nand2_1 _17424_ (.Y(_10604_),
    .A(net746),
    .B(net745));
 sg13g2_nor2b_1 _17425_ (.A(net1010),
    .B_N(_10562_),
    .Y(_10605_));
 sg13g2_buf_2 _17426_ (.A(_10605_),
    .X(_10606_));
 sg13g2_buf_8 _17427_ (.A(_10562_),
    .X(_10607_));
 sg13g2_inv_2 _17428_ (.Y(_10608_),
    .A(net1006));
 sg13g2_mux2_1 _17429_ (.A0(_10474_),
    .A1(\cpu.ex.r_mult[18] ),
    .S(_10608_),
    .X(_10609_));
 sg13g2_a22oi_1 _17430_ (.Y(_10610_),
    .B1(_10609_),
    .B2(net665),
    .A2(_10606_),
    .A1(\cpu.ex.r_14[2] ));
 sg13g2_nor2_1 _17431_ (.A(_10604_),
    .B(_10610_),
    .Y(_10611_));
 sg13g2_buf_8 _17432_ (.A(net1007),
    .X(_10612_));
 sg13g2_buf_8 _17433_ (.A(net868),
    .X(_10613_));
 sg13g2_buf_8 _17434_ (.A(_10607_),
    .X(_10614_));
 sg13g2_nor2_1 _17435_ (.A(net744),
    .B(net867),
    .Y(_10615_));
 sg13g2_and2_1 _17436_ (.A(net868),
    .B(net1009),
    .X(_10616_));
 sg13g2_buf_1 _17437_ (.A(_10616_),
    .X(_10617_));
 sg13g2_a22oi_1 _17438_ (.Y(_10618_),
    .B1(_10617_),
    .B2(\cpu.ex.r_11[2] ),
    .A2(_10615_),
    .A1(\cpu.ex.r_lr[2] ));
 sg13g2_inv_1 _17439_ (.Y(_10619_),
    .A(net1010));
 sg13g2_buf_1 _17440_ (.A(_10619_),
    .X(_10620_));
 sg13g2_buf_1 _17441_ (.A(_10563_),
    .X(_10621_));
 sg13g2_buf_1 _17442_ (.A(net1005),
    .X(_10622_));
 sg13g2_nor2_1 _17443_ (.A(net743),
    .B(net866),
    .Y(_10623_));
 sg13g2_nand2b_1 _17444_ (.Y(_10624_),
    .B(_10623_),
    .A_N(_10618_));
 sg13g2_and2_1 _17445_ (.A(net1010),
    .B(_10567_),
    .X(_10625_));
 sg13g2_buf_2 _17446_ (.A(_10625_),
    .X(_10626_));
 sg13g2_and2_1 _17447_ (.A(net872),
    .B(_10626_),
    .X(_10627_));
 sg13g2_buf_1 _17448_ (.A(_10627_),
    .X(_10628_));
 sg13g2_nand2_1 _17449_ (.Y(_10629_),
    .A(\cpu.ex.r_epc[2] ),
    .B(_10628_));
 sg13g2_buf_8 _17450_ (.A(net869),
    .X(_10630_));
 sg13g2_buf_1 _17451_ (.A(net742),
    .X(_10631_));
 sg13g2_nor2b_1 _17452_ (.A(_10567_),
    .B_N(net1010),
    .Y(_10632_));
 sg13g2_buf_2 _17453_ (.A(_10632_),
    .X(_10633_));
 sg13g2_buf_1 _17454_ (.A(_10633_),
    .X(_10634_));
 sg13g2_buf_1 _17455_ (.A(_10607_),
    .X(_10635_));
 sg13g2_inv_1 _17456_ (.Y(_10636_),
    .A(_10472_));
 sg13g2_buf_1 _17457_ (.A(_10636_),
    .X(_10637_));
 sg13g2_nand2_1 _17458_ (.Y(_10638_),
    .A(_10614_),
    .B(\cpu.ex.r_13[2] ));
 sg13g2_o21ai_1 _17459_ (.B1(_10638_),
    .Y(_10639_),
    .A1(_10635_),
    .A2(_10637_));
 sg13g2_nand3_1 _17460_ (.B(net663),
    .C(_10639_),
    .A(_10631_),
    .Y(_10640_));
 sg13g2_nand3_1 _17461_ (.B(_10629_),
    .C(_10640_),
    .A(_10624_),
    .Y(_10641_));
 sg13g2_xor2_1 _17462_ (.B(_10563_),
    .A(net1110),
    .X(_10642_));
 sg13g2_xor2_1 _17463_ (.B(_10567_),
    .A(net1019),
    .X(_10643_));
 sg13g2_xor2_1 _17464_ (.B(_10562_),
    .A(net1111),
    .X(_10644_));
 sg13g2_xor2_1 _17465_ (.B(_10566_),
    .A(net1018),
    .X(_10645_));
 sg13g2_nor4_2 _17466_ (.A(_10642_),
    .B(_10643_),
    .C(_10644_),
    .Y(_10646_),
    .D(_10645_));
 sg13g2_nand2_1 _17467_ (.Y(_10647_),
    .A(_10332_),
    .B(_10646_));
 sg13g2_buf_1 _17468_ (.A(_10647_),
    .X(_10648_));
 sg13g2_nand3_1 _17469_ (.B(\cpu.ex.r_9[2] ),
    .C(_10633_),
    .A(net865),
    .Y(_10649_));
 sg13g2_nor2b_1 _17470_ (.A(_10583_),
    .B_N(_10595_),
    .Y(_10650_));
 sg13g2_buf_1 _17471_ (.A(_10650_),
    .X(_10651_));
 sg13g2_nand3_1 _17472_ (.B(_10482_),
    .C(_10651_),
    .A(_10608_),
    .Y(_10652_));
 sg13g2_a21o_1 _17473_ (.A2(_10652_),
    .A1(_10649_),
    .B1(net664),
    .X(_10653_));
 sg13g2_and2_1 _17474_ (.A(net1009),
    .B(_10569_),
    .X(_10654_));
 sg13g2_buf_1 _17475_ (.A(_10654_),
    .X(_10655_));
 sg13g2_nand3_1 _17476_ (.B(\cpu.ex.r_12[2] ),
    .C(_10655_),
    .A(net664),
    .Y(_10656_));
 sg13g2_nand3_1 _17477_ (.B(_10653_),
    .C(_10656_),
    .A(net608),
    .Y(_10657_));
 sg13g2_nor4_2 _17478_ (.A(_10599_),
    .B(_10611_),
    .C(_10641_),
    .Y(_10658_),
    .D(_10657_));
 sg13g2_buf_8 _17479_ (.A(net608),
    .X(_10659_));
 sg13g2_nor2_1 _17480_ (.A(_09268_),
    .B(net532),
    .Y(_10660_));
 sg13g2_nor4_1 _17481_ (.A(_10582_),
    .B(_10575_),
    .C(_10658_),
    .D(_10660_),
    .Y(_10661_));
 sg13g2_buf_1 _17482_ (.A(_10578_),
    .X(_10662_));
 sg13g2_nor3_1 _17483_ (.A(net1004),
    .B(_10658_),
    .C(_10660_),
    .Y(_10663_));
 sg13g2_a221oi_1 _17484_ (.B2(_08613_),
    .C1(_10663_),
    .B1(_10661_),
    .A1(_10577_),
    .Y(_10664_),
    .A2(_10580_));
 sg13g2_buf_8 _17485_ (.A(_10664_),
    .X(_10665_));
 sg13g2_nor3_1 _17486_ (.A(net471),
    .B(\cpu.ex.c_mult_off[3] ),
    .C(_10665_),
    .Y(_10666_));
 sg13g2_inv_1 _17487_ (.Y(_10667_),
    .A(_10563_));
 sg13g2_buf_2 _17488_ (.A(_10667_),
    .X(_10668_));
 sg13g2_buf_1 _17489_ (.A(_10668_),
    .X(_10669_));
 sg13g2_and2_1 _17490_ (.A(net1010),
    .B(_10562_),
    .X(_10670_));
 sg13g2_buf_1 _17491_ (.A(_10670_),
    .X(_10671_));
 sg13g2_nand3_1 _17492_ (.B(\cpu.ex.r_11[8] ),
    .C(_10671_),
    .A(net741),
    .Y(_10672_));
 sg13g2_nand3_1 _17493_ (.B(\cpu.ex.r_stmp[8] ),
    .C(_10590_),
    .A(net743),
    .Y(_10673_));
 sg13g2_a21oi_1 _17494_ (.A1(_10672_),
    .A2(_10673_),
    .Y(_10674_),
    .B1(_10597_));
 sg13g2_nor2b_1 _17495_ (.A(_00264_),
    .B_N(_10613_),
    .Y(_10675_));
 sg13g2_nor2b_1 _17496_ (.A(_10601_),
    .B_N(\cpu.ex.r_13[8] ),
    .Y(_10676_));
 sg13g2_and3_1 _17497_ (.X(_10677_),
    .A(net871),
    .B(net1009),
    .C(_10621_));
 sg13g2_buf_1 _17498_ (.A(_10677_),
    .X(_10678_));
 sg13g2_o21ai_1 _17499_ (.B1(_10678_),
    .Y(_10679_),
    .A1(_10675_),
    .A2(_10676_));
 sg13g2_nor2b_1 _17500_ (.A(net1006),
    .B_N(net868),
    .Y(_10680_));
 sg13g2_buf_2 _17501_ (.A(_10680_),
    .X(_10681_));
 sg13g2_buf_1 _17502_ (.A(\cpu.ex.r_sp[8] ),
    .X(_10682_));
 sg13g2_buf_1 _17503_ (.A(net871),
    .X(_10683_));
 sg13g2_mux2_1 _17504_ (.A0(_10682_),
    .A1(\cpu.ex.r_epc[8] ),
    .S(net740),
    .X(_10684_));
 sg13g2_nand3_1 _17505_ (.B(_10681_),
    .C(_10684_),
    .A(net741),
    .Y(_10685_));
 sg13g2_buf_1 _17506_ (.A(_10651_),
    .X(_10686_));
 sg13g2_nand3_1 _17507_ (.B(_10686_),
    .C(_10592_),
    .A(\cpu.ex.r_10[8] ),
    .Y(_10687_));
 sg13g2_buf_8 _17508_ (.A(net1009),
    .X(_10688_));
 sg13g2_mux2_1 _17509_ (.A0(\cpu.ex.r_lr[8] ),
    .A1(\cpu.ex.r_9[8] ),
    .S(net863),
    .X(_10689_));
 sg13g2_nand3_1 _17510_ (.B(_10634_),
    .C(_10689_),
    .A(net741),
    .Y(_10690_));
 sg13g2_nand4_1 _17511_ (.B(_10685_),
    .C(_10687_),
    .A(_10679_),
    .Y(_10691_),
    .D(_10690_));
 sg13g2_nor2b_1 _17512_ (.A(_10562_),
    .B_N(net1010),
    .Y(_10692_));
 sg13g2_buf_2 _17513_ (.A(_10692_),
    .X(_10693_));
 sg13g2_a22oi_1 _17514_ (.Y(_10694_),
    .B1(_10693_),
    .B2(\cpu.ex.r_mult[24] ),
    .A2(_10606_),
    .A1(\cpu.ex.r_14[8] ));
 sg13g2_buf_1 _17515_ (.A(net867),
    .X(_10695_));
 sg13g2_mux2_1 _17516_ (.A0(\cpu.ex.r_8[8] ),
    .A1(\cpu.ex.r_12[8] ),
    .S(net866),
    .X(_10696_));
 sg13g2_nand3_1 _17517_ (.B(_10569_),
    .C(_10696_),
    .A(_10695_),
    .Y(_10697_));
 sg13g2_o21ai_1 _17518_ (.B1(_10697_),
    .Y(_10698_),
    .A1(_10604_),
    .A2(_10694_));
 sg13g2_nor3_1 _17519_ (.A(_10674_),
    .B(_10691_),
    .C(_10698_),
    .Y(_10699_));
 sg13g2_nor2_1 _17520_ (.A(_09202_),
    .B(net608),
    .Y(_10700_));
 sg13g2_a21oi_2 _17521_ (.B1(_10700_),
    .Y(_10701_),
    .A2(_10699_),
    .A1(net532));
 sg13g2_nand2_1 _17522_ (.Y(_10702_),
    .A(_10557_),
    .B(_10701_));
 sg13g2_inv_1 _17523_ (.Y(\cpu.ex.c_mult_off[1] ),
    .A(_10557_));
 sg13g2_buf_1 _17524_ (.A(\cpu.addr[10] ),
    .X(_10703_));
 sg13g2_nor2b_1 _17525_ (.A(net868),
    .B_N(net1005),
    .Y(_10704_));
 sg13g2_mux2_1 _17526_ (.A0(\cpu.ex.r_12[10] ),
    .A1(\cpu.ex.r_13[10] ),
    .S(net740),
    .X(_10705_));
 sg13g2_nor2b_1 _17527_ (.A(net1005),
    .B_N(net1007),
    .Y(_10706_));
 sg13g2_mux2_1 _17528_ (.A0(\cpu.ex.r_10[10] ),
    .A1(\cpu.ex.r_11[10] ),
    .S(net748),
    .X(_10707_));
 sg13g2_a22oi_1 _17529_ (.Y(_10708_),
    .B1(_10706_),
    .B2(_10707_),
    .A2(_10705_),
    .A1(_10704_));
 sg13g2_nand2b_1 _17530_ (.Y(_10709_),
    .B(net739),
    .A_N(_10708_));
 sg13g2_nand2b_1 _17531_ (.Y(_10710_),
    .B(net1007),
    .A_N(net1010));
 sg13g2_buf_2 _17532_ (.A(_10710_),
    .X(_10711_));
 sg13g2_nor2_1 _17533_ (.A(net741),
    .B(_10711_),
    .Y(_10712_));
 sg13g2_mux2_1 _17534_ (.A0(\cpu.ex.r_stmp[10] ),
    .A1(\cpu.ex.r_14[10] ),
    .S(net865),
    .X(_10713_));
 sg13g2_buf_8 _17535_ (.A(_10612_),
    .X(_10714_));
 sg13g2_nand3b_1 _17536_ (.B(net865),
    .C(\cpu.ex.r_8[10] ),
    .Y(_10715_),
    .A_N(net738));
 sg13g2_buf_1 _17537_ (.A(\cpu.ex.r_sp[10] ),
    .X(_10716_));
 sg13g2_nand3b_1 _17538_ (.B(_10716_),
    .C(net738),
    .Y(_10717_),
    .A_N(net867));
 sg13g2_or2_1 _17539_ (.X(_10718_),
    .B(_10588_),
    .A(net1010));
 sg13g2_buf_1 _17540_ (.A(_10718_),
    .X(_10719_));
 sg13g2_a21oi_1 _17541_ (.A1(_10715_),
    .A2(_10717_),
    .Y(_10720_),
    .B1(_10719_));
 sg13g2_a221oi_1 _17542_ (.B2(_10713_),
    .C1(_10720_),
    .B1(_10712_),
    .A1(\cpu.ex.r_epc[10] ),
    .Y(_10721_),
    .A2(_10628_));
 sg13g2_nor2_1 _17543_ (.A(net868),
    .B(_10602_),
    .Y(_10722_));
 sg13g2_and2_1 _17544_ (.A(net1007),
    .B(net1008),
    .X(_10723_));
 sg13g2_buf_1 _17545_ (.A(_10723_),
    .X(_10724_));
 sg13g2_a221oi_1 _17546_ (.B2(net1106),
    .C1(net865),
    .B1(_10724_),
    .A1(\cpu.ex.r_lr[10] ),
    .Y(_10725_),
    .A2(_10722_));
 sg13g2_inv_1 _17547_ (.Y(_10726_),
    .A(_00266_));
 sg13g2_a221oi_1 _17548_ (.B2(_10726_),
    .C1(_10608_),
    .B1(_10724_),
    .A1(\cpu.ex.r_9[10] ),
    .Y(_10727_),
    .A2(_10722_));
 sg13g2_or3_1 _17549_ (.A(net743),
    .B(_10725_),
    .C(_10727_),
    .X(_10728_));
 sg13g2_nand3_1 _17550_ (.B(_10721_),
    .C(_10728_),
    .A(_10709_),
    .Y(_10729_));
 sg13g2_mux2_1 _17551_ (.A0(net1104),
    .A1(_10729_),
    .S(net608),
    .X(_10730_));
 sg13g2_nand2_1 _17552_ (.Y(_10731_),
    .A(\cpu.ex.c_mult_off[1] ),
    .B(_10730_));
 sg13g2_a221oi_1 _17553_ (.B2(_10731_),
    .C1(_10561_),
    .B1(_10702_),
    .A1(net1004),
    .Y(_10732_),
    .A2(_10577_));
 sg13g2_a21o_1 _17554_ (.A2(_08577_),
    .A1(_08574_),
    .B1(_08612_),
    .X(_10733_));
 sg13g2_buf_1 _17555_ (.A(_10733_),
    .X(_10734_));
 sg13g2_nor3_1 _17556_ (.A(_10582_),
    .B(_10734_),
    .C(_10575_),
    .Y(_10735_));
 sg13g2_buf_8 _17557_ (.A(_10735_),
    .X(_10736_));
 sg13g2_inv_1 _17558_ (.Y(_10737_),
    .A(_00291_));
 sg13g2_buf_1 _17559_ (.A(_00289_),
    .X(_10738_));
 sg13g2_nor2_1 _17560_ (.A(_10738_),
    .B(net471),
    .Y(_10739_));
 sg13g2_a21oi_1 _17561_ (.A1(_10737_),
    .A2(net471),
    .Y(_10740_),
    .B1(_10739_));
 sg13g2_nor4_1 _17562_ (.A(_10579_),
    .B(_10736_),
    .C(net609),
    .D(_10740_),
    .Y(_10741_));
 sg13g2_nand2_1 _17563_ (.Y(_10742_),
    .A(_10556_),
    .B(net609));
 sg13g2_nand2_1 _17564_ (.Y(_10743_),
    .A(_10572_),
    .B(_10573_));
 sg13g2_nor2_1 _17565_ (.A(_08476_),
    .B(_10579_),
    .Y(_10744_));
 sg13g2_and2_1 _17566_ (.A(_10743_),
    .B(_10744_),
    .X(_10745_));
 sg13g2_and2_1 _17567_ (.A(_10332_),
    .B(_10646_),
    .X(_10746_));
 sg13g2_buf_8 _17568_ (.A(_10746_),
    .X(_10747_));
 sg13g2_buf_8 _17569_ (.A(_10747_),
    .X(_10748_));
 sg13g2_inv_1 _17570_ (.Y(_10749_),
    .A(net1126));
 sg13g2_mux2_1 _17571_ (.A0(\cpu.ex.r_12[0] ),
    .A1(\cpu.ex.r_14[0] ),
    .S(net1007),
    .X(_10750_));
 sg13g2_nand2_1 _17572_ (.Y(_10751_),
    .A(net866),
    .B(_10750_));
 sg13g2_nand3_1 _17573_ (.B(_10668_),
    .C(\cpu.ex.r_8[0] ),
    .A(_10596_),
    .Y(_10752_));
 sg13g2_nand2b_1 _17574_ (.Y(_10753_),
    .B(net1006),
    .A_N(net871));
 sg13g2_a21oi_1 _17575_ (.A1(_10751_),
    .A2(_10752_),
    .Y(_10754_),
    .B1(_10753_));
 sg13g2_mux2_1 _17576_ (.A0(\cpu.ex.r_11[0] ),
    .A1(\cpu.ex.r_15[0] ),
    .S(_10563_),
    .X(_10755_));
 sg13g2_nor2b_1 _17577_ (.A(net1005),
    .B_N(\cpu.ex.r_9[0] ),
    .Y(_10756_));
 sg13g2_mux2_1 _17578_ (.A0(_10755_),
    .A1(_10756_),
    .S(_10596_),
    .X(_10757_));
 sg13g2_nand3b_1 _17579_ (.B(net1005),
    .C(\cpu.ex.r_stmp[0] ),
    .Y(_10758_),
    .A_N(_10587_));
 sg13g2_nand3b_1 _17580_ (.B(\cpu.ex.r_10[0] ),
    .C(_10587_),
    .Y(_10759_),
    .A_N(net1005));
 sg13g2_a21oi_1 _17581_ (.A1(_10758_),
    .A2(_10759_),
    .Y(_10760_),
    .B1(_10711_));
 sg13g2_a21o_1 _17582_ (.A2(_10757_),
    .A1(_10671_),
    .B1(_10760_),
    .X(_10761_));
 sg13g2_buf_1 _17583_ (.A(\cpu.ex.genblk3.r_prev_supmode ),
    .X(_10762_));
 sg13g2_and2_1 _17584_ (.A(_10762_),
    .B(net871),
    .X(_10763_));
 sg13g2_nor2b_1 _17585_ (.A(net871),
    .B_N(_09257_),
    .Y(_10764_));
 sg13g2_a22oi_1 _17586_ (.Y(_10765_),
    .B1(_10764_),
    .B2(_10704_),
    .A2(_10763_),
    .A1(_10706_));
 sg13g2_nand3b_1 _17587_ (.B(net1006),
    .C(\cpu.ex.r_13[0] ),
    .Y(_10766_),
    .A_N(net868));
 sg13g2_nand3b_1 _17588_ (.B(\cpu.ex.r_mult[16] ),
    .C(_10612_),
    .Y(_10767_),
    .A_N(net1009));
 sg13g2_nand2_1 _17589_ (.Y(_10768_),
    .A(net871),
    .B(_10621_));
 sg13g2_a21o_1 _17590_ (.A2(_10767_),
    .A1(_10766_),
    .B1(_10768_),
    .X(_10769_));
 sg13g2_o21ai_1 _17591_ (.B1(_10769_),
    .Y(_10770_),
    .A1(net865),
    .A2(_10765_));
 sg13g2_nor4_1 _17592_ (.A(_10747_),
    .B(_10754_),
    .C(_10761_),
    .D(_10770_),
    .Y(_10771_));
 sg13g2_a221oi_1 _17593_ (.B2(_10749_),
    .C1(_10771_),
    .B1(net531),
    .A1(net1004),
    .Y(_10772_),
    .A2(_10575_));
 sg13g2_nor4_2 _17594_ (.A(_10582_),
    .B(_10734_),
    .C(_10745_),
    .Y(_10773_),
    .D(_10772_));
 sg13g2_a21oi_1 _17595_ (.A1(_10749_),
    .A2(_10747_),
    .Y(_10774_),
    .B1(_10771_));
 sg13g2_a221oi_1 _17596_ (.B2(_10579_),
    .C1(_10744_),
    .B1(_10774_),
    .A1(_08537_),
    .Y(_10775_),
    .A2(_08613_));
 sg13g2_buf_1 _17597_ (.A(_10775_),
    .X(_10776_));
 sg13g2_nor3_1 _17598_ (.A(_10742_),
    .B(_10773_),
    .C(_10776_),
    .Y(_10777_));
 sg13g2_or4_1 _17599_ (.A(\cpu.ex.c_mult_off[0] ),
    .B(_10732_),
    .C(_10741_),
    .D(_10777_),
    .X(_10778_));
 sg13g2_buf_1 _17600_ (.A(_10778_),
    .X(_10779_));
 sg13g2_nand3_1 _17601_ (.B(\cpu.ex.r_stmp[6] ),
    .C(net662),
    .A(_10603_),
    .Y(_10780_));
 sg13g2_nand3_1 _17602_ (.B(\cpu.ex.r_lr[6] ),
    .C(_10633_),
    .A(net741),
    .Y(_10781_));
 sg13g2_a21o_1 _17603_ (.A2(_10781_),
    .A1(_10780_),
    .B1(net739),
    .X(_10782_));
 sg13g2_nand3_1 _17604_ (.B(\cpu.ex.r_8[6] ),
    .C(_10569_),
    .A(net865),
    .Y(_10783_));
 sg13g2_nand3_1 _17605_ (.B(\cpu.ex.r_epc[6] ),
    .C(_10626_),
    .A(_10608_),
    .Y(_10784_));
 sg13g2_a21o_1 _17606_ (.A2(_10784_),
    .A1(_10783_),
    .B1(net664),
    .X(_10785_));
 sg13g2_nor2_1 _17607_ (.A(_10668_),
    .B(_10753_),
    .Y(_10786_));
 sg13g2_mux2_1 _17608_ (.A0(\cpu.ex.r_12[6] ),
    .A1(\cpu.ex.r_14[6] ),
    .S(_10613_),
    .X(_10787_));
 sg13g2_buf_1 _17609_ (.A(\cpu.ex.r_sp[6] ),
    .X(_10788_));
 sg13g2_nor2_2 _17610_ (.A(_10584_),
    .B(net1009),
    .Y(_10789_));
 sg13g2_and3_1 _17611_ (.X(_10790_),
    .A(_10584_),
    .B(net1006),
    .C(\cpu.ex.r_11[6] ));
 sg13g2_a21o_1 _17612_ (.A2(_10789_),
    .A1(_10788_),
    .B1(_10790_),
    .X(_10791_));
 sg13g2_inv_1 _17613_ (.Y(_10792_),
    .A(\cpu.ex.r_10[6] ));
 sg13g2_nand2b_1 _17614_ (.Y(_10793_),
    .B(_10688_),
    .A_N(net869));
 sg13g2_nor3_1 _17615_ (.A(_10792_),
    .B(_10711_),
    .C(_10793_),
    .Y(_10794_));
 sg13g2_a221oi_1 _17616_ (.B2(_10706_),
    .C1(_10794_),
    .B1(_10791_),
    .A1(_10786_),
    .Y(_10795_),
    .A2(_10787_));
 sg13g2_inv_1 _17617_ (.Y(_10796_),
    .A(\cpu.ex.r_9[6] ));
 sg13g2_or2_1 _17618_ (.X(_10797_),
    .B(_10588_),
    .A(net1007));
 sg13g2_buf_1 _17619_ (.A(_10797_),
    .X(_10798_));
 sg13g2_nand3b_1 _17620_ (.B(net742),
    .C(net744),
    .Y(_10799_),
    .A_N(_00262_));
 sg13g2_o21ai_1 _17621_ (.B1(_10799_),
    .Y(_10800_),
    .A1(_10796_),
    .A2(_10798_));
 sg13g2_nand3b_1 _17622_ (.B(net867),
    .C(\cpu.ex.r_13[6] ),
    .Y(_10801_),
    .A_N(net744));
 sg13g2_buf_1 _17623_ (.A(\cpu.ex.r_mult[22] ),
    .X(_10802_));
 sg13g2_nand3b_1 _17624_ (.B(_10802_),
    .C(net744),
    .Y(_10803_),
    .A_N(_10614_));
 sg13g2_a21oi_1 _17625_ (.A1(_10801_),
    .A2(_10803_),
    .Y(_10804_),
    .B1(_10768_));
 sg13g2_a21oi_1 _17626_ (.A1(_10671_),
    .A2(_10800_),
    .Y(_10805_),
    .B1(_10804_));
 sg13g2_nand4_1 _17627_ (.B(_10785_),
    .C(_10795_),
    .A(_10782_),
    .Y(_10806_),
    .D(_10805_));
 sg13g2_nor4_1 _17628_ (.A(net471),
    .B(\cpu.ex.c_mult_off[3] ),
    .C(net531),
    .D(_10806_),
    .Y(_10807_));
 sg13g2_mux2_1 _17629_ (.A0(net922),
    .A1(_09206_),
    .S(net609),
    .X(_10808_));
 sg13g2_nor3_1 _17630_ (.A(net471),
    .B(net532),
    .C(_10808_),
    .Y(_10809_));
 sg13g2_and2_1 _17631_ (.A(_09374_),
    .B(_09376_),
    .X(_10810_));
 sg13g2_xnor2_1 _17632_ (.Y(_10811_),
    .A(_09375_),
    .B(_09376_));
 sg13g2_nor2_1 _17633_ (.A(_09362_),
    .B(_09374_),
    .Y(_10812_));
 sg13g2_a22oi_1 _17634_ (.Y(_10813_),
    .B1(_10811_),
    .B2(_10812_),
    .A2(_10810_),
    .A1(_09362_));
 sg13g2_nand2b_1 _17635_ (.Y(_10814_),
    .B(net1008),
    .A_N(net1007));
 sg13g2_buf_1 _17636_ (.A(\cpu.ex.mmu_read[14] ),
    .X(_10815_));
 sg13g2_a22oi_1 _17637_ (.Y(_10816_),
    .B1(_10693_),
    .B2(_10815_),
    .A2(_10606_),
    .A1(\cpu.ex.r_12[14] ));
 sg13g2_buf_1 _17638_ (.A(_10668_),
    .X(_10817_));
 sg13g2_mux2_1 _17639_ (.A0(\cpu.ex.r_8[14] ),
    .A1(\cpu.ex.r_10[14] ),
    .S(net744),
    .X(_10818_));
 sg13g2_nand3_1 _17640_ (.B(_10606_),
    .C(_10818_),
    .A(net737),
    .Y(_10819_));
 sg13g2_o21ai_1 _17641_ (.B1(_10819_),
    .Y(_10820_),
    .A1(_10814_),
    .A2(_10816_));
 sg13g2_a21oi_1 _17642_ (.A1(\cpu.ex.r_mult[30] ),
    .A2(_10590_),
    .Y(_10821_),
    .B1(net747));
 sg13g2_mux2_1 _17643_ (.A0(\cpu.ex.r_9[14] ),
    .A1(\cpu.ex.r_13[14] ),
    .S(net869),
    .X(_10822_));
 sg13g2_a221oi_1 _17644_ (.B2(net739),
    .C1(net746),
    .B1(_10822_),
    .A1(\cpu.ex.r_lr[14] ),
    .Y(_10823_),
    .A2(net872));
 sg13g2_nor3_1 _17645_ (.A(net743),
    .B(_10821_),
    .C(_10823_),
    .Y(_10824_));
 sg13g2_buf_1 _17646_ (.A(\cpu.ex.r_sp[14] ),
    .X(_10825_));
 sg13g2_mux2_1 _17647_ (.A0(\cpu.ex.r_epc[14] ),
    .A1(\cpu.ex.r_11[14] ),
    .S(net863),
    .X(_10826_));
 sg13g2_a221oi_1 _17648_ (.B2(net748),
    .C1(net664),
    .B1(_10826_),
    .A1(_10825_),
    .Y(_10827_),
    .A2(_10789_));
 sg13g2_inv_1 _17649_ (.Y(_10828_),
    .A(_00270_));
 sg13g2_mux2_1 _17650_ (.A0(\cpu.ex.r_stmp[14] ),
    .A1(\cpu.ex.r_14[14] ),
    .S(net863),
    .X(_10829_));
 sg13g2_a221oi_1 _17651_ (.B2(net743),
    .C1(net741),
    .B1(_10829_),
    .A1(_10828_),
    .Y(_10830_),
    .A2(_10671_));
 sg13g2_nor3_1 _17652_ (.A(net747),
    .B(_10827_),
    .C(_10830_),
    .Y(_10831_));
 sg13g2_or3_1 _17653_ (.A(_10820_),
    .B(_10824_),
    .C(_10831_),
    .X(_10832_));
 sg13g2_a221oi_1 _17654_ (.B2(_09371_),
    .C1(_10832_),
    .B1(_10813_),
    .A1(_10332_),
    .Y(_10833_),
    .A2(_10646_));
 sg13g2_nor4_1 _17655_ (.A(\cpu.ex.c_mult_off[0] ),
    .B(_10807_),
    .C(_10809_),
    .D(_10833_),
    .Y(_10834_));
 sg13g2_and2_1 _17656_ (.A(_09376_),
    .B(_10556_),
    .X(_10835_));
 sg13g2_mux2_1 _17657_ (.A0(\cpu.ex.r_8[12] ),
    .A1(\cpu.ex.r_12[12] ),
    .S(net869),
    .X(_10836_));
 sg13g2_mux2_1 _17658_ (.A0(\cpu.ex.r_lr[12] ),
    .A1(\cpu.ex.r_9[12] ),
    .S(net863),
    .X(_10837_));
 sg13g2_nor2_1 _17659_ (.A(net743),
    .B(_10798_),
    .Y(_10838_));
 sg13g2_a22oi_1 _17660_ (.Y(_10839_),
    .B1(_10837_),
    .B2(_10838_),
    .A2(_10836_),
    .A1(_10655_));
 sg13g2_a22oi_1 _17661_ (.Y(_10840_),
    .B1(_10693_),
    .B2(_10338_),
    .A2(_10606_),
    .A1(\cpu.ex.r_14[12] ));
 sg13g2_nand2b_1 _17662_ (.Y(_10841_),
    .B(_10724_),
    .A_N(_10840_));
 sg13g2_nor2_1 _17663_ (.A(net866),
    .B(_10711_),
    .Y(_10842_));
 sg13g2_and2_1 _17664_ (.A(net1006),
    .B(\cpu.ex.r_10[12] ),
    .X(_10843_));
 sg13g2_inv_1 _17665_ (.Y(_10844_),
    .A(_10371_));
 sg13g2_nand3b_1 _17666_ (.B(\cpu.ex.r_epc[12] ),
    .C(net868),
    .Y(_10845_),
    .A_N(net1005));
 sg13g2_o21ai_1 _17667_ (.B1(_10845_),
    .Y(_10846_),
    .A1(_10844_),
    .A2(_10814_));
 sg13g2_and4_1 _17668_ (.A(net863),
    .B(net869),
    .C(\cpu.ex.r_13[12] ),
    .D(_10633_),
    .X(_10847_));
 sg13g2_a221oi_1 _17669_ (.B2(_10693_),
    .C1(_10847_),
    .B1(_10846_),
    .A1(_10842_),
    .Y(_10848_),
    .A2(_10843_));
 sg13g2_nor2b_1 _17670_ (.A(_00268_),
    .B_N(net1008),
    .Y(_10849_));
 sg13g2_nor2b_1 _17671_ (.A(net1005),
    .B_N(\cpu.ex.r_11[12] ),
    .Y(_10850_));
 sg13g2_o21ai_1 _17672_ (.B1(_10671_),
    .Y(_10851_),
    .A1(_10849_),
    .A2(_10850_));
 sg13g2_mux2_1 _17673_ (.A0(_10373_),
    .A1(\cpu.ex.r_stmp[12] ),
    .S(net1008),
    .X(_10852_));
 sg13g2_nand2_1 _17674_ (.Y(_10853_),
    .A(_10789_),
    .B(_10852_));
 sg13g2_a21o_1 _17675_ (.A2(_10853_),
    .A1(_10851_),
    .B1(_10596_),
    .X(_10854_));
 sg13g2_and4_1 _17676_ (.A(_10839_),
    .B(_10841_),
    .C(_10848_),
    .D(_10854_),
    .X(_10855_));
 sg13g2_nor2_1 _17677_ (.A(_09539_),
    .B(net608),
    .Y(_10856_));
 sg13g2_a21o_1 _17678_ (.A2(_10855_),
    .A1(net608),
    .B1(_10856_),
    .X(_10857_));
 sg13g2_buf_1 _17679_ (.A(_10857_),
    .X(_10858_));
 sg13g2_nand2_1 _17680_ (.Y(_10859_),
    .A(net893),
    .B(net531));
 sg13g2_nor2_1 _17681_ (.A(net665),
    .B(_10817_),
    .Y(_10860_));
 sg13g2_inv_1 _17682_ (.Y(_10861_),
    .A(_08475_));
 sg13g2_or2_1 _17683_ (.X(_10862_),
    .B(net863),
    .A(net870));
 sg13g2_nand3_1 _17684_ (.B(net865),
    .C(\cpu.ex.r_14[4] ),
    .A(net746),
    .Y(_10863_));
 sg13g2_o21ai_1 _17685_ (.B1(_10863_),
    .Y(_10864_),
    .A1(_10861_),
    .A2(_10862_));
 sg13g2_inv_1 _17686_ (.Y(_10865_),
    .A(\cpu.ex.r_lr[4] ));
 sg13g2_nand3_1 _17687_ (.B(net745),
    .C(\cpu.ex.r_mult[20] ),
    .A(net746),
    .Y(_10866_));
 sg13g2_o21ai_1 _17688_ (.B1(_10866_),
    .Y(_10867_),
    .A1(_10865_),
    .A2(_10798_));
 sg13g2_a22oi_1 _17689_ (.Y(_10868_),
    .B1(_10867_),
    .B2(_10693_),
    .A2(_10864_),
    .A1(_10860_));
 sg13g2_mux2_1 _17690_ (.A0(\cpu.ex.r_epc[4] ),
    .A1(\cpu.ex.r_11[4] ),
    .S(_10635_),
    .X(_10869_));
 sg13g2_and2_1 _17691_ (.A(net741),
    .B(_10626_),
    .X(_10870_));
 sg13g2_buf_1 _17692_ (.A(\cpu.ex.r_sp[4] ),
    .X(_10871_));
 sg13g2_mux2_1 _17693_ (.A0(_10871_),
    .A1(\cpu.ex.r_stmp[4] ),
    .S(net745),
    .X(_10872_));
 sg13g2_nor2_1 _17694_ (.A(net739),
    .B(_10711_),
    .Y(_10873_));
 sg13g2_mux2_1 _17695_ (.A0(\cpu.ex.r_9[4] ),
    .A1(\cpu.ex.r_13[4] ),
    .S(_10602_),
    .X(_10874_));
 sg13g2_and3_1 _17696_ (.X(_10875_),
    .A(net739),
    .B(net663),
    .C(_10874_));
 sg13g2_a221oi_1 _17697_ (.B2(_10873_),
    .C1(_10875_),
    .B1(_10872_),
    .A1(_10869_),
    .Y(_10876_),
    .A2(_10870_));
 sg13g2_nor2b_1 _17698_ (.A(_00260_),
    .B_N(net742),
    .Y(_10877_));
 sg13g2_nor2b_1 _17699_ (.A(net745),
    .B_N(\cpu.ex.r_8[4] ),
    .Y(_10878_));
 sg13g2_a22oi_1 _17700_ (.Y(_10879_),
    .B1(_10878_),
    .B2(_10569_),
    .A2(_10877_),
    .A1(_10626_));
 sg13g2_nand3b_1 _17701_ (.B(_10630_),
    .C(\cpu.ex.r_12[4] ),
    .Y(_10880_),
    .A_N(_10600_));
 sg13g2_nand3b_1 _17702_ (.B(\cpu.ex.r_10[4] ),
    .C(net744),
    .Y(_10881_),
    .A_N(_10622_));
 sg13g2_a21o_1 _17703_ (.A2(_10881_),
    .A1(_10880_),
    .B1(net665),
    .X(_10882_));
 sg13g2_buf_1 _17704_ (.A(_10608_),
    .X(_10883_));
 sg13g2_a21o_1 _17705_ (.A2(_10882_),
    .A1(_10879_),
    .B1(net736),
    .X(_10884_));
 sg13g2_nand4_1 _17706_ (.B(_10868_),
    .C(_10876_),
    .A(_10648_),
    .Y(_10885_),
    .D(_10884_));
 sg13g2_a21oi_1 _17707_ (.A1(_10859_),
    .A2(_10885_),
    .Y(_10886_),
    .B1(_10742_));
 sg13g2_a21oi_1 _17708_ (.A1(_10835_),
    .A2(_10858_),
    .Y(_10887_),
    .B1(_10886_));
 sg13g2_inv_1 _17709_ (.Y(_10888_),
    .A(_09998_));
 sg13g2_buf_1 _17710_ (.A(_10888_),
    .X(_10889_));
 sg13g2_nand2_1 _17711_ (.Y(_10890_),
    .A(_10889_),
    .B(_10747_));
 sg13g2_and2_1 _17712_ (.A(net1009),
    .B(net1008),
    .X(_10891_));
 sg13g2_buf_2 _17713_ (.A(_10891_),
    .X(_10892_));
 sg13g2_a221oi_1 _17714_ (.B2(\cpu.ex.r_13[5] ),
    .C1(net746),
    .B1(_10892_),
    .A1(\cpu.ex.r_lr[5] ),
    .Y(_10893_),
    .A2(net872));
 sg13g2_inv_1 _17715_ (.Y(_10894_),
    .A(_00261_));
 sg13g2_a221oi_1 _17716_ (.B2(_10894_),
    .C1(_10596_),
    .B1(_10892_),
    .A1(\cpu.ex.r_epc[5] ),
    .Y(_10895_),
    .A2(net872));
 sg13g2_nor3_1 _17717_ (.A(_10620_),
    .B(_10893_),
    .C(_10895_),
    .Y(_10896_));
 sg13g2_nor2b_1 _17718_ (.A(net870),
    .B_N(net1006),
    .Y(_10897_));
 sg13g2_buf_1 _17719_ (.A(\cpu.ex.r_sp[5] ),
    .X(_10898_));
 sg13g2_a22oi_1 _17720_ (.Y(_10899_),
    .B1(_10681_),
    .B2(_10898_),
    .A2(_10897_),
    .A1(\cpu.ex.r_8[5] ));
 sg13g2_nand3b_1 _17721_ (.B(net742),
    .C(\cpu.ex.r_12[5] ),
    .Y(_10900_),
    .A_N(_10683_));
 sg13g2_nand3b_1 _17722_ (.B(\cpu.ex.r_9[5] ),
    .C(net748),
    .Y(_10901_),
    .A_N(_10622_));
 sg13g2_nand2b_1 _17723_ (.Y(_10902_),
    .B(net867),
    .A_N(net870));
 sg13g2_a21o_1 _17724_ (.A2(_10901_),
    .A1(_10900_),
    .B1(_10902_),
    .X(_10903_));
 sg13g2_o21ai_1 _17725_ (.B1(_10903_),
    .Y(_10904_),
    .A1(_10719_),
    .A2(_10899_));
 sg13g2_nand3_1 _17726_ (.B(net662),
    .C(_10892_),
    .A(\cpu.ex.r_14[5] ),
    .Y(_10905_));
 sg13g2_mux2_1 _17727_ (.A0(\cpu.ex.r_stmp[5] ),
    .A1(\cpu.ex.r_mult[21] ),
    .S(net740),
    .X(_10906_));
 sg13g2_nand3_1 _17728_ (.B(_10681_),
    .C(_10906_),
    .A(net664),
    .Y(_10907_));
 sg13g2_mux2_1 _17729_ (.A0(\cpu.ex.r_10[5] ),
    .A1(\cpu.ex.r_11[5] ),
    .S(_10683_),
    .X(_10908_));
 sg13g2_nand3_1 _17730_ (.B(_10592_),
    .C(_10908_),
    .A(_10601_),
    .Y(_10909_));
 sg13g2_nand3_1 _17731_ (.B(_10907_),
    .C(_10909_),
    .A(_10905_),
    .Y(_10910_));
 sg13g2_or4_1 _17732_ (.A(_10747_),
    .B(_10896_),
    .C(_10904_),
    .D(_10910_),
    .X(_10911_));
 sg13g2_a21oi_1 _17733_ (.A1(_10890_),
    .A2(_10911_),
    .Y(_10912_),
    .B1(_10742_));
 sg13g2_inv_1 _17734_ (.Y(_10913_),
    .A(_00269_));
 sg13g2_mux4_1 _17735_ (.S0(_10668_),
    .A0(_10913_),
    .A1(\cpu.ex.r_11[13] ),
    .A2(_10269_),
    .A3(\cpu.ex.r_epc[13] ),
    .S1(net736),
    .X(_10914_));
 sg13g2_mux2_1 _17736_ (.A0(\cpu.ex.r_sp[13] ),
    .A1(\cpu.ex.r_stmp[13] ),
    .S(net866),
    .X(_10915_));
 sg13g2_a22oi_1 _17737_ (.Y(_10916_),
    .B1(_10915_),
    .B2(net736),
    .A2(_10592_),
    .A1(\cpu.ex.r_10[13] ));
 sg13g2_a21oi_1 _17738_ (.A1(net743),
    .A2(_10916_),
    .Y(_10917_),
    .B1(net747));
 sg13g2_o21ai_1 _17739_ (.B1(_10917_),
    .Y(_10918_),
    .A1(net743),
    .A2(_10914_));
 sg13g2_nor2_1 _17740_ (.A(net741),
    .B(_10902_),
    .Y(_10919_));
 sg13g2_mux2_1 _17741_ (.A0(\cpu.ex.r_12[13] ),
    .A1(\cpu.ex.r_13[13] ),
    .S(net748),
    .X(_10920_));
 sg13g2_mux2_1 _17742_ (.A0(\cpu.ex.r_lr[13] ),
    .A1(_10304_),
    .S(net869),
    .X(_10921_));
 sg13g2_a22oi_1 _17743_ (.Y(_10922_),
    .B1(_10921_),
    .B2(_10608_),
    .A2(_10592_),
    .A1(\cpu.ex.r_9[13] ));
 sg13g2_inv_1 _17744_ (.Y(_10923_),
    .A(_10922_));
 sg13g2_a22oi_1 _17745_ (.Y(_10924_),
    .B1(_10724_),
    .B2(\cpu.ex.r_14[13] ),
    .A2(_10722_),
    .A1(\cpu.ex.r_8[13] ));
 sg13g2_nor2_1 _17746_ (.A(_10753_),
    .B(_10924_),
    .Y(_10925_));
 sg13g2_a221oi_1 _17747_ (.B2(net663),
    .C1(_10925_),
    .B1(_10923_),
    .A1(_10919_),
    .Y(_10926_),
    .A2(_10920_));
 sg13g2_and4_1 _17748_ (.A(net532),
    .B(_10835_),
    .C(_10918_),
    .D(_10926_),
    .X(_10927_));
 sg13g2_nand4_1 _17749_ (.B(_09376_),
    .C(_10556_),
    .A(_08489_),
    .Y(_10928_),
    .D(net531));
 sg13g2_nand2_1 _17750_ (.Y(_10929_),
    .A(\cpu.ex.c_mult_off[0] ),
    .B(_10928_));
 sg13g2_nor2_1 _17751_ (.A(_10711_),
    .B(_10793_),
    .Y(_10930_));
 sg13g2_mux4_1 _17752_ (.S0(net871),
    .A0(\cpu.ex.r_12[15] ),
    .A1(\cpu.ex.r_13[15] ),
    .A2(\cpu.ex.r_14[15] ),
    .A3(\cpu.ex.r_15[15] ),
    .S1(net868),
    .X(_10931_));
 sg13g2_and2_1 _17753_ (.A(_10892_),
    .B(_10931_),
    .X(_10932_));
 sg13g2_a21o_1 _17754_ (.A2(_10930_),
    .A1(\cpu.ex.r_10[15] ),
    .B1(_10932_),
    .X(_10933_));
 sg13g2_and2_1 _17755_ (.A(net866),
    .B(\cpu.ex.r_stmp[15] ),
    .X(_10934_));
 sg13g2_nor2b_1 _17756_ (.A(net742),
    .B_N(\cpu.ex.r_8[15] ),
    .Y(_10935_));
 sg13g2_a22oi_1 _17757_ (.Y(_10936_),
    .B1(_10935_),
    .B2(_10897_),
    .A2(_10934_),
    .A1(_10681_));
 sg13g2_buf_1 _17758_ (.A(\cpu.ex.r_sp[15] ),
    .X(_10937_));
 sg13g2_nand3b_1 _17759_ (.B(net744),
    .C(_10937_),
    .Y(_10938_),
    .A_N(net740));
 sg13g2_nand3b_1 _17760_ (.B(\cpu.ex.r_lr[15] ),
    .C(net740),
    .Y(_10939_),
    .A_N(net870));
 sg13g2_or2_1 _17761_ (.X(_10940_),
    .B(net866),
    .A(net863));
 sg13g2_a21o_1 _17762_ (.A2(_10939_),
    .A1(_10938_),
    .B1(_10940_),
    .X(_10941_));
 sg13g2_o21ai_1 _17763_ (.B1(_10941_),
    .Y(_10942_),
    .A1(net665),
    .A2(_10936_));
 sg13g2_nand3_1 _17764_ (.B(net872),
    .C(_10626_),
    .A(\cpu.ex.r_epc[15] ),
    .Y(_10943_));
 sg13g2_nand3b_1 _17765_ (.B(net863),
    .C(net740),
    .Y(_10944_),
    .A_N(net866));
 sg13g2_mux2_1 _17766_ (.A0(\cpu.ex.r_9[15] ),
    .A1(\cpu.ex.r_11[15] ),
    .S(net744),
    .X(_10945_));
 sg13g2_nand2b_1 _17767_ (.Y(_10946_),
    .B(_10945_),
    .A_N(_10944_));
 sg13g2_buf_1 _17768_ (.A(\cpu.ex.mmu_read[15] ),
    .X(_10947_));
 sg13g2_mux2_1 _17769_ (.A0(_10947_),
    .A1(\cpu.ex.r_mult[31] ),
    .S(_10600_),
    .X(_10948_));
 sg13g2_nand3_1 _17770_ (.B(_10693_),
    .C(_10948_),
    .A(_10631_),
    .Y(_10949_));
 sg13g2_nand3_1 _17771_ (.B(_10946_),
    .C(_10949_),
    .A(_10943_),
    .Y(_10950_));
 sg13g2_or4_1 _17772_ (.A(_10747_),
    .B(_10933_),
    .C(_10942_),
    .D(_10950_),
    .X(_10951_));
 sg13g2_a21oi_1 _17773_ (.A1(_09456_),
    .A2(_10747_),
    .Y(_10952_),
    .B1(net609));
 sg13g2_inv_1 _17774_ (.Y(_10953_),
    .A(\cpu.ex.r_sp[7] ));
 sg13g2_nand3_1 _17775_ (.B(net742),
    .C(\cpu.ex.r_mult[23] ),
    .A(net748),
    .Y(_10954_));
 sg13g2_o21ai_1 _17776_ (.B1(_10954_),
    .Y(_10955_),
    .A1(_10953_),
    .A2(_10719_));
 sg13g2_inv_1 _17777_ (.Y(_10956_),
    .A(\cpu.ex.r_lr[7] ));
 sg13g2_nand3_1 _17778_ (.B(net867),
    .C(\cpu.ex.r_11[7] ),
    .A(net738),
    .Y(_10957_));
 sg13g2_o21ai_1 _17779_ (.B1(_10957_),
    .Y(_10958_),
    .A1(_10956_),
    .A2(_10862_));
 sg13g2_nand3b_1 _17780_ (.B(net738),
    .C(\cpu.ex.r_10[7] ),
    .Y(_10959_),
    .A_N(_10585_));
 sg13g2_nand3b_1 _17781_ (.B(\cpu.ex.r_9[7] ),
    .C(net748),
    .Y(_10960_),
    .A_N(_10714_));
 sg13g2_a21oi_1 _17782_ (.A1(_10959_),
    .A2(_10960_),
    .Y(_10961_),
    .B1(_10793_));
 sg13g2_a221oi_1 _17783_ (.B2(_10623_),
    .C1(_10961_),
    .B1(_10958_),
    .A1(_10681_),
    .Y(_10962_),
    .A2(_10955_));
 sg13g2_nand3_1 _17784_ (.B(\cpu.ex.r_14[7] ),
    .C(_10606_),
    .A(_10603_),
    .Y(_10963_));
 sg13g2_nand3_1 _17785_ (.B(\cpu.ex.r_epc[7] ),
    .C(_10565_),
    .A(_10586_),
    .Y(_10964_));
 sg13g2_a21o_1 _17786_ (.A2(_10964_),
    .A1(_10963_),
    .B1(net747),
    .X(_10965_));
 sg13g2_mux2_1 _17787_ (.A0(\cpu.ex.r_8[7] ),
    .A1(\cpu.ex.r_12[7] ),
    .S(_10630_),
    .X(_10966_));
 sg13g2_nand2b_1 _17788_ (.Y(_10967_),
    .B(\cpu.ex.r_13[7] ),
    .A_N(_10714_));
 sg13g2_o21ai_1 _17789_ (.B1(_10967_),
    .Y(_10968_),
    .A1(_10596_),
    .A2(_00263_));
 sg13g2_buf_1 _17790_ (.A(\cpu.dec.user_io ),
    .X(_10969_));
 sg13g2_mux2_1 _17791_ (.A0(_10969_),
    .A1(\cpu.ex.r_stmp[7] ),
    .S(net870),
    .X(_10970_));
 sg13g2_and3_1 _17792_ (.X(_10971_),
    .A(net745),
    .B(_10789_),
    .C(_10970_));
 sg13g2_a221oi_1 _17793_ (.B2(_10678_),
    .C1(_10971_),
    .B1(_10968_),
    .A1(_10655_),
    .Y(_10972_),
    .A2(_10966_));
 sg13g2_nand4_1 _17794_ (.B(_10962_),
    .C(_10965_),
    .A(net608),
    .Y(_10973_),
    .D(_10972_));
 sg13g2_inv_1 _17795_ (.Y(_10974_),
    .A(_09204_));
 sg13g2_a21oi_1 _17796_ (.A1(_10974_),
    .A2(net531),
    .Y(_10975_),
    .B1(\cpu.ex.c_mult_off[3] ));
 sg13g2_a221oi_1 _17797_ (.B2(_10975_),
    .C1(net471),
    .B1(_10973_),
    .A1(_10951_),
    .Y(_10976_),
    .A2(_10952_));
 sg13g2_nor4_1 _17798_ (.A(_10912_),
    .B(_10927_),
    .C(_10929_),
    .D(_10976_),
    .Y(_10977_));
 sg13g2_a221oi_1 _17799_ (.B2(_10887_),
    .C1(_10977_),
    .B1(_10834_),
    .A1(net1004),
    .Y(_10978_),
    .A2(_10577_));
 sg13g2_buf_1 _17800_ (.A(_10978_),
    .X(_10979_));
 sg13g2_mux4_1 _17801_ (.S0(_10556_),
    .A0(_00195_),
    .A1(_00287_),
    .A2(_00293_),
    .A3(net1130),
    .S1(net609),
    .X(_10980_));
 sg13g2_buf_1 _17802_ (.A(_00294_),
    .X(_10981_));
 sg13g2_mux4_1 _17803_ (.S0(_10556_),
    .A0(_00194_),
    .A1(_00196_),
    .A2(_00292_),
    .A3(_10981_),
    .S1(net609),
    .X(_10982_));
 sg13g2_mux2_1 _17804_ (.A0(_10980_),
    .A1(_10982_),
    .S(\cpu.ex.c_mult_off[0] ),
    .X(_10983_));
 sg13g2_nand2_1 _17805_ (.Y(_10984_),
    .A(net1004),
    .B(_10983_));
 sg13g2_o21ai_1 _17806_ (.B1(_09375_),
    .Y(_10985_),
    .A1(_09362_),
    .A2(_09374_));
 sg13g2_nand3b_1 _17807_ (.B(_10985_),
    .C(_09371_),
    .Y(_10986_),
    .A_N(_10558_));
 sg13g2_buf_1 _17808_ (.A(_10986_),
    .X(\cpu.ex.c_mult_off[2] ));
 sg13g2_o21ai_1 _17809_ (.B1(\cpu.ex.c_mult_off[2] ),
    .Y(_10987_),
    .A1(_10736_),
    .A2(_10984_));
 sg13g2_nand2_1 _17810_ (.Y(_10988_),
    .A(net1126),
    .B(net613));
 sg13g2_a22oi_1 _17811_ (.Y(_10989_),
    .B1(_10344_),
    .B2(\cpu.ex.r_12[0] ),
    .A2(net875),
    .A1(\cpu.ex.r_stmp[0] ));
 sg13g2_and2_1 _17812_ (.A(\cpu.ex.r_10[0] ),
    .B(net1017),
    .X(_10990_));
 sg13g2_nor2b_1 _17813_ (.A(net881),
    .B_N(_09257_),
    .Y(_10991_));
 sg13g2_a22oi_1 _17814_ (.Y(_10992_),
    .B1(net880),
    .B2(_10991_),
    .A2(_10990_),
    .A1(_10265_));
 sg13g2_o21ai_1 _17815_ (.B1(_10992_),
    .Y(_10993_),
    .A1(net752),
    .A2(_10989_));
 sg13g2_mux2_1 _17816_ (.A0(\cpu.ex.r_9[0] ),
    .A1(\cpu.ex.r_13[0] ),
    .S(net1014),
    .X(_10994_));
 sg13g2_a22oi_1 _17817_ (.Y(_10995_),
    .B1(_10994_),
    .B2(_10340_),
    .A2(_10368_),
    .A1(\cpu.ex.r_11[0] ));
 sg13g2_nand3_1 _17818_ (.B(net881),
    .C(net880),
    .A(\cpu.ex.r_mult[16] ),
    .Y(_10996_));
 sg13g2_o21ai_1 _17819_ (.B1(_10996_),
    .Y(_10997_),
    .A1(_10355_),
    .A2(_10995_));
 sg13g2_mux2_1 _17820_ (.A0(_10993_),
    .A1(_10997_),
    .S(net759),
    .X(_10998_));
 sg13g2_a22oi_1 _17821_ (.Y(_10999_),
    .B1(_10388_),
    .B2(\cpu.ex.r_15[0] ),
    .A2(_10308_),
    .A1(_10762_));
 sg13g2_nor2_1 _17822_ (.A(net1017),
    .B(net1014),
    .Y(_11000_));
 sg13g2_a22oi_1 _17823_ (.Y(_11001_),
    .B1(_11000_),
    .B2(\cpu.ex.r_8[0] ),
    .A2(_10458_),
    .A1(\cpu.ex.r_14[0] ));
 sg13g2_nand2b_1 _17824_ (.Y(_11002_),
    .B(_10299_),
    .A_N(_11001_));
 sg13g2_o21ai_1 _17825_ (.B1(_11002_),
    .Y(_11003_),
    .A1(_10448_),
    .A2(_10999_));
 sg13g2_o21ai_1 _17826_ (.B1(_10335_),
    .Y(_11004_),
    .A1(_10998_),
    .A2(_11003_));
 sg13g2_nor2_1 _17827_ (.A(_10408_),
    .B(_10322_),
    .Y(_11005_));
 sg13g2_and3_1 _17828_ (.X(_11006_),
    .A(_10988_),
    .B(_11004_),
    .C(_11005_));
 sg13g2_buf_1 _17829_ (.A(_11006_),
    .X(_11007_));
 sg13g2_buf_1 _17830_ (.A(\cpu.dec.imm[0] ),
    .X(_11008_));
 sg13g2_nor3_1 _17831_ (.A(_11008_),
    .B(net1109),
    .C(_10322_),
    .Y(_11009_));
 sg13g2_or2_1 _17832_ (.X(_11010_),
    .B(_11009_),
    .A(net1012));
 sg13g2_buf_1 _17833_ (.A(_11010_),
    .X(_11011_));
 sg13g2_nor3_1 _17834_ (.A(_11007_),
    .B(_11011_),
    .C(_10519_),
    .Y(_11012_));
 sg13g2_o21ai_1 _17835_ (.B1(_11012_),
    .Y(_11013_),
    .A1(_10979_),
    .A2(_10987_));
 sg13g2_nor3_1 _17836_ (.A(_10666_),
    .B(_10779_),
    .C(_11013_),
    .Y(_11014_));
 sg13g2_nand3_1 _17837_ (.B(_11004_),
    .C(_11005_),
    .A(_10988_),
    .Y(_11015_));
 sg13g2_buf_1 _17838_ (.A(_11015_),
    .X(_11016_));
 sg13g2_nor2_1 _17839_ (.A(net1012),
    .B(_11009_),
    .Y(_11017_));
 sg13g2_and4_1 _17840_ (.A(_11016_),
    .B(_11017_),
    .C(_10549_),
    .D(_10550_),
    .X(_11018_));
 sg13g2_buf_8 _17841_ (.A(_11018_),
    .X(_11019_));
 sg13g2_o21ai_1 _17842_ (.B1(_11019_),
    .Y(_11020_),
    .A1(_10979_),
    .A2(_10987_));
 sg13g2_nand3_1 _17843_ (.B(_10444_),
    .C(net663),
    .A(net664),
    .Y(_11021_));
 sg13g2_nand3_1 _17844_ (.B(_10436_),
    .C(net662),
    .A(net737),
    .Y(_11022_));
 sg13g2_a21oi_1 _17845_ (.A1(_11021_),
    .A2(_11022_),
    .Y(_11023_),
    .B1(net739));
 sg13g2_nand3_1 _17846_ (.B(\cpu.ex.r_10[3] ),
    .C(_10606_),
    .A(net737),
    .Y(_11024_));
 sg13g2_nand3_1 _17847_ (.B(\cpu.ex.r_mult[19] ),
    .C(_10590_),
    .A(net665),
    .Y(_11025_));
 sg13g2_a21oi_1 _17848_ (.A1(_11024_),
    .A2(_11025_),
    .Y(_11026_),
    .B1(net747));
 sg13g2_nand3_1 _17849_ (.B(\cpu.ex.r_13[3] ),
    .C(net663),
    .A(net739),
    .Y(_11027_));
 sg13g2_nand3_1 _17850_ (.B(\cpu.ex.r_stmp[3] ),
    .C(net662),
    .A(net736),
    .Y(_11028_));
 sg13g2_a21oi_1 _17851_ (.A1(_11027_),
    .A2(_11028_),
    .Y(_11029_),
    .B1(net737));
 sg13g2_nor3_1 _17852_ (.A(_11023_),
    .B(_11026_),
    .C(_11029_),
    .Y(_11030_));
 sg13g2_mux2_1 _17853_ (.A0(\cpu.ex.r_12[3] ),
    .A1(\cpu.ex.r_14[3] ),
    .S(net746),
    .X(_11031_));
 sg13g2_nand2_1 _17854_ (.Y(_11032_),
    .A(net746),
    .B(\cpu.ex.r_11[3] ));
 sg13g2_nand2b_1 _17855_ (.Y(_11033_),
    .B(\cpu.ex.r_9[3] ),
    .A_N(net738));
 sg13g2_a21oi_1 _17856_ (.A1(_11032_),
    .A2(_11033_),
    .Y(_11034_),
    .B1(_10944_));
 sg13g2_a221oi_1 _17857_ (.B2(_11031_),
    .C1(_11034_),
    .B1(_10786_),
    .A1(\cpu.ex.r_epc[3] ),
    .Y(_11035_),
    .A2(_10628_));
 sg13g2_a22oi_1 _17858_ (.Y(_11036_),
    .B1(_10592_),
    .B2(\cpu.ex.r_8[3] ),
    .A2(_10590_),
    .A1(net1129));
 sg13g2_nand2b_1 _17859_ (.Y(_11037_),
    .B(_10569_),
    .A_N(_11036_));
 sg13g2_nor2b_1 _17860_ (.A(net738),
    .B_N(\cpu.ex.r_lr[3] ),
    .Y(_11038_));
 sg13g2_nor2b_1 _17861_ (.A(_00259_),
    .B_N(net742),
    .Y(_11039_));
 sg13g2_a22oi_1 _17862_ (.Y(_11040_),
    .B1(_10617_),
    .B2(_11039_),
    .A2(_11038_),
    .A1(net872));
 sg13g2_nand2b_1 _17863_ (.Y(_11041_),
    .B(net665),
    .A_N(_11040_));
 sg13g2_and4_1 _17864_ (.A(net608),
    .B(_11035_),
    .C(_11037_),
    .D(_11041_),
    .X(_11042_));
 sg13g2_a22oi_1 _17865_ (.Y(_11043_),
    .B1(_11030_),
    .B2(_11042_),
    .A2(net531),
    .A1(_09341_));
 sg13g2_buf_2 _17866_ (.A(_11043_),
    .X(_11044_));
 sg13g2_mux2_1 _17867_ (.A0(\cpu.ex.r_12[11] ),
    .A1(\cpu.ex.r_13[11] ),
    .S(net748),
    .X(_11045_));
 sg13g2_nand3b_1 _17868_ (.B(net865),
    .C(\cpu.ex.r_8[11] ),
    .Y(_11046_),
    .A_N(net738));
 sg13g2_nand3b_1 _17869_ (.B(_10395_),
    .C(net746),
    .Y(_11047_),
    .A_N(net867));
 sg13g2_a21oi_1 _17870_ (.A1(_11046_),
    .A2(_11047_),
    .Y(_11048_),
    .B1(_10719_));
 sg13g2_a221oi_1 _17871_ (.B2(_11045_),
    .C1(_11048_),
    .B1(_10919_),
    .A1(\cpu.ex.r_10[11] ),
    .Y(_11049_),
    .A2(_10930_));
 sg13g2_inv_1 _17872_ (.Y(_11050_),
    .A(_00267_));
 sg13g2_mux4_1 _17873_ (.S0(_10668_),
    .A0(_11050_),
    .A1(\cpu.ex.r_11[11] ),
    .A2(\cpu.ex.r_mult[27] ),
    .A3(\cpu.ex.r_epc[11] ),
    .S1(net736),
    .X(_11051_));
 sg13g2_nand2_1 _17874_ (.Y(_11052_),
    .A(_10626_),
    .B(_11051_));
 sg13g2_nand3_1 _17875_ (.B(\cpu.ex.r_9[11] ),
    .C(_10634_),
    .A(_10669_),
    .Y(_11053_));
 sg13g2_nand3_1 _17876_ (.B(\cpu.ex.r_14[11] ),
    .C(_10686_),
    .A(net745),
    .Y(_11054_));
 sg13g2_a21o_1 _17877_ (.A2(_11054_),
    .A1(_11053_),
    .B1(net736),
    .X(_11055_));
 sg13g2_nand3_1 _17878_ (.B(\cpu.ex.r_lr[11] ),
    .C(net663),
    .A(_10669_),
    .Y(_11056_));
 sg13g2_nand3_1 _17879_ (.B(\cpu.ex.r_stmp[11] ),
    .C(net662),
    .A(net745),
    .Y(_11057_));
 sg13g2_a21o_1 _17880_ (.A2(_11057_),
    .A1(_11056_),
    .B1(_10695_),
    .X(_11058_));
 sg13g2_nand4_1 _17881_ (.B(_11052_),
    .C(_11055_),
    .A(_11049_),
    .Y(_11059_),
    .D(_11058_));
 sg13g2_mux2_1 _17882_ (.A0(net1107),
    .A1(_11059_),
    .S(_10659_),
    .X(_11060_));
 sg13g2_buf_2 _17883_ (.A(_11060_),
    .X(_11061_));
 sg13g2_a22oi_1 _17884_ (.Y(_11062_),
    .B1(_10693_),
    .B2(\cpu.ex.mmu_read[1] ),
    .A2(_10606_),
    .A1(\cpu.ex.r_12[1] ));
 sg13g2_o21ai_1 _17885_ (.B1(net747),
    .Y(_11063_),
    .A1(net737),
    .A2(_11062_));
 sg13g2_a22oi_1 _17886_ (.Y(_11064_),
    .B1(_10592_),
    .B2(\cpu.ex.r_11[1] ),
    .A2(_10590_),
    .A1(\cpu.ex.r_mult[17] ));
 sg13g2_inv_1 _17887_ (.Y(_11065_),
    .A(_00257_));
 sg13g2_nor2b_1 _17888_ (.A(_10585_),
    .B_N(_10539_),
    .Y(_11066_));
 sg13g2_a221oi_1 _17889_ (.B2(_10565_),
    .C1(_10597_),
    .B1(_11066_),
    .A1(_11065_),
    .Y(_11067_),
    .A2(_10678_));
 sg13g2_o21ai_1 _17890_ (.B1(_11067_),
    .Y(_11068_),
    .A1(_10620_),
    .A2(_11064_));
 sg13g2_nand3_1 _17891_ (.B(\cpu.ex.r_8[1] ),
    .C(_10569_),
    .A(net739),
    .Y(_11069_));
 sg13g2_nand3_1 _17892_ (.B(\cpu.ex.r_epc[1] ),
    .C(_10626_),
    .A(_10883_),
    .Y(_11070_));
 sg13g2_nand2_1 _17893_ (.Y(_11071_),
    .A(_11069_),
    .B(_11070_));
 sg13g2_mux2_1 _17894_ (.A0(_10526_),
    .A1(\cpu.ex.r_stmp[1] ),
    .S(net738),
    .X(_11072_));
 sg13g2_nand3_1 _17895_ (.B(_10789_),
    .C(_11072_),
    .A(net664),
    .Y(_11073_));
 sg13g2_mux2_1 _17896_ (.A0(\cpu.ex.r_lr[1] ),
    .A1(\cpu.ex.r_9[1] ),
    .S(net867),
    .X(_11074_));
 sg13g2_nand3_1 _17897_ (.B(net663),
    .C(_11074_),
    .A(net737),
    .Y(_11075_));
 sg13g2_nand3_1 _17898_ (.B(net662),
    .C(_10892_),
    .A(\cpu.ex.r_14[1] ),
    .Y(_11076_));
 sg13g2_nand3_1 _17899_ (.B(_11075_),
    .C(_11076_),
    .A(_11073_),
    .Y(_11077_));
 sg13g2_a221oi_1 _17900_ (.B2(net737),
    .C1(_11077_),
    .B1(_11071_),
    .A1(_11063_),
    .Y(_11078_),
    .A2(_11068_));
 sg13g2_nand3_1 _17901_ (.B(\cpu.ex.r_13[1] ),
    .C(net663),
    .A(net664),
    .Y(_11079_));
 sg13g2_nand3_1 _17902_ (.B(\cpu.ex.r_10[1] ),
    .C(net662),
    .A(_10817_),
    .Y(_11080_));
 sg13g2_a21oi_1 _17903_ (.A1(_11079_),
    .A2(_11080_),
    .Y(_11081_),
    .B1(net736));
 sg13g2_nor2_1 _17904_ (.A(net531),
    .B(_11081_),
    .Y(_11082_));
 sg13g2_a22oi_1 _17905_ (.Y(_11083_),
    .B1(_11078_),
    .B2(_11082_),
    .A2(net531),
    .A1(_10050_));
 sg13g2_buf_2 _17906_ (.A(_11083_),
    .X(_11084_));
 sg13g2_buf_2 _17907_ (.A(\cpu.addr[9] ),
    .X(_11085_));
 sg13g2_a221oi_1 _17908_ (.B2(\cpu.ex.r_11[9] ),
    .C1(net745),
    .B1(_10626_),
    .A1(\cpu.ex.r_8[9] ),
    .Y(_11086_),
    .A2(_10569_));
 sg13g2_a221oi_1 _17909_ (.B2(\cpu.ex.r_14[9] ),
    .C1(_10668_),
    .B1(_10651_),
    .A1(\cpu.ex.r_13[9] ),
    .Y(_11087_),
    .A2(_10633_));
 sg13g2_nor3_1 _17910_ (.A(_10883_),
    .B(_11086_),
    .C(_11087_),
    .Y(_11088_));
 sg13g2_a22oi_1 _17911_ (.Y(_11089_),
    .B1(_10681_),
    .B2(\cpu.ex.r_epc[9] ),
    .A2(_10897_),
    .A1(\cpu.ex.r_9[9] ));
 sg13g2_nor2b_1 _17912_ (.A(_11089_),
    .B_N(_10623_),
    .Y(_11090_));
 sg13g2_inv_1 _17913_ (.Y(_11091_),
    .A(\cpu.ex.r_10[9] ));
 sg13g2_nand3b_1 _17914_ (.B(net869),
    .C(net740),
    .Y(_11092_),
    .A_N(_00265_));
 sg13g2_o21ai_1 _17915_ (.B1(_11092_),
    .Y(_11093_),
    .A1(_11091_),
    .A2(_10719_));
 sg13g2_nand3b_1 _17916_ (.B(_10688_),
    .C(\cpu.ex.r_12[9] ),
    .Y(_11094_),
    .A_N(net870));
 sg13g2_nand3b_1 _17917_ (.B(\cpu.ex.r_stmp[9] ),
    .C(net870),
    .Y(_11095_),
    .A_N(net1006));
 sg13g2_nand2b_1 _17918_ (.Y(_11096_),
    .B(net742),
    .A_N(net740));
 sg13g2_a21oi_1 _17919_ (.A1(_11094_),
    .A2(_11095_),
    .Y(_11097_),
    .B1(_11096_));
 sg13g2_a21o_1 _17920_ (.A2(_11093_),
    .A1(_10617_),
    .B1(_11097_),
    .X(_11098_));
 sg13g2_nand2_1 _17921_ (.Y(_11099_),
    .A(net665),
    .B(_10608_));
 sg13g2_a22oi_1 _17922_ (.Y(_11100_),
    .B1(_10724_),
    .B2(\cpu.ex.r_mult[25] ),
    .A2(_10722_),
    .A1(\cpu.ex.r_lr[9] ));
 sg13g2_buf_1 _17923_ (.A(\cpu.ex.r_sp[9] ),
    .X(_11101_));
 sg13g2_nand3_1 _17924_ (.B(net872),
    .C(net662),
    .A(_11101_),
    .Y(_11102_));
 sg13g2_o21ai_1 _17925_ (.B1(_11102_),
    .Y(_11103_),
    .A1(_11099_),
    .A2(_11100_));
 sg13g2_or4_1 _17926_ (.A(_11088_),
    .B(_11090_),
    .C(_11098_),
    .D(_11103_),
    .X(_11104_));
 sg13g2_mux2_1 _17927_ (.A0(_11085_),
    .A1(_11104_),
    .S(_10659_),
    .X(_11105_));
 sg13g2_buf_2 _17928_ (.A(_11105_),
    .X(_11106_));
 sg13g2_mux4_1 _17929_ (.S0(\cpu.ex.c_mult_off[3] ),
    .A0(_11044_),
    .A1(_11061_),
    .A2(_11084_),
    .A3(_11106_),
    .S1(net471),
    .X(_11107_));
 sg13g2_a21oi_1 _17930_ (.A1(net1004),
    .A2(_10577_),
    .Y(_11108_),
    .B1(_11107_));
 sg13g2_buf_2 _17931_ (.A(_00290_),
    .X(_11109_));
 sg13g2_buf_1 _17932_ (.A(_00200_),
    .X(_11110_));
 sg13g2_mux4_1 _17933_ (.S0(net471),
    .A0(_00288_),
    .A1(_11109_),
    .A2(_00191_),
    .A3(_11110_),
    .S1(net609),
    .X(_11111_));
 sg13g2_and2_1 _17934_ (.A(\cpu.ex.c_mult_off[0] ),
    .B(_11111_),
    .X(_11112_));
 sg13g2_nor2_1 _17935_ (.A(_10579_),
    .B(_10736_),
    .Y(_11113_));
 sg13g2_buf_2 _17936_ (.A(_11113_),
    .X(_11114_));
 sg13g2_a221oi_1 _17937_ (.B2(_11114_),
    .C1(\cpu.ex.c_mult_off[2] ),
    .B1(_11112_),
    .A1(\cpu.ex.c_mult_off[0] ),
    .Y(_11115_),
    .A2(_11108_));
 sg13g2_a21oi_1 _17938_ (.A1(_11013_),
    .A2(_11020_),
    .Y(_11116_),
    .B1(_11115_));
 sg13g2_nor3_1 _17939_ (.A(_10666_),
    .B(_10779_),
    .C(_11020_),
    .Y(_11117_));
 sg13g2_nor4_2 _17940_ (.A(_10553_),
    .B(_11014_),
    .C(_11116_),
    .Y(_11118_),
    .D(_11117_));
 sg13g2_o21ai_1 _17941_ (.B1(_11118_),
    .Y(_11119_),
    .A1(_10507_),
    .A2(_10517_));
 sg13g2_nor3_1 _17942_ (.A(net1105),
    .B(net694),
    .C(_10505_),
    .Y(_11120_));
 sg13g2_nor2_1 _17943_ (.A(net694),
    .B(_10505_),
    .Y(_11121_));
 sg13g2_buf_1 _17944_ (.A(_10513_),
    .X(_11122_));
 sg13g2_nor3_1 _17945_ (.A(_10508_),
    .B(net694),
    .C(net240),
    .Y(_11123_));
 sg13g2_a221oi_1 _17946_ (.B2(_10515_),
    .C1(_11123_),
    .B1(_11121_),
    .A1(_11118_),
    .Y(_11124_),
    .A2(_11120_));
 sg13g2_buf_1 _17947_ (.A(_11124_),
    .X(_11125_));
 sg13g2_and2_1 _17948_ (.A(_11119_),
    .B(_11125_),
    .X(_11126_));
 sg13g2_nand2_1 _17949_ (.Y(_11127_),
    .A(_08819_),
    .B(net1012));
 sg13g2_a22oi_1 _17950_ (.Y(_11128_),
    .B1(_10454_),
    .B2(\cpu.ex.r_11[8] ),
    .A2(_10452_),
    .A1(_10682_));
 sg13g2_nand2b_1 _17951_ (.Y(_11129_),
    .B(_10368_),
    .A_N(_11128_));
 sg13g2_nand3_1 _17952_ (.B(_10355_),
    .C(_10357_),
    .A(\cpu.ex.r_epc[8] ),
    .Y(_11130_));
 sg13g2_nand3_1 _17953_ (.B(net760),
    .C(_10345_),
    .A(\cpu.ex.r_8[8] ),
    .Y(_11131_));
 sg13g2_a21oi_1 _17954_ (.A1(_11130_),
    .A2(_11131_),
    .Y(_11132_),
    .B1(_10287_));
 sg13g2_nand3_1 _17955_ (.B(_10341_),
    .C(_10266_),
    .A(\cpu.ex.r_9[8] ),
    .Y(_11133_));
 sg13g2_nand3_1 _17956_ (.B(_10279_),
    .C(net875),
    .A(\cpu.ex.r_mult[24] ),
    .Y(_11134_));
 sg13g2_a21oi_1 _17957_ (.A1(_11133_),
    .A2(_11134_),
    .Y(_11135_),
    .B1(net760));
 sg13g2_nand3_1 _17958_ (.B(net752),
    .C(_10360_),
    .A(\cpu.ex.r_lr[8] ),
    .Y(_11136_));
 sg13g2_nand3_1 _17959_ (.B(net758),
    .C(_10290_),
    .A(\cpu.ex.r_stmp[8] ),
    .Y(_11137_));
 sg13g2_a21oi_1 _17960_ (.A1(_11136_),
    .A2(_11137_),
    .Y(_11138_),
    .B1(net757));
 sg13g2_nor2b_1 _17961_ (.A(_00264_),
    .B_N(net761),
    .Y(_11139_));
 sg13g2_nor2b_1 _17962_ (.A(_10256_),
    .B_N(\cpu.ex.r_13[8] ),
    .Y(_11140_));
 sg13g2_and3_1 _17963_ (.X(_11141_),
    .A(_10277_),
    .B(net757),
    .C(net878));
 sg13g2_o21ai_1 _17964_ (.B1(_11141_),
    .Y(_11142_),
    .A1(_11139_),
    .A2(_11140_));
 sg13g2_nand3_1 _17965_ (.B(_10388_),
    .C(_10290_),
    .A(\cpu.ex.r_14[8] ),
    .Y(_11143_));
 sg13g2_nand3b_1 _17966_ (.B(net878),
    .C(\cpu.ex.r_12[8] ),
    .Y(_11144_),
    .A_N(net881));
 sg13g2_nand3b_1 _17967_ (.B(net761),
    .C(\cpu.ex.r_10[8] ),
    .Y(_11145_),
    .A_N(net878));
 sg13g2_nand2b_1 _17968_ (.Y(_11146_),
    .B(net877),
    .A_N(net879));
 sg13g2_buf_2 _17969_ (.A(_11146_),
    .X(_11147_));
 sg13g2_a21o_1 _17970_ (.A2(_11145_),
    .A1(_11144_),
    .B1(_11147_),
    .X(_11148_));
 sg13g2_nand3_1 _17971_ (.B(_11143_),
    .C(_11148_),
    .A(_11142_),
    .Y(_11149_));
 sg13g2_nor4_1 _17972_ (.A(_11132_),
    .B(_11135_),
    .C(_11138_),
    .D(_11149_),
    .Y(_11150_));
 sg13g2_a21oi_1 _17973_ (.A1(_11129_),
    .A2(_11150_),
    .Y(_11151_),
    .B1(_10315_));
 sg13g2_and2_1 _17974_ (.A(_09202_),
    .B(net613),
    .X(_11152_));
 sg13g2_nor3_1 _17975_ (.A(_10408_),
    .B(_11151_),
    .C(_11152_),
    .Y(_11153_));
 sg13g2_nor2_1 _17976_ (.A(net1013),
    .B(\cpu.dec.imm[8] ),
    .Y(_11154_));
 sg13g2_o21ai_1 _17977_ (.B1(_10413_),
    .Y(_11155_),
    .A1(_11153_),
    .A2(_11154_));
 sg13g2_buf_1 _17978_ (.A(_11155_),
    .X(_11156_));
 sg13g2_nand2_1 _17979_ (.Y(_11157_),
    .A(_11127_),
    .B(_11156_));
 sg13g2_buf_2 _17980_ (.A(_11157_),
    .X(_11158_));
 sg13g2_buf_1 _17981_ (.A(_00301_),
    .X(_11159_));
 sg13g2_nor2_1 _17982_ (.A(net1102),
    .B(_09370_),
    .Y(_11160_));
 sg13g2_and2_1 _17983_ (.A(_11127_),
    .B(_11156_),
    .X(_11161_));
 sg13g2_buf_1 _17984_ (.A(_11161_),
    .X(_11162_));
 sg13g2_mux2_1 _17985_ (.A0(net1102),
    .A1(_11160_),
    .S(_11162_),
    .X(_11163_));
 sg13g2_buf_2 _17986_ (.A(_00299_),
    .X(_11164_));
 sg13g2_nand2b_1 _17987_ (.Y(_11165_),
    .B(_10325_),
    .A_N(_08807_));
 sg13g2_buf_1 _17988_ (.A(_11165_),
    .X(_11166_));
 sg13g2_nor2_1 _17989_ (.A(net666),
    .B(_11147_),
    .Y(_11167_));
 sg13g2_mux2_1 _17990_ (.A0(\cpu.ex.r_12[10] ),
    .A1(\cpu.ex.r_14[10] ),
    .S(net672),
    .X(_11168_));
 sg13g2_inv_1 _17991_ (.Y(_11169_),
    .A(\cpu.ex.r_8[10] ));
 sg13g2_nand3b_1 _17992_ (.B(net667),
    .C(\cpu.ex.r_lr[10] ),
    .Y(_11170_),
    .A_N(net669));
 sg13g2_o21ai_1 _17993_ (.B1(_11170_),
    .Y(_11171_),
    .A1(_11169_),
    .A2(_11147_));
 sg13g2_nand2b_1 _17994_ (.Y(_11172_),
    .B(net669),
    .A_N(_00266_));
 sg13g2_nand2b_1 _17995_ (.Y(_11173_),
    .B(net1106),
    .A_N(net669));
 sg13g2_a21oi_1 _17996_ (.A1(_11172_),
    .A2(_11173_),
    .Y(_11174_),
    .B1(_10275_));
 sg13g2_a221oi_1 _17997_ (.B2(_11000_),
    .C1(_11174_),
    .B1(_11171_),
    .A1(_11167_),
    .Y(_11175_),
    .A2(_11168_));
 sg13g2_a22oi_1 _17998_ (.Y(_11176_),
    .B1(net751),
    .B2(\cpu.ex.r_9[10] ),
    .A2(net755),
    .A1(\cpu.ex.r_10[10] ));
 sg13g2_nand2b_1 _17999_ (.Y(_11177_),
    .B(net670),
    .A_N(_11176_));
 sg13g2_mux2_1 _18000_ (.A0(_10716_),
    .A1(\cpu.ex.r_stmp[10] ),
    .S(net756),
    .X(_11178_));
 sg13g2_and2_1 _18001_ (.A(\cpu.ex.r_11[10] ),
    .B(net667),
    .X(_11179_));
 sg13g2_a22oi_1 _18002_ (.Y(_11180_),
    .B1(_11179_),
    .B2(net670),
    .A2(_11178_),
    .A1(_10452_));
 sg13g2_nand2b_1 _18003_ (.Y(_11181_),
    .B(net612),
    .A_N(_11180_));
 sg13g2_nand3_1 _18004_ (.B(net668),
    .C(net753),
    .A(\cpu.ex.r_13[10] ),
    .Y(_11182_));
 sg13g2_nand3_1 _18005_ (.B(net666),
    .C(net875),
    .A(\cpu.ex.r_epc[10] ),
    .Y(_11183_));
 sg13g2_a21o_1 _18006_ (.A2(_11183_),
    .A1(_11182_),
    .B1(net671),
    .X(_11184_));
 sg13g2_nand4_1 _18007_ (.B(_11177_),
    .C(_11181_),
    .A(_11175_),
    .Y(_11185_),
    .D(_11184_));
 sg13g2_a221oi_1 _18008_ (.B2(_11185_),
    .C1(net873),
    .B1(net533),
    .A1(net1104),
    .Y(_11186_),
    .A2(net534));
 sg13g2_nor2_1 _18009_ (.A(_10319_),
    .B(\cpu.dec.imm[10] ),
    .Y(_11187_));
 sg13g2_o21ai_1 _18010_ (.B1(_10414_),
    .Y(_11188_),
    .A1(_11186_),
    .A2(_11187_));
 sg13g2_buf_2 _18011_ (.A(_11188_),
    .X(_11189_));
 sg13g2_and2_1 _18012_ (.A(_11166_),
    .B(_11189_),
    .X(_11190_));
 sg13g2_buf_2 _18013_ (.A(_11190_),
    .X(_11191_));
 sg13g2_a221oi_1 _18014_ (.B2(_11164_),
    .C1(_11191_),
    .B1(_11163_),
    .A1(net694),
    .Y(_11192_),
    .A2(_11158_));
 sg13g2_xnor2_1 _18015_ (.Y(_11193_),
    .A(net1102),
    .B(_11158_));
 sg13g2_nor2_1 _18016_ (.A(_11164_),
    .B(net694),
    .Y(_11194_));
 sg13g2_nand2_1 _18017_ (.Y(_11195_),
    .A(_11166_),
    .B(_11189_));
 sg13g2_a21oi_1 _18018_ (.A1(_11193_),
    .A2(_11194_),
    .Y(_11196_),
    .B1(_11195_));
 sg13g2_nand2_1 _18019_ (.Y(_11197_),
    .A(_08787_),
    .B(_10326_));
 sg13g2_nand2_1 _18020_ (.Y(_11198_),
    .A(\cpu.ex.r_13[9] ),
    .B(_10369_));
 sg13g2_nor2b_1 _18021_ (.A(_00265_),
    .B_N(net758),
    .Y(_11199_));
 sg13g2_nor2b_1 _18022_ (.A(net758),
    .B_N(\cpu.ex.r_11[9] ),
    .Y(_11200_));
 sg13g2_o21ai_1 _18023_ (.B1(_10257_),
    .Y(_11201_),
    .A1(_11199_),
    .A2(_11200_));
 sg13g2_a21oi_1 _18024_ (.A1(_11198_),
    .A2(_11201_),
    .Y(_11202_),
    .B1(_10262_));
 sg13g2_and2_1 _18025_ (.A(\cpu.ex.r_8[9] ),
    .B(_10280_),
    .X(_11203_));
 sg13g2_o21ai_1 _18026_ (.B1(_10286_),
    .Y(_11204_),
    .A1(_11202_),
    .A2(_11203_));
 sg13g2_nand3_1 _18027_ (.B(net752),
    .C(net875),
    .A(_11101_),
    .Y(_11205_));
 sg13g2_nand3_1 _18028_ (.B(net756),
    .C(net753),
    .A(\cpu.ex.r_12[9] ),
    .Y(_11206_));
 sg13g2_nand3_1 _18029_ (.B(_11205_),
    .C(_11206_),
    .A(net760),
    .Y(_11207_));
 sg13g2_nand3_1 _18030_ (.B(net754),
    .C(net670),
    .A(\cpu.ex.r_9[9] ),
    .Y(_11208_));
 sg13g2_nand3_1 _18031_ (.B(_10257_),
    .C(net880),
    .A(\cpu.ex.r_mult[25] ),
    .Y(_11209_));
 sg13g2_nand3_1 _18032_ (.B(_11208_),
    .C(_11209_),
    .A(net667),
    .Y(_11210_));
 sg13g2_and2_1 _18033_ (.A(\cpu.ex.r_14[9] ),
    .B(net758),
    .X(_11211_));
 sg13g2_a21oi_1 _18034_ (.A1(\cpu.ex.r_10[9] ),
    .A2(net752),
    .Y(_11212_),
    .B1(_11211_));
 sg13g2_nand3_1 _18035_ (.B(_10295_),
    .C(_10308_),
    .A(\cpu.ex.r_epc[9] ),
    .Y(_11213_));
 sg13g2_o21ai_1 _18036_ (.B1(_11213_),
    .Y(_11214_),
    .A1(_11147_),
    .A2(_11212_));
 sg13g2_nand3_1 _18037_ (.B(net756),
    .C(net755),
    .A(\cpu.ex.r_stmp[9] ),
    .Y(_11215_));
 sg13g2_nand3_1 _18038_ (.B(_10352_),
    .C(net751),
    .A(\cpu.ex.r_lr[9] ),
    .Y(_11216_));
 sg13g2_a21oi_1 _18039_ (.A1(_11215_),
    .A2(_11216_),
    .Y(_11217_),
    .B1(_10286_));
 sg13g2_a221oi_1 _18040_ (.B2(net612),
    .C1(_11217_),
    .B1(_11214_),
    .A1(_11207_),
    .Y(_11218_),
    .A2(_11210_));
 sg13g2_a21oi_1 _18041_ (.A1(_11204_),
    .A2(_11218_),
    .Y(_11219_),
    .B1(_10315_));
 sg13g2_nand2_1 _18042_ (.Y(_11220_),
    .A(_11085_),
    .B(_10252_));
 sg13g2_inv_1 _18043_ (.Y(_11221_),
    .A(_11220_));
 sg13g2_o21ai_1 _18044_ (.B1(net1013),
    .Y(_11222_),
    .A1(_11219_),
    .A2(_11221_));
 sg13g2_nand2_1 _18045_ (.Y(_11223_),
    .A(net873),
    .B(\cpu.dec.imm[9] ));
 sg13g2_nand3_1 _18046_ (.B(_11222_),
    .C(_11223_),
    .A(_10414_),
    .Y(_11224_));
 sg13g2_buf_1 _18047_ (.A(_11224_),
    .X(_11225_));
 sg13g2_nand2_1 _18048_ (.Y(_11226_),
    .A(_11197_),
    .B(_11225_));
 sg13g2_buf_1 _18049_ (.A(_11226_),
    .X(_11227_));
 sg13g2_buf_1 _18050_ (.A(_00300_),
    .X(_11228_));
 sg13g2_nor2_1 _18051_ (.A(_11228_),
    .B(_09370_),
    .Y(_11229_));
 sg13g2_xnor2_1 _18052_ (.Y(_11230_),
    .A(net217),
    .B(_11229_));
 sg13g2_nor3_1 _18053_ (.A(_11192_),
    .B(_11196_),
    .C(_11230_),
    .Y(_11231_));
 sg13g2_buf_1 _18054_ (.A(_00302_),
    .X(_11232_));
 sg13g2_nand2b_1 _18055_ (.Y(_11233_),
    .B(_10325_),
    .A_N(_08777_));
 sg13g2_buf_1 _18056_ (.A(_11233_),
    .X(_11234_));
 sg13g2_nand3_1 _18057_ (.B(_10279_),
    .C(net753),
    .A(\cpu.ex.r_12[6] ),
    .Y(_11235_));
 sg13g2_nand3_1 _18058_ (.B(net752),
    .C(net875),
    .A(_10788_),
    .Y(_11236_));
 sg13g2_nand3_1 _18059_ (.B(net754),
    .C(net670),
    .A(\cpu.ex.r_8[6] ),
    .Y(_11237_));
 sg13g2_nand3_1 _18060_ (.B(net761),
    .C(_10268_),
    .A(\cpu.ex.r_stmp[6] ),
    .Y(_11238_));
 sg13g2_and4_1 _18061_ (.A(_11235_),
    .B(_11236_),
    .C(_11237_),
    .D(_11238_),
    .X(_11239_));
 sg13g2_and2_1 _18062_ (.A(_10255_),
    .B(_10268_),
    .X(_11240_));
 sg13g2_nor2_2 _18063_ (.A(net761),
    .B(_10478_),
    .Y(_11241_));
 sg13g2_a221oi_1 _18064_ (.B2(\cpu.ex.r_9[6] ),
    .C1(net760),
    .B1(_11241_),
    .A1(_10802_),
    .Y(_11242_),
    .A2(_11240_));
 sg13g2_a21o_1 _18065_ (.A2(_11239_),
    .A1(net760),
    .B1(_11242_),
    .X(_11243_));
 sg13g2_and2_1 _18066_ (.A(\cpu.ex.r_14[6] ),
    .B(_10290_),
    .X(_11244_));
 sg13g2_nand2b_1 _18067_ (.Y(_11245_),
    .B(net761),
    .A_N(_00262_));
 sg13g2_nand2b_1 _18068_ (.Y(_11246_),
    .B(\cpu.ex.r_13[6] ),
    .A_N(net761));
 sg13g2_a21oi_1 _18069_ (.A1(_11245_),
    .A2(_11246_),
    .Y(_11247_),
    .B1(_10261_));
 sg13g2_o21ai_1 _18070_ (.B1(_10284_),
    .Y(_11248_),
    .A1(_11244_),
    .A2(_11247_));
 sg13g2_nand3b_1 _18071_ (.B(net759),
    .C(\cpu.ex.r_epc[6] ),
    .Y(_11249_),
    .A_N(_10283_));
 sg13g2_o21ai_1 _18072_ (.B1(_11249_),
    .Y(_11250_),
    .A1(_10792_),
    .A2(_11147_));
 sg13g2_and3_1 _18073_ (.X(_11251_),
    .A(\cpu.ex.r_11[6] ),
    .B(net881),
    .C(net877));
 sg13g2_a21o_1 _18074_ (.A2(_10294_),
    .A1(\cpu.ex.r_lr[6] ),
    .B1(_11251_),
    .X(_11252_));
 sg13g2_a221oi_1 _18075_ (.B2(_10277_),
    .C1(net756),
    .B1(_11252_),
    .A1(net672),
    .Y(_11253_),
    .A2(_11250_));
 sg13g2_a21o_1 _18076_ (.A2(_11248_),
    .A1(net756),
    .B1(_11253_),
    .X(_11254_));
 sg13g2_a21oi_1 _18077_ (.A1(_11243_),
    .A2(_11254_),
    .Y(_11255_),
    .B1(_10315_));
 sg13g2_and2_1 _18078_ (.A(_09206_),
    .B(_10252_),
    .X(_11256_));
 sg13g2_nor3_1 _18079_ (.A(_10408_),
    .B(_11255_),
    .C(_11256_),
    .Y(_11257_));
 sg13g2_nor2_1 _18080_ (.A(net1013),
    .B(\cpu.dec.imm[6] ),
    .Y(_11258_));
 sg13g2_o21ai_1 _18081_ (.B1(net750),
    .Y(_11259_),
    .A1(_11257_),
    .A2(_11258_));
 sg13g2_buf_1 _18082_ (.A(_11259_),
    .X(_11260_));
 sg13g2_nand2_1 _18083_ (.Y(_11261_),
    .A(_11234_),
    .B(_11260_));
 sg13g2_buf_1 _18084_ (.A(_11261_),
    .X(_11262_));
 sg13g2_xnor2_1 _18085_ (.Y(_11263_),
    .A(net1101),
    .B(_11262_));
 sg13g2_buf_1 _18086_ (.A(_10802_),
    .X(_11264_));
 sg13g2_inv_1 _18087_ (.Y(_11265_),
    .A(net1003));
 sg13g2_a221oi_1 _18088_ (.B2(\cpu.ex.r_13[7] ),
    .C1(net672),
    .B1(_10454_),
    .A1(_10969_),
    .Y(_11266_),
    .A2(_10452_));
 sg13g2_nor2b_1 _18089_ (.A(_10284_),
    .B_N(net759),
    .Y(_11267_));
 sg13g2_a221oi_1 _18090_ (.B2(\cpu.ex.r_mult[23] ),
    .C1(net754),
    .B1(_11267_),
    .A1(\cpu.ex.r_14[7] ),
    .Y(_11268_),
    .A2(_10299_));
 sg13g2_o21ai_1 _18091_ (.B1(net756),
    .Y(_11269_),
    .A1(_11266_),
    .A2(_11268_));
 sg13g2_nand3_1 _18092_ (.B(net757),
    .C(net755),
    .A(\cpu.ex.r_10[7] ),
    .Y(_11270_));
 sg13g2_mux2_1 _18093_ (.A0(\cpu.ex.r_9[7] ),
    .A1(\cpu.ex.r_11[7] ),
    .S(net761),
    .X(_11271_));
 sg13g2_nand2_1 _18094_ (.Y(_11272_),
    .A(_10454_),
    .B(_11271_));
 sg13g2_nand3_1 _18095_ (.B(net759),
    .C(_10294_),
    .A(\cpu.ex.r_lr[7] ),
    .Y(_11273_));
 sg13g2_nand4_1 _18096_ (.B(_11270_),
    .C(_11272_),
    .A(net666),
    .Y(_11274_),
    .D(_11273_));
 sg13g2_nor2b_1 _18097_ (.A(_00263_),
    .B_N(_10454_),
    .Y(_11275_));
 sg13g2_a21o_1 _18098_ (.A2(_10452_),
    .A1(\cpu.ex.r_stmp[7] ),
    .B1(_11275_),
    .X(_11276_));
 sg13g2_and2_1 _18099_ (.A(\cpu.ex.r_epc[7] ),
    .B(net759),
    .X(_11277_));
 sg13g2_a21oi_1 _18100_ (.A1(\cpu.ex.r_sp[7] ),
    .A2(net760),
    .Y(_11278_),
    .B1(_11277_));
 sg13g2_mux2_1 _18101_ (.A0(\cpu.ex.r_8[7] ),
    .A1(\cpu.ex.r_12[7] ),
    .S(net878),
    .X(_11279_));
 sg13g2_nand3_1 _18102_ (.B(_10345_),
    .C(_11279_),
    .A(net760),
    .Y(_11280_));
 sg13g2_o21ai_1 _18103_ (.B1(_11280_),
    .Y(_11281_),
    .A1(_10481_),
    .A2(_11278_));
 sg13g2_a221oi_1 _18104_ (.B2(_10458_),
    .C1(_11281_),
    .B1(_11276_),
    .A1(_11269_),
    .Y(_11282_),
    .A2(_11274_));
 sg13g2_nand2_1 _18105_ (.Y(_11283_),
    .A(_09204_),
    .B(net613));
 sg13g2_o21ai_1 _18106_ (.B1(_11283_),
    .Y(_11284_),
    .A1(_10315_),
    .A2(_11282_));
 sg13g2_inv_1 _18107_ (.Y(_11285_),
    .A(\cpu.dec.imm[7] ));
 sg13g2_a21oi_1 _18108_ (.A1(net873),
    .A2(_11285_),
    .Y(_11286_),
    .B1(net1012));
 sg13g2_o21ai_1 _18109_ (.B1(_11286_),
    .Y(_11287_),
    .A1(_10409_),
    .A2(_11284_));
 sg13g2_buf_1 _18110_ (.A(_11287_),
    .X(_11288_));
 sg13g2_and2_1 _18111_ (.A(_08797_),
    .B(net1012),
    .X(_11289_));
 sg13g2_a21oi_1 _18112_ (.A1(_10467_),
    .A2(_10322_),
    .Y(_11290_),
    .B1(_11289_));
 sg13g2_and2_1 _18113_ (.A(_11288_),
    .B(_11290_),
    .X(_11291_));
 sg13g2_buf_1 _18114_ (.A(_11291_),
    .X(_11292_));
 sg13g2_nor2_1 _18115_ (.A(_11265_),
    .B(_11292_),
    .Y(_11293_));
 sg13g2_nor3_1 _18116_ (.A(net1003),
    .B(net1101),
    .C(_11262_),
    .Y(_11294_));
 sg13g2_buf_1 _18117_ (.A(_11292_),
    .X(_11295_));
 sg13g2_a22oi_1 _18118_ (.Y(_11296_),
    .B1(_11294_),
    .B2(net216),
    .A2(_11293_),
    .A1(_11263_));
 sg13g2_a21oi_1 _18119_ (.A1(_11265_),
    .A2(net1101),
    .Y(_11297_),
    .B1(_09378_));
 sg13g2_and2_1 _18120_ (.A(_11234_),
    .B(_11260_),
    .X(_11298_));
 sg13g2_buf_1 _18121_ (.A(_11298_),
    .X(_11299_));
 sg13g2_nand2_1 _18122_ (.Y(_11300_),
    .A(_11288_),
    .B(_11290_));
 sg13g2_buf_1 _18123_ (.A(_11300_),
    .X(_11301_));
 sg13g2_nor2_1 _18124_ (.A(_11299_),
    .B(net239),
    .Y(_11302_));
 sg13g2_nand2b_1 _18125_ (.Y(_11303_),
    .B(_11302_),
    .A_N(_11297_));
 sg13g2_o21ai_1 _18126_ (.B1(_11303_),
    .Y(_11304_),
    .A1(_09378_),
    .A2(_11296_));
 sg13g2_nor3_1 _18127_ (.A(_09811_),
    .B(_10240_),
    .C(_10250_),
    .Y(_11305_));
 sg13g2_nor2b_1 _18128_ (.A(_10259_),
    .B_N(net874),
    .Y(_11306_));
 sg13g2_nor2b_1 _18129_ (.A(_10390_),
    .B_N(_10259_),
    .Y(_11307_));
 sg13g2_a221oi_1 _18130_ (.B2(\cpu.ex.r_lr[4] ),
    .C1(net757),
    .B1(_11307_),
    .A1(_08475_),
    .Y(_11308_),
    .A2(_11306_));
 sg13g2_a221oi_1 _18131_ (.B2(\cpu.ex.r_9[4] ),
    .C1(_10355_),
    .B1(_11307_),
    .A1(\cpu.ex.r_12[4] ),
    .Y(_11309_),
    .A2(_11306_));
 sg13g2_o21ai_1 _18132_ (.B1(net754),
    .Y(_11310_),
    .A1(_11308_),
    .A2(_11309_));
 sg13g2_mux2_1 _18133_ (.A0(\cpu.ex.r_10[4] ),
    .A1(\cpu.ex.r_14[4] ),
    .S(_10390_),
    .X(_11311_));
 sg13g2_a22oi_1 _18134_ (.Y(_11312_),
    .B1(_11311_),
    .B2(_10260_),
    .A2(_11307_),
    .A1(\cpu.ex.r_11[4] ));
 sg13g2_nor2b_1 _18135_ (.A(_10276_),
    .B_N(_10871_),
    .Y(_11313_));
 sg13g2_nor2b_1 _18136_ (.A(_00260_),
    .B_N(_10276_),
    .Y(_11314_));
 sg13g2_a221oi_1 _18137_ (.B2(_10388_),
    .C1(_10340_),
    .B1(_11314_),
    .A1(_10308_),
    .Y(_11315_),
    .A2(_11313_));
 sg13g2_o21ai_1 _18138_ (.B1(_11315_),
    .Y(_11316_),
    .A1(_10355_),
    .A2(_11312_));
 sg13g2_and3_1 _18139_ (.X(_11317_),
    .A(_10335_),
    .B(_11310_),
    .C(_11316_));
 sg13g2_a221oi_1 _18140_ (.B2(\cpu.ex.r_8[4] ),
    .C1(net759),
    .B1(_11241_),
    .A1(\cpu.ex.r_stmp[4] ),
    .Y(_11318_),
    .A2(_11240_));
 sg13g2_mux2_1 _18141_ (.A0(\cpu.ex.r_epc[4] ),
    .A1(\cpu.ex.r_mult[20] ),
    .S(_10278_),
    .X(_11319_));
 sg13g2_a221oi_1 _18142_ (.B2(net875),
    .C1(_10261_),
    .B1(_11319_),
    .A1(\cpu.ex.r_13[4] ),
    .Y(_11320_),
    .A2(_10392_));
 sg13g2_nor3_1 _18143_ (.A(_10315_),
    .B(_11318_),
    .C(_11320_),
    .Y(_11321_));
 sg13g2_or4_1 _18144_ (.A(_10497_),
    .B(_11305_),
    .C(_11317_),
    .D(_11321_),
    .X(_11322_));
 sg13g2_buf_1 _18145_ (.A(_11322_),
    .X(_11323_));
 sg13g2_nor4_1 _18146_ (.A(net1109),
    .B(_10321_),
    .C(_10322_),
    .D(\cpu.dec.imm[4] ),
    .Y(_11324_));
 sg13g2_a21oi_2 _18147_ (.B1(_11324_),
    .Y(_11325_),
    .A2(net1012),
    .A1(_08817_));
 sg13g2_nand2_1 _18148_ (.Y(_11326_),
    .A(_11323_),
    .B(_11325_));
 sg13g2_buf_2 _18149_ (.A(_11326_),
    .X(_11327_));
 sg13g2_buf_1 _18150_ (.A(_00304_),
    .X(_11328_));
 sg13g2_nor2_2 _18151_ (.A(_11328_),
    .B(_09370_),
    .Y(_11329_));
 sg13g2_nand2_1 _18152_ (.Y(_11330_),
    .A(_11327_),
    .B(_11329_));
 sg13g2_and2_1 _18153_ (.A(_11323_),
    .B(_11325_),
    .X(_11331_));
 sg13g2_buf_8 _18154_ (.A(_11331_),
    .X(_11332_));
 sg13g2_nand2b_1 _18155_ (.Y(_11333_),
    .B(net287),
    .A_N(_11329_));
 sg13g2_buf_1 _18156_ (.A(_11333_),
    .X(_11334_));
 sg13g2_and2_1 _18157_ (.A(_11330_),
    .B(_11334_),
    .X(_11335_));
 sg13g2_nor2_1 _18158_ (.A(_08829_),
    .B(_10467_),
    .Y(_11336_));
 sg13g2_mux2_1 _18159_ (.A0(\cpu.ex.r_stmp[5] ),
    .A1(\cpu.ex.r_14[5] ),
    .S(net757),
    .X(_11337_));
 sg13g2_a22oi_1 _18160_ (.Y(_11338_),
    .B1(_11337_),
    .B2(net672),
    .A2(net753),
    .A1(\cpu.ex.r_12[5] ));
 sg13g2_nor2_1 _18161_ (.A(net666),
    .B(_11338_),
    .Y(_11339_));
 sg13g2_and2_1 _18162_ (.A(\cpu.ex.r_8[5] ),
    .B(_11241_),
    .X(_11340_));
 sg13g2_o21ai_1 _18163_ (.B1(_10262_),
    .Y(_11341_),
    .A1(_11339_),
    .A2(_11340_));
 sg13g2_a22oi_1 _18164_ (.Y(_11342_),
    .B1(net751),
    .B2(\cpu.ex.r_9[5] ),
    .A2(_10291_),
    .A1(\cpu.ex.r_10[5] ));
 sg13g2_a221oi_1 _18165_ (.B2(\cpu.ex.r_lr[5] ),
    .C1(net757),
    .B1(net751),
    .A1(_10898_),
    .Y(_11343_),
    .A2(net755));
 sg13g2_a21oi_1 _18166_ (.A1(net669),
    .A2(_11342_),
    .Y(_11344_),
    .B1(_11343_));
 sg13g2_nand2b_1 _18167_ (.Y(_11345_),
    .B(net758),
    .A_N(_00261_));
 sg13g2_nand2b_1 _18168_ (.Y(_11346_),
    .B(\cpu.ex.r_11[5] ),
    .A_N(net878));
 sg13g2_a21oi_1 _18169_ (.A1(_11345_),
    .A2(_11346_),
    .Y(_11347_),
    .B1(_10341_));
 sg13g2_a21o_1 _18170_ (.A2(_10369_),
    .A1(\cpu.ex.r_13[5] ),
    .B1(_11347_),
    .X(_11348_));
 sg13g2_and2_1 _18171_ (.A(\cpu.ex.r_mult[21] ),
    .B(net758),
    .X(_11349_));
 sg13g2_a21oi_1 _18172_ (.A1(\cpu.ex.r_epc[5] ),
    .A2(_10352_),
    .Y(_11350_),
    .B1(_11349_));
 sg13g2_nor3_1 _18173_ (.A(_10285_),
    .B(_10448_),
    .C(_11350_),
    .Y(_11351_));
 sg13g2_a221oi_1 _18174_ (.B2(_10454_),
    .C1(_11351_),
    .B1(_11348_),
    .A1(_10353_),
    .Y(_11352_),
    .A2(_11344_));
 sg13g2_a21o_1 _18175_ (.A2(_11352_),
    .A1(_11341_),
    .B1(_10315_),
    .X(_11353_));
 sg13g2_buf_1 _18176_ (.A(_11353_),
    .X(_11354_));
 sg13g2_nand2_1 _18177_ (.Y(_11355_),
    .A(_09998_),
    .B(net613));
 sg13g2_a21o_1 _18178_ (.A2(_11355_),
    .A1(_11354_),
    .B1(net873),
    .X(_11356_));
 sg13g2_nand2_1 _18179_ (.Y(_11357_),
    .A(net873),
    .B(\cpu.dec.imm[5] ));
 sg13g2_and3_1 _18180_ (.X(_11358_),
    .A(net750),
    .B(_11356_),
    .C(_11357_));
 sg13g2_buf_1 _18181_ (.A(_11358_),
    .X(_11359_));
 sg13g2_nor2_1 _18182_ (.A(_11336_),
    .B(_11359_),
    .Y(_11360_));
 sg13g2_buf_2 _18183_ (.A(_11360_),
    .X(_11361_));
 sg13g2_buf_2 _18184_ (.A(_00303_),
    .X(_11362_));
 sg13g2_nor2_2 _18185_ (.A(_11362_),
    .B(_09370_),
    .Y(_11363_));
 sg13g2_xnor2_1 _18186_ (.Y(_11364_),
    .A(_11361_),
    .B(_11363_));
 sg13g2_nand4_1 _18187_ (.B(_11304_),
    .C(_11335_),
    .A(_11231_),
    .Y(_11365_),
    .D(_11364_));
 sg13g2_and2_1 _18188_ (.A(_11164_),
    .B(_11191_),
    .X(_11366_));
 sg13g2_inv_1 _18189_ (.Y(_11367_),
    .A(_11228_));
 sg13g2_nor2_1 _18190_ (.A(_08786_),
    .B(_10467_),
    .Y(_11368_));
 sg13g2_and3_1 _18191_ (.X(_11369_),
    .A(net750),
    .B(_11222_),
    .C(_11223_));
 sg13g2_buf_1 _18192_ (.A(_11369_),
    .X(_11370_));
 sg13g2_nor2_1 _18193_ (.A(_11368_),
    .B(_11370_),
    .Y(_11371_));
 sg13g2_buf_1 _18194_ (.A(_11371_),
    .X(_11372_));
 sg13g2_o21ai_1 _18195_ (.B1(net215),
    .Y(_11373_),
    .A1(net1102),
    .A2(_11162_));
 sg13g2_nor3_1 _18196_ (.A(net1102),
    .B(_11371_),
    .C(_11162_),
    .Y(_11374_));
 sg13g2_a21oi_1 _18197_ (.A1(_11367_),
    .A2(_11373_),
    .Y(_11375_),
    .B1(_11374_));
 sg13g2_buf_1 _18198_ (.A(_11195_),
    .X(_11376_));
 sg13g2_nand2b_1 _18199_ (.Y(_11377_),
    .B(net214),
    .A_N(_11164_));
 sg13g2_o21ai_1 _18200_ (.B1(_11377_),
    .Y(_11378_),
    .A1(_11366_),
    .A2(_11375_));
 sg13g2_buf_1 _18201_ (.A(_11299_),
    .X(_11379_));
 sg13g2_nand2_1 _18202_ (.Y(_11380_),
    .A(net1003),
    .B(net749));
 sg13g2_nor2_1 _18203_ (.A(net194),
    .B(_11380_),
    .Y(_11381_));
 sg13g2_and2_1 _18204_ (.A(_11327_),
    .B(_11329_),
    .X(_11382_));
 sg13g2_buf_1 _18205_ (.A(_11382_),
    .X(_11383_));
 sg13g2_nor3_1 _18206_ (.A(_11383_),
    .B(_11336_),
    .C(_11359_),
    .Y(_11384_));
 sg13g2_inv_1 _18207_ (.Y(_11385_),
    .A(_11363_));
 sg13g2_o21ai_1 _18208_ (.B1(_11383_),
    .Y(_11386_),
    .A1(_11336_),
    .A2(_11359_));
 sg13g2_o21ai_1 _18209_ (.B1(_11386_),
    .Y(_11387_),
    .A1(_11384_),
    .A2(_11385_));
 sg13g2_o21ai_1 _18210_ (.B1(_11387_),
    .Y(_11388_),
    .A1(_11302_),
    .A2(_11381_));
 sg13g2_nor2_1 _18211_ (.A(_00302_),
    .B(_09370_),
    .Y(_11389_));
 sg13g2_and2_1 _18212_ (.A(_11292_),
    .B(_11389_),
    .X(_11390_));
 sg13g2_nor3_1 _18213_ (.A(_11265_),
    .B(net1101),
    .C(net694),
    .Y(_11391_));
 sg13g2_o21ai_1 _18214_ (.B1(_11387_),
    .Y(_11392_),
    .A1(_11390_),
    .A2(_11391_));
 sg13g2_buf_1 _18215_ (.A(_11262_),
    .X(_11393_));
 sg13g2_o21ai_1 _18216_ (.B1(net193),
    .Y(_11394_),
    .A1(_11390_),
    .A2(_11391_));
 sg13g2_or2_1 _18217_ (.X(_11395_),
    .B(_11380_),
    .A(net239));
 sg13g2_nand4_1 _18218_ (.B(_11392_),
    .C(_11394_),
    .A(_11388_),
    .Y(_11396_),
    .D(_11395_));
 sg13g2_a22oi_1 _18219_ (.Y(_11397_),
    .B1(_11231_),
    .B2(_11396_),
    .A2(_11378_),
    .A1(_10428_));
 sg13g2_o21ai_1 _18220_ (.B1(_11397_),
    .Y(_11398_),
    .A1(_11126_),
    .A2(_11365_));
 sg13g2_buf_8 _18221_ (.A(_11398_),
    .X(_11399_));
 sg13g2_buf_1 _18222_ (.A(_10382_),
    .X(_11400_));
 sg13g2_xnor2_1 _18223_ (.Y(_11401_),
    .A(_10331_),
    .B(net213));
 sg13g2_inv_1 _18224_ (.Y(_11402_),
    .A(net1011));
 sg13g2_nor2_1 _18225_ (.A(_11402_),
    .B(net170),
    .Y(_11403_));
 sg13g2_nor3_1 _18226_ (.A(_10424_),
    .B(_10331_),
    .C(net213),
    .Y(_11404_));
 sg13g2_a22oi_1 _18227_ (.Y(_11405_),
    .B1(_11404_),
    .B2(net170),
    .A2(_11403_),
    .A1(_11401_));
 sg13g2_o21ai_1 _18228_ (.B1(net749),
    .Y(_11406_),
    .A1(_10424_),
    .A2(_10384_));
 sg13g2_nand3_1 _18229_ (.B(net213),
    .C(_11406_),
    .A(net170),
    .Y(_11407_));
 sg13g2_o21ai_1 _18230_ (.B1(_11407_),
    .Y(_11408_),
    .A1(_09379_),
    .A2(_11405_));
 sg13g2_and2_1 _18231_ (.A(_10385_),
    .B(_10415_),
    .X(_11409_));
 sg13g2_buf_2 _18232_ (.A(_11409_),
    .X(_11410_));
 sg13g2_buf_1 _18233_ (.A(_11410_),
    .X(_11411_));
 sg13g2_nand2_1 _18234_ (.Y(_11412_),
    .A(net1106),
    .B(net749));
 sg13g2_nand2_1 _18235_ (.Y(_11413_),
    .A(net212),
    .B(_11412_));
 sg13g2_nand3_1 _18236_ (.B(_11408_),
    .C(_11413_),
    .A(_11399_),
    .Y(_11414_));
 sg13g2_buf_1 _18237_ (.A(_11414_),
    .X(_11415_));
 sg13g2_buf_1 _18238_ (.A(net749),
    .X(_11416_));
 sg13g2_inv_1 _18239_ (.Y(_11417_),
    .A(\cpu.dec.imm[15] ));
 sg13g2_nand3_1 _18240_ (.B(net670),
    .C(_10357_),
    .A(\cpu.ex.r_11[15] ),
    .Y(_11418_));
 sg13g2_nand3_1 _18241_ (.B(_11000_),
    .C(_10454_),
    .A(\cpu.ex.r_9[15] ),
    .Y(_11419_));
 sg13g2_nand2_1 _18242_ (.Y(_11420_),
    .A(_11418_),
    .B(_11419_));
 sg13g2_a22oi_1 _18243_ (.Y(_11421_),
    .B1(_10434_),
    .B2(_10937_),
    .A2(_10392_),
    .A1(\cpu.ex.r_12[15] ));
 sg13g2_mux2_1 _18244_ (.A0(\cpu.ex.r_stmp[15] ),
    .A1(\cpu.ex.r_14[15] ),
    .S(_10285_),
    .X(_11422_));
 sg13g2_mux2_1 _18245_ (.A0(_10947_),
    .A1(\cpu.ex.r_mult[31] ),
    .S(net672),
    .X(_11423_));
 sg13g2_a22oi_1 _18246_ (.Y(_11424_),
    .B1(_11423_),
    .B2(_11267_),
    .A2(_11422_),
    .A1(net755));
 sg13g2_nand2b_1 _18247_ (.Y(_11425_),
    .B(_10288_),
    .A_N(_11424_));
 sg13g2_o21ai_1 _18248_ (.B1(_11425_),
    .Y(_11426_),
    .A1(net610),
    .A2(_11421_));
 sg13g2_inv_1 _18249_ (.Y(_11427_),
    .A(\cpu.ex.r_epc[15] ));
 sg13g2_nand3_1 _18250_ (.B(net611),
    .C(net668),
    .A(\cpu.ex.r_15[15] ),
    .Y(_11428_));
 sg13g2_o21ai_1 _18251_ (.B1(_11428_),
    .Y(_11429_),
    .A1(_11427_),
    .A2(_10433_));
 sg13g2_nor2_1 _18252_ (.A(net610),
    .B(_10478_),
    .Y(_11430_));
 sg13g2_a22oi_1 _18253_ (.Y(_11431_),
    .B1(_11430_),
    .B2(\cpu.ex.r_10[15] ),
    .A2(_11429_),
    .A1(_10296_));
 sg13g2_inv_1 _18254_ (.Y(_11432_),
    .A(\cpu.ex.r_lr[15] ));
 sg13g2_nand3_1 _18255_ (.B(net611),
    .C(_10288_),
    .A(\cpu.ex.r_13[15] ),
    .Y(_11433_));
 sg13g2_o21ai_1 _18256_ (.B1(_11433_),
    .Y(_11434_),
    .A1(_11432_),
    .A2(_10433_));
 sg13g2_a221oi_1 _18257_ (.B2(net610),
    .C1(_10258_),
    .B1(_11434_),
    .A1(\cpu.ex.r_8[15] ),
    .Y(_11435_),
    .A2(_11430_));
 sg13g2_a21oi_1 _18258_ (.A1(_10258_),
    .A2(_11431_),
    .Y(_11436_),
    .B1(_11435_));
 sg13g2_or3_1 _18259_ (.A(_11420_),
    .B(_11426_),
    .C(_11436_),
    .X(_11437_));
 sg13g2_a22oi_1 _18260_ (.Y(_11438_),
    .B1(net533),
    .B2(_11437_),
    .A2(net534),
    .A1(net1059));
 sg13g2_mux2_1 _18261_ (.A0(_11417_),
    .A1(_11438_),
    .S(net1013),
    .X(_11439_));
 sg13g2_a22oi_1 _18262_ (.Y(_11440_),
    .B1(net750),
    .B2(_11439_),
    .A2(net876),
    .A1(_08703_));
 sg13g2_buf_1 _18263_ (.A(_11440_),
    .X(_11441_));
 sg13g2_buf_1 _18264_ (.A(_11441_),
    .X(_11442_));
 sg13g2_inv_1 _18265_ (.Y(_11443_),
    .A(_10269_));
 sg13g2_a21oi_1 _18266_ (.A1(_00297_),
    .A2(net169),
    .Y(_11444_),
    .B1(_11443_));
 sg13g2_nand2_1 _18267_ (.Y(_11445_),
    .A(net661),
    .B(_11444_));
 sg13g2_inv_1 _18268_ (.Y(_11446_),
    .A(\cpu.dec.imm[14] ));
 sg13g2_a22oi_1 _18269_ (.Y(_11447_),
    .B1(net751),
    .B2(\cpu.ex.r_lr[14] ),
    .A2(net755),
    .A1(_10825_));
 sg13g2_mux2_1 _18270_ (.A0(\cpu.ex.r_12[14] ),
    .A1(\cpu.ex.r_14[14] ),
    .S(net612),
    .X(_11448_));
 sg13g2_mux2_1 _18271_ (.A0(\cpu.ex.r_8[14] ),
    .A1(\cpu.ex.r_9[14] ),
    .S(net610),
    .X(_11449_));
 sg13g2_a22oi_1 _18272_ (.Y(_11450_),
    .B1(_11449_),
    .B2(_11241_),
    .A2(_11448_),
    .A1(_11167_));
 sg13g2_o21ai_1 _18273_ (.B1(_11450_),
    .Y(_11451_),
    .A1(_10433_),
    .A2(_11447_));
 sg13g2_inv_1 _18274_ (.Y(_11452_),
    .A(\cpu.ex.r_11[14] ));
 sg13g2_nand2_1 _18275_ (.Y(_11453_),
    .A(\cpu.ex.r_mult[30] ),
    .B(net880));
 sg13g2_o21ai_1 _18276_ (.B1(_11453_),
    .Y(_11454_),
    .A1(_11452_),
    .A2(_10478_));
 sg13g2_inv_1 _18277_ (.Y(_11455_),
    .A(\cpu.ex.r_10[14] ));
 sg13g2_nand2_1 _18278_ (.Y(_11456_),
    .A(\cpu.ex.r_epc[14] ),
    .B(_11267_));
 sg13g2_o21ai_1 _18279_ (.B1(_11456_),
    .Y(_11457_),
    .A1(_11455_),
    .A2(_11147_));
 sg13g2_a22oi_1 _18280_ (.Y(_11458_),
    .B1(_11457_),
    .B2(_10368_),
    .A2(_11454_),
    .A1(_10357_));
 sg13g2_nand3_1 _18281_ (.B(net671),
    .C(net875),
    .A(\cpu.ex.r_stmp[14] ),
    .Y(_11459_));
 sg13g2_nand3_1 _18282_ (.B(net610),
    .C(net753),
    .A(\cpu.ex.r_13[14] ),
    .Y(_11460_));
 sg13g2_a21oi_1 _18283_ (.A1(_11459_),
    .A2(_11460_),
    .Y(_11461_),
    .B1(net666));
 sg13g2_a22oi_1 _18284_ (.Y(_11462_),
    .B1(_10473_),
    .B2(_10828_),
    .A2(_10294_),
    .A1(_10815_));
 sg13g2_nor2_1 _18285_ (.A(_10471_),
    .B(_11462_),
    .Y(_11463_));
 sg13g2_nor2_1 _18286_ (.A(_11461_),
    .B(_11463_),
    .Y(_11464_));
 sg13g2_nand3b_1 _18287_ (.B(_11458_),
    .C(_11464_),
    .Y(_11465_),
    .A_N(_11451_));
 sg13g2_a22oi_1 _18288_ (.Y(_11466_),
    .B1(net533),
    .B2(_11465_),
    .A2(net534),
    .A1(net678));
 sg13g2_mux2_1 _18289_ (.A0(_11446_),
    .A1(_11466_),
    .S(net1013),
    .X(_11467_));
 sg13g2_a22oi_1 _18290_ (.Y(_11468_),
    .B1(net750),
    .B2(_11467_),
    .A2(net876),
    .A1(_08871_));
 sg13g2_buf_2 _18291_ (.A(_11468_),
    .X(_11469_));
 sg13g2_buf_1 _18292_ (.A(_11469_),
    .X(_11470_));
 sg13g2_nand2b_1 _18293_ (.Y(_11471_),
    .B(_10428_),
    .A_N(_00297_));
 sg13g2_or2_1 _18294_ (.X(_11472_),
    .B(_11471_),
    .A(net192));
 sg13g2_a22oi_1 _18295_ (.Y(_11473_),
    .B1(_11445_),
    .B2(_11472_),
    .A2(_11415_),
    .A1(_10430_));
 sg13g2_or2_1 _18296_ (.X(_11474_),
    .B(_11469_),
    .A(_11441_));
 sg13g2_a21oi_1 _18297_ (.A1(_10430_),
    .A2(_11415_),
    .Y(_11475_),
    .B1(_11474_));
 sg13g2_inv_2 _18298_ (.Y(_11476_),
    .A(_11469_));
 sg13g2_nand3_1 _18299_ (.B(_11444_),
    .C(_11476_),
    .A(net661),
    .Y(_11477_));
 sg13g2_o21ai_1 _18300_ (.B1(_11477_),
    .Y(_11478_),
    .A1(net169),
    .A2(_11471_));
 sg13g2_or3_1 _18301_ (.A(_11473_),
    .B(_11475_),
    .C(_11478_),
    .X(_11479_));
 sg13g2_buf_8 _18302_ (.A(_11479_),
    .X(_11480_));
 sg13g2_buf_8 _18303_ (.A(_11480_),
    .X(_11481_));
 sg13g2_nor2_1 _18304_ (.A(_11191_),
    .B(net215),
    .Y(_11482_));
 sg13g2_a21oi_1 _18305_ (.A1(_10523_),
    .A2(_10547_),
    .Y(_11483_),
    .B1(_10324_));
 sg13g2_a221oi_1 _18306_ (.B2(_11017_),
    .C1(_11483_),
    .B1(_11016_),
    .A1(net1072),
    .Y(_11484_),
    .A2(net876));
 sg13g2_buf_1 _18307_ (.A(_11484_),
    .X(_11485_));
 sg13g2_and2_1 _18308_ (.A(_10507_),
    .B(_11485_),
    .X(_11486_));
 sg13g2_buf_1 _18309_ (.A(_11486_),
    .X(_11487_));
 sg13g2_nand2_1 _18310_ (.Y(_11488_),
    .A(_10382_),
    .B(_10417_));
 sg13g2_nor3_1 _18311_ (.A(net287),
    .B(_11361_),
    .C(_11488_),
    .Y(_11489_));
 sg13g2_and3_1 _18312_ (.X(_11490_),
    .A(_11482_),
    .B(_11487_),
    .C(_11489_));
 sg13g2_nand4_1 _18313_ (.B(_11158_),
    .C(net193),
    .A(_10329_),
    .Y(_11491_),
    .D(net216));
 sg13g2_nor2_1 _18314_ (.A(_11474_),
    .B(_11491_),
    .Y(_11492_));
 sg13g2_buf_1 _18315_ (.A(_09367_),
    .X(_11493_));
 sg13g2_buf_1 _18316_ (.A(_11493_),
    .X(_11494_));
 sg13g2_nor2_1 _18317_ (.A(net1120),
    .B(net607),
    .Y(_11495_));
 sg13g2_buf_1 _18318_ (.A(_11495_),
    .X(_11496_));
 sg13g2_o21ai_1 _18319_ (.B1(_11496_),
    .Y(_11497_),
    .A1(_09373_),
    .A2(net694));
 sg13g2_a21oi_1 _18320_ (.A1(_11490_),
    .A2(_11492_),
    .Y(_11498_),
    .B1(_11497_));
 sg13g2_buf_2 _18321_ (.A(_11498_),
    .X(_11499_));
 sg13g2_buf_1 _18322_ (.A(_11499_),
    .X(_11500_));
 sg13g2_o21ai_1 _18323_ (.B1(_11115_),
    .Y(_11501_),
    .A1(_10666_),
    .A2(_10779_));
 sg13g2_buf_1 _18324_ (.A(_11501_),
    .X(_11502_));
 sg13g2_or2_1 _18325_ (.X(_11503_),
    .B(_10987_),
    .A(_10979_));
 sg13g2_buf_1 _18326_ (.A(_11503_),
    .X(_11504_));
 sg13g2_and2_1 _18327_ (.A(_11502_),
    .B(_11504_),
    .X(_11505_));
 sg13g2_buf_1 _18328_ (.A(_11505_),
    .X(_11506_));
 sg13g2_buf_1 _18329_ (.A(_11506_),
    .X(_11507_));
 sg13g2_buf_1 _18330_ (.A(net99),
    .X(_11508_));
 sg13g2_nand2_1 _18331_ (.Y(_11509_),
    .A(_11016_),
    .B(_11017_));
 sg13g2_buf_1 _18332_ (.A(_11509_),
    .X(_11510_));
 sg13g2_nor3_1 _18333_ (.A(_11496_),
    .B(net84),
    .C(net286),
    .Y(_11511_));
 sg13g2_a21oi_1 _18334_ (.A1(_11481_),
    .A2(net85),
    .Y(_11512_),
    .B1(_11511_));
 sg13g2_buf_1 _18335_ (.A(\cpu.ex.r_mult[0] ),
    .X(_11513_));
 sg13g2_a21oi_1 _18336_ (.A1(net1112),
    .A2(_10223_),
    .Y(_11514_),
    .B1(_10234_));
 sg13g2_buf_2 _18337_ (.A(_11514_),
    .X(_11515_));
 sg13g2_nor2_2 _18338_ (.A(_09373_),
    .B(net1120),
    .Y(_11516_));
 sg13g2_nand2_2 _18339_ (.Y(_11517_),
    .A(_09371_),
    .B(_11516_));
 sg13g2_nand2_1 _18340_ (.Y(_11518_),
    .A(_11515_),
    .B(_11517_));
 sg13g2_buf_1 _18341_ (.A(_11518_),
    .X(_11519_));
 sg13g2_nand2_1 _18342_ (.Y(_11520_),
    .A(_11513_),
    .B(_11519_));
 sg13g2_o21ai_1 _18343_ (.B1(_11520_),
    .Y(\cpu.ex.c_mult[0] ),
    .A1(net535),
    .A2(_11512_));
 sg13g2_buf_1 _18344_ (.A(\cpu.dec.load ),
    .X(_11521_));
 sg13g2_nand2_2 _18345_ (.Y(_11522_),
    .A(_08473_),
    .B(net294));
 sg13g2_nor2_1 _18346_ (.A(\cpu.ex.c_div_running ),
    .B(\cpu.ex.c_mult_running ),
    .Y(_11523_));
 sg13g2_buf_1 _18347_ (.A(_00256_),
    .X(_11524_));
 sg13g2_buf_1 _18348_ (.A(net1004),
    .X(_11525_));
 sg13g2_nand2_1 _18349_ (.Y(_11526_),
    .A(net861),
    .B(\cpu.cond[2] ));
 sg13g2_inv_2 _18350_ (.Y(_11527_),
    .A(net1125));
 sg13g2_a21oi_1 _18351_ (.A1(_11524_),
    .A2(_11526_),
    .Y(_11528_),
    .B1(_11527_));
 sg13g2_nor2_1 _18352_ (.A(net861),
    .B(\cpu.dec.jmp ),
    .Y(_11529_));
 sg13g2_nor3_1 _18353_ (.A(net1060),
    .B(_09292_),
    .C(net1036),
    .Y(_11530_));
 sg13g2_o21ai_1 _18354_ (.B1(_11530_),
    .Y(_11531_),
    .A1(_11528_),
    .A2(_11529_));
 sg13g2_a21oi_1 _18355_ (.A1(_10762_),
    .A2(\cpu.dec.r_swapsp ),
    .Y(_11532_),
    .B1(_11531_));
 sg13g2_nor2_1 _18356_ (.A(net899),
    .B(_09377_),
    .Y(_11533_));
 sg13g2_nor2_2 _18357_ (.A(_11516_),
    .B(_11533_),
    .Y(_11534_));
 sg13g2_a21oi_1 _18358_ (.A1(_11523_),
    .A2(_11532_),
    .Y(_11535_),
    .B1(_11534_));
 sg13g2_a21oi_1 _18359_ (.A1(_11522_),
    .A2(_11535_),
    .Y(_11536_),
    .B1(net899));
 sg13g2_buf_1 _18360_ (.A(_11536_),
    .X(_11537_));
 sg13g2_nand2_1 _18361_ (.Y(_11538_),
    .A(_00308_),
    .B(net191));
 sg13g2_a21o_1 _18362_ (.A2(_11535_),
    .A1(_11522_),
    .B1(net899),
    .X(_11539_));
 sg13g2_buf_2 _18363_ (.A(_11539_),
    .X(_11540_));
 sg13g2_nor2_1 _18364_ (.A(net1041),
    .B(_09274_),
    .Y(_11541_));
 sg13g2_nor2_1 _18365_ (.A(_09823_),
    .B(_09815_),
    .Y(_11542_));
 sg13g2_o21ai_1 _18366_ (.B1(_11542_),
    .Y(_11543_),
    .A1(_09824_),
    .A2(_09819_));
 sg13g2_a21oi_2 _18367_ (.B1(_09281_),
    .Y(_11544_),
    .A2(_11543_),
    .A1(_11541_));
 sg13g2_nand2_1 _18368_ (.Y(_11545_),
    .A(_11540_),
    .B(_11544_));
 sg13g2_a21o_1 _18369_ (.A2(_11545_),
    .A1(_11538_),
    .B1(_08576_),
    .X(_11546_));
 sg13g2_o21ai_1 _18370_ (.B1(_11546_),
    .Y(_00054_),
    .A1(_11521_),
    .A2(_11538_));
 sg13g2_nand2_1 _18371_ (.Y(_11547_),
    .A(_11502_),
    .B(_11504_));
 sg13g2_buf_1 _18372_ (.A(_11547_),
    .X(_11548_));
 sg13g2_and2_1 _18373_ (.A(_10549_),
    .B(_10550_),
    .X(_11549_));
 sg13g2_buf_1 _18374_ (.A(_11549_),
    .X(_11550_));
 sg13g2_buf_1 _18375_ (.A(_11550_),
    .X(_11551_));
 sg13g2_nand2_1 _18376_ (.Y(_11552_),
    .A(net115),
    .B(net238));
 sg13g2_buf_1 _18377_ (.A(net693),
    .X(_11553_));
 sg13g2_and2_1 _18378_ (.A(_11513_),
    .B(net606),
    .X(_11554_));
 sg13g2_o21ai_1 _18379_ (.B1(_11554_),
    .Y(_11555_),
    .A1(net99),
    .A2(_10552_));
 sg13g2_o21ai_1 _18380_ (.B1(_11555_),
    .Y(_11556_),
    .A1(_11513_),
    .A2(_11552_));
 sg13g2_nor2_1 _18381_ (.A(net606),
    .B(_11552_),
    .Y(_11557_));
 sg13g2_a221oi_1 _18382_ (.B2(net1120),
    .C1(_11557_),
    .B1(_11556_),
    .A1(_11513_),
    .Y(_11558_),
    .A2(_11499_));
 sg13g2_buf_1 _18383_ (.A(\cpu.ex.r_mult[1] ),
    .X(_11559_));
 sg13g2_nand2_1 _18384_ (.Y(_11560_),
    .A(_11559_),
    .B(net470));
 sg13g2_o21ai_1 _18385_ (.B1(_11560_),
    .Y(\cpu.ex.c_mult[1] ),
    .A1(_10236_),
    .A2(_11558_));
 sg13g2_or2_1 _18386_ (.X(_11561_),
    .B(_10503_),
    .A(_10499_));
 sg13g2_buf_2 _18387_ (.A(_11561_),
    .X(_11562_));
 sg13g2_buf_1 _18388_ (.A(_11562_),
    .X(_11563_));
 sg13g2_and3_1 _18389_ (.X(_11564_),
    .A(_11513_),
    .B(net693),
    .C(_10550_));
 sg13g2_buf_1 _18390_ (.A(_11564_),
    .X(_11565_));
 sg13g2_nand2_1 _18391_ (.Y(_11566_),
    .A(_10549_),
    .B(_11565_));
 sg13g2_xnor2_1 _18392_ (.Y(_11567_),
    .A(net285),
    .B(_11566_));
 sg13g2_nor2_1 _18393_ (.A(net99),
    .B(_11567_),
    .Y(_11568_));
 sg13g2_nand2_1 _18394_ (.Y(_11569_),
    .A(_11559_),
    .B(net606));
 sg13g2_xnor2_1 _18395_ (.Y(_11570_),
    .A(_11568_),
    .B(_11569_));
 sg13g2_a22oi_1 _18396_ (.Y(_11571_),
    .B1(_11570_),
    .B2(_09388_),
    .A2(net85),
    .A1(_11559_));
 sg13g2_inv_1 _18397_ (.Y(_11572_),
    .A(_11571_));
 sg13g2_a22oi_1 _18398_ (.Y(_11573_),
    .B1(_11572_),
    .B2(_11515_),
    .A2(net470),
    .A1(\cpu.ex.r_mult[2] ));
 sg13g2_inv_1 _18399_ (.Y(\cpu.ex.c_mult[2] ),
    .A(_11573_));
 sg13g2_buf_2 _18400_ (.A(_00120_),
    .X(_11574_));
 sg13g2_inv_1 _18401_ (.Y(_11575_),
    .A(_11574_));
 sg13g2_nand3_1 _18402_ (.B(net693),
    .C(_10505_),
    .A(_11559_),
    .Y(_11576_));
 sg13g2_buf_1 _18403_ (.A(_11576_),
    .X(_11577_));
 sg13g2_inv_1 _18404_ (.Y(_11578_),
    .A(_11559_));
 sg13g2_o21ai_1 _18405_ (.B1(_11578_),
    .Y(_11579_),
    .A1(_10499_),
    .A2(_10503_));
 sg13g2_nand3_1 _18406_ (.B(_11565_),
    .C(_11579_),
    .A(_10549_),
    .Y(_11580_));
 sg13g2_buf_1 _18407_ (.A(_11580_),
    .X(_11581_));
 sg13g2_nand2_1 _18408_ (.Y(_11582_),
    .A(_11577_),
    .B(_11581_));
 sg13g2_xnor2_1 _18409_ (.Y(_11583_),
    .A(net240),
    .B(_11582_));
 sg13g2_nor2_1 _18410_ (.A(net99),
    .B(_11583_),
    .Y(_11584_));
 sg13g2_buf_1 _18411_ (.A(_11494_),
    .X(_11585_));
 sg13g2_a22oi_1 _18412_ (.Y(_11586_),
    .B1(_11584_),
    .B2(net530),
    .A2(_11499_),
    .A1(_11575_));
 sg13g2_nor2_1 _18413_ (.A(_11574_),
    .B(net607),
    .Y(_11587_));
 sg13g2_mux2_1 _18414_ (.A0(_11587_),
    .A1(_11574_),
    .S(_11584_),
    .X(_11588_));
 sg13g2_nand2_1 _18415_ (.Y(_11589_),
    .A(net1120),
    .B(_11588_));
 sg13g2_a21oi_1 _18416_ (.A1(_11586_),
    .A2(_11589_),
    .Y(_11590_),
    .B1(_10236_));
 sg13g2_a21o_1 _18417_ (.A2(net470),
    .A1(\cpu.ex.r_mult[3] ),
    .B1(_11590_),
    .X(\cpu.ex.c_mult[3] ));
 sg13g2_buf_1 _18418_ (.A(_00127_),
    .X(_11591_));
 sg13g2_nor2_1 _18419_ (.A(_11591_),
    .B(_09367_),
    .Y(_11592_));
 sg13g2_nand2_1 _18420_ (.Y(_11593_),
    .A(_10464_),
    .B(_10470_));
 sg13g2_buf_1 _18421_ (.A(_11593_),
    .X(_11594_));
 sg13g2_o21ai_1 _18422_ (.B1(net237),
    .Y(_11595_),
    .A1(net285),
    .A2(_11566_));
 sg13g2_a221oi_1 _18423_ (.B2(_11566_),
    .C1(_11578_),
    .B1(net285),
    .A1(_11574_),
    .Y(_11596_),
    .A2(net237));
 sg13g2_a21oi_1 _18424_ (.A1(_11575_),
    .A2(_11595_),
    .Y(_11597_),
    .B1(_11596_));
 sg13g2_nor3_1 _18425_ (.A(_10510_),
    .B(_10512_),
    .C(_11562_),
    .Y(_11598_));
 sg13g2_buf_2 _18426_ (.A(_11598_),
    .X(_11599_));
 sg13g2_nand2b_1 _18427_ (.Y(_11600_),
    .B(_11599_),
    .A_N(_11566_));
 sg13g2_o21ai_1 _18428_ (.B1(_11600_),
    .Y(_11601_),
    .A1(net607),
    .A2(_11597_));
 sg13g2_xnor2_1 _18429_ (.Y(_11602_),
    .A(net287),
    .B(_11601_));
 sg13g2_nor2_1 _18430_ (.A(net99),
    .B(_11602_),
    .Y(_11603_));
 sg13g2_mux2_1 _18431_ (.A0(_11592_),
    .A1(_11591_),
    .S(_11603_),
    .X(_11604_));
 sg13g2_and2_1 _18432_ (.A(net1120),
    .B(_11515_),
    .X(_11605_));
 sg13g2_inv_1 _18433_ (.Y(_11606_),
    .A(_11591_));
 sg13g2_a22oi_1 _18434_ (.Y(_11607_),
    .B1(_11603_),
    .B2(net530),
    .A2(_11500_),
    .A1(_11606_));
 sg13g2_nor2_1 _18435_ (.A(_10236_),
    .B(_11607_),
    .Y(_11608_));
 sg13g2_a221oi_1 _18436_ (.B2(_11605_),
    .C1(_11608_),
    .B1(_11604_),
    .A1(\cpu.ex.r_mult[4] ),
    .Y(_11609_),
    .A2(net470));
 sg13g2_inv_1 _18437_ (.Y(\cpu.ex.c_mult[4] ),
    .A(_11609_));
 sg13g2_buf_1 _18438_ (.A(_00139_),
    .X(_11610_));
 sg13g2_inv_1 _18439_ (.Y(_11611_),
    .A(_11610_));
 sg13g2_nor2_1 _18440_ (.A(_11610_),
    .B(net660),
    .Y(_11612_));
 sg13g2_buf_1 _18441_ (.A(_11612_),
    .X(_11613_));
 sg13g2_buf_1 _18442_ (.A(_11361_),
    .X(_11614_));
 sg13g2_nand3_1 _18443_ (.B(_10464_),
    .C(_10470_),
    .A(net287),
    .Y(_11615_));
 sg13g2_a21oi_2 _18444_ (.B1(_11606_),
    .Y(_11616_),
    .A2(_11325_),
    .A1(_11323_));
 sg13g2_or3_1 _18445_ (.A(_11574_),
    .B(_09367_),
    .C(_11616_),
    .X(_11617_));
 sg13g2_a22oi_1 _18446_ (.Y(_11618_),
    .B1(_11615_),
    .B2(_11617_),
    .A2(_11581_),
    .A1(_11577_));
 sg13g2_buf_1 _18447_ (.A(_11618_),
    .X(_11619_));
 sg13g2_nand3_1 _18448_ (.B(_10470_),
    .C(_11592_),
    .A(_10464_),
    .Y(_11620_));
 sg13g2_a21oi_1 _18449_ (.A1(_11577_),
    .A2(_11581_),
    .Y(_11621_),
    .B1(_11620_));
 sg13g2_nor2_1 _18450_ (.A(_11574_),
    .B(_11616_),
    .Y(_11622_));
 sg13g2_nor3_1 _18451_ (.A(_09367_),
    .B(_10510_),
    .C(_10512_),
    .Y(_11623_));
 sg13g2_and2_1 _18452_ (.A(net287),
    .B(_11592_),
    .X(_11624_));
 sg13g2_a21o_1 _18453_ (.A2(_11623_),
    .A1(_11622_),
    .B1(_11624_),
    .X(_11625_));
 sg13g2_buf_1 _18454_ (.A(_11625_),
    .X(_11626_));
 sg13g2_nor3_1 _18455_ (.A(_11619_),
    .B(_11621_),
    .C(_11626_),
    .Y(_11627_));
 sg13g2_xnor2_1 _18456_ (.Y(_11628_),
    .A(net168),
    .B(_11627_));
 sg13g2_nand2_1 _18457_ (.Y(_11629_),
    .A(net115),
    .B(_11628_));
 sg13g2_xnor2_1 _18458_ (.Y(_11630_),
    .A(_11613_),
    .B(_11629_));
 sg13g2_a22oi_1 _18459_ (.Y(_11631_),
    .B1(_11630_),
    .B2(_09388_),
    .A2(_11499_),
    .A1(_11611_));
 sg13g2_nand2_1 _18460_ (.Y(_11632_),
    .A(\cpu.ex.r_mult[5] ),
    .B(net470));
 sg13g2_o21ai_1 _18461_ (.B1(_11632_),
    .Y(\cpu.ex.c_mult[5] ),
    .A1(_10236_),
    .A2(_11631_));
 sg13g2_or3_1 _18462_ (.A(_11619_),
    .B(_11621_),
    .C(_11626_),
    .X(_11633_));
 sg13g2_nand2_1 _18463_ (.Y(_11634_),
    .A(_11613_),
    .B(_11633_));
 sg13g2_nor4_2 _18464_ (.A(_11613_),
    .B(_11619_),
    .C(_11621_),
    .Y(_11635_),
    .D(_11626_));
 sg13g2_nand2b_1 _18465_ (.Y(_11636_),
    .B(_11361_),
    .A_N(_11635_));
 sg13g2_buf_1 _18466_ (.A(_11636_),
    .X(_11637_));
 sg13g2_and3_1 _18467_ (.X(_11638_),
    .A(net193),
    .B(_11634_),
    .C(_11637_));
 sg13g2_a21oi_1 _18468_ (.A1(_11634_),
    .A2(_11637_),
    .Y(_11639_),
    .B1(net193));
 sg13g2_nor3_1 _18469_ (.A(net99),
    .B(_11638_),
    .C(_11639_),
    .Y(_11640_));
 sg13g2_buf_2 _18470_ (.A(_00151_),
    .X(_11641_));
 sg13g2_nor2_1 _18471_ (.A(_11641_),
    .B(net660),
    .Y(_11642_));
 sg13g2_mux2_1 _18472_ (.A0(_11642_),
    .A1(_11641_),
    .S(_11640_),
    .X(_11643_));
 sg13g2_a22oi_1 _18473_ (.Y(_11644_),
    .B1(_11643_),
    .B2(net1120),
    .A2(_11640_),
    .A1(net530));
 sg13g2_inv_1 _18474_ (.Y(_11645_),
    .A(_11499_));
 sg13g2_nor2_1 _18475_ (.A(_10236_),
    .B(_11645_),
    .Y(_11646_));
 sg13g2_buf_1 _18476_ (.A(_11646_),
    .X(_11647_));
 sg13g2_inv_1 _18477_ (.Y(_11648_),
    .A(_11641_));
 sg13g2_a22oi_1 _18478_ (.Y(_11649_),
    .B1(_11647_),
    .B2(_11648_),
    .A2(net470),
    .A1(\cpu.ex.r_mult[6] ));
 sg13g2_o21ai_1 _18479_ (.B1(_11649_),
    .Y(\cpu.ex.c_mult[6] ),
    .A1(_10237_),
    .A2(_11644_));
 sg13g2_buf_1 _18480_ (.A(_00163_),
    .X(_11650_));
 sg13g2_inv_1 _18481_ (.Y(_11651_),
    .A(_11650_));
 sg13g2_nor2_1 _18482_ (.A(_11650_),
    .B(_09367_),
    .Y(_11652_));
 sg13g2_nand3_1 _18483_ (.B(_11634_),
    .C(_11637_),
    .A(net193),
    .Y(_11653_));
 sg13g2_a21oi_1 _18484_ (.A1(_11653_),
    .A2(_11642_),
    .Y(_11654_),
    .B1(_11639_));
 sg13g2_xnor2_1 _18485_ (.Y(_11655_),
    .A(net216),
    .B(_11654_));
 sg13g2_nor2_1 _18486_ (.A(net84),
    .B(_11655_),
    .Y(_11656_));
 sg13g2_mux2_1 _18487_ (.A0(_11652_),
    .A1(_11650_),
    .S(_11656_),
    .X(_11657_));
 sg13g2_nor3_1 _18488_ (.A(net606),
    .B(net84),
    .C(_11655_),
    .Y(_11658_));
 sg13g2_a221oi_1 _18489_ (.B2(_09383_),
    .C1(_11658_),
    .B1(_11657_),
    .A1(_11651_),
    .Y(_11659_),
    .A2(_11500_));
 sg13g2_buf_1 _18490_ (.A(_11519_),
    .X(_11660_));
 sg13g2_nand2_1 _18491_ (.Y(_11661_),
    .A(\cpu.ex.r_mult[7] ),
    .B(net411));
 sg13g2_o21ai_1 _18492_ (.B1(_11661_),
    .Y(\cpu.ex.c_mult[7] ),
    .A1(_10237_),
    .A2(_11659_));
 sg13g2_nand2_1 _18493_ (.Y(_11662_),
    .A(_09388_),
    .B(_11515_));
 sg13g2_buf_2 _18494_ (.A(_11662_),
    .X(_11663_));
 sg13g2_buf_1 _18495_ (.A(_00164_),
    .X(_11664_));
 sg13g2_nor2_1 _18496_ (.A(_11664_),
    .B(_09367_),
    .Y(_11665_));
 sg13g2_buf_1 _18497_ (.A(_11665_),
    .X(_11666_));
 sg13g2_buf_1 _18498_ (.A(_11158_),
    .X(_11667_));
 sg13g2_nor2_1 _18499_ (.A(_11648_),
    .B(_11651_),
    .Y(_11668_));
 sg13g2_or2_1 _18500_ (.X(_11669_),
    .B(_11668_),
    .A(net660));
 sg13g2_a21o_1 _18501_ (.A2(_11668_),
    .A1(_11610_),
    .B1(net660),
    .X(_11670_));
 sg13g2_nand2b_1 _18502_ (.Y(_11671_),
    .B(net876),
    .A_N(_08829_));
 sg13g2_nand3_1 _18503_ (.B(_11356_),
    .C(_11357_),
    .A(net750),
    .Y(_11672_));
 sg13g2_buf_1 _18504_ (.A(_11672_),
    .X(_11673_));
 sg13g2_nand2_1 _18505_ (.Y(_11674_),
    .A(_11671_),
    .B(_11673_));
 sg13g2_buf_2 _18506_ (.A(_11674_),
    .X(_11675_));
 sg13g2_a221oi_1 _18507_ (.B2(_11675_),
    .C1(_11295_),
    .B1(_11670_),
    .A1(_11393_),
    .Y(_11676_),
    .A2(_11669_));
 sg13g2_buf_1 _18508_ (.A(_11676_),
    .X(_11677_));
 sg13g2_inv_1 _18509_ (.Y(_11678_),
    .A(_11677_));
 sg13g2_or4_1 _18510_ (.A(_11610_),
    .B(_10510_),
    .C(_10512_),
    .D(_11616_),
    .X(_11679_));
 sg13g2_nand2_1 _18511_ (.Y(_11680_),
    .A(_11575_),
    .B(_11611_));
 sg13g2_or2_1 _18512_ (.X(_11681_),
    .B(_11680_),
    .A(_11616_));
 sg13g2_a22oi_1 _18513_ (.Y(_11682_),
    .B1(_11679_),
    .B2(_11681_),
    .A2(_11581_),
    .A1(_11577_));
 sg13g2_nand3_1 _18514_ (.B(_11323_),
    .C(_11325_),
    .A(_11606_),
    .Y(_11683_));
 sg13g2_buf_1 _18515_ (.A(_11683_),
    .X(_11684_));
 sg13g2_nor2_1 _18516_ (.A(_11610_),
    .B(_11684_),
    .Y(_11685_));
 sg13g2_nor4_1 _18517_ (.A(_10510_),
    .B(_10512_),
    .C(_11616_),
    .D(_11680_),
    .Y(_11686_));
 sg13g2_or2_1 _18518_ (.X(_11687_),
    .B(_11686_),
    .A(_11685_));
 sg13g2_or4_1 _18519_ (.A(_11651_),
    .B(net194),
    .C(_11682_),
    .D(_11687_),
    .X(_11688_));
 sg13g2_nor2_1 _18520_ (.A(_11578_),
    .B(_11562_),
    .Y(_11689_));
 sg13g2_o21ai_1 _18521_ (.B1(_11684_),
    .Y(_11690_),
    .A1(_10510_),
    .A2(_10512_));
 sg13g2_nand2_1 _18522_ (.Y(_11691_),
    .A(_11574_),
    .B(_11684_));
 sg13g2_and3_1 _18523_ (.X(_11692_),
    .A(_10549_),
    .B(_11565_),
    .C(_11579_));
 sg13g2_a221oi_1 _18524_ (.B2(_11691_),
    .C1(_11692_),
    .B1(_11690_),
    .A1(net693),
    .Y(_11693_),
    .A2(_11689_));
 sg13g2_nand2_1 _18525_ (.Y(_11694_),
    .A(_11591_),
    .B(_11327_));
 sg13g2_o21ai_1 _18526_ (.B1(_11694_),
    .Y(_11695_),
    .A1(_11575_),
    .A2(_11690_));
 sg13g2_o21ai_1 _18527_ (.B1(_11668_),
    .Y(_11696_),
    .A1(_11693_),
    .A2(_11695_));
 sg13g2_nand4_1 _18528_ (.B(_11688_),
    .C(_11696_),
    .A(_11553_),
    .Y(_11697_),
    .D(_11677_));
 sg13g2_o21ai_1 _18529_ (.B1(_11697_),
    .Y(_11698_),
    .A1(_11637_),
    .A2(_11678_));
 sg13g2_nand2_1 _18530_ (.Y(_11699_),
    .A(_11361_),
    .B(_11652_));
 sg13g2_nand2_1 _18531_ (.Y(_11700_),
    .A(_11613_),
    .B(_11652_));
 sg13g2_a221oi_1 _18532_ (.B2(_11700_),
    .C1(_11627_),
    .B1(_11699_),
    .A1(_11641_),
    .Y(_11701_),
    .A2(net193));
 sg13g2_nor3_1 _18533_ (.A(_11641_),
    .B(_11650_),
    .C(net607),
    .Y(_11702_));
 sg13g2_nor2_1 _18534_ (.A(_11641_),
    .B(_11700_),
    .Y(_11703_));
 sg13g2_nor3_1 _18535_ (.A(net193),
    .B(_11675_),
    .C(_11700_),
    .Y(_11704_));
 sg13g2_a221oi_1 _18536_ (.B2(_11361_),
    .C1(_11704_),
    .B1(_11703_),
    .A1(net194),
    .Y(_11705_),
    .A2(_11702_));
 sg13g2_nand2b_1 _18537_ (.Y(_11706_),
    .B(_11705_),
    .A_N(_11701_));
 sg13g2_nor2_1 _18538_ (.A(_11698_),
    .B(_11706_),
    .Y(_11707_));
 sg13g2_xnor2_1 _18539_ (.Y(_11708_),
    .A(net190),
    .B(_11707_));
 sg13g2_nor2_1 _18540_ (.A(net84),
    .B(_11708_),
    .Y(_11709_));
 sg13g2_xnor2_1 _18541_ (.Y(_11710_),
    .A(_11666_),
    .B(_11709_));
 sg13g2_inv_1 _18542_ (.Y(_11711_),
    .A(_11664_));
 sg13g2_a22oi_1 _18543_ (.Y(_11712_),
    .B1(_11647_),
    .B2(_11711_),
    .A2(net470),
    .A1(\cpu.ex.r_mult[8] ));
 sg13g2_o21ai_1 _18544_ (.B1(_11712_),
    .Y(\cpu.ex.c_mult[8] ),
    .A1(_11663_),
    .A2(_11710_));
 sg13g2_buf_1 _18545_ (.A(_00165_),
    .X(_11713_));
 sg13g2_inv_1 _18546_ (.Y(_11714_),
    .A(_11713_));
 sg13g2_nand2_1 _18547_ (.Y(_11715_),
    .A(_11714_),
    .B(_09386_));
 sg13g2_or2_1 _18548_ (.X(_11716_),
    .B(_11715_),
    .A(_11663_));
 sg13g2_nor2_1 _18549_ (.A(_11496_),
    .B(_10236_),
    .Y(_11717_));
 sg13g2_nand2_1 _18550_ (.Y(_11718_),
    .A(_11717_),
    .B(_11715_));
 sg13g2_buf_1 _18551_ (.A(_11162_),
    .X(_11719_));
 sg13g2_nor2_1 _18552_ (.A(net189),
    .B(_11666_),
    .Y(_11720_));
 sg13g2_nand3_1 _18553_ (.B(_11156_),
    .C(_11666_),
    .A(_11127_),
    .Y(_11721_));
 sg13g2_buf_1 _18554_ (.A(_11721_),
    .X(_11722_));
 sg13g2_o21ai_1 _18555_ (.B1(_11722_),
    .Y(_11723_),
    .A1(_11707_),
    .A2(_11720_));
 sg13g2_xnor2_1 _18556_ (.Y(_11724_),
    .A(net215),
    .B(_11723_));
 sg13g2_nor2_1 _18557_ (.A(_11508_),
    .B(_11724_),
    .Y(_11725_));
 sg13g2_mux2_1 _18558_ (.A0(_11716_),
    .A1(_11718_),
    .S(_11725_),
    .X(_11726_));
 sg13g2_buf_1 _18559_ (.A(_11647_),
    .X(_11727_));
 sg13g2_a22oi_1 _18560_ (.Y(_11728_),
    .B1(net58),
    .B2(_11714_),
    .A2(net411),
    .A1(\cpu.ex.r_mult[9] ));
 sg13g2_nand2_1 _18561_ (.Y(\cpu.ex.c_mult[9] ),
    .A(_11726_),
    .B(_11728_));
 sg13g2_buf_1 _18562_ (.A(_00166_),
    .X(_11729_));
 sg13g2_inv_1 _18563_ (.Y(_11730_),
    .A(_11729_));
 sg13g2_buf_1 _18564_ (.A(_11191_),
    .X(_11731_));
 sg13g2_a21oi_1 _18565_ (.A1(_11613_),
    .A2(_11633_),
    .Y(_11732_),
    .B1(_11361_));
 sg13g2_a21oi_1 _18566_ (.A1(_11197_),
    .A2(_11225_),
    .Y(_11733_),
    .B1(_11715_));
 sg13g2_nand2_1 _18567_ (.Y(_11734_),
    .A(_11664_),
    .B(_11713_));
 sg13g2_a221oi_1 _18568_ (.B2(_11734_),
    .C1(_11370_),
    .B1(net693),
    .A1(_08788_),
    .Y(_11735_),
    .A2(_10326_));
 sg13g2_a21o_1 _18569_ (.A2(_11733_),
    .A1(_11664_),
    .B1(_11735_),
    .X(_11736_));
 sg13g2_nor3_1 _18570_ (.A(_11713_),
    .B(_11368_),
    .C(_11370_),
    .Y(_11737_));
 sg13g2_a21oi_1 _18571_ (.A1(_11197_),
    .A2(_11225_),
    .Y(_11738_),
    .B1(_11714_));
 sg13g2_nor2_1 _18572_ (.A(_11737_),
    .B(_11738_),
    .Y(_11739_));
 sg13g2_and2_1 _18573_ (.A(_11158_),
    .B(_11666_),
    .X(_11740_));
 sg13g2_a22oi_1 _18574_ (.Y(_11741_),
    .B1(_11739_),
    .B2(_11740_),
    .A2(_11736_),
    .A1(net189));
 sg13g2_mux2_1 _18575_ (.A0(_11650_),
    .A1(_11652_),
    .S(_11292_),
    .X(_11742_));
 sg13g2_a22oi_1 _18576_ (.Y(_11743_),
    .B1(_11742_),
    .B2(_11641_),
    .A2(net239),
    .A1(net660));
 sg13g2_nand2_1 _18577_ (.Y(_11744_),
    .A(_11651_),
    .B(_11300_));
 sg13g2_nand3_1 _18578_ (.B(_11288_),
    .C(_11290_),
    .A(_11650_),
    .Y(_11745_));
 sg13g2_buf_1 _18579_ (.A(_11745_),
    .X(_11746_));
 sg13g2_nand3_1 _18580_ (.B(_11744_),
    .C(_11746_),
    .A(_11642_),
    .Y(_11747_));
 sg13g2_mux2_1 _18581_ (.A0(_11743_),
    .A1(_11747_),
    .S(_11262_),
    .X(_11748_));
 sg13g2_or4_1 _18582_ (.A(_11635_),
    .B(_11732_),
    .C(_11741_),
    .D(_11748_),
    .X(_11749_));
 sg13g2_buf_1 _18583_ (.A(_11749_),
    .X(_11750_));
 sg13g2_nand3_1 _18584_ (.B(_11234_),
    .C(_11260_),
    .A(_11648_),
    .Y(_11751_));
 sg13g2_nand3_1 _18585_ (.B(_11156_),
    .C(_11746_),
    .A(_11127_),
    .Y(_11752_));
 sg13g2_nand2_1 _18586_ (.Y(_11753_),
    .A(_11711_),
    .B(_11746_));
 sg13g2_a221oi_1 _18587_ (.B2(_11753_),
    .C1(_11738_),
    .B1(_11752_),
    .A1(_11744_),
    .Y(_11754_),
    .A2(_11751_));
 sg13g2_nor3_1 _18588_ (.A(_11664_),
    .B(_11158_),
    .C(_11738_),
    .Y(_11755_));
 sg13g2_nor3_1 _18589_ (.A(_11737_),
    .B(_11754_),
    .C(_11755_),
    .Y(_11756_));
 sg13g2_or2_1 _18590_ (.X(_11757_),
    .B(_11756_),
    .A(net607));
 sg13g2_buf_1 _18591_ (.A(_11757_),
    .X(_11758_));
 sg13g2_nand2_1 _18592_ (.Y(_11759_),
    .A(_11750_),
    .B(_11758_));
 sg13g2_xnor2_1 _18593_ (.Y(_11760_),
    .A(net188),
    .B(_11759_));
 sg13g2_nor2_1 _18594_ (.A(net84),
    .B(_11760_),
    .Y(_11761_));
 sg13g2_nor2_1 _18595_ (.A(_11729_),
    .B(net660),
    .Y(_11762_));
 sg13g2_xor2_1 _18596_ (.B(_11762_),
    .A(_11761_),
    .X(_11763_));
 sg13g2_a22oi_1 _18597_ (.Y(_11764_),
    .B1(_11763_),
    .B2(_09388_),
    .A2(net85),
    .A1(_11730_));
 sg13g2_nand2_1 _18598_ (.Y(_11765_),
    .A(\cpu.ex.r_mult[10] ),
    .B(net411));
 sg13g2_o21ai_1 _18599_ (.B1(_11765_),
    .Y(\cpu.ex.c_mult[10] ),
    .A1(net535),
    .A2(_11764_));
 sg13g2_inv_1 _18600_ (.Y(_11766_),
    .A(_00167_));
 sg13g2_buf_1 _18601_ (.A(_10417_),
    .X(_11767_));
 sg13g2_nor2_1 _18602_ (.A(_11729_),
    .B(_11715_),
    .Y(_11768_));
 sg13g2_o21ai_1 _18603_ (.B1(_11768_),
    .Y(_11769_),
    .A1(net99),
    .A2(_11482_));
 sg13g2_nor2_1 _18604_ (.A(_11730_),
    .B(net214),
    .Y(_11770_));
 sg13g2_nand3_1 _18605_ (.B(_11166_),
    .C(_11189_),
    .A(net607),
    .Y(_11771_));
 sg13g2_nand3_1 _18606_ (.B(_11730_),
    .C(net693),
    .A(_11713_),
    .Y(_11772_));
 sg13g2_a21o_1 _18607_ (.A2(_11189_),
    .A1(_11166_),
    .B1(_11772_),
    .X(_11773_));
 sg13g2_nand4_1 _18608_ (.B(_11729_),
    .C(_11166_),
    .A(_11713_),
    .Y(_11774_),
    .D(_11189_));
 sg13g2_nand3_1 _18609_ (.B(_11773_),
    .C(_11774_),
    .A(_11771_),
    .Y(_11775_));
 sg13g2_a22oi_1 _18610_ (.Y(_11776_),
    .B1(_11775_),
    .B2(net215),
    .A2(_11770_),
    .A1(_11733_));
 sg13g2_nand2_1 _18611_ (.Y(_11777_),
    .A(_11769_),
    .B(_11776_));
 sg13g2_nor2_1 _18612_ (.A(_11729_),
    .B(_11376_),
    .Y(_11778_));
 sg13g2_a21oi_1 _18613_ (.A1(_11166_),
    .A2(_11189_),
    .Y(_11779_),
    .B1(_11730_));
 sg13g2_nor4_1 _18614_ (.A(_11713_),
    .B(_11368_),
    .C(_11370_),
    .D(_11779_),
    .Y(_11780_));
 sg13g2_nor2_1 _18615_ (.A(_11778_),
    .B(_11780_),
    .Y(_11781_));
 sg13g2_nor2_1 _18616_ (.A(net530),
    .B(_11781_),
    .Y(_11782_));
 sg13g2_a21oi_1 _18617_ (.A1(_11723_),
    .A2(_11777_),
    .Y(_11783_),
    .B1(_11782_));
 sg13g2_xnor2_1 _18618_ (.Y(_11784_),
    .A(net211),
    .B(_11783_));
 sg13g2_nor2_1 _18619_ (.A(_11508_),
    .B(_11784_),
    .Y(_11785_));
 sg13g2_nand2_1 _18620_ (.Y(_11786_),
    .A(_11766_),
    .B(_11553_));
 sg13g2_xnor2_1 _18621_ (.Y(_11787_),
    .A(_11785_),
    .B(_11786_));
 sg13g2_a22oi_1 _18622_ (.Y(_11788_),
    .B1(_11787_),
    .B2(_09388_),
    .A2(net85),
    .A1(_11766_));
 sg13g2_nand2_1 _18623_ (.Y(_11789_),
    .A(\cpu.ex.r_mult[11] ),
    .B(_11660_));
 sg13g2_o21ai_1 _18624_ (.B1(_11789_),
    .Y(\cpu.ex.c_mult[11] ),
    .A1(net535),
    .A2(_11788_));
 sg13g2_nor2_1 _18625_ (.A(_00167_),
    .B(net660),
    .Y(_11790_));
 sg13g2_buf_2 _18626_ (.A(_11790_),
    .X(_11791_));
 sg13g2_o21ai_1 _18627_ (.B1(net214),
    .Y(_11792_),
    .A1(net217),
    .A2(_11722_));
 sg13g2_a221oi_1 _18628_ (.B2(_11722_),
    .C1(_11713_),
    .B1(net217),
    .A1(_11729_),
    .Y(_11793_),
    .A2(_11376_));
 sg13g2_a21oi_1 _18629_ (.A1(_11730_),
    .A2(_11792_),
    .Y(_11794_),
    .B1(_11793_));
 sg13g2_and2_1 _18630_ (.A(net189),
    .B(_11666_),
    .X(_11795_));
 sg13g2_nand3_1 _18631_ (.B(net215),
    .C(_11795_),
    .A(net188),
    .Y(_11796_));
 sg13g2_o21ai_1 _18632_ (.B1(_11796_),
    .Y(_11797_),
    .A1(net607),
    .A2(_11794_));
 sg13g2_nor2_1 _18633_ (.A(_11791_),
    .B(_11797_),
    .Y(_11798_));
 sg13g2_a21oi_1 _18634_ (.A1(_11791_),
    .A2(_11797_),
    .Y(_11799_),
    .B1(net212));
 sg13g2_xnor2_1 _18635_ (.Y(_11800_),
    .A(_11410_),
    .B(_11791_));
 sg13g2_xnor2_1 _18636_ (.Y(_11801_),
    .A(_11195_),
    .B(_11762_));
 sg13g2_nand2b_1 _18637_ (.Y(_11802_),
    .B(_11801_),
    .A_N(_11800_));
 sg13g2_nor2_1 _18638_ (.A(_11741_),
    .B(_11802_),
    .Y(_11803_));
 sg13g2_o21ai_1 _18639_ (.B1(_11803_),
    .Y(_11804_),
    .A1(_11698_),
    .A2(_11706_));
 sg13g2_o21ai_1 _18640_ (.B1(_11804_),
    .Y(_11805_),
    .A1(_11798_),
    .A2(_11799_));
 sg13g2_xnor2_1 _18641_ (.Y(_11806_),
    .A(net213),
    .B(_11805_));
 sg13g2_nand2_1 _18642_ (.Y(_11807_),
    .A(net115),
    .B(_11806_));
 sg13g2_inv_1 _18643_ (.Y(_11808_),
    .A(_00168_));
 sg13g2_nand2_1 _18644_ (.Y(_11809_),
    .A(_11808_),
    .B(_09386_));
 sg13g2_xnor2_1 _18645_ (.Y(_11810_),
    .A(_11807_),
    .B(_11809_));
 sg13g2_a22oi_1 _18646_ (.Y(_11811_),
    .B1(net58),
    .B2(_11808_),
    .A2(net411),
    .A1(\cpu.ex.r_mult[12] ));
 sg13g2_o21ai_1 _18647_ (.B1(_11811_),
    .Y(\cpu.ex.c_mult[12] ),
    .A1(_11663_),
    .A2(_11810_));
 sg13g2_nor2_1 _18648_ (.A(_11675_),
    .B(_11635_),
    .Y(_11812_));
 sg13g2_and3_1 _18649_ (.X(_11813_),
    .A(net606),
    .B(_11688_),
    .C(_11677_));
 sg13g2_a22oi_1 _18650_ (.Y(_11814_),
    .B1(_11813_),
    .B2(_11696_),
    .A2(_11677_),
    .A1(_11812_));
 sg13g2_nor2b_1 _18651_ (.A(_11701_),
    .B_N(_11705_),
    .Y(_11815_));
 sg13g2_nor2_1 _18652_ (.A(_00168_),
    .B(net660),
    .Y(_11816_));
 sg13g2_xnor2_1 _18653_ (.Y(_11817_),
    .A(_10382_),
    .B(_11816_));
 sg13g2_nand3_1 _18654_ (.B(_11227_),
    .C(_11768_),
    .A(net214),
    .Y(_11818_));
 sg13g2_a21oi_1 _18655_ (.A1(_11776_),
    .A2(_11818_),
    .Y(_11819_),
    .B1(_11800_));
 sg13g2_nand4_1 _18656_ (.B(_11666_),
    .C(_11817_),
    .A(net115),
    .Y(_11820_),
    .D(_11819_));
 sg13g2_nand4_1 _18657_ (.B(net189),
    .C(_11817_),
    .A(net115),
    .Y(_11821_),
    .D(_11819_));
 sg13g2_a22oi_1 _18658_ (.Y(_11822_),
    .B1(_11820_),
    .B2(_11821_),
    .A2(_11815_),
    .A1(_11814_));
 sg13g2_o21ai_1 _18659_ (.B1(net606),
    .Y(_11823_),
    .A1(_11778_),
    .A2(_11780_));
 sg13g2_o21ai_1 _18660_ (.B1(_11823_),
    .Y(_11824_),
    .A1(_11767_),
    .A2(_11786_));
 sg13g2_nor2_1 _18661_ (.A(_11410_),
    .B(_11791_),
    .Y(_11825_));
 sg13g2_a21oi_1 _18662_ (.A1(_11400_),
    .A2(_11809_),
    .Y(_11826_),
    .B1(_11825_));
 sg13g2_a22oi_1 _18663_ (.Y(_11827_),
    .B1(_11824_),
    .B2(_11826_),
    .A2(_11816_),
    .A1(_10383_));
 sg13g2_nand4_1 _18664_ (.B(_11795_),
    .C(_11817_),
    .A(_11548_),
    .Y(_11828_),
    .D(_11819_));
 sg13g2_o21ai_1 _18665_ (.B1(_11828_),
    .Y(_11829_),
    .A1(net99),
    .A2(_11827_));
 sg13g2_nor2_1 _18666_ (.A(_11822_),
    .B(_11829_),
    .Y(_11830_));
 sg13g2_buf_1 _18667_ (.A(_00169_),
    .X(_11831_));
 sg13g2_nor2_2 _18668_ (.A(_11831_),
    .B(_11493_),
    .Y(_11832_));
 sg13g2_buf_1 _18669_ (.A(net170),
    .X(_11833_));
 sg13g2_nor2_1 _18670_ (.A(net84),
    .B(net141),
    .Y(_11834_));
 sg13g2_xnor2_1 _18671_ (.Y(_11835_),
    .A(_11832_),
    .B(_11834_));
 sg13g2_xor2_1 _18672_ (.B(_11835_),
    .A(_11830_),
    .X(_11836_));
 sg13g2_nand2_1 _18673_ (.Y(_11837_),
    .A(_11717_),
    .B(_11836_));
 sg13g2_inv_1 _18674_ (.Y(_11838_),
    .A(_11831_));
 sg13g2_a22oi_1 _18675_ (.Y(_11839_),
    .B1(_11647_),
    .B2(_11838_),
    .A2(net470),
    .A1(\cpu.ex.r_mult[13] ));
 sg13g2_and2_1 _18676_ (.A(_11837_),
    .B(_11839_),
    .X(_11840_));
 sg13g2_inv_1 _18677_ (.Y(\cpu.ex.c_mult[13] ),
    .A(_11840_));
 sg13g2_xor2_1 _18678_ (.B(_11832_),
    .A(_10329_),
    .X(_11841_));
 sg13g2_nor2_1 _18679_ (.A(_11802_),
    .B(_11841_),
    .Y(_11842_));
 sg13g2_nand3_1 _18680_ (.B(_11817_),
    .C(_11842_),
    .A(net115),
    .Y(_11843_));
 sg13g2_a21oi_1 _18681_ (.A1(_11750_),
    .A2(_11758_),
    .Y(_11844_),
    .B1(_11843_));
 sg13g2_a22oi_1 _18682_ (.Y(_11845_),
    .B1(_11191_),
    .B2(_11730_),
    .A2(_11410_),
    .A1(_11766_));
 sg13g2_o21ai_1 _18683_ (.B1(_11816_),
    .Y(_11846_),
    .A1(_11766_),
    .A2(net212));
 sg13g2_o21ai_1 _18684_ (.B1(_10382_),
    .Y(_11847_),
    .A1(_11845_),
    .A2(_11846_));
 sg13g2_a22oi_1 _18685_ (.Y(_11848_),
    .B1(_11791_),
    .B2(net212),
    .A2(_11762_),
    .A1(_11191_));
 sg13g2_o21ai_1 _18686_ (.B1(_11809_),
    .Y(_11849_),
    .A1(_11825_),
    .A2(_11848_));
 sg13g2_nor2b_1 _18687_ (.A(_10329_),
    .B_N(_11832_),
    .Y(_11850_));
 sg13g2_a21oi_1 _18688_ (.A1(_11847_),
    .A2(_11849_),
    .Y(_11851_),
    .B1(_11850_));
 sg13g2_nor2b_1 _18689_ (.A(_11832_),
    .B_N(_10329_),
    .Y(_11852_));
 sg13g2_or3_1 _18690_ (.A(_11506_),
    .B(_11851_),
    .C(_11852_),
    .X(_11853_));
 sg13g2_nand2b_1 _18691_ (.Y(_11854_),
    .B(_11853_),
    .A_N(_11844_));
 sg13g2_nor2_2 _18692_ (.A(_00170_),
    .B(net607),
    .Y(_11855_));
 sg13g2_a21oi_1 _18693_ (.A1(_11502_),
    .A2(_11504_),
    .Y(_11856_),
    .B1(_11476_));
 sg13g2_xnor2_1 _18694_ (.Y(_11857_),
    .A(_11855_),
    .B(_11856_));
 sg13g2_xor2_1 _18695_ (.B(_11857_),
    .A(_11854_),
    .X(_11858_));
 sg13g2_inv_1 _18696_ (.Y(_11859_),
    .A(_00170_));
 sg13g2_a22oi_1 _18697_ (.Y(_11860_),
    .B1(net58),
    .B2(_11859_),
    .A2(net411),
    .A1(\cpu.ex.r_mult[14] ));
 sg13g2_o21ai_1 _18698_ (.B1(_11860_),
    .Y(\cpu.ex.c_mult[14] ),
    .A1(_11663_),
    .A2(_11858_));
 sg13g2_buf_1 _18699_ (.A(\cpu.ex.r_mult[15] ),
    .X(_11861_));
 sg13g2_and2_1 _18700_ (.A(_11469_),
    .B(_11855_),
    .X(_11862_));
 sg13g2_buf_1 _18701_ (.A(_11862_),
    .X(_11863_));
 sg13g2_nor2_1 _18702_ (.A(_11469_),
    .B(_11855_),
    .Y(_11864_));
 sg13g2_nor4_1 _18703_ (.A(_11831_),
    .B(_11585_),
    .C(net141),
    .D(_11864_),
    .Y(_11865_));
 sg13g2_o21ai_1 _18704_ (.B1(net115),
    .Y(_11866_),
    .A1(_11863_),
    .A2(_11865_));
 sg13g2_nor4_1 _18705_ (.A(_11831_),
    .B(_11585_),
    .C(_11507_),
    .D(_11864_),
    .Y(_11867_));
 sg13g2_o21ai_1 _18706_ (.B1(_11867_),
    .Y(_11868_),
    .A1(_11822_),
    .A2(_11829_));
 sg13g2_nor3_1 _18707_ (.A(net84),
    .B(net141),
    .C(_11864_),
    .Y(_11869_));
 sg13g2_o21ai_1 _18708_ (.B1(_11869_),
    .Y(_11870_),
    .A1(_11822_),
    .A2(_11829_));
 sg13g2_nand3_1 _18709_ (.B(_11868_),
    .C(_11870_),
    .A(_11866_),
    .Y(_11871_));
 sg13g2_inv_1 _18710_ (.Y(_11872_),
    .A(_11441_));
 sg13g2_a21oi_1 _18711_ (.A1(_11502_),
    .A2(_11504_),
    .Y(_11873_),
    .B1(_11872_));
 sg13g2_nor2_1 _18712_ (.A(_00171_),
    .B(_11494_),
    .Y(_11874_));
 sg13g2_xnor2_1 _18713_ (.Y(_11875_),
    .A(_11873_),
    .B(_11874_));
 sg13g2_xnor2_1 _18714_ (.Y(_11876_),
    .A(_11871_),
    .B(_11875_));
 sg13g2_nand2_1 _18715_ (.Y(_11877_),
    .A(_09388_),
    .B(_11876_));
 sg13g2_o21ai_1 _18716_ (.B1(_11877_),
    .Y(_11878_),
    .A1(_00171_),
    .A2(_11645_));
 sg13g2_a22oi_1 _18717_ (.Y(_11879_),
    .B1(_11878_),
    .B2(_11515_),
    .A2(net411),
    .A1(_11861_));
 sg13g2_inv_1 _18718_ (.Y(\cpu.ex.c_mult[15] ),
    .A(_11879_));
 sg13g2_inv_1 _18719_ (.Y(_00000_),
    .A(net2));
 sg13g2_inv_1 _18720_ (.Y(_11880_),
    .A(\cpu.qspi.r_state[11] ));
 sg13g2_nor2_1 _18721_ (.A(_11880_),
    .B(net631),
    .Y(_00004_));
 sg13g2_inv_1 _18722_ (.Y(_11881_),
    .A(_09851_));
 sg13g2_nor3_1 _18723_ (.A(_11881_),
    .B(net629),
    .C(net142),
    .Y(_00008_));
 sg13g2_buf_1 _18724_ (.A(\cpu.qspi.r_state[10] ),
    .X(_11882_));
 sg13g2_inv_1 _18725_ (.Y(_11883_),
    .A(_11882_));
 sg13g2_nor2_1 _18726_ (.A(_11883_),
    .B(net631),
    .Y(_00003_));
 sg13g2_buf_1 _18727_ (.A(\cpu.qspi.r_state[15] ),
    .X(_11884_));
 sg13g2_buf_1 _18728_ (.A(net764),
    .X(_11885_));
 sg13g2_and2_1 _18729_ (.A(_11884_),
    .B(_11885_),
    .X(_00002_));
 sg13g2_and3_1 _18730_ (.X(_00001_),
    .A(net1118),
    .B(net659),
    .C(_09842_));
 sg13g2_and2_1 _18731_ (.A(_10859_),
    .B(_10885_),
    .X(_11886_));
 sg13g2_buf_1 _18732_ (.A(_11886_),
    .X(_11887_));
 sg13g2_nor4_1 _18733_ (.A(_11061_),
    .B(_10701_),
    .C(_10730_),
    .D(_11887_),
    .Y(_11888_));
 sg13g2_mux2_1 _18734_ (.A0(_09206_),
    .A1(_10806_),
    .S(net532),
    .X(_11889_));
 sg13g2_nand2_1 _18735_ (.Y(_11890_),
    .A(_10890_),
    .B(_10911_));
 sg13g2_o21ai_1 _18736_ (.B1(_10973_),
    .Y(_11891_),
    .A1(net1042),
    .A2(net532));
 sg13g2_nand2_1 _18737_ (.Y(_11892_),
    .A(_11890_),
    .B(_11891_));
 sg13g2_nor3_1 _18738_ (.A(_11084_),
    .B(_11889_),
    .C(_11892_),
    .Y(_11893_));
 sg13g2_nand2_1 _18739_ (.Y(_11894_),
    .A(_11888_),
    .B(_11893_));
 sg13g2_buf_1 _18740_ (.A(net678),
    .X(_11895_));
 sg13g2_nand2b_1 _18741_ (.Y(_11896_),
    .B(_10748_),
    .A_N(net605));
 sg13g2_o21ai_1 _18742_ (.B1(_11896_),
    .Y(_11897_),
    .A1(_10748_),
    .A2(_10832_));
 sg13g2_nor2_1 _18743_ (.A(_10658_),
    .B(_10660_),
    .Y(_11898_));
 sg13g2_nand2_1 _18744_ (.Y(_11899_),
    .A(_10918_),
    .B(_10926_));
 sg13g2_mux2_1 _18745_ (.A0(net614),
    .A1(_11899_),
    .S(net532),
    .X(_11900_));
 sg13g2_nor2_1 _18746_ (.A(_11898_),
    .B(_11900_),
    .Y(_11901_));
 sg13g2_nor3_1 _18747_ (.A(_11044_),
    .B(_11106_),
    .C(_10774_),
    .Y(_11902_));
 sg13g2_nand4_1 _18748_ (.B(_11897_),
    .C(_11901_),
    .A(_10858_),
    .Y(_11903_),
    .D(_11902_));
 sg13g2_nor2_1 _18749_ (.A(_11894_),
    .B(_11903_),
    .Y(_11904_));
 sg13g2_buf_1 _18750_ (.A(_08588_),
    .X(_11905_));
 sg13g2_o21ai_1 _18751_ (.B1(_10951_),
    .Y(_11906_),
    .A1(net860),
    .A2(net532));
 sg13g2_o21ai_1 _18752_ (.B1(_11906_),
    .Y(_11907_),
    .A1(\cpu.cond[1] ),
    .A2(_11904_));
 sg13g2_xnor2_1 _18753_ (.Y(_11908_),
    .A(_11527_),
    .B(_11907_));
 sg13g2_buf_1 _18754_ (.A(_10579_),
    .X(_11909_));
 sg13g2_a21oi_1 _18755_ (.A1(_00271_),
    .A2(_11908_),
    .Y(_11910_),
    .B1(_11909_));
 sg13g2_nor2_1 _18756_ (.A(\cpu.dec.jmp ),
    .B(_11910_),
    .Y(_11911_));
 sg13g2_nor2_1 _18757_ (.A(_09293_),
    .B(net1036),
    .Y(_11912_));
 sg13g2_buf_1 _18758_ (.A(_11912_),
    .X(_11913_));
 sg13g2_nor2b_1 _18759_ (.A(_11911_),
    .B_N(net658),
    .Y(_00053_));
 sg13g2_nor4_1 _18760_ (.A(_09870_),
    .B(net618),
    .C(_09830_),
    .D(_09869_),
    .Y(_00007_));
 sg13g2_buf_1 _18761_ (.A(\cpu.qspi.r_state[3] ),
    .X(_11914_));
 sg13g2_inv_1 _18762_ (.Y(_11915_),
    .A(_11914_));
 sg13g2_nor2_1 _18763_ (.A(_11915_),
    .B(net631),
    .Y(_00009_));
 sg13g2_buf_2 _18764_ (.A(\cpu.qspi.r_state[6] ),
    .X(_11916_));
 sg13g2_and2_1 _18765_ (.A(_11916_),
    .B(net659),
    .X(_00010_));
 sg13g2_and3_1 _18766_ (.X(_00005_),
    .A(_09901_),
    .B(_09878_),
    .C(_09842_));
 sg13g2_buf_2 _18767_ (.A(\cpu.qspi.r_state[13] ),
    .X(_11917_));
 sg13g2_and2_1 _18768_ (.A(_11917_),
    .B(net659),
    .X(_00006_));
 sg13g2_and2_1 _18769_ (.A(_09104_),
    .B(_11885_),
    .X(_00052_));
 sg13g2_or2_1 _18770_ (.X(_11918_),
    .B(net1122),
    .A(_09331_));
 sg13g2_buf_1 _18771_ (.A(_11918_),
    .X(_11919_));
 sg13g2_nor3_1 _18772_ (.A(_09285_),
    .B(net1121),
    .C(_11919_),
    .Y(_11920_));
 sg13g2_a21oi_1 _18773_ (.A1(net419),
    .A2(_11919_),
    .Y(_11921_),
    .B1(_11920_));
 sg13g2_nand2_1 _18774_ (.Y(_11922_),
    .A(_09295_),
    .B(_11921_));
 sg13g2_inv_1 _18775_ (.Y(_11923_),
    .A(_00224_));
 sg13g2_nor3_2 _18776_ (.A(net1122),
    .B(net1121),
    .C(_11923_),
    .Y(_11924_));
 sg13g2_buf_1 _18777_ (.A(net1030),
    .X(_11925_));
 sg13g2_buf_1 _18778_ (.A(net858),
    .X(_11926_));
 sg13g2_buf_1 _18779_ (.A(net894),
    .X(_11927_));
 sg13g2_inv_1 _18780_ (.Y(_11928_),
    .A(_00280_));
 sg13g2_nand2_1 _18781_ (.Y(_11929_),
    .A(net894),
    .B(_00281_));
 sg13g2_o21ai_1 _18782_ (.B1(_11929_),
    .Y(_11930_),
    .A1(net734),
    .A2(_11928_));
 sg13g2_buf_1 _18783_ (.A(net893),
    .X(_11931_));
 sg13g2_buf_1 _18784_ (.A(\cpu.spi.r_src[2] ),
    .X(_11932_));
 sg13g2_nand3_1 _18785_ (.B(net733),
    .C(_11932_),
    .A(net858),
    .Y(_11933_));
 sg13g2_o21ai_1 _18786_ (.B1(_11933_),
    .Y(_11934_),
    .A1(net735),
    .A2(_11930_));
 sg13g2_and2_1 _18787_ (.A(_11924_),
    .B(_11934_),
    .X(_11935_));
 sg13g2_buf_1 _18788_ (.A(net735),
    .X(_11936_));
 sg13g2_buf_1 _18789_ (.A(net734),
    .X(_11937_));
 sg13g2_buf_1 _18790_ (.A(\cpu.spi.r_mode[2][1] ),
    .X(_11938_));
 sg13g2_buf_1 _18791_ (.A(\cpu.spi.r_mode[0][1] ),
    .X(_11939_));
 sg13g2_nand2b_1 _18792_ (.Y(_11940_),
    .B(_11937_),
    .A_N(_11939_));
 sg13g2_o21ai_1 _18793_ (.B1(_11940_),
    .Y(_11941_),
    .A1(net656),
    .A2(_11938_));
 sg13g2_buf_1 _18794_ (.A(\cpu.spi.r_mode[1][1] ),
    .X(_11942_));
 sg13g2_buf_1 _18795_ (.A(net734),
    .X(_11943_));
 sg13g2_mux2_1 _18796_ (.A0(_11939_),
    .A1(_11942_),
    .S(_11943_),
    .X(_11944_));
 sg13g2_nor2_1 _18797_ (.A(net657),
    .B(_11944_),
    .Y(_11945_));
 sg13g2_a21oi_1 _18798_ (.A1(net657),
    .A2(_11941_),
    .Y(_11946_),
    .B1(_11945_));
 sg13g2_buf_1 _18799_ (.A(\cpu.spi.r_sel[1] ),
    .X(_11947_));
 sg13g2_buf_1 _18800_ (.A(_11947_),
    .X(_11948_));
 sg13g2_buf_1 _18801_ (.A(net1002),
    .X(_11949_));
 sg13g2_buf_1 _18802_ (.A(\cpu.spi.r_sel[0] ),
    .X(_11950_));
 sg13g2_inv_1 _18803_ (.Y(_11951_),
    .A(_11950_));
 sg13g2_mux2_1 _18804_ (.A0(_11928_),
    .A1(_11932_),
    .S(_11951_),
    .X(_11952_));
 sg13g2_buf_1 _18805_ (.A(_11950_),
    .X(_11953_));
 sg13g2_buf_1 _18806_ (.A(net1001),
    .X(_11954_));
 sg13g2_buf_1 _18807_ (.A(net1001),
    .X(_11955_));
 sg13g2_nand2_1 _18808_ (.Y(_11956_),
    .A(net855),
    .B(_00281_));
 sg13g2_o21ai_1 _18809_ (.B1(_11956_),
    .Y(_11957_),
    .A1(_11954_),
    .A2(_11928_));
 sg13g2_nor2_1 _18810_ (.A(net1002),
    .B(_11957_),
    .Y(_11958_));
 sg13g2_a21oi_2 _18811_ (.B1(_11958_),
    .Y(_11959_),
    .A2(_11952_),
    .A1(net857));
 sg13g2_nor2_1 _18812_ (.A(_11924_),
    .B(_11959_),
    .Y(_11960_));
 sg13g2_nor2_1 _18813_ (.A(net1038),
    .B(_09347_),
    .Y(_11961_));
 sg13g2_inv_1 _18814_ (.Y(_11962_),
    .A(_11947_));
 sg13g2_buf_1 _18815_ (.A(net855),
    .X(_11963_));
 sg13g2_mux2_1 _18816_ (.A0(_11939_),
    .A1(_11942_),
    .S(net732),
    .X(_11964_));
 sg13g2_nor2_1 _18817_ (.A(_11962_),
    .B(_11950_),
    .Y(_11965_));
 sg13g2_a22oi_1 _18818_ (.Y(_11966_),
    .B1(_11965_),
    .B2(_11938_),
    .A2(_11964_),
    .A1(_11962_));
 sg13g2_xnor2_1 _18819_ (.Y(_11967_),
    .A(_11961_),
    .B(_11966_));
 sg13g2_a22oi_1 _18820_ (.Y(_11968_),
    .B1(_11960_),
    .B2(_11967_),
    .A2(_11946_),
    .A1(_11935_));
 sg13g2_nor2_1 _18821_ (.A(_11935_),
    .B(_11960_),
    .Y(_11969_));
 sg13g2_buf_1 _18822_ (.A(\cpu.gpio.genblk1[3].srcs_o[5] ),
    .X(_11970_));
 sg13g2_o21ai_1 _18823_ (.B1(_11970_),
    .Y(_11971_),
    .A1(_11922_),
    .A2(_11969_));
 sg13g2_o21ai_1 _18824_ (.B1(_11971_),
    .Y(_00316_),
    .A1(_11922_),
    .A2(_11968_));
 sg13g2_nor2b_1 _18825_ (.A(_11922_),
    .B_N(_11969_),
    .Y(_11972_));
 sg13g2_or3_1 _18826_ (.A(net1122),
    .B(net1121),
    .C(_11923_),
    .X(_11973_));
 sg13g2_buf_1 _18827_ (.A(_11973_),
    .X(_11974_));
 sg13g2_and2_1 _18828_ (.A(_11924_),
    .B(_11946_),
    .X(_11975_));
 sg13g2_a21oi_1 _18829_ (.A1(_11974_),
    .A2(_11967_),
    .Y(_11976_),
    .B1(_11975_));
 sg13g2_buf_1 _18830_ (.A(\cpu.gpio.genblk1[3].srcs_o[4] ),
    .X(_11977_));
 sg13g2_nor2_1 _18831_ (.A(_11977_),
    .B(_11972_),
    .Y(_11978_));
 sg13g2_a21oi_1 _18832_ (.A1(_11972_),
    .A2(_11976_),
    .Y(_00317_),
    .B1(_11978_));
 sg13g2_buf_1 _18833_ (.A(\cpu.gpio.genblk1[3].srcs_o[3] ),
    .X(_11979_));
 sg13g2_mux2_1 _18834_ (.A0(\cpu.spi.r_out[7] ),
    .A1(_10103_),
    .S(net897),
    .X(_11980_));
 sg13g2_nor2_1 _18835_ (.A(net899),
    .B(_09265_),
    .Y(_11981_));
 sg13g2_inv_1 _18836_ (.Y(_11982_),
    .A(_00222_));
 sg13g2_mux2_1 _18837_ (.A0(\cpu.spi.r_mode[1][0] ),
    .A1(_11982_),
    .S(_11951_),
    .X(_11983_));
 sg13g2_a22oi_1 _18838_ (.Y(_11984_),
    .B1(_11983_),
    .B2(_11962_),
    .A2(_11965_),
    .A1(\cpu.spi.r_mode[2][0] ));
 sg13g2_buf_1 _18839_ (.A(_11984_),
    .X(_11985_));
 sg13g2_nand2_1 _18840_ (.Y(_11986_),
    .A(net473),
    .B(_11985_));
 sg13g2_a21o_1 _18841_ (.A2(_09301_),
    .A1(_00219_),
    .B1(net1122),
    .X(_11987_));
 sg13g2_inv_1 _18842_ (.Y(_11988_),
    .A(_09331_));
 sg13g2_o21ai_1 _18843_ (.B1(_09339_),
    .Y(_11989_),
    .A1(_09193_),
    .A2(_11985_));
 sg13g2_nand2_1 _18844_ (.Y(_11990_),
    .A(_11988_),
    .B(_11989_));
 sg13g2_o21ai_1 _18845_ (.B1(_11990_),
    .Y(_11991_),
    .A1(_11986_),
    .A2(_11987_));
 sg13g2_nor2_1 _18846_ (.A(net1121),
    .B(_11919_),
    .Y(_11992_));
 sg13g2_buf_1 _18847_ (.A(_11985_),
    .X(_11993_));
 sg13g2_nor2_1 _18848_ (.A(_09196_),
    .B(net604),
    .Y(_11994_));
 sg13g2_a22oi_1 _18849_ (.Y(_11995_),
    .B1(_11994_),
    .B2(_09354_),
    .A2(_11992_),
    .A1(_09196_));
 sg13g2_and3_1 _18850_ (.X(_11996_),
    .A(_11981_),
    .B(_11991_),
    .C(_11995_));
 sg13g2_nor2b_1 _18851_ (.A(_11959_),
    .B_N(_11996_),
    .Y(_11997_));
 sg13g2_mux2_1 _18852_ (.A0(_11979_),
    .A1(_11980_),
    .S(_11997_),
    .X(_00318_));
 sg13g2_buf_1 _18853_ (.A(\cpu.gpio.genblk1[3].srcs_o[2] ),
    .X(_11998_));
 sg13g2_nand2_1 _18854_ (.Y(_11999_),
    .A(_11959_),
    .B(_11996_));
 sg13g2_mux2_1 _18855_ (.A0(_11980_),
    .A1(_11998_),
    .S(_11999_),
    .X(_00319_));
 sg13g2_nand2_1 _18856_ (.Y(_12000_),
    .A(net780),
    .B(_09405_));
 sg13g2_nor3_1 _18857_ (.A(_09391_),
    .B(_08468_),
    .C(_09826_),
    .Y(_12001_));
 sg13g2_buf_1 _18858_ (.A(\cpu.dcache.r_offset[2] ),
    .X(_12002_));
 sg13g2_buf_1 _18859_ (.A(\cpu.dcache.r_offset[1] ),
    .X(_12003_));
 sg13g2_inv_2 _18860_ (.Y(_12004_),
    .A(_12003_));
 sg13g2_buf_1 _18861_ (.A(\cpu.dcache.r_offset[0] ),
    .X(_12005_));
 sg13g2_inv_2 _18862_ (.Y(_12006_),
    .A(net1096));
 sg13g2_nor2_2 _18863_ (.A(_12004_),
    .B(_12006_),
    .Y(_12007_));
 sg13g2_nand3_1 _18864_ (.B(\cpu.d_wstrobe_d ),
    .C(_12007_),
    .A(_12002_),
    .Y(_12008_));
 sg13g2_buf_1 _18865_ (.A(_12008_),
    .X(_12009_));
 sg13g2_o21ai_1 _18866_ (.B1(_12009_),
    .Y(_12010_),
    .A1(_09823_),
    .A2(_09815_));
 sg13g2_and2_1 _18867_ (.A(_12001_),
    .B(_12010_),
    .X(_12011_));
 sg13g2_buf_1 _18868_ (.A(_12011_),
    .X(_12012_));
 sg13g2_nand2b_1 _18869_ (.Y(_12013_),
    .B(_12012_),
    .A_N(_12000_));
 sg13g2_buf_1 _18870_ (.A(_12013_),
    .X(_12014_));
 sg13g2_nand2_1 _18871_ (.Y(_12015_),
    .A(_08466_),
    .B(net1058));
 sg13g2_buf_2 _18872_ (.A(_00273_),
    .X(_12016_));
 sg13g2_o21ai_1 _18873_ (.B1(_12016_),
    .Y(_12017_),
    .A1(net1123),
    .A2(_12015_));
 sg13g2_nor2_1 _18874_ (.A(_12014_),
    .B(_12017_),
    .Y(_12018_));
 sg13g2_buf_2 _18875_ (.A(_12018_),
    .X(_12019_));
 sg13g2_buf_1 _18876_ (.A(_12019_),
    .X(_12020_));
 sg13g2_buf_1 _18877_ (.A(uio_in[0]),
    .X(_12021_));
 sg13g2_buf_1 _18878_ (.A(_12021_),
    .X(_12022_));
 sg13g2_buf_2 _18879_ (.A(net1095),
    .X(_12023_));
 sg13g2_buf_1 _18880_ (.A(_12000_),
    .X(_12024_));
 sg13g2_buf_1 _18881_ (.A(\cpu.d_wstrobe_d ),
    .X(_12025_));
 sg13g2_buf_1 _18882_ (.A(_00274_),
    .X(_12026_));
 sg13g2_buf_1 _18883_ (.A(_12026_),
    .X(_12027_));
 sg13g2_buf_1 _18884_ (.A(_12003_),
    .X(_12028_));
 sg13g2_nor2_1 _18885_ (.A(_12028_),
    .B(_12006_),
    .Y(_12029_));
 sg13g2_buf_2 _18886_ (.A(_12029_),
    .X(_12030_));
 sg13g2_nand3_1 _18887_ (.B(net999),
    .C(_12030_),
    .A(net1094),
    .Y(_12031_));
 sg13g2_buf_2 _18888_ (.A(_12031_),
    .X(_12032_));
 sg13g2_nor2_1 _18889_ (.A(net603),
    .B(_12032_),
    .Y(_12033_));
 sg13g2_buf_2 _18890_ (.A(_12033_),
    .X(_12034_));
 sg13g2_nor2b_1 _18891_ (.A(_12034_),
    .B_N(\cpu.dcache.r_data[0][0] ),
    .Y(_12035_));
 sg13g2_a21oi_1 _18892_ (.A1(net1000),
    .A2(_12034_),
    .Y(_12036_),
    .B1(_12035_));
 sg13g2_buf_1 _18893_ (.A(_10048_),
    .X(_12037_));
 sg13g2_nand2_1 _18894_ (.Y(_12038_),
    .A(net853),
    .B(net57));
 sg13g2_o21ai_1 _18895_ (.B1(_12038_),
    .Y(_00320_),
    .A1(net57),
    .A2(_12036_));
 sg13g2_inv_1 _18896_ (.Y(_12039_),
    .A(_12016_));
 sg13g2_mux2_1 _18897_ (.A0(net997),
    .A1(net674),
    .S(net1123),
    .X(_12040_));
 sg13g2_nor3_1 _18898_ (.A(_12014_),
    .B(_12015_),
    .C(_12040_),
    .Y(_12041_));
 sg13g2_buf_1 _18899_ (.A(_12041_),
    .X(_12042_));
 sg13g2_buf_1 _18900_ (.A(_12042_),
    .X(_12043_));
 sg13g2_buf_1 _18901_ (.A(uio_in[2]),
    .X(_12044_));
 sg13g2_buf_1 _18902_ (.A(_12044_),
    .X(_12045_));
 sg13g2_buf_2 _18903_ (.A(net1093),
    .X(_12046_));
 sg13g2_nand3_1 _18904_ (.B(net999),
    .C(_12007_),
    .A(net1094),
    .Y(_12047_));
 sg13g2_buf_2 _18905_ (.A(_12047_),
    .X(_12048_));
 sg13g2_nor2_1 _18906_ (.A(net603),
    .B(_12048_),
    .Y(_12049_));
 sg13g2_buf_2 _18907_ (.A(_12049_),
    .X(_12050_));
 sg13g2_nor2b_1 _18908_ (.A(_12050_),
    .B_N(\cpu.dcache.r_data[0][10] ),
    .Y(_12051_));
 sg13g2_a21oi_1 _18909_ (.A1(net996),
    .A2(_12050_),
    .Y(_12052_),
    .B1(_12051_));
 sg13g2_nor2b_1 _18910_ (.A(net1041),
    .B_N(_08466_),
    .Y(_12053_));
 sg13g2_buf_1 _18911_ (.A(_12053_),
    .X(_12054_));
 sg13g2_and2_1 _18912_ (.A(net1123),
    .B(_12054_),
    .X(_12055_));
 sg13g2_buf_1 _18913_ (.A(_12055_),
    .X(_12056_));
 sg13g2_mux2_1 _18914_ (.A0(_10074_),
    .A1(_10191_),
    .S(net602),
    .X(_12057_));
 sg13g2_buf_2 _18915_ (.A(_12057_),
    .X(_12058_));
 sg13g2_buf_1 _18916_ (.A(_12058_),
    .X(_12059_));
 sg13g2_nand2_1 _18917_ (.Y(_12060_),
    .A(net410),
    .B(_12042_));
 sg13g2_o21ai_1 _18918_ (.B1(_12060_),
    .Y(_00321_),
    .A1(net56),
    .A2(_12052_));
 sg13g2_buf_1 _18919_ (.A(uio_in[3]),
    .X(_12061_));
 sg13g2_buf_1 _18920_ (.A(_12061_),
    .X(_12062_));
 sg13g2_buf_2 _18921_ (.A(net1092),
    .X(_12063_));
 sg13g2_nor2b_1 _18922_ (.A(_12050_),
    .B_N(\cpu.dcache.r_data[0][11] ),
    .Y(_12064_));
 sg13g2_a21oi_1 _18923_ (.A1(net995),
    .A2(_12050_),
    .Y(_12065_),
    .B1(_12064_));
 sg13g2_mux2_1 _18924_ (.A0(net1113),
    .A1(_10198_),
    .S(net602),
    .X(_12066_));
 sg13g2_buf_2 _18925_ (.A(_12066_),
    .X(_12067_));
 sg13g2_nand2_1 _18926_ (.Y(_12068_),
    .A(net56),
    .B(_12067_));
 sg13g2_o21ai_1 _18927_ (.B1(_12068_),
    .Y(_00322_),
    .A1(net56),
    .A2(_12065_));
 sg13g2_nand2_1 _18928_ (.Y(_12069_),
    .A(net1123),
    .B(_12054_));
 sg13g2_and2_1 _18929_ (.A(_10203_),
    .B(net602),
    .X(_12070_));
 sg13g2_a21oi_1 _18930_ (.A1(_10085_),
    .A2(_12069_),
    .Y(_12071_),
    .B1(_12070_));
 sg13g2_buf_2 _18931_ (.A(_12071_),
    .X(_12072_));
 sg13g2_buf_2 _18932_ (.A(_12021_),
    .X(_12073_));
 sg13g2_nor2_1 _18933_ (.A(_12004_),
    .B(_12005_),
    .Y(_12074_));
 sg13g2_nand3_1 _18934_ (.B(_12027_),
    .C(_12074_),
    .A(net1094),
    .Y(_12075_));
 sg13g2_buf_4 _18935_ (.X(_12076_),
    .A(_12075_));
 sg13g2_nor2_2 _18936_ (.A(net603),
    .B(_12076_),
    .Y(_12077_));
 sg13g2_mux2_1 _18937_ (.A0(\cpu.dcache.r_data[0][12] ),
    .A1(net1091),
    .S(_12077_),
    .X(_12078_));
 sg13g2_nor2_1 _18938_ (.A(_12042_),
    .B(_12078_),
    .Y(_12079_));
 sg13g2_a21oi_1 _18939_ (.A1(net56),
    .A2(_12072_),
    .Y(_00323_),
    .B1(_12079_));
 sg13g2_and2_1 _18940_ (.A(_10205_),
    .B(net602),
    .X(_12080_));
 sg13g2_a21oi_1 _18941_ (.A1(_10091_),
    .A2(_12069_),
    .Y(_12081_),
    .B1(_12080_));
 sg13g2_buf_2 _18942_ (.A(_12081_),
    .X(_12082_));
 sg13g2_buf_1 _18943_ (.A(uio_in[1]),
    .X(_12083_));
 sg13g2_buf_1 _18944_ (.A(_12083_),
    .X(_12084_));
 sg13g2_mux2_1 _18945_ (.A0(\cpu.dcache.r_data[0][13] ),
    .A1(net1090),
    .S(_12077_),
    .X(_12085_));
 sg13g2_nor2_1 _18946_ (.A(_12042_),
    .B(_12085_),
    .Y(_12086_));
 sg13g2_a21oi_1 _18947_ (.A1(net56),
    .A2(_12082_),
    .Y(_00324_),
    .B1(_12086_));
 sg13g2_and2_1 _18948_ (.A(_10215_),
    .B(_12056_),
    .X(_12087_));
 sg13g2_a21oi_1 _18949_ (.A1(_10097_),
    .A2(_12069_),
    .Y(_12088_),
    .B1(_12087_));
 sg13g2_buf_2 _18950_ (.A(_12088_),
    .X(_12089_));
 sg13g2_buf_2 _18951_ (.A(_12044_),
    .X(_12090_));
 sg13g2_mux2_1 _18952_ (.A0(\cpu.dcache.r_data[0][14] ),
    .A1(net1089),
    .S(_12077_),
    .X(_12091_));
 sg13g2_nor2_1 _18953_ (.A(_12042_),
    .B(_12091_),
    .Y(_12092_));
 sg13g2_a21oi_1 _18954_ (.A1(_12043_),
    .A2(_12089_),
    .Y(_00325_),
    .B1(_12092_));
 sg13g2_and2_1 _18955_ (.A(_10220_),
    .B(net602),
    .X(_12093_));
 sg13g2_a21oi_1 _18956_ (.A1(_10103_),
    .A2(_12069_),
    .Y(_12094_),
    .B1(_12093_));
 sg13g2_buf_2 _18957_ (.A(_12094_),
    .X(_12095_));
 sg13g2_buf_2 _18958_ (.A(_12061_),
    .X(_12096_));
 sg13g2_mux2_1 _18959_ (.A0(\cpu.dcache.r_data[0][15] ),
    .A1(net1088),
    .S(_12077_),
    .X(_12097_));
 sg13g2_nor2_1 _18960_ (.A(_12042_),
    .B(_12097_),
    .Y(_12098_));
 sg13g2_a21oi_1 _18961_ (.A1(_12043_),
    .A2(_12095_),
    .Y(_00326_),
    .B1(_12098_));
 sg13g2_o21ai_1 _18962_ (.B1(net674),
    .Y(_12099_),
    .A1(net1123),
    .A2(_12015_));
 sg13g2_nor2_1 _18963_ (.A(_12014_),
    .B(_12099_),
    .Y(_12100_));
 sg13g2_buf_2 _18964_ (.A(_12100_),
    .X(_12101_));
 sg13g2_buf_1 _18965_ (.A(_12101_),
    .X(_12102_));
 sg13g2_buf_1 _18966_ (.A(_12002_),
    .X(_12103_));
 sg13g2_nand3_1 _18967_ (.B(net1094),
    .C(_12030_),
    .A(net994),
    .Y(_12104_));
 sg13g2_buf_2 _18968_ (.A(_12104_),
    .X(_12105_));
 sg13g2_nor2_1 _18969_ (.A(net603),
    .B(_12105_),
    .Y(_12106_));
 sg13g2_buf_2 _18970_ (.A(_12106_),
    .X(_12107_));
 sg13g2_nor2b_1 _18971_ (.A(_12107_),
    .B_N(\cpu.dcache.r_data[0][16] ),
    .Y(_12108_));
 sg13g2_a21oi_1 _18972_ (.A1(net1000),
    .A2(_12107_),
    .Y(_12109_),
    .B1(_12108_));
 sg13g2_nand2_1 _18973_ (.Y(_12110_),
    .A(net853),
    .B(net55));
 sg13g2_o21ai_1 _18974_ (.B1(_12110_),
    .Y(_00327_),
    .A1(_12102_),
    .A2(_12109_));
 sg13g2_buf_1 _18975_ (.A(_10115_),
    .X(_12111_));
 sg13g2_mux2_1 _18976_ (.A0(\cpu.dcache.r_data[0][17] ),
    .A1(net1090),
    .S(_12107_),
    .X(_12112_));
 sg13g2_nor2_1 _18977_ (.A(_12101_),
    .B(_12112_),
    .Y(_12113_));
 sg13g2_a21oi_1 _18978_ (.A1(net731),
    .A2(net55),
    .Y(_00328_),
    .B1(_12113_));
 sg13g2_nor2b_1 _18979_ (.A(_12107_),
    .B_N(\cpu.dcache.r_data[0][18] ),
    .Y(_12114_));
 sg13g2_a21oi_1 _18980_ (.A1(net996),
    .A2(_12107_),
    .Y(_12115_),
    .B1(_12114_));
 sg13g2_nand2_1 _18981_ (.Y(_12116_),
    .A(_10133_),
    .B(net55));
 sg13g2_o21ai_1 _18982_ (.B1(_12116_),
    .Y(_00329_),
    .A1(net55),
    .A2(_12115_));
 sg13g2_nor2b_1 _18983_ (.A(_12107_),
    .B_N(\cpu.dcache.r_data[0][19] ),
    .Y(_12117_));
 sg13g2_a21oi_1 _18984_ (.A1(net995),
    .A2(_12107_),
    .Y(_12118_),
    .B1(_12117_));
 sg13g2_buf_1 _18985_ (.A(net1113),
    .X(_12119_));
 sg13g2_nand2_1 _18986_ (.Y(_12120_),
    .A(net993),
    .B(_12101_));
 sg13g2_o21ai_1 _18987_ (.B1(_12120_),
    .Y(_00330_),
    .A1(net55),
    .A2(_12118_));
 sg13g2_mux2_1 _18988_ (.A0(\cpu.dcache.r_data[0][1] ),
    .A1(net1090),
    .S(_12034_),
    .X(_12121_));
 sg13g2_nor2_1 _18989_ (.A(_12019_),
    .B(_12121_),
    .Y(_12122_));
 sg13g2_a21oi_1 _18990_ (.A1(net731),
    .A2(net57),
    .Y(_00331_),
    .B1(_12122_));
 sg13g2_nor2_1 _18991_ (.A(net998),
    .B(net1096),
    .Y(_12123_));
 sg13g2_nand3_1 _18992_ (.B(net1094),
    .C(_12123_),
    .A(net994),
    .Y(_12124_));
 sg13g2_buf_2 _18993_ (.A(_12124_),
    .X(_12125_));
 sg13g2_nor2_1 _18994_ (.A(net603),
    .B(_12125_),
    .Y(_12126_));
 sg13g2_buf_2 _18995_ (.A(_12126_),
    .X(_12127_));
 sg13g2_nor2b_1 _18996_ (.A(_12127_),
    .B_N(\cpu.dcache.r_data[0][20] ),
    .Y(_12128_));
 sg13g2_a21oi_1 _18997_ (.A1(net1000),
    .A2(_12127_),
    .Y(_12129_),
    .B1(_12128_));
 sg13g2_buf_1 _18998_ (.A(_10085_),
    .X(_12130_));
 sg13g2_nand2_1 _18999_ (.Y(_12131_),
    .A(net992),
    .B(_12101_));
 sg13g2_o21ai_1 _19000_ (.B1(_12131_),
    .Y(_00332_),
    .A1(net55),
    .A2(_12129_));
 sg13g2_buf_1 _19001_ (.A(_12083_),
    .X(_12132_));
 sg13g2_buf_2 _19002_ (.A(net1087),
    .X(_12133_));
 sg13g2_nor2b_1 _19003_ (.A(_12127_),
    .B_N(\cpu.dcache.r_data[0][21] ),
    .Y(_12134_));
 sg13g2_a21oi_1 _19004_ (.A1(net991),
    .A2(_12127_),
    .Y(_12135_),
    .B1(_12134_));
 sg13g2_buf_1 _19005_ (.A(_10091_),
    .X(_12136_));
 sg13g2_nand2_1 _19006_ (.Y(_12137_),
    .A(net990),
    .B(_12101_));
 sg13g2_o21ai_1 _19007_ (.B1(_12137_),
    .Y(_00333_),
    .A1(net55),
    .A2(_12135_));
 sg13g2_nor2b_1 _19008_ (.A(_12127_),
    .B_N(\cpu.dcache.r_data[0][22] ),
    .Y(_12138_));
 sg13g2_a21oi_1 _19009_ (.A1(net996),
    .A2(_12127_),
    .Y(_12139_),
    .B1(_12138_));
 sg13g2_buf_1 _19010_ (.A(_10097_),
    .X(_12140_));
 sg13g2_nand2_1 _19011_ (.Y(_12141_),
    .A(net989),
    .B(_12101_));
 sg13g2_o21ai_1 _19012_ (.B1(_12141_),
    .Y(_00334_),
    .A1(net55),
    .A2(_12139_));
 sg13g2_nor2b_1 _19013_ (.A(_12127_),
    .B_N(\cpu.dcache.r_data[0][23] ),
    .Y(_12142_));
 sg13g2_a21oi_1 _19014_ (.A1(net995),
    .A2(_12127_),
    .Y(_12143_),
    .B1(_12142_));
 sg13g2_buf_1 _19015_ (.A(_10103_),
    .X(_12144_));
 sg13g2_nand2_1 _19016_ (.Y(_12145_),
    .A(_12144_),
    .B(_12101_));
 sg13g2_o21ai_1 _19017_ (.B1(_12145_),
    .Y(_00335_),
    .A1(_12102_),
    .A2(_12143_));
 sg13g2_or2_1 _19018_ (.X(_12146_),
    .B(net654),
    .A(_12024_));
 sg13g2_buf_1 _19019_ (.A(_12146_),
    .X(_12147_));
 sg13g2_mux2_1 _19020_ (.A0(net1091),
    .A1(\cpu.dcache.r_data[0][24] ),
    .S(net469),
    .X(_12148_));
 sg13g2_mux2_1 _19021_ (.A0(_10047_),
    .A1(_10181_),
    .S(net602),
    .X(_12149_));
 sg13g2_buf_2 _19022_ (.A(_12149_),
    .X(_12150_));
 sg13g2_buf_1 _19023_ (.A(_12150_),
    .X(_12151_));
 sg13g2_nand2_1 _19024_ (.Y(_12152_),
    .A(net1123),
    .B(_12016_));
 sg13g2_o21ai_1 _19025_ (.B1(_12152_),
    .Y(_12153_),
    .A1(net1123),
    .A2(_09992_));
 sg13g2_nor3_1 _19026_ (.A(_12014_),
    .B(_12015_),
    .C(_12153_),
    .Y(_12154_));
 sg13g2_buf_1 _19027_ (.A(_12154_),
    .X(_12155_));
 sg13g2_mux2_1 _19028_ (.A0(_12148_),
    .A1(net409),
    .S(net67),
    .X(_00336_));
 sg13g2_buf_4 _19029_ (.X(_12156_),
    .A(net1087));
 sg13g2_mux2_1 _19030_ (.A0(_12156_),
    .A1(\cpu.dcache.r_data[0][25] ),
    .S(net469),
    .X(_12157_));
 sg13g2_nand2_1 _19031_ (.Y(_12158_),
    .A(_10186_),
    .B(net602));
 sg13g2_o21ai_1 _19032_ (.B1(_12158_),
    .Y(_12159_),
    .A1(_10114_),
    .A2(net602));
 sg13g2_buf_2 _19033_ (.A(_12159_),
    .X(_12160_));
 sg13g2_buf_1 _19034_ (.A(_12160_),
    .X(_12161_));
 sg13g2_mux2_1 _19035_ (.A0(_12157_),
    .A1(net372),
    .S(net67),
    .X(_00337_));
 sg13g2_mux2_1 _19036_ (.A0(net1089),
    .A1(\cpu.dcache.r_data[0][26] ),
    .S(net469),
    .X(_12162_));
 sg13g2_mux2_1 _19037_ (.A0(_12162_),
    .A1(_12059_),
    .S(_12155_),
    .X(_00338_));
 sg13g2_mux2_1 _19038_ (.A0(net1088),
    .A1(\cpu.dcache.r_data[0][27] ),
    .S(net469),
    .X(_12163_));
 sg13g2_buf_1 _19039_ (.A(_12067_),
    .X(_12164_));
 sg13g2_mux2_1 _19040_ (.A0(_12163_),
    .A1(net408),
    .S(net67),
    .X(_00339_));
 sg13g2_buf_1 _19041_ (.A(_12072_),
    .X(_12165_));
 sg13g2_nand3_1 _19042_ (.B(net1094),
    .C(_12074_),
    .A(net994),
    .Y(_12166_));
 sg13g2_buf_4 _19043_ (.X(_12167_),
    .A(_12166_));
 sg13g2_nor2_2 _19044_ (.A(_12024_),
    .B(_12167_),
    .Y(_12168_));
 sg13g2_mux2_1 _19045_ (.A0(\cpu.dcache.r_data[0][28] ),
    .A1(net1091),
    .S(_12168_),
    .X(_12169_));
 sg13g2_nor2_1 _19046_ (.A(net67),
    .B(_12169_),
    .Y(_12170_));
 sg13g2_a21oi_1 _19047_ (.A1(net371),
    .A2(net67),
    .Y(_00340_),
    .B1(_12170_));
 sg13g2_buf_1 _19048_ (.A(_12082_),
    .X(_12171_));
 sg13g2_mux2_1 _19049_ (.A0(\cpu.dcache.r_data[0][29] ),
    .A1(_12084_),
    .S(_12168_),
    .X(_12172_));
 sg13g2_nor2_1 _19050_ (.A(net67),
    .B(_12172_),
    .Y(_12173_));
 sg13g2_a21oi_1 _19051_ (.A1(_12171_),
    .A2(net67),
    .Y(_00341_),
    .B1(_12173_));
 sg13g2_nor2b_1 _19052_ (.A(_12034_),
    .B_N(\cpu.dcache.r_data[0][2] ),
    .Y(_12174_));
 sg13g2_a21oi_1 _19053_ (.A1(net996),
    .A2(_12034_),
    .Y(_12175_),
    .B1(_12174_));
 sg13g2_buf_1 _19054_ (.A(_10132_),
    .X(_12176_));
 sg13g2_nand2_1 _19055_ (.Y(_12177_),
    .A(net852),
    .B(net57));
 sg13g2_o21ai_1 _19056_ (.B1(_12177_),
    .Y(_00342_),
    .A1(_12020_),
    .A2(_12175_));
 sg13g2_buf_1 _19057_ (.A(_12089_),
    .X(_12178_));
 sg13g2_mux2_1 _19058_ (.A0(\cpu.dcache.r_data[0][30] ),
    .A1(net1089),
    .S(_12168_),
    .X(_12179_));
 sg13g2_nor2_1 _19059_ (.A(_12154_),
    .B(_12179_),
    .Y(_12180_));
 sg13g2_a21oi_1 _19060_ (.A1(net369),
    .A2(_12155_),
    .Y(_00343_),
    .B1(_12180_));
 sg13g2_buf_1 _19061_ (.A(_12095_),
    .X(_12181_));
 sg13g2_mux2_1 _19062_ (.A0(\cpu.dcache.r_data[0][31] ),
    .A1(net1088),
    .S(_12168_),
    .X(_12182_));
 sg13g2_nor2_1 _19063_ (.A(_12154_),
    .B(_12182_),
    .Y(_12183_));
 sg13g2_a21oi_1 _19064_ (.A1(_12181_),
    .A2(net67),
    .Y(_00344_),
    .B1(_12183_));
 sg13g2_nor2b_1 _19065_ (.A(_12034_),
    .B_N(\cpu.dcache.r_data[0][3] ),
    .Y(_12184_));
 sg13g2_a21oi_1 _19066_ (.A1(net995),
    .A2(_12034_),
    .Y(_12185_),
    .B1(_12184_));
 sg13g2_nand2_1 _19067_ (.Y(_12186_),
    .A(net993),
    .B(_12019_));
 sg13g2_o21ai_1 _19068_ (.B1(_12186_),
    .Y(_00345_),
    .A1(_12020_),
    .A2(_12185_));
 sg13g2_nand3_1 _19069_ (.B(net999),
    .C(_12123_),
    .A(net1094),
    .Y(_12187_));
 sg13g2_buf_2 _19070_ (.A(_12187_),
    .X(_12188_));
 sg13g2_nor2_1 _19071_ (.A(net603),
    .B(_12188_),
    .Y(_12189_));
 sg13g2_buf_2 _19072_ (.A(_12189_),
    .X(_12190_));
 sg13g2_nor2b_1 _19073_ (.A(_12190_),
    .B_N(\cpu.dcache.r_data[0][4] ),
    .Y(_12191_));
 sg13g2_a21oi_1 _19074_ (.A1(net1000),
    .A2(_12190_),
    .Y(_12192_),
    .B1(_12191_));
 sg13g2_buf_1 _19075_ (.A(_10085_),
    .X(_12193_));
 sg13g2_nand2_1 _19076_ (.Y(_12194_),
    .A(net987),
    .B(_12019_));
 sg13g2_o21ai_1 _19077_ (.B1(_12194_),
    .Y(_00346_),
    .A1(net57),
    .A2(_12192_));
 sg13g2_nor2b_1 _19078_ (.A(_12190_),
    .B_N(\cpu.dcache.r_data[0][5] ),
    .Y(_12195_));
 sg13g2_a21oi_1 _19079_ (.A1(net991),
    .A2(_12190_),
    .Y(_12196_),
    .B1(_12195_));
 sg13g2_nand2_1 _19080_ (.Y(_12197_),
    .A(net990),
    .B(_12019_));
 sg13g2_o21ai_1 _19081_ (.B1(_12197_),
    .Y(_00347_),
    .A1(net57),
    .A2(_12196_));
 sg13g2_nor2b_1 _19082_ (.A(_12190_),
    .B_N(\cpu.dcache.r_data[0][6] ),
    .Y(_12198_));
 sg13g2_a21oi_1 _19083_ (.A1(net996),
    .A2(_12190_),
    .Y(_12199_),
    .B1(_12198_));
 sg13g2_nand2_1 _19084_ (.Y(_12200_),
    .A(_12140_),
    .B(_12019_));
 sg13g2_o21ai_1 _19085_ (.B1(_12200_),
    .Y(_00348_),
    .A1(net57),
    .A2(_12199_));
 sg13g2_nor2b_1 _19086_ (.A(_12190_),
    .B_N(\cpu.dcache.r_data[0][7] ),
    .Y(_12201_));
 sg13g2_a21oi_1 _19087_ (.A1(net995),
    .A2(_12190_),
    .Y(_12202_),
    .B1(_12201_));
 sg13g2_nand2_1 _19088_ (.Y(_12203_),
    .A(net988),
    .B(_12019_));
 sg13g2_o21ai_1 _19089_ (.B1(_12203_),
    .Y(_00349_),
    .A1(net57),
    .A2(_12202_));
 sg13g2_nor2b_1 _19090_ (.A(_12050_),
    .B_N(\cpu.dcache.r_data[0][8] ),
    .Y(_12204_));
 sg13g2_a21oi_1 _19091_ (.A1(net1000),
    .A2(_12050_),
    .Y(_12205_),
    .B1(_12204_));
 sg13g2_nand2_1 _19092_ (.Y(_12206_),
    .A(net56),
    .B(_12150_));
 sg13g2_o21ai_1 _19093_ (.B1(_12206_),
    .Y(_00350_),
    .A1(net56),
    .A2(_12205_));
 sg13g2_nor2b_1 _19094_ (.A(_12050_),
    .B_N(\cpu.dcache.r_data[0][9] ),
    .Y(_12207_));
 sg13g2_a21oi_1 _19095_ (.A1(net991),
    .A2(_12050_),
    .Y(_12208_),
    .B1(_12207_));
 sg13g2_nand2_1 _19096_ (.Y(_12209_),
    .A(_12042_),
    .B(_12160_));
 sg13g2_o21ai_1 _19097_ (.B1(_12209_),
    .Y(_00351_),
    .A1(net56),
    .A2(_12208_));
 sg13g2_nand2_1 _19098_ (.Y(_12210_),
    .A(net1119),
    .B(_09421_));
 sg13g2_buf_2 _19099_ (.A(_12210_),
    .X(_12211_));
 sg13g2_buf_1 _19100_ (.A(_12211_),
    .X(_12212_));
 sg13g2_inv_1 _19101_ (.Y(_12213_),
    .A(_12017_));
 sg13g2_nand2_1 _19102_ (.Y(_12214_),
    .A(_12012_),
    .B(_12213_));
 sg13g2_buf_2 _19103_ (.A(_12214_),
    .X(_12215_));
 sg13g2_nor2_1 _19104_ (.A(net601),
    .B(_12215_),
    .Y(_12216_));
 sg13g2_buf_2 _19105_ (.A(_12216_),
    .X(_12217_));
 sg13g2_buf_1 _19106_ (.A(_12217_),
    .X(_12218_));
 sg13g2_nor2_1 _19107_ (.A(_12211_),
    .B(_12032_),
    .Y(_12219_));
 sg13g2_buf_2 _19108_ (.A(_12219_),
    .X(_12220_));
 sg13g2_nor2b_1 _19109_ (.A(_12220_),
    .B_N(\cpu.dcache.r_data[1][0] ),
    .Y(_12221_));
 sg13g2_a21oi_1 _19110_ (.A1(net1000),
    .A2(_12220_),
    .Y(_12222_),
    .B1(_12221_));
 sg13g2_nand2_1 _19111_ (.Y(_12223_),
    .A(net853),
    .B(_12218_));
 sg13g2_o21ai_1 _19112_ (.B1(_12223_),
    .Y(_00352_),
    .A1(net54),
    .A2(_12222_));
 sg13g2_nand3b_1 _19113_ (.B(_12054_),
    .C(_12012_),
    .Y(_12224_),
    .A_N(_12040_));
 sg13g2_buf_2 _19114_ (.A(_12224_),
    .X(_12225_));
 sg13g2_nor2_1 _19115_ (.A(net601),
    .B(_12225_),
    .Y(_12226_));
 sg13g2_buf_2 _19116_ (.A(_12226_),
    .X(_12227_));
 sg13g2_buf_1 _19117_ (.A(_12227_),
    .X(_12228_));
 sg13g2_nor2_1 _19118_ (.A(net601),
    .B(_12048_),
    .Y(_12229_));
 sg13g2_buf_2 _19119_ (.A(_12229_),
    .X(_12230_));
 sg13g2_nor2b_1 _19120_ (.A(_12230_),
    .B_N(\cpu.dcache.r_data[1][10] ),
    .Y(_12231_));
 sg13g2_a21oi_1 _19121_ (.A1(net996),
    .A2(_12230_),
    .Y(_12232_),
    .B1(_12231_));
 sg13g2_nand2_1 _19122_ (.Y(_12233_),
    .A(net410),
    .B(net53));
 sg13g2_o21ai_1 _19123_ (.B1(_12233_),
    .Y(_00353_),
    .A1(net53),
    .A2(_12232_));
 sg13g2_nor2b_1 _19124_ (.A(_12230_),
    .B_N(\cpu.dcache.r_data[1][11] ),
    .Y(_12234_));
 sg13g2_a21oi_1 _19125_ (.A1(net995),
    .A2(_12230_),
    .Y(_12235_),
    .B1(_12234_));
 sg13g2_nand2_1 _19126_ (.Y(_12236_),
    .A(net408),
    .B(net53));
 sg13g2_o21ai_1 _19127_ (.B1(_12236_),
    .Y(_00354_),
    .A1(net53),
    .A2(_12235_));
 sg13g2_buf_1 _19128_ (.A(_12021_),
    .X(_12237_));
 sg13g2_nor2_2 _19129_ (.A(net601),
    .B(_12076_),
    .Y(_12238_));
 sg13g2_mux2_1 _19130_ (.A0(\cpu.dcache.r_data[1][12] ),
    .A1(net1086),
    .S(_12238_),
    .X(_12239_));
 sg13g2_nor2_1 _19131_ (.A(_12227_),
    .B(_12239_),
    .Y(_12240_));
 sg13g2_a21oi_1 _19132_ (.A1(net371),
    .A2(net53),
    .Y(_00355_),
    .B1(_12240_));
 sg13g2_mux2_1 _19133_ (.A0(\cpu.dcache.r_data[1][13] ),
    .A1(net1090),
    .S(_12238_),
    .X(_12241_));
 sg13g2_nor2_1 _19134_ (.A(_12227_),
    .B(_12241_),
    .Y(_12242_));
 sg13g2_a21oi_1 _19135_ (.A1(net370),
    .A2(net53),
    .Y(_00356_),
    .B1(_12242_));
 sg13g2_buf_1 _19136_ (.A(_12044_),
    .X(_12243_));
 sg13g2_mux2_1 _19137_ (.A0(\cpu.dcache.r_data[1][14] ),
    .A1(net1085),
    .S(_12238_),
    .X(_12244_));
 sg13g2_nor2_1 _19138_ (.A(_12227_),
    .B(_12244_),
    .Y(_12245_));
 sg13g2_a21oi_1 _19139_ (.A1(net369),
    .A2(_12228_),
    .Y(_00357_),
    .B1(_12245_));
 sg13g2_buf_1 _19140_ (.A(_12061_),
    .X(_12246_));
 sg13g2_mux2_1 _19141_ (.A0(\cpu.dcache.r_data[1][15] ),
    .A1(net1084),
    .S(_12238_),
    .X(_12247_));
 sg13g2_nor2_1 _19142_ (.A(_12227_),
    .B(_12247_),
    .Y(_12248_));
 sg13g2_a21oi_1 _19143_ (.A1(net368),
    .A2(_12228_),
    .Y(_00358_),
    .B1(_12248_));
 sg13g2_inv_1 _19144_ (.Y(_12249_),
    .A(_12099_));
 sg13g2_nand2_1 _19145_ (.Y(_12250_),
    .A(_12012_),
    .B(_12249_));
 sg13g2_buf_2 _19146_ (.A(_12250_),
    .X(_12251_));
 sg13g2_nor2_1 _19147_ (.A(net601),
    .B(_12251_),
    .Y(_12252_));
 sg13g2_buf_2 _19148_ (.A(_12252_),
    .X(_12253_));
 sg13g2_buf_1 _19149_ (.A(_12253_),
    .X(_12254_));
 sg13g2_buf_1 _19150_ (.A(net1095),
    .X(_12255_));
 sg13g2_nor2_1 _19151_ (.A(_12211_),
    .B(_12105_),
    .Y(_12256_));
 sg13g2_buf_2 _19152_ (.A(_12256_),
    .X(_12257_));
 sg13g2_nor2b_1 _19153_ (.A(_12257_),
    .B_N(\cpu.dcache.r_data[1][16] ),
    .Y(_12258_));
 sg13g2_a21oi_1 _19154_ (.A1(net986),
    .A2(_12257_),
    .Y(_12259_),
    .B1(_12258_));
 sg13g2_nand2_1 _19155_ (.Y(_12260_),
    .A(net853),
    .B(_12254_));
 sg13g2_o21ai_1 _19156_ (.B1(_12260_),
    .Y(_00359_),
    .A1(net52),
    .A2(_12259_));
 sg13g2_mux2_1 _19157_ (.A0(\cpu.dcache.r_data[1][17] ),
    .A1(net1090),
    .S(_12257_),
    .X(_12261_));
 sg13g2_nor2_1 _19158_ (.A(_12253_),
    .B(_12261_),
    .Y(_12262_));
 sg13g2_a21oi_1 _19159_ (.A1(net731),
    .A2(net52),
    .Y(_00360_),
    .B1(_12262_));
 sg13g2_buf_1 _19160_ (.A(net1093),
    .X(_12263_));
 sg13g2_nor2b_1 _19161_ (.A(_12257_),
    .B_N(\cpu.dcache.r_data[1][18] ),
    .Y(_12264_));
 sg13g2_a21oi_1 _19162_ (.A1(net985),
    .A2(_12257_),
    .Y(_12265_),
    .B1(_12264_));
 sg13g2_nand2_1 _19163_ (.Y(_12266_),
    .A(net852),
    .B(net52));
 sg13g2_o21ai_1 _19164_ (.B1(_12266_),
    .Y(_00361_),
    .A1(net52),
    .A2(_12265_));
 sg13g2_buf_1 _19165_ (.A(net1092),
    .X(_12267_));
 sg13g2_nor2b_1 _19166_ (.A(_12257_),
    .B_N(\cpu.dcache.r_data[1][19] ),
    .Y(_12268_));
 sg13g2_a21oi_1 _19167_ (.A1(net984),
    .A2(_12257_),
    .Y(_12269_),
    .B1(_12268_));
 sg13g2_nand2_1 _19168_ (.Y(_12270_),
    .A(net993),
    .B(_12253_));
 sg13g2_o21ai_1 _19169_ (.B1(_12270_),
    .Y(_00362_),
    .A1(net52),
    .A2(_12269_));
 sg13g2_buf_1 _19170_ (.A(_12083_),
    .X(_12271_));
 sg13g2_mux2_1 _19171_ (.A0(\cpu.dcache.r_data[1][1] ),
    .A1(net1083),
    .S(_12220_),
    .X(_12272_));
 sg13g2_nor2_1 _19172_ (.A(_12217_),
    .B(_12272_),
    .Y(_12273_));
 sg13g2_a21oi_1 _19173_ (.A1(net731),
    .A2(net54),
    .Y(_00363_),
    .B1(_12273_));
 sg13g2_nor2_1 _19174_ (.A(net601),
    .B(_12125_),
    .Y(_12274_));
 sg13g2_buf_2 _19175_ (.A(_12274_),
    .X(_12275_));
 sg13g2_nor2b_1 _19176_ (.A(_12275_),
    .B_N(\cpu.dcache.r_data[1][20] ),
    .Y(_12276_));
 sg13g2_a21oi_1 _19177_ (.A1(net986),
    .A2(_12275_),
    .Y(_12277_),
    .B1(_12276_));
 sg13g2_nand2_1 _19178_ (.Y(_12278_),
    .A(net987),
    .B(_12253_));
 sg13g2_o21ai_1 _19179_ (.B1(_12278_),
    .Y(_00364_),
    .A1(net52),
    .A2(_12277_));
 sg13g2_nor2b_1 _19180_ (.A(_12275_),
    .B_N(\cpu.dcache.r_data[1][21] ),
    .Y(_12279_));
 sg13g2_a21oi_1 _19181_ (.A1(net991),
    .A2(_12275_),
    .Y(_12280_),
    .B1(_12279_));
 sg13g2_buf_1 _19182_ (.A(_10091_),
    .X(_12281_));
 sg13g2_nand2_1 _19183_ (.Y(_12282_),
    .A(_12281_),
    .B(_12253_));
 sg13g2_o21ai_1 _19184_ (.B1(_12282_),
    .Y(_00365_),
    .A1(net52),
    .A2(_12280_));
 sg13g2_nor2b_1 _19185_ (.A(_12275_),
    .B_N(\cpu.dcache.r_data[1][22] ),
    .Y(_12283_));
 sg13g2_a21oi_1 _19186_ (.A1(net985),
    .A2(_12275_),
    .Y(_12284_),
    .B1(_12283_));
 sg13g2_nand2_1 _19187_ (.Y(_12285_),
    .A(net989),
    .B(_12253_));
 sg13g2_o21ai_1 _19188_ (.B1(_12285_),
    .Y(_00366_),
    .A1(net52),
    .A2(_12284_));
 sg13g2_nor2b_1 _19189_ (.A(_12275_),
    .B_N(\cpu.dcache.r_data[1][23] ),
    .Y(_12286_));
 sg13g2_a21oi_1 _19190_ (.A1(net984),
    .A2(_12275_),
    .Y(_12287_),
    .B1(_12286_));
 sg13g2_nand2_1 _19191_ (.Y(_12288_),
    .A(net988),
    .B(_12253_));
 sg13g2_o21ai_1 _19192_ (.B1(_12288_),
    .Y(_00367_),
    .A1(_12254_),
    .A2(_12287_));
 sg13g2_nand3b_1 _19193_ (.B(_12054_),
    .C(_12012_),
    .Y(_12289_),
    .A_N(_12153_));
 sg13g2_buf_2 _19194_ (.A(_12289_),
    .X(_12290_));
 sg13g2_nor2_1 _19195_ (.A(_12212_),
    .B(_12290_),
    .Y(_12291_));
 sg13g2_buf_2 _19196_ (.A(_12291_),
    .X(_12292_));
 sg13g2_buf_1 _19197_ (.A(_12292_),
    .X(_12293_));
 sg13g2_nor2_1 _19198_ (.A(_12211_),
    .B(net654),
    .Y(_12294_));
 sg13g2_buf_1 _19199_ (.A(_12294_),
    .X(_12295_));
 sg13g2_nor2b_1 _19200_ (.A(net529),
    .B_N(\cpu.dcache.r_data[1][24] ),
    .Y(_12296_));
 sg13g2_a21oi_1 _19201_ (.A1(_12255_),
    .A2(net529),
    .Y(_12297_),
    .B1(_12296_));
 sg13g2_nand2_1 _19202_ (.Y(_12298_),
    .A(net409),
    .B(net51));
 sg13g2_o21ai_1 _19203_ (.B1(_12298_),
    .Y(_00368_),
    .A1(net51),
    .A2(_12297_));
 sg13g2_nor2b_1 _19204_ (.A(net529),
    .B_N(\cpu.dcache.r_data[1][25] ),
    .Y(_12299_));
 sg13g2_a21oi_1 _19205_ (.A1(net991),
    .A2(net529),
    .Y(_12300_),
    .B1(_12299_));
 sg13g2_nand2_1 _19206_ (.Y(_12301_),
    .A(net372),
    .B(net51));
 sg13g2_o21ai_1 _19207_ (.B1(_12301_),
    .Y(_00369_),
    .A1(net51),
    .A2(_12300_));
 sg13g2_nor2b_1 _19208_ (.A(net529),
    .B_N(\cpu.dcache.r_data[1][26] ),
    .Y(_12302_));
 sg13g2_a21oi_1 _19209_ (.A1(_12263_),
    .A2(net529),
    .Y(_12303_),
    .B1(_12302_));
 sg13g2_nand2_1 _19210_ (.Y(_12304_),
    .A(net410),
    .B(_12292_));
 sg13g2_o21ai_1 _19211_ (.B1(_12304_),
    .Y(_00370_),
    .A1(_12293_),
    .A2(_12303_));
 sg13g2_nor2b_1 _19212_ (.A(_12295_),
    .B_N(\cpu.dcache.r_data[1][27] ),
    .Y(_12305_));
 sg13g2_a21oi_1 _19213_ (.A1(_12267_),
    .A2(_12295_),
    .Y(_12306_),
    .B1(_12305_));
 sg13g2_nand2_1 _19214_ (.Y(_12307_),
    .A(net408),
    .B(_12292_));
 sg13g2_o21ai_1 _19215_ (.B1(_12307_),
    .Y(_00371_),
    .A1(_12293_),
    .A2(_12306_));
 sg13g2_nor2_2 _19216_ (.A(net601),
    .B(_12167_),
    .Y(_12308_));
 sg13g2_mux2_1 _19217_ (.A0(\cpu.dcache.r_data[1][28] ),
    .A1(_12237_),
    .S(_12308_),
    .X(_12309_));
 sg13g2_nor2_1 _19218_ (.A(_12292_),
    .B(_12309_),
    .Y(_12310_));
 sg13g2_a21oi_1 _19219_ (.A1(net371),
    .A2(net51),
    .Y(_00372_),
    .B1(_12310_));
 sg13g2_mux2_1 _19220_ (.A0(\cpu.dcache.r_data[1][29] ),
    .A1(net1083),
    .S(_12308_),
    .X(_12311_));
 sg13g2_nor2_1 _19221_ (.A(_12292_),
    .B(_12311_),
    .Y(_12312_));
 sg13g2_a21oi_1 _19222_ (.A1(net370),
    .A2(net51),
    .Y(_00373_),
    .B1(_12312_));
 sg13g2_nor2b_1 _19223_ (.A(_12220_),
    .B_N(\cpu.dcache.r_data[1][2] ),
    .Y(_12313_));
 sg13g2_a21oi_1 _19224_ (.A1(net985),
    .A2(_12220_),
    .Y(_12314_),
    .B1(_12313_));
 sg13g2_nand2_1 _19225_ (.Y(_12315_),
    .A(net852),
    .B(net54));
 sg13g2_o21ai_1 _19226_ (.B1(_12315_),
    .Y(_00374_),
    .A1(_12218_),
    .A2(_12314_));
 sg13g2_mux2_1 _19227_ (.A0(\cpu.dcache.r_data[1][30] ),
    .A1(net1085),
    .S(_12308_),
    .X(_12316_));
 sg13g2_nor2_1 _19228_ (.A(_12292_),
    .B(_12316_),
    .Y(_12317_));
 sg13g2_a21oi_1 _19229_ (.A1(net369),
    .A2(net51),
    .Y(_00375_),
    .B1(_12317_));
 sg13g2_mux2_1 _19230_ (.A0(\cpu.dcache.r_data[1][31] ),
    .A1(net1084),
    .S(_12308_),
    .X(_12318_));
 sg13g2_nor2_1 _19231_ (.A(_12292_),
    .B(_12318_),
    .Y(_12319_));
 sg13g2_a21oi_1 _19232_ (.A1(net368),
    .A2(net51),
    .Y(_00376_),
    .B1(_12319_));
 sg13g2_nor2b_1 _19233_ (.A(_12220_),
    .B_N(\cpu.dcache.r_data[1][3] ),
    .Y(_12320_));
 sg13g2_a21oi_1 _19234_ (.A1(net984),
    .A2(_12220_),
    .Y(_12321_),
    .B1(_12320_));
 sg13g2_nand2_1 _19235_ (.Y(_12322_),
    .A(net993),
    .B(_12217_));
 sg13g2_o21ai_1 _19236_ (.B1(_12322_),
    .Y(_00377_),
    .A1(net54),
    .A2(_12321_));
 sg13g2_nor2_1 _19237_ (.A(_12211_),
    .B(_12188_),
    .Y(_12323_));
 sg13g2_buf_2 _19238_ (.A(_12323_),
    .X(_12324_));
 sg13g2_nor2b_1 _19239_ (.A(_12324_),
    .B_N(\cpu.dcache.r_data[1][4] ),
    .Y(_12325_));
 sg13g2_a21oi_1 _19240_ (.A1(net986),
    .A2(_12324_),
    .Y(_12326_),
    .B1(_12325_));
 sg13g2_nand2_1 _19241_ (.Y(_12327_),
    .A(net987),
    .B(_12217_));
 sg13g2_o21ai_1 _19242_ (.B1(_12327_),
    .Y(_00378_),
    .A1(net54),
    .A2(_12326_));
 sg13g2_nor2b_1 _19243_ (.A(_12324_),
    .B_N(\cpu.dcache.r_data[1][5] ),
    .Y(_12328_));
 sg13g2_a21oi_1 _19244_ (.A1(net991),
    .A2(_12324_),
    .Y(_12329_),
    .B1(_12328_));
 sg13g2_nand2_1 _19245_ (.Y(_12330_),
    .A(net983),
    .B(_12217_));
 sg13g2_o21ai_1 _19246_ (.B1(_12330_),
    .Y(_00379_),
    .A1(net54),
    .A2(_12329_));
 sg13g2_nor2b_1 _19247_ (.A(_12324_),
    .B_N(\cpu.dcache.r_data[1][6] ),
    .Y(_12331_));
 sg13g2_a21oi_1 _19248_ (.A1(net985),
    .A2(_12324_),
    .Y(_12332_),
    .B1(_12331_));
 sg13g2_buf_1 _19249_ (.A(_10097_),
    .X(_12333_));
 sg13g2_nand2_1 _19250_ (.Y(_12334_),
    .A(net982),
    .B(_12217_));
 sg13g2_o21ai_1 _19251_ (.B1(_12334_),
    .Y(_00380_),
    .A1(net54),
    .A2(_12332_));
 sg13g2_nor2b_1 _19252_ (.A(_12324_),
    .B_N(\cpu.dcache.r_data[1][7] ),
    .Y(_12335_));
 sg13g2_a21oi_1 _19253_ (.A1(net984),
    .A2(_12324_),
    .Y(_12336_),
    .B1(_12335_));
 sg13g2_nand2_1 _19254_ (.Y(_12337_),
    .A(net988),
    .B(_12217_));
 sg13g2_o21ai_1 _19255_ (.B1(_12337_),
    .Y(_00381_),
    .A1(net54),
    .A2(_12336_));
 sg13g2_nor2b_1 _19256_ (.A(_12230_),
    .B_N(\cpu.dcache.r_data[1][8] ),
    .Y(_12338_));
 sg13g2_a21oi_1 _19257_ (.A1(net986),
    .A2(_12230_),
    .Y(_12339_),
    .B1(_12338_));
 sg13g2_nand2_1 _19258_ (.Y(_12340_),
    .A(net409),
    .B(_12227_));
 sg13g2_o21ai_1 _19259_ (.B1(_12340_),
    .Y(_00382_),
    .A1(net53),
    .A2(_12339_));
 sg13g2_buf_1 _19260_ (.A(_12132_),
    .X(_12341_));
 sg13g2_nor2b_1 _19261_ (.A(_12230_),
    .B_N(\cpu.dcache.r_data[1][9] ),
    .Y(_12342_));
 sg13g2_a21oi_1 _19262_ (.A1(net981),
    .A2(_12230_),
    .Y(_12343_),
    .B1(_12342_));
 sg13g2_nand2_1 _19263_ (.Y(_12344_),
    .A(net372),
    .B(_12227_));
 sg13g2_o21ai_1 _19264_ (.B1(_12344_),
    .Y(_00383_),
    .A1(net53),
    .A2(_12343_));
 sg13g2_nand2_1 _19265_ (.Y(_12345_),
    .A(net632),
    .B(_09405_));
 sg13g2_buf_1 _19266_ (.A(_12345_),
    .X(_12346_));
 sg13g2_buf_1 _19267_ (.A(_12346_),
    .X(_12347_));
 sg13g2_nor2_1 _19268_ (.A(net407),
    .B(_12215_),
    .Y(_12348_));
 sg13g2_buf_2 _19269_ (.A(_12348_),
    .X(_12349_));
 sg13g2_buf_1 _19270_ (.A(_12349_),
    .X(_12350_));
 sg13g2_nor2_1 _19271_ (.A(_12346_),
    .B(_12032_),
    .Y(_12351_));
 sg13g2_buf_2 _19272_ (.A(_12351_),
    .X(_12352_));
 sg13g2_nor2b_1 _19273_ (.A(_12352_),
    .B_N(\cpu.dcache.r_data[2][0] ),
    .Y(_12353_));
 sg13g2_a21oi_1 _19274_ (.A1(net986),
    .A2(_12352_),
    .Y(_12354_),
    .B1(_12353_));
 sg13g2_nand2_1 _19275_ (.Y(_12355_),
    .A(net853),
    .B(_12350_));
 sg13g2_o21ai_1 _19276_ (.B1(_12355_),
    .Y(_00384_),
    .A1(net50),
    .A2(_12354_));
 sg13g2_nor2_1 _19277_ (.A(net407),
    .B(_12225_),
    .Y(_12356_));
 sg13g2_buf_1 _19278_ (.A(_12356_),
    .X(_12357_));
 sg13g2_buf_1 _19279_ (.A(_12357_),
    .X(_12358_));
 sg13g2_nor2_1 _19280_ (.A(net407),
    .B(_12048_),
    .Y(_12359_));
 sg13g2_buf_2 _19281_ (.A(_12359_),
    .X(_12360_));
 sg13g2_nor2b_1 _19282_ (.A(_12360_),
    .B_N(\cpu.dcache.r_data[2][10] ),
    .Y(_12361_));
 sg13g2_a21oi_1 _19283_ (.A1(net985),
    .A2(_12360_),
    .Y(_12362_),
    .B1(_12361_));
 sg13g2_nand2_1 _19284_ (.Y(_12363_),
    .A(net410),
    .B(net49));
 sg13g2_o21ai_1 _19285_ (.B1(_12363_),
    .Y(_00385_),
    .A1(net49),
    .A2(_12362_));
 sg13g2_nor2b_1 _19286_ (.A(_12360_),
    .B_N(\cpu.dcache.r_data[2][11] ),
    .Y(_12364_));
 sg13g2_a21oi_1 _19287_ (.A1(net984),
    .A2(_12360_),
    .Y(_12365_),
    .B1(_12364_));
 sg13g2_nand2_1 _19288_ (.Y(_12366_),
    .A(net408),
    .B(net49));
 sg13g2_o21ai_1 _19289_ (.B1(_12366_),
    .Y(_00386_),
    .A1(net49),
    .A2(_12365_));
 sg13g2_nor2_2 _19290_ (.A(net407),
    .B(_12076_),
    .Y(_12367_));
 sg13g2_mux2_1 _19291_ (.A0(\cpu.dcache.r_data[2][12] ),
    .A1(net1086),
    .S(_12367_),
    .X(_12368_));
 sg13g2_nor2_1 _19292_ (.A(_12357_),
    .B(_12368_),
    .Y(_12369_));
 sg13g2_a21oi_1 _19293_ (.A1(net371),
    .A2(net49),
    .Y(_00387_),
    .B1(_12369_));
 sg13g2_mux2_1 _19294_ (.A0(\cpu.dcache.r_data[2][13] ),
    .A1(net1083),
    .S(_12367_),
    .X(_12370_));
 sg13g2_nor2_1 _19295_ (.A(_12357_),
    .B(_12370_),
    .Y(_12371_));
 sg13g2_a21oi_1 _19296_ (.A1(net370),
    .A2(net49),
    .Y(_00388_),
    .B1(_12371_));
 sg13g2_mux2_1 _19297_ (.A0(\cpu.dcache.r_data[2][14] ),
    .A1(net1085),
    .S(_12367_),
    .X(_12372_));
 sg13g2_nor2_1 _19298_ (.A(_12357_),
    .B(_12372_),
    .Y(_12373_));
 sg13g2_a21oi_1 _19299_ (.A1(net369),
    .A2(_12358_),
    .Y(_00389_),
    .B1(_12373_));
 sg13g2_mux2_1 _19300_ (.A0(\cpu.dcache.r_data[2][15] ),
    .A1(net1084),
    .S(_12367_),
    .X(_12374_));
 sg13g2_nor2_1 _19301_ (.A(_12357_),
    .B(_12374_),
    .Y(_12375_));
 sg13g2_a21oi_1 _19302_ (.A1(net368),
    .A2(_12358_),
    .Y(_00390_),
    .B1(_12375_));
 sg13g2_nor2_1 _19303_ (.A(net407),
    .B(_12251_),
    .Y(_12376_));
 sg13g2_buf_2 _19304_ (.A(_12376_),
    .X(_12377_));
 sg13g2_buf_1 _19305_ (.A(_12377_),
    .X(_12378_));
 sg13g2_nor2_1 _19306_ (.A(_12346_),
    .B(_12105_),
    .Y(_12379_));
 sg13g2_buf_2 _19307_ (.A(_12379_),
    .X(_12380_));
 sg13g2_nor2b_1 _19308_ (.A(_12380_),
    .B_N(\cpu.dcache.r_data[2][16] ),
    .Y(_12381_));
 sg13g2_a21oi_1 _19309_ (.A1(net986),
    .A2(_12380_),
    .Y(_12382_),
    .B1(_12381_));
 sg13g2_nand2_1 _19310_ (.Y(_12383_),
    .A(net853),
    .B(net48));
 sg13g2_o21ai_1 _19311_ (.B1(_12383_),
    .Y(_00391_),
    .A1(net48),
    .A2(_12382_));
 sg13g2_mux2_1 _19312_ (.A0(\cpu.dcache.r_data[2][17] ),
    .A1(net1083),
    .S(_12380_),
    .X(_12384_));
 sg13g2_nor2_1 _19313_ (.A(_12377_),
    .B(_12384_),
    .Y(_12385_));
 sg13g2_a21oi_1 _19314_ (.A1(net731),
    .A2(net48),
    .Y(_00392_),
    .B1(_12385_));
 sg13g2_nor2b_1 _19315_ (.A(_12380_),
    .B_N(\cpu.dcache.r_data[2][18] ),
    .Y(_12386_));
 sg13g2_a21oi_1 _19316_ (.A1(net985),
    .A2(_12380_),
    .Y(_12387_),
    .B1(_12386_));
 sg13g2_nand2_1 _19317_ (.Y(_12388_),
    .A(net852),
    .B(net48));
 sg13g2_o21ai_1 _19318_ (.B1(_12388_),
    .Y(_00393_),
    .A1(net48),
    .A2(_12387_));
 sg13g2_nor2b_1 _19319_ (.A(_12380_),
    .B_N(\cpu.dcache.r_data[2][19] ),
    .Y(_12389_));
 sg13g2_a21oi_1 _19320_ (.A1(net984),
    .A2(_12380_),
    .Y(_12390_),
    .B1(_12389_));
 sg13g2_nand2_1 _19321_ (.Y(_12391_),
    .A(net993),
    .B(_12377_));
 sg13g2_o21ai_1 _19322_ (.B1(_12391_),
    .Y(_00394_),
    .A1(net48),
    .A2(_12390_));
 sg13g2_mux2_1 _19323_ (.A0(\cpu.dcache.r_data[2][1] ),
    .A1(net1083),
    .S(_12352_),
    .X(_12392_));
 sg13g2_nor2_1 _19324_ (.A(_12349_),
    .B(_12392_),
    .Y(_12393_));
 sg13g2_a21oi_1 _19325_ (.A1(net731),
    .A2(net50),
    .Y(_00395_),
    .B1(_12393_));
 sg13g2_nor2_1 _19326_ (.A(net407),
    .B(_12125_),
    .Y(_12394_));
 sg13g2_buf_2 _19327_ (.A(_12394_),
    .X(_12395_));
 sg13g2_nor2b_1 _19328_ (.A(_12395_),
    .B_N(\cpu.dcache.r_data[2][20] ),
    .Y(_12396_));
 sg13g2_a21oi_1 _19329_ (.A1(net986),
    .A2(_12395_),
    .Y(_12397_),
    .B1(_12396_));
 sg13g2_nand2_1 _19330_ (.Y(_12398_),
    .A(net987),
    .B(_12377_));
 sg13g2_o21ai_1 _19331_ (.B1(_12398_),
    .Y(_00396_),
    .A1(_12378_),
    .A2(_12397_));
 sg13g2_nor2b_1 _19332_ (.A(_12395_),
    .B_N(\cpu.dcache.r_data[2][21] ),
    .Y(_12399_));
 sg13g2_a21oi_1 _19333_ (.A1(net981),
    .A2(_12395_),
    .Y(_12400_),
    .B1(_12399_));
 sg13g2_nand2_1 _19334_ (.Y(_12401_),
    .A(net983),
    .B(_12377_));
 sg13g2_o21ai_1 _19335_ (.B1(_12401_),
    .Y(_00397_),
    .A1(net48),
    .A2(_12400_));
 sg13g2_nor2b_1 _19336_ (.A(_12395_),
    .B_N(\cpu.dcache.r_data[2][22] ),
    .Y(_12402_));
 sg13g2_a21oi_1 _19337_ (.A1(net985),
    .A2(_12395_),
    .Y(_12403_),
    .B1(_12402_));
 sg13g2_nand2_1 _19338_ (.Y(_12404_),
    .A(net982),
    .B(_12377_));
 sg13g2_o21ai_1 _19339_ (.B1(_12404_),
    .Y(_00398_),
    .A1(_12378_),
    .A2(_12403_));
 sg13g2_nor2b_1 _19340_ (.A(_12395_),
    .B_N(\cpu.dcache.r_data[2][23] ),
    .Y(_12405_));
 sg13g2_a21oi_1 _19341_ (.A1(net984),
    .A2(_12395_),
    .Y(_12406_),
    .B1(_12405_));
 sg13g2_nand2_1 _19342_ (.Y(_12407_),
    .A(net988),
    .B(_12377_));
 sg13g2_o21ai_1 _19343_ (.B1(_12407_),
    .Y(_00399_),
    .A1(net48),
    .A2(_12406_));
 sg13g2_nor2_1 _19344_ (.A(_12347_),
    .B(_12290_),
    .Y(_12408_));
 sg13g2_buf_1 _19345_ (.A(_12408_),
    .X(_12409_));
 sg13g2_buf_1 _19346_ (.A(_12409_),
    .X(_12410_));
 sg13g2_nor2_1 _19347_ (.A(_12346_),
    .B(net654),
    .Y(_12411_));
 sg13g2_buf_1 _19348_ (.A(_12411_),
    .X(_12412_));
 sg13g2_nor2b_1 _19349_ (.A(net367),
    .B_N(\cpu.dcache.r_data[2][24] ),
    .Y(_12413_));
 sg13g2_a21oi_1 _19350_ (.A1(_12255_),
    .A2(net367),
    .Y(_12414_),
    .B1(_12413_));
 sg13g2_nand2_1 _19351_ (.Y(_12415_),
    .A(net409),
    .B(net47));
 sg13g2_o21ai_1 _19352_ (.B1(_12415_),
    .Y(_00400_),
    .A1(net47),
    .A2(_12414_));
 sg13g2_nor2b_1 _19353_ (.A(net367),
    .B_N(\cpu.dcache.r_data[2][25] ),
    .Y(_12416_));
 sg13g2_a21oi_1 _19354_ (.A1(_12341_),
    .A2(net367),
    .Y(_12417_),
    .B1(_12416_));
 sg13g2_nand2_1 _19355_ (.Y(_12418_),
    .A(net372),
    .B(net47));
 sg13g2_o21ai_1 _19356_ (.B1(_12418_),
    .Y(_00401_),
    .A1(net47),
    .A2(_12417_));
 sg13g2_nor2b_1 _19357_ (.A(net367),
    .B_N(\cpu.dcache.r_data[2][26] ),
    .Y(_12419_));
 sg13g2_a21oi_1 _19358_ (.A1(_12263_),
    .A2(net367),
    .Y(_12420_),
    .B1(_12419_));
 sg13g2_nand2_1 _19359_ (.Y(_12421_),
    .A(net410),
    .B(_12409_));
 sg13g2_o21ai_1 _19360_ (.B1(_12421_),
    .Y(_00402_),
    .A1(net47),
    .A2(_12420_));
 sg13g2_nor2b_1 _19361_ (.A(_12412_),
    .B_N(\cpu.dcache.r_data[2][27] ),
    .Y(_12422_));
 sg13g2_a21oi_1 _19362_ (.A1(_12267_),
    .A2(_12412_),
    .Y(_12423_),
    .B1(_12422_));
 sg13g2_nand2_1 _19363_ (.Y(_12424_),
    .A(_12164_),
    .B(_12409_));
 sg13g2_o21ai_1 _19364_ (.B1(_12424_),
    .Y(_00403_),
    .A1(_12410_),
    .A2(_12423_));
 sg13g2_nor2_2 _19365_ (.A(net407),
    .B(_12167_),
    .Y(_12425_));
 sg13g2_mux2_1 _19366_ (.A0(\cpu.dcache.r_data[2][28] ),
    .A1(net1086),
    .S(_12425_),
    .X(_12426_));
 sg13g2_nor2_1 _19367_ (.A(_12409_),
    .B(_12426_),
    .Y(_12427_));
 sg13g2_a21oi_1 _19368_ (.A1(_12165_),
    .A2(net47),
    .Y(_00404_),
    .B1(_12427_));
 sg13g2_mux2_1 _19369_ (.A0(\cpu.dcache.r_data[2][29] ),
    .A1(net1083),
    .S(_12425_),
    .X(_12428_));
 sg13g2_nor2_1 _19370_ (.A(_12409_),
    .B(_12428_),
    .Y(_12429_));
 sg13g2_a21oi_1 _19371_ (.A1(net370),
    .A2(net47),
    .Y(_00405_),
    .B1(_12429_));
 sg13g2_nor2b_1 _19372_ (.A(_12352_),
    .B_N(\cpu.dcache.r_data[2][2] ),
    .Y(_12430_));
 sg13g2_a21oi_1 _19373_ (.A1(net985),
    .A2(_12352_),
    .Y(_12431_),
    .B1(_12430_));
 sg13g2_nand2_1 _19374_ (.Y(_12432_),
    .A(net852),
    .B(_12350_));
 sg13g2_o21ai_1 _19375_ (.B1(_12432_),
    .Y(_00406_),
    .A1(net50),
    .A2(_12431_));
 sg13g2_mux2_1 _19376_ (.A0(\cpu.dcache.r_data[2][30] ),
    .A1(net1085),
    .S(_12425_),
    .X(_12433_));
 sg13g2_nor2_1 _19377_ (.A(_12409_),
    .B(_12433_),
    .Y(_12434_));
 sg13g2_a21oi_1 _19378_ (.A1(_12178_),
    .A2(_12410_),
    .Y(_00407_),
    .B1(_12434_));
 sg13g2_mux2_1 _19379_ (.A0(\cpu.dcache.r_data[2][31] ),
    .A1(net1084),
    .S(_12425_),
    .X(_12435_));
 sg13g2_nor2_1 _19380_ (.A(_12409_),
    .B(_12435_),
    .Y(_12436_));
 sg13g2_a21oi_1 _19381_ (.A1(net368),
    .A2(net47),
    .Y(_00408_),
    .B1(_12436_));
 sg13g2_nor2b_1 _19382_ (.A(_12352_),
    .B_N(\cpu.dcache.r_data[2][3] ),
    .Y(_12437_));
 sg13g2_a21oi_1 _19383_ (.A1(net984),
    .A2(_12352_),
    .Y(_12438_),
    .B1(_12437_));
 sg13g2_nand2_1 _19384_ (.Y(_12439_),
    .A(net993),
    .B(_12349_));
 sg13g2_o21ai_1 _19385_ (.B1(_12439_),
    .Y(_00409_),
    .A1(net50),
    .A2(_12438_));
 sg13g2_nor2_1 _19386_ (.A(_12346_),
    .B(_12188_),
    .Y(_12440_));
 sg13g2_buf_2 _19387_ (.A(_12440_),
    .X(_12441_));
 sg13g2_nor2b_1 _19388_ (.A(_12441_),
    .B_N(\cpu.dcache.r_data[2][4] ),
    .Y(_12442_));
 sg13g2_a21oi_1 _19389_ (.A1(net986),
    .A2(_12441_),
    .Y(_12443_),
    .B1(_12442_));
 sg13g2_nand2_1 _19390_ (.Y(_12444_),
    .A(net987),
    .B(_12349_));
 sg13g2_o21ai_1 _19391_ (.B1(_12444_),
    .Y(_00410_),
    .A1(net50),
    .A2(_12443_));
 sg13g2_nor2b_1 _19392_ (.A(_12441_),
    .B_N(\cpu.dcache.r_data[2][5] ),
    .Y(_12445_));
 sg13g2_a21oi_1 _19393_ (.A1(net981),
    .A2(_12441_),
    .Y(_12446_),
    .B1(_12445_));
 sg13g2_nand2_1 _19394_ (.Y(_12447_),
    .A(net983),
    .B(_12349_));
 sg13g2_o21ai_1 _19395_ (.B1(_12447_),
    .Y(_00411_),
    .A1(net50),
    .A2(_12446_));
 sg13g2_buf_1 _19396_ (.A(net1093),
    .X(_12448_));
 sg13g2_nor2b_1 _19397_ (.A(_12441_),
    .B_N(\cpu.dcache.r_data[2][6] ),
    .Y(_12449_));
 sg13g2_a21oi_1 _19398_ (.A1(net980),
    .A2(_12441_),
    .Y(_12450_),
    .B1(_12449_));
 sg13g2_nand2_1 _19399_ (.Y(_12451_),
    .A(net982),
    .B(_12349_));
 sg13g2_o21ai_1 _19400_ (.B1(_12451_),
    .Y(_00412_),
    .A1(net50),
    .A2(_12450_));
 sg13g2_buf_1 _19401_ (.A(net1092),
    .X(_12452_));
 sg13g2_nor2b_1 _19402_ (.A(_12441_),
    .B_N(\cpu.dcache.r_data[2][7] ),
    .Y(_12453_));
 sg13g2_a21oi_1 _19403_ (.A1(net979),
    .A2(_12441_),
    .Y(_12454_),
    .B1(_12453_));
 sg13g2_nand2_1 _19404_ (.Y(_12455_),
    .A(net988),
    .B(_12349_));
 sg13g2_o21ai_1 _19405_ (.B1(_12455_),
    .Y(_00413_),
    .A1(net50),
    .A2(_12454_));
 sg13g2_buf_1 _19406_ (.A(net1095),
    .X(_12456_));
 sg13g2_nor2b_1 _19407_ (.A(_12360_),
    .B_N(\cpu.dcache.r_data[2][8] ),
    .Y(_12457_));
 sg13g2_a21oi_1 _19408_ (.A1(_12456_),
    .A2(_12360_),
    .Y(_12458_),
    .B1(_12457_));
 sg13g2_nand2_1 _19409_ (.Y(_12459_),
    .A(net409),
    .B(_12357_));
 sg13g2_o21ai_1 _19410_ (.B1(_12459_),
    .Y(_00414_),
    .A1(net49),
    .A2(_12458_));
 sg13g2_nor2b_1 _19411_ (.A(_12360_),
    .B_N(\cpu.dcache.r_data[2][9] ),
    .Y(_12460_));
 sg13g2_a21oi_1 _19412_ (.A1(net981),
    .A2(_12360_),
    .Y(_12461_),
    .B1(_12460_));
 sg13g2_nand2_1 _19413_ (.Y(_12462_),
    .A(net372),
    .B(_12357_));
 sg13g2_o21ai_1 _19414_ (.B1(_12462_),
    .Y(_00415_),
    .A1(net49),
    .A2(_12461_));
 sg13g2_nand2_1 _19415_ (.Y(_12463_),
    .A(net1119),
    .B(_09521_));
 sg13g2_buf_1 _19416_ (.A(_12463_),
    .X(_12464_));
 sg13g2_buf_1 _19417_ (.A(_12464_),
    .X(_12465_));
 sg13g2_nor2_1 _19418_ (.A(net528),
    .B(_12215_),
    .Y(_12466_));
 sg13g2_buf_1 _19419_ (.A(_12466_),
    .X(_12467_));
 sg13g2_nor2_1 _19420_ (.A(_12464_),
    .B(_12032_),
    .Y(_12468_));
 sg13g2_buf_2 _19421_ (.A(_12468_),
    .X(_12469_));
 sg13g2_nor2b_1 _19422_ (.A(_12469_),
    .B_N(\cpu.dcache.r_data[3][0] ),
    .Y(_12470_));
 sg13g2_a21oi_1 _19423_ (.A1(net978),
    .A2(_12469_),
    .Y(_12471_),
    .B1(_12470_));
 sg13g2_nand2_1 _19424_ (.Y(_12472_),
    .A(_12037_),
    .B(net66));
 sg13g2_o21ai_1 _19425_ (.B1(_12472_),
    .Y(_00416_),
    .A1(net66),
    .A2(_12471_));
 sg13g2_nor2_1 _19426_ (.A(net528),
    .B(_12225_),
    .Y(_12473_));
 sg13g2_buf_1 _19427_ (.A(_12473_),
    .X(_12474_));
 sg13g2_buf_1 _19428_ (.A(_12474_),
    .X(_12475_));
 sg13g2_nor2_1 _19429_ (.A(_12464_),
    .B(_12048_),
    .Y(_12476_));
 sg13g2_buf_2 _19430_ (.A(_12476_),
    .X(_12477_));
 sg13g2_nor2b_1 _19431_ (.A(_12477_),
    .B_N(\cpu.dcache.r_data[3][10] ),
    .Y(_12478_));
 sg13g2_a21oi_1 _19432_ (.A1(_12448_),
    .A2(_12477_),
    .Y(_12479_),
    .B1(_12478_));
 sg13g2_nand2_1 _19433_ (.Y(_12480_),
    .A(net410),
    .B(net46));
 sg13g2_o21ai_1 _19434_ (.B1(_12480_),
    .Y(_00417_),
    .A1(net46),
    .A2(_12479_));
 sg13g2_nor2b_1 _19435_ (.A(_12477_),
    .B_N(\cpu.dcache.r_data[3][11] ),
    .Y(_12481_));
 sg13g2_a21oi_1 _19436_ (.A1(net979),
    .A2(_12477_),
    .Y(_12482_),
    .B1(_12481_));
 sg13g2_nand2_1 _19437_ (.Y(_12483_),
    .A(net408),
    .B(net46));
 sg13g2_o21ai_1 _19438_ (.B1(_12483_),
    .Y(_00418_),
    .A1(net46),
    .A2(_12482_));
 sg13g2_nor2_2 _19439_ (.A(net528),
    .B(_12076_),
    .Y(_12484_));
 sg13g2_mux2_1 _19440_ (.A0(\cpu.dcache.r_data[3][12] ),
    .A1(net1086),
    .S(_12484_),
    .X(_12485_));
 sg13g2_nor2_1 _19441_ (.A(_12474_),
    .B(_12485_),
    .Y(_12486_));
 sg13g2_a21oi_1 _19442_ (.A1(net371),
    .A2(net46),
    .Y(_00419_),
    .B1(_12486_));
 sg13g2_mux2_1 _19443_ (.A0(\cpu.dcache.r_data[3][13] ),
    .A1(_12271_),
    .S(_12484_),
    .X(_12487_));
 sg13g2_nor2_1 _19444_ (.A(_12474_),
    .B(_12487_),
    .Y(_12488_));
 sg13g2_a21oi_1 _19445_ (.A1(net370),
    .A2(net46),
    .Y(_00420_),
    .B1(_12488_));
 sg13g2_mux2_1 _19446_ (.A0(\cpu.dcache.r_data[3][14] ),
    .A1(_12243_),
    .S(_12484_),
    .X(_12489_));
 sg13g2_nor2_1 _19447_ (.A(_12474_),
    .B(_12489_),
    .Y(_12490_));
 sg13g2_a21oi_1 _19448_ (.A1(net369),
    .A2(_12475_),
    .Y(_00421_),
    .B1(_12490_));
 sg13g2_mux2_1 _19449_ (.A0(\cpu.dcache.r_data[3][15] ),
    .A1(net1084),
    .S(_12484_),
    .X(_12491_));
 sg13g2_nor2_1 _19450_ (.A(_12474_),
    .B(_12491_),
    .Y(_12492_));
 sg13g2_a21oi_1 _19451_ (.A1(net368),
    .A2(_12475_),
    .Y(_00422_),
    .B1(_12492_));
 sg13g2_nor2_1 _19452_ (.A(net528),
    .B(_12251_),
    .Y(_12493_));
 sg13g2_buf_1 _19453_ (.A(_12493_),
    .X(_12494_));
 sg13g2_nor2_1 _19454_ (.A(_12464_),
    .B(_12105_),
    .Y(_12495_));
 sg13g2_buf_2 _19455_ (.A(_12495_),
    .X(_12496_));
 sg13g2_nor2b_1 _19456_ (.A(_12496_),
    .B_N(\cpu.dcache.r_data[3][16] ),
    .Y(_12497_));
 sg13g2_a21oi_1 _19457_ (.A1(net978),
    .A2(_12496_),
    .Y(_12498_),
    .B1(_12497_));
 sg13g2_nand2_1 _19458_ (.Y(_12499_),
    .A(net853),
    .B(net65));
 sg13g2_o21ai_1 _19459_ (.B1(_12499_),
    .Y(_00423_),
    .A1(net65),
    .A2(_12498_));
 sg13g2_mux2_1 _19460_ (.A0(\cpu.dcache.r_data[3][17] ),
    .A1(net1083),
    .S(_12496_),
    .X(_12500_));
 sg13g2_nor2_1 _19461_ (.A(_12493_),
    .B(_12500_),
    .Y(_12501_));
 sg13g2_a21oi_1 _19462_ (.A1(_12111_),
    .A2(net65),
    .Y(_00424_),
    .B1(_12501_));
 sg13g2_nor2b_1 _19463_ (.A(_12496_),
    .B_N(\cpu.dcache.r_data[3][18] ),
    .Y(_12502_));
 sg13g2_a21oi_1 _19464_ (.A1(net980),
    .A2(_12496_),
    .Y(_12503_),
    .B1(_12502_));
 sg13g2_nand2_1 _19465_ (.Y(_12504_),
    .A(_12176_),
    .B(net65));
 sg13g2_o21ai_1 _19466_ (.B1(_12504_),
    .Y(_00425_),
    .A1(_12494_),
    .A2(_12503_));
 sg13g2_nor2b_1 _19467_ (.A(_12496_),
    .B_N(\cpu.dcache.r_data[3][19] ),
    .Y(_12505_));
 sg13g2_a21oi_1 _19468_ (.A1(net979),
    .A2(_12496_),
    .Y(_12506_),
    .B1(_12505_));
 sg13g2_nand2_1 _19469_ (.Y(_12507_),
    .A(_12119_),
    .B(_12493_));
 sg13g2_o21ai_1 _19470_ (.B1(_12507_),
    .Y(_00426_),
    .A1(_12494_),
    .A2(_12506_));
 sg13g2_mux2_1 _19471_ (.A0(\cpu.dcache.r_data[3][1] ),
    .A1(net1083),
    .S(_12469_),
    .X(_12508_));
 sg13g2_nor2_1 _19472_ (.A(_12466_),
    .B(_12508_),
    .Y(_12509_));
 sg13g2_a21oi_1 _19473_ (.A1(net731),
    .A2(net66),
    .Y(_00427_),
    .B1(_12509_));
 sg13g2_or2_1 _19474_ (.X(_12510_),
    .B(_12125_),
    .A(net528));
 sg13g2_buf_1 _19475_ (.A(_12510_),
    .X(_12511_));
 sg13g2_mux2_1 _19476_ (.A0(net1091),
    .A1(\cpu.dcache.r_data[3][20] ),
    .S(_12511_),
    .X(_12512_));
 sg13g2_mux2_1 _19477_ (.A0(_12512_),
    .A1(_10152_),
    .S(net65),
    .X(_00428_));
 sg13g2_mux2_1 _19478_ (.A0(_12156_),
    .A1(\cpu.dcache.r_data[3][21] ),
    .S(_12511_),
    .X(_12513_));
 sg13g2_mux2_1 _19479_ (.A0(_12513_),
    .A1(_10158_),
    .S(net65),
    .X(_00429_));
 sg13g2_mux2_1 _19480_ (.A0(net1089),
    .A1(\cpu.dcache.r_data[3][22] ),
    .S(_12511_),
    .X(_12514_));
 sg13g2_mux2_1 _19481_ (.A0(_12514_),
    .A1(_10164_),
    .S(net65),
    .X(_00430_));
 sg13g2_mux2_1 _19482_ (.A0(net1088),
    .A1(\cpu.dcache.r_data[3][23] ),
    .S(_12511_),
    .X(_12515_));
 sg13g2_buf_1 _19483_ (.A(net1021),
    .X(_12516_));
 sg13g2_mux2_1 _19484_ (.A0(_12515_),
    .A1(net851),
    .S(net65),
    .X(_00431_));
 sg13g2_nor2_1 _19485_ (.A(_12465_),
    .B(_12290_),
    .Y(_12517_));
 sg13g2_buf_1 _19486_ (.A(_12517_),
    .X(_12518_));
 sg13g2_buf_1 _19487_ (.A(_12518_),
    .X(_12519_));
 sg13g2_nor2_1 _19488_ (.A(_12464_),
    .B(net654),
    .Y(_12520_));
 sg13g2_buf_1 _19489_ (.A(_12520_),
    .X(_12521_));
 sg13g2_nor2b_1 _19490_ (.A(net468),
    .B_N(\cpu.dcache.r_data[3][24] ),
    .Y(_12522_));
 sg13g2_a21oi_1 _19491_ (.A1(_12456_),
    .A2(net468),
    .Y(_12523_),
    .B1(_12522_));
 sg13g2_nand2_1 _19492_ (.Y(_12524_),
    .A(_12151_),
    .B(net45));
 sg13g2_o21ai_1 _19493_ (.B1(_12524_),
    .Y(_00432_),
    .A1(net45),
    .A2(_12523_));
 sg13g2_nor2b_1 _19494_ (.A(net468),
    .B_N(\cpu.dcache.r_data[3][25] ),
    .Y(_12525_));
 sg13g2_a21oi_1 _19495_ (.A1(_12341_),
    .A2(net468),
    .Y(_12526_),
    .B1(_12525_));
 sg13g2_nand2_1 _19496_ (.Y(_12527_),
    .A(net372),
    .B(net45));
 sg13g2_o21ai_1 _19497_ (.B1(_12527_),
    .Y(_00433_),
    .A1(net45),
    .A2(_12526_));
 sg13g2_nor2b_1 _19498_ (.A(net468),
    .B_N(\cpu.dcache.r_data[3][26] ),
    .Y(_12528_));
 sg13g2_a21oi_1 _19499_ (.A1(_12448_),
    .A2(net468),
    .Y(_12529_),
    .B1(_12528_));
 sg13g2_nand2_1 _19500_ (.Y(_12530_),
    .A(net410),
    .B(_12518_));
 sg13g2_o21ai_1 _19501_ (.B1(_12530_),
    .Y(_00434_),
    .A1(_12519_),
    .A2(_12529_));
 sg13g2_nor2b_1 _19502_ (.A(net468),
    .B_N(\cpu.dcache.r_data[3][27] ),
    .Y(_12531_));
 sg13g2_a21oi_1 _19503_ (.A1(_12452_),
    .A2(net468),
    .Y(_12532_),
    .B1(_12531_));
 sg13g2_nand2_1 _19504_ (.Y(_12533_),
    .A(_12164_),
    .B(_12518_));
 sg13g2_o21ai_1 _19505_ (.B1(_12533_),
    .Y(_00435_),
    .A1(_12519_),
    .A2(_12532_));
 sg13g2_nor2_2 _19506_ (.A(_12465_),
    .B(_12167_),
    .Y(_12534_));
 sg13g2_mux2_1 _19507_ (.A0(\cpu.dcache.r_data[3][28] ),
    .A1(net1086),
    .S(_12534_),
    .X(_12535_));
 sg13g2_nor2_1 _19508_ (.A(_12518_),
    .B(_12535_),
    .Y(_12536_));
 sg13g2_a21oi_1 _19509_ (.A1(_12165_),
    .A2(net45),
    .Y(_00436_),
    .B1(_12536_));
 sg13g2_mux2_1 _19510_ (.A0(\cpu.dcache.r_data[3][29] ),
    .A1(_12271_),
    .S(_12534_),
    .X(_12537_));
 sg13g2_nor2_1 _19511_ (.A(_12518_),
    .B(_12537_),
    .Y(_12538_));
 sg13g2_a21oi_1 _19512_ (.A1(net370),
    .A2(net45),
    .Y(_00437_),
    .B1(_12538_));
 sg13g2_nor2b_1 _19513_ (.A(_12469_),
    .B_N(\cpu.dcache.r_data[3][2] ),
    .Y(_12539_));
 sg13g2_a21oi_1 _19514_ (.A1(net980),
    .A2(_12469_),
    .Y(_12540_),
    .B1(_12539_));
 sg13g2_nand2_1 _19515_ (.Y(_12541_),
    .A(net852),
    .B(net66));
 sg13g2_o21ai_1 _19516_ (.B1(_12541_),
    .Y(_00438_),
    .A1(_12467_),
    .A2(_12540_));
 sg13g2_mux2_1 _19517_ (.A0(\cpu.dcache.r_data[3][30] ),
    .A1(net1085),
    .S(_12534_),
    .X(_12542_));
 sg13g2_nor2_1 _19518_ (.A(_12518_),
    .B(_12542_),
    .Y(_12543_));
 sg13g2_a21oi_1 _19519_ (.A1(_12178_),
    .A2(net45),
    .Y(_00439_),
    .B1(_12543_));
 sg13g2_mux2_1 _19520_ (.A0(\cpu.dcache.r_data[3][31] ),
    .A1(net1084),
    .S(_12534_),
    .X(_12544_));
 sg13g2_nor2_1 _19521_ (.A(_12518_),
    .B(_12544_),
    .Y(_12545_));
 sg13g2_a21oi_1 _19522_ (.A1(net368),
    .A2(net45),
    .Y(_00440_),
    .B1(_12545_));
 sg13g2_nor2b_1 _19523_ (.A(_12469_),
    .B_N(\cpu.dcache.r_data[3][3] ),
    .Y(_12546_));
 sg13g2_a21oi_1 _19524_ (.A1(net979),
    .A2(_12469_),
    .Y(_12547_),
    .B1(_12546_));
 sg13g2_nand2_1 _19525_ (.Y(_12548_),
    .A(net993),
    .B(_12466_));
 sg13g2_o21ai_1 _19526_ (.B1(_12548_),
    .Y(_00441_),
    .A1(_12467_),
    .A2(_12547_));
 sg13g2_or2_1 _19527_ (.X(_12549_),
    .B(_12188_),
    .A(net528));
 sg13g2_buf_1 _19528_ (.A(_12549_),
    .X(_12550_));
 sg13g2_mux2_1 _19529_ (.A0(net1091),
    .A1(\cpu.dcache.r_data[3][4] ),
    .S(_12550_),
    .X(_12551_));
 sg13g2_mux2_1 _19530_ (.A0(_12551_),
    .A1(net992),
    .S(net66),
    .X(_00442_));
 sg13g2_mux2_1 _19531_ (.A0(net1090),
    .A1(\cpu.dcache.r_data[3][5] ),
    .S(_12550_),
    .X(_12552_));
 sg13g2_mux2_1 _19532_ (.A0(_12552_),
    .A1(net990),
    .S(net66),
    .X(_00443_));
 sg13g2_mux2_1 _19533_ (.A0(net1089),
    .A1(\cpu.dcache.r_data[3][6] ),
    .S(_12550_),
    .X(_12553_));
 sg13g2_mux2_1 _19534_ (.A0(_12553_),
    .A1(net882),
    .S(net66),
    .X(_00444_));
 sg13g2_mux2_1 _19535_ (.A0(net1088),
    .A1(\cpu.dcache.r_data[3][7] ),
    .S(_12550_),
    .X(_12554_));
 sg13g2_mux2_1 _19536_ (.A0(_12554_),
    .A1(_12516_),
    .S(net66),
    .X(_00445_));
 sg13g2_nor2b_1 _19537_ (.A(_12477_),
    .B_N(\cpu.dcache.r_data[3][8] ),
    .Y(_12555_));
 sg13g2_a21oi_1 _19538_ (.A1(net978),
    .A2(_12477_),
    .Y(_12556_),
    .B1(_12555_));
 sg13g2_nand2_1 _19539_ (.Y(_12557_),
    .A(net409),
    .B(_12474_));
 sg13g2_o21ai_1 _19540_ (.B1(_12557_),
    .Y(_00446_),
    .A1(net46),
    .A2(_12556_));
 sg13g2_nor2b_1 _19541_ (.A(_12477_),
    .B_N(\cpu.dcache.r_data[3][9] ),
    .Y(_12558_));
 sg13g2_a21oi_1 _19542_ (.A1(net981),
    .A2(_12477_),
    .Y(_12559_),
    .B1(_12558_));
 sg13g2_nand2_1 _19543_ (.Y(_12560_),
    .A(_12161_),
    .B(_12474_));
 sg13g2_o21ai_1 _19544_ (.B1(_12560_),
    .Y(_00447_),
    .A1(net46),
    .A2(_12559_));
 sg13g2_buf_1 _19545_ (.A(_10110_),
    .X(_12561_));
 sg13g2_nor2_1 _19546_ (.A(net600),
    .B(_12215_),
    .Y(_12562_));
 sg13g2_buf_2 _19547_ (.A(_12562_),
    .X(_12563_));
 sg13g2_buf_1 _19548_ (.A(_12563_),
    .X(_12564_));
 sg13g2_nor2_1 _19549_ (.A(_10110_),
    .B(_12032_),
    .Y(_12565_));
 sg13g2_buf_2 _19550_ (.A(_12565_),
    .X(_12566_));
 sg13g2_nor2b_1 _19551_ (.A(_12566_),
    .B_N(\cpu.dcache.r_data[4][0] ),
    .Y(_12567_));
 sg13g2_a21oi_1 _19552_ (.A1(net978),
    .A2(_12566_),
    .Y(_12568_),
    .B1(_12567_));
 sg13g2_nand2_1 _19553_ (.Y(_12569_),
    .A(net853),
    .B(_12564_));
 sg13g2_o21ai_1 _19554_ (.B1(_12569_),
    .Y(_00448_),
    .A1(_12564_),
    .A2(_12568_));
 sg13g2_nor2_1 _19555_ (.A(_12561_),
    .B(_12225_),
    .Y(_12570_));
 sg13g2_buf_1 _19556_ (.A(_12570_),
    .X(_12571_));
 sg13g2_buf_1 _19557_ (.A(_12571_),
    .X(_12572_));
 sg13g2_nor2_1 _19558_ (.A(net600),
    .B(_12048_),
    .Y(_12573_));
 sg13g2_buf_2 _19559_ (.A(_12573_),
    .X(_12574_));
 sg13g2_nor2b_1 _19560_ (.A(_12574_),
    .B_N(\cpu.dcache.r_data[4][10] ),
    .Y(_12575_));
 sg13g2_a21oi_1 _19561_ (.A1(net980),
    .A2(_12574_),
    .Y(_12576_),
    .B1(_12575_));
 sg13g2_nand2_1 _19562_ (.Y(_12577_),
    .A(net410),
    .B(net43));
 sg13g2_o21ai_1 _19563_ (.B1(_12577_),
    .Y(_00449_),
    .A1(net43),
    .A2(_12576_));
 sg13g2_nor2b_1 _19564_ (.A(_12574_),
    .B_N(\cpu.dcache.r_data[4][11] ),
    .Y(_12578_));
 sg13g2_a21oi_1 _19565_ (.A1(_12452_),
    .A2(_12574_),
    .Y(_12579_),
    .B1(_12578_));
 sg13g2_nand2_1 _19566_ (.Y(_12580_),
    .A(net408),
    .B(net43));
 sg13g2_o21ai_1 _19567_ (.B1(_12580_),
    .Y(_00450_),
    .A1(net43),
    .A2(_12579_));
 sg13g2_nor2_2 _19568_ (.A(net600),
    .B(_12076_),
    .Y(_12581_));
 sg13g2_mux2_1 _19569_ (.A0(\cpu.dcache.r_data[4][12] ),
    .A1(net1086),
    .S(_12581_),
    .X(_12582_));
 sg13g2_nor2_1 _19570_ (.A(_12571_),
    .B(_12582_),
    .Y(_12583_));
 sg13g2_a21oi_1 _19571_ (.A1(net371),
    .A2(net43),
    .Y(_00451_),
    .B1(_12583_));
 sg13g2_buf_1 _19572_ (.A(_12083_),
    .X(_12584_));
 sg13g2_mux2_1 _19573_ (.A0(\cpu.dcache.r_data[4][13] ),
    .A1(net1082),
    .S(_12581_),
    .X(_12585_));
 sg13g2_nor2_1 _19574_ (.A(_12571_),
    .B(_12585_),
    .Y(_12586_));
 sg13g2_a21oi_1 _19575_ (.A1(net370),
    .A2(net43),
    .Y(_00452_),
    .B1(_12586_));
 sg13g2_mux2_1 _19576_ (.A0(\cpu.dcache.r_data[4][14] ),
    .A1(_12243_),
    .S(_12581_),
    .X(_12587_));
 sg13g2_nor2_1 _19577_ (.A(_12571_),
    .B(_12587_),
    .Y(_12588_));
 sg13g2_a21oi_1 _19578_ (.A1(net369),
    .A2(_12572_),
    .Y(_00453_),
    .B1(_12588_));
 sg13g2_mux2_1 _19579_ (.A0(\cpu.dcache.r_data[4][15] ),
    .A1(net1084),
    .S(_12581_),
    .X(_12589_));
 sg13g2_nor2_1 _19580_ (.A(_12571_),
    .B(_12589_),
    .Y(_12590_));
 sg13g2_a21oi_1 _19581_ (.A1(net368),
    .A2(_12572_),
    .Y(_00454_),
    .B1(_12590_));
 sg13g2_nor2_1 _19582_ (.A(net600),
    .B(_12251_),
    .Y(_12591_));
 sg13g2_buf_2 _19583_ (.A(_12591_),
    .X(_12592_));
 sg13g2_buf_1 _19584_ (.A(_12592_),
    .X(_12593_));
 sg13g2_nor2_1 _19585_ (.A(_10110_),
    .B(_12105_),
    .Y(_12594_));
 sg13g2_buf_2 _19586_ (.A(_12594_),
    .X(_12595_));
 sg13g2_nor2b_1 _19587_ (.A(_12595_),
    .B_N(\cpu.dcache.r_data[4][16] ),
    .Y(_12596_));
 sg13g2_a21oi_1 _19588_ (.A1(net978),
    .A2(_12595_),
    .Y(_12597_),
    .B1(_12596_));
 sg13g2_nand2_1 _19589_ (.Y(_12598_),
    .A(_12037_),
    .B(net42));
 sg13g2_o21ai_1 _19590_ (.B1(_12598_),
    .Y(_00455_),
    .A1(net42),
    .A2(_12597_));
 sg13g2_mux2_1 _19591_ (.A0(\cpu.dcache.r_data[4][17] ),
    .A1(net1082),
    .S(_12595_),
    .X(_12599_));
 sg13g2_nor2_1 _19592_ (.A(_12592_),
    .B(_12599_),
    .Y(_12600_));
 sg13g2_a21oi_1 _19593_ (.A1(_12111_),
    .A2(net42),
    .Y(_00456_),
    .B1(_12600_));
 sg13g2_nor2b_1 _19594_ (.A(_12595_),
    .B_N(\cpu.dcache.r_data[4][18] ),
    .Y(_12601_));
 sg13g2_a21oi_1 _19595_ (.A1(net980),
    .A2(_12595_),
    .Y(_12602_),
    .B1(_12601_));
 sg13g2_nand2_1 _19596_ (.Y(_12603_),
    .A(_12176_),
    .B(net42));
 sg13g2_o21ai_1 _19597_ (.B1(_12603_),
    .Y(_00457_),
    .A1(net42),
    .A2(_12602_));
 sg13g2_nor2b_1 _19598_ (.A(_12595_),
    .B_N(\cpu.dcache.r_data[4][19] ),
    .Y(_12604_));
 sg13g2_a21oi_1 _19599_ (.A1(net979),
    .A2(_12595_),
    .Y(_12605_),
    .B1(_12604_));
 sg13g2_nand2_1 _19600_ (.Y(_12606_),
    .A(_12119_),
    .B(_12592_));
 sg13g2_o21ai_1 _19601_ (.B1(_12606_),
    .Y(_00458_),
    .A1(net42),
    .A2(_12605_));
 sg13g2_mux2_1 _19602_ (.A0(\cpu.dcache.r_data[4][1] ),
    .A1(net1082),
    .S(_12566_),
    .X(_12607_));
 sg13g2_nor2_1 _19603_ (.A(_12563_),
    .B(_12607_),
    .Y(_12608_));
 sg13g2_a21oi_1 _19604_ (.A1(net731),
    .A2(net44),
    .Y(_00459_),
    .B1(_12608_));
 sg13g2_nor2_1 _19605_ (.A(net600),
    .B(_12125_),
    .Y(_12609_));
 sg13g2_buf_2 _19606_ (.A(_12609_),
    .X(_12610_));
 sg13g2_nor2b_1 _19607_ (.A(_12610_),
    .B_N(\cpu.dcache.r_data[4][20] ),
    .Y(_12611_));
 sg13g2_a21oi_1 _19608_ (.A1(net978),
    .A2(_12610_),
    .Y(_12612_),
    .B1(_12611_));
 sg13g2_nand2_1 _19609_ (.Y(_12613_),
    .A(net987),
    .B(_12592_));
 sg13g2_o21ai_1 _19610_ (.B1(_12613_),
    .Y(_00460_),
    .A1(net42),
    .A2(_12612_));
 sg13g2_nor2b_1 _19611_ (.A(_12610_),
    .B_N(\cpu.dcache.r_data[4][21] ),
    .Y(_12614_));
 sg13g2_a21oi_1 _19612_ (.A1(net981),
    .A2(_12610_),
    .Y(_12615_),
    .B1(_12614_));
 sg13g2_nand2_1 _19613_ (.Y(_12616_),
    .A(net983),
    .B(_12592_));
 sg13g2_o21ai_1 _19614_ (.B1(_12616_),
    .Y(_00461_),
    .A1(net42),
    .A2(_12615_));
 sg13g2_nor2b_1 _19615_ (.A(_12610_),
    .B_N(\cpu.dcache.r_data[4][22] ),
    .Y(_12617_));
 sg13g2_a21oi_1 _19616_ (.A1(net980),
    .A2(_12610_),
    .Y(_12618_),
    .B1(_12617_));
 sg13g2_nand2_1 _19617_ (.Y(_12619_),
    .A(net982),
    .B(_12592_));
 sg13g2_o21ai_1 _19618_ (.B1(_12619_),
    .Y(_00462_),
    .A1(_12593_),
    .A2(_12618_));
 sg13g2_nor2b_1 _19619_ (.A(_12610_),
    .B_N(\cpu.dcache.r_data[4][23] ),
    .Y(_12620_));
 sg13g2_a21oi_1 _19620_ (.A1(net979),
    .A2(_12610_),
    .Y(_12621_),
    .B1(_12620_));
 sg13g2_nand2_1 _19621_ (.Y(_12622_),
    .A(net988),
    .B(_12592_));
 sg13g2_o21ai_1 _19622_ (.B1(_12622_),
    .Y(_00463_),
    .A1(_12593_),
    .A2(_12621_));
 sg13g2_or2_1 _19623_ (.X(_12623_),
    .B(net654),
    .A(_10110_));
 sg13g2_buf_1 _19624_ (.A(_12623_),
    .X(_12624_));
 sg13g2_mux2_1 _19625_ (.A0(net1091),
    .A1(\cpu.dcache.r_data[4][24] ),
    .S(net527),
    .X(_12625_));
 sg13g2_nor2_1 _19626_ (.A(net600),
    .B(_12290_),
    .Y(_12626_));
 sg13g2_buf_1 _19627_ (.A(_12626_),
    .X(_12627_));
 sg13g2_mux2_1 _19628_ (.A0(_12625_),
    .A1(net409),
    .S(net64),
    .X(_00464_));
 sg13g2_mux2_1 _19629_ (.A0(_12084_),
    .A1(\cpu.dcache.r_data[4][25] ),
    .S(net527),
    .X(_12628_));
 sg13g2_mux2_1 _19630_ (.A0(_12628_),
    .A1(net372),
    .S(net64),
    .X(_00465_));
 sg13g2_mux2_1 _19631_ (.A0(net1089),
    .A1(\cpu.dcache.r_data[4][26] ),
    .S(net527),
    .X(_12629_));
 sg13g2_mux2_1 _19632_ (.A0(_12629_),
    .A1(_12059_),
    .S(net64),
    .X(_00466_));
 sg13g2_mux2_1 _19633_ (.A0(net1088),
    .A1(\cpu.dcache.r_data[4][27] ),
    .S(net527),
    .X(_12630_));
 sg13g2_mux2_1 _19634_ (.A0(_12630_),
    .A1(net408),
    .S(net64),
    .X(_00467_));
 sg13g2_nor2_2 _19635_ (.A(_12561_),
    .B(_12167_),
    .Y(_12631_));
 sg13g2_mux2_1 _19636_ (.A0(\cpu.dcache.r_data[4][28] ),
    .A1(_12237_),
    .S(_12631_),
    .X(_12632_));
 sg13g2_nor2_1 _19637_ (.A(net64),
    .B(_12632_),
    .Y(_12633_));
 sg13g2_a21oi_1 _19638_ (.A1(net371),
    .A2(net64),
    .Y(_00468_),
    .B1(_12633_));
 sg13g2_mux2_1 _19639_ (.A0(\cpu.dcache.r_data[4][29] ),
    .A1(net1082),
    .S(_12631_),
    .X(_12634_));
 sg13g2_nor2_1 _19640_ (.A(net64),
    .B(_12634_),
    .Y(_12635_));
 sg13g2_a21oi_1 _19641_ (.A1(_12171_),
    .A2(net64),
    .Y(_00469_),
    .B1(_12635_));
 sg13g2_nor2b_1 _19642_ (.A(_12566_),
    .B_N(\cpu.dcache.r_data[4][2] ),
    .Y(_12636_));
 sg13g2_a21oi_1 _19643_ (.A1(net980),
    .A2(_12566_),
    .Y(_12637_),
    .B1(_12636_));
 sg13g2_nand2_1 _19644_ (.Y(_12638_),
    .A(net852),
    .B(net44));
 sg13g2_o21ai_1 _19645_ (.B1(_12638_),
    .Y(_00470_),
    .A1(net44),
    .A2(_12637_));
 sg13g2_mux2_1 _19646_ (.A0(\cpu.dcache.r_data[4][30] ),
    .A1(net1085),
    .S(_12631_),
    .X(_12639_));
 sg13g2_nor2_1 _19647_ (.A(_12626_),
    .B(_12639_),
    .Y(_12640_));
 sg13g2_a21oi_1 _19648_ (.A1(net369),
    .A2(_12627_),
    .Y(_00471_),
    .B1(_12640_));
 sg13g2_mux2_1 _19649_ (.A0(\cpu.dcache.r_data[4][31] ),
    .A1(_12246_),
    .S(_12631_),
    .X(_12641_));
 sg13g2_nor2_1 _19650_ (.A(_12626_),
    .B(_12641_),
    .Y(_12642_));
 sg13g2_a21oi_1 _19651_ (.A1(_12181_),
    .A2(_12627_),
    .Y(_00472_),
    .B1(_12642_));
 sg13g2_nor2b_1 _19652_ (.A(_12566_),
    .B_N(\cpu.dcache.r_data[4][3] ),
    .Y(_12643_));
 sg13g2_a21oi_1 _19653_ (.A1(net979),
    .A2(_12566_),
    .Y(_12644_),
    .B1(_12643_));
 sg13g2_nand2_1 _19654_ (.Y(_12645_),
    .A(net993),
    .B(_12563_));
 sg13g2_o21ai_1 _19655_ (.B1(_12645_),
    .Y(_00473_),
    .A1(net44),
    .A2(_12644_));
 sg13g2_nor2_1 _19656_ (.A(net600),
    .B(_12188_),
    .Y(_12646_));
 sg13g2_buf_2 _19657_ (.A(_12646_),
    .X(_12647_));
 sg13g2_nor2b_1 _19658_ (.A(_12647_),
    .B_N(\cpu.dcache.r_data[4][4] ),
    .Y(_12648_));
 sg13g2_a21oi_1 _19659_ (.A1(net978),
    .A2(_12647_),
    .Y(_12649_),
    .B1(_12648_));
 sg13g2_nand2_1 _19660_ (.Y(_12650_),
    .A(net987),
    .B(_12563_));
 sg13g2_o21ai_1 _19661_ (.B1(_12650_),
    .Y(_00474_),
    .A1(net44),
    .A2(_12649_));
 sg13g2_nor2b_1 _19662_ (.A(_12647_),
    .B_N(\cpu.dcache.r_data[4][5] ),
    .Y(_12651_));
 sg13g2_a21oi_1 _19663_ (.A1(net981),
    .A2(_12647_),
    .Y(_12652_),
    .B1(_12651_));
 sg13g2_nand2_1 _19664_ (.Y(_12653_),
    .A(net983),
    .B(_12563_));
 sg13g2_o21ai_1 _19665_ (.B1(_12653_),
    .Y(_00475_),
    .A1(net44),
    .A2(_12652_));
 sg13g2_nor2b_1 _19666_ (.A(_12647_),
    .B_N(\cpu.dcache.r_data[4][6] ),
    .Y(_12654_));
 sg13g2_a21oi_1 _19667_ (.A1(net980),
    .A2(_12647_),
    .Y(_12655_),
    .B1(_12654_));
 sg13g2_nand2_1 _19668_ (.Y(_12656_),
    .A(net982),
    .B(_12563_));
 sg13g2_o21ai_1 _19669_ (.B1(_12656_),
    .Y(_00476_),
    .A1(net44),
    .A2(_12655_));
 sg13g2_nor2b_1 _19670_ (.A(_12647_),
    .B_N(\cpu.dcache.r_data[4][7] ),
    .Y(_12657_));
 sg13g2_a21oi_1 _19671_ (.A1(net979),
    .A2(_12647_),
    .Y(_12658_),
    .B1(_12657_));
 sg13g2_nand2_1 _19672_ (.Y(_12659_),
    .A(net988),
    .B(_12563_));
 sg13g2_o21ai_1 _19673_ (.B1(_12659_),
    .Y(_00477_),
    .A1(net44),
    .A2(_12658_));
 sg13g2_nor2b_1 _19674_ (.A(_12574_),
    .B_N(\cpu.dcache.r_data[4][8] ),
    .Y(_12660_));
 sg13g2_a21oi_1 _19675_ (.A1(net978),
    .A2(_12574_),
    .Y(_12661_),
    .B1(_12660_));
 sg13g2_nand2_1 _19676_ (.Y(_12662_),
    .A(_12151_),
    .B(_12571_));
 sg13g2_o21ai_1 _19677_ (.B1(_12662_),
    .Y(_00478_),
    .A1(net43),
    .A2(_12661_));
 sg13g2_nor2b_1 _19678_ (.A(_12574_),
    .B_N(\cpu.dcache.r_data[4][9] ),
    .Y(_12663_));
 sg13g2_a21oi_1 _19679_ (.A1(net981),
    .A2(_12574_),
    .Y(_12664_),
    .B1(_12663_));
 sg13g2_nand2_1 _19680_ (.Y(_12665_),
    .A(_12161_),
    .B(_12571_));
 sg13g2_o21ai_1 _19681_ (.B1(_12665_),
    .Y(_00479_),
    .A1(net43),
    .A2(_12664_));
 sg13g2_nand2_1 _19682_ (.Y(_12666_),
    .A(net894),
    .B(_09421_));
 sg13g2_buf_1 _19683_ (.A(_12666_),
    .X(_12667_));
 sg13g2_buf_1 _19684_ (.A(net653),
    .X(_12668_));
 sg13g2_nor2_1 _19685_ (.A(net599),
    .B(_12215_),
    .Y(_12669_));
 sg13g2_buf_2 _19686_ (.A(_12669_),
    .X(_12670_));
 sg13g2_buf_1 _19687_ (.A(_12670_),
    .X(_12671_));
 sg13g2_buf_1 _19688_ (.A(_12022_),
    .X(_12672_));
 sg13g2_nor2_1 _19689_ (.A(net653),
    .B(_12032_),
    .Y(_12673_));
 sg13g2_buf_2 _19690_ (.A(_12673_),
    .X(_12674_));
 sg13g2_nor2b_1 _19691_ (.A(_12674_),
    .B_N(\cpu.dcache.r_data[5][0] ),
    .Y(_12675_));
 sg13g2_a21oi_1 _19692_ (.A1(net977),
    .A2(_12674_),
    .Y(_12676_),
    .B1(_12675_));
 sg13g2_buf_1 _19693_ (.A(net1029),
    .X(_12677_));
 sg13g2_nand2_1 _19694_ (.Y(_12678_),
    .A(net850),
    .B(net41));
 sg13g2_o21ai_1 _19695_ (.B1(_12678_),
    .Y(_00480_),
    .A1(net41),
    .A2(_12676_));
 sg13g2_nor2_1 _19696_ (.A(_12668_),
    .B(_12225_),
    .Y(_12679_));
 sg13g2_buf_2 _19697_ (.A(_12679_),
    .X(_12680_));
 sg13g2_buf_1 _19698_ (.A(_12680_),
    .X(_12681_));
 sg13g2_buf_1 _19699_ (.A(net1093),
    .X(_12682_));
 sg13g2_nor2_1 _19700_ (.A(net599),
    .B(_12048_),
    .Y(_12683_));
 sg13g2_buf_2 _19701_ (.A(_12683_),
    .X(_12684_));
 sg13g2_nor2b_1 _19702_ (.A(_12684_),
    .B_N(\cpu.dcache.r_data[5][10] ),
    .Y(_12685_));
 sg13g2_a21oi_1 _19703_ (.A1(net976),
    .A2(_12684_),
    .Y(_12686_),
    .B1(_12685_));
 sg13g2_nand2_1 _19704_ (.Y(_12687_),
    .A(_12058_),
    .B(net40));
 sg13g2_o21ai_1 _19705_ (.B1(_12687_),
    .Y(_00481_),
    .A1(net40),
    .A2(_12686_));
 sg13g2_buf_1 _19706_ (.A(net1092),
    .X(_12688_));
 sg13g2_nor2b_1 _19707_ (.A(_12684_),
    .B_N(\cpu.dcache.r_data[5][11] ),
    .Y(_12689_));
 sg13g2_a21oi_1 _19708_ (.A1(net975),
    .A2(_12684_),
    .Y(_12690_),
    .B1(_12689_));
 sg13g2_nand2_1 _19709_ (.Y(_12691_),
    .A(net408),
    .B(net40));
 sg13g2_o21ai_1 _19710_ (.B1(_12691_),
    .Y(_00482_),
    .A1(net40),
    .A2(_12690_));
 sg13g2_nor2_2 _19711_ (.A(net599),
    .B(_12076_),
    .Y(_12692_));
 sg13g2_mux2_1 _19712_ (.A0(\cpu.dcache.r_data[5][12] ),
    .A1(net1086),
    .S(_12692_),
    .X(_12693_));
 sg13g2_nor2_1 _19713_ (.A(_12680_),
    .B(_12693_),
    .Y(_12694_));
 sg13g2_a21oi_1 _19714_ (.A1(net371),
    .A2(net40),
    .Y(_00483_),
    .B1(_12694_));
 sg13g2_mux2_1 _19715_ (.A0(\cpu.dcache.r_data[5][13] ),
    .A1(net1082),
    .S(_12692_),
    .X(_12695_));
 sg13g2_nor2_1 _19716_ (.A(_12680_),
    .B(_12695_),
    .Y(_12696_));
 sg13g2_a21oi_1 _19717_ (.A1(net370),
    .A2(net40),
    .Y(_00484_),
    .B1(_12696_));
 sg13g2_mux2_1 _19718_ (.A0(\cpu.dcache.r_data[5][14] ),
    .A1(net1085),
    .S(_12692_),
    .X(_12697_));
 sg13g2_nor2_1 _19719_ (.A(_12680_),
    .B(_12697_),
    .Y(_12698_));
 sg13g2_a21oi_1 _19720_ (.A1(net369),
    .A2(_12681_),
    .Y(_00485_),
    .B1(_12698_));
 sg13g2_mux2_1 _19721_ (.A0(\cpu.dcache.r_data[5][15] ),
    .A1(net1084),
    .S(_12692_),
    .X(_12699_));
 sg13g2_nor2_1 _19722_ (.A(_12680_),
    .B(_12699_),
    .Y(_12700_));
 sg13g2_a21oi_1 _19723_ (.A1(net368),
    .A2(_12681_),
    .Y(_00486_),
    .B1(_12700_));
 sg13g2_nor2_1 _19724_ (.A(net599),
    .B(_12251_),
    .Y(_12701_));
 sg13g2_buf_2 _19725_ (.A(_12701_),
    .X(_12702_));
 sg13g2_buf_1 _19726_ (.A(_12702_),
    .X(_12703_));
 sg13g2_nor2_1 _19727_ (.A(net653),
    .B(_12105_),
    .Y(_12704_));
 sg13g2_buf_2 _19728_ (.A(_12704_),
    .X(_12705_));
 sg13g2_nor2b_1 _19729_ (.A(_12705_),
    .B_N(\cpu.dcache.r_data[5][16] ),
    .Y(_12706_));
 sg13g2_a21oi_1 _19730_ (.A1(net977),
    .A2(_12705_),
    .Y(_12707_),
    .B1(_12706_));
 sg13g2_nand2_1 _19731_ (.Y(_12708_),
    .A(net850),
    .B(net39));
 sg13g2_o21ai_1 _19732_ (.B1(_12708_),
    .Y(_00487_),
    .A1(net39),
    .A2(_12707_));
 sg13g2_mux2_1 _19733_ (.A0(\cpu.dcache.r_data[5][17] ),
    .A1(net1082),
    .S(_12705_),
    .X(_12709_));
 sg13g2_nor2_1 _19734_ (.A(_12702_),
    .B(_12709_),
    .Y(_12710_));
 sg13g2_a21oi_1 _19735_ (.A1(net762),
    .A2(net39),
    .Y(_00488_),
    .B1(_12710_));
 sg13g2_nor2b_1 _19736_ (.A(_12705_),
    .B_N(\cpu.dcache.r_data[5][18] ),
    .Y(_12711_));
 sg13g2_a21oi_1 _19737_ (.A1(net976),
    .A2(_12705_),
    .Y(_12712_),
    .B1(_12711_));
 sg13g2_nand2_1 _19738_ (.Y(_12713_),
    .A(net852),
    .B(net39));
 sg13g2_o21ai_1 _19739_ (.B1(_12713_),
    .Y(_00489_),
    .A1(net39),
    .A2(_12712_));
 sg13g2_nor2b_1 _19740_ (.A(_12705_),
    .B_N(\cpu.dcache.r_data[5][19] ),
    .Y(_12714_));
 sg13g2_a21oi_1 _19741_ (.A1(net975),
    .A2(_12705_),
    .Y(_12715_),
    .B1(_12714_));
 sg13g2_buf_1 _19742_ (.A(net1113),
    .X(_12716_));
 sg13g2_nand2_1 _19743_ (.Y(_12717_),
    .A(net974),
    .B(_12702_));
 sg13g2_o21ai_1 _19744_ (.B1(_12717_),
    .Y(_00490_),
    .A1(net39),
    .A2(_12715_));
 sg13g2_mux2_1 _19745_ (.A0(\cpu.dcache.r_data[5][1] ),
    .A1(net1082),
    .S(_12674_),
    .X(_12718_));
 sg13g2_nor2_1 _19746_ (.A(_12670_),
    .B(_12718_),
    .Y(_12719_));
 sg13g2_a21oi_1 _19747_ (.A1(net762),
    .A2(net41),
    .Y(_00491_),
    .B1(_12719_));
 sg13g2_nor2_1 _19748_ (.A(net599),
    .B(_12125_),
    .Y(_12720_));
 sg13g2_buf_2 _19749_ (.A(_12720_),
    .X(_12721_));
 sg13g2_nor2b_1 _19750_ (.A(_12721_),
    .B_N(\cpu.dcache.r_data[5][20] ),
    .Y(_12722_));
 sg13g2_a21oi_1 _19751_ (.A1(net977),
    .A2(_12721_),
    .Y(_12723_),
    .B1(_12722_));
 sg13g2_nand2_1 _19752_ (.Y(_12724_),
    .A(_12193_),
    .B(_12702_));
 sg13g2_o21ai_1 _19753_ (.B1(_12724_),
    .Y(_00492_),
    .A1(net39),
    .A2(_12723_));
 sg13g2_buf_1 _19754_ (.A(net1087),
    .X(_12725_));
 sg13g2_nor2b_1 _19755_ (.A(_12721_),
    .B_N(\cpu.dcache.r_data[5][21] ),
    .Y(_12726_));
 sg13g2_a21oi_1 _19756_ (.A1(net973),
    .A2(_12721_),
    .Y(_12727_),
    .B1(_12726_));
 sg13g2_nand2_1 _19757_ (.Y(_12728_),
    .A(net983),
    .B(_12702_));
 sg13g2_o21ai_1 _19758_ (.B1(_12728_),
    .Y(_00493_),
    .A1(_12703_),
    .A2(_12727_));
 sg13g2_nor2b_1 _19759_ (.A(_12721_),
    .B_N(\cpu.dcache.r_data[5][22] ),
    .Y(_12729_));
 sg13g2_a21oi_1 _19760_ (.A1(net976),
    .A2(_12721_),
    .Y(_12730_),
    .B1(_12729_));
 sg13g2_nand2_1 _19761_ (.Y(_12731_),
    .A(_12333_),
    .B(_12702_));
 sg13g2_o21ai_1 _19762_ (.B1(_12731_),
    .Y(_00494_),
    .A1(_12703_),
    .A2(_12730_));
 sg13g2_nor2b_1 _19763_ (.A(_12721_),
    .B_N(\cpu.dcache.r_data[5][23] ),
    .Y(_02682_));
 sg13g2_a21oi_1 _19764_ (.A1(net975),
    .A2(_12721_),
    .Y(_02683_),
    .B1(_02682_));
 sg13g2_nand2_1 _19765_ (.Y(_02684_),
    .A(_12144_),
    .B(_12702_));
 sg13g2_o21ai_1 _19766_ (.B1(_02684_),
    .Y(_00495_),
    .A1(net39),
    .A2(_02683_));
 sg13g2_nor2_1 _19767_ (.A(net599),
    .B(_12290_),
    .Y(_02685_));
 sg13g2_buf_2 _19768_ (.A(_02685_),
    .X(_02686_));
 sg13g2_buf_1 _19769_ (.A(_02686_),
    .X(_02687_));
 sg13g2_nor2_1 _19770_ (.A(_12667_),
    .B(net654),
    .Y(_02688_));
 sg13g2_buf_1 _19771_ (.A(_02688_),
    .X(_02689_));
 sg13g2_nor2b_1 _19772_ (.A(net526),
    .B_N(\cpu.dcache.r_data[5][24] ),
    .Y(_02690_));
 sg13g2_a21oi_1 _19773_ (.A1(_12672_),
    .A2(net526),
    .Y(_02691_),
    .B1(_02690_));
 sg13g2_nand2_1 _19774_ (.Y(_02692_),
    .A(net409),
    .B(net38));
 sg13g2_o21ai_1 _19775_ (.B1(_02692_),
    .Y(_00496_),
    .A1(net38),
    .A2(_02691_));
 sg13g2_nor2b_1 _19776_ (.A(net526),
    .B_N(\cpu.dcache.r_data[5][25] ),
    .Y(_02693_));
 sg13g2_a21oi_1 _19777_ (.A1(net973),
    .A2(net526),
    .Y(_02694_),
    .B1(_02693_));
 sg13g2_nand2_1 _19778_ (.Y(_02695_),
    .A(net372),
    .B(net38));
 sg13g2_o21ai_1 _19779_ (.B1(_02695_),
    .Y(_00497_),
    .A1(net38),
    .A2(_02694_));
 sg13g2_nor2b_1 _19780_ (.A(net526),
    .B_N(\cpu.dcache.r_data[5][26] ),
    .Y(_02696_));
 sg13g2_a21oi_1 _19781_ (.A1(_12682_),
    .A2(net526),
    .Y(_02697_),
    .B1(_02696_));
 sg13g2_nand2_1 _19782_ (.Y(_02698_),
    .A(_12058_),
    .B(_02686_));
 sg13g2_o21ai_1 _19783_ (.B1(_02698_),
    .Y(_00498_),
    .A1(net38),
    .A2(_02697_));
 sg13g2_nor2b_1 _19784_ (.A(net526),
    .B_N(\cpu.dcache.r_data[5][27] ),
    .Y(_02699_));
 sg13g2_a21oi_1 _19785_ (.A1(_12688_),
    .A2(net526),
    .Y(_02700_),
    .B1(_02699_));
 sg13g2_nand2_1 _19786_ (.Y(_02701_),
    .A(_12067_),
    .B(_02686_));
 sg13g2_o21ai_1 _19787_ (.B1(_02701_),
    .Y(_00499_),
    .A1(net38),
    .A2(_02700_));
 sg13g2_nor2_2 _19788_ (.A(net599),
    .B(_12167_),
    .Y(_02702_));
 sg13g2_mux2_1 _19789_ (.A0(\cpu.dcache.r_data[5][28] ),
    .A1(net1086),
    .S(_02702_),
    .X(_02703_));
 sg13g2_nor2_1 _19790_ (.A(_02686_),
    .B(_02703_),
    .Y(_02704_));
 sg13g2_a21oi_1 _19791_ (.A1(_12072_),
    .A2(net38),
    .Y(_00500_),
    .B1(_02704_));
 sg13g2_mux2_1 _19792_ (.A0(\cpu.dcache.r_data[5][29] ),
    .A1(_12584_),
    .S(_02702_),
    .X(_02705_));
 sg13g2_nor2_1 _19793_ (.A(_02686_),
    .B(_02705_),
    .Y(_02706_));
 sg13g2_a21oi_1 _19794_ (.A1(_12082_),
    .A2(net38),
    .Y(_00501_),
    .B1(_02706_));
 sg13g2_nor2b_1 _19795_ (.A(_12674_),
    .B_N(\cpu.dcache.r_data[5][2] ),
    .Y(_02707_));
 sg13g2_a21oi_1 _19796_ (.A1(net976),
    .A2(_12674_),
    .Y(_02708_),
    .B1(_02707_));
 sg13g2_buf_1 _19797_ (.A(_10132_),
    .X(_02709_));
 sg13g2_nand2_1 _19798_ (.Y(_02710_),
    .A(net849),
    .B(net41));
 sg13g2_o21ai_1 _19799_ (.B1(_02710_),
    .Y(_00502_),
    .A1(_12671_),
    .A2(_02708_));
 sg13g2_mux2_1 _19800_ (.A0(\cpu.dcache.r_data[5][30] ),
    .A1(net1085),
    .S(_02702_),
    .X(_02711_));
 sg13g2_nor2_1 _19801_ (.A(_02686_),
    .B(_02711_),
    .Y(_02712_));
 sg13g2_a21oi_1 _19802_ (.A1(_12089_),
    .A2(_02687_),
    .Y(_00503_),
    .B1(_02712_));
 sg13g2_mux2_1 _19803_ (.A0(\cpu.dcache.r_data[5][31] ),
    .A1(_12246_),
    .S(_02702_),
    .X(_02713_));
 sg13g2_nor2_1 _19804_ (.A(_02686_),
    .B(_02713_),
    .Y(_02714_));
 sg13g2_a21oi_1 _19805_ (.A1(_12095_),
    .A2(_02687_),
    .Y(_00504_),
    .B1(_02714_));
 sg13g2_nor2b_1 _19806_ (.A(_12674_),
    .B_N(\cpu.dcache.r_data[5][3] ),
    .Y(_02715_));
 sg13g2_a21oi_1 _19807_ (.A1(net975),
    .A2(_12674_),
    .Y(_02716_),
    .B1(_02715_));
 sg13g2_nand2_1 _19808_ (.Y(_02717_),
    .A(net974),
    .B(_12670_));
 sg13g2_o21ai_1 _19809_ (.B1(_02717_),
    .Y(_00505_),
    .A1(_12671_),
    .A2(_02716_));
 sg13g2_nor2_1 _19810_ (.A(net653),
    .B(_12188_),
    .Y(_02718_));
 sg13g2_buf_2 _19811_ (.A(_02718_),
    .X(_02719_));
 sg13g2_nor2b_1 _19812_ (.A(_02719_),
    .B_N(\cpu.dcache.r_data[5][4] ),
    .Y(_02720_));
 sg13g2_a21oi_1 _19813_ (.A1(net977),
    .A2(_02719_),
    .Y(_02721_),
    .B1(_02720_));
 sg13g2_nand2_1 _19814_ (.Y(_02722_),
    .A(net987),
    .B(_12670_));
 sg13g2_o21ai_1 _19815_ (.B1(_02722_),
    .Y(_00506_),
    .A1(net41),
    .A2(_02721_));
 sg13g2_nor2b_1 _19816_ (.A(_02719_),
    .B_N(\cpu.dcache.r_data[5][5] ),
    .Y(_02723_));
 sg13g2_a21oi_1 _19817_ (.A1(net973),
    .A2(_02719_),
    .Y(_02724_),
    .B1(_02723_));
 sg13g2_nand2_1 _19818_ (.Y(_02725_),
    .A(net983),
    .B(_12670_));
 sg13g2_o21ai_1 _19819_ (.B1(_02725_),
    .Y(_00507_),
    .A1(net41),
    .A2(_02724_));
 sg13g2_nor2b_1 _19820_ (.A(_02719_),
    .B_N(\cpu.dcache.r_data[5][6] ),
    .Y(_02726_));
 sg13g2_a21oi_1 _19821_ (.A1(net976),
    .A2(_02719_),
    .Y(_02727_),
    .B1(_02726_));
 sg13g2_nand2_1 _19822_ (.Y(_02728_),
    .A(net982),
    .B(_12670_));
 sg13g2_o21ai_1 _19823_ (.B1(_02728_),
    .Y(_00508_),
    .A1(net41),
    .A2(_02727_));
 sg13g2_nor2b_1 _19824_ (.A(_02719_),
    .B_N(\cpu.dcache.r_data[5][7] ),
    .Y(_02729_));
 sg13g2_a21oi_1 _19825_ (.A1(net975),
    .A2(_02719_),
    .Y(_02730_),
    .B1(_02729_));
 sg13g2_nand2_1 _19826_ (.Y(_02731_),
    .A(net988),
    .B(_12670_));
 sg13g2_o21ai_1 _19827_ (.B1(_02731_),
    .Y(_00509_),
    .A1(net41),
    .A2(_02730_));
 sg13g2_nor2b_1 _19828_ (.A(_12684_),
    .B_N(\cpu.dcache.r_data[5][8] ),
    .Y(_02732_));
 sg13g2_a21oi_1 _19829_ (.A1(_12672_),
    .A2(_12684_),
    .Y(_02733_),
    .B1(_02732_));
 sg13g2_nand2_1 _19830_ (.Y(_02734_),
    .A(_12150_),
    .B(_12680_));
 sg13g2_o21ai_1 _19831_ (.B1(_02734_),
    .Y(_00510_),
    .A1(net40),
    .A2(_02733_));
 sg13g2_nor2b_1 _19832_ (.A(_12684_),
    .B_N(\cpu.dcache.r_data[5][9] ),
    .Y(_02735_));
 sg13g2_a21oi_1 _19833_ (.A1(net973),
    .A2(_12684_),
    .Y(_02736_),
    .B1(_02735_));
 sg13g2_nand2_1 _19834_ (.Y(_02737_),
    .A(_12160_),
    .B(_12680_));
 sg13g2_o21ai_1 _19835_ (.B1(_02737_),
    .Y(_00511_),
    .A1(net40),
    .A2(_02736_));
 sg13g2_nand2_1 _19836_ (.Y(_02738_),
    .A(net784),
    .B(_09416_));
 sg13g2_buf_2 _19837_ (.A(_02738_),
    .X(_02739_));
 sg13g2_buf_1 _19838_ (.A(_02739_),
    .X(_02740_));
 sg13g2_nor2_1 _19839_ (.A(net525),
    .B(_12215_),
    .Y(_02741_));
 sg13g2_buf_2 _19840_ (.A(_02741_),
    .X(_02742_));
 sg13g2_buf_1 _19841_ (.A(_02742_),
    .X(_02743_));
 sg13g2_nor2_1 _19842_ (.A(_02739_),
    .B(_12032_),
    .Y(_02744_));
 sg13g2_buf_2 _19843_ (.A(_02744_),
    .X(_02745_));
 sg13g2_nor2b_1 _19844_ (.A(_02745_),
    .B_N(\cpu.dcache.r_data[6][0] ),
    .Y(_02746_));
 sg13g2_a21oi_1 _19845_ (.A1(net977),
    .A2(_02745_),
    .Y(_02747_),
    .B1(_02746_));
 sg13g2_nand2_1 _19846_ (.Y(_02748_),
    .A(net850),
    .B(net37));
 sg13g2_o21ai_1 _19847_ (.B1(_02748_),
    .Y(_00512_),
    .A1(net37),
    .A2(_02747_));
 sg13g2_nor2_1 _19848_ (.A(net525),
    .B(_12225_),
    .Y(_02749_));
 sg13g2_buf_2 _19849_ (.A(_02749_),
    .X(_02750_));
 sg13g2_buf_1 _19850_ (.A(_02750_),
    .X(_02751_));
 sg13g2_nor2_1 _19851_ (.A(net525),
    .B(_12048_),
    .Y(_02752_));
 sg13g2_buf_2 _19852_ (.A(_02752_),
    .X(_02753_));
 sg13g2_nor2b_1 _19853_ (.A(_02753_),
    .B_N(\cpu.dcache.r_data[6][10] ),
    .Y(_02754_));
 sg13g2_a21oi_1 _19854_ (.A1(net976),
    .A2(_02753_),
    .Y(_02755_),
    .B1(_02754_));
 sg13g2_nand2_1 _19855_ (.Y(_02756_),
    .A(_12058_),
    .B(net36));
 sg13g2_o21ai_1 _19856_ (.B1(_02756_),
    .Y(_00513_),
    .A1(net36),
    .A2(_02755_));
 sg13g2_nor2b_1 _19857_ (.A(_02753_),
    .B_N(\cpu.dcache.r_data[6][11] ),
    .Y(_02757_));
 sg13g2_a21oi_1 _19858_ (.A1(net975),
    .A2(_02753_),
    .Y(_02758_),
    .B1(_02757_));
 sg13g2_nand2_1 _19859_ (.Y(_02759_),
    .A(_12067_),
    .B(net36));
 sg13g2_o21ai_1 _19860_ (.B1(_02759_),
    .Y(_00514_),
    .A1(net36),
    .A2(_02758_));
 sg13g2_nor2_2 _19861_ (.A(net525),
    .B(_12076_),
    .Y(_02760_));
 sg13g2_mux2_1 _19862_ (.A0(\cpu.dcache.r_data[6][12] ),
    .A1(net1095),
    .S(_02760_),
    .X(_02761_));
 sg13g2_nor2_1 _19863_ (.A(_02750_),
    .B(_02761_),
    .Y(_02762_));
 sg13g2_a21oi_1 _19864_ (.A1(_12072_),
    .A2(_02751_),
    .Y(_00515_),
    .B1(_02762_));
 sg13g2_mux2_1 _19865_ (.A0(\cpu.dcache.r_data[6][13] ),
    .A1(_12584_),
    .S(_02760_),
    .X(_02763_));
 sg13g2_nor2_1 _19866_ (.A(_02750_),
    .B(_02763_),
    .Y(_02764_));
 sg13g2_a21oi_1 _19867_ (.A1(_12082_),
    .A2(net36),
    .Y(_00516_),
    .B1(_02764_));
 sg13g2_mux2_1 _19868_ (.A0(\cpu.dcache.r_data[6][14] ),
    .A1(net1093),
    .S(_02760_),
    .X(_02765_));
 sg13g2_nor2_1 _19869_ (.A(_02750_),
    .B(_02765_),
    .Y(_02766_));
 sg13g2_a21oi_1 _19870_ (.A1(_12089_),
    .A2(_02751_),
    .Y(_00517_),
    .B1(_02766_));
 sg13g2_mux2_1 _19871_ (.A0(\cpu.dcache.r_data[6][15] ),
    .A1(net1092),
    .S(_02760_),
    .X(_02767_));
 sg13g2_nor2_1 _19872_ (.A(_02750_),
    .B(_02767_),
    .Y(_02768_));
 sg13g2_a21oi_1 _19873_ (.A1(_12095_),
    .A2(net36),
    .Y(_00518_),
    .B1(_02768_));
 sg13g2_nor2_1 _19874_ (.A(net525),
    .B(_12251_),
    .Y(_02769_));
 sg13g2_buf_2 _19875_ (.A(_02769_),
    .X(_02770_));
 sg13g2_buf_1 _19876_ (.A(_02770_),
    .X(_02771_));
 sg13g2_nor2_1 _19877_ (.A(_02739_),
    .B(_12105_),
    .Y(_02772_));
 sg13g2_buf_2 _19878_ (.A(_02772_),
    .X(_02773_));
 sg13g2_nor2b_1 _19879_ (.A(_02773_),
    .B_N(\cpu.dcache.r_data[6][16] ),
    .Y(_02774_));
 sg13g2_a21oi_1 _19880_ (.A1(net977),
    .A2(_02773_),
    .Y(_02775_),
    .B1(_02774_));
 sg13g2_nand2_1 _19881_ (.Y(_02776_),
    .A(_12677_),
    .B(net35));
 sg13g2_o21ai_1 _19882_ (.B1(_02776_),
    .Y(_00519_),
    .A1(_02771_),
    .A2(_02775_));
 sg13g2_mux2_1 _19883_ (.A0(\cpu.dcache.r_data[6][17] ),
    .A1(net1082),
    .S(_02773_),
    .X(_02777_));
 sg13g2_nor2_1 _19884_ (.A(_02770_),
    .B(_02777_),
    .Y(_02778_));
 sg13g2_a21oi_1 _19885_ (.A1(_10116_),
    .A2(_02771_),
    .Y(_00520_),
    .B1(_02778_));
 sg13g2_nor2b_1 _19886_ (.A(_02773_),
    .B_N(\cpu.dcache.r_data[6][18] ),
    .Y(_02779_));
 sg13g2_a21oi_1 _19887_ (.A1(net976),
    .A2(_02773_),
    .Y(_02780_),
    .B1(_02779_));
 sg13g2_nand2_1 _19888_ (.Y(_02781_),
    .A(net849),
    .B(net35));
 sg13g2_o21ai_1 _19889_ (.B1(_02781_),
    .Y(_00521_),
    .A1(net35),
    .A2(_02780_));
 sg13g2_nor2b_1 _19890_ (.A(_02773_),
    .B_N(\cpu.dcache.r_data[6][19] ),
    .Y(_02782_));
 sg13g2_a21oi_1 _19891_ (.A1(net975),
    .A2(_02773_),
    .Y(_02783_),
    .B1(_02782_));
 sg13g2_nand2_1 _19892_ (.Y(_02784_),
    .A(net974),
    .B(_02770_));
 sg13g2_o21ai_1 _19893_ (.B1(_02784_),
    .Y(_00522_),
    .A1(net35),
    .A2(_02783_));
 sg13g2_mux2_1 _19894_ (.A0(\cpu.dcache.r_data[6][1] ),
    .A1(net1087),
    .S(_02745_),
    .X(_02785_));
 sg13g2_nor2_1 _19895_ (.A(_02742_),
    .B(_02785_),
    .Y(_02786_));
 sg13g2_a21oi_1 _19896_ (.A1(net762),
    .A2(_02743_),
    .Y(_00523_),
    .B1(_02786_));
 sg13g2_nor2_1 _19897_ (.A(net525),
    .B(_12125_),
    .Y(_02787_));
 sg13g2_buf_2 _19898_ (.A(_02787_),
    .X(_02788_));
 sg13g2_nor2b_1 _19899_ (.A(_02788_),
    .B_N(\cpu.dcache.r_data[6][20] ),
    .Y(_02789_));
 sg13g2_a21oi_1 _19900_ (.A1(net977),
    .A2(_02788_),
    .Y(_02790_),
    .B1(_02789_));
 sg13g2_nand2_1 _19901_ (.Y(_02791_),
    .A(_12193_),
    .B(_02770_));
 sg13g2_o21ai_1 _19902_ (.B1(_02791_),
    .Y(_00524_),
    .A1(net35),
    .A2(_02790_));
 sg13g2_nor2b_1 _19903_ (.A(_02788_),
    .B_N(\cpu.dcache.r_data[6][21] ),
    .Y(_02792_));
 sg13g2_a21oi_1 _19904_ (.A1(net973),
    .A2(_02788_),
    .Y(_02793_),
    .B1(_02792_));
 sg13g2_nand2_1 _19905_ (.Y(_02794_),
    .A(_12281_),
    .B(_02770_));
 sg13g2_o21ai_1 _19906_ (.B1(_02794_),
    .Y(_00525_),
    .A1(net35),
    .A2(_02793_));
 sg13g2_nor2b_1 _19907_ (.A(_02788_),
    .B_N(\cpu.dcache.r_data[6][22] ),
    .Y(_02795_));
 sg13g2_a21oi_1 _19908_ (.A1(net976),
    .A2(_02788_),
    .Y(_02796_),
    .B1(_02795_));
 sg13g2_nand2_1 _19909_ (.Y(_02797_),
    .A(_12333_),
    .B(_02770_));
 sg13g2_o21ai_1 _19910_ (.B1(_02797_),
    .Y(_00526_),
    .A1(net35),
    .A2(_02796_));
 sg13g2_nor2b_1 _19911_ (.A(_02788_),
    .B_N(\cpu.dcache.r_data[6][23] ),
    .Y(_02798_));
 sg13g2_a21oi_1 _19912_ (.A1(net975),
    .A2(_02788_),
    .Y(_02799_),
    .B1(_02798_));
 sg13g2_nand2_1 _19913_ (.Y(_02800_),
    .A(_10104_),
    .B(_02770_));
 sg13g2_o21ai_1 _19914_ (.B1(_02800_),
    .Y(_00527_),
    .A1(net35),
    .A2(_02799_));
 sg13g2_nor2_1 _19915_ (.A(_02740_),
    .B(_12290_),
    .Y(_02801_));
 sg13g2_buf_2 _19916_ (.A(_02801_),
    .X(_02802_));
 sg13g2_buf_1 _19917_ (.A(_02802_),
    .X(_02803_));
 sg13g2_nor2_1 _19918_ (.A(_02739_),
    .B(net654),
    .Y(_02804_));
 sg13g2_buf_1 _19919_ (.A(_02804_),
    .X(_02805_));
 sg13g2_nor2b_1 _19920_ (.A(net467),
    .B_N(\cpu.dcache.r_data[6][24] ),
    .Y(_02806_));
 sg13g2_a21oi_1 _19921_ (.A1(net977),
    .A2(net467),
    .Y(_02807_),
    .B1(_02806_));
 sg13g2_nand2_1 _19922_ (.Y(_02808_),
    .A(_12150_),
    .B(net34));
 sg13g2_o21ai_1 _19923_ (.B1(_02808_),
    .Y(_00528_),
    .A1(net34),
    .A2(_02807_));
 sg13g2_nor2b_1 _19924_ (.A(net467),
    .B_N(\cpu.dcache.r_data[6][25] ),
    .Y(_02809_));
 sg13g2_a21oi_1 _19925_ (.A1(_12725_),
    .A2(net467),
    .Y(_02810_),
    .B1(_02809_));
 sg13g2_nand2_1 _19926_ (.Y(_02811_),
    .A(_12160_),
    .B(net34));
 sg13g2_o21ai_1 _19927_ (.B1(_02811_),
    .Y(_00529_),
    .A1(net34),
    .A2(_02810_));
 sg13g2_nor2b_1 _19928_ (.A(net467),
    .B_N(\cpu.dcache.r_data[6][26] ),
    .Y(_02812_));
 sg13g2_a21oi_1 _19929_ (.A1(_12682_),
    .A2(net467),
    .Y(_02813_),
    .B1(_02812_));
 sg13g2_nand2_1 _19930_ (.Y(_02814_),
    .A(_12058_),
    .B(_02802_));
 sg13g2_o21ai_1 _19931_ (.B1(_02814_),
    .Y(_00530_),
    .A1(_02803_),
    .A2(_02813_));
 sg13g2_nor2b_1 _19932_ (.A(net467),
    .B_N(\cpu.dcache.r_data[6][27] ),
    .Y(_02815_));
 sg13g2_a21oi_1 _19933_ (.A1(_12688_),
    .A2(net467),
    .Y(_02816_),
    .B1(_02815_));
 sg13g2_nand2_1 _19934_ (.Y(_02817_),
    .A(_12067_),
    .B(_02802_));
 sg13g2_o21ai_1 _19935_ (.B1(_02817_),
    .Y(_00531_),
    .A1(net34),
    .A2(_02816_));
 sg13g2_nor2_2 _19936_ (.A(net525),
    .B(_12167_),
    .Y(_02818_));
 sg13g2_mux2_1 _19937_ (.A0(\cpu.dcache.r_data[6][28] ),
    .A1(net1095),
    .S(_02818_),
    .X(_02819_));
 sg13g2_nor2_1 _19938_ (.A(_02802_),
    .B(_02819_),
    .Y(_02820_));
 sg13g2_a21oi_1 _19939_ (.A1(_12072_),
    .A2(net34),
    .Y(_00532_),
    .B1(_02820_));
 sg13g2_mux2_1 _19940_ (.A0(\cpu.dcache.r_data[6][29] ),
    .A1(net1087),
    .S(_02818_),
    .X(_02821_));
 sg13g2_nor2_1 _19941_ (.A(_02802_),
    .B(_02821_),
    .Y(_02822_));
 sg13g2_a21oi_1 _19942_ (.A1(_12082_),
    .A2(net34),
    .Y(_00533_),
    .B1(_02822_));
 sg13g2_buf_2 _19943_ (.A(net1093),
    .X(_02823_));
 sg13g2_nor2b_1 _19944_ (.A(_02745_),
    .B_N(\cpu.dcache.r_data[6][2] ),
    .Y(_02824_));
 sg13g2_a21oi_1 _19945_ (.A1(net972),
    .A2(_02745_),
    .Y(_02825_),
    .B1(_02824_));
 sg13g2_nand2_1 _19946_ (.Y(_02826_),
    .A(net849),
    .B(net37));
 sg13g2_o21ai_1 _19947_ (.B1(_02826_),
    .Y(_00534_),
    .A1(net37),
    .A2(_02825_));
 sg13g2_mux2_1 _19948_ (.A0(\cpu.dcache.r_data[6][30] ),
    .A1(net1093),
    .S(_02818_),
    .X(_02827_));
 sg13g2_nor2_1 _19949_ (.A(_02802_),
    .B(_02827_),
    .Y(_02828_));
 sg13g2_a21oi_1 _19950_ (.A1(_12089_),
    .A2(_02803_),
    .Y(_00535_),
    .B1(_02828_));
 sg13g2_mux2_1 _19951_ (.A0(\cpu.dcache.r_data[6][31] ),
    .A1(net1092),
    .S(_02818_),
    .X(_02829_));
 sg13g2_nor2_1 _19952_ (.A(_02802_),
    .B(_02829_),
    .Y(_02830_));
 sg13g2_a21oi_1 _19953_ (.A1(_12095_),
    .A2(net34),
    .Y(_00536_),
    .B1(_02830_));
 sg13g2_buf_2 _19954_ (.A(net1092),
    .X(_02831_));
 sg13g2_nor2b_1 _19955_ (.A(_02745_),
    .B_N(\cpu.dcache.r_data[6][3] ),
    .Y(_02832_));
 sg13g2_a21oi_1 _19956_ (.A1(net971),
    .A2(_02745_),
    .Y(_02833_),
    .B1(_02832_));
 sg13g2_nand2_1 _19957_ (.Y(_02834_),
    .A(net974),
    .B(_02742_));
 sg13g2_o21ai_1 _19958_ (.B1(_02834_),
    .Y(_00537_),
    .A1(_02743_),
    .A2(_02833_));
 sg13g2_buf_2 _19959_ (.A(net1095),
    .X(_02835_));
 sg13g2_nor2_1 _19960_ (.A(_02739_),
    .B(_12188_),
    .Y(_02836_));
 sg13g2_buf_2 _19961_ (.A(_02836_),
    .X(_02837_));
 sg13g2_nor2b_1 _19962_ (.A(_02837_),
    .B_N(\cpu.dcache.r_data[6][4] ),
    .Y(_02838_));
 sg13g2_a21oi_1 _19963_ (.A1(net970),
    .A2(_02837_),
    .Y(_02839_),
    .B1(_02838_));
 sg13g2_nand2_1 _19964_ (.Y(_02840_),
    .A(net1024),
    .B(_02742_));
 sg13g2_o21ai_1 _19965_ (.B1(_02840_),
    .Y(_00538_),
    .A1(net37),
    .A2(_02839_));
 sg13g2_nor2b_1 _19966_ (.A(_02837_),
    .B_N(\cpu.dcache.r_data[6][5] ),
    .Y(_02841_));
 sg13g2_a21oi_1 _19967_ (.A1(net973),
    .A2(_02837_),
    .Y(_02842_),
    .B1(_02841_));
 sg13g2_nand2_1 _19968_ (.Y(_02843_),
    .A(net983),
    .B(_02742_));
 sg13g2_o21ai_1 _19969_ (.B1(_02843_),
    .Y(_00539_),
    .A1(net37),
    .A2(_02842_));
 sg13g2_nor2b_1 _19970_ (.A(_02837_),
    .B_N(\cpu.dcache.r_data[6][6] ),
    .Y(_02844_));
 sg13g2_a21oi_1 _19971_ (.A1(net972),
    .A2(_02837_),
    .Y(_02845_),
    .B1(_02844_));
 sg13g2_nand2_1 _19972_ (.Y(_02846_),
    .A(net982),
    .B(_02742_));
 sg13g2_o21ai_1 _19973_ (.B1(_02846_),
    .Y(_00540_),
    .A1(net37),
    .A2(_02845_));
 sg13g2_nor2b_1 _19974_ (.A(_02837_),
    .B_N(\cpu.dcache.r_data[6][7] ),
    .Y(_02847_));
 sg13g2_a21oi_1 _19975_ (.A1(net971),
    .A2(_02837_),
    .Y(_02848_),
    .B1(_02847_));
 sg13g2_nand2_1 _19976_ (.Y(_02849_),
    .A(net1021),
    .B(_02742_));
 sg13g2_o21ai_1 _19977_ (.B1(_02849_),
    .Y(_00541_),
    .A1(net37),
    .A2(_02848_));
 sg13g2_nor2b_1 _19978_ (.A(_02753_),
    .B_N(\cpu.dcache.r_data[6][8] ),
    .Y(_02850_));
 sg13g2_a21oi_1 _19979_ (.A1(net970),
    .A2(_02753_),
    .Y(_02851_),
    .B1(_02850_));
 sg13g2_nand2_1 _19980_ (.Y(_02852_),
    .A(_12150_),
    .B(_02750_));
 sg13g2_o21ai_1 _19981_ (.B1(_02852_),
    .Y(_00542_),
    .A1(net36),
    .A2(_02851_));
 sg13g2_nor2b_1 _19982_ (.A(_02753_),
    .B_N(\cpu.dcache.r_data[6][9] ),
    .Y(_02853_));
 sg13g2_a21oi_1 _19983_ (.A1(net973),
    .A2(_02753_),
    .Y(_02854_),
    .B1(_02853_));
 sg13g2_nand2_1 _19984_ (.Y(_02855_),
    .A(_12160_),
    .B(_02750_));
 sg13g2_o21ai_1 _19985_ (.B1(_02855_),
    .Y(_00543_),
    .A1(net36),
    .A2(_02854_));
 sg13g2_buf_1 _19986_ (.A(net539),
    .X(_02856_));
 sg13g2_nor2_1 _19987_ (.A(net466),
    .B(_12215_),
    .Y(_02857_));
 sg13g2_buf_1 _19988_ (.A(_02857_),
    .X(_02858_));
 sg13g2_nor2_1 _19989_ (.A(net539),
    .B(_12032_),
    .Y(_02859_));
 sg13g2_buf_2 _19990_ (.A(_02859_),
    .X(_02860_));
 sg13g2_nor2b_1 _19991_ (.A(_02860_),
    .B_N(\cpu.dcache.r_data[7][0] ),
    .Y(_02861_));
 sg13g2_a21oi_1 _19992_ (.A1(net970),
    .A2(_02860_),
    .Y(_02862_),
    .B1(_02861_));
 sg13g2_nand2_1 _19993_ (.Y(_02863_),
    .A(net850),
    .B(net63));
 sg13g2_o21ai_1 _19994_ (.B1(_02863_),
    .Y(_00544_),
    .A1(net63),
    .A2(_02862_));
 sg13g2_nor2_1 _19995_ (.A(net466),
    .B(_12225_),
    .Y(_02864_));
 sg13g2_buf_2 _19996_ (.A(_02864_),
    .X(_02865_));
 sg13g2_buf_1 _19997_ (.A(_02865_),
    .X(_02866_));
 sg13g2_nor2_1 _19998_ (.A(net539),
    .B(_12048_),
    .Y(_02867_));
 sg13g2_buf_2 _19999_ (.A(_02867_),
    .X(_02868_));
 sg13g2_nor2b_1 _20000_ (.A(_02868_),
    .B_N(\cpu.dcache.r_data[7][10] ),
    .Y(_02869_));
 sg13g2_a21oi_1 _20001_ (.A1(net972),
    .A2(_02868_),
    .Y(_02870_),
    .B1(_02869_));
 sg13g2_nand2_1 _20002_ (.Y(_02871_),
    .A(_12058_),
    .B(net33));
 sg13g2_o21ai_1 _20003_ (.B1(_02871_),
    .Y(_00545_),
    .A1(net33),
    .A2(_02870_));
 sg13g2_nor2b_1 _20004_ (.A(_02868_),
    .B_N(\cpu.dcache.r_data[7][11] ),
    .Y(_02872_));
 sg13g2_a21oi_1 _20005_ (.A1(net971),
    .A2(_02868_),
    .Y(_02873_),
    .B1(_02872_));
 sg13g2_nand2_1 _20006_ (.Y(_02874_),
    .A(_12067_),
    .B(net33));
 sg13g2_o21ai_1 _20007_ (.B1(_02874_),
    .Y(_00546_),
    .A1(net33),
    .A2(_02873_));
 sg13g2_nor2_2 _20008_ (.A(net466),
    .B(_12076_),
    .Y(_02875_));
 sg13g2_mux2_1 _20009_ (.A0(\cpu.dcache.r_data[7][12] ),
    .A1(net1095),
    .S(_02875_),
    .X(_02876_));
 sg13g2_nor2_1 _20010_ (.A(_02865_),
    .B(_02876_),
    .Y(_02877_));
 sg13g2_a21oi_1 _20011_ (.A1(_12072_),
    .A2(net33),
    .Y(_00547_),
    .B1(_02877_));
 sg13g2_mux2_1 _20012_ (.A0(\cpu.dcache.r_data[7][13] ),
    .A1(net1087),
    .S(_02875_),
    .X(_02878_));
 sg13g2_nor2_1 _20013_ (.A(_02865_),
    .B(_02878_),
    .Y(_02879_));
 sg13g2_a21oi_1 _20014_ (.A1(_12082_),
    .A2(net33),
    .Y(_00548_),
    .B1(_02879_));
 sg13g2_mux2_1 _20015_ (.A0(\cpu.dcache.r_data[7][14] ),
    .A1(net1093),
    .S(_02875_),
    .X(_02880_));
 sg13g2_nor2_1 _20016_ (.A(_02865_),
    .B(_02880_),
    .Y(_02881_));
 sg13g2_a21oi_1 _20017_ (.A1(_12089_),
    .A2(_02866_),
    .Y(_00549_),
    .B1(_02881_));
 sg13g2_mux2_1 _20018_ (.A0(\cpu.dcache.r_data[7][15] ),
    .A1(net1092),
    .S(_02875_),
    .X(_02882_));
 sg13g2_nor2_1 _20019_ (.A(_02865_),
    .B(_02882_),
    .Y(_02883_));
 sg13g2_a21oi_1 _20020_ (.A1(_12095_),
    .A2(_02866_),
    .Y(_00550_),
    .B1(_02883_));
 sg13g2_nor2_1 _20021_ (.A(net466),
    .B(_12251_),
    .Y(_02884_));
 sg13g2_buf_1 _20022_ (.A(_02884_),
    .X(_02885_));
 sg13g2_nor2_1 _20023_ (.A(net539),
    .B(_12105_),
    .Y(_02886_));
 sg13g2_buf_2 _20024_ (.A(_02886_),
    .X(_02887_));
 sg13g2_nor2b_1 _20025_ (.A(_02887_),
    .B_N(\cpu.dcache.r_data[7][16] ),
    .Y(_02888_));
 sg13g2_a21oi_1 _20026_ (.A1(net970),
    .A2(_02887_),
    .Y(_02889_),
    .B1(_02888_));
 sg13g2_nand2_1 _20027_ (.Y(_02890_),
    .A(_12677_),
    .B(net62));
 sg13g2_o21ai_1 _20028_ (.B1(_02890_),
    .Y(_00551_),
    .A1(net62),
    .A2(_02889_));
 sg13g2_mux2_1 _20029_ (.A0(\cpu.dcache.r_data[7][17] ),
    .A1(net1087),
    .S(_02887_),
    .X(_02891_));
 sg13g2_nor2_1 _20030_ (.A(_02884_),
    .B(_02891_),
    .Y(_02892_));
 sg13g2_a21oi_1 _20031_ (.A1(net762),
    .A2(_02885_),
    .Y(_00552_),
    .B1(_02892_));
 sg13g2_nor2b_1 _20032_ (.A(_02887_),
    .B_N(\cpu.dcache.r_data[7][18] ),
    .Y(_02893_));
 sg13g2_a21oi_1 _20033_ (.A1(net972),
    .A2(_02887_),
    .Y(_02894_),
    .B1(_02893_));
 sg13g2_nand2_1 _20034_ (.Y(_02895_),
    .A(net849),
    .B(net62));
 sg13g2_o21ai_1 _20035_ (.B1(_02895_),
    .Y(_00553_),
    .A1(_02885_),
    .A2(_02894_));
 sg13g2_nor2b_1 _20036_ (.A(_02887_),
    .B_N(\cpu.dcache.r_data[7][19] ),
    .Y(_02896_));
 sg13g2_a21oi_1 _20037_ (.A1(net971),
    .A2(_02887_),
    .Y(_02897_),
    .B1(_02896_));
 sg13g2_nand2_1 _20038_ (.Y(_02898_),
    .A(_12716_),
    .B(_02884_));
 sg13g2_o21ai_1 _20039_ (.B1(_02898_),
    .Y(_00554_),
    .A1(net62),
    .A2(_02897_));
 sg13g2_mux2_1 _20040_ (.A0(\cpu.dcache.r_data[7][1] ),
    .A1(net1087),
    .S(_02860_),
    .X(_02899_));
 sg13g2_nor2_1 _20041_ (.A(_02857_),
    .B(_02899_),
    .Y(_02900_));
 sg13g2_a21oi_1 _20042_ (.A1(_10116_),
    .A2(net63),
    .Y(_00555_),
    .B1(_02900_));
 sg13g2_or2_1 _20043_ (.X(_02901_),
    .B(_12125_),
    .A(net466));
 sg13g2_buf_1 _20044_ (.A(_02901_),
    .X(_02902_));
 sg13g2_mux2_1 _20045_ (.A0(net1091),
    .A1(\cpu.dcache.r_data[7][20] ),
    .S(_02902_),
    .X(_02903_));
 sg13g2_mux2_1 _20046_ (.A0(_02903_),
    .A1(net992),
    .S(net62),
    .X(_00556_));
 sg13g2_mux2_1 _20047_ (.A0(net1090),
    .A1(\cpu.dcache.r_data[7][21] ),
    .S(_02902_),
    .X(_02904_));
 sg13g2_mux2_1 _20048_ (.A0(_02904_),
    .A1(net990),
    .S(net62),
    .X(_00557_));
 sg13g2_mux2_1 _20049_ (.A0(net1089),
    .A1(\cpu.dcache.r_data[7][22] ),
    .S(_02902_),
    .X(_02905_));
 sg13g2_mux2_1 _20050_ (.A0(_02905_),
    .A1(_12140_),
    .S(net62),
    .X(_00558_));
 sg13g2_mux2_1 _20051_ (.A0(net1088),
    .A1(\cpu.dcache.r_data[7][23] ),
    .S(_02902_),
    .X(_02906_));
 sg13g2_mux2_1 _20052_ (.A0(_02906_),
    .A1(_12516_),
    .S(net62),
    .X(_00559_));
 sg13g2_nor2_1 _20053_ (.A(_02856_),
    .B(_12290_),
    .Y(_02907_));
 sg13g2_buf_2 _20054_ (.A(_02907_),
    .X(_02908_));
 sg13g2_buf_1 _20055_ (.A(_02908_),
    .X(_02909_));
 sg13g2_nor2_1 _20056_ (.A(_10056_),
    .B(net654),
    .Y(_02910_));
 sg13g2_buf_1 _20057_ (.A(_02910_),
    .X(_02911_));
 sg13g2_nor2b_1 _20058_ (.A(net406),
    .B_N(\cpu.dcache.r_data[7][24] ),
    .Y(_02912_));
 sg13g2_a21oi_1 _20059_ (.A1(net970),
    .A2(net406),
    .Y(_02913_),
    .B1(_02912_));
 sg13g2_nand2_1 _20060_ (.Y(_02914_),
    .A(_12150_),
    .B(net32));
 sg13g2_o21ai_1 _20061_ (.B1(_02914_),
    .Y(_00560_),
    .A1(_02909_),
    .A2(_02913_));
 sg13g2_nor2b_1 _20062_ (.A(net406),
    .B_N(\cpu.dcache.r_data[7][25] ),
    .Y(_02915_));
 sg13g2_a21oi_1 _20063_ (.A1(_12725_),
    .A2(net406),
    .Y(_02916_),
    .B1(_02915_));
 sg13g2_nand2_1 _20064_ (.Y(_02917_),
    .A(_12160_),
    .B(net32));
 sg13g2_o21ai_1 _20065_ (.B1(_02917_),
    .Y(_00561_),
    .A1(net32),
    .A2(_02916_));
 sg13g2_nor2b_1 _20066_ (.A(net406),
    .B_N(\cpu.dcache.r_data[7][26] ),
    .Y(_02918_));
 sg13g2_a21oi_1 _20067_ (.A1(net972),
    .A2(net406),
    .Y(_02919_),
    .B1(_02918_));
 sg13g2_nand2_1 _20068_ (.Y(_02920_),
    .A(_12058_),
    .B(_02908_));
 sg13g2_o21ai_1 _20069_ (.B1(_02920_),
    .Y(_00562_),
    .A1(net32),
    .A2(_02919_));
 sg13g2_nor2b_1 _20070_ (.A(net406),
    .B_N(\cpu.dcache.r_data[7][27] ),
    .Y(_02921_));
 sg13g2_a21oi_1 _20071_ (.A1(net971),
    .A2(net406),
    .Y(_02922_),
    .B1(_02921_));
 sg13g2_nand2_1 _20072_ (.Y(_02923_),
    .A(_12067_),
    .B(_02908_));
 sg13g2_o21ai_1 _20073_ (.B1(_02923_),
    .Y(_00563_),
    .A1(_02909_),
    .A2(_02922_));
 sg13g2_nor2_2 _20074_ (.A(net466),
    .B(_12167_),
    .Y(_02924_));
 sg13g2_mux2_1 _20075_ (.A0(\cpu.dcache.r_data[7][28] ),
    .A1(net1095),
    .S(_02924_),
    .X(_02925_));
 sg13g2_nor2_1 _20076_ (.A(_02908_),
    .B(_02925_),
    .Y(_02926_));
 sg13g2_a21oi_1 _20077_ (.A1(_12072_),
    .A2(net32),
    .Y(_00564_),
    .B1(_02926_));
 sg13g2_mux2_1 _20078_ (.A0(\cpu.dcache.r_data[7][29] ),
    .A1(_12132_),
    .S(_02924_),
    .X(_02927_));
 sg13g2_nor2_1 _20079_ (.A(_02908_),
    .B(_02927_),
    .Y(_02928_));
 sg13g2_a21oi_1 _20080_ (.A1(_12082_),
    .A2(net32),
    .Y(_00565_),
    .B1(_02928_));
 sg13g2_nor2b_1 _20081_ (.A(_02860_),
    .B_N(\cpu.dcache.r_data[7][2] ),
    .Y(_02929_));
 sg13g2_a21oi_1 _20082_ (.A1(net972),
    .A2(_02860_),
    .Y(_02930_),
    .B1(_02929_));
 sg13g2_nand2_1 _20083_ (.Y(_02931_),
    .A(_02709_),
    .B(net63));
 sg13g2_o21ai_1 _20084_ (.B1(_02931_),
    .Y(_00566_),
    .A1(_02858_),
    .A2(_02930_));
 sg13g2_mux2_1 _20085_ (.A0(\cpu.dcache.r_data[7][30] ),
    .A1(_12045_),
    .S(_02924_),
    .X(_02932_));
 sg13g2_nor2_1 _20086_ (.A(_02908_),
    .B(_02932_),
    .Y(_02933_));
 sg13g2_a21oi_1 _20087_ (.A1(_12089_),
    .A2(net32),
    .Y(_00567_),
    .B1(_02933_));
 sg13g2_mux2_1 _20088_ (.A0(\cpu.dcache.r_data[7][31] ),
    .A1(_12062_),
    .S(_02924_),
    .X(_02934_));
 sg13g2_nor2_1 _20089_ (.A(_02908_),
    .B(_02934_),
    .Y(_02935_));
 sg13g2_a21oi_1 _20090_ (.A1(_12095_),
    .A2(net32),
    .Y(_00568_),
    .B1(_02935_));
 sg13g2_nor2b_1 _20091_ (.A(_02860_),
    .B_N(\cpu.dcache.r_data[7][3] ),
    .Y(_02936_));
 sg13g2_a21oi_1 _20092_ (.A1(net971),
    .A2(_02860_),
    .Y(_02937_),
    .B1(_02936_));
 sg13g2_nand2_1 _20093_ (.Y(_02938_),
    .A(_12716_),
    .B(_02857_));
 sg13g2_o21ai_1 _20094_ (.B1(_02938_),
    .Y(_00569_),
    .A1(_02858_),
    .A2(_02937_));
 sg13g2_or2_1 _20095_ (.X(_02939_),
    .B(_12188_),
    .A(net466));
 sg13g2_buf_1 _20096_ (.A(_02939_),
    .X(_02940_));
 sg13g2_mux2_1 _20097_ (.A0(net1091),
    .A1(\cpu.dcache.r_data[7][4] ),
    .S(_02940_),
    .X(_02941_));
 sg13g2_mux2_1 _20098_ (.A0(_02941_),
    .A1(_12130_),
    .S(net63),
    .X(_00570_));
 sg13g2_mux2_1 _20099_ (.A0(net1090),
    .A1(\cpu.dcache.r_data[7][5] ),
    .S(_02940_),
    .X(_02942_));
 sg13g2_mux2_1 _20100_ (.A0(_02942_),
    .A1(net990),
    .S(net63),
    .X(_00571_));
 sg13g2_mux2_1 _20101_ (.A0(net1089),
    .A1(\cpu.dcache.r_data[7][6] ),
    .S(_02940_),
    .X(_02943_));
 sg13g2_mux2_1 _20102_ (.A0(_02943_),
    .A1(net989),
    .S(net63),
    .X(_00572_));
 sg13g2_mux2_1 _20103_ (.A0(net1088),
    .A1(\cpu.dcache.r_data[7][7] ),
    .S(_02940_),
    .X(_02944_));
 sg13g2_mux2_1 _20104_ (.A0(_02944_),
    .A1(net851),
    .S(net63),
    .X(_00573_));
 sg13g2_nor2b_1 _20105_ (.A(_02868_),
    .B_N(\cpu.dcache.r_data[7][8] ),
    .Y(_02945_));
 sg13g2_a21oi_1 _20106_ (.A1(net970),
    .A2(_02868_),
    .Y(_02946_),
    .B1(_02945_));
 sg13g2_nand2_1 _20107_ (.Y(_02947_),
    .A(_12150_),
    .B(_02865_));
 sg13g2_o21ai_1 _20108_ (.B1(_02947_),
    .Y(_00574_),
    .A1(net33),
    .A2(_02946_));
 sg13g2_nor2b_1 _20109_ (.A(_02868_),
    .B_N(\cpu.dcache.r_data[7][9] ),
    .Y(_02948_));
 sg13g2_a21oi_1 _20110_ (.A1(net973),
    .A2(_02868_),
    .Y(_02949_),
    .B1(_02948_));
 sg13g2_nand2_1 _20111_ (.Y(_02950_),
    .A(_12160_),
    .B(_02865_));
 sg13g2_o21ai_1 _20112_ (.B1(_02950_),
    .Y(_00575_),
    .A1(net33),
    .A2(_02949_));
 sg13g2_and2_1 _20113_ (.A(_11542_),
    .B(_12001_),
    .X(_02951_));
 sg13g2_buf_1 _20114_ (.A(_09209_),
    .X(_02952_));
 sg13g2_buf_1 _20115_ (.A(\cpu.d_rstrobe_d ),
    .X(_02953_));
 sg13g2_nor2_1 _20116_ (.A(_02952_),
    .B(_02953_),
    .Y(_02954_));
 sg13g2_nand4_1 _20117_ (.B(_12025_),
    .C(_09211_),
    .A(_09824_),
    .Y(_02955_),
    .D(_02954_));
 sg13g2_nand2b_1 _20118_ (.Y(_02956_),
    .B(_02955_),
    .A_N(_02951_));
 sg13g2_buf_2 _20119_ (.A(_02956_),
    .X(_02957_));
 sg13g2_and2_1 _20120_ (.A(net994),
    .B(_12007_),
    .X(_02958_));
 sg13g2_xor2_1 _20121_ (.B(_12025_),
    .A(_02953_),
    .X(_02959_));
 sg13g2_a21oi_1 _20122_ (.A1(_02958_),
    .A2(_02959_),
    .Y(_02960_),
    .B1(_02951_));
 sg13g2_buf_2 _20123_ (.A(_02960_),
    .X(_02961_));
 sg13g2_nor2_1 _20124_ (.A(net603),
    .B(_02961_),
    .Y(_02962_));
 sg13g2_mux2_1 _20125_ (.A0(\cpu.dcache.r_dirty[0] ),
    .A1(_02957_),
    .S(_02962_),
    .X(_00576_));
 sg13g2_nor2_1 _20126_ (.A(_12212_),
    .B(_02961_),
    .Y(_02963_));
 sg13g2_mux2_1 _20127_ (.A0(\cpu.dcache.r_dirty[1] ),
    .A1(_02957_),
    .S(_02963_),
    .X(_00577_));
 sg13g2_nor2_1 _20128_ (.A(_12347_),
    .B(_02961_),
    .Y(_02964_));
 sg13g2_mux2_1 _20129_ (.A0(\cpu.dcache.r_dirty[2] ),
    .A1(_02957_),
    .S(_02964_),
    .X(_00578_));
 sg13g2_nor2_1 _20130_ (.A(net528),
    .B(_02961_),
    .Y(_02965_));
 sg13g2_mux2_1 _20131_ (.A0(\cpu.dcache.r_dirty[3] ),
    .A1(_02957_),
    .S(_02965_),
    .X(_00579_));
 sg13g2_nor2_1 _20132_ (.A(net600),
    .B(_02961_),
    .Y(_02966_));
 sg13g2_mux2_1 _20133_ (.A0(\cpu.dcache.r_dirty[4] ),
    .A1(_02957_),
    .S(_02966_),
    .X(_00580_));
 sg13g2_nor2_1 _20134_ (.A(_12668_),
    .B(_02961_),
    .Y(_02967_));
 sg13g2_mux2_1 _20135_ (.A0(\cpu.dcache.r_dirty[5] ),
    .A1(_02957_),
    .S(_02967_),
    .X(_00581_));
 sg13g2_nor2_1 _20136_ (.A(_02740_),
    .B(_02961_),
    .Y(_02968_));
 sg13g2_mux2_1 _20137_ (.A0(\cpu.dcache.r_dirty[6] ),
    .A1(_02957_),
    .S(_02968_),
    .X(_00582_));
 sg13g2_nor2_1 _20138_ (.A(_02856_),
    .B(_02961_),
    .Y(_02969_));
 sg13g2_mux2_1 _20139_ (.A0(\cpu.dcache.r_dirty[7] ),
    .A1(_02957_),
    .S(_02969_),
    .X(_00583_));
 sg13g2_buf_1 _20140_ (.A(net862),
    .X(_02970_));
 sg13g2_buf_1 _20141_ (.A(net730),
    .X(_02971_));
 sg13g2_buf_1 _20142_ (.A(net469),
    .X(_02972_));
 sg13g2_buf_1 _20143_ (.A(net469),
    .X(_02973_));
 sg13g2_nand2_1 _20144_ (.Y(_02974_),
    .A(\cpu.dcache.r_tag[0][5] ),
    .B(net404));
 sg13g2_o21ai_1 _20145_ (.B1(_02974_),
    .Y(_00587_),
    .A1(net652),
    .A2(net405));
 sg13g2_mux2_1 _20146_ (.A0(net415),
    .A1(\cpu.dcache.r_tag[0][15] ),
    .S(net405),
    .X(_00588_));
 sg13g2_mux2_1 _20147_ (.A0(net416),
    .A1(\cpu.dcache.r_tag[0][16] ),
    .S(_02972_),
    .X(_00589_));
 sg13g2_mux2_1 _20148_ (.A0(net380),
    .A1(\cpu.dcache.r_tag[0][17] ),
    .S(net405),
    .X(_00590_));
 sg13g2_mux2_1 _20149_ (.A0(net377),
    .A1(\cpu.dcache.r_tag[0][18] ),
    .S(net405),
    .X(_00591_));
 sg13g2_mux2_1 _20150_ (.A0(net417),
    .A1(\cpu.dcache.r_tag[0][19] ),
    .S(_02972_),
    .X(_00592_));
 sg13g2_mux2_1 _20151_ (.A0(_09728_),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .S(net405),
    .X(_00593_));
 sg13g2_mux2_1 _20152_ (.A0(_09799_),
    .A1(\cpu.dcache.r_tag[0][21] ),
    .S(net405),
    .X(_00594_));
 sg13g2_mux2_1 _20153_ (.A0(net376),
    .A1(\cpu.dcache.r_tag[0][22] ),
    .S(net404),
    .X(_00595_));
 sg13g2_inv_1 _20154_ (.Y(_02975_),
    .A(net378));
 sg13g2_nand2_1 _20155_ (.Y(_02976_),
    .A(\cpu.dcache.r_tag[0][23] ),
    .B(net469));
 sg13g2_o21ai_1 _20156_ (.B1(_02976_),
    .Y(_00596_),
    .A1(_02975_),
    .A2(net405));
 sg13g2_buf_1 _20157_ (.A(net1028),
    .X(_02977_));
 sg13g2_buf_1 _20158_ (.A(net847),
    .X(_02978_));
 sg13g2_mux2_1 _20159_ (.A0(net729),
    .A1(\cpu.dcache.r_tag[0][6] ),
    .S(_02973_),
    .X(_00597_));
 sg13g2_buf_1 _20160_ (.A(_10974_),
    .X(_02979_));
 sg13g2_buf_1 _20161_ (.A(net846),
    .X(_02980_));
 sg13g2_nand2_1 _20162_ (.Y(_02981_),
    .A(\cpu.dcache.r_tag[0][7] ),
    .B(_12147_));
 sg13g2_o21ai_1 _20163_ (.B1(_02981_),
    .Y(_00598_),
    .A1(_02980_),
    .A2(net405));
 sg13g2_buf_1 _20164_ (.A(net1043),
    .X(_02982_));
 sg13g2_buf_1 _20165_ (.A(net845),
    .X(_02983_));
 sg13g2_mux2_1 _20166_ (.A0(_02983_),
    .A1(\cpu.dcache.r_tag[0][8] ),
    .S(net404),
    .X(_00599_));
 sg13g2_buf_1 _20167_ (.A(_11085_),
    .X(_02984_));
 sg13g2_buf_1 _20168_ (.A(net969),
    .X(_02985_));
 sg13g2_mux2_1 _20169_ (.A0(_02985_),
    .A1(\cpu.dcache.r_tag[0][9] ),
    .S(net404),
    .X(_00600_));
 sg13g2_buf_1 _20170_ (.A(net1104),
    .X(_02986_));
 sg13g2_buf_1 _20171_ (.A(net968),
    .X(_02987_));
 sg13g2_mux2_1 _20172_ (.A0(_02987_),
    .A1(\cpu.dcache.r_tag[0][10] ),
    .S(net404),
    .X(_00601_));
 sg13g2_buf_1 _20173_ (.A(net1107),
    .X(_02988_));
 sg13g2_buf_1 _20174_ (.A(net967),
    .X(_02989_));
 sg13g2_mux2_1 _20175_ (.A0(_02989_),
    .A1(\cpu.dcache.r_tag[0][11] ),
    .S(net404),
    .X(_00602_));
 sg13g2_mux2_1 _20176_ (.A0(_09464_),
    .A1(\cpu.dcache.r_tag[0][12] ),
    .S(net404),
    .X(_00603_));
 sg13g2_mux2_1 _20177_ (.A0(net381),
    .A1(\cpu.dcache.r_tag[0][13] ),
    .S(_02973_),
    .X(_00604_));
 sg13g2_mux2_1 _20178_ (.A0(_09553_),
    .A1(\cpu.dcache.r_tag[0][14] ),
    .S(net404),
    .X(_00605_));
 sg13g2_buf_2 _20179_ (.A(net735),
    .X(_02990_));
 sg13g2_buf_1 _20180_ (.A(net651),
    .X(_02991_));
 sg13g2_buf_1 _20181_ (.A(net598),
    .X(_02992_));
 sg13g2_buf_1 _20182_ (.A(net529),
    .X(_02993_));
 sg13g2_mux2_1 _20183_ (.A0(\cpu.dcache.r_tag[1][5] ),
    .A1(net524),
    .S(net465),
    .X(_00606_));
 sg13g2_mux2_1 _20184_ (.A0(\cpu.dcache.r_tag[1][15] ),
    .A1(net415),
    .S(net465),
    .X(_00607_));
 sg13g2_mux2_1 _20185_ (.A0(\cpu.dcache.r_tag[1][16] ),
    .A1(net416),
    .S(_02993_),
    .X(_00608_));
 sg13g2_mux2_1 _20186_ (.A0(\cpu.dcache.r_tag[1][17] ),
    .A1(_09513_),
    .S(net465),
    .X(_00609_));
 sg13g2_mux2_1 _20187_ (.A0(\cpu.dcache.r_tag[1][18] ),
    .A1(net377),
    .S(net465),
    .X(_00610_));
 sg13g2_mux2_1 _20188_ (.A0(\cpu.dcache.r_tag[1][19] ),
    .A1(net417),
    .S(net465),
    .X(_00611_));
 sg13g2_mux2_1 _20189_ (.A0(\cpu.dcache.r_tag[1][20] ),
    .A1(net414),
    .S(net465),
    .X(_00612_));
 sg13g2_mux2_1 _20190_ (.A0(\cpu.dcache.r_tag[1][21] ),
    .A1(net375),
    .S(net465),
    .X(_00613_));
 sg13g2_mux2_1 _20191_ (.A0(\cpu.dcache.r_tag[1][22] ),
    .A1(net376),
    .S(_02993_),
    .X(_00614_));
 sg13g2_mux2_1 _20192_ (.A0(\cpu.dcache.r_tag[1][23] ),
    .A1(net378),
    .S(net465),
    .X(_00615_));
 sg13g2_buf_1 _20193_ (.A(net847),
    .X(_02994_));
 sg13g2_buf_1 _20194_ (.A(net529),
    .X(_02995_));
 sg13g2_mux2_1 _20195_ (.A0(\cpu.dcache.r_tag[1][6] ),
    .A1(net726),
    .S(_02995_),
    .X(_00616_));
 sg13g2_buf_1 _20196_ (.A(net1042),
    .X(_02996_));
 sg13g2_buf_1 _20197_ (.A(net841),
    .X(_02997_));
 sg13g2_mux2_1 _20198_ (.A0(\cpu.dcache.r_tag[1][7] ),
    .A1(net725),
    .S(net464),
    .X(_00617_));
 sg13g2_buf_1 _20199_ (.A(net845),
    .X(_02998_));
 sg13g2_mux2_1 _20200_ (.A0(\cpu.dcache.r_tag[1][8] ),
    .A1(net724),
    .S(net464),
    .X(_00618_));
 sg13g2_buf_1 _20201_ (.A(net969),
    .X(_02999_));
 sg13g2_mux2_1 _20202_ (.A0(\cpu.dcache.r_tag[1][9] ),
    .A1(net840),
    .S(net464),
    .X(_00619_));
 sg13g2_buf_1 _20203_ (.A(net968),
    .X(_03000_));
 sg13g2_mux2_1 _20204_ (.A0(\cpu.dcache.r_tag[1][10] ),
    .A1(net839),
    .S(net464),
    .X(_00620_));
 sg13g2_buf_1 _20205_ (.A(net967),
    .X(_03001_));
 sg13g2_mux2_1 _20206_ (.A0(\cpu.dcache.r_tag[1][11] ),
    .A1(net838),
    .S(net464),
    .X(_00621_));
 sg13g2_mux2_1 _20207_ (.A0(\cpu.dcache.r_tag[1][12] ),
    .A1(net382),
    .S(net464),
    .X(_00622_));
 sg13g2_mux2_1 _20208_ (.A0(\cpu.dcache.r_tag[1][13] ),
    .A1(net381),
    .S(_02995_),
    .X(_00623_));
 sg13g2_mux2_1 _20209_ (.A0(\cpu.dcache.r_tag[1][14] ),
    .A1(net379),
    .S(net464),
    .X(_00624_));
 sg13g2_buf_1 _20210_ (.A(net367),
    .X(_03002_));
 sg13g2_mux2_1 _20211_ (.A0(\cpu.dcache.r_tag[2][5] ),
    .A1(net524),
    .S(net334),
    .X(_00625_));
 sg13g2_mux2_1 _20212_ (.A0(\cpu.dcache.r_tag[2][15] ),
    .A1(net415),
    .S(net334),
    .X(_00626_));
 sg13g2_mux2_1 _20213_ (.A0(\cpu.dcache.r_tag[2][16] ),
    .A1(net416),
    .S(_03002_),
    .X(_00627_));
 sg13g2_mux2_1 _20214_ (.A0(\cpu.dcache.r_tag[2][17] ),
    .A1(net380),
    .S(net334),
    .X(_00628_));
 sg13g2_mux2_1 _20215_ (.A0(\cpu.dcache.r_tag[2][18] ),
    .A1(net377),
    .S(net334),
    .X(_00629_));
 sg13g2_mux2_1 _20216_ (.A0(\cpu.dcache.r_tag[2][19] ),
    .A1(net417),
    .S(_03002_),
    .X(_00630_));
 sg13g2_mux2_1 _20217_ (.A0(\cpu.dcache.r_tag[2][20] ),
    .A1(net414),
    .S(net334),
    .X(_00631_));
 sg13g2_mux2_1 _20218_ (.A0(\cpu.dcache.r_tag[2][21] ),
    .A1(net375),
    .S(net334),
    .X(_00632_));
 sg13g2_mux2_1 _20219_ (.A0(\cpu.dcache.r_tag[2][22] ),
    .A1(net376),
    .S(net334),
    .X(_00633_));
 sg13g2_mux2_1 _20220_ (.A0(\cpu.dcache.r_tag[2][23] ),
    .A1(net378),
    .S(net334),
    .X(_00634_));
 sg13g2_buf_1 _20221_ (.A(net367),
    .X(_03003_));
 sg13g2_mux2_1 _20222_ (.A0(\cpu.dcache.r_tag[2][6] ),
    .A1(net726),
    .S(_03003_),
    .X(_00635_));
 sg13g2_mux2_1 _20223_ (.A0(\cpu.dcache.r_tag[2][7] ),
    .A1(net725),
    .S(net333),
    .X(_00636_));
 sg13g2_mux2_1 _20224_ (.A0(\cpu.dcache.r_tag[2][8] ),
    .A1(net724),
    .S(net333),
    .X(_00637_));
 sg13g2_mux2_1 _20225_ (.A0(\cpu.dcache.r_tag[2][9] ),
    .A1(net840),
    .S(net333),
    .X(_00638_));
 sg13g2_mux2_1 _20226_ (.A0(\cpu.dcache.r_tag[2][10] ),
    .A1(net839),
    .S(net333),
    .X(_00639_));
 sg13g2_mux2_1 _20227_ (.A0(\cpu.dcache.r_tag[2][11] ),
    .A1(net838),
    .S(net333),
    .X(_00640_));
 sg13g2_mux2_1 _20228_ (.A0(\cpu.dcache.r_tag[2][12] ),
    .A1(net382),
    .S(net333),
    .X(_00641_));
 sg13g2_mux2_1 _20229_ (.A0(\cpu.dcache.r_tag[2][13] ),
    .A1(net381),
    .S(_03003_),
    .X(_00642_));
 sg13g2_mux2_1 _20230_ (.A0(\cpu.dcache.r_tag[2][14] ),
    .A1(net379),
    .S(net333),
    .X(_00643_));
 sg13g2_buf_1 _20231_ (.A(_12521_),
    .X(_03004_));
 sg13g2_mux2_1 _20232_ (.A0(\cpu.dcache.r_tag[3][5] ),
    .A1(net524),
    .S(net403),
    .X(_00644_));
 sg13g2_mux2_1 _20233_ (.A0(\cpu.dcache.r_tag[3][15] ),
    .A1(net415),
    .S(net403),
    .X(_00645_));
 sg13g2_mux2_1 _20234_ (.A0(\cpu.dcache.r_tag[3][16] ),
    .A1(net416),
    .S(net403),
    .X(_00646_));
 sg13g2_mux2_1 _20235_ (.A0(\cpu.dcache.r_tag[3][17] ),
    .A1(net380),
    .S(net403),
    .X(_00647_));
 sg13g2_mux2_1 _20236_ (.A0(\cpu.dcache.r_tag[3][18] ),
    .A1(_09754_),
    .S(net403),
    .X(_00648_));
 sg13g2_mux2_1 _20237_ (.A0(\cpu.dcache.r_tag[3][19] ),
    .A1(net417),
    .S(_03004_),
    .X(_00649_));
 sg13g2_mux2_1 _20238_ (.A0(\cpu.dcache.r_tag[3][20] ),
    .A1(net414),
    .S(net403),
    .X(_00650_));
 sg13g2_mux2_1 _20239_ (.A0(\cpu.dcache.r_tag[3][21] ),
    .A1(net375),
    .S(net403),
    .X(_00651_));
 sg13g2_mux2_1 _20240_ (.A0(\cpu.dcache.r_tag[3][22] ),
    .A1(net376),
    .S(_03004_),
    .X(_00652_));
 sg13g2_mux2_1 _20241_ (.A0(\cpu.dcache.r_tag[3][23] ),
    .A1(_09640_),
    .S(net403),
    .X(_00653_));
 sg13g2_buf_1 _20242_ (.A(_12521_),
    .X(_03005_));
 sg13g2_mux2_1 _20243_ (.A0(\cpu.dcache.r_tag[3][6] ),
    .A1(net726),
    .S(_03005_),
    .X(_00654_));
 sg13g2_mux2_1 _20244_ (.A0(\cpu.dcache.r_tag[3][7] ),
    .A1(net725),
    .S(net402),
    .X(_00655_));
 sg13g2_mux2_1 _20245_ (.A0(\cpu.dcache.r_tag[3][8] ),
    .A1(net724),
    .S(net402),
    .X(_00656_));
 sg13g2_mux2_1 _20246_ (.A0(\cpu.dcache.r_tag[3][9] ),
    .A1(_02999_),
    .S(_03005_),
    .X(_00657_));
 sg13g2_mux2_1 _20247_ (.A0(\cpu.dcache.r_tag[3][10] ),
    .A1(net839),
    .S(net402),
    .X(_00658_));
 sg13g2_mux2_1 _20248_ (.A0(\cpu.dcache.r_tag[3][11] ),
    .A1(net838),
    .S(net402),
    .X(_00659_));
 sg13g2_mux2_1 _20249_ (.A0(\cpu.dcache.r_tag[3][12] ),
    .A1(net382),
    .S(net402),
    .X(_00660_));
 sg13g2_mux2_1 _20250_ (.A0(\cpu.dcache.r_tag[3][13] ),
    .A1(_09489_),
    .S(net402),
    .X(_00661_));
 sg13g2_mux2_1 _20251_ (.A0(\cpu.dcache.r_tag[3][14] ),
    .A1(net379),
    .S(net402),
    .X(_00662_));
 sg13g2_buf_1 _20252_ (.A(net527),
    .X(_03006_));
 sg13g2_nand2_1 _20253_ (.Y(_03007_),
    .A(\cpu.dcache.r_tag[4][5] ),
    .B(net527));
 sg13g2_o21ai_1 _20254_ (.B1(_03007_),
    .Y(_00663_),
    .A1(_02971_),
    .A2(net463));
 sg13g2_mux2_1 _20255_ (.A0(net415),
    .A1(\cpu.dcache.r_tag[4][15] ),
    .S(net463),
    .X(_00664_));
 sg13g2_mux2_1 _20256_ (.A0(net416),
    .A1(\cpu.dcache.r_tag[4][16] ),
    .S(net463),
    .X(_00665_));
 sg13g2_mux2_1 _20257_ (.A0(net380),
    .A1(\cpu.dcache.r_tag[4][17] ),
    .S(net463),
    .X(_00666_));
 sg13g2_mux2_1 _20258_ (.A0(net377),
    .A1(\cpu.dcache.r_tag[4][18] ),
    .S(net463),
    .X(_00667_));
 sg13g2_mux2_1 _20259_ (.A0(net417),
    .A1(\cpu.dcache.r_tag[4][19] ),
    .S(net463),
    .X(_00668_));
 sg13g2_mux2_1 _20260_ (.A0(net414),
    .A1(\cpu.dcache.r_tag[4][20] ),
    .S(_03006_),
    .X(_00669_));
 sg13g2_buf_1 _20261_ (.A(net527),
    .X(_03008_));
 sg13g2_mux2_1 _20262_ (.A0(net375),
    .A1(\cpu.dcache.r_tag[4][21] ),
    .S(net462),
    .X(_00670_));
 sg13g2_mux2_1 _20263_ (.A0(net376),
    .A1(\cpu.dcache.r_tag[4][22] ),
    .S(net462),
    .X(_00671_));
 sg13g2_nand2_1 _20264_ (.Y(_03009_),
    .A(\cpu.dcache.r_tag[4][23] ),
    .B(net527));
 sg13g2_o21ai_1 _20265_ (.B1(_03009_),
    .Y(_00672_),
    .A1(_02975_),
    .A2(_03006_));
 sg13g2_mux2_1 _20266_ (.A0(_02978_),
    .A1(\cpu.dcache.r_tag[4][6] ),
    .S(_03008_),
    .X(_00673_));
 sg13g2_nand2_1 _20267_ (.Y(_03010_),
    .A(\cpu.dcache.r_tag[4][7] ),
    .B(_12624_));
 sg13g2_o21ai_1 _20268_ (.B1(_03010_),
    .Y(_00674_),
    .A1(_02980_),
    .A2(net463));
 sg13g2_mux2_1 _20269_ (.A0(net727),
    .A1(\cpu.dcache.r_tag[4][8] ),
    .S(net462),
    .X(_00675_));
 sg13g2_mux2_1 _20270_ (.A0(_02985_),
    .A1(\cpu.dcache.r_tag[4][9] ),
    .S(net462),
    .X(_00676_));
 sg13g2_mux2_1 _20271_ (.A0(_02987_),
    .A1(\cpu.dcache.r_tag[4][10] ),
    .S(_03008_),
    .X(_00677_));
 sg13g2_mux2_1 _20272_ (.A0(net842),
    .A1(\cpu.dcache.r_tag[4][11] ),
    .S(net462),
    .X(_00678_));
 sg13g2_mux2_1 _20273_ (.A0(net382),
    .A1(\cpu.dcache.r_tag[4][12] ),
    .S(net462),
    .X(_00679_));
 sg13g2_mux2_1 _20274_ (.A0(net381),
    .A1(\cpu.dcache.r_tag[4][13] ),
    .S(net462),
    .X(_00680_));
 sg13g2_mux2_1 _20275_ (.A0(net379),
    .A1(\cpu.dcache.r_tag[4][14] ),
    .S(net462),
    .X(_00681_));
 sg13g2_buf_1 _20276_ (.A(_02689_),
    .X(_03011_));
 sg13g2_mux2_1 _20277_ (.A0(\cpu.dcache.r_tag[5][5] ),
    .A1(net524),
    .S(net461),
    .X(_00682_));
 sg13g2_mux2_1 _20278_ (.A0(\cpu.dcache.r_tag[5][15] ),
    .A1(_09713_),
    .S(net461),
    .X(_00683_));
 sg13g2_mux2_1 _20279_ (.A0(\cpu.dcache.r_tag[5][16] ),
    .A1(_09686_),
    .S(net461),
    .X(_00684_));
 sg13g2_mux2_1 _20280_ (.A0(\cpu.dcache.r_tag[5][17] ),
    .A1(_09513_),
    .S(net461),
    .X(_00685_));
 sg13g2_mux2_1 _20281_ (.A0(\cpu.dcache.r_tag[5][18] ),
    .A1(net377),
    .S(net461),
    .X(_00686_));
 sg13g2_mux2_1 _20282_ (.A0(\cpu.dcache.r_tag[5][19] ),
    .A1(_09665_),
    .S(_03011_),
    .X(_00687_));
 sg13g2_mux2_1 _20283_ (.A0(\cpu.dcache.r_tag[5][20] ),
    .A1(net414),
    .S(net461),
    .X(_00688_));
 sg13g2_mux2_1 _20284_ (.A0(\cpu.dcache.r_tag[5][21] ),
    .A1(net375),
    .S(net461),
    .X(_00689_));
 sg13g2_mux2_1 _20285_ (.A0(\cpu.dcache.r_tag[5][22] ),
    .A1(net376),
    .S(_03011_),
    .X(_00690_));
 sg13g2_mux2_1 _20286_ (.A0(\cpu.dcache.r_tag[5][23] ),
    .A1(net378),
    .S(net461),
    .X(_00691_));
 sg13g2_buf_1 _20287_ (.A(_02689_),
    .X(_03012_));
 sg13g2_mux2_1 _20288_ (.A0(\cpu.dcache.r_tag[5][6] ),
    .A1(_02994_),
    .S(_03012_),
    .X(_00692_));
 sg13g2_mux2_1 _20289_ (.A0(\cpu.dcache.r_tag[5][7] ),
    .A1(net725),
    .S(net460),
    .X(_00693_));
 sg13g2_mux2_1 _20290_ (.A0(\cpu.dcache.r_tag[5][8] ),
    .A1(_02998_),
    .S(net460),
    .X(_00694_));
 sg13g2_mux2_1 _20291_ (.A0(\cpu.dcache.r_tag[5][9] ),
    .A1(_02999_),
    .S(net460),
    .X(_00695_));
 sg13g2_mux2_1 _20292_ (.A0(\cpu.dcache.r_tag[5][10] ),
    .A1(_03000_),
    .S(net460),
    .X(_00696_));
 sg13g2_mux2_1 _20293_ (.A0(\cpu.dcache.r_tag[5][11] ),
    .A1(_03001_),
    .S(net460),
    .X(_00697_));
 sg13g2_mux2_1 _20294_ (.A0(\cpu.dcache.r_tag[5][12] ),
    .A1(_09464_),
    .S(net460),
    .X(_00698_));
 sg13g2_mux2_1 _20295_ (.A0(\cpu.dcache.r_tag[5][13] ),
    .A1(net381),
    .S(_03012_),
    .X(_00699_));
 sg13g2_mux2_1 _20296_ (.A0(\cpu.dcache.r_tag[5][14] ),
    .A1(net379),
    .S(net460),
    .X(_00700_));
 sg13g2_buf_1 _20297_ (.A(_02805_),
    .X(_03013_));
 sg13g2_mux2_1 _20298_ (.A0(\cpu.dcache.r_tag[6][5] ),
    .A1(net524),
    .S(net401),
    .X(_00701_));
 sg13g2_mux2_1 _20299_ (.A0(\cpu.dcache.r_tag[6][15] ),
    .A1(net415),
    .S(net401),
    .X(_00702_));
 sg13g2_mux2_1 _20300_ (.A0(\cpu.dcache.r_tag[6][16] ),
    .A1(net416),
    .S(net401),
    .X(_00703_));
 sg13g2_mux2_1 _20301_ (.A0(\cpu.dcache.r_tag[6][17] ),
    .A1(net380),
    .S(net401),
    .X(_00704_));
 sg13g2_mux2_1 _20302_ (.A0(\cpu.dcache.r_tag[6][18] ),
    .A1(net377),
    .S(net401),
    .X(_00705_));
 sg13g2_mux2_1 _20303_ (.A0(\cpu.dcache.r_tag[6][19] ),
    .A1(net417),
    .S(_03013_),
    .X(_00706_));
 sg13g2_mux2_1 _20304_ (.A0(\cpu.dcache.r_tag[6][20] ),
    .A1(net414),
    .S(net401),
    .X(_00707_));
 sg13g2_mux2_1 _20305_ (.A0(\cpu.dcache.r_tag[6][21] ),
    .A1(net375),
    .S(net401),
    .X(_00708_));
 sg13g2_mux2_1 _20306_ (.A0(\cpu.dcache.r_tag[6][22] ),
    .A1(_09776_),
    .S(_03013_),
    .X(_00709_));
 sg13g2_mux2_1 _20307_ (.A0(\cpu.dcache.r_tag[6][23] ),
    .A1(net378),
    .S(net401),
    .X(_00710_));
 sg13g2_buf_1 _20308_ (.A(_02805_),
    .X(_03014_));
 sg13g2_mux2_1 _20309_ (.A0(\cpu.dcache.r_tag[6][6] ),
    .A1(_02994_),
    .S(net400),
    .X(_00711_));
 sg13g2_mux2_1 _20310_ (.A0(\cpu.dcache.r_tag[6][7] ),
    .A1(net725),
    .S(net400),
    .X(_00712_));
 sg13g2_mux2_1 _20311_ (.A0(\cpu.dcache.r_tag[6][8] ),
    .A1(net724),
    .S(net400),
    .X(_00713_));
 sg13g2_mux2_1 _20312_ (.A0(\cpu.dcache.r_tag[6][9] ),
    .A1(net840),
    .S(_03014_),
    .X(_00714_));
 sg13g2_mux2_1 _20313_ (.A0(\cpu.dcache.r_tag[6][10] ),
    .A1(_03000_),
    .S(_03014_),
    .X(_00715_));
 sg13g2_mux2_1 _20314_ (.A0(\cpu.dcache.r_tag[6][11] ),
    .A1(_03001_),
    .S(net400),
    .X(_00716_));
 sg13g2_mux2_1 _20315_ (.A0(\cpu.dcache.r_tag[6][12] ),
    .A1(net382),
    .S(net400),
    .X(_00717_));
 sg13g2_mux2_1 _20316_ (.A0(\cpu.dcache.r_tag[6][13] ),
    .A1(_09489_),
    .S(net400),
    .X(_00718_));
 sg13g2_mux2_1 _20317_ (.A0(\cpu.dcache.r_tag[6][14] ),
    .A1(net379),
    .S(net400),
    .X(_00719_));
 sg13g2_buf_1 _20318_ (.A(_02911_),
    .X(_03015_));
 sg13g2_mux2_1 _20319_ (.A0(\cpu.dcache.r_tag[7][5] ),
    .A1(net524),
    .S(net366),
    .X(_00720_));
 sg13g2_mux2_1 _20320_ (.A0(\cpu.dcache.r_tag[7][15] ),
    .A1(net415),
    .S(net366),
    .X(_00721_));
 sg13g2_mux2_1 _20321_ (.A0(\cpu.dcache.r_tag[7][16] ),
    .A1(net416),
    .S(net366),
    .X(_00722_));
 sg13g2_mux2_1 _20322_ (.A0(\cpu.dcache.r_tag[7][17] ),
    .A1(net380),
    .S(net366),
    .X(_00723_));
 sg13g2_mux2_1 _20323_ (.A0(\cpu.dcache.r_tag[7][18] ),
    .A1(net377),
    .S(net366),
    .X(_00724_));
 sg13g2_mux2_1 _20324_ (.A0(\cpu.dcache.r_tag[7][19] ),
    .A1(net417),
    .S(_03015_),
    .X(_00725_));
 sg13g2_mux2_1 _20325_ (.A0(\cpu.dcache.r_tag[7][20] ),
    .A1(net414),
    .S(net366),
    .X(_00726_));
 sg13g2_mux2_1 _20326_ (.A0(\cpu.dcache.r_tag[7][21] ),
    .A1(net375),
    .S(net366),
    .X(_00727_));
 sg13g2_mux2_1 _20327_ (.A0(\cpu.dcache.r_tag[7][22] ),
    .A1(net376),
    .S(_03015_),
    .X(_00728_));
 sg13g2_mux2_1 _20328_ (.A0(\cpu.dcache.r_tag[7][23] ),
    .A1(_09640_),
    .S(net366),
    .X(_00729_));
 sg13g2_buf_1 _20329_ (.A(_02977_),
    .X(_03016_));
 sg13g2_buf_1 _20330_ (.A(_02911_),
    .X(_03017_));
 sg13g2_mux2_1 _20331_ (.A0(\cpu.dcache.r_tag[7][6] ),
    .A1(net723),
    .S(net365),
    .X(_00730_));
 sg13g2_mux2_1 _20332_ (.A0(\cpu.dcache.r_tag[7][7] ),
    .A1(net725),
    .S(net365),
    .X(_00731_));
 sg13g2_buf_1 _20333_ (.A(net845),
    .X(_03018_));
 sg13g2_mux2_1 _20334_ (.A0(\cpu.dcache.r_tag[7][8] ),
    .A1(net722),
    .S(net365),
    .X(_00732_));
 sg13g2_buf_1 _20335_ (.A(net969),
    .X(_03019_));
 sg13g2_mux2_1 _20336_ (.A0(\cpu.dcache.r_tag[7][9] ),
    .A1(net837),
    .S(net365),
    .X(_00733_));
 sg13g2_buf_1 _20337_ (.A(net968),
    .X(_03020_));
 sg13g2_mux2_1 _20338_ (.A0(\cpu.dcache.r_tag[7][10] ),
    .A1(net836),
    .S(net365),
    .X(_00734_));
 sg13g2_buf_1 _20339_ (.A(net967),
    .X(_03021_));
 sg13g2_mux2_1 _20340_ (.A0(\cpu.dcache.r_tag[7][11] ),
    .A1(net835),
    .S(_03017_),
    .X(_00735_));
 sg13g2_mux2_1 _20341_ (.A0(\cpu.dcache.r_tag[7][12] ),
    .A1(net382),
    .S(net365),
    .X(_00736_));
 sg13g2_mux2_1 _20342_ (.A0(\cpu.dcache.r_tag[7][13] ),
    .A1(net381),
    .S(net365),
    .X(_00737_));
 sg13g2_mux2_1 _20343_ (.A0(\cpu.dcache.r_tag[7][14] ),
    .A1(_09553_),
    .S(_03017_),
    .X(_00738_));
 sg13g2_buf_1 _20344_ (.A(net223),
    .X(_03022_));
 sg13g2_buf_1 _20345_ (.A(_08420_),
    .X(_03023_));
 sg13g2_nand2_1 _20346_ (.Y(_03024_),
    .A(net284),
    .B(net291));
 sg13g2_buf_2 _20347_ (.A(_03024_),
    .X(_03025_));
 sg13g2_nand2_1 _20348_ (.Y(_03026_),
    .A(_09040_),
    .B(_09042_));
 sg13g2_buf_2 _20349_ (.A(_03026_),
    .X(_03027_));
 sg13g2_o21ai_1 _20350_ (.B1(_03027_),
    .Y(_03028_),
    .A1(net187),
    .A2(_03025_));
 sg13g2_buf_1 _20351_ (.A(_08377_),
    .X(_03029_));
 sg13g2_nand2_2 _20352_ (.Y(_03030_),
    .A(_08354_),
    .B(net236));
 sg13g2_nor2_1 _20353_ (.A(_09048_),
    .B(_03030_),
    .Y(_03031_));
 sg13g2_a21oi_1 _20354_ (.A1(net195),
    .A2(_03028_),
    .Y(_03032_),
    .B1(_03031_));
 sg13g2_nor2_1 _20355_ (.A(_11525_),
    .B(_09000_),
    .Y(_03033_));
 sg13g2_a21oi_1 _20356_ (.A1(net107),
    .A2(_03032_),
    .Y(_00747_),
    .B1(_03033_));
 sg13g2_buf_1 _20357_ (.A(net1125),
    .X(_03034_));
 sg13g2_buf_1 _20358_ (.A(net966),
    .X(_03035_));
 sg13g2_a21oi_1 _20359_ (.A1(_08313_),
    .A2(_09025_),
    .Y(_03036_),
    .B1(_09033_));
 sg13g2_buf_1 _20360_ (.A(_03036_),
    .X(_03037_));
 sg13g2_buf_1 _20361_ (.A(_03037_),
    .X(_03038_));
 sg13g2_buf_1 _20362_ (.A(_09042_),
    .X(_03039_));
 sg13g2_nor2_2 _20363_ (.A(net236),
    .B(net282),
    .Y(_03040_));
 sg13g2_nor2_1 _20364_ (.A(net284),
    .B(_08437_),
    .Y(_03041_));
 sg13g2_a21oi_1 _20365_ (.A1(net283),
    .A2(_03040_),
    .Y(_03042_),
    .B1(_03041_));
 sg13g2_buf_1 _20366_ (.A(net291),
    .X(_03043_));
 sg13g2_buf_2 _20367_ (.A(net236),
    .X(_03044_));
 sg13g2_buf_1 _20368_ (.A(net284),
    .X(_03045_));
 sg13g2_buf_1 _20369_ (.A(net234),
    .X(_03046_));
 sg13g2_buf_1 _20370_ (.A(net209),
    .X(_03047_));
 sg13g2_buf_1 _20371_ (.A(net292),
    .X(_03048_));
 sg13g2_nor2_1 _20372_ (.A(net236),
    .B(net233),
    .Y(_03049_));
 sg13g2_a21oi_1 _20373_ (.A1(net210),
    .A2(net186),
    .Y(_03050_),
    .B1(_03049_));
 sg13g2_buf_1 _20374_ (.A(_08354_),
    .X(_03051_));
 sg13g2_buf_1 _20375_ (.A(net208),
    .X(_03052_));
 sg13g2_buf_1 _20376_ (.A(net233),
    .X(_03053_));
 sg13g2_buf_1 _20377_ (.A(_08438_),
    .X(_03054_));
 sg13g2_o21ai_1 _20378_ (.B1(net206),
    .Y(_03055_),
    .A1(net185),
    .A2(net207));
 sg13g2_a22oi_1 _20379_ (.Y(_03056_),
    .B1(_03055_),
    .B2(net210),
    .A2(_03050_),
    .A1(net235));
 sg13g2_o21ai_1 _20380_ (.B1(_03056_),
    .Y(_03057_),
    .A1(net195),
    .A2(_03042_));
 sg13g2_mux2_1 _20381_ (.A0(_03035_),
    .A1(_03057_),
    .S(net119),
    .X(_00748_));
 sg13g2_inv_1 _20382_ (.Y(_03058_),
    .A(\cpu.cond[1] ));
 sg13g2_nor2_2 _20383_ (.A(_08354_),
    .B(_08377_),
    .Y(_03059_));
 sg13g2_nor2_1 _20384_ (.A(_08404_),
    .B(net284),
    .Y(_03060_));
 sg13g2_buf_1 _20385_ (.A(_03060_),
    .X(_03061_));
 sg13g2_nand3_1 _20386_ (.B(_03059_),
    .C(net205),
    .A(net118),
    .Y(_03062_));
 sg13g2_o21ai_1 _20387_ (.B1(_03062_),
    .Y(_00749_),
    .A1(_03058_),
    .A2(net106));
 sg13g2_buf_1 _20388_ (.A(_09046_),
    .X(_03063_));
 sg13g2_nor2_1 _20389_ (.A(net195),
    .B(net184),
    .Y(_03064_));
 sg13g2_o21ai_1 _20390_ (.B1(net210),
    .Y(_03065_),
    .A1(net185),
    .A2(_03027_));
 sg13g2_nor2_1 _20391_ (.A(_03064_),
    .B(_03065_),
    .Y(_03066_));
 sg13g2_mux2_1 _20392_ (.A0(\cpu.cond[2] ),
    .A1(_03066_),
    .S(net119),
    .X(_00750_));
 sg13g2_or3_1 _20393_ (.A(net89),
    .B(_09106_),
    .C(_09916_),
    .X(_03067_));
 sg13g2_o21ai_1 _20394_ (.B1(_03067_),
    .Y(_00751_),
    .A1(_09368_),
    .A2(net106));
 sg13g2_buf_1 _20395_ (.A(_08404_),
    .X(_03068_));
 sg13g2_nand2_2 _20396_ (.Y(_03069_),
    .A(net232),
    .B(_09046_));
 sg13g2_nand2b_1 _20397_ (.Y(_03070_),
    .B(_08344_),
    .A_N(_00177_));
 sg13g2_mux2_1 _20398_ (.A0(\cpu.icache.r_data[7][25] ),
    .A1(\cpu.icache.r_data[3][25] ),
    .S(_08366_),
    .X(_03071_));
 sg13g2_a22oi_1 _20399_ (.Y(_03072_),
    .B1(_03071_),
    .B2(net792),
    .A2(net697),
    .A1(\cpu.icache.r_data[6][25] ));
 sg13g2_nand2b_1 _20400_ (.Y(_03073_),
    .B(_08338_),
    .A_N(_03072_));
 sg13g2_a22oi_1 _20401_ (.Y(_03074_),
    .B1(net547),
    .B2(\cpu.icache.r_data[2][25] ),
    .A2(net633),
    .A1(\cpu.icache.r_data[4][25] ));
 sg13g2_a22oi_1 _20402_ (.Y(_03075_),
    .B1(net555),
    .B2(\cpu.icache.r_data[5][25] ),
    .A2(net635),
    .A1(\cpu.icache.r_data[1][25] ));
 sg13g2_nand4_1 _20403_ (.B(_03073_),
    .C(_03074_),
    .A(_03070_),
    .Y(_03076_),
    .D(_03075_));
 sg13g2_nand2_1 _20404_ (.Y(_03077_),
    .A(_00176_),
    .B(_08344_));
 sg13g2_mux2_1 _20405_ (.A0(\cpu.icache.r_data[7][9] ),
    .A1(\cpu.icache.r_data[3][9] ),
    .S(net924),
    .X(_03078_));
 sg13g2_a22oi_1 _20406_ (.Y(_03079_),
    .B1(net704),
    .B2(_03078_),
    .A2(_08314_),
    .A1(\cpu.icache.r_data[4][9] ));
 sg13g2_a22oi_1 _20407_ (.Y(_03080_),
    .B1(_08348_),
    .B2(\cpu.icache.r_data[2][9] ),
    .A2(net641),
    .A1(\cpu.icache.r_data[1][9] ));
 sg13g2_a22oi_1 _20408_ (.Y(_03081_),
    .B1(net634),
    .B2(\cpu.icache.r_data[5][9] ),
    .A2(_08326_),
    .A1(\cpu.icache.r_data[6][9] ));
 sg13g2_nand4_1 _20409_ (.B(_03079_),
    .C(_03080_),
    .A(net549),
    .Y(_03082_),
    .D(_03081_));
 sg13g2_a21o_1 _20410_ (.A2(_03082_),
    .A1(_03077_),
    .B1(_08312_),
    .X(_03083_));
 sg13g2_o21ai_1 _20411_ (.B1(_03083_),
    .Y(_03084_),
    .A1(net923),
    .A2(_03076_));
 sg13g2_buf_1 _20412_ (.A(_03084_),
    .X(_03085_));
 sg13g2_a22oi_1 _20413_ (.Y(_03086_),
    .B1(net638),
    .B2(\cpu.icache.r_data[5][7] ),
    .A2(net699),
    .A1(\cpu.icache.r_data[4][7] ));
 sg13g2_a22oi_1 _20414_ (.Y(_03087_),
    .B1(net640),
    .B2(\cpu.icache.r_data[2][7] ),
    .A2(net700),
    .A1(\cpu.icache.r_data[1][7] ));
 sg13g2_mux2_1 _20415_ (.A0(\cpu.icache.r_data[7][7] ),
    .A1(\cpu.icache.r_data[3][7] ),
    .S(net1071),
    .X(_03088_));
 sg13g2_a22oi_1 _20416_ (.Y(_03089_),
    .B1(_03088_),
    .B2(_08397_),
    .A2(net795),
    .A1(\cpu.icache.r_data[6][7] ));
 sg13g2_nand2b_1 _20417_ (.Y(_03090_),
    .B(net698),
    .A_N(_03089_));
 sg13g2_and4_1 _20418_ (.A(net550),
    .B(_03086_),
    .C(_03087_),
    .D(_03090_),
    .X(_03091_));
 sg13g2_a21oi_1 _20419_ (.A1(_00172_),
    .A2(net483),
    .Y(_03092_),
    .B1(_03091_));
 sg13g2_nor2_1 _20420_ (.A(_00173_),
    .B(net550),
    .Y(_03093_));
 sg13g2_mux2_1 _20421_ (.A0(\cpu.icache.r_data[4][23] ),
    .A1(\cpu.icache.r_data[6][23] ),
    .S(net797),
    .X(_03094_));
 sg13g2_a22oi_1 _20422_ (.Y(_03095_),
    .B1(_03094_),
    .B2(net930),
    .A2(net704),
    .A1(\cpu.icache.r_data[7][23] ));
 sg13g2_nor2_1 _20423_ (.A(net786),
    .B(_03095_),
    .Y(_03096_));
 sg13g2_a22oi_1 _20424_ (.Y(_03097_),
    .B1(net481),
    .B2(\cpu.icache.r_data[3][23] ),
    .A2(net552),
    .A1(\cpu.icache.r_data[2][23] ));
 sg13g2_a22oi_1 _20425_ (.Y(_03098_),
    .B1(net634),
    .B2(\cpu.icache.r_data[5][23] ),
    .A2(net641),
    .A1(\cpu.icache.r_data[1][23] ));
 sg13g2_nand2_1 _20426_ (.Y(_03099_),
    .A(_03097_),
    .B(_03098_));
 sg13g2_or4_1 _20427_ (.A(net923),
    .B(_03093_),
    .C(_03096_),
    .D(_03099_),
    .X(_03100_));
 sg13g2_o21ai_1 _20428_ (.B1(_03100_),
    .Y(_03101_),
    .A1(net926),
    .A2(_03092_));
 sg13g2_buf_1 _20429_ (.A(_03101_),
    .X(_03102_));
 sg13g2_nand3_1 _20430_ (.B(_03085_),
    .C(_03102_),
    .A(_08311_),
    .Y(_03103_));
 sg13g2_buf_1 _20431_ (.A(_03103_),
    .X(_03104_));
 sg13g2_inv_1 _20432_ (.Y(_03105_),
    .A(_00174_));
 sg13g2_a22oi_1 _20433_ (.Y(_03106_),
    .B1(net555),
    .B2(\cpu.icache.r_data[5][8] ),
    .A2(net635),
    .A1(\cpu.icache.r_data[1][8] ));
 sg13g2_a22oi_1 _20434_ (.Y(_03107_),
    .B1(net481),
    .B2(\cpu.icache.r_data[3][8] ),
    .A2(net556),
    .A1(\cpu.icache.r_data[2][8] ));
 sg13g2_mux2_1 _20435_ (.A0(\cpu.icache.r_data[4][8] ),
    .A1(\cpu.icache.r_data[6][8] ),
    .S(net931),
    .X(_03108_));
 sg13g2_a22oi_1 _20436_ (.Y(_03109_),
    .B1(_03108_),
    .B2(net930),
    .A2(_08315_),
    .A1(\cpu.icache.r_data[7][8] ));
 sg13g2_or2_1 _20437_ (.X(_03110_),
    .B(_03109_),
    .A(net786));
 sg13g2_nand4_1 _20438_ (.B(_03106_),
    .C(_03107_),
    .A(net554),
    .Y(_03111_),
    .D(_03110_));
 sg13g2_o21ai_1 _20439_ (.B1(_03111_),
    .Y(_03112_),
    .A1(_03105_),
    .A2(net482));
 sg13g2_nor2_1 _20440_ (.A(_00175_),
    .B(_08333_),
    .Y(_03113_));
 sg13g2_mux2_1 _20441_ (.A0(\cpu.icache.r_data[4][24] ),
    .A1(\cpu.icache.r_data[6][24] ),
    .S(net793),
    .X(_03114_));
 sg13g2_a22oi_1 _20442_ (.Y(_03115_),
    .B1(_03114_),
    .B2(net930),
    .A2(_08315_),
    .A1(\cpu.icache.r_data[7][24] ));
 sg13g2_nor2_1 _20443_ (.A(net786),
    .B(_03115_),
    .Y(_03116_));
 sg13g2_a22oi_1 _20444_ (.Y(_03117_),
    .B1(net547),
    .B2(\cpu.icache.r_data[2][24] ),
    .A2(net548),
    .A1(\cpu.icache.r_data[1][24] ));
 sg13g2_a22oi_1 _20445_ (.Y(_03118_),
    .B1(net555),
    .B2(\cpu.icache.r_data[5][24] ),
    .A2(net481),
    .A1(\cpu.icache.r_data[3][24] ));
 sg13g2_nand2_1 _20446_ (.Y(_03119_),
    .A(_03117_),
    .B(_03118_));
 sg13g2_nor4_1 _20447_ (.A(_08390_),
    .B(_03113_),
    .C(_03116_),
    .D(_03119_),
    .Y(_03120_));
 sg13g2_a21oi_1 _20448_ (.A1(_08390_),
    .A2(_03112_),
    .Y(_03121_),
    .B1(_03120_));
 sg13g2_buf_1 _20449_ (.A(_03121_),
    .X(_03122_));
 sg13g2_or3_1 _20450_ (.A(_08458_),
    .B(_03104_),
    .C(net231),
    .X(_03123_));
 sg13g2_or2_1 _20451_ (.X(_03124_),
    .B(_03123_),
    .A(_09051_));
 sg13g2_buf_1 _20452_ (.A(_03124_),
    .X(_03125_));
 sg13g2_or3_1 _20453_ (.A(_09106_),
    .B(_03069_),
    .C(_03125_),
    .X(_03126_));
 sg13g2_buf_1 _20454_ (.A(_03126_),
    .X(_03127_));
 sg13g2_nor3_1 _20455_ (.A(_09093_),
    .B(net221),
    .C(_03127_),
    .Y(_03128_));
 sg13g2_mux2_1 _20456_ (.A0(\cpu.dec.do_flush_all ),
    .A1(_03128_),
    .S(net105),
    .X(_00752_));
 sg13g2_nand2_1 _20457_ (.Y(_03129_),
    .A(net221),
    .B(_09905_));
 sg13g2_nor2_1 _20458_ (.A(_09109_),
    .B(_03129_),
    .Y(_03130_));
 sg13g2_mux2_1 _20459_ (.A0(\cpu.dec.do_flush_write ),
    .A1(_03130_),
    .S(_09918_),
    .X(_00753_));
 sg13g2_nand2_1 _20460_ (.Y(_03131_),
    .A(_03059_),
    .B(_03069_));
 sg13g2_buf_2 _20461_ (.A(_03131_),
    .X(_03132_));
 sg13g2_nor2_1 _20462_ (.A(_09177_),
    .B(_03129_),
    .Y(_03133_));
 sg13g2_nor2_1 _20463_ (.A(_09048_),
    .B(_03133_),
    .Y(_03134_));
 sg13g2_nor2_2 _20464_ (.A(_08404_),
    .B(_03025_),
    .Y(_03135_));
 sg13g2_a22oi_1 _20465_ (.Y(_03136_),
    .B1(_03135_),
    .B2(net290),
    .A2(_03134_),
    .A1(net244));
 sg13g2_buf_1 _20466_ (.A(_08437_),
    .X(_03137_));
 sg13g2_buf_1 _20467_ (.A(net230),
    .X(_03138_));
 sg13g2_buf_1 _20468_ (.A(net204),
    .X(_03139_));
 sg13g2_and4_1 _20469_ (.A(net172),
    .B(net183),
    .C(net244),
    .D(_03027_),
    .X(_03140_));
 sg13g2_buf_1 _20470_ (.A(net232),
    .X(_03141_));
 sg13g2_nand2_1 _20471_ (.Y(_03142_),
    .A(net203),
    .B(_03059_));
 sg13g2_nor3_1 _20472_ (.A(net206),
    .B(net243),
    .C(_03142_),
    .Y(_03143_));
 sg13g2_nor2_1 _20473_ (.A(net209),
    .B(_09092_),
    .Y(_03144_));
 sg13g2_buf_1 _20474_ (.A(net232),
    .X(_03145_));
 sg13g2_nand3_1 _20475_ (.B(net209),
    .C(net290),
    .A(net202),
    .Y(_03146_));
 sg13g2_nor2b_1 _20476_ (.A(_03144_),
    .B_N(_03146_),
    .Y(_03147_));
 sg13g2_nor3_1 _20477_ (.A(net183),
    .B(_03030_),
    .C(_03147_),
    .Y(_03148_));
 sg13g2_buf_1 _20478_ (.A(_03039_),
    .X(_03149_));
 sg13g2_nor2_1 _20479_ (.A(_08437_),
    .B(_09171_),
    .Y(_03150_));
 sg13g2_nand2_1 _20480_ (.Y(_03151_),
    .A(net229),
    .B(_03150_));
 sg13g2_nand2_1 _20481_ (.Y(_03152_),
    .A(net292),
    .B(net291));
 sg13g2_nand3_1 _20482_ (.B(net289),
    .C(_03152_),
    .A(net209),
    .Y(_03153_));
 sg13g2_nand2_1 _20483_ (.Y(_03154_),
    .A(_08354_),
    .B(_08379_));
 sg13g2_buf_1 _20484_ (.A(_03154_),
    .X(_03155_));
 sg13g2_a21oi_1 _20485_ (.A1(_03151_),
    .A2(_03153_),
    .Y(_03156_),
    .B1(_03155_));
 sg13g2_nor4_1 _20486_ (.A(_03140_),
    .B(_03143_),
    .C(_03148_),
    .D(_03156_),
    .Y(_03157_));
 sg13g2_o21ai_1 _20487_ (.B1(_03157_),
    .Y(_03158_),
    .A1(_03132_),
    .A2(_03136_));
 sg13g2_mux2_1 _20488_ (.A0(_11008_),
    .A1(_03158_),
    .S(_09918_),
    .X(_00754_));
 sg13g2_nand2_1 _20489_ (.Y(_03159_),
    .A(net284),
    .B(_03150_));
 sg13g2_inv_1 _20490_ (.Y(_03160_),
    .A(_03159_));
 sg13g2_nand2_1 _20491_ (.Y(_03161_),
    .A(_03137_),
    .B(_09126_));
 sg13g2_nand2_1 _20492_ (.Y(_03162_),
    .A(net291),
    .B(net246));
 sg13g2_a21oi_1 _20493_ (.A1(_03161_),
    .A2(_03162_),
    .Y(_03163_),
    .B1(_03023_));
 sg13g2_o21ai_1 _20494_ (.B1(net232),
    .Y(_03164_),
    .A1(_03160_),
    .A2(_03163_));
 sg13g2_nor2_1 _20495_ (.A(net230),
    .B(_03085_),
    .Y(_03165_));
 sg13g2_nor2_1 _20496_ (.A(_08404_),
    .B(_09042_),
    .Y(_03166_));
 sg13g2_nand2_1 _20497_ (.Y(_03167_),
    .A(_03165_),
    .B(_03166_));
 sg13g2_nand3_1 _20498_ (.B(_03164_),
    .C(_03167_),
    .A(net223),
    .Y(_03168_));
 sg13g2_nand2_2 _20499_ (.Y(_03169_),
    .A(_08440_),
    .B(net221));
 sg13g2_nor2_1 _20500_ (.A(net291),
    .B(_09091_),
    .Y(_03170_));
 sg13g2_a21oi_1 _20501_ (.A1(_09044_),
    .A2(_09035_),
    .Y(_03171_),
    .B1(_03170_));
 sg13g2_nand2_1 _20502_ (.Y(_03172_),
    .A(_09042_),
    .B(_03171_));
 sg13g2_nand2_1 _20503_ (.Y(_03173_),
    .A(net284),
    .B(_03165_));
 sg13g2_nand4_1 _20504_ (.B(_03169_),
    .C(_03172_),
    .A(_08377_),
    .Y(_03174_),
    .D(_03173_));
 sg13g2_and3_1 _20505_ (.X(_03175_),
    .A(_03051_),
    .B(_03168_),
    .C(_03174_));
 sg13g2_buf_2 _20506_ (.A(_03175_),
    .X(_03176_));
 sg13g2_nor2_1 _20507_ (.A(_03132_),
    .B(_03167_),
    .Y(_03177_));
 sg13g2_nand2_1 _20508_ (.Y(_03178_),
    .A(_08404_),
    .B(_08437_));
 sg13g2_buf_2 _20509_ (.A(_03178_),
    .X(_03179_));
 sg13g2_o21ai_1 _20510_ (.B1(_08380_),
    .Y(_03180_),
    .A1(_09126_),
    .A2(_03179_));
 sg13g2_buf_1 _20511_ (.A(_03180_),
    .X(_03181_));
 sg13g2_nor2_2 _20512_ (.A(net282),
    .B(net204),
    .Y(_03182_));
 sg13g2_inv_1 _20513_ (.Y(_03183_),
    .A(_03179_));
 sg13g2_a21oi_1 _20514_ (.A1(_03182_),
    .A2(_03122_),
    .Y(_03184_),
    .B1(_03183_));
 sg13g2_nor2_1 _20515_ (.A(net140),
    .B(_03184_),
    .Y(_03185_));
 sg13g2_nand2_1 _20516_ (.Y(_03186_),
    .A(_03037_),
    .B(_03060_));
 sg13g2_nor3_1 _20517_ (.A(net292),
    .B(net284),
    .C(_03137_),
    .Y(_03187_));
 sg13g2_buf_2 _20518_ (.A(_03187_),
    .X(_03188_));
 sg13g2_nand2_1 _20519_ (.Y(_03189_),
    .A(net221),
    .B(_03188_));
 sg13g2_a22oi_1 _20520_ (.Y(_03190_),
    .B1(_03186_),
    .B2(_03189_),
    .A2(_03181_),
    .A1(_03132_));
 sg13g2_nor4_1 _20521_ (.A(_03176_),
    .B(_03177_),
    .C(_03185_),
    .D(_03190_),
    .Y(_03191_));
 sg13g2_nor2_1 _20522_ (.A(\cpu.dec.imm[10] ),
    .B(net118),
    .Y(_03192_));
 sg13g2_a21oi_1 _20523_ (.A1(net107),
    .A2(_03191_),
    .Y(_00755_),
    .B1(_03192_));
 sg13g2_and2_1 _20524_ (.A(_03167_),
    .B(_03186_),
    .X(_03193_));
 sg13g2_buf_2 _20525_ (.A(_03193_),
    .X(_03194_));
 sg13g2_nand2_1 _20526_ (.Y(_03195_),
    .A(net244),
    .B(_03188_));
 sg13g2_a21oi_1 _20527_ (.A1(_03194_),
    .A2(_03195_),
    .Y(_03196_),
    .B1(_09175_));
 sg13g2_nor2_2 _20528_ (.A(net292),
    .B(_03023_),
    .Y(_03197_));
 sg13g2_o21ai_1 _20529_ (.B1(net235),
    .Y(_03198_),
    .A1(net293),
    .A2(_03197_));
 sg13g2_buf_1 _20530_ (.A(net292),
    .X(_03199_));
 sg13g2_o21ai_1 _20531_ (.B1(net228),
    .Y(_03200_),
    .A1(_09046_),
    .A2(net293));
 sg13g2_nand2_1 _20532_ (.Y(_03201_),
    .A(_03198_),
    .B(_03200_));
 sg13g2_inv_2 _20533_ (.Y(_03202_),
    .A(net231));
 sg13g2_nor2_1 _20534_ (.A(_03104_),
    .B(_03202_),
    .Y(_03203_));
 sg13g2_buf_1 _20535_ (.A(_03203_),
    .X(_03204_));
 sg13g2_nand2_1 _20536_ (.Y(_03205_),
    .A(net291),
    .B(_03197_));
 sg13g2_buf_1 _20537_ (.A(_03205_),
    .X(_03206_));
 sg13g2_a21oi_1 _20538_ (.A1(net220),
    .A2(_03203_),
    .Y(_03207_),
    .B1(_03206_));
 sg13g2_buf_1 _20539_ (.A(_03207_),
    .X(_03208_));
 sg13g2_o21ai_1 _20540_ (.B1(_03208_),
    .Y(_03209_),
    .A1(net244),
    .A2(net139));
 sg13g2_a21oi_1 _20541_ (.A1(_03201_),
    .A2(_03209_),
    .Y(_03210_),
    .B1(net140));
 sg13g2_nor3_1 _20542_ (.A(_03176_),
    .B(_03196_),
    .C(_03210_),
    .Y(_03211_));
 sg13g2_nor2_1 _20543_ (.A(\cpu.dec.imm[11] ),
    .B(net118),
    .Y(_03212_));
 sg13g2_a21oi_1 _20544_ (.A1(net107),
    .A2(_03211_),
    .Y(_00756_),
    .B1(_03212_));
 sg13g2_nand2_1 _20545_ (.Y(_03213_),
    .A(net290),
    .B(_03188_));
 sg13g2_a21oi_1 _20546_ (.A1(_03194_),
    .A2(_03213_),
    .Y(_03214_),
    .B1(_03132_));
 sg13g2_o21ai_1 _20547_ (.B1(_03208_),
    .Y(_03215_),
    .A1(net290),
    .A2(net139));
 sg13g2_a21oi_1 _20548_ (.A1(_03201_),
    .A2(_03215_),
    .Y(_03216_),
    .B1(net140));
 sg13g2_nor3_1 _20549_ (.A(_03176_),
    .B(_03214_),
    .C(_03216_),
    .Y(_03217_));
 sg13g2_nor2_1 _20550_ (.A(\cpu.dec.imm[12] ),
    .B(net118),
    .Y(_03218_));
 sg13g2_a21oi_1 _20551_ (.A1(net107),
    .A2(_03217_),
    .Y(_00757_),
    .B1(_03218_));
 sg13g2_nor2_1 _20552_ (.A(_09051_),
    .B(_09897_),
    .Y(_03219_));
 sg13g2_buf_1 _20553_ (.A(_03219_),
    .X(_03220_));
 sg13g2_o21ai_1 _20554_ (.B1(_03194_),
    .Y(_03221_),
    .A1(net293),
    .A2(_03206_));
 sg13g2_a21oi_1 _20555_ (.A1(_03220_),
    .A2(_03221_),
    .Y(_03222_),
    .B1(_03176_));
 sg13g2_o21ai_1 _20556_ (.B1(_03208_),
    .Y(_03223_),
    .A1(_03038_),
    .A2(net139));
 sg13g2_a21o_1 _20557_ (.A2(_03223_),
    .A1(_03201_),
    .B1(net140),
    .X(_03224_));
 sg13g2_a21oi_1 _20558_ (.A1(_03222_),
    .A2(_03224_),
    .Y(_03225_),
    .B1(net89));
 sg13g2_a21o_1 _20559_ (.A2(net79),
    .A1(\cpu.dec.imm[13] ),
    .B1(_03225_),
    .X(_00758_));
 sg13g2_nand2_1 _20560_ (.Y(_03226_),
    .A(net295),
    .B(_03188_));
 sg13g2_a21o_1 _20561_ (.A2(_03226_),
    .A1(_03194_),
    .B1(_03132_),
    .X(_03227_));
 sg13g2_o21ai_1 _20562_ (.B1(_03208_),
    .Y(_03228_),
    .A1(_08460_),
    .A2(net139));
 sg13g2_a21oi_1 _20563_ (.A1(_03201_),
    .A2(_03228_),
    .Y(_03229_),
    .B1(net140));
 sg13g2_nor3_1 _20564_ (.A(_09015_),
    .B(_03176_),
    .C(_03229_),
    .Y(_03230_));
 sg13g2_a22oi_1 _20565_ (.Y(_00759_),
    .B1(_03227_),
    .B2(_03230_),
    .A2(net79),
    .A1(_11446_));
 sg13g2_o21ai_1 _20566_ (.B1(_03194_),
    .Y(_03231_),
    .A1(_08460_),
    .A2(_03206_));
 sg13g2_nand2_1 _20567_ (.Y(_03232_),
    .A(_03220_),
    .B(_03231_));
 sg13g2_a22oi_1 _20568_ (.Y(_00760_),
    .B1(_03230_),
    .B2(_03232_),
    .A2(net79),
    .A1(_11417_));
 sg13g2_buf_2 _20569_ (.A(_09014_),
    .X(_03233_));
 sg13g2_nor2_1 _20570_ (.A(net292),
    .B(_03025_),
    .Y(_03234_));
 sg13g2_buf_2 _20571_ (.A(_03234_),
    .X(_03235_));
 sg13g2_nand2_1 _20572_ (.Y(_03236_),
    .A(net236),
    .B(_03235_));
 sg13g2_mux2_1 _20573_ (.A0(_08311_),
    .A1(_09072_),
    .S(_03236_),
    .X(_03237_));
 sg13g2_a21oi_1 _20574_ (.A1(_09042_),
    .A2(_03203_),
    .Y(_03238_),
    .B1(net230));
 sg13g2_o21ai_1 _20575_ (.B1(net206),
    .Y(_03239_),
    .A1(net233),
    .A2(_03238_));
 sg13g2_nand2_1 _20576_ (.Y(_03240_),
    .A(_03027_),
    .B(_03025_));
 sg13g2_a22oi_1 _20577_ (.Y(_03241_),
    .B1(_03240_),
    .B2(net219),
    .A2(_03239_),
    .A1(net290));
 sg13g2_nor2_1 _20578_ (.A(net291),
    .B(_09072_),
    .Y(_03242_));
 sg13g2_nor2_1 _20579_ (.A(_08310_),
    .B(net230),
    .Y(_03243_));
 sg13g2_a21oi_1 _20580_ (.A1(net230),
    .A2(_09072_),
    .Y(_03244_),
    .B1(_03243_));
 sg13g2_nand2_1 _20581_ (.Y(_03245_),
    .A(net230),
    .B(net246));
 sg13g2_o21ai_1 _20582_ (.B1(_03245_),
    .Y(_03246_),
    .A1(net230),
    .A2(_09072_));
 sg13g2_mux4_1 _20583_ (.S0(_03068_),
    .A0(_09162_),
    .A1(_03242_),
    .A2(_03244_),
    .A3(_03246_),
    .S1(_03045_),
    .X(_03247_));
 sg13g2_nand2_1 _20584_ (.Y(_03248_),
    .A(net223),
    .B(_03247_));
 sg13g2_o21ai_1 _20585_ (.B1(_03248_),
    .Y(_03249_),
    .A1(_03022_),
    .A2(_03241_));
 sg13g2_nand2_1 _20586_ (.Y(_03250_),
    .A(_09893_),
    .B(_03249_));
 sg13g2_o21ai_1 _20587_ (.B1(_03250_),
    .Y(_03251_),
    .A1(_09893_),
    .A2(_03237_));
 sg13g2_nand2_1 _20588_ (.Y(_03252_),
    .A(net98),
    .B(_03251_));
 sg13g2_o21ai_1 _20589_ (.B1(_03252_),
    .Y(_00761_),
    .A1(_10521_),
    .A2(net106));
 sg13g2_nor2_1 _20590_ (.A(_03043_),
    .B(net219),
    .Y(_03253_));
 sg13g2_nor3_1 _20591_ (.A(net229),
    .B(_03243_),
    .C(_03253_),
    .Y(_03254_));
 sg13g2_nor2_1 _20592_ (.A(_03144_),
    .B(_03254_),
    .Y(_03255_));
 sg13g2_nand2b_1 _20593_ (.Y(_03256_),
    .B(_03235_),
    .A_N(net295));
 sg13g2_o21ai_1 _20594_ (.B1(_03256_),
    .Y(_03257_),
    .A1(net288),
    .A2(_03235_));
 sg13g2_o21ai_1 _20595_ (.B1(_03045_),
    .Y(_03258_),
    .A1(net204),
    .A2(net336));
 sg13g2_nand2_1 _20596_ (.Y(_03259_),
    .A(net282),
    .B(_09127_));
 sg13g2_o21ai_1 _20597_ (.B1(_03259_),
    .Y(_03260_),
    .A1(_03253_),
    .A2(_03258_));
 sg13g2_inv_1 _20598_ (.Y(_03261_),
    .A(_03161_));
 sg13g2_or2_1 _20599_ (.X(_03262_),
    .B(_03041_),
    .A(_09046_));
 sg13g2_buf_1 _20600_ (.A(_03262_),
    .X(_03263_));
 sg13g2_inv_1 _20601_ (.Y(_03264_),
    .A(_03263_));
 sg13g2_a22oi_1 _20602_ (.Y(_03265_),
    .B1(_03264_),
    .B2(net288),
    .A2(_03261_),
    .A1(net209));
 sg13g2_nor2_1 _20603_ (.A(net207),
    .B(_03265_),
    .Y(_03266_));
 sg13g2_a21oi_1 _20604_ (.A1(net207),
    .A2(_03260_),
    .Y(_03267_),
    .B1(_03266_));
 sg13g2_nor2_1 _20605_ (.A(net222),
    .B(_03206_),
    .Y(_03268_));
 sg13g2_o21ai_1 _20606_ (.B1(_03259_),
    .Y(_03269_),
    .A1(net229),
    .A2(_03245_));
 sg13g2_o21ai_1 _20607_ (.B1(_03159_),
    .Y(_03270_),
    .A1(_08311_),
    .A2(_03179_));
 sg13g2_a221oi_1 _20608_ (.B2(_03053_),
    .C1(_03270_),
    .B1(_03269_),
    .A1(_03268_),
    .Y(_03271_),
    .A2(net139));
 sg13g2_mux4_1 _20609_ (.S0(_03044_),
    .A0(_03255_),
    .A1(_03257_),
    .A2(_03267_),
    .A3(_03271_),
    .S1(net195),
    .X(_03272_));
 sg13g2_nand2_1 _20610_ (.Y(_03273_),
    .A(_10500_),
    .B(net89));
 sg13g2_o21ai_1 _20611_ (.B1(_03273_),
    .Y(_00762_),
    .A1(net79),
    .A2(_03272_));
 sg13g2_nor2b_1 _20612_ (.A(_09177_),
    .B_N(_09905_),
    .Y(_03274_));
 sg13g2_nand3_1 _20613_ (.B(net235),
    .C(_03037_),
    .A(net234),
    .Y(_03275_));
 sg13g2_o21ai_1 _20614_ (.B1(_03275_),
    .Y(_03276_),
    .A1(_08311_),
    .A2(net209));
 sg13g2_nand2_1 _20615_ (.Y(_03277_),
    .A(net204),
    .B(net336));
 sg13g2_a21oi_1 _20616_ (.A1(_03258_),
    .A2(_03277_),
    .Y(_03278_),
    .B1(net228));
 sg13g2_a21oi_1 _20617_ (.A1(net207),
    .A2(_03276_),
    .Y(_03279_),
    .B1(_03278_));
 sg13g2_o21ai_1 _20618_ (.B1(_03279_),
    .Y(_03280_),
    .A1(_03169_),
    .A2(_03274_));
 sg13g2_nand2_1 _20619_ (.Y(_03281_),
    .A(net222),
    .B(_09897_));
 sg13g2_nand3_1 _20620_ (.B(_03280_),
    .C(_03281_),
    .A(_03059_),
    .Y(_03282_));
 sg13g2_nor2_1 _20621_ (.A(net195),
    .B(net223),
    .Y(_03283_));
 sg13g2_buf_2 _20622_ (.A(_03283_),
    .X(_03284_));
 sg13g2_nor2_1 _20623_ (.A(net336),
    .B(_03235_),
    .Y(_03285_));
 sg13g2_a21oi_1 _20624_ (.A1(net293),
    .A2(_03235_),
    .Y(_03286_),
    .B1(_03285_));
 sg13g2_nand2_1 _20625_ (.Y(_03287_),
    .A(net172),
    .B(_03183_));
 sg13g2_o21ai_1 _20626_ (.B1(_03287_),
    .Y(_03288_),
    .A1(net184),
    .A2(_03155_));
 sg13g2_nor3_1 _20627_ (.A(_03054_),
    .B(net220),
    .C(_03155_),
    .Y(_03289_));
 sg13g2_a221oi_1 _20628_ (.B2(net295),
    .C1(_03289_),
    .B1(_03288_),
    .A1(_03284_),
    .Y(_03290_),
    .A2(_03286_));
 sg13g2_a22oi_1 _20629_ (.Y(_03291_),
    .B1(_03182_),
    .B2(net244),
    .A2(_03060_),
    .A1(_09097_));
 sg13g2_nand3_1 _20630_ (.B(_03188_),
    .C(net139),
    .A(net295),
    .Y(_03292_));
 sg13g2_nand3_1 _20631_ (.B(_03291_),
    .C(_03292_),
    .A(_03169_),
    .Y(_03293_));
 sg13g2_nand3_1 _20632_ (.B(_03179_),
    .C(_03293_),
    .A(_08381_),
    .Y(_03294_));
 sg13g2_nand3_1 _20633_ (.B(_03290_),
    .C(_03294_),
    .A(_03282_),
    .Y(_03295_));
 sg13g2_mux2_1 _20634_ (.A0(_10465_),
    .A1(_03295_),
    .S(net105),
    .X(_00763_));
 sg13g2_mux2_1 _20635_ (.A0(net293),
    .A1(net222),
    .S(_03235_),
    .X(_03296_));
 sg13g2_a22oi_1 _20636_ (.Y(_03297_),
    .B1(net289),
    .B2(_03182_),
    .A2(net336),
    .A1(net282));
 sg13g2_nand2_1 _20637_ (.Y(_03298_),
    .A(net283),
    .B(_03134_));
 sg13g2_o21ai_1 _20638_ (.B1(_03298_),
    .Y(_03299_),
    .A1(_03141_),
    .A2(_03297_));
 sg13g2_nand2_1 _20639_ (.Y(_03300_),
    .A(net187),
    .B(net293));
 sg13g2_nand2_1 _20640_ (.Y(_03301_),
    .A(_03138_),
    .B(net293));
 sg13g2_o21ai_1 _20641_ (.B1(_03301_),
    .Y(_03302_),
    .A1(_03139_),
    .A2(net336));
 sg13g2_o21ai_1 _20642_ (.B1(net283),
    .Y(_03303_),
    .A1(net183),
    .A2(net139));
 sg13g2_o21ai_1 _20643_ (.B1(net172),
    .Y(_03304_),
    .A1(net336),
    .A2(_03027_));
 sg13g2_a221oi_1 _20644_ (.B2(_03197_),
    .C1(_03304_),
    .B1(_03303_),
    .A1(net186),
    .Y(_03305_),
    .A2(_03302_));
 sg13g2_a221oi_1 _20645_ (.B2(_03052_),
    .C1(_03305_),
    .B1(_03300_),
    .A1(_03220_),
    .Y(_03306_),
    .A2(_03299_));
 sg13g2_a21oi_1 _20646_ (.A1(_03284_),
    .A2(_03296_),
    .Y(_03307_),
    .B1(_03306_));
 sg13g2_mux2_1 _20647_ (.A0(\cpu.dec.imm[4] ),
    .A1(_03307_),
    .S(net105),
    .X(_00764_));
 sg13g2_nand2_1 _20648_ (.Y(_03308_),
    .A(_03069_),
    .B(_03172_));
 sg13g2_mux2_1 _20649_ (.A0(net222),
    .A1(net243),
    .S(_03138_),
    .X(_03309_));
 sg13g2_nor2_2 _20650_ (.A(net230),
    .B(_03102_),
    .Y(_03310_));
 sg13g2_o21ai_1 _20651_ (.B1(_03047_),
    .Y(_03311_),
    .A1(_03199_),
    .A2(_03310_));
 sg13g2_a21oi_1 _20652_ (.A1(_03053_),
    .A2(_03309_),
    .Y(_03312_),
    .B1(_03311_));
 sg13g2_o21ai_1 _20653_ (.B1(_03281_),
    .Y(_03313_),
    .A1(_03308_),
    .A2(_03312_));
 sg13g2_nor2_1 _20654_ (.A(net243),
    .B(_03135_),
    .Y(_03314_));
 sg13g2_a21oi_1 _20655_ (.A1(net289),
    .A2(_03135_),
    .Y(_03315_),
    .B1(_03314_));
 sg13g2_nand2_1 _20656_ (.Y(_03316_),
    .A(_03029_),
    .B(_09145_));
 sg13g2_a21oi_1 _20657_ (.A1(_03051_),
    .A2(_08440_),
    .Y(_03317_),
    .B1(_03316_));
 sg13g2_o21ai_1 _20658_ (.B1(_03317_),
    .Y(_03318_),
    .A1(_03206_),
    .A2(net139));
 sg13g2_o21ai_1 _20659_ (.B1(_03318_),
    .Y(_03319_),
    .A1(_03155_),
    .A2(_03315_));
 sg13g2_nand2_1 _20660_ (.Y(_03320_),
    .A(net234),
    .B(_03310_));
 sg13g2_o21ai_1 _20661_ (.B1(_03320_),
    .Y(_03321_),
    .A1(net209),
    .A2(net243));
 sg13g2_a22oi_1 _20662_ (.Y(_03322_),
    .B1(_03321_),
    .B2(net207),
    .A2(_03134_),
    .A1(_09145_));
 sg13g2_nor2_1 _20663_ (.A(_03132_),
    .B(_03322_),
    .Y(_03323_));
 sg13g2_nor3_1 _20664_ (.A(_03284_),
    .B(_03319_),
    .C(_03323_),
    .Y(_03324_));
 sg13g2_a21oi_1 _20665_ (.A1(_03284_),
    .A2(_03313_),
    .Y(_03325_),
    .B1(_03324_));
 sg13g2_mux2_1 _20666_ (.A0(\cpu.dec.imm[5] ),
    .A1(_03325_),
    .S(_03233_),
    .X(_00765_));
 sg13g2_nand2_1 _20667_ (.Y(_03326_),
    .A(net203),
    .B(net219));
 sg13g2_a22oi_1 _20668_ (.Y(_03327_),
    .B1(_03310_),
    .B2(net186),
    .A2(_03061_),
    .A1(net244));
 sg13g2_o21ai_1 _20669_ (.B1(_03327_),
    .Y(_03328_),
    .A1(_03238_),
    .A2(_03326_));
 sg13g2_nand2_1 _20670_ (.Y(_03329_),
    .A(net172),
    .B(_03328_));
 sg13g2_inv_1 _20671_ (.Y(_03330_),
    .A(_03245_));
 sg13g2_nor3_1 _20672_ (.A(net203),
    .B(_03330_),
    .C(_03310_),
    .Y(_03331_));
 sg13g2_a21oi_1 _20673_ (.A1(net235),
    .A2(net231),
    .Y(_03332_),
    .B1(net228));
 sg13g2_nor3_1 _20674_ (.A(net229),
    .B(_03331_),
    .C(_03332_),
    .Y(_03333_));
 sg13g2_buf_1 _20675_ (.A(_03102_),
    .X(_03334_));
 sg13g2_a21oi_1 _20676_ (.A1(_09897_),
    .A2(_03334_),
    .Y(_03335_),
    .B1(_03030_));
 sg13g2_o21ai_1 _20677_ (.B1(_03335_),
    .Y(_03336_),
    .A1(_03308_),
    .A2(_03333_));
 sg13g2_nor3_1 _20678_ (.A(_03145_),
    .B(_03025_),
    .C(_03202_),
    .Y(_03337_));
 sg13g2_a21o_1 _20679_ (.A2(net205),
    .A1(net244),
    .B1(_03337_),
    .X(_03338_));
 sg13g2_nor2_1 _20680_ (.A(net202),
    .B(_03334_),
    .Y(_03339_));
 sg13g2_a22oi_1 _20681_ (.Y(_03340_),
    .B1(_03339_),
    .B2(_03046_),
    .A2(net219),
    .A1(net203));
 sg13g2_nand2_1 _20682_ (.Y(_03341_),
    .A(net282),
    .B(net246));
 sg13g2_o21ai_1 _20683_ (.B1(_03341_),
    .Y(_03342_),
    .A1(net183),
    .A2(_03340_));
 sg13g2_a22oi_1 _20684_ (.Y(_03343_),
    .B1(_03342_),
    .B2(_09895_),
    .A2(_03338_),
    .A1(_03220_));
 sg13g2_nand3_1 _20685_ (.B(_03336_),
    .C(_03343_),
    .A(_03329_),
    .Y(_03344_));
 sg13g2_mux2_1 _20686_ (.A0(\cpu.dec.imm[6] ),
    .A1(_03344_),
    .S(net98),
    .X(_00766_));
 sg13g2_buf_1 _20687_ (.A(_09014_),
    .X(_03345_));
 sg13g2_a21oi_1 _20688_ (.A1(_09127_),
    .A2(_03203_),
    .Y(_03346_),
    .B1(net228));
 sg13g2_nor2_1 _20689_ (.A(net229),
    .B(net290),
    .Y(_03347_));
 sg13g2_a21oi_1 _20690_ (.A1(_03149_),
    .A2(_03346_),
    .Y(_03348_),
    .B1(_03347_));
 sg13g2_o21ai_1 _20691_ (.B1(net140),
    .Y(_03349_),
    .A1(net232),
    .A2(_09051_));
 sg13g2_a22oi_1 _20692_ (.Y(_03350_),
    .B1(_03349_),
    .B2(_03149_),
    .A2(net235),
    .A1(net172));
 sg13g2_or2_1 _20693_ (.X(_03351_),
    .B(net140),
    .A(net228));
 sg13g2_o21ai_1 _20694_ (.B1(_03351_),
    .Y(_03352_),
    .A1(_09072_),
    .A2(_03350_));
 sg13g2_o21ai_1 _20695_ (.B1(_03352_),
    .Y(_03353_),
    .A1(net183),
    .A2(_03348_));
 sg13g2_o21ai_1 _20696_ (.B1(_03341_),
    .Y(_03354_),
    .A1(_03039_),
    .A2(_09904_));
 sg13g2_nand2_1 _20697_ (.Y(_03355_),
    .A(net234),
    .B(net231));
 sg13g2_a21oi_1 _20698_ (.A1(net233),
    .A2(_03355_),
    .Y(_03356_),
    .B1(net204));
 sg13g2_o21ai_1 _20699_ (.B1(_03356_),
    .Y(_03357_),
    .A1(net228),
    .A2(_03354_));
 sg13g2_o21ai_1 _20700_ (.B1(_03357_),
    .Y(_03358_),
    .A1(_03047_),
    .A2(_03161_));
 sg13g2_a21oi_1 _20701_ (.A1(_09895_),
    .A2(_03358_),
    .Y(_03359_),
    .B1(_03177_));
 sg13g2_buf_1 _20702_ (.A(_03085_),
    .X(_03360_));
 sg13g2_nand2_1 _20703_ (.Y(_03361_),
    .A(_03068_),
    .B(net234));
 sg13g2_o21ai_1 _20704_ (.B1(_03169_),
    .Y(_03362_),
    .A1(_03360_),
    .A2(_03361_));
 sg13g2_nor2_1 _20705_ (.A(_03308_),
    .B(_03362_),
    .Y(_03363_));
 sg13g2_a21oi_1 _20706_ (.A1(_09897_),
    .A2(_03202_),
    .Y(_03364_),
    .B1(_03363_));
 sg13g2_o21ai_1 _20707_ (.B1(_03284_),
    .Y(_03365_),
    .A1(_03337_),
    .A2(_03364_));
 sg13g2_nand3_1 _20708_ (.B(_03359_),
    .C(_03365_),
    .A(_03353_),
    .Y(_03366_));
 sg13g2_nand2_1 _20709_ (.Y(_03367_),
    .A(net97),
    .B(_03366_));
 sg13g2_o21ai_1 _20710_ (.B1(_03367_),
    .Y(_00767_),
    .A1(_11285_),
    .A2(_09892_));
 sg13g2_o21ai_1 _20711_ (.B1(_03194_),
    .Y(_03368_),
    .A1(_09913_),
    .A2(_03206_));
 sg13g2_nor2_1 _20712_ (.A(_03199_),
    .B(_03030_),
    .Y(_03369_));
 sg13g2_nor2_1 _20713_ (.A(_03054_),
    .B(_03360_),
    .Y(_03370_));
 sg13g2_a221oi_1 _20714_ (.B2(_03370_),
    .C1(_03176_),
    .B1(_03369_),
    .A1(_03220_),
    .Y(_03371_),
    .A2(_03368_));
 sg13g2_o21ai_1 _20715_ (.B1(_03208_),
    .Y(_03372_),
    .A1(_09145_),
    .A2(_03204_));
 sg13g2_nand4_1 _20716_ (.B(_03179_),
    .C(_03186_),
    .A(_03173_),
    .Y(_03373_),
    .D(_03372_));
 sg13g2_nand2b_1 _20717_ (.Y(_03374_),
    .B(_03373_),
    .A_N(net140));
 sg13g2_nand3_1 _20718_ (.B(_03371_),
    .C(_03374_),
    .A(_08999_),
    .Y(_03375_));
 sg13g2_o21ai_1 _20719_ (.B1(_03375_),
    .Y(_03376_),
    .A1(\cpu.dec.imm[8] ),
    .A2(net97));
 sg13g2_inv_1 _20720_ (.Y(_00768_),
    .A(_03376_));
 sg13g2_nand2_1 _20721_ (.Y(_03377_),
    .A(_09914_),
    .B(_03188_));
 sg13g2_a21oi_1 _20722_ (.A1(_03194_),
    .A2(_03377_),
    .Y(_03378_),
    .B1(_03132_));
 sg13g2_o21ai_1 _20723_ (.B1(_03208_),
    .Y(_03379_),
    .A1(_09914_),
    .A2(_03204_));
 sg13g2_a221oi_1 _20724_ (.B2(_09097_),
    .C1(_03183_),
    .B1(_03182_),
    .A1(_03038_),
    .Y(_03380_),
    .A2(net205));
 sg13g2_a21oi_1 _20725_ (.A1(_03379_),
    .A2(_03380_),
    .Y(_03381_),
    .B1(_03181_));
 sg13g2_nor3_1 _20726_ (.A(_03176_),
    .B(_03378_),
    .C(_03381_),
    .Y(_03382_));
 sg13g2_nor2_1 _20727_ (.A(\cpu.dec.imm[9] ),
    .B(_09103_),
    .Y(_03383_));
 sg13g2_a21oi_1 _20728_ (.A1(net107),
    .A2(_03382_),
    .Y(_00769_),
    .B1(_03383_));
 sg13g2_buf_1 _20729_ (.A(\cpu.dec.do_inv_mmu ),
    .X(_03384_));
 sg13g2_buf_1 _20730_ (.A(net920),
    .X(_03385_));
 sg13g2_nand2_1 _20731_ (.Y(_03386_),
    .A(_03385_),
    .B(_09897_));
 sg13g2_nor4_1 _20732_ (.A(_09015_),
    .B(_09096_),
    .C(_03125_),
    .D(_03386_),
    .Y(_03387_));
 sg13g2_a21o_1 _20733_ (.A2(net79),
    .A1(_03384_),
    .B1(_03387_),
    .X(_00770_));
 sg13g2_nor3_1 _20734_ (.A(net89),
    .B(_03142_),
    .C(_03263_),
    .Y(_03388_));
 sg13g2_a21o_1 _20735_ (.A2(net79),
    .A1(\cpu.dec.io ),
    .B1(_03388_),
    .X(_00771_));
 sg13g2_nor2_2 _20736_ (.A(_09126_),
    .B(_09173_),
    .Y(_03389_));
 sg13g2_nand2_2 _20737_ (.Y(_03390_),
    .A(_09169_),
    .B(_03389_));
 sg13g2_nor4_1 _20738_ (.A(_09015_),
    .B(_09048_),
    .C(_03155_),
    .D(_03390_),
    .Y(_03391_));
 sg13g2_a21o_1 _20739_ (.A2(net79),
    .A1(\cpu.dec.jmp ),
    .B1(_03391_),
    .X(_00772_));
 sg13g2_o21ai_1 _20740_ (.B1(net186),
    .Y(_03392_),
    .A1(net187),
    .A2(net183));
 sg13g2_nor2_1 _20741_ (.A(net284),
    .B(net291),
    .Y(_03393_));
 sg13g2_a22oi_1 _20742_ (.Y(_03394_),
    .B1(_03393_),
    .B2(net187),
    .A2(_03392_),
    .A1(net185));
 sg13g2_nand2_1 _20743_ (.Y(_03395_),
    .A(_03059_),
    .B(_03135_));
 sg13g2_o21ai_1 _20744_ (.B1(_03395_),
    .Y(_03396_),
    .A1(net207),
    .A2(_03394_));
 sg13g2_mux2_1 _20745_ (.A0(_11521_),
    .A1(_03396_),
    .S(net119),
    .X(_00773_));
 sg13g2_nor3_1 _20746_ (.A(net283),
    .B(_09053_),
    .C(_09094_),
    .Y(_03397_));
 sg13g2_mux2_1 _20747_ (.A0(\cpu.dec.mult ),
    .A1(_03397_),
    .S(net98),
    .X(_00774_));
 sg13g2_nand2_1 _20748_ (.Y(_03398_),
    .A(net208),
    .B(net203));
 sg13g2_nor2_1 _20749_ (.A(net283),
    .B(_03398_),
    .Y(_03399_));
 sg13g2_nor3_1 _20750_ (.A(net208),
    .B(net203),
    .C(_09038_),
    .Y(_03400_));
 sg13g2_nor4_1 _20751_ (.A(net210),
    .B(net206),
    .C(_03399_),
    .D(_03400_),
    .Y(_03401_));
 sg13g2_nor2_1 _20752_ (.A(_08459_),
    .B(_03037_),
    .Y(_03402_));
 sg13g2_nor3_1 _20753_ (.A(_08441_),
    .B(_09884_),
    .C(_03402_),
    .Y(_03403_));
 sg13g2_o21ai_1 _20754_ (.B1(net118),
    .Y(_03404_),
    .A1(_03401_),
    .A2(_03403_));
 sg13g2_o21ai_1 _20755_ (.B1(_03404_),
    .Y(_00775_),
    .A1(net873),
    .A2(net119));
 sg13g2_a21oi_1 _20756_ (.A1(net232),
    .A2(_03393_),
    .Y(_03405_),
    .B1(_03135_));
 sg13g2_nor3_1 _20757_ (.A(_08377_),
    .B(net243),
    .C(_03405_),
    .Y(_03406_));
 sg13g2_nor4_1 _20758_ (.A(net232),
    .B(net282),
    .C(net235),
    .D(_03102_),
    .Y(_03407_));
 sg13g2_nor3_1 _20759_ (.A(net208),
    .B(_03406_),
    .C(_03407_),
    .Y(_03408_));
 sg13g2_nand2_1 _20760_ (.Y(_03409_),
    .A(_03025_),
    .B(net201));
 sg13g2_a22oi_1 _20761_ (.Y(_03410_),
    .B1(_03409_),
    .B2(_03044_),
    .A2(_03310_),
    .A1(net229));
 sg13g2_a21oi_1 _20762_ (.A1(net206),
    .A2(_03284_),
    .Y(_03411_),
    .B1(_03408_));
 sg13g2_o21ai_1 _20763_ (.B1(_09895_),
    .Y(_03412_),
    .A1(net228),
    .A2(net201));
 sg13g2_a21oi_1 _20764_ (.A1(_09169_),
    .A2(_03389_),
    .Y(_03413_),
    .B1(net201));
 sg13g2_nor3_1 _20765_ (.A(net202),
    .B(net293),
    .C(_03390_),
    .Y(_03414_));
 sg13g2_o21ai_1 _20766_ (.B1(_03063_),
    .Y(_03415_),
    .A1(_03413_),
    .A2(_03414_));
 sg13g2_nand2b_1 _20767_ (.Y(_03416_),
    .B(_03415_),
    .A_N(_03412_));
 sg13g2_o21ai_1 _20768_ (.B1(_03416_),
    .Y(_03417_),
    .A1(net203),
    .A2(_03411_));
 sg13g2_a221oi_1 _20769_ (.B2(_03410_),
    .C1(_03417_),
    .B1(_03408_),
    .A1(net243),
    .Y(_03418_),
    .A2(_03369_));
 sg13g2_mux2_1 _20770_ (.A0(\cpu.dec.r_rd[0] ),
    .A1(_03418_),
    .S(net98),
    .X(_00776_));
 sg13g2_nor2_1 _20771_ (.A(_03061_),
    .B(_03182_),
    .Y(_03419_));
 sg13g2_a21o_1 _20772_ (.A2(_03390_),
    .A1(_03063_),
    .B1(_03141_),
    .X(_03420_));
 sg13g2_a22oi_1 _20773_ (.Y(_03421_),
    .B1(_03420_),
    .B2(_09895_),
    .A2(_03419_),
    .A1(_08381_));
 sg13g2_nand4_1 _20774_ (.B(net243),
    .C(net221),
    .A(_09092_),
    .Y(_03422_),
    .D(net246));
 sg13g2_or3_1 _20775_ (.A(_09106_),
    .B(_03125_),
    .C(_03422_),
    .X(_03423_));
 sg13g2_nand3_1 _20776_ (.B(net282),
    .C(net231),
    .A(net202),
    .Y(_03424_));
 sg13g2_nand3_1 _20777_ (.B(net234),
    .C(net246),
    .A(_03048_),
    .Y(_03425_));
 sg13g2_nand3_1 _20778_ (.B(_03424_),
    .C(_03425_),
    .A(_03043_),
    .Y(_03426_));
 sg13g2_o21ai_1 _20779_ (.B1(net202),
    .Y(_03427_),
    .A1(net234),
    .A2(_09162_));
 sg13g2_nand3_1 _20780_ (.B(_03355_),
    .C(_03427_),
    .A(_03139_),
    .Y(_03428_));
 sg13g2_nand2_1 _20781_ (.Y(_03429_),
    .A(_03426_),
    .B(_03428_));
 sg13g2_a21oi_1 _20782_ (.A1(_03132_),
    .A2(_03423_),
    .Y(_03430_),
    .B1(_03429_));
 sg13g2_a21oi_1 _20783_ (.A1(net219),
    .A2(_03369_),
    .Y(_03431_),
    .B1(_03430_));
 sg13g2_o21ai_1 _20784_ (.B1(_03431_),
    .Y(_03432_),
    .A1(_03202_),
    .A2(_03421_));
 sg13g2_mux2_1 _20785_ (.A0(\cpu.dec.r_rd[1] ),
    .A1(_03432_),
    .S(net98),
    .X(_00777_));
 sg13g2_o21ai_1 _20786_ (.B1(_03197_),
    .Y(_03433_),
    .A1(_03261_),
    .A2(_03165_));
 sg13g2_nor2_1 _20787_ (.A(net235),
    .B(net227),
    .Y(_03434_));
 sg13g2_o21ai_1 _20788_ (.B1(_03166_),
    .Y(_03435_),
    .A1(_03150_),
    .A2(_03434_));
 sg13g2_nand2_1 _20789_ (.Y(_03436_),
    .A(_03433_),
    .B(_03435_));
 sg13g2_a22oi_1 _20790_ (.Y(_03437_),
    .B1(_03436_),
    .B2(_03220_),
    .A2(_03369_),
    .A1(net221));
 sg13g2_o21ai_1 _20791_ (.B1(_03437_),
    .Y(_03438_),
    .A1(net227),
    .A2(_03421_));
 sg13g2_mux2_1 _20792_ (.A0(\cpu.dec.r_rd[2] ),
    .A1(_03438_),
    .S(net98),
    .X(_00778_));
 sg13g2_nor3_1 _20793_ (.A(_03048_),
    .B(_03046_),
    .C(_03243_),
    .Y(_03439_));
 sg13g2_a21o_1 _20794_ (.A2(_03166_),
    .A1(_03022_),
    .B1(_03439_),
    .X(_03440_));
 sg13g2_o21ai_1 _20795_ (.B1(_03398_),
    .Y(_03441_),
    .A1(net208),
    .A2(net206));
 sg13g2_a22oi_1 _20796_ (.Y(_03442_),
    .B1(_03441_),
    .B2(net210),
    .A2(_03440_),
    .A1(net195));
 sg13g2_a21oi_1 _20797_ (.A1(net184),
    .A2(_03390_),
    .Y(_03443_),
    .B1(_03197_));
 sg13g2_o21ai_1 _20798_ (.B1(_03069_),
    .Y(_03444_),
    .A1(_08311_),
    .A2(_03443_));
 sg13g2_nand2_1 _20799_ (.Y(_03445_),
    .A(_09895_),
    .B(_03444_));
 sg13g2_nand3_1 _20800_ (.B(_03442_),
    .C(_03445_),
    .A(_08999_),
    .Y(_03446_));
 sg13g2_o21ai_1 _20801_ (.B1(_03446_),
    .Y(_03447_),
    .A1(\cpu.dec.r_rd[3] ),
    .A2(net97));
 sg13g2_inv_1 _20802_ (.Y(_00779_),
    .A(_03447_));
 sg13g2_nand2b_1 _20803_ (.Y(_03448_),
    .B(_09174_),
    .A_N(_09177_));
 sg13g2_inv_1 _20804_ (.Y(_03449_),
    .A(_03448_));
 sg13g2_a221oi_1 _20805_ (.B2(net184),
    .C1(net144),
    .B1(_03449_),
    .A1(net202),
    .Y(_03450_),
    .A2(_03263_));
 sg13g2_nand2_1 _20806_ (.Y(_03451_),
    .A(net206),
    .B(_03027_));
 sg13g2_nand2_1 _20807_ (.Y(_03452_),
    .A(_09035_),
    .B(_03390_));
 sg13g2_nor2_1 _20808_ (.A(_09048_),
    .B(_03155_),
    .Y(_03453_));
 sg13g2_a22oi_1 _20809_ (.Y(_03454_),
    .B1(_03452_),
    .B2(_03453_),
    .A2(_03451_),
    .A1(_08380_));
 sg13g2_o21ai_1 _20810_ (.B1(_03454_),
    .Y(_03455_),
    .A1(_09897_),
    .A2(_03030_));
 sg13g2_nand2_1 _20811_ (.Y(_03456_),
    .A(net201),
    .B(_03395_));
 sg13g2_o21ai_1 _20812_ (.B1(_03456_),
    .Y(_03457_),
    .A1(_03450_),
    .A2(_03455_));
 sg13g2_nand3_1 _20813_ (.B(net203),
    .C(net201),
    .A(net187),
    .Y(_03458_));
 sg13g2_nor2_1 _20814_ (.A(net223),
    .B(net202),
    .Y(_03459_));
 sg13g2_or3_1 _20815_ (.A(net235),
    .B(_03049_),
    .C(_03459_),
    .X(_03460_));
 sg13g2_nand4_1 _20816_ (.B(net186),
    .C(_03458_),
    .A(net185),
    .Y(_03461_),
    .D(_03460_));
 sg13g2_nand3_1 _20817_ (.B(_03457_),
    .C(_03461_),
    .A(_08999_),
    .Y(_03462_));
 sg13g2_o21ai_1 _20818_ (.B1(_03462_),
    .Y(_03463_),
    .A1(_10586_),
    .A2(net97));
 sg13g2_inv_1 _20819_ (.Y(_00780_),
    .A(_03463_));
 sg13g2_o21ai_1 _20820_ (.B1(_09048_),
    .Y(_03464_),
    .A1(net186),
    .A2(net231));
 sg13g2_o21ai_1 _20821_ (.B1(net231),
    .Y(_03465_),
    .A1(net202),
    .A2(_03452_));
 sg13g2_nand3_1 _20822_ (.B(_03152_),
    .C(_03465_),
    .A(_03040_),
    .Y(_03466_));
 sg13g2_a21oi_1 _20823_ (.A1(net204),
    .A2(_03448_),
    .Y(_03467_),
    .B1(net282));
 sg13g2_nor2_1 _20824_ (.A(net232),
    .B(_03467_),
    .Y(_03468_));
 sg13g2_nor3_1 _20825_ (.A(_03235_),
    .B(_03393_),
    .C(_03468_),
    .Y(_03469_));
 sg13g2_nor2_1 _20826_ (.A(net144),
    .B(_03469_),
    .Y(_03470_));
 sg13g2_o21ai_1 _20827_ (.B1(_03145_),
    .Y(_03471_),
    .A1(net204),
    .A2(_03104_));
 sg13g2_nor2_1 _20828_ (.A(net223),
    .B(_03202_),
    .Y(_03472_));
 sg13g2_nand3_1 _20829_ (.B(_03471_),
    .C(_03472_),
    .A(net229),
    .Y(_03473_));
 sg13g2_a21oi_1 _20830_ (.A1(_03152_),
    .A2(_03179_),
    .Y(_03474_),
    .B1(_03029_));
 sg13g2_a22oi_1 _20831_ (.Y(_03475_),
    .B1(_03474_),
    .B2(net209),
    .A2(_03472_),
    .A1(_09046_));
 sg13g2_a21oi_1 _20832_ (.A1(_03473_),
    .A2(_03475_),
    .Y(_03476_),
    .B1(net208));
 sg13g2_a221oi_1 _20833_ (.B2(net231),
    .C1(_03476_),
    .B1(_03470_),
    .A1(net185),
    .Y(_03477_),
    .A2(_03466_));
 sg13g2_a21oi_1 _20834_ (.A1(_03284_),
    .A2(_03464_),
    .Y(_03478_),
    .B1(_03477_));
 sg13g2_nand2_1 _20835_ (.Y(_03479_),
    .A(net97),
    .B(_03478_));
 sg13g2_o21ai_1 _20836_ (.B1(_03479_),
    .Y(_00781_),
    .A1(net747),
    .A2(net106));
 sg13g2_nor2b_1 _20837_ (.A(_03470_),
    .B_N(_03454_),
    .Y(_03480_));
 sg13g2_o21ai_1 _20838_ (.B1(_03025_),
    .Y(_03481_),
    .A1(net234),
    .A2(net227));
 sg13g2_nor2_1 _20839_ (.A(net233),
    .B(net227),
    .Y(_03482_));
 sg13g2_a22oi_1 _20840_ (.Y(_03483_),
    .B1(_03482_),
    .B2(_03040_),
    .A2(_03481_),
    .A1(net236));
 sg13g2_inv_1 _20841_ (.Y(_03484_),
    .A(_03483_));
 sg13g2_o21ai_1 _20842_ (.B1(_03152_),
    .Y(_03485_),
    .A1(net208),
    .A2(_03179_));
 sg13g2_a22oi_1 _20843_ (.Y(_03486_),
    .B1(_03485_),
    .B2(_03040_),
    .A2(_03484_),
    .A1(_03052_));
 sg13g2_o21ai_1 _20844_ (.B1(_03486_),
    .Y(_03487_),
    .A1(net227),
    .A2(_03480_));
 sg13g2_nand2_1 _20845_ (.Y(_03488_),
    .A(net97),
    .B(_03487_));
 sg13g2_o21ai_1 _20846_ (.B1(_03488_),
    .Y(_00782_),
    .A1(net737),
    .A2(net106));
 sg13g2_nand2_1 _20847_ (.Y(_03489_),
    .A(net184),
    .B(_03284_));
 sg13g2_nand2_1 _20848_ (.Y(_03490_),
    .A(net233),
    .B(net204));
 sg13g2_a21oi_1 _20849_ (.A1(net288),
    .A2(_03452_),
    .Y(_03491_),
    .B1(_03490_));
 sg13g2_o21ai_1 _20850_ (.B1(net186),
    .Y(_03492_),
    .A1(net228),
    .A2(net183));
 sg13g2_o21ai_1 _20851_ (.B1(net187),
    .Y(_03493_),
    .A1(_03491_),
    .A2(_03492_));
 sg13g2_a21o_1 _20852_ (.A2(_03451_),
    .A1(net236),
    .B1(net208),
    .X(_03494_));
 sg13g2_a21o_1 _20853_ (.A2(_03494_),
    .A1(_03493_),
    .B1(_03450_),
    .X(_03495_));
 sg13g2_nand3_1 _20854_ (.B(_03489_),
    .C(_03495_),
    .A(_09014_),
    .Y(_03496_));
 sg13g2_o21ai_1 _20855_ (.B1(_03496_),
    .Y(_00783_),
    .A1(net736),
    .A2(net106));
 sg13g2_nand3_1 _20856_ (.B(net205),
    .C(net201),
    .A(net187),
    .Y(_03497_));
 sg13g2_o21ai_1 _20857_ (.B1(_03497_),
    .Y(_03498_),
    .A1(_09145_),
    .A2(net205));
 sg13g2_o21ai_1 _20858_ (.B1(_09163_),
    .Y(_03499_),
    .A1(_09173_),
    .A2(net201));
 sg13g2_nor2_1 _20859_ (.A(_09177_),
    .B(_03169_),
    .Y(_03500_));
 sg13g2_a21o_1 _20860_ (.A2(_09177_),
    .A1(_08440_),
    .B1(_03235_),
    .X(_03501_));
 sg13g2_buf_1 _20861_ (.A(_03501_),
    .X(_03502_));
 sg13g2_a221oi_1 _20862_ (.B2(_09145_),
    .C1(net144),
    .B1(_03502_),
    .A1(_03499_),
    .Y(_03503_),
    .A2(_03500_));
 sg13g2_a221oi_1 _20863_ (.B2(net185),
    .C1(_03503_),
    .B1(_03498_),
    .A1(net210),
    .Y(_03504_),
    .A2(net243));
 sg13g2_nand2_1 _20864_ (.Y(_03505_),
    .A(net97),
    .B(_03504_));
 sg13g2_o21ai_1 _20865_ (.B1(_03505_),
    .Y(_00784_),
    .A1(net671),
    .A2(net106));
 sg13g2_nand3_1 _20866_ (.B(net205),
    .C(_03202_),
    .A(net187),
    .Y(_03506_));
 sg13g2_o21ai_1 _20867_ (.B1(_03506_),
    .Y(_03507_),
    .A1(net219),
    .A2(net205));
 sg13g2_o21ai_1 _20868_ (.B1(_09173_),
    .Y(_03508_),
    .A1(net220),
    .A2(_09172_));
 sg13g2_nand2_1 _20869_ (.Y(_03509_),
    .A(_08440_),
    .B(_03508_));
 sg13g2_nor3_1 _20870_ (.A(_09177_),
    .B(_03389_),
    .C(_03509_),
    .Y(_03510_));
 sg13g2_nand2_1 _20871_ (.Y(_03511_),
    .A(_09174_),
    .B(_03202_));
 sg13g2_a221oi_1 _20872_ (.B2(_03511_),
    .C1(net144),
    .B1(_03510_),
    .A1(net219),
    .Y(_03512_),
    .A2(_03502_));
 sg13g2_a221oi_1 _20873_ (.B2(net185),
    .C1(_03512_),
    .B1(_03507_),
    .A1(net210),
    .Y(_03513_),
    .A2(_09172_));
 sg13g2_nand2_1 _20874_ (.Y(_03514_),
    .A(_03345_),
    .B(_03513_));
 sg13g2_o21ai_1 _20875_ (.B1(_03514_),
    .Y(_00785_),
    .A1(net754),
    .A2(net106));
 sg13g2_a21oi_1 _20876_ (.A1(net195),
    .A2(_03502_),
    .Y(_03515_),
    .B1(net210));
 sg13g2_a21oi_1 _20877_ (.A1(_09174_),
    .A2(net227),
    .Y(_03516_),
    .B1(net144));
 sg13g2_or3_1 _20878_ (.A(net236),
    .B(_03027_),
    .C(net227),
    .X(_03517_));
 sg13g2_o21ai_1 _20879_ (.B1(_03517_),
    .Y(_03518_),
    .A1(net220),
    .A2(net205));
 sg13g2_a22oi_1 _20880_ (.Y(_03519_),
    .B1(_03518_),
    .B2(net185),
    .A2(_03516_),
    .A1(_03510_));
 sg13g2_o21ai_1 _20881_ (.B1(_03519_),
    .Y(_03520_),
    .A1(net220),
    .A2(_03515_));
 sg13g2_nand2_1 _20882_ (.Y(_03521_),
    .A(_03345_),
    .B(_03520_));
 sg13g2_o21ai_1 _20883_ (.B1(_03521_),
    .Y(_00786_),
    .A1(net666),
    .A2(net105));
 sg13g2_nor2_1 _20884_ (.A(net207),
    .B(net184),
    .Y(_03522_));
 sg13g2_o21ai_1 _20885_ (.B1(net222),
    .Y(_03523_),
    .A1(_08440_),
    .A2(_03522_));
 sg13g2_o21ai_1 _20886_ (.B1(_03523_),
    .Y(_03524_),
    .A1(net288),
    .A2(_03027_));
 sg13g2_inv_1 _20887_ (.Y(_03525_),
    .A(_03509_));
 sg13g2_nor3_1 _20888_ (.A(_09175_),
    .B(_03502_),
    .C(_03525_),
    .Y(_03526_));
 sg13g2_a21oi_1 _20889_ (.A1(_09895_),
    .A2(_03524_),
    .Y(_03527_),
    .B1(_03526_));
 sg13g2_mux2_1 _20890_ (.A0(net611),
    .A1(_03527_),
    .S(_03233_),
    .X(_00787_));
 sg13g2_mux2_1 _20891_ (.A0(_10322_),
    .A1(_09164_),
    .S(net98),
    .X(_00788_));
 sg13g2_nand3_1 _20892_ (.B(_09178_),
    .C(_03389_),
    .A(net118),
    .Y(_03528_));
 sg13g2_o21ai_1 _20893_ (.B1(_03528_),
    .Y(_00789_),
    .A1(_10467_),
    .A2(net105));
 sg13g2_inv_1 _20894_ (.Y(_03529_),
    .A(\cpu.dec.r_set_cc ));
 sg13g2_nand3_1 _20895_ (.B(_09108_),
    .C(_09105_),
    .A(net118),
    .Y(_03530_));
 sg13g2_o21ai_1 _20896_ (.B1(_03530_),
    .Y(_00790_),
    .A1(_03529_),
    .A2(net105));
 sg13g2_inv_1 _20897_ (.Y(_03531_),
    .A(\cpu.dec.r_store ));
 sg13g2_nor3_1 _20898_ (.A(net206),
    .B(net144),
    .C(_03134_),
    .Y(_03532_));
 sg13g2_o21ai_1 _20899_ (.B1(net207),
    .Y(_03533_),
    .A1(_03064_),
    .A2(_03532_));
 sg13g2_o21ai_1 _20900_ (.B1(_03533_),
    .Y(_03534_),
    .A1(_03025_),
    .A2(_03142_));
 sg13g2_nand2_1 _20901_ (.Y(_03535_),
    .A(net97),
    .B(_03534_));
 sg13g2_o21ai_1 _20902_ (.B1(_03535_),
    .Y(_00791_),
    .A1(_03531_),
    .A2(net105));
 sg13g2_nor3_1 _20903_ (.A(net89),
    .B(_03127_),
    .C(_03422_),
    .Y(_03536_));
 sg13g2_a21o_1 _20904_ (.A2(_09016_),
    .A1(\cpu.dec.r_swapsp ),
    .B1(_03536_),
    .X(_00792_));
 sg13g2_nor4_1 _20905_ (.A(_09015_),
    .B(_09882_),
    .C(_03127_),
    .D(_03129_),
    .Y(_03537_));
 sg13g2_a21o_1 _20906_ (.A2(_09016_),
    .A1(\cpu.dec.r_sys_call ),
    .B1(_03537_),
    .X(_00793_));
 sg13g2_nor2_1 _20907_ (.A(net283),
    .B(_09145_),
    .Y(_03538_));
 sg13g2_a21oi_1 _20908_ (.A1(net283),
    .A2(_09169_),
    .Y(_03539_),
    .B1(_03538_));
 sg13g2_o21ai_1 _20909_ (.B1(_09895_),
    .Y(_03540_),
    .A1(_03069_),
    .A2(_03539_));
 sg13g2_xnor2_1 _20910_ (.Y(_03541_),
    .A(net220),
    .B(_09163_));
 sg13g2_nand2_1 _20911_ (.Y(_03542_),
    .A(_08476_),
    .B(_09035_));
 sg13g2_o21ai_1 _20912_ (.B1(_03542_),
    .Y(_03543_),
    .A1(net920),
    .A2(_09035_));
 sg13g2_nand2_1 _20913_ (.Y(_03544_),
    .A(_03170_),
    .B(_03543_));
 sg13g2_o21ai_1 _20914_ (.B1(net233),
    .Y(_03545_),
    .A1(_03541_),
    .A2(_03544_));
 sg13g2_a21oi_1 _20915_ (.A1(net183),
    .A2(_03452_),
    .Y(_03546_),
    .B1(net229));
 sg13g2_nand2_1 _20916_ (.Y(_03547_),
    .A(net186),
    .B(_03545_));
 sg13g2_o21ai_1 _20917_ (.B1(_03547_),
    .Y(_03548_),
    .A1(net288),
    .A2(_03546_));
 sg13g2_nand2b_1 _20918_ (.Y(_03549_),
    .B(_03122_),
    .A_N(_03102_));
 sg13g2_xnor2_1 _20919_ (.Y(_03550_),
    .A(_03085_),
    .B(_03549_));
 sg13g2_nor2_1 _20920_ (.A(net721),
    .B(_03550_),
    .Y(_03551_));
 sg13g2_a22oi_1 _20921_ (.Y(_03552_),
    .B1(_03548_),
    .B2(_03551_),
    .A2(_03545_),
    .A1(net184));
 sg13g2_nand2_1 _20922_ (.Y(_03553_),
    .A(_08310_),
    .B(_09071_));
 sg13g2_o21ai_1 _20923_ (.B1(_03553_),
    .Y(_03554_),
    .A1(net336),
    .A2(_09169_));
 sg13g2_a22oi_1 _20924_ (.Y(_03555_),
    .B1(_03554_),
    .B2(_03037_),
    .A2(_03402_),
    .A1(_09145_));
 sg13g2_nand3_1 _20925_ (.B(_03188_),
    .C(_03551_),
    .A(_08311_),
    .Y(_03556_));
 sg13g2_o21ai_1 _20926_ (.B1(_03556_),
    .Y(_03557_),
    .A1(_09048_),
    .A2(_03555_));
 sg13g2_nand4_1 _20927_ (.B(net227),
    .C(net201),
    .A(_09093_),
    .Y(_03558_),
    .D(_03202_));
 sg13g2_nor4_1 _20928_ (.A(_03385_),
    .B(_10969_),
    .C(net292),
    .D(_03041_),
    .Y(_03559_));
 sg13g2_o21ai_1 _20929_ (.B1(_09172_),
    .Y(_03560_),
    .A1(net920),
    .A2(_09144_));
 sg13g2_nand3_1 _20930_ (.B(net221),
    .C(_03560_),
    .A(_09091_),
    .Y(_03561_));
 sg13g2_nand2_1 _20931_ (.Y(_03562_),
    .A(_09072_),
    .B(_03561_));
 sg13g2_nand3_1 _20932_ (.B(_03037_),
    .C(_03562_),
    .A(_08310_),
    .Y(_03563_));
 sg13g2_nand3_1 _20933_ (.B(_08459_),
    .C(_03563_),
    .A(net233),
    .Y(_03564_));
 sg13g2_o21ai_1 _20934_ (.B1(_03564_),
    .Y(_03565_),
    .A1(net184),
    .A2(_03559_));
 sg13g2_nor2_1 _20935_ (.A(net283),
    .B(_03386_),
    .Y(_03566_));
 sg13g2_a21oi_1 _20936_ (.A1(net289),
    .A2(_09904_),
    .Y(_03567_),
    .B1(net290));
 sg13g2_a21oi_1 _20937_ (.A1(_03422_),
    .A2(_03567_),
    .Y(_03568_),
    .B1(_03123_));
 sg13g2_a221oi_1 _20938_ (.B2(_03568_),
    .C1(net144),
    .B1(_03566_),
    .A1(_03556_),
    .Y(_03569_),
    .A2(_03565_));
 sg13g2_a221oi_1 _20939_ (.B2(_03031_),
    .C1(_03569_),
    .B1(_03558_),
    .A1(net172),
    .Y(_03570_),
    .A2(_03557_));
 sg13g2_o21ai_1 _20940_ (.B1(_03570_),
    .Y(_03571_),
    .A1(_03540_),
    .A2(_03552_));
 sg13g2_mux2_1 _20941_ (.A0(_09212_),
    .A1(_03571_),
    .S(net98),
    .X(_00794_));
 sg13g2_buf_1 _20942_ (.A(net1126),
    .X(_03572_));
 sg13g2_buf_1 _20943_ (.A(_03572_),
    .X(_03573_));
 sg13g2_nand2b_1 _20944_ (.Y(_03574_),
    .B(net1019),
    .A_N(net1018));
 sg13g2_buf_1 _20945_ (.A(_03574_),
    .X(_03575_));
 sg13g2_inv_1 _20946_ (.Y(_03576_),
    .A(_10227_));
 sg13g2_nand3_1 _20947_ (.B(_03576_),
    .C(net1112),
    .A(_10225_),
    .Y(_03577_));
 sg13g2_buf_1 _20948_ (.A(_03577_),
    .X(_03578_));
 sg13g2_nor2_1 _20949_ (.A(_03575_),
    .B(_03578_),
    .Y(_03579_));
 sg13g2_buf_1 _20950_ (.A(_03579_),
    .X(_03580_));
 sg13g2_buf_1 _20951_ (.A(net597),
    .X(_03581_));
 sg13g2_mux2_1 _20952_ (.A0(\cpu.ex.r_10[0] ),
    .A1(net833),
    .S(net523),
    .X(_00799_));
 sg13g2_mux2_1 _20953_ (.A0(\cpu.ex.r_10[10] ),
    .A1(net836),
    .S(net523),
    .X(_00800_));
 sg13g2_mux2_1 _20954_ (.A0(\cpu.ex.r_10[11] ),
    .A1(net835),
    .S(_03581_),
    .X(_00801_));
 sg13g2_buf_1 _20955_ (.A(net620),
    .X(_03582_));
 sg13g2_buf_1 _20956_ (.A(net522),
    .X(_03583_));
 sg13g2_mux2_1 _20957_ (.A0(\cpu.ex.r_10[12] ),
    .A1(net459),
    .S(net523),
    .X(_00802_));
 sg13g2_buf_1 _20958_ (.A(net614),
    .X(_03584_));
 sg13g2_buf_1 _20959_ (.A(net521),
    .X(_03585_));
 sg13g2_mux2_1 _20960_ (.A0(\cpu.ex.r_10[13] ),
    .A1(net458),
    .S(net523),
    .X(_00803_));
 sg13g2_buf_1 _20961_ (.A(_11895_),
    .X(_03586_));
 sg13g2_nand2_1 _20962_ (.Y(_03587_),
    .A(net520),
    .B(net597));
 sg13g2_o21ai_1 _20963_ (.B1(_03587_),
    .Y(_00804_),
    .A1(_11455_),
    .A2(net523));
 sg13g2_buf_1 _20964_ (.A(_11905_),
    .X(_03588_));
 sg13g2_mux2_1 _20965_ (.A0(\cpu.ex.r_10[15] ),
    .A1(net720),
    .S(net523),
    .X(_00805_));
 sg13g2_buf_1 _20966_ (.A(net538),
    .X(_03589_));
 sg13g2_mux2_1 _20967_ (.A0(\cpu.ex.r_10[1] ),
    .A1(net457),
    .S(_03581_),
    .X(_00806_));
 sg13g2_buf_1 _20968_ (.A(_09286_),
    .X(_03590_));
 sg13g2_buf_1 _20969_ (.A(net596),
    .X(_03591_));
 sg13g2_mux2_1 _20970_ (.A0(\cpu.ex.r_10[2] ),
    .A1(net519),
    .S(net597),
    .X(_00807_));
 sg13g2_buf_1 _20971_ (.A(net632),
    .X(_03592_));
 sg13g2_mux2_1 _20972_ (.A0(\cpu.ex.r_10[3] ),
    .A1(net518),
    .S(net597),
    .X(_00808_));
 sg13g2_buf_2 _20973_ (.A(net656),
    .X(_03593_));
 sg13g2_buf_1 _20974_ (.A(net595),
    .X(_03594_));
 sg13g2_mux2_1 _20975_ (.A0(\cpu.ex.r_10[4] ),
    .A1(net517),
    .S(net597),
    .X(_00809_));
 sg13g2_mux2_1 _20976_ (.A0(\cpu.ex.r_10[5] ),
    .A1(_02992_),
    .S(net597),
    .X(_00810_));
 sg13g2_nand2_1 _20977_ (.Y(_03595_),
    .A(net847),
    .B(net597));
 sg13g2_o21ai_1 _20978_ (.B1(_03595_),
    .Y(_00811_),
    .A1(_10792_),
    .A2(net523));
 sg13g2_mux2_1 _20979_ (.A0(\cpu.ex.r_10[7] ),
    .A1(net725),
    .S(_03580_),
    .X(_00812_));
 sg13g2_mux2_1 _20980_ (.A0(\cpu.ex.r_10[8] ),
    .A1(_03018_),
    .S(_03580_),
    .X(_00813_));
 sg13g2_nand2_1 _20981_ (.Y(_03596_),
    .A(net969),
    .B(net597));
 sg13g2_o21ai_1 _20982_ (.B1(_03596_),
    .Y(_00814_),
    .A1(_11091_),
    .A2(net523));
 sg13g2_nor2_1 _20983_ (.A(_10233_),
    .B(_03578_),
    .Y(_03597_));
 sg13g2_buf_4 _20984_ (.X(_03598_),
    .A(_03597_));
 sg13g2_buf_1 _20985_ (.A(_03598_),
    .X(_03599_));
 sg13g2_mux2_1 _20986_ (.A0(\cpu.ex.r_11[0] ),
    .A1(net833),
    .S(net516),
    .X(_00815_));
 sg13g2_mux2_1 _20987_ (.A0(\cpu.ex.r_11[10] ),
    .A1(_03020_),
    .S(net516),
    .X(_00816_));
 sg13g2_mux2_1 _20988_ (.A0(\cpu.ex.r_11[11] ),
    .A1(net835),
    .S(net516),
    .X(_00817_));
 sg13g2_mux2_1 _20989_ (.A0(\cpu.ex.r_11[12] ),
    .A1(net459),
    .S(net516),
    .X(_00818_));
 sg13g2_mux2_1 _20990_ (.A0(\cpu.ex.r_11[13] ),
    .A1(net458),
    .S(net516),
    .X(_00819_));
 sg13g2_nand2_1 _20991_ (.Y(_03600_),
    .A(net520),
    .B(_03598_));
 sg13g2_o21ai_1 _20992_ (.B1(_03600_),
    .Y(_00820_),
    .A1(_11452_),
    .A2(net516));
 sg13g2_mux2_1 _20993_ (.A0(\cpu.ex.r_11[15] ),
    .A1(net720),
    .S(net516),
    .X(_00821_));
 sg13g2_mux2_1 _20994_ (.A0(\cpu.ex.r_11[1] ),
    .A1(net457),
    .S(net516),
    .X(_00822_));
 sg13g2_mux2_1 _20995_ (.A0(\cpu.ex.r_11[2] ),
    .A1(net519),
    .S(_03599_),
    .X(_00823_));
 sg13g2_mux2_1 _20996_ (.A0(\cpu.ex.r_11[3] ),
    .A1(_03592_),
    .S(_03599_),
    .X(_00824_));
 sg13g2_mux2_1 _20997_ (.A0(\cpu.ex.r_11[4] ),
    .A1(net517),
    .S(_03598_),
    .X(_00825_));
 sg13g2_mux2_1 _20998_ (.A0(\cpu.ex.r_11[5] ),
    .A1(net524),
    .S(_03598_),
    .X(_00826_));
 sg13g2_mux2_1 _20999_ (.A0(\cpu.ex.r_11[6] ),
    .A1(net723),
    .S(_03598_),
    .X(_00827_));
 sg13g2_mux2_1 _21000_ (.A0(\cpu.ex.r_11[7] ),
    .A1(net725),
    .S(_03598_),
    .X(_00828_));
 sg13g2_mux2_1 _21001_ (.A0(\cpu.ex.r_11[8] ),
    .A1(net722),
    .S(_03598_),
    .X(_00829_));
 sg13g2_mux2_1 _21002_ (.A0(\cpu.ex.r_11[9] ),
    .A1(net837),
    .S(_03598_),
    .X(_00830_));
 sg13g2_nand3_1 _21003_ (.B(net1110),
    .C(net1112),
    .A(net1111),
    .Y(_03601_));
 sg13g2_buf_1 _21004_ (.A(_03601_),
    .X(_03602_));
 sg13g2_nor3_1 _21005_ (.A(_10230_),
    .B(_10232_),
    .C(_03602_),
    .Y(_03603_));
 sg13g2_buf_2 _21006_ (.A(_03603_),
    .X(_03604_));
 sg13g2_buf_1 _21007_ (.A(_03604_),
    .X(_03605_));
 sg13g2_mux2_1 _21008_ (.A0(\cpu.ex.r_12[0] ),
    .A1(net833),
    .S(net594),
    .X(_00831_));
 sg13g2_mux2_1 _21009_ (.A0(\cpu.ex.r_12[10] ),
    .A1(net836),
    .S(net594),
    .X(_00832_));
 sg13g2_mux2_1 _21010_ (.A0(\cpu.ex.r_12[11] ),
    .A1(net835),
    .S(_03605_),
    .X(_00833_));
 sg13g2_mux2_1 _21011_ (.A0(\cpu.ex.r_12[12] ),
    .A1(net459),
    .S(net594),
    .X(_00834_));
 sg13g2_mux2_1 _21012_ (.A0(\cpu.ex.r_12[13] ),
    .A1(net458),
    .S(net594),
    .X(_00835_));
 sg13g2_buf_1 _21013_ (.A(net520),
    .X(_03606_));
 sg13g2_mux2_1 _21014_ (.A0(\cpu.ex.r_12[14] ),
    .A1(net456),
    .S(net594),
    .X(_00836_));
 sg13g2_inv_1 _21015_ (.Y(_03607_),
    .A(\cpu.ex.r_12[15] ));
 sg13g2_nand2_1 _21016_ (.Y(_03608_),
    .A(net860),
    .B(_03604_));
 sg13g2_o21ai_1 _21017_ (.B1(_03608_),
    .Y(_00837_),
    .A1(_03607_),
    .A2(net594));
 sg13g2_mux2_1 _21018_ (.A0(\cpu.ex.r_12[1] ),
    .A1(net457),
    .S(_03605_),
    .X(_00838_));
 sg13g2_mux2_1 _21019_ (.A0(\cpu.ex.r_12[2] ),
    .A1(net519),
    .S(net594),
    .X(_00839_));
 sg13g2_mux2_1 _21020_ (.A0(\cpu.ex.r_12[3] ),
    .A1(net518),
    .S(net594),
    .X(_00840_));
 sg13g2_mux2_1 _21021_ (.A0(\cpu.ex.r_12[4] ),
    .A1(net517),
    .S(_03604_),
    .X(_00841_));
 sg13g2_mux2_1 _21022_ (.A0(\cpu.ex.r_12[5] ),
    .A1(_02992_),
    .S(_03604_),
    .X(_00842_));
 sg13g2_mux2_1 _21023_ (.A0(\cpu.ex.r_12[6] ),
    .A1(net723),
    .S(_03604_),
    .X(_00843_));
 sg13g2_mux2_1 _21024_ (.A0(\cpu.ex.r_12[7] ),
    .A1(_02997_),
    .S(_03604_),
    .X(_00844_));
 sg13g2_mux2_1 _21025_ (.A0(\cpu.ex.r_12[8] ),
    .A1(net722),
    .S(_03604_),
    .X(_00845_));
 sg13g2_mux2_1 _21026_ (.A0(\cpu.ex.r_12[9] ),
    .A1(net837),
    .S(_03604_),
    .X(_00846_));
 sg13g2_inv_1 _21027_ (.Y(_03609_),
    .A(net1019));
 sg13g2_nand2_1 _21028_ (.Y(_03610_),
    .A(_03609_),
    .B(net1018));
 sg13g2_nor2_1 _21029_ (.A(_03602_),
    .B(_03610_),
    .Y(_03611_));
 sg13g2_buf_2 _21030_ (.A(_03611_),
    .X(_03612_));
 sg13g2_buf_1 _21031_ (.A(_03612_),
    .X(_03613_));
 sg13g2_mux2_1 _21032_ (.A0(\cpu.ex.r_13[0] ),
    .A1(net833),
    .S(net515),
    .X(_00847_));
 sg13g2_mux2_1 _21033_ (.A0(\cpu.ex.r_13[10] ),
    .A1(_03020_),
    .S(net515),
    .X(_00848_));
 sg13g2_mux2_1 _21034_ (.A0(\cpu.ex.r_13[11] ),
    .A1(_03021_),
    .S(_03613_),
    .X(_00849_));
 sg13g2_mux2_1 _21035_ (.A0(\cpu.ex.r_13[12] ),
    .A1(net459),
    .S(net515),
    .X(_00850_));
 sg13g2_mux2_1 _21036_ (.A0(\cpu.ex.r_13[13] ),
    .A1(net458),
    .S(net515),
    .X(_00851_));
 sg13g2_mux2_1 _21037_ (.A0(\cpu.ex.r_13[14] ),
    .A1(net456),
    .S(net515),
    .X(_00852_));
 sg13g2_mux2_1 _21038_ (.A0(\cpu.ex.r_13[15] ),
    .A1(net720),
    .S(net515),
    .X(_00853_));
 sg13g2_mux2_1 _21039_ (.A0(\cpu.ex.r_13[1] ),
    .A1(net457),
    .S(net515),
    .X(_00854_));
 sg13g2_mux2_1 _21040_ (.A0(\cpu.ex.r_13[2] ),
    .A1(net519),
    .S(net515),
    .X(_00855_));
 sg13g2_mux2_1 _21041_ (.A0(\cpu.ex.r_13[3] ),
    .A1(net518),
    .S(_03613_),
    .X(_00856_));
 sg13g2_mux2_1 _21042_ (.A0(\cpu.ex.r_13[4] ),
    .A1(net517),
    .S(_03612_),
    .X(_00857_));
 sg13g2_mux2_1 _21043_ (.A0(\cpu.ex.r_13[5] ),
    .A1(net524),
    .S(_03612_),
    .X(_00858_));
 sg13g2_mux2_1 _21044_ (.A0(\cpu.ex.r_13[6] ),
    .A1(net723),
    .S(_03612_),
    .X(_00859_));
 sg13g2_mux2_1 _21045_ (.A0(\cpu.ex.r_13[7] ),
    .A1(_02997_),
    .S(_03612_),
    .X(_00860_));
 sg13g2_mux2_1 _21046_ (.A0(\cpu.ex.r_13[8] ),
    .A1(net722),
    .S(_03612_),
    .X(_00861_));
 sg13g2_mux2_1 _21047_ (.A0(\cpu.ex.r_13[9] ),
    .A1(net837),
    .S(_03612_),
    .X(_00862_));
 sg13g2_nor2_1 _21048_ (.A(_03575_),
    .B(_03602_),
    .Y(_03614_));
 sg13g2_buf_2 _21049_ (.A(_03614_),
    .X(_03615_));
 sg13g2_buf_1 _21050_ (.A(_03615_),
    .X(_03616_));
 sg13g2_mux2_1 _21051_ (.A0(\cpu.ex.r_14[0] ),
    .A1(net833),
    .S(net514),
    .X(_00863_));
 sg13g2_mux2_1 _21052_ (.A0(\cpu.ex.r_14[10] ),
    .A1(net836),
    .S(net514),
    .X(_00864_));
 sg13g2_mux2_1 _21053_ (.A0(\cpu.ex.r_14[11] ),
    .A1(net835),
    .S(_03616_),
    .X(_00865_));
 sg13g2_mux2_1 _21054_ (.A0(\cpu.ex.r_14[12] ),
    .A1(net459),
    .S(net514),
    .X(_00866_));
 sg13g2_mux2_1 _21055_ (.A0(\cpu.ex.r_14[13] ),
    .A1(net458),
    .S(net514),
    .X(_00867_));
 sg13g2_mux2_1 _21056_ (.A0(\cpu.ex.r_14[14] ),
    .A1(net456),
    .S(net514),
    .X(_00868_));
 sg13g2_mux2_1 _21057_ (.A0(\cpu.ex.r_14[15] ),
    .A1(net720),
    .S(net514),
    .X(_00869_));
 sg13g2_mux2_1 _21058_ (.A0(\cpu.ex.r_14[1] ),
    .A1(net457),
    .S(net514),
    .X(_00870_));
 sg13g2_mux2_1 _21059_ (.A0(\cpu.ex.r_14[2] ),
    .A1(_03591_),
    .S(_03616_),
    .X(_00871_));
 sg13g2_mux2_1 _21060_ (.A0(\cpu.ex.r_14[3] ),
    .A1(net518),
    .S(net514),
    .X(_00872_));
 sg13g2_mux2_1 _21061_ (.A0(\cpu.ex.r_14[4] ),
    .A1(_03594_),
    .S(_03615_),
    .X(_00873_));
 sg13g2_buf_1 _21062_ (.A(net651),
    .X(_03617_));
 sg13g2_mux2_1 _21063_ (.A0(\cpu.ex.r_14[5] ),
    .A1(net593),
    .S(_03615_),
    .X(_00874_));
 sg13g2_mux2_1 _21064_ (.A0(\cpu.ex.r_14[6] ),
    .A1(_03016_),
    .S(_03615_),
    .X(_00875_));
 sg13g2_buf_1 _21065_ (.A(net841),
    .X(_03618_));
 sg13g2_mux2_1 _21066_ (.A0(\cpu.ex.r_14[7] ),
    .A1(net719),
    .S(_03615_),
    .X(_00876_));
 sg13g2_mux2_1 _21067_ (.A0(\cpu.ex.r_14[8] ),
    .A1(net722),
    .S(_03615_),
    .X(_00877_));
 sg13g2_mux2_1 _21068_ (.A0(\cpu.ex.r_14[9] ),
    .A1(_03019_),
    .S(_03615_),
    .X(_00878_));
 sg13g2_nor2_1 _21069_ (.A(_10233_),
    .B(_03602_),
    .Y(_03619_));
 sg13g2_buf_2 _21070_ (.A(_03619_),
    .X(_03620_));
 sg13g2_buf_1 _21071_ (.A(_03620_),
    .X(_03621_));
 sg13g2_mux2_1 _21072_ (.A0(\cpu.ex.r_15[0] ),
    .A1(_03573_),
    .S(_03621_),
    .X(_00879_));
 sg13g2_mux2_1 _21073_ (.A0(\cpu.ex.r_15[10] ),
    .A1(net836),
    .S(net592),
    .X(_00880_));
 sg13g2_mux2_1 _21074_ (.A0(\cpu.ex.r_15[11] ),
    .A1(net835),
    .S(net592),
    .X(_00881_));
 sg13g2_mux2_1 _21075_ (.A0(\cpu.ex.r_15[12] ),
    .A1(_03583_),
    .S(net592),
    .X(_00882_));
 sg13g2_mux2_1 _21076_ (.A0(\cpu.ex.r_15[13] ),
    .A1(net458),
    .S(net592),
    .X(_00883_));
 sg13g2_mux2_1 _21077_ (.A0(\cpu.ex.r_15[14] ),
    .A1(net456),
    .S(net592),
    .X(_00884_));
 sg13g2_mux2_1 _21078_ (.A0(\cpu.ex.r_15[15] ),
    .A1(net720),
    .S(net592),
    .X(_00885_));
 sg13g2_mux2_1 _21079_ (.A0(\cpu.ex.r_15[1] ),
    .A1(net457),
    .S(_03621_),
    .X(_00886_));
 sg13g2_mux2_1 _21080_ (.A0(\cpu.ex.r_15[2] ),
    .A1(net519),
    .S(net592),
    .X(_00887_));
 sg13g2_mux2_1 _21081_ (.A0(\cpu.ex.r_15[3] ),
    .A1(net518),
    .S(net592),
    .X(_00888_));
 sg13g2_mux2_1 _21082_ (.A0(\cpu.ex.r_15[4] ),
    .A1(_03594_),
    .S(_03620_),
    .X(_00889_));
 sg13g2_mux2_1 _21083_ (.A0(\cpu.ex.r_15[5] ),
    .A1(net593),
    .S(_03620_),
    .X(_00890_));
 sg13g2_mux2_1 _21084_ (.A0(\cpu.ex.r_15[6] ),
    .A1(net723),
    .S(_03620_),
    .X(_00891_));
 sg13g2_mux2_1 _21085_ (.A0(\cpu.ex.r_15[7] ),
    .A1(net719),
    .S(_03620_),
    .X(_00892_));
 sg13g2_mux2_1 _21086_ (.A0(\cpu.ex.r_15[8] ),
    .A1(net722),
    .S(_03620_),
    .X(_00893_));
 sg13g2_mux2_1 _21087_ (.A0(\cpu.ex.r_15[9] ),
    .A1(net837),
    .S(_03620_),
    .X(_00894_));
 sg13g2_nor3_1 _21088_ (.A(net1019),
    .B(net1018),
    .C(_03578_),
    .Y(_03622_));
 sg13g2_buf_4 _21089_ (.X(_03623_),
    .A(_03622_));
 sg13g2_buf_1 _21090_ (.A(_03623_),
    .X(_03624_));
 sg13g2_mux2_1 _21091_ (.A0(\cpu.ex.r_8[0] ),
    .A1(net833),
    .S(net513),
    .X(_00895_));
 sg13g2_nand2_1 _21092_ (.Y(_03625_),
    .A(net968),
    .B(_03623_));
 sg13g2_o21ai_1 _21093_ (.B1(_03625_),
    .Y(_00896_),
    .A1(_11169_),
    .A2(net513));
 sg13g2_mux2_1 _21094_ (.A0(\cpu.ex.r_8[11] ),
    .A1(net835),
    .S(net513),
    .X(_00897_));
 sg13g2_mux2_1 _21095_ (.A0(\cpu.ex.r_8[12] ),
    .A1(_03583_),
    .S(_03624_),
    .X(_00898_));
 sg13g2_mux2_1 _21096_ (.A0(\cpu.ex.r_8[13] ),
    .A1(net458),
    .S(net513),
    .X(_00899_));
 sg13g2_mux2_1 _21097_ (.A0(\cpu.ex.r_8[14] ),
    .A1(net456),
    .S(net513),
    .X(_00900_));
 sg13g2_mux2_1 _21098_ (.A0(\cpu.ex.r_8[15] ),
    .A1(net720),
    .S(net513),
    .X(_00901_));
 sg13g2_mux2_1 _21099_ (.A0(\cpu.ex.r_8[1] ),
    .A1(net457),
    .S(_03624_),
    .X(_00902_));
 sg13g2_mux2_1 _21100_ (.A0(\cpu.ex.r_8[2] ),
    .A1(net519),
    .S(net513),
    .X(_00903_));
 sg13g2_mux2_1 _21101_ (.A0(\cpu.ex.r_8[3] ),
    .A1(net518),
    .S(net513),
    .X(_00904_));
 sg13g2_mux2_1 _21102_ (.A0(\cpu.ex.r_8[4] ),
    .A1(net517),
    .S(_03623_),
    .X(_00905_));
 sg13g2_mux2_1 _21103_ (.A0(\cpu.ex.r_8[5] ),
    .A1(net593),
    .S(_03623_),
    .X(_00906_));
 sg13g2_mux2_1 _21104_ (.A0(\cpu.ex.r_8[6] ),
    .A1(net723),
    .S(_03623_),
    .X(_00907_));
 sg13g2_mux2_1 _21105_ (.A0(\cpu.ex.r_8[7] ),
    .A1(net719),
    .S(_03623_),
    .X(_00908_));
 sg13g2_mux2_1 _21106_ (.A0(\cpu.ex.r_8[8] ),
    .A1(_03018_),
    .S(_03623_),
    .X(_00909_));
 sg13g2_mux2_1 _21107_ (.A0(\cpu.ex.r_8[9] ),
    .A1(net837),
    .S(_03623_),
    .X(_00910_));
 sg13g2_nor2_1 _21108_ (.A(_03578_),
    .B(_03610_),
    .Y(_03626_));
 sg13g2_buf_1 _21109_ (.A(_03626_),
    .X(_03627_));
 sg13g2_buf_1 _21110_ (.A(net591),
    .X(_03628_));
 sg13g2_mux2_1 _21111_ (.A0(\cpu.ex.r_9[0] ),
    .A1(net833),
    .S(net512),
    .X(_00911_));
 sg13g2_mux2_1 _21112_ (.A0(\cpu.ex.r_9[10] ),
    .A1(net836),
    .S(net512),
    .X(_00912_));
 sg13g2_mux2_1 _21113_ (.A0(\cpu.ex.r_9[11] ),
    .A1(_03021_),
    .S(_03628_),
    .X(_00913_));
 sg13g2_buf_1 _21114_ (.A(net522),
    .X(_03629_));
 sg13g2_mux2_1 _21115_ (.A0(\cpu.ex.r_9[12] ),
    .A1(net455),
    .S(net512),
    .X(_00914_));
 sg13g2_buf_1 _21116_ (.A(net521),
    .X(_03630_));
 sg13g2_mux2_1 _21117_ (.A0(\cpu.ex.r_9[13] ),
    .A1(net454),
    .S(net512),
    .X(_00915_));
 sg13g2_mux2_1 _21118_ (.A0(\cpu.ex.r_9[14] ),
    .A1(_03606_),
    .S(net512),
    .X(_00916_));
 sg13g2_mux2_1 _21119_ (.A0(\cpu.ex.r_9[15] ),
    .A1(net720),
    .S(net512),
    .X(_00917_));
 sg13g2_mux2_1 _21120_ (.A0(\cpu.ex.r_9[1] ),
    .A1(net457),
    .S(_03628_),
    .X(_00918_));
 sg13g2_mux2_1 _21121_ (.A0(\cpu.ex.r_9[2] ),
    .A1(net519),
    .S(net591),
    .X(_00919_));
 sg13g2_mux2_1 _21122_ (.A0(\cpu.ex.r_9[3] ),
    .A1(net518),
    .S(net591),
    .X(_00920_));
 sg13g2_mux2_1 _21123_ (.A0(\cpu.ex.r_9[4] ),
    .A1(net517),
    .S(_03627_),
    .X(_00921_));
 sg13g2_mux2_1 _21124_ (.A0(\cpu.ex.r_9[5] ),
    .A1(net593),
    .S(net591),
    .X(_00922_));
 sg13g2_nand2_1 _21125_ (.Y(_03631_),
    .A(net847),
    .B(net591));
 sg13g2_o21ai_1 _21126_ (.B1(_03631_),
    .Y(_00923_),
    .A1(_10796_),
    .A2(net512));
 sg13g2_mux2_1 _21127_ (.A0(\cpu.ex.r_9[7] ),
    .A1(net719),
    .S(net591),
    .X(_00924_));
 sg13g2_mux2_1 _21128_ (.A0(\cpu.ex.r_9[8] ),
    .A1(net722),
    .S(net591),
    .X(_00925_));
 sg13g2_inv_1 _21129_ (.Y(_03632_),
    .A(\cpu.ex.r_9[9] ));
 sg13g2_nand2_1 _21130_ (.Y(_03633_),
    .A(net969),
    .B(net591));
 sg13g2_o21ai_1 _21131_ (.B1(_03633_),
    .Y(_00926_),
    .A1(_03632_),
    .A2(net512));
 sg13g2_a21oi_1 _21132_ (.A1(_08579_),
    .A2(_11544_),
    .Y(_03634_),
    .B1(_11537_));
 sg13g2_buf_1 _21133_ (.A(_03634_),
    .X(_03635_));
 sg13g2_inv_1 _21134_ (.Y(_03636_),
    .A(_00194_));
 sg13g2_inv_1 _21135_ (.Y(_03637_),
    .A(_11906_));
 sg13g2_buf_8 _21136_ (.A(_10577_),
    .X(_03638_));
 sg13g2_nand2_1 _21137_ (.Y(_03639_),
    .A(net1004),
    .B(net281));
 sg13g2_buf_1 _21138_ (.A(_03639_),
    .X(_03640_));
 sg13g2_mux2_1 _21139_ (.A0(_03636_),
    .A1(_03637_),
    .S(net200),
    .X(_03641_));
 sg13g2_buf_1 _21140_ (.A(_03641_),
    .X(_03642_));
 sg13g2_buf_1 _21141_ (.A(_03642_),
    .X(_03643_));
 sg13g2_buf_1 _21142_ (.A(net138),
    .X(_03644_));
 sg13g2_inv_2 _21143_ (.Y(_03645_),
    .A(_00292_));
 sg13g2_a21oi_1 _21144_ (.A1(net861),
    .A2(net281),
    .Y(_03646_),
    .B1(_11891_));
 sg13g2_a21o_1 _21145_ (.A2(_11114_),
    .A1(_03645_),
    .B1(_03646_),
    .X(_03647_));
 sg13g2_buf_1 _21146_ (.A(_03647_),
    .X(_03648_));
 sg13g2_nand2_1 _21147_ (.Y(_03649_),
    .A(net239),
    .B(_03648_));
 sg13g2_buf_1 _21148_ (.A(_03649_),
    .X(_03650_));
 sg13g2_inv_1 _21149_ (.Y(_03651_),
    .A(_00293_));
 sg13g2_nand3_1 _21150_ (.B(_03651_),
    .C(net281),
    .A(net861),
    .Y(_03652_));
 sg13g2_buf_1 _21151_ (.A(_03652_),
    .X(_03653_));
 sg13g2_buf_1 _21152_ (.A(_10736_),
    .X(_03654_));
 sg13g2_o21ai_1 _21153_ (.B1(_11889_),
    .Y(_03655_),
    .A1(net859),
    .A2(net280));
 sg13g2_nand2_1 _21154_ (.Y(_03656_),
    .A(_03653_),
    .B(_03655_));
 sg13g2_buf_2 _21155_ (.A(_03656_),
    .X(_03657_));
 sg13g2_nand2b_1 _21156_ (.Y(_03658_),
    .B(_11393_),
    .A_N(_03657_));
 sg13g2_a21oi_2 _21157_ (.B1(_03646_),
    .Y(_03659_),
    .A2(_11114_),
    .A1(_03645_));
 sg13g2_nand2_1 _21158_ (.Y(_03660_),
    .A(net216),
    .B(_03659_));
 sg13g2_nand2_1 _21159_ (.Y(_03661_),
    .A(_03658_),
    .B(_03660_));
 sg13g2_nand3b_1 _21160_ (.B(_03638_),
    .C(net861),
    .Y(_03662_),
    .A_N(_10981_));
 sg13g2_buf_1 _21161_ (.A(_03662_),
    .X(_03663_));
 sg13g2_inv_1 _21162_ (.Y(_03664_),
    .A(_11890_));
 sg13g2_o21ai_1 _21163_ (.B1(_03664_),
    .Y(_03665_),
    .A1(net859),
    .A2(net280));
 sg13g2_buf_1 _21164_ (.A(_03665_),
    .X(_03666_));
 sg13g2_nand2_1 _21165_ (.Y(_03667_),
    .A(_03663_),
    .B(_03666_));
 sg13g2_buf_2 _21166_ (.A(_03667_),
    .X(_03668_));
 sg13g2_nor2_1 _21167_ (.A(net168),
    .B(_03668_),
    .Y(_03669_));
 sg13g2_nand2_1 _21168_ (.Y(_03670_),
    .A(net194),
    .B(_03657_));
 sg13g2_buf_2 _21169_ (.A(_03670_),
    .X(_03671_));
 sg13g2_and2_1 _21170_ (.A(_03650_),
    .B(_03671_),
    .X(_03672_));
 sg13g2_a22oi_1 _21171_ (.Y(_03673_),
    .B1(_03669_),
    .B2(_03672_),
    .A2(_03661_),
    .A1(_03650_));
 sg13g2_buf_1 _21172_ (.A(_03673_),
    .X(_03674_));
 sg13g2_nand4_1 _21173_ (.B(_03671_),
    .C(_03663_),
    .A(_03650_),
    .Y(_03675_),
    .D(_03666_));
 sg13g2_nand3_1 _21174_ (.B(_03650_),
    .C(_03671_),
    .A(_11675_),
    .Y(_03676_));
 sg13g2_nand3b_1 _21175_ (.B(net281),
    .C(_10662_),
    .Y(_03677_),
    .A_N(_00191_));
 sg13g2_buf_2 _21176_ (.A(_03677_),
    .X(_03678_));
 sg13g2_o21ai_1 _21177_ (.B1(_11044_),
    .Y(_03679_),
    .A1(_10579_),
    .A2(_10736_));
 sg13g2_buf_1 _21178_ (.A(_03679_),
    .X(_03680_));
 sg13g2_nand2_1 _21179_ (.Y(_03681_),
    .A(_03678_),
    .B(_03680_));
 sg13g2_buf_1 _21180_ (.A(_03681_),
    .X(_03682_));
 sg13g2_nand2_1 _21181_ (.Y(_03683_),
    .A(net241),
    .B(_11562_));
 sg13g2_nand3b_1 _21182_ (.B(_11525_),
    .C(net281),
    .Y(_03684_),
    .A_N(net1130));
 sg13g2_buf_2 _21183_ (.A(_03684_),
    .X(_03685_));
 sg13g2_o21ai_1 _21184_ (.B1(_11887_),
    .Y(_03686_),
    .A1(_11909_),
    .A2(net280));
 sg13g2_buf_2 _21185_ (.A(_03686_),
    .X(_03687_));
 sg13g2_a21oi_2 _21186_ (.B1(_11327_),
    .Y(_03688_),
    .A2(_03687_),
    .A1(_03685_));
 sg13g2_a21oi_1 _21187_ (.A1(net167),
    .A2(_03683_),
    .Y(_03689_),
    .B1(_03688_));
 sg13g2_nor3_1 _21188_ (.A(net859),
    .B(_11110_),
    .C(net280),
    .Y(_03690_));
 sg13g2_inv_1 _21189_ (.Y(_03691_),
    .A(_11084_));
 sg13g2_a21oi_1 _21190_ (.A1(net861),
    .A2(net281),
    .Y(_03692_),
    .B1(_03691_));
 sg13g2_nor4_2 _21191_ (.A(_10773_),
    .B(_10776_),
    .C(_11007_),
    .Y(_03693_),
    .D(_11011_));
 sg13g2_o21ai_1 _21192_ (.B1(_03693_),
    .Y(_03694_),
    .A1(_03690_),
    .A2(_03692_));
 sg13g2_nor3_1 _21193_ (.A(_03690_),
    .B(_03692_),
    .C(_03693_),
    .Y(_03695_));
 sg13g2_a21o_1 _21194_ (.A2(_03694_),
    .A1(_10552_),
    .B1(_03695_),
    .X(_03696_));
 sg13g2_o21ai_1 _21195_ (.B1(_11898_),
    .Y(_03697_),
    .A1(net859),
    .A2(net280));
 sg13g2_o21ai_1 _21196_ (.B1(_03697_),
    .Y(_03698_),
    .A1(_00295_),
    .A2(net200));
 sg13g2_buf_2 _21197_ (.A(_03698_),
    .X(_03699_));
 sg13g2_a221oi_1 _21198_ (.B2(net240),
    .C1(_03688_),
    .B1(net167),
    .A1(_03699_),
    .Y(_03700_),
    .A2(_10505_));
 sg13g2_nand4_1 _21199_ (.B(_11562_),
    .C(_03678_),
    .A(_10665_),
    .Y(_03701_),
    .D(_03680_));
 sg13g2_nand3_1 _21200_ (.B(_03685_),
    .C(_03687_),
    .A(_11327_),
    .Y(_03702_));
 sg13g2_buf_1 _21201_ (.A(_03702_),
    .X(_03703_));
 sg13g2_o21ai_1 _21202_ (.B1(_03703_),
    .Y(_03704_),
    .A1(_03688_),
    .A2(_03701_));
 sg13g2_a221oi_1 _21203_ (.B2(_03700_),
    .C1(_03704_),
    .B1(_03696_),
    .A1(net237),
    .Y(_03705_),
    .A2(_03689_));
 sg13g2_buf_2 _21204_ (.A(_03705_),
    .X(_03706_));
 sg13g2_a21o_1 _21205_ (.A2(_03676_),
    .A1(_03675_),
    .B1(_03706_),
    .X(_03707_));
 sg13g2_buf_1 _21206_ (.A(_03707_),
    .X(_03708_));
 sg13g2_nor3_1 _21207_ (.A(net859),
    .B(_11109_),
    .C(net280),
    .Y(_03709_));
 sg13g2_a21o_1 _21208_ (.A2(_11106_),
    .A1(net200),
    .B1(_03709_),
    .X(_03710_));
 sg13g2_buf_1 _21209_ (.A(_03710_),
    .X(_03711_));
 sg13g2_nand2_2 _21210_ (.Y(_03712_),
    .A(net215),
    .B(_03711_));
 sg13g2_nor3_1 _21211_ (.A(net859),
    .B(_00291_),
    .C(_03654_),
    .Y(_03713_));
 sg13g2_a21oi_2 _21212_ (.B1(_03713_),
    .Y(_03714_),
    .A2(_10701_),
    .A1(net200));
 sg13g2_nand2_1 _21213_ (.Y(_03715_),
    .A(_03712_),
    .B(_03714_));
 sg13g2_nand2_1 _21214_ (.Y(_03716_),
    .A(net190),
    .B(_03712_));
 sg13g2_a22oi_1 _21215_ (.Y(_03717_),
    .B1(_03715_),
    .B2(_03716_),
    .A2(_03708_),
    .A1(_03674_));
 sg13g2_inv_1 _21216_ (.Y(_03718_),
    .A(_03712_));
 sg13g2_nand2_1 _21217_ (.Y(_03719_),
    .A(net190),
    .B(_03714_));
 sg13g2_a21oi_2 _21218_ (.B1(_03709_),
    .Y(_03720_),
    .A2(_11106_),
    .A1(net200));
 sg13g2_nand2_1 _21219_ (.Y(_03721_),
    .A(net217),
    .B(_03720_));
 sg13g2_o21ai_1 _21220_ (.B1(_03721_),
    .Y(_03722_),
    .A1(_03718_),
    .A2(_03719_));
 sg13g2_inv_1 _21221_ (.Y(_03723_),
    .A(_00287_));
 sg13g2_a21oi_1 _21222_ (.A1(net861),
    .A2(_03638_),
    .Y(_03724_),
    .B1(_10858_));
 sg13g2_a21o_1 _21223_ (.A2(_11114_),
    .A1(_03723_),
    .B1(_03724_),
    .X(_03725_));
 sg13g2_buf_1 _21224_ (.A(_03725_),
    .X(_03726_));
 sg13g2_nand2b_1 _21225_ (.Y(_03727_),
    .B(net213),
    .A_N(_03726_));
 sg13g2_buf_1 _21226_ (.A(_03727_),
    .X(_03728_));
 sg13g2_nand3b_1 _21227_ (.B(net281),
    .C(net861),
    .Y(_03729_),
    .A_N(_10738_));
 sg13g2_buf_1 _21228_ (.A(_03729_),
    .X(_03730_));
 sg13g2_o21ai_1 _21229_ (.B1(_10730_),
    .Y(_03731_),
    .A1(net859),
    .A2(net280));
 sg13g2_and2_1 _21230_ (.A(_03730_),
    .B(_03731_),
    .X(_03732_));
 sg13g2_buf_1 _21231_ (.A(_03732_),
    .X(_03733_));
 sg13g2_nand2_1 _21232_ (.Y(_03734_),
    .A(net214),
    .B(_03733_));
 sg13g2_nor3_1 _21233_ (.A(net859),
    .B(_00288_),
    .C(_03654_),
    .Y(_03735_));
 sg13g2_a21oi_2 _21234_ (.B1(_03735_),
    .Y(_03736_),
    .A2(_11061_),
    .A1(net200));
 sg13g2_nand2_2 _21235_ (.Y(_03737_),
    .A(net211),
    .B(_03736_));
 sg13g2_nand3_1 _21236_ (.B(_03734_),
    .C(_03737_),
    .A(_03728_),
    .Y(_03738_));
 sg13g2_nor3_2 _21237_ (.A(_03717_),
    .B(_03722_),
    .C(_03738_),
    .Y(_03739_));
 sg13g2_inv_1 _21238_ (.Y(_03740_),
    .A(_03728_));
 sg13g2_a21o_1 _21239_ (.A2(_11061_),
    .A1(_03640_),
    .B1(_03735_),
    .X(_03741_));
 sg13g2_buf_2 _21240_ (.A(_03741_),
    .X(_03742_));
 sg13g2_nand2_1 _21241_ (.Y(_03743_),
    .A(net212),
    .B(_03742_));
 sg13g2_nor2_1 _21242_ (.A(net214),
    .B(_03733_),
    .Y(_03744_));
 sg13g2_nand3_1 _21243_ (.B(_03744_),
    .C(_03737_),
    .A(_03728_),
    .Y(_03745_));
 sg13g2_o21ai_1 _21244_ (.B1(_03745_),
    .Y(_03746_),
    .A1(_03740_),
    .A2(_03743_));
 sg13g2_buf_1 _21245_ (.A(_03746_),
    .X(_03747_));
 sg13g2_inv_1 _21246_ (.Y(_03748_),
    .A(_00195_));
 sg13g2_inv_1 _21247_ (.Y(_03749_),
    .A(_11897_));
 sg13g2_mux2_1 _21248_ (.A0(_03748_),
    .A1(_03749_),
    .S(net200),
    .X(_03750_));
 sg13g2_buf_1 _21249_ (.A(_03750_),
    .X(_03751_));
 sg13g2_buf_1 _21250_ (.A(_03751_),
    .X(_03752_));
 sg13g2_buf_1 _21251_ (.A(_03726_),
    .X(_03753_));
 sg13g2_nand2_1 _21252_ (.Y(_03754_),
    .A(_10383_),
    .B(net165));
 sg13g2_inv_1 _21253_ (.Y(_03755_),
    .A(_00196_));
 sg13g2_mux2_1 _21254_ (.A0(_03755_),
    .A1(_11900_),
    .S(net200),
    .X(_03756_));
 sg13g2_buf_1 _21255_ (.A(_03756_),
    .X(_03757_));
 sg13g2_nand2b_1 _21256_ (.Y(_03758_),
    .B(net164),
    .A_N(net170));
 sg13g2_buf_1 _21257_ (.A(_03758_),
    .X(_03759_));
 sg13g2_nand2_1 _21258_ (.Y(_03760_),
    .A(_03754_),
    .B(_03759_));
 sg13g2_nor4_1 _21259_ (.A(_03739_),
    .B(_03747_),
    .C(net137),
    .D(_03760_),
    .Y(_03761_));
 sg13g2_nor4_1 _21260_ (.A(net192),
    .B(_03739_),
    .C(_03747_),
    .D(_03760_),
    .Y(_03762_));
 sg13g2_inv_1 _21261_ (.Y(_03763_),
    .A(net164));
 sg13g2_nand2_1 _21262_ (.Y(_03764_),
    .A(net170),
    .B(_03763_));
 sg13g2_a21oi_1 _21263_ (.A1(_11470_),
    .A2(net137),
    .Y(_03765_),
    .B1(_03764_));
 sg13g2_nor2_1 _21264_ (.A(_11114_),
    .B(_11897_),
    .Y(_03766_));
 sg13g2_a21oi_2 _21265_ (.B1(_03766_),
    .Y(_03767_),
    .A2(_11114_),
    .A1(_03748_));
 sg13g2_nand2_2 _21266_ (.Y(_03768_),
    .A(_11476_),
    .B(_03767_));
 sg13g2_nand2b_1 _21267_ (.Y(_03769_),
    .B(_03768_),
    .A_N(_03765_));
 sg13g2_nor3_2 _21268_ (.A(_03761_),
    .B(_03762_),
    .C(_03769_),
    .Y(_03770_));
 sg13g2_o21ai_1 _21269_ (.B1(net169),
    .Y(_03771_),
    .A1(net114),
    .A2(_03770_));
 sg13g2_a21oi_1 _21270_ (.A1(net114),
    .A2(_03770_),
    .Y(_03772_),
    .B1(net1045));
 sg13g2_inv_1 _21271_ (.Y(_03773_),
    .A(_03642_));
 sg13g2_buf_1 _21272_ (.A(_03757_),
    .X(_03774_));
 sg13g2_or2_1 _21273_ (.X(_03775_),
    .B(net136),
    .A(_10330_));
 sg13g2_buf_1 _21274_ (.A(_03775_),
    .X(_03776_));
 sg13g2_nand2_1 _21275_ (.Y(_03777_),
    .A(_10330_),
    .B(net136));
 sg13g2_nand3b_1 _21276_ (.B(net281),
    .C(_10662_),
    .Y(_03778_),
    .A_N(_11110_));
 sg13g2_buf_1 _21277_ (.A(_03778_),
    .X(_03779_));
 sg13g2_o21ai_1 _21278_ (.B1(_11084_),
    .Y(_03780_),
    .A1(_10579_),
    .A2(net280));
 sg13g2_buf_1 _21279_ (.A(_03780_),
    .X(_03781_));
 sg13g2_nand3_1 _21280_ (.B(_03779_),
    .C(_03781_),
    .A(_11550_),
    .Y(_03782_));
 sg13g2_nor2_1 _21281_ (.A(_10773_),
    .B(_10776_),
    .Y(_03783_));
 sg13g2_nor2_2 _21282_ (.A(_11007_),
    .B(_11011_),
    .Y(_03784_));
 sg13g2_nand2b_1 _21283_ (.Y(_03785_),
    .B(_03784_),
    .A_N(_03783_));
 sg13g2_a21oi_1 _21284_ (.A1(_03779_),
    .A2(_03781_),
    .Y(_03786_),
    .B1(_11550_));
 sg13g2_a221oi_1 _21285_ (.B2(_03785_),
    .C1(_03786_),
    .B1(_03782_),
    .A1(_03699_),
    .Y(_03787_),
    .A2(_11562_));
 sg13g2_buf_1 _21286_ (.A(_03787_),
    .X(_03788_));
 sg13g2_a21oi_1 _21287_ (.A1(_03685_),
    .A2(_03687_),
    .Y(_03789_),
    .B1(_11332_));
 sg13g2_a21o_1 _21288_ (.A2(_11327_),
    .A1(_11887_),
    .B1(_11044_),
    .X(_03790_));
 sg13g2_o21ai_1 _21289_ (.B1(_00191_),
    .Y(_03791_),
    .A1(_08316_),
    .A2(net287));
 sg13g2_mux2_1 _21290_ (.A0(_03790_),
    .A1(_03791_),
    .S(_11114_),
    .X(_03792_));
 sg13g2_o21ai_1 _21291_ (.B1(_03792_),
    .Y(_03793_),
    .A1(_11593_),
    .A2(_03789_));
 sg13g2_nand3_1 _21292_ (.B(_03685_),
    .C(_03687_),
    .A(_11332_),
    .Y(_03794_));
 sg13g2_nand3_1 _21293_ (.B(_03678_),
    .C(_03680_),
    .A(_10513_),
    .Y(_03795_));
 sg13g2_nand4_1 _21294_ (.B(_10505_),
    .C(_03678_),
    .A(net241),
    .Y(_03796_),
    .D(_03680_));
 sg13g2_nand3_1 _21295_ (.B(_10513_),
    .C(_10505_),
    .A(net241),
    .Y(_03797_));
 sg13g2_nand4_1 _21296_ (.B(_03795_),
    .C(_03796_),
    .A(_03794_),
    .Y(_03798_),
    .D(_03797_));
 sg13g2_buf_1 _21297_ (.A(_03798_),
    .X(_03799_));
 sg13g2_nand2_1 _21298_ (.Y(_03800_),
    .A(_03685_),
    .B(_03687_));
 sg13g2_buf_1 _21299_ (.A(_03800_),
    .X(_03801_));
 sg13g2_nand2_1 _21300_ (.Y(_03802_),
    .A(_11327_),
    .B(_03801_));
 sg13g2_buf_1 _21301_ (.A(_03648_),
    .X(_03803_));
 sg13g2_nand4_1 _21302_ (.B(_11260_),
    .C(_03653_),
    .A(_11234_),
    .Y(_03804_),
    .D(_03655_));
 sg13g2_buf_1 _21303_ (.A(_03804_),
    .X(_03805_));
 sg13g2_nand4_1 _21304_ (.B(_11673_),
    .C(_03663_),
    .A(_11671_),
    .Y(_03806_),
    .D(_03666_));
 sg13g2_buf_1 _21305_ (.A(_03806_),
    .X(_03807_));
 sg13g2_nand3_1 _21306_ (.B(_03805_),
    .C(_03807_),
    .A(_03803_),
    .Y(_03808_));
 sg13g2_a221oi_1 _21307_ (.B2(_03802_),
    .C1(_03808_),
    .B1(_03799_),
    .A1(_03788_),
    .Y(_03809_),
    .A2(_03793_));
 sg13g2_nand3_1 _21308_ (.B(_03805_),
    .C(_03807_),
    .A(_11295_),
    .Y(_03810_));
 sg13g2_a221oi_1 _21309_ (.B2(_03802_),
    .C1(_03810_),
    .B1(_03799_),
    .A1(_03788_),
    .Y(_03811_),
    .A2(_03793_));
 sg13g2_nor2_1 _21310_ (.A(net239),
    .B(_03659_),
    .Y(_03812_));
 sg13g2_a22oi_1 _21311_ (.Y(_03813_),
    .B1(_03663_),
    .B2(_03666_),
    .A2(_11673_),
    .A1(_11671_));
 sg13g2_a22oi_1 _21312_ (.Y(_03814_),
    .B1(_03653_),
    .B2(_03655_),
    .A2(_11260_),
    .A1(_11234_));
 sg13g2_o21ai_1 _21313_ (.B1(_03805_),
    .Y(_03815_),
    .A1(_03813_),
    .A2(_03814_));
 sg13g2_a21oi_1 _21314_ (.A1(_11301_),
    .A2(_03659_),
    .Y(_03816_),
    .B1(_03815_));
 sg13g2_nor4_1 _21315_ (.A(_03809_),
    .B(_03811_),
    .C(_03812_),
    .D(_03816_),
    .Y(_03817_));
 sg13g2_buf_2 _21316_ (.A(_03817_),
    .X(_03818_));
 sg13g2_a21oi_1 _21317_ (.A1(_03730_),
    .A2(_03731_),
    .Y(_03819_),
    .B1(_11191_));
 sg13g2_nand2_1 _21318_ (.Y(_03820_),
    .A(_03742_),
    .B(_03819_));
 sg13g2_o21ai_1 _21319_ (.B1(_10417_),
    .Y(_03821_),
    .A1(_03742_),
    .A2(_03819_));
 sg13g2_and2_1 _21320_ (.A(_03820_),
    .B(_03821_),
    .X(_03822_));
 sg13g2_buf_1 _21321_ (.A(_03822_),
    .X(_03823_));
 sg13g2_nand2_1 _21322_ (.Y(_03824_),
    .A(net217),
    .B(_03711_));
 sg13g2_a21o_1 _21323_ (.A2(_10701_),
    .A1(_03640_),
    .B1(_03713_),
    .X(_03825_));
 sg13g2_buf_1 _21324_ (.A(_03825_),
    .X(_03826_));
 sg13g2_nand2_1 _21325_ (.Y(_03827_),
    .A(net190),
    .B(_03826_));
 sg13g2_buf_1 _21326_ (.A(_03827_),
    .X(_03828_));
 sg13g2_and3_1 _21327_ (.X(_03829_),
    .A(_03823_),
    .B(_03824_),
    .C(_03828_));
 sg13g2_nor2_1 _21328_ (.A(net215),
    .B(_03720_),
    .Y(_03830_));
 sg13g2_a22oi_1 _21329_ (.Y(_03831_),
    .B1(_03714_),
    .B2(_11719_),
    .A2(_03720_),
    .A1(_11372_));
 sg13g2_a22oi_1 _21330_ (.Y(_03832_),
    .B1(_03733_),
    .B2(net188),
    .A2(_03736_),
    .A1(net212));
 sg13g2_o21ai_1 _21331_ (.B1(_03832_),
    .Y(_03833_),
    .A1(_03830_),
    .A2(_03831_));
 sg13g2_nor2_2 _21332_ (.A(net213),
    .B(_03726_),
    .Y(_03834_));
 sg13g2_a21o_1 _21333_ (.A2(_03833_),
    .A1(_03823_),
    .B1(_03834_),
    .X(_03835_));
 sg13g2_a21o_1 _21334_ (.A2(_03829_),
    .A1(_03818_),
    .B1(_03835_),
    .X(_03836_));
 sg13g2_nand2_1 _21335_ (.Y(_03837_),
    .A(_11400_),
    .B(net165));
 sg13g2_nand3_1 _21336_ (.B(_03836_),
    .C(_03837_),
    .A(_03777_),
    .Y(_03838_));
 sg13g2_a22oi_1 _21337_ (.Y(_03839_),
    .B1(_03776_),
    .B2(_03838_),
    .A2(net137),
    .A1(_11476_));
 sg13g2_nor2_1 _21338_ (.A(_11476_),
    .B(net137),
    .Y(_03840_));
 sg13g2_or2_1 _21339_ (.X(_03841_),
    .B(_03840_),
    .A(_03839_));
 sg13g2_o21ai_1 _21340_ (.B1(net169),
    .Y(_03842_),
    .A1(_03773_),
    .A2(_03841_));
 sg13g2_inv_1 _21341_ (.Y(_03843_),
    .A(_09180_));
 sg13g2_buf_1 _21342_ (.A(_03843_),
    .X(_03844_));
 sg13g2_a21oi_1 _21343_ (.A1(_03773_),
    .A2(_03841_),
    .Y(_03845_),
    .B1(net832));
 sg13g2_a221oi_1 _21344_ (.B2(_03845_),
    .C1(_03635_),
    .B1(_03842_),
    .A1(_03771_),
    .Y(_03846_),
    .A2(_03772_));
 sg13g2_a21o_1 _21345_ (.A2(net83),
    .A1(\cpu.ex.r_cc ),
    .B1(_03846_),
    .X(_00927_));
 sg13g2_nor2_1 _21346_ (.A(net1111),
    .B(net1110),
    .Y(_03847_));
 sg13g2_nand4_1 _21347_ (.B(_10232_),
    .C(net1112),
    .A(net1019),
    .Y(_03848_),
    .D(_03847_));
 sg13g2_nor2_1 _21348_ (.A(_08476_),
    .B(_03848_),
    .Y(_03849_));
 sg13g2_buf_2 _21349_ (.A(_03849_),
    .X(_03850_));
 sg13g2_buf_1 _21350_ (.A(_03850_),
    .X(_03851_));
 sg13g2_mux2_1 _21351_ (.A0(\cpu.ex.r_epc[1] ),
    .A1(_03589_),
    .S(net590),
    .X(_00929_));
 sg13g2_mux2_1 _21352_ (.A0(\cpu.ex.r_epc[11] ),
    .A1(net835),
    .S(net590),
    .X(_00930_));
 sg13g2_mux2_1 _21353_ (.A0(\cpu.ex.r_epc[12] ),
    .A1(net455),
    .S(net590),
    .X(_00931_));
 sg13g2_mux2_1 _21354_ (.A0(\cpu.ex.r_epc[13] ),
    .A1(net454),
    .S(net590),
    .X(_00932_));
 sg13g2_mux2_1 _21355_ (.A0(\cpu.ex.r_epc[14] ),
    .A1(_03606_),
    .S(net590),
    .X(_00933_));
 sg13g2_nand2_1 _21356_ (.Y(_03852_),
    .A(net860),
    .B(_03850_));
 sg13g2_o21ai_1 _21357_ (.B1(_03852_),
    .Y(_00934_),
    .A1(_11427_),
    .A2(_03851_));
 sg13g2_mux2_1 _21358_ (.A0(\cpu.ex.r_epc[2] ),
    .A1(net519),
    .S(net590),
    .X(_00935_));
 sg13g2_mux2_1 _21359_ (.A0(\cpu.ex.r_epc[3] ),
    .A1(_03592_),
    .S(_03851_),
    .X(_00936_));
 sg13g2_mux2_1 _21360_ (.A0(\cpu.ex.r_epc[4] ),
    .A1(net517),
    .S(net590),
    .X(_00937_));
 sg13g2_mux2_1 _21361_ (.A0(\cpu.ex.r_epc[5] ),
    .A1(net593),
    .S(net590),
    .X(_00938_));
 sg13g2_mux2_1 _21362_ (.A0(\cpu.ex.r_epc[6] ),
    .A1(net723),
    .S(_03850_),
    .X(_00939_));
 sg13g2_mux2_1 _21363_ (.A0(\cpu.ex.r_epc[7] ),
    .A1(net719),
    .S(_03850_),
    .X(_00940_));
 sg13g2_mux2_1 _21364_ (.A0(\cpu.ex.r_epc[8] ),
    .A1(net722),
    .S(_03850_),
    .X(_00941_));
 sg13g2_mux2_1 _21365_ (.A0(\cpu.ex.r_epc[9] ),
    .A1(net837),
    .S(_03850_),
    .X(_00942_));
 sg13g2_mux2_1 _21366_ (.A0(\cpu.ex.r_epc[10] ),
    .A1(net836),
    .S(_03850_),
    .X(_00943_));
 sg13g2_nand4_1 _21367_ (.B(net1018),
    .C(net1112),
    .A(_03609_),
    .Y(_03853_),
    .D(_03847_));
 sg13g2_buf_1 _21368_ (.A(_03853_),
    .X(_03854_));
 sg13g2_buf_1 _21369_ (.A(_03854_),
    .X(_03855_));
 sg13g2_buf_1 _21370_ (.A(_03854_),
    .X(_03856_));
 sg13g2_nand2_1 _21371_ (.Y(_03857_),
    .A(\cpu.ex.r_lr[1] ),
    .B(net588));
 sg13g2_o21ai_1 _21372_ (.B1(_03857_),
    .Y(_00949_),
    .A1(net536),
    .A2(net589));
 sg13g2_mux2_1 _21373_ (.A0(_02989_),
    .A1(\cpu.ex.r_lr[11] ),
    .S(_03855_),
    .X(_00950_));
 sg13g2_buf_1 _21374_ (.A(net522),
    .X(_03858_));
 sg13g2_mux2_1 _21375_ (.A0(_03858_),
    .A1(\cpu.ex.r_lr[12] ),
    .S(net589),
    .X(_00951_));
 sg13g2_buf_1 _21376_ (.A(net521),
    .X(_03859_));
 sg13g2_mux2_1 _21377_ (.A0(net452),
    .A1(\cpu.ex.r_lr[13] ),
    .S(net589),
    .X(_00952_));
 sg13g2_buf_1 _21378_ (.A(net520),
    .X(_03860_));
 sg13g2_mux2_1 _21379_ (.A0(_03860_),
    .A1(\cpu.ex.r_lr[14] ),
    .S(net588),
    .X(_00953_));
 sg13g2_buf_1 _21380_ (.A(net676),
    .X(_03861_));
 sg13g2_nand2_1 _21381_ (.Y(_03862_),
    .A(\cpu.ex.r_lr[15] ),
    .B(net588));
 sg13g2_o21ai_1 _21382_ (.B1(_03862_),
    .Y(_00954_),
    .A1(net587),
    .A2(net589));
 sg13g2_nand2_1 _21383_ (.Y(_03863_),
    .A(\cpu.ex.r_lr[2] ),
    .B(_03856_));
 sg13g2_o21ai_1 _21384_ (.B1(_03863_),
    .Y(_00955_),
    .A1(net767),
    .A2(net589));
 sg13g2_nand2_1 _21385_ (.Y(_03864_),
    .A(\cpu.ex.r_lr[3] ),
    .B(net588));
 sg13g2_o21ai_1 _21386_ (.B1(_03864_),
    .Y(_00956_),
    .A1(net780),
    .A2(net589));
 sg13g2_buf_1 _21387_ (.A(net733),
    .X(_03865_));
 sg13g2_buf_1 _21388_ (.A(net650),
    .X(_03866_));
 sg13g2_nand2_1 _21389_ (.Y(_03867_),
    .A(\cpu.ex.r_lr[4] ),
    .B(net588));
 sg13g2_o21ai_1 _21390_ (.B1(_03867_),
    .Y(_00957_),
    .A1(net586),
    .A2(net589));
 sg13g2_nand2_1 _21391_ (.Y(_03868_),
    .A(\cpu.ex.r_lr[5] ),
    .B(_03854_));
 sg13g2_o21ai_1 _21392_ (.B1(_03868_),
    .Y(_00958_),
    .A1(_02971_),
    .A2(_03855_));
 sg13g2_mux2_1 _21393_ (.A0(_02978_),
    .A1(\cpu.ex.r_lr[6] ),
    .S(net588),
    .X(_00959_));
 sg13g2_nand2_1 _21394_ (.Y(_03869_),
    .A(\cpu.ex.r_lr[7] ),
    .B(_03854_));
 sg13g2_o21ai_1 _21395_ (.B1(_03869_),
    .Y(_00960_),
    .A1(net728),
    .A2(net589));
 sg13g2_mux2_1 _21396_ (.A0(_02983_),
    .A1(\cpu.ex.r_lr[8] ),
    .S(_03856_),
    .X(_00961_));
 sg13g2_mux2_1 _21397_ (.A0(net844),
    .A1(\cpu.ex.r_lr[9] ),
    .S(net588),
    .X(_00962_));
 sg13g2_mux2_1 _21398_ (.A0(net843),
    .A1(\cpu.ex.r_lr[10] ),
    .S(net588),
    .X(_00963_));
 sg13g2_nor3_1 _21399_ (.A(_11473_),
    .B(_11475_),
    .C(_11478_),
    .Y(_03870_));
 sg13g2_buf_2 _21400_ (.A(_03870_),
    .X(_03871_));
 sg13g2_buf_8 _21401_ (.A(_03871_),
    .X(_03872_));
 sg13g2_nor2_1 _21402_ (.A(net286),
    .B(net27),
    .Y(_03873_));
 sg13g2_xnor2_1 _21403_ (.Y(_03874_),
    .A(net84),
    .B(_03873_));
 sg13g2_o21ai_1 _21404_ (.B1(_11874_),
    .Y(_03875_),
    .A1(net169),
    .A2(_11863_));
 sg13g2_nand2_1 _21405_ (.Y(_03876_),
    .A(net169),
    .B(_11863_));
 sg13g2_a21oi_1 _21406_ (.A1(_03875_),
    .A2(_03876_),
    .Y(_03877_),
    .B1(_11507_));
 sg13g2_inv_1 _21407_ (.Y(_03878_),
    .A(_00171_));
 sg13g2_o21ai_1 _21408_ (.B1(_11855_),
    .Y(_03879_),
    .A1(_03878_),
    .A2(_11873_));
 sg13g2_o21ai_1 _21409_ (.B1(_11856_),
    .Y(_03880_),
    .A1(net169),
    .A2(_11874_));
 sg13g2_a221oi_1 _21410_ (.B2(_03880_),
    .C1(_11843_),
    .B1(_03879_),
    .A1(_11750_),
    .Y(_03881_),
    .A2(_11758_));
 sg13g2_a21oi_1 _21411_ (.A1(_03879_),
    .A2(_03880_),
    .Y(_03882_),
    .B1(_11853_));
 sg13g2_nor3_1 _21412_ (.A(_03877_),
    .B(_03881_),
    .C(_03882_),
    .Y(_03883_));
 sg13g2_buf_2 _21413_ (.A(_03883_),
    .X(_03884_));
 sg13g2_nand2_1 _21414_ (.Y(_03885_),
    .A(_11861_),
    .B(net606));
 sg13g2_xnor2_1 _21415_ (.Y(_03886_),
    .A(_03884_),
    .B(_03885_));
 sg13g2_buf_1 _21416_ (.A(_10234_),
    .X(_03887_));
 sg13g2_buf_1 _21417_ (.A(_03887_),
    .X(_03888_));
 sg13g2_nor2_1 _21418_ (.A(net535),
    .B(_11517_),
    .Y(_03889_));
 sg13g2_buf_1 _21419_ (.A(_03889_),
    .X(_03890_));
 sg13g2_nand3_1 _21420_ (.B(_10223_),
    .C(\cpu.ex.r_cc ),
    .A(_10222_),
    .Y(_03891_));
 sg13g2_nor2_1 _21421_ (.A(net649),
    .B(_03891_),
    .Y(_03892_));
 sg13g2_a221oi_1 _21422_ (.B2(\cpu.ex.r_mult[16] ),
    .C1(_03892_),
    .B1(_03890_),
    .A1(_03572_),
    .Y(_03893_),
    .A2(net585));
 sg13g2_o21ai_1 _21423_ (.B1(_03893_),
    .Y(_03894_),
    .A1(_11663_),
    .A2(_03886_));
 sg13g2_a21o_1 _21424_ (.A2(_03874_),
    .A1(net58),
    .B1(_03894_),
    .X(_00964_));
 sg13g2_nand2_1 _21425_ (.Y(_03895_),
    .A(_11515_),
    .B(net85));
 sg13g2_buf_1 _21426_ (.A(_03895_),
    .X(_03896_));
 sg13g2_buf_1 _21427_ (.A(_03896_),
    .X(_03897_));
 sg13g2_nor2_1 _21428_ (.A(net115),
    .B(net286),
    .Y(_03898_));
 sg13g2_xnor2_1 _21429_ (.Y(_03899_),
    .A(net238),
    .B(_03898_));
 sg13g2_nor2_1 _21430_ (.A(net27),
    .B(_03899_),
    .Y(_03900_));
 sg13g2_xnor2_1 _21431_ (.Y(_03901_),
    .A(_10519_),
    .B(_03900_));
 sg13g2_nor2_1 _21432_ (.A(net530),
    .B(_11663_),
    .Y(_03902_));
 sg13g2_buf_1 _21433_ (.A(_03902_),
    .X(_03903_));
 sg13g2_nor2_2 _21434_ (.A(_03884_),
    .B(_03885_),
    .Y(_03904_));
 sg13g2_xnor2_1 _21435_ (.Y(_03905_),
    .A(_10518_),
    .B(_03904_));
 sg13g2_or2_1 _21436_ (.X(_03906_),
    .B(_03891_),
    .A(_03844_));
 sg13g2_or2_1 _21437_ (.X(_03907_),
    .B(_11517_),
    .A(_10236_));
 sg13g2_o21ai_1 _21438_ (.B1(_03907_),
    .Y(_03908_),
    .A1(net649),
    .A2(_03906_));
 sg13g2_buf_2 _21439_ (.A(_03908_),
    .X(_03909_));
 sg13g2_buf_1 _21440_ (.A(_03909_),
    .X(_03910_));
 sg13g2_a21oi_1 _21441_ (.A1(net538),
    .A2(net649),
    .Y(_03911_),
    .B1(net364));
 sg13g2_a21oi_1 _21442_ (.A1(_10524_),
    .A2(_03890_),
    .Y(_03912_),
    .B1(_03911_));
 sg13g2_a21oi_1 _21443_ (.A1(net332),
    .A2(_03905_),
    .Y(_03913_),
    .B1(_03912_));
 sg13g2_o21ai_1 _21444_ (.B1(_03913_),
    .Y(_00965_),
    .A1(net31),
    .A2(_03901_));
 sg13g2_or4_1 _21445_ (.A(_10553_),
    .B(_11014_),
    .C(_11116_),
    .D(_11117_),
    .X(_03914_));
 sg13g2_buf_1 _21446_ (.A(_10505_),
    .X(_03915_));
 sg13g2_nand2_1 _21447_ (.Y(_03916_),
    .A(_03914_),
    .B(net279));
 sg13g2_nand2_1 _21448_ (.Y(_03917_),
    .A(_11118_),
    .B(net285));
 sg13g2_nand3_1 _21449_ (.B(_03917_),
    .C(net28),
    .A(_03916_),
    .Y(_03918_));
 sg13g2_nor2_1 _21450_ (.A(_10514_),
    .B(net628),
    .Y(_03919_));
 sg13g2_xor2_1 _21451_ (.B(_03919_),
    .A(_03918_),
    .X(_03920_));
 sg13g2_buf_1 _21452_ (.A(_03890_),
    .X(_03921_));
 sg13g2_nand2b_1 _21453_ (.Y(_03922_),
    .B(net363),
    .A_N(\cpu.ex.r_mult[18] ));
 sg13g2_a21o_1 _21454_ (.A2(net585),
    .A1(net596),
    .B1(net364),
    .X(_03923_));
 sg13g2_nor3_1 _21455_ (.A(_10518_),
    .B(_03884_),
    .C(_03885_),
    .Y(_03924_));
 sg13g2_xnor2_1 _21456_ (.Y(_03925_),
    .A(_10514_),
    .B(_03924_));
 sg13g2_a22oi_1 _21457_ (.Y(_03926_),
    .B1(_03925_),
    .B2(net332),
    .A2(_03923_),
    .A1(_03922_));
 sg13g2_o21ai_1 _21458_ (.B1(_03926_),
    .Y(_00966_),
    .A1(net31),
    .A2(_03920_));
 sg13g2_a21oi_1 _21459_ (.A1(net632),
    .A2(net649),
    .Y(_03927_),
    .B1(_03909_));
 sg13g2_nor2_2 _21460_ (.A(net530),
    .B(_11496_),
    .Y(_03928_));
 sg13g2_nor2_1 _21461_ (.A(_10514_),
    .B(_10518_),
    .Y(_03929_));
 sg13g2_nand2_2 _21462_ (.Y(_03930_),
    .A(_03904_),
    .B(_03929_));
 sg13g2_and2_1 _21463_ (.A(_03928_),
    .B(_03930_),
    .X(_03931_));
 sg13g2_nor2_1 _21464_ (.A(_03914_),
    .B(net279),
    .Y(_03932_));
 sg13g2_o21ai_1 _21465_ (.B1(_03916_),
    .Y(_03933_),
    .A1(_03932_),
    .A2(_03919_));
 sg13g2_xnor2_1 _21466_ (.Y(_03934_),
    .A(net237),
    .B(_03933_));
 sg13g2_a221oi_1 _21467_ (.B2(_03934_),
    .C1(_11645_),
    .B1(net28),
    .A1(\cpu.dec.div ),
    .Y(_03935_),
    .A2(_11913_));
 sg13g2_inv_1 _21468_ (.Y(_03936_),
    .A(net1105));
 sg13g2_o21ai_1 _21469_ (.B1(_03936_),
    .Y(_03937_),
    .A1(_03931_),
    .A2(_03935_));
 sg13g2_nand2_1 _21470_ (.Y(_03938_),
    .A(net1105),
    .B(_03928_));
 sg13g2_o21ai_1 _21471_ (.B1(_03927_),
    .Y(_03939_),
    .A1(_03930_),
    .A2(_03938_));
 sg13g2_and4_1 _21472_ (.A(net1105),
    .B(net28),
    .C(net85),
    .D(_03934_),
    .X(_03940_));
 sg13g2_nor2_1 _21473_ (.A(_03939_),
    .B(_03940_),
    .Y(_03941_));
 sg13g2_nor2_1 _21474_ (.A(\cpu.ex.r_mult[19] ),
    .B(_03907_),
    .Y(_03942_));
 sg13g2_a221oi_1 _21475_ (.B2(_03941_),
    .C1(_03942_),
    .B1(_03937_),
    .A1(net535),
    .Y(_00967_),
    .A2(_03927_));
 sg13g2_xnor2_1 _21476_ (.Y(_03943_),
    .A(net287),
    .B(_11126_));
 sg13g2_nor2_1 _21477_ (.A(net27),
    .B(_03943_),
    .Y(_03944_));
 sg13g2_xnor2_1 _21478_ (.Y(_03945_),
    .A(_11329_),
    .B(_03944_));
 sg13g2_nor2_1 _21479_ (.A(_11328_),
    .B(net530),
    .Y(_03946_));
 sg13g2_nor2_1 _21480_ (.A(net1105),
    .B(_03930_),
    .Y(_03947_));
 sg13g2_mux2_1 _21481_ (.A0(_03946_),
    .A1(_11328_),
    .S(_03947_),
    .X(_03948_));
 sg13g2_nand2b_1 _21482_ (.Y(_03949_),
    .B(net363),
    .A_N(\cpu.ex.r_mult[20] ));
 sg13g2_a21o_1 _21483_ (.A2(net585),
    .A1(net595),
    .B1(net364),
    .X(_03950_));
 sg13g2_a22oi_1 _21484_ (.Y(_03951_),
    .B1(_03949_),
    .B2(_03950_),
    .A2(_03948_),
    .A1(_11605_));
 sg13g2_o21ai_1 _21485_ (.B1(_03951_),
    .Y(_00968_),
    .A1(net31),
    .A2(_03945_));
 sg13g2_nand2_1 _21486_ (.Y(_03952_),
    .A(_11119_),
    .B(_11125_));
 sg13g2_a21oi_1 _21487_ (.A1(_03952_),
    .A2(_11334_),
    .Y(_03953_),
    .B1(_11383_));
 sg13g2_xnor2_1 _21488_ (.Y(_03954_),
    .A(net168),
    .B(_03953_));
 sg13g2_nor2_1 _21489_ (.A(net27),
    .B(_03954_),
    .Y(_03955_));
 sg13g2_xnor2_1 _21490_ (.Y(_03956_),
    .A(_11363_),
    .B(_03955_));
 sg13g2_nand2b_1 _21491_ (.Y(_03957_),
    .B(net363),
    .A_N(\cpu.ex.r_mult[21] ));
 sg13g2_a21o_1 _21492_ (.A2(net585),
    .A1(net651),
    .B1(net364),
    .X(_03958_));
 sg13g2_or3_1 _21493_ (.A(_11328_),
    .B(net1105),
    .C(_03930_),
    .X(_03959_));
 sg13g2_xor2_1 _21494_ (.B(_03959_),
    .A(_11362_),
    .X(_03960_));
 sg13g2_a22oi_1 _21495_ (.Y(_03961_),
    .B1(_03960_),
    .B2(net332),
    .A2(_03958_),
    .A1(_03957_));
 sg13g2_o21ai_1 _21496_ (.B1(_03961_),
    .Y(_00969_),
    .A1(net31),
    .A2(_03956_));
 sg13g2_nand2_1 _21497_ (.Y(_03962_),
    .A(net168),
    .B(_03953_));
 sg13g2_nor2_1 _21498_ (.A(net168),
    .B(_03953_),
    .Y(_03963_));
 sg13g2_a21oi_1 _21499_ (.A1(_11363_),
    .A2(_03962_),
    .Y(_03964_),
    .B1(_03963_));
 sg13g2_xnor2_1 _21500_ (.Y(_03965_),
    .A(net194),
    .B(_03964_));
 sg13g2_nor2_1 _21501_ (.A(net27),
    .B(_03965_),
    .Y(_03966_));
 sg13g2_xnor2_1 _21502_ (.Y(_03967_),
    .A(_11389_),
    .B(_03966_));
 sg13g2_nor3_1 _21503_ (.A(_11362_),
    .B(_11328_),
    .C(net1105),
    .Y(_03968_));
 sg13g2_nor2b_1 _21504_ (.A(_03930_),
    .B_N(_03968_),
    .Y(_03969_));
 sg13g2_xnor2_1 _21505_ (.Y(_03970_),
    .A(net1101),
    .B(_03969_));
 sg13g2_a21oi_1 _21506_ (.A1(net1028),
    .A2(net649),
    .Y(_03971_),
    .B1(_03909_));
 sg13g2_a21oi_1 _21507_ (.A1(_11265_),
    .A2(_03890_),
    .Y(_03972_),
    .B1(_03971_));
 sg13g2_a21oi_1 _21508_ (.A1(net332),
    .A2(_03970_),
    .Y(_03973_),
    .B1(_03972_));
 sg13g2_o21ai_1 _21509_ (.B1(_03973_),
    .Y(_00970_),
    .A1(net31),
    .A2(_03967_));
 sg13g2_nand2_1 _21510_ (.Y(_03974_),
    .A(net1101),
    .B(net194));
 sg13g2_nand3_1 _21511_ (.B(_11334_),
    .C(_03974_),
    .A(_11675_),
    .Y(_03975_));
 sg13g2_nand3b_1 _21512_ (.B(_11334_),
    .C(_03974_),
    .Y(_03976_),
    .A_N(_11362_));
 sg13g2_a22oi_1 _21513_ (.Y(_03977_),
    .B1(_03975_),
    .B2(_03976_),
    .A2(_11125_),
    .A1(_11119_));
 sg13g2_nor2_1 _21514_ (.A(_11362_),
    .B(net168),
    .Y(_03978_));
 sg13g2_a221oi_1 _21515_ (.B2(_11362_),
    .C1(_11330_),
    .B1(net168),
    .A1(_11232_),
    .Y(_03979_),
    .A2(net194));
 sg13g2_a21oi_1 _21516_ (.A1(_03974_),
    .A2(_03978_),
    .Y(_03980_),
    .B1(_03979_));
 sg13g2_inv_1 _21517_ (.Y(_03981_),
    .A(_03980_));
 sg13g2_nor2_1 _21518_ (.A(_11232_),
    .B(net194),
    .Y(_03982_));
 sg13g2_nor3_2 _21519_ (.A(_03977_),
    .B(_03981_),
    .C(_03982_),
    .Y(_03983_));
 sg13g2_nand2_1 _21520_ (.Y(_03984_),
    .A(_11118_),
    .B(_10507_));
 sg13g2_nand3_1 _21521_ (.B(_11327_),
    .C(_11675_),
    .A(net193),
    .Y(_03985_));
 sg13g2_o21ai_1 _21522_ (.B1(net628),
    .Y(_03986_),
    .A1(_03984_),
    .A2(_03985_));
 sg13g2_buf_1 _21523_ (.A(_03986_),
    .X(_03987_));
 sg13g2_inv_1 _21524_ (.Y(_03988_),
    .A(_03987_));
 sg13g2_nor3_1 _21525_ (.A(net239),
    .B(_03983_),
    .C(_03988_),
    .Y(_03989_));
 sg13g2_o21ai_1 _21526_ (.B1(net239),
    .Y(_03990_),
    .A1(_03983_),
    .A2(_03988_));
 sg13g2_nor2b_1 _21527_ (.A(_03989_),
    .B_N(_03990_),
    .Y(_03991_));
 sg13g2_nand2_1 _21528_ (.Y(_03992_),
    .A(net28),
    .B(_03991_));
 sg13g2_xnor2_1 _21529_ (.Y(_03993_),
    .A(_11380_),
    .B(_03992_));
 sg13g2_nand2b_1 _21530_ (.Y(_03994_),
    .B(net363),
    .A_N(\cpu.ex.r_mult[23] ));
 sg13g2_a21o_1 _21531_ (.A2(net585),
    .A1(net1042),
    .B1(net364),
    .X(_03995_));
 sg13g2_nor3_1 _21532_ (.A(net1101),
    .B(_10514_),
    .C(_10518_),
    .Y(_03996_));
 sg13g2_nand4_1 _21533_ (.B(net606),
    .C(_03968_),
    .A(_11861_),
    .Y(_03997_),
    .D(_03996_));
 sg13g2_nor2_1 _21534_ (.A(_03884_),
    .B(_03997_),
    .Y(_03998_));
 sg13g2_xnor2_1 _21535_ (.Y(_03999_),
    .A(_11265_),
    .B(_03998_));
 sg13g2_a22oi_1 _21536_ (.Y(_04000_),
    .B1(_03999_),
    .B2(net332),
    .A2(_03995_),
    .A1(_03994_));
 sg13g2_o21ai_1 _21537_ (.B1(_04000_),
    .Y(_00971_),
    .A1(net31),
    .A2(_03993_));
 sg13g2_inv_1 _21538_ (.Y(_04001_),
    .A(\cpu.ex.r_mult[24] ));
 sg13g2_inv_2 _21539_ (.Y(_04002_),
    .A(net1102));
 sg13g2_nor2b_1 _21540_ (.A(net1101),
    .B_N(_03968_),
    .Y(_04003_));
 sg13g2_nand4_1 _21541_ (.B(_03904_),
    .C(_03929_),
    .A(net1003),
    .Y(_04004_),
    .D(_04003_));
 sg13g2_xnor2_1 _21542_ (.Y(_04005_),
    .A(_04002_),
    .B(_04004_));
 sg13g2_a221oi_1 _21543_ (.B2(_04005_),
    .C1(_03909_),
    .B1(_03903_),
    .A1(net1043),
    .Y(_04006_),
    .A2(net649));
 sg13g2_and3_1 _21544_ (.X(_04007_),
    .A(_11304_),
    .B(_11335_),
    .C(_11364_));
 sg13g2_a21oi_1 _21545_ (.A1(_03952_),
    .A2(_04007_),
    .Y(_04008_),
    .B1(_11396_));
 sg13g2_xnor2_1 _21546_ (.Y(_04009_),
    .A(net189),
    .B(_04008_));
 sg13g2_nor2_1 _21547_ (.A(net27),
    .B(_04009_),
    .Y(_04010_));
 sg13g2_xnor2_1 _21548_ (.Y(_04011_),
    .A(_11160_),
    .B(_04010_));
 sg13g2_and2_1 _21549_ (.A(_03897_),
    .B(_04006_),
    .X(_04012_));
 sg13g2_a221oi_1 _21550_ (.B2(_04011_),
    .C1(_04012_),
    .B1(_04006_),
    .A1(_04001_),
    .Y(_00972_),
    .A2(net363));
 sg13g2_nand2_1 _21551_ (.Y(_04013_),
    .A(net1102),
    .B(net189));
 sg13g2_and3_1 _21552_ (.X(_04014_),
    .A(net1003),
    .B(net661),
    .C(_04013_));
 sg13g2_nand3_1 _21553_ (.B(net216),
    .C(_03987_),
    .A(_04002_),
    .Y(_04015_));
 sg13g2_nand2_1 _21554_ (.Y(_04016_),
    .A(_04002_),
    .B(net190));
 sg13g2_o21ai_1 _21555_ (.B1(_04016_),
    .Y(_04017_),
    .A1(_03983_),
    .A2(_04015_));
 sg13g2_nor4_1 _21556_ (.A(net189),
    .B(net239),
    .C(_03983_),
    .D(_03988_),
    .Y(_04018_));
 sg13g2_a221oi_1 _21557_ (.B2(net661),
    .C1(_04018_),
    .B1(_04017_),
    .A1(_03990_),
    .Y(_04019_),
    .A2(_04014_));
 sg13g2_xnor2_1 _21558_ (.Y(_04020_),
    .A(net215),
    .B(_04019_));
 sg13g2_nor2_1 _21559_ (.A(net27),
    .B(_04020_),
    .Y(_04021_));
 sg13g2_xnor2_1 _21560_ (.Y(_04022_),
    .A(_11229_),
    .B(_04021_));
 sg13g2_nand2b_1 _21561_ (.Y(_04023_),
    .B(net363),
    .A_N(\cpu.ex.r_mult[25] ));
 sg13g2_a21o_1 _21562_ (.A2(net585),
    .A1(_11085_),
    .B1(net364),
    .X(_04024_));
 sg13g2_nand3_1 _21563_ (.B(_04002_),
    .C(_03998_),
    .A(net1003),
    .Y(_04025_));
 sg13g2_nor3_1 _21564_ (.A(_11228_),
    .B(net1102),
    .C(_04004_),
    .Y(_04026_));
 sg13g2_a21oi_1 _21565_ (.A1(_11228_),
    .A2(_04025_),
    .Y(_04027_),
    .B1(_04026_));
 sg13g2_a22oi_1 _21566_ (.Y(_04028_),
    .B1(_04027_),
    .B2(net332),
    .A2(_04024_),
    .A1(_04023_));
 sg13g2_o21ai_1 _21567_ (.B1(_04028_),
    .Y(_00973_),
    .A1(net31),
    .A2(_04022_));
 sg13g2_xnor2_1 _21568_ (.Y(_04029_),
    .A(_11164_),
    .B(_04026_));
 sg13g2_inv_2 _21569_ (.Y(_04030_),
    .A(net1106));
 sg13g2_a21oi_1 _21570_ (.A1(net1104),
    .A2(_03887_),
    .Y(_04031_),
    .B1(_03909_));
 sg13g2_a21oi_1 _21571_ (.A1(_04030_),
    .A2(_03890_),
    .Y(_04032_),
    .B1(_04031_));
 sg13g2_a21oi_1 _21572_ (.A1(_03903_),
    .A2(_04029_),
    .Y(_04033_),
    .B1(_04032_));
 sg13g2_nand3_1 _21573_ (.B(net190),
    .C(_03989_),
    .A(net217),
    .Y(_04034_));
 sg13g2_nand2_1 _21574_ (.Y(_04035_),
    .A(_11367_),
    .B(net217));
 sg13g2_nor2_1 _21575_ (.A(_11159_),
    .B(net189),
    .Y(_04036_));
 sg13g2_nor3_1 _21576_ (.A(_04036_),
    .B(net216),
    .C(_03982_),
    .Y(_04037_));
 sg13g2_nor3_1 _21577_ (.A(net1003),
    .B(_04036_),
    .C(_03982_),
    .Y(_04038_));
 sg13g2_nor2_1 _21578_ (.A(_03977_),
    .B(_03981_),
    .Y(_04039_));
 sg13g2_o21ai_1 _21579_ (.B1(_04039_),
    .Y(_04040_),
    .A1(_04037_),
    .A2(_04038_));
 sg13g2_a221oi_1 _21580_ (.B2(_11264_),
    .C1(_03987_),
    .B1(net216),
    .A1(_04002_),
    .Y(_04041_),
    .A2(net190));
 sg13g2_nor3_1 _21581_ (.A(_11264_),
    .B(_04036_),
    .C(net216),
    .Y(_04042_));
 sg13g2_nor2_1 _21582_ (.A(_04041_),
    .B(_04042_),
    .Y(_04043_));
 sg13g2_and3_1 _21583_ (.X(_04044_),
    .A(_04013_),
    .B(_04040_),
    .C(_04043_));
 sg13g2_o21ai_1 _21584_ (.B1(_04044_),
    .Y(_04045_),
    .A1(_11367_),
    .A2(net217));
 sg13g2_a22oi_1 _21585_ (.Y(_04046_),
    .B1(_04035_),
    .B2(_04045_),
    .A2(_04034_),
    .A1(_09379_));
 sg13g2_nor4_1 _21586_ (.A(net188),
    .B(_11194_),
    .C(_03872_),
    .D(net31),
    .Y(_04047_));
 sg13g2_nand2b_1 _21587_ (.Y(_04048_),
    .B(_04047_),
    .A_N(_04046_));
 sg13g2_nand3_1 _21588_ (.B(_11194_),
    .C(net58),
    .A(net188),
    .Y(_04049_));
 sg13g2_or4_1 _21589_ (.A(net214),
    .B(_11194_),
    .C(_03871_),
    .D(_03896_),
    .X(_04050_));
 sg13g2_mux2_1 _21590_ (.A0(_04049_),
    .A1(_04050_),
    .S(_04046_),
    .X(_04051_));
 sg13g2_nor4_1 _21591_ (.A(_11164_),
    .B(net628),
    .C(net188),
    .D(_03896_),
    .Y(_04052_));
 sg13g2_nor3_1 _21592_ (.A(_11164_),
    .B(net628),
    .C(_03896_),
    .Y(_04053_));
 sg13g2_a22oi_1 _21593_ (.Y(_04054_),
    .B1(_04053_),
    .B2(_03872_),
    .A2(_04052_),
    .A1(_04046_));
 sg13g2_nand4_1 _21594_ (.B(_04048_),
    .C(_04051_),
    .A(_04033_),
    .Y(_00974_),
    .D(_04054_));
 sg13g2_nand2_1 _21595_ (.Y(_04055_),
    .A(_11367_),
    .B(_04002_));
 sg13g2_nand2b_1 _21596_ (.Y(_04056_),
    .B(net1003),
    .A_N(_11164_));
 sg13g2_nor4_2 _21597_ (.A(_03884_),
    .B(_03997_),
    .C(_04055_),
    .Y(_04057_),
    .D(_04056_));
 sg13g2_xnor2_1 _21598_ (.Y(_04058_),
    .A(_04030_),
    .B(_04057_));
 sg13g2_a221oi_1 _21599_ (.B2(_04058_),
    .C1(_03910_),
    .B1(net332),
    .A1(net1107),
    .Y(_04059_),
    .A2(net585));
 sg13g2_xnor2_1 _21600_ (.Y(_04060_),
    .A(net212),
    .B(_11399_));
 sg13g2_a21oi_1 _21601_ (.A1(net28),
    .A2(_04060_),
    .Y(_04061_),
    .B1(_11412_));
 sg13g2_and3_1 _21602_ (.X(_04062_),
    .A(_11412_),
    .B(net28),
    .C(_04060_));
 sg13g2_o21ai_1 _21603_ (.B1(net58),
    .Y(_04063_),
    .A1(_04061_),
    .A2(_04062_));
 sg13g2_a22oi_1 _21604_ (.Y(_00975_),
    .B1(_04059_),
    .B2(_04063_),
    .A2(net363),
    .A1(_10402_));
 sg13g2_nand2_1 _21605_ (.Y(_04064_),
    .A(net1106),
    .B(_04057_));
 sg13g2_xnor2_1 _21606_ (.Y(_04065_),
    .A(_10384_),
    .B(_04064_));
 sg13g2_a221oi_1 _21607_ (.B2(_04065_),
    .C1(_03909_),
    .B1(_03902_),
    .A1(net620),
    .Y(_04066_),
    .A2(net649));
 sg13g2_nor2_1 _21608_ (.A(net211),
    .B(_11399_),
    .Y(_04067_));
 sg13g2_nand2_1 _21609_ (.Y(_04068_),
    .A(net211),
    .B(_11399_));
 sg13g2_o21ai_1 _21610_ (.B1(_04068_),
    .Y(_04069_),
    .A1(_11412_),
    .A2(_04067_));
 sg13g2_xnor2_1 _21611_ (.Y(_04070_),
    .A(net213),
    .B(_04069_));
 sg13g2_nor2_1 _21612_ (.A(_03871_),
    .B(_04070_),
    .Y(_04071_));
 sg13g2_nor2_1 _21613_ (.A(_10331_),
    .B(net628),
    .Y(_04072_));
 sg13g2_xnor2_1 _21614_ (.Y(_04073_),
    .A(_04071_),
    .B(_04072_));
 sg13g2_and2_1 _21615_ (.A(_03897_),
    .B(_04066_),
    .X(_04074_));
 sg13g2_a221oi_1 _21616_ (.B2(_04073_),
    .C1(_04074_),
    .B1(_04066_),
    .A1(_11402_),
    .Y(_00976_),
    .A2(_03921_));
 sg13g2_a21oi_1 _21617_ (.A1(net614),
    .A2(net649),
    .Y(_04075_),
    .B1(_03909_));
 sg13g2_a22oi_1 _21618_ (.Y(_04076_),
    .B1(_04075_),
    .B2(net535),
    .A2(net363),
    .A1(_11443_));
 sg13g2_nor4_1 _21619_ (.A(net1011),
    .B(net141),
    .C(_10421_),
    .D(_03871_),
    .Y(_04077_));
 sg13g2_nand2_1 _21620_ (.Y(_04078_),
    .A(net1106),
    .B(net212));
 sg13g2_nand2b_1 _21621_ (.Y(_04079_),
    .B(_11401_),
    .A_N(_04078_));
 sg13g2_nand4_1 _21622_ (.B(_10384_),
    .C(_10383_),
    .A(_04030_),
    .Y(_04080_),
    .D(net211));
 sg13g2_a21oi_1 _21623_ (.A1(_04079_),
    .A2(_04080_),
    .Y(_04081_),
    .B1(net628));
 sg13g2_a21oi_1 _21624_ (.A1(_04030_),
    .A2(_10331_),
    .Y(_04082_),
    .B1(net628));
 sg13g2_nor2_1 _21625_ (.A(_11488_),
    .B(_04082_),
    .Y(_04083_));
 sg13g2_o21ai_1 _21626_ (.B1(_11399_),
    .Y(_04084_),
    .A1(_04081_),
    .A2(_04083_));
 sg13g2_buf_1 _21627_ (.A(_04084_),
    .X(_04085_));
 sg13g2_nand2b_1 _21628_ (.Y(_04086_),
    .B(_04085_),
    .A_N(_10425_));
 sg13g2_nand2_1 _21629_ (.Y(_04087_),
    .A(net1011),
    .B(net661));
 sg13g2_a21oi_1 _21630_ (.A1(_11481_),
    .A2(_04086_),
    .Y(_04088_),
    .B1(_04087_));
 sg13g2_o21ai_1 _21631_ (.B1(net661),
    .Y(_04089_),
    .A1(net1011),
    .A2(_10422_));
 sg13g2_and4_1 _21632_ (.A(net141),
    .B(_11480_),
    .C(_04085_),
    .D(_04089_),
    .X(_04090_));
 sg13g2_nor2_1 _21633_ (.A(net141),
    .B(_11645_),
    .Y(_04091_));
 sg13g2_nand3b_1 _21634_ (.B(_04087_),
    .C(_04091_),
    .Y(_04092_),
    .A_N(_04085_));
 sg13g2_nand4_1 _21635_ (.B(net661),
    .C(net141),
    .A(net1011),
    .Y(_04093_),
    .D(net85));
 sg13g2_a21oi_1 _21636_ (.A1(_10421_),
    .A2(_04085_),
    .Y(_04094_),
    .B1(_04093_));
 sg13g2_nor4_1 _21637_ (.A(_11402_),
    .B(net530),
    .C(_11496_),
    .D(_04057_),
    .Y(_04095_));
 sg13g2_nor3_1 _21638_ (.A(_04030_),
    .B(net1011),
    .C(_10331_),
    .Y(_04096_));
 sg13g2_and3_1 _21639_ (.X(_04097_),
    .A(_03928_),
    .B(_04057_),
    .C(_04096_));
 sg13g2_nand2_1 _21640_ (.Y(_04098_),
    .A(net1106),
    .B(_10384_));
 sg13g2_nand3_1 _21641_ (.B(_03928_),
    .C(_04098_),
    .A(net1011),
    .Y(_04099_));
 sg13g2_nand2_1 _21642_ (.Y(_04100_),
    .A(_04075_),
    .B(_04099_));
 sg13g2_nor4_1 _21643_ (.A(_04094_),
    .B(_04095_),
    .C(_04097_),
    .D(_04100_),
    .Y(_04101_));
 sg13g2_o21ai_1 _21644_ (.B1(_04101_),
    .Y(_04102_),
    .A1(_03871_),
    .A2(_04092_));
 sg13g2_or4_1 _21645_ (.A(_04077_),
    .B(_04088_),
    .C(_04090_),
    .D(_04102_),
    .X(_04103_));
 sg13g2_nand2_1 _21646_ (.Y(_04104_),
    .A(_11645_),
    .B(_04101_));
 sg13g2_and3_1 _21647_ (.X(_00977_),
    .A(_04076_),
    .B(_04103_),
    .C(_04104_));
 sg13g2_a21oi_1 _21648_ (.A1(net605),
    .A2(net585),
    .Y(_04105_),
    .B1(net364));
 sg13g2_nand2_1 _21649_ (.Y(_04106_),
    .A(_10430_),
    .B(_11415_));
 sg13g2_xnor2_1 _21650_ (.Y(_04107_),
    .A(_04106_),
    .B(net192));
 sg13g2_nand2_1 _21651_ (.Y(_04108_),
    .A(_10269_),
    .B(net661));
 sg13g2_a21oi_1 _21652_ (.A1(net28),
    .A2(_04107_),
    .Y(_04109_),
    .B1(_04108_));
 sg13g2_and3_1 _21653_ (.X(_04110_),
    .A(net28),
    .B(_04107_),
    .C(_04108_));
 sg13g2_o21ai_1 _21654_ (.B1(net85),
    .Y(_04111_),
    .A1(_04109_),
    .A2(_04110_));
 sg13g2_nor3_1 _21655_ (.A(_11402_),
    .B(_10331_),
    .C(_04064_),
    .Y(_04112_));
 sg13g2_xnor2_1 _21656_ (.Y(_04113_),
    .A(_11443_),
    .B(_04112_));
 sg13g2_a221oi_1 _21657_ (.B2(_04113_),
    .C1(_03910_),
    .B1(_03928_),
    .A1(net605),
    .Y(_04114_),
    .A2(_03888_));
 sg13g2_nor3_1 _21658_ (.A(\cpu.ex.r_mult[30] ),
    .B(net535),
    .C(_11517_),
    .Y(_04115_));
 sg13g2_a221oi_1 _21659_ (.B2(_04114_),
    .C1(_04115_),
    .B1(_04111_),
    .A1(net535),
    .Y(_00978_),
    .A2(_04105_));
 sg13g2_nand2_1 _21660_ (.Y(_04116_),
    .A(_10269_),
    .B(_04112_));
 sg13g2_xor2_1 _21661_ (.B(_04116_),
    .A(_00297_),
    .X(_04117_));
 sg13g2_inv_1 _21662_ (.Y(_04118_),
    .A(\cpu.ex.r_mult[31] ));
 sg13g2_o21ai_1 _21663_ (.B1(_11416_),
    .Y(_04119_),
    .A1(_10418_),
    .A2(_10269_));
 sg13g2_nand2_1 _21664_ (.Y(_04120_),
    .A(net211),
    .B(_04119_));
 sg13g2_xnor2_1 _21665_ (.Y(_04121_),
    .A(_11443_),
    .B(net192));
 sg13g2_nand4_1 _21666_ (.B(_10269_),
    .C(net211),
    .A(_04030_),
    .Y(_04122_),
    .D(net192));
 sg13g2_o21ai_1 _21667_ (.B1(_04122_),
    .Y(_04123_),
    .A1(_04078_),
    .A2(_04121_));
 sg13g2_nand2_1 _21668_ (.Y(_04124_),
    .A(_11416_),
    .B(_04123_));
 sg13g2_o21ai_1 _21669_ (.B1(_04124_),
    .Y(_04125_),
    .A1(net192),
    .A2(_04120_));
 sg13g2_nand3_1 _21670_ (.B(_11408_),
    .C(_04125_),
    .A(_11399_),
    .Y(_04126_));
 sg13g2_nand2_1 _21671_ (.Y(_04127_),
    .A(_10430_),
    .B(net192));
 sg13g2_o21ai_1 _21672_ (.B1(_04108_),
    .Y(_04128_),
    .A1(_10430_),
    .A2(net192));
 sg13g2_nand2_1 _21673_ (.Y(_04129_),
    .A(_04127_),
    .B(_04128_));
 sg13g2_a21oi_1 _21674_ (.A1(_04126_),
    .A2(_04129_),
    .Y(_04130_),
    .B1(net169));
 sg13g2_nor2_1 _21675_ (.A(_11471_),
    .B(_03896_),
    .Y(_04131_));
 sg13g2_o21ai_1 _21676_ (.B1(_04131_),
    .Y(_04132_),
    .A1(net27),
    .A2(_04130_));
 sg13g2_a21oi_1 _21677_ (.A1(net860),
    .A2(_03888_),
    .Y(_04133_),
    .B1(net364));
 sg13g2_a22oi_1 _21678_ (.Y(_04134_),
    .B1(_04132_),
    .B2(_04133_),
    .A2(_03921_),
    .A1(_04118_));
 sg13g2_a21o_1 _21679_ (.A2(_04117_),
    .A1(net332),
    .B1(_04134_),
    .X(_00979_));
 sg13g2_nor2_1 _21680_ (.A(_09276_),
    .B(_11524_),
    .Y(_04135_));
 sg13g2_mux2_1 _21681_ (.A0(_04135_),
    .A1(_08576_),
    .S(_11910_),
    .X(_04136_));
 sg13g2_nor2_1 _21682_ (.A(_08615_),
    .B(_10743_),
    .Y(_04137_));
 sg13g2_buf_1 _21683_ (.A(_04137_),
    .X(_04138_));
 sg13g2_nand3_1 _21684_ (.B(_04136_),
    .C(net226),
    .A(net658),
    .Y(_04139_));
 sg13g2_buf_2 _21685_ (.A(_04139_),
    .X(_04140_));
 sg13g2_buf_1 _21686_ (.A(_04140_),
    .X(_04141_));
 sg13g2_or2_1 _21687_ (.X(_04142_),
    .B(_11533_),
    .A(_11516_));
 sg13g2_buf_2 _21688_ (.A(_04142_),
    .X(_04143_));
 sg13g2_and2_1 _21689_ (.A(_08255_),
    .B(_03642_),
    .X(_04144_));
 sg13g2_buf_2 _21690_ (.A(_04144_),
    .X(_04145_));
 sg13g2_a21o_1 _21691_ (.A2(_11599_),
    .A1(_11019_),
    .B1(_11487_),
    .X(_04146_));
 sg13g2_and2_1 _21692_ (.A(_11019_),
    .B(_10507_),
    .X(_04147_));
 sg13g2_buf_2 _21693_ (.A(_04147_),
    .X(_04148_));
 sg13g2_buf_1 _21694_ (.A(_04148_),
    .X(_04149_));
 sg13g2_nor4_1 _21695_ (.A(net286),
    .B(net238),
    .C(net240),
    .D(net279),
    .Y(_04150_));
 sg13g2_buf_1 _21696_ (.A(_04150_),
    .X(_04151_));
 sg13g2_buf_1 _21697_ (.A(_04151_),
    .X(_04152_));
 sg13g2_a21o_1 _21698_ (.A2(net162),
    .A1(_03801_),
    .B1(net161),
    .X(_04153_));
 sg13g2_a21oi_1 _21699_ (.A1(_04145_),
    .A2(_04146_),
    .Y(_04154_),
    .B1(_04153_));
 sg13g2_buf_1 _21700_ (.A(_03826_),
    .X(_04155_));
 sg13g2_a21oi_2 _21701_ (.B1(_11562_),
    .Y(_04156_),
    .A2(_10470_),
    .A1(_10464_));
 sg13g2_and2_1 _21702_ (.A(_11019_),
    .B(_04156_),
    .X(_04157_));
 sg13g2_buf_1 _21703_ (.A(_04157_),
    .X(_04158_));
 sg13g2_buf_1 _21704_ (.A(net199),
    .X(_04159_));
 sg13g2_nor4_1 _21705_ (.A(net286),
    .B(net238),
    .C(net240),
    .D(net285),
    .Y(_04160_));
 sg13g2_buf_1 _21706_ (.A(_04160_),
    .X(_04161_));
 sg13g2_buf_1 _21707_ (.A(net181),
    .X(_04162_));
 sg13g2_buf_1 _21708_ (.A(_03657_),
    .X(_04163_));
 sg13g2_a22oi_1 _21709_ (.Y(_04164_),
    .B1(net160),
    .B2(net134),
    .A2(net182),
    .A1(net135));
 sg13g2_nand2_1 _21710_ (.Y(_04165_),
    .A(_10520_),
    .B(net873));
 sg13g2_o21ai_1 _21711_ (.B1(_04165_),
    .Y(_04166_),
    .A1(_10409_),
    .A2(_10522_));
 sg13g2_a21oi_1 _21712_ (.A1(_10537_),
    .A2(_10545_),
    .Y(_04167_),
    .B1(_10546_));
 sg13g2_o21ai_1 _21713_ (.B1(net750),
    .Y(_04168_),
    .A1(_04166_),
    .A2(_04167_));
 sg13g2_nand2_1 _21714_ (.Y(_04169_),
    .A(net1072),
    .B(net876));
 sg13g2_a22oi_1 _21715_ (.Y(_04170_),
    .B1(_04168_),
    .B2(_04169_),
    .A2(_11017_),
    .A1(_11016_));
 sg13g2_buf_1 _21716_ (.A(_04170_),
    .X(_04171_));
 sg13g2_and2_1 _21717_ (.A(_04156_),
    .B(_04171_),
    .X(_04172_));
 sg13g2_buf_1 _21718_ (.A(_04172_),
    .X(_04173_));
 sg13g2_buf_1 _21719_ (.A(_04173_),
    .X(_04174_));
 sg13g2_buf_1 _21720_ (.A(net180),
    .X(_04175_));
 sg13g2_nor4_1 _21721_ (.A(net286),
    .B(net238),
    .C(_11594_),
    .D(net279),
    .Y(_04176_));
 sg13g2_buf_2 _21722_ (.A(_04176_),
    .X(_04177_));
 sg13g2_nand2_1 _21723_ (.Y(_04178_),
    .A(_03730_),
    .B(_03731_));
 sg13g2_buf_1 _21724_ (.A(_04178_),
    .X(_04179_));
 sg13g2_buf_1 _21725_ (.A(_04179_),
    .X(_04180_));
 sg13g2_a22oi_1 _21726_ (.Y(_04181_),
    .B1(_04177_),
    .B2(net133),
    .A2(net159),
    .A1(net163));
 sg13g2_and2_1 _21727_ (.A(_11599_),
    .B(_04171_),
    .X(_04182_));
 sg13g2_buf_1 _21728_ (.A(_04182_),
    .X(_04183_));
 sg13g2_nor3_1 _21729_ (.A(_10510_),
    .B(_10512_),
    .C(net279),
    .Y(_04184_));
 sg13g2_and2_1 _21730_ (.A(_11485_),
    .B(_04184_),
    .X(_04185_));
 sg13g2_buf_2 _21731_ (.A(_04185_),
    .X(_04186_));
 sg13g2_buf_1 _21732_ (.A(_03711_),
    .X(_04187_));
 sg13g2_a22oi_1 _21733_ (.Y(_04188_),
    .B1(_04186_),
    .B2(net132),
    .A2(_04183_),
    .A1(net138));
 sg13g2_buf_1 _21734_ (.A(_03668_),
    .X(_04189_));
 sg13g2_and2_1 _21735_ (.A(_11485_),
    .B(_04156_),
    .X(_04190_));
 sg13g2_buf_1 _21736_ (.A(_04190_),
    .X(_04191_));
 sg13g2_buf_1 _21737_ (.A(_04191_),
    .X(_04192_));
 sg13g2_and2_1 _21738_ (.A(_04171_),
    .B(_04184_),
    .X(_04193_));
 sg13g2_buf_1 _21739_ (.A(_04193_),
    .X(_04194_));
 sg13g2_buf_1 _21740_ (.A(_04194_),
    .X(_04195_));
 sg13g2_buf_1 _21741_ (.A(_03742_),
    .X(_04196_));
 sg13g2_a22oi_1 _21742_ (.Y(_04197_),
    .B1(net158),
    .B2(net130),
    .A2(net179),
    .A1(net131));
 sg13g2_and2_1 _21743_ (.A(_11019_),
    .B(_04184_),
    .X(_04198_));
 sg13g2_buf_1 _21744_ (.A(_04198_),
    .X(_04199_));
 sg13g2_buf_1 _21745_ (.A(_04199_),
    .X(_04200_));
 sg13g2_and2_1 _21746_ (.A(_11485_),
    .B(_11599_),
    .X(_04201_));
 sg13g2_buf_2 _21747_ (.A(_04201_),
    .X(_04202_));
 sg13g2_a22oi_1 _21748_ (.Y(_04203_),
    .B1(_04202_),
    .B2(net164),
    .A2(net157),
    .A1(net165));
 sg13g2_nor4_1 _21749_ (.A(_11509_),
    .B(_11550_),
    .C(net237),
    .D(_11562_),
    .Y(_04204_));
 sg13g2_buf_2 _21750_ (.A(_04204_),
    .X(_04205_));
 sg13g2_and2_1 _21751_ (.A(_10507_),
    .B(_04171_),
    .X(_04206_));
 sg13g2_buf_1 _21752_ (.A(_04206_),
    .X(_04207_));
 sg13g2_buf_1 _21753_ (.A(_04207_),
    .X(_04208_));
 sg13g2_a22oi_1 _21754_ (.Y(_04209_),
    .B1(net156),
    .B2(net167),
    .A2(_04205_),
    .A1(net166));
 sg13g2_and4_1 _21755_ (.A(_04188_),
    .B(_04197_),
    .C(_04203_),
    .D(_04209_),
    .X(_04210_));
 sg13g2_nand4_1 _21756_ (.B(_04164_),
    .C(_04181_),
    .A(_04154_),
    .Y(_04211_),
    .D(_04210_));
 sg13g2_or2_1 _21757_ (.X(_04212_),
    .B(net1116),
    .A(_08255_));
 sg13g2_buf_2 _21758_ (.A(_04212_),
    .X(_04213_));
 sg13g2_buf_1 _21759_ (.A(net161),
    .X(_04214_));
 sg13g2_nand2_1 _21760_ (.Y(_04215_),
    .A(net241),
    .B(net129));
 sg13g2_nand3_1 _21761_ (.B(_04213_),
    .C(_04215_),
    .A(_04211_),
    .Y(_04216_));
 sg13g2_nor2_1 _21762_ (.A(_09908_),
    .B(\cpu.dec.r_op[7] ),
    .Y(_04217_));
 sg13g2_nor2_1 _21763_ (.A(_08255_),
    .B(net1116),
    .Y(_04218_));
 sg13g2_nor4_1 _21764_ (.A(_09001_),
    .B(net1124),
    .C(\cpu.dec.r_op[9] ),
    .D(_09889_),
    .Y(_04219_));
 sg13g2_nor2_1 _21765_ (.A(_09166_),
    .B(_09180_),
    .Y(_04220_));
 sg13g2_nand4_1 _21766_ (.B(_04217_),
    .C(_04219_),
    .A(_04218_),
    .Y(_04221_),
    .D(_04220_));
 sg13g2_buf_1 _21767_ (.A(_04221_),
    .X(_04222_));
 sg13g2_and2_1 _21768_ (.A(_04217_),
    .B(_04222_),
    .X(_04223_));
 sg13g2_buf_1 _21769_ (.A(_04223_),
    .X(_04224_));
 sg13g2_nand3_1 _21770_ (.B(_03779_),
    .C(_03781_),
    .A(_10552_),
    .Y(_04225_));
 sg13g2_buf_1 _21771_ (.A(_04225_),
    .X(_04226_));
 sg13g2_nand2_1 _21772_ (.Y(_04227_),
    .A(_03779_),
    .B(_03781_));
 sg13g2_buf_2 _21773_ (.A(_04227_),
    .X(_04228_));
 sg13g2_nand2_1 _21774_ (.Y(_04229_),
    .A(net238),
    .B(_04228_));
 sg13g2_buf_1 _21775_ (.A(_03783_),
    .X(_04230_));
 sg13g2_buf_1 _21776_ (.A(net225),
    .X(_04231_));
 sg13g2_a21oi_1 _21777_ (.A1(_04226_),
    .A2(_04229_),
    .Y(_04232_),
    .B1(net198));
 sg13g2_nor2_1 _21778_ (.A(_04224_),
    .B(_04232_),
    .Y(_04233_));
 sg13g2_nand2_1 _21779_ (.Y(_04234_),
    .A(_04226_),
    .B(_04229_));
 sg13g2_a21o_1 _21780_ (.A2(_04224_),
    .A1(net225),
    .B1(net286),
    .X(_04235_));
 sg13g2_nand2_1 _21781_ (.Y(_04236_),
    .A(_04217_),
    .B(_04222_));
 sg13g2_buf_2 _21782_ (.A(_04236_),
    .X(_04237_));
 sg13g2_nor2_1 _21783_ (.A(_03783_),
    .B(_04237_),
    .Y(_04238_));
 sg13g2_a21oi_1 _21784_ (.A1(net832),
    .A2(net225),
    .Y(_04239_),
    .B1(_04238_));
 sg13g2_nor3_1 _21785_ (.A(net286),
    .B(_04234_),
    .C(_04239_),
    .Y(_04240_));
 sg13g2_a21oi_1 _21786_ (.A1(_04234_),
    .A2(_04235_),
    .Y(_04241_),
    .B1(_04240_));
 sg13g2_o21ai_1 _21787_ (.B1(_04241_),
    .Y(_04242_),
    .A1(_09180_),
    .A2(_04233_));
 sg13g2_mux2_1 _21788_ (.A0(net1047),
    .A1(net1046),
    .S(_04229_),
    .X(_04243_));
 sg13g2_o21ai_1 _21789_ (.B1(_04226_),
    .Y(_04244_),
    .A1(net1033),
    .A2(_04243_));
 sg13g2_and2_1 _21790_ (.A(_09889_),
    .B(net198),
    .X(_04245_));
 sg13g2_buf_1 _21791_ (.A(_11534_),
    .X(_04246_));
 sg13g2_a221oi_1 _21792_ (.B2(_04245_),
    .C1(net331),
    .B1(net129),
    .A1(_09001_),
    .Y(_04247_),
    .A2(_11372_));
 sg13g2_nand4_1 _21793_ (.B(_04242_),
    .C(_04244_),
    .A(_04216_),
    .Y(_04248_),
    .D(_04247_));
 sg13g2_o21ai_1 _21794_ (.B1(_04248_),
    .Y(_04249_),
    .A1(_04143_),
    .A2(\cpu.ex.c_mult[1] ));
 sg13g2_or2_1 _21795_ (.X(_04250_),
    .B(_10743_),
    .A(_08615_));
 sg13g2_buf_1 _21796_ (.A(_04250_),
    .X(_04251_));
 sg13g2_nand2_1 _21797_ (.Y(_04252_),
    .A(_08580_),
    .B(net658));
 sg13g2_nor2_1 _21798_ (.A(_04251_),
    .B(_04252_),
    .Y(_04253_));
 sg13g2_and2_1 _21799_ (.A(_11911_),
    .B(_04253_),
    .X(_04254_));
 sg13g2_buf_1 _21800_ (.A(_04254_),
    .X(_04255_));
 sg13g2_nor2_1 _21801_ (.A(_10582_),
    .B(_10734_),
    .Y(_04256_));
 sg13g2_buf_1 _21802_ (.A(_04256_),
    .X(_04257_));
 sg13g2_nand2_1 _21803_ (.Y(_04258_),
    .A(\cpu.dec.iready ),
    .B(_00199_));
 sg13g2_nor2_1 _21804_ (.A(\cpu.ex.r_branch_stall ),
    .B(_04258_),
    .Y(_04259_));
 sg13g2_buf_2 _21805_ (.A(_04259_),
    .X(_04260_));
 sg13g2_nand3_1 _21806_ (.B(net330),
    .C(_04260_),
    .A(_09212_),
    .Y(_04261_));
 sg13g2_o21ai_1 _21807_ (.B1(_04261_),
    .Y(_04262_),
    .A1(net330),
    .A2(_04260_));
 sg13g2_nand4_1 _21808_ (.B(_09213_),
    .C(_09258_),
    .A(_08580_),
    .Y(_04263_),
    .D(net658));
 sg13g2_nand2_1 _21809_ (.Y(_04264_),
    .A(_09381_),
    .B(_04263_));
 sg13g2_a221oi_1 _21810_ (.B2(_08576_),
    .C1(_04264_),
    .B1(_04262_),
    .A1(_11911_),
    .Y(_04265_),
    .A2(_04253_));
 sg13g2_and2_1 _21811_ (.A(_04140_),
    .B(_04265_),
    .X(_04266_));
 sg13g2_buf_1 _21812_ (.A(_04266_),
    .X(_04267_));
 sg13g2_buf_1 _21813_ (.A(_04267_),
    .X(_04268_));
 sg13g2_a22oi_1 _21814_ (.Y(_04269_),
    .B1(net61),
    .B2(net794),
    .A2(net96),
    .A1(_11110_));
 sg13g2_o21ai_1 _21815_ (.B1(_04269_),
    .Y(_00980_),
    .A1(net82),
    .A2(_04249_));
 sg13g2_buf_1 _21816_ (.A(_04143_),
    .X(_04270_));
 sg13g2_a221oi_1 _21817_ (.B2(_11766_),
    .C1(net278),
    .B1(net58),
    .A1(\cpu.ex.r_mult[11] ),
    .Y(_04271_),
    .A2(_11660_));
 sg13g2_nand2_1 _21818_ (.Y(_04272_),
    .A(_11717_),
    .B(_11791_));
 sg13g2_nand2_1 _21819_ (.Y(_04273_),
    .A(_11717_),
    .B(_11786_));
 sg13g2_mux2_1 _21820_ (.A0(_04272_),
    .A1(_04273_),
    .S(_11785_),
    .X(_04274_));
 sg13g2_nand2_1 _21821_ (.Y(_04275_),
    .A(_03743_),
    .B(_03737_));
 sg13g2_nand2_1 _21822_ (.Y(_04276_),
    .A(net188),
    .B(_03733_));
 sg13g2_nand4_1 _21823_ (.B(_03824_),
    .C(_03818_),
    .A(_03733_),
    .Y(_04277_),
    .D(_03828_));
 sg13g2_nand4_1 _21824_ (.B(_03824_),
    .C(_03818_),
    .A(net188),
    .Y(_04278_),
    .D(_03828_));
 sg13g2_or2_1 _21825_ (.X(_04279_),
    .B(_03831_),
    .A(_03830_));
 sg13g2_a21o_1 _21826_ (.A2(_04179_),
    .A1(net214),
    .B1(_04279_),
    .X(_04280_));
 sg13g2_nand4_1 _21827_ (.B(_04277_),
    .C(_04278_),
    .A(_04276_),
    .Y(_04281_),
    .D(_04280_));
 sg13g2_buf_1 _21828_ (.A(_04281_),
    .X(_04282_));
 sg13g2_xnor2_1 _21829_ (.Y(_04283_),
    .A(_04275_),
    .B(_04282_));
 sg13g2_nor2_1 _21830_ (.A(_03717_),
    .B(_03722_),
    .Y(_04284_));
 sg13g2_o21ai_1 _21831_ (.B1(_03734_),
    .Y(_04285_),
    .A1(_04284_),
    .A2(_03744_));
 sg13g2_xor2_1 _21832_ (.B(_04275_),
    .A(_04285_),
    .X(_04286_));
 sg13g2_and4_1 _21833_ (.A(_04218_),
    .B(_04217_),
    .C(_04219_),
    .D(_04220_),
    .X(_04287_));
 sg13g2_buf_1 _21834_ (.A(_04287_),
    .X(_04288_));
 sg13g2_nand2_1 _21835_ (.Y(_04289_),
    .A(_03668_),
    .B(_03706_));
 sg13g2_o21ai_1 _21836_ (.B1(net168),
    .Y(_04290_),
    .A1(_03668_),
    .A2(_03706_));
 sg13g2_nor2_1 _21837_ (.A(_11379_),
    .B(_03657_),
    .Y(_04291_));
 sg13g2_a21o_1 _21838_ (.A2(_04290_),
    .A1(_04289_),
    .B1(_04291_),
    .X(_04292_));
 sg13g2_buf_1 _21839_ (.A(_04292_),
    .X(_04293_));
 sg13g2_and2_1 _21840_ (.A(_03650_),
    .B(_03660_),
    .X(_04294_));
 sg13g2_buf_1 _21841_ (.A(_04294_),
    .X(_04295_));
 sg13g2_nand2b_1 _21842_ (.Y(_04296_),
    .B(_09908_),
    .A_N(_04295_));
 sg13g2_a21oi_1 _21843_ (.A1(_03671_),
    .A2(_04293_),
    .Y(_04297_),
    .B1(_04296_));
 sg13g2_and4_1 _21844_ (.A(_09908_),
    .B(_03671_),
    .C(_04293_),
    .D(_04295_),
    .X(_04298_));
 sg13g2_buf_1 _21845_ (.A(_04298_),
    .X(_04299_));
 sg13g2_nor3_2 _21846_ (.A(net331),
    .B(_04297_),
    .C(_04299_),
    .Y(_04300_));
 sg13g2_buf_1 _21847_ (.A(net165),
    .X(_04301_));
 sg13g2_nand3_1 _21848_ (.B(_10552_),
    .C(_10507_),
    .A(_03784_),
    .Y(_04302_));
 sg13g2_buf_2 _21849_ (.A(_04302_),
    .X(_04303_));
 sg13g2_nand2_1 _21850_ (.Y(_04304_),
    .A(_11019_),
    .B(_10507_));
 sg13g2_a21oi_1 _21851_ (.A1(net164),
    .A2(net156),
    .Y(_04305_),
    .B1(net161));
 sg13g2_o21ai_1 _21852_ (.B1(_04305_),
    .Y(_04306_),
    .A1(_03767_),
    .A2(_04304_));
 sg13g2_buf_1 _21853_ (.A(net179),
    .X(_04307_));
 sg13g2_and2_1 _21854_ (.A(net114),
    .B(net155),
    .X(_04308_));
 sg13g2_o21ai_1 _21855_ (.B1(net1116),
    .Y(_04309_),
    .A1(_04306_),
    .A2(_04308_));
 sg13g2_a21oi_1 _21856_ (.A1(net285),
    .A2(_11485_),
    .Y(_04310_),
    .B1(net240));
 sg13g2_nor2_1 _21857_ (.A(_03773_),
    .B(_04310_),
    .Y(_04311_));
 sg13g2_a21o_1 _21858_ (.A2(_04156_),
    .A1(net114),
    .B1(_04311_),
    .X(_04312_));
 sg13g2_o21ai_1 _21859_ (.B1(net1073),
    .Y(_04313_),
    .A1(_04306_),
    .A2(_04312_));
 sg13g2_nand2_1 _21860_ (.Y(_04314_),
    .A(_04309_),
    .B(_04313_));
 sg13g2_o21ai_1 _21861_ (.B1(_04314_),
    .Y(_04315_),
    .A1(net128),
    .A2(_04303_));
 sg13g2_buf_1 _21862_ (.A(_03699_),
    .X(_04316_));
 sg13g2_o21ai_1 _21863_ (.B1(_04303_),
    .Y(_04317_),
    .A1(_03714_),
    .A2(_04304_));
 sg13g2_a21oi_1 _21864_ (.A1(_04316_),
    .A2(_04177_),
    .Y(_04318_),
    .B1(_04317_));
 sg13g2_buf_1 _21865_ (.A(net156),
    .X(_04319_));
 sg13g2_a22oi_1 _21866_ (.Y(_04320_),
    .B1(_04319_),
    .B2(_04187_),
    .A2(_04307_),
    .A1(net163));
 sg13g2_buf_1 _21867_ (.A(_04186_),
    .X(_04321_));
 sg13g2_buf_1 _21868_ (.A(net167),
    .X(_04322_));
 sg13g2_a22oi_1 _21869_ (.Y(_04323_),
    .B1(_04321_),
    .B2(net125),
    .A2(net159),
    .A1(net131));
 sg13g2_buf_1 _21870_ (.A(_04228_),
    .X(_04324_));
 sg13g2_a22oi_1 _21871_ (.Y(_04325_),
    .B1(net157),
    .B2(_04231_),
    .A2(net158),
    .A1(net124));
 sg13g2_buf_1 _21872_ (.A(_03801_),
    .X(_04326_));
 sg13g2_a22oi_1 _21873_ (.Y(_04327_),
    .B1(_04162_),
    .B2(net134),
    .A2(net182),
    .A1(net123));
 sg13g2_and4_1 _21874_ (.A(_04320_),
    .B(_04323_),
    .C(_04325_),
    .D(_04327_),
    .X(_04328_));
 sg13g2_nand2_1 _21875_ (.Y(_04329_),
    .A(_04318_),
    .B(_04328_));
 sg13g2_nand2_1 _21876_ (.Y(_04330_),
    .A(_03733_),
    .B(net129));
 sg13g2_nand3_1 _21877_ (.B(_04329_),
    .C(_04330_),
    .A(net1032),
    .Y(_04331_));
 sg13g2_mux2_1 _21878_ (.A0(net1047),
    .A1(net1046),
    .S(_03743_),
    .X(_04332_));
 sg13g2_or2_1 _21879_ (.X(_04333_),
    .B(_04332_),
    .A(net1033));
 sg13g2_a22oi_1 _21880_ (.Y(_04334_),
    .B1(_03737_),
    .B2(_04333_),
    .A2(net240),
    .A1(_09002_));
 sg13g2_nand4_1 _21881_ (.B(_04315_),
    .C(_04331_),
    .A(_04300_),
    .Y(_04335_),
    .D(_04334_));
 sg13g2_a221oi_1 _21882_ (.B2(_04288_),
    .C1(_04335_),
    .B1(_04286_),
    .A1(net1045),
    .Y(_04336_),
    .A2(_04283_));
 sg13g2_a21o_1 _21883_ (.A2(_04274_),
    .A1(_04271_),
    .B1(_04336_),
    .X(_04337_));
 sg13g2_inv_1 _21884_ (.Y(_04338_),
    .A(_00288_));
 sg13g2_nand2_1 _21885_ (.Y(_04339_),
    .A(net928),
    .B(net704));
 sg13g2_nor2_2 _21886_ (.A(_08817_),
    .B(_04339_),
    .Y(_04340_));
 sg13g2_nand4_1 _21887_ (.B(_08777_),
    .C(_08797_),
    .A(_08829_),
    .Y(_04341_),
    .D(_04340_));
 sg13g2_nor2_1 _21888_ (.A(_08820_),
    .B(_04341_),
    .Y(_04342_));
 sg13g2_nand3_1 _21889_ (.B(_08807_),
    .C(_04342_),
    .A(_08786_),
    .Y(_04343_));
 sg13g2_xnor2_1 _21890_ (.Y(_04344_),
    .A(_04338_),
    .B(_04343_));
 sg13g2_buf_1 _21891_ (.A(_04255_),
    .X(_04345_));
 sg13g2_a22oi_1 _21892_ (.Y(_04346_),
    .B1(_04344_),
    .B2(net81),
    .A2(net61),
    .A1(\cpu.ex.pc[11] ));
 sg13g2_o21ai_1 _21893_ (.B1(_04346_),
    .Y(_00981_),
    .A1(net82),
    .A2(_04337_));
 sg13g2_inv_1 _21894_ (.Y(_04347_),
    .A(_03737_));
 sg13g2_a21oi_1 _21895_ (.A1(_03743_),
    .A2(_04285_),
    .Y(_04348_),
    .B1(_04347_));
 sg13g2_nand2_1 _21896_ (.Y(_04349_),
    .A(_03728_),
    .B(_03754_));
 sg13g2_xor2_1 _21897_ (.B(_04349_),
    .A(_04348_),
    .X(_04350_));
 sg13g2_or3_1 _21898_ (.A(net331),
    .B(_04297_),
    .C(_04299_),
    .X(_04351_));
 sg13g2_and3_1 _21899_ (.X(_04352_),
    .A(_03824_),
    .B(_03818_),
    .C(_03828_));
 sg13g2_o21ai_1 _21900_ (.B1(_03823_),
    .Y(_04353_),
    .A1(_04352_),
    .A2(_03833_));
 sg13g2_xnor2_1 _21901_ (.Y(_04354_),
    .A(_04353_),
    .B(_04349_));
 sg13g2_nor2_1 _21902_ (.A(net832),
    .B(_04354_),
    .Y(_04355_));
 sg13g2_nand2_1 _21903_ (.Y(_04356_),
    .A(net135),
    .B(_04192_));
 sg13g2_nand2_1 _21904_ (.Y(_04357_),
    .A(net132),
    .B(_04148_));
 sg13g2_nor4_1 _21905_ (.A(_11510_),
    .B(net238),
    .C(_11594_),
    .D(net279),
    .Y(_04358_));
 sg13g2_buf_2 _21906_ (.A(_04358_),
    .X(_04359_));
 sg13g2_a22oi_1 _21907_ (.Y(_04360_),
    .B1(_04359_),
    .B2(net125),
    .A2(net157),
    .A1(net124));
 sg13g2_and2_1 _21908_ (.A(net163),
    .B(_04160_),
    .X(_04361_));
 sg13g2_a221oi_1 _21909_ (.B2(net133),
    .C1(_04361_),
    .B1(_04319_),
    .A1(_04189_),
    .Y(_04362_),
    .A2(net182));
 sg13g2_nand4_1 _21910_ (.B(_04357_),
    .C(_04360_),
    .A(_04356_),
    .Y(_04363_),
    .D(_04362_));
 sg13g2_buf_1 _21911_ (.A(net161),
    .X(_04364_));
 sg13g2_a21oi_1 _21912_ (.A1(_04163_),
    .A2(net159),
    .Y(_04365_),
    .B1(net122));
 sg13g2_nand2_1 _21913_ (.Y(_04366_),
    .A(net127),
    .B(_04195_));
 sg13g2_a22oi_1 _21914_ (.Y(_04367_),
    .B1(_04202_),
    .B2(_04231_),
    .A2(net154),
    .A1(net123));
 sg13g2_nand3_1 _21915_ (.B(_04366_),
    .C(_04367_),
    .A(_04365_),
    .Y(_04368_));
 sg13g2_nor2_1 _21916_ (.A(_04363_),
    .B(_04368_),
    .Y(_04369_));
 sg13g2_nand2_1 _21917_ (.Y(_04370_),
    .A(_03736_),
    .B(net129));
 sg13g2_nand2_1 _21918_ (.Y(_04371_),
    .A(net1032),
    .B(_04370_));
 sg13g2_mux2_1 _21919_ (.A0(net1124),
    .A1(_09166_),
    .S(_03754_),
    .X(_04372_));
 sg13g2_or2_1 _21920_ (.X(_04373_),
    .B(_04372_),
    .A(net1115));
 sg13g2_a22oi_1 _21921_ (.Y(_04374_),
    .B1(_03728_),
    .B2(_04373_),
    .A2(net287),
    .A1(net1048));
 sg13g2_o21ai_1 _21922_ (.B1(_04374_),
    .Y(_04375_),
    .A1(_04369_),
    .A2(_04371_));
 sg13g2_nor2_1 _21923_ (.A(_03774_),
    .B(_04303_),
    .Y(_04376_));
 sg13g2_a22oi_1 _21924_ (.Y(_04377_),
    .B1(_04208_),
    .B2(_03752_),
    .A2(net162),
    .A1(net138));
 sg13g2_nand2_1 _21925_ (.Y(_04378_),
    .A(_04303_),
    .B(_04377_));
 sg13g2_or2_1 _21926_ (.X(_04379_),
    .B(_04378_),
    .A(_04312_));
 sg13g2_a22oi_1 _21927_ (.Y(_04380_),
    .B1(_04379_),
    .B2(net1073),
    .A2(_04378_),
    .A1(_09880_));
 sg13g2_nor2_1 _21928_ (.A(_04376_),
    .B(_04380_),
    .Y(_04381_));
 sg13g2_nor4_1 _21929_ (.A(_04351_),
    .B(_04355_),
    .C(_04375_),
    .D(_04381_),
    .Y(_04382_));
 sg13g2_o21ai_1 _21930_ (.B1(_04382_),
    .Y(_04383_),
    .A1(_04222_),
    .A2(_04350_));
 sg13g2_o21ai_1 _21931_ (.B1(_04383_),
    .Y(_04384_),
    .A1(net278),
    .A2(\cpu.ex.c_mult[12] ));
 sg13g2_nor2_1 _21932_ (.A(_08769_),
    .B(_04343_),
    .Y(_04385_));
 sg13g2_xnor2_1 _21933_ (.Y(_04386_),
    .A(_00287_),
    .B(_04385_));
 sg13g2_a22oi_1 _21934_ (.Y(_04387_),
    .B1(_04386_),
    .B2(net81),
    .A2(net61),
    .A1(net790));
 sg13g2_o21ai_1 _21935_ (.B1(_04387_),
    .Y(_00982_),
    .A1(net82),
    .A2(_04384_));
 sg13g2_and2_1 _21936_ (.A(_03759_),
    .B(_03764_),
    .X(_04388_));
 sg13g2_buf_1 _21937_ (.A(_04388_),
    .X(_04389_));
 sg13g2_nor2_1 _21938_ (.A(net211),
    .B(net130),
    .Y(_04390_));
 sg13g2_or3_1 _21939_ (.A(_03834_),
    .B(_04390_),
    .C(_04282_),
    .X(_04391_));
 sg13g2_a221oi_1 _21940_ (.B2(_04391_),
    .C1(net832),
    .B1(_04389_),
    .A1(net213),
    .Y(_04392_),
    .A2(net128));
 sg13g2_o21ai_1 _21941_ (.B1(_03736_),
    .Y(_04393_),
    .A1(_04282_),
    .A2(_04389_));
 sg13g2_nor2_1 _21942_ (.A(_11411_),
    .B(_03834_),
    .Y(_04394_));
 sg13g2_nor4_1 _21943_ (.A(_03736_),
    .B(_03834_),
    .C(_04282_),
    .D(_04389_),
    .Y(_04395_));
 sg13g2_a21oi_1 _21944_ (.A1(_04393_),
    .A2(_04394_),
    .Y(_04396_),
    .B1(_04395_));
 sg13g2_and2_1 _21945_ (.A(_10383_),
    .B(net128),
    .X(_04397_));
 sg13g2_nor3_2 _21946_ (.A(_03739_),
    .B(_03747_),
    .C(_04397_),
    .Y(_04398_));
 sg13g2_xnor2_1 _21947_ (.Y(_04399_),
    .A(_04398_),
    .B(_04389_));
 sg13g2_o21ai_1 _21948_ (.B1(net1032),
    .Y(_04400_),
    .A1(net128),
    .A2(_04303_));
 sg13g2_a21oi_1 _21949_ (.A1(net133),
    .A2(_04149_),
    .Y(_04401_),
    .B1(net129));
 sg13g2_nand2_1 _21950_ (.Y(_04402_),
    .A(net127),
    .B(net157));
 sg13g2_a22oi_1 _21951_ (.Y(_04403_),
    .B1(net158),
    .B2(_04322_),
    .A2(net154),
    .A1(_04189_));
 sg13g2_a22oi_1 _21952_ (.Y(_04404_),
    .B1(_04205_),
    .B2(net225),
    .A2(_04202_),
    .A1(_04228_));
 sg13g2_a22oi_1 _21953_ (.Y(_04405_),
    .B1(_04359_),
    .B2(net123),
    .A2(net160),
    .A1(net135));
 sg13g2_and4_1 _21954_ (.A(_04402_),
    .B(_04403_),
    .C(_04404_),
    .D(_04405_),
    .X(_04406_));
 sg13g2_a22oi_1 _21955_ (.Y(_04407_),
    .B1(net182),
    .B2(net134),
    .A2(_04175_),
    .A1(_03803_));
 sg13g2_a22oi_1 _21956_ (.Y(_04408_),
    .B1(net126),
    .B2(net130),
    .A2(net155),
    .A1(_04187_));
 sg13g2_nand4_1 _21957_ (.B(_04406_),
    .C(_04407_),
    .A(_04401_),
    .Y(_04409_),
    .D(_04408_));
 sg13g2_nand2b_1 _21958_ (.Y(_04410_),
    .B(_04409_),
    .A_N(_04400_));
 sg13g2_nand2_1 _21959_ (.Y(_04411_),
    .A(_11767_),
    .B(net130));
 sg13g2_o21ai_1 _21960_ (.B1(_03837_),
    .Y(_04412_),
    .A1(_03834_),
    .A2(_04411_));
 sg13g2_a21o_1 _21961_ (.A2(_04412_),
    .A1(_09180_),
    .B1(net1046),
    .X(_04413_));
 sg13g2_nor2b_1 _21962_ (.A(_11833_),
    .B_N(net1115),
    .Y(_04414_));
 sg13g2_a21oi_1 _21963_ (.A1(_09001_),
    .A2(_11614_),
    .Y(_04415_),
    .B1(_04414_));
 sg13g2_nor2b_1 _21964_ (.A(_11833_),
    .B_N(net1124),
    .Y(_04416_));
 sg13g2_o21ai_1 _21965_ (.B1(_03774_),
    .Y(_04417_),
    .A1(_09886_),
    .A2(_04416_));
 sg13g2_o21ai_1 _21966_ (.B1(net1073),
    .Y(_04418_),
    .A1(_03644_),
    .A2(_04364_));
 sg13g2_nand2_1 _21967_ (.Y(_04419_),
    .A(_03767_),
    .B(net122));
 sg13g2_nand2b_1 _21968_ (.Y(_04420_),
    .B(_04419_),
    .A_N(_04418_));
 sg13g2_a22oi_1 _21969_ (.Y(_04421_),
    .B1(net126),
    .B2(net114),
    .A2(_04364_),
    .A1(_03752_));
 sg13g2_nand2b_1 _21970_ (.Y(_04422_),
    .B(net1116),
    .A_N(_04421_));
 sg13g2_nand4_1 _21971_ (.B(_04417_),
    .C(_04420_),
    .A(_04415_),
    .Y(_04423_),
    .D(_04422_));
 sg13g2_a21oi_1 _21972_ (.A1(_04389_),
    .A2(_04413_),
    .Y(_04424_),
    .B1(_04423_));
 sg13g2_nand3_1 _21973_ (.B(_04410_),
    .C(_04424_),
    .A(_04300_),
    .Y(_04425_));
 sg13g2_a221oi_1 _21974_ (.B2(_04288_),
    .C1(_04425_),
    .B1(_04399_),
    .A1(_04392_),
    .Y(_04426_),
    .A2(_04396_));
 sg13g2_a21o_1 _21975_ (.A2(_11840_),
    .A1(_04246_),
    .B1(_04426_),
    .X(_04427_));
 sg13g2_nand2_1 _21976_ (.Y(_04428_),
    .A(net790),
    .B(_04385_));
 sg13g2_xnor2_1 _21977_ (.Y(_04429_),
    .A(_03755_),
    .B(_04428_));
 sg13g2_a22oi_1 _21978_ (.Y(_04430_),
    .B1(_04429_),
    .B2(net81),
    .A2(net61),
    .A1(net912));
 sg13g2_o21ai_1 _21979_ (.B1(_04430_),
    .Y(_00983_),
    .A1(net82),
    .A2(_04427_));
 sg13g2_nand2_1 _21980_ (.Y(_04431_),
    .A(_11469_),
    .B(net166));
 sg13g2_nand2_2 _21981_ (.Y(_04432_),
    .A(_03768_),
    .B(_04431_));
 sg13g2_nor2b_1 _21982_ (.A(_04432_),
    .B_N(_03759_),
    .Y(_04433_));
 sg13g2_nand2_1 _21983_ (.Y(_04434_),
    .A(_03764_),
    .B(_04432_));
 sg13g2_nor2_1 _21984_ (.A(_04398_),
    .B(_04434_),
    .Y(_04435_));
 sg13g2_a21oi_1 _21985_ (.A1(_04398_),
    .A2(_04433_),
    .Y(_04436_),
    .B1(_04435_));
 sg13g2_nand2b_1 _21986_ (.Y(_04437_),
    .B(_04432_),
    .A_N(_03838_));
 sg13g2_nand2_1 _21987_ (.Y(_04438_),
    .A(_03836_),
    .B(_03837_));
 sg13g2_nand4_1 _21988_ (.B(_04431_),
    .C(_03776_),
    .A(_03768_),
    .Y(_04439_),
    .D(_04438_));
 sg13g2_a21oi_1 _21989_ (.A1(_04437_),
    .A2(_04439_),
    .Y(_04440_),
    .B1(net832));
 sg13g2_mux2_1 _21990_ (.A0(_03777_),
    .A1(_03776_),
    .S(_04432_),
    .X(_04441_));
 sg13g2_a21o_1 _21991_ (.A2(_04214_),
    .A1(net1116),
    .B1(_08256_),
    .X(_04442_));
 sg13g2_a22oi_1 _21992_ (.Y(_04443_),
    .B1(_03644_),
    .B2(_04442_),
    .A2(_11379_),
    .A1(net1048));
 sg13g2_o21ai_1 _21993_ (.B1(_04443_),
    .Y(_04444_),
    .A1(_03844_),
    .A2(_04441_));
 sg13g2_mux2_1 _21994_ (.A0(net1047),
    .A1(net1046),
    .S(_04431_),
    .X(_04445_));
 sg13g2_o21ai_1 _21995_ (.B1(_03768_),
    .Y(_04446_),
    .A1(_09887_),
    .A2(_04445_));
 sg13g2_nand2b_1 _21996_ (.Y(_04447_),
    .B(_04446_),
    .A_N(_04444_));
 sg13g2_mux2_1 _21997_ (.A0(_03764_),
    .A1(_03759_),
    .S(_04432_),
    .X(_04448_));
 sg13g2_a21oi_1 _21998_ (.A1(_03742_),
    .A2(_04148_),
    .Y(_04449_),
    .B1(_04151_));
 sg13g2_a22oi_1 _21999_ (.Y(_04450_),
    .B1(_04321_),
    .B2(net134),
    .A2(_04183_),
    .A1(net198));
 sg13g2_a22oi_1 _22000_ (.Y(_04451_),
    .B1(_04359_),
    .B2(net131),
    .A2(net157),
    .A1(net125));
 sg13g2_a22oi_1 _22001_ (.Y(_04452_),
    .B1(net126),
    .B2(net128),
    .A2(net159),
    .A1(net135));
 sg13g2_nand4_1 _22002_ (.B(_04450_),
    .C(_04451_),
    .A(_04449_),
    .Y(_04453_),
    .D(_04452_));
 sg13g2_nand2_1 _22003_ (.Y(_04454_),
    .A(net133),
    .B(net179));
 sg13g2_nand2_1 _22004_ (.Y(_04455_),
    .A(net163),
    .B(net182));
 sg13g2_a22oi_1 _22005_ (.Y(_04456_),
    .B1(_04205_),
    .B2(net124),
    .A2(net160),
    .A1(net132));
 sg13g2_a22oi_1 _22006_ (.Y(_04457_),
    .B1(_04202_),
    .B2(net127),
    .A2(net158),
    .A1(_04326_));
 sg13g2_nand4_1 _22007_ (.B(_04455_),
    .C(_04456_),
    .A(_04454_),
    .Y(_04458_),
    .D(_04457_));
 sg13g2_nor2b_1 _22008_ (.A(_04376_),
    .B_N(_09890_),
    .Y(_04459_));
 sg13g2_o21ai_1 _22009_ (.B1(_04459_),
    .Y(_04460_),
    .A1(_04453_),
    .A2(_04458_));
 sg13g2_o21ai_1 _22010_ (.B1(_04460_),
    .Y(_04461_),
    .A1(_04222_),
    .A2(_04448_));
 sg13g2_nor4_1 _22011_ (.A(_04351_),
    .B(_04440_),
    .C(_04447_),
    .D(_04461_),
    .Y(_04462_));
 sg13g2_o21ai_1 _22012_ (.B1(_04462_),
    .Y(_04463_),
    .A1(_04222_),
    .A2(_04436_));
 sg13g2_o21ai_1 _22013_ (.B1(_04463_),
    .Y(_04464_),
    .A1(net278),
    .A2(\cpu.ex.c_mult[14] ));
 sg13g2_nand3_1 _22014_ (.B(net912),
    .C(_04385_),
    .A(net790),
    .Y(_04465_));
 sg13g2_xnor2_1 _22015_ (.Y(_04466_),
    .A(_03748_),
    .B(_04465_));
 sg13g2_a22oi_1 _22016_ (.Y(_04467_),
    .B1(_04466_),
    .B2(net81),
    .A2(net61),
    .A1(net915));
 sg13g2_o21ai_1 _22017_ (.B1(_04467_),
    .Y(_00984_),
    .A1(net82),
    .A2(_04464_));
 sg13g2_nand2_1 _22018_ (.Y(_04468_),
    .A(_11442_),
    .B(net114));
 sg13g2_nand2_1 _22019_ (.Y(_04469_),
    .A(_11872_),
    .B(_03773_));
 sg13g2_a21oi_1 _22020_ (.A1(_04468_),
    .A2(_04469_),
    .Y(_04470_),
    .B1(net832));
 sg13g2_nand2_1 _22021_ (.Y(_04471_),
    .A(_04468_),
    .B(_04469_));
 sg13g2_nor4_1 _22022_ (.A(net832),
    .B(_03839_),
    .C(_03840_),
    .D(_04471_),
    .Y(_04472_));
 sg13g2_a21oi_1 _22023_ (.A1(_03839_),
    .A2(_04470_),
    .Y(_04473_),
    .B1(_04472_));
 sg13g2_a22oi_1 _22024_ (.Y(_04474_),
    .B1(_04200_),
    .B2(_04326_),
    .A2(_04177_),
    .A1(net134));
 sg13g2_a22oi_1 _22025_ (.Y(_04475_),
    .B1(_04202_),
    .B2(net125),
    .A2(net182),
    .A1(_04155_));
 sg13g2_and2_1 _22026_ (.A(net130),
    .B(net155),
    .X(_04476_));
 sg13g2_a221oi_1 _22027_ (.B2(_04324_),
    .C1(_04476_),
    .B1(_04183_),
    .A1(net128),
    .Y(_04477_),
    .A2(_04149_));
 sg13g2_a22oi_1 _22028_ (.Y(_04478_),
    .B1(_04195_),
    .B2(net131),
    .A2(net180),
    .A1(net132));
 sg13g2_a22oi_1 _22029_ (.Y(_04479_),
    .B1(net154),
    .B2(net163),
    .A2(_04161_),
    .A1(net133));
 sg13g2_nand2_1 _22030_ (.Y(_04480_),
    .A(_03783_),
    .B(_11551_));
 sg13g2_o21ai_1 _22031_ (.B1(_04480_),
    .Y(_04481_),
    .A1(net241),
    .A2(_11551_));
 sg13g2_nand3_1 _22032_ (.B(_11599_),
    .C(_04481_),
    .A(_03784_),
    .Y(_04482_));
 sg13g2_and4_1 _22033_ (.A(_04305_),
    .B(_04478_),
    .C(_04479_),
    .D(_04482_),
    .X(_04483_));
 sg13g2_nand4_1 _22034_ (.B(_04475_),
    .C(_04477_),
    .A(_04474_),
    .Y(_04484_),
    .D(_04483_));
 sg13g2_nand3_1 _22035_ (.B(_04419_),
    .C(_04484_),
    .A(net1032),
    .Y(_04485_));
 sg13g2_mux2_1 _22036_ (.A0(net1047),
    .A1(_09167_),
    .S(_04468_),
    .X(_04486_));
 sg13g2_o21ai_1 _22037_ (.B1(_04469_),
    .Y(_04487_),
    .A1(_09887_),
    .A2(_04486_));
 sg13g2_nand3_1 _22038_ (.B(_03840_),
    .C(_04471_),
    .A(net1045),
    .Y(_04488_));
 sg13g2_a21oi_1 _22039_ (.A1(net1048),
    .A2(_11301_),
    .Y(_04489_),
    .B1(_04145_));
 sg13g2_and4_1 _22040_ (.A(_04485_),
    .B(_04487_),
    .C(_04488_),
    .D(_04489_),
    .X(_04490_));
 sg13g2_nand3_1 _22041_ (.B(_04473_),
    .C(_04490_),
    .A(_04300_),
    .Y(_04491_));
 sg13g2_xor2_1 _22042_ (.B(_04471_),
    .A(_03770_),
    .X(_04492_));
 sg13g2_nor2_1 _22043_ (.A(_04222_),
    .B(_04492_),
    .Y(_04493_));
 sg13g2_nor2_1 _22044_ (.A(_11861_),
    .B(_11515_),
    .Y(_04494_));
 sg13g2_a221oi_1 _22045_ (.B2(_03878_),
    .C1(net278),
    .B1(_11727_),
    .A1(_11861_),
    .Y(_04495_),
    .A2(net411));
 sg13g2_o21ai_1 _22046_ (.B1(_04495_),
    .Y(_04496_),
    .A1(_11877_),
    .A2(_04494_));
 sg13g2_o21ai_1 _22047_ (.B1(_04496_),
    .Y(_04497_),
    .A1(_04491_),
    .A2(_04493_));
 sg13g2_or2_1 _22048_ (.X(_04498_),
    .B(_04465_),
    .A(_08871_));
 sg13g2_xnor2_1 _22049_ (.Y(_04499_),
    .A(_03636_),
    .B(_04498_));
 sg13g2_a22oi_1 _22050_ (.Y(_04500_),
    .B1(_04499_),
    .B2(net81),
    .A2(net61),
    .A1(_08538_));
 sg13g2_o21ai_1 _22051_ (.B1(_04500_),
    .Y(_00985_),
    .A1(net82),
    .A2(_04497_));
 sg13g2_nand3_1 _22052_ (.B(net330),
    .C(_11530_),
    .A(_09212_),
    .Y(_04501_));
 sg13g2_a21oi_1 _22053_ (.A1(net923),
    .A2(net96),
    .Y(_04502_),
    .B1(_04267_));
 sg13g2_a21oi_1 _22054_ (.A1(net794),
    .A2(net96),
    .Y(_04503_),
    .B1(net701));
 sg13g2_a21o_1 _22055_ (.A2(_04502_),
    .A1(net701),
    .B1(_04503_),
    .X(_04504_));
 sg13g2_a21oi_2 _22056_ (.B1(_03786_),
    .Y(_04505_),
    .A2(_03785_),
    .A1(_03782_));
 sg13g2_xnor2_1 _22057_ (.Y(_04506_),
    .A(net241),
    .B(net285));
 sg13g2_xnor2_1 _22058_ (.Y(_04507_),
    .A(_04505_),
    .B(_04506_));
 sg13g2_nand2b_1 _22059_ (.Y(_04508_),
    .B(net122),
    .A_N(net125));
 sg13g2_a21oi_1 _22060_ (.A1(_03657_),
    .A2(net179),
    .Y(_04509_),
    .B1(_04151_));
 sg13g2_a22oi_1 _22061_ (.Y(_04510_),
    .B1(net156),
    .B2(_03801_),
    .A2(net180),
    .A1(_03826_));
 sg13g2_a21oi_1 _22062_ (.A1(net130),
    .A2(_04177_),
    .Y(_04511_),
    .B1(_04361_));
 sg13g2_nand2_1 _22063_ (.Y(_04512_),
    .A(net164),
    .B(_04199_));
 sg13g2_a22oi_1 _22064_ (.Y(_04513_),
    .B1(_04186_),
    .B2(_04179_),
    .A2(net199),
    .A1(_03711_));
 sg13g2_a22oi_1 _22065_ (.Y(_04514_),
    .B1(_04205_),
    .B2(_03642_),
    .A2(_04148_),
    .A1(_03668_));
 sg13g2_a22oi_1 _22066_ (.Y(_04515_),
    .B1(_04202_),
    .B2(net166),
    .A2(_04194_),
    .A1(net165));
 sg13g2_and4_1 _22067_ (.A(_04512_),
    .B(_04513_),
    .C(_04514_),
    .D(_04515_),
    .X(_04516_));
 sg13g2_nand4_1 _22068_ (.B(_04510_),
    .C(_04511_),
    .A(_04509_),
    .Y(_04517_),
    .D(_04516_));
 sg13g2_nand2_1 _22069_ (.Y(_04518_),
    .A(net240),
    .B(net279));
 sg13g2_nor2_1 _22070_ (.A(_10552_),
    .B(_04518_),
    .Y(_04519_));
 sg13g2_o21ai_1 _22071_ (.B1(net138),
    .Y(_04520_),
    .A1(_11487_),
    .A2(_04519_));
 sg13g2_nand2b_1 _22072_ (.Y(_04521_),
    .B(_04520_),
    .A_N(_04517_));
 sg13g2_a22oi_1 _22073_ (.Y(_04522_),
    .B1(_04521_),
    .B2(net1073),
    .A2(_04517_),
    .A1(net1116));
 sg13g2_inv_1 _22074_ (.Y(_04523_),
    .A(_04522_));
 sg13g2_a21oi_1 _22075_ (.A1(_10552_),
    .A2(_03694_),
    .Y(_04524_),
    .B1(_03695_));
 sg13g2_xnor2_1 _22076_ (.Y(_04525_),
    .A(_04524_),
    .B(_04506_));
 sg13g2_nand2_1 _22077_ (.Y(_04526_),
    .A(_04237_),
    .B(_04525_));
 sg13g2_a21oi_1 _22078_ (.A1(_09001_),
    .A2(_11731_),
    .Y(_04527_),
    .B1(_11534_));
 sg13g2_a22oi_1 _22079_ (.Y(_04528_),
    .B1(net126),
    .B2(net198),
    .A2(net122),
    .A1(net124));
 sg13g2_nand2b_1 _22080_ (.Y(_04529_),
    .B(net1032),
    .A_N(_04528_));
 sg13g2_nor2_1 _22081_ (.A(net241),
    .B(net285),
    .Y(_04530_));
 sg13g2_mux2_1 _22082_ (.A0(_09166_),
    .A1(net1124),
    .S(_04530_),
    .X(_04531_));
 sg13g2_o21ai_1 _22083_ (.B1(_03683_),
    .Y(_04532_),
    .A1(net1115),
    .A2(_04531_));
 sg13g2_nand4_1 _22084_ (.B(_04527_),
    .C(_04529_),
    .A(_04526_),
    .Y(_04533_),
    .D(_04532_));
 sg13g2_a221oi_1 _22085_ (.B2(_04523_),
    .C1(_04533_),
    .B1(_04508_),
    .A1(net1045),
    .Y(_04534_),
    .A2(_04507_));
 sg13g2_a21oi_1 _22086_ (.A1(net331),
    .A2(_11573_),
    .Y(_04535_),
    .B1(_04534_));
 sg13g2_nand2b_1 _22087_ (.Y(_04536_),
    .B(_04535_),
    .A_N(_04140_));
 sg13g2_nand3_1 _22088_ (.B(_04504_),
    .C(_04536_),
    .A(_04501_),
    .Y(_00986_));
 sg13g2_nand2b_1 _22089_ (.Y(_04537_),
    .B(net161),
    .A_N(net123));
 sg13g2_nand2_1 _22090_ (.Y(_04538_),
    .A(net114),
    .B(_04205_));
 sg13g2_a22oi_1 _22091_ (.Y(_04539_),
    .B1(net181),
    .B2(_03826_),
    .A2(_04173_),
    .A1(_03711_));
 sg13g2_a22oi_1 _22092_ (.Y(_04540_),
    .B1(_04200_),
    .B2(net166),
    .A2(net199),
    .A1(_04179_));
 sg13g2_a21oi_1 _22093_ (.A1(_03657_),
    .A2(_04148_),
    .Y(_04541_),
    .B1(_04151_));
 sg13g2_a22oi_1 _22094_ (.Y(_04542_),
    .B1(_04194_),
    .B2(net164),
    .A2(_04191_),
    .A1(net163));
 sg13g2_nand4_1 _22095_ (.B(_04540_),
    .C(_04541_),
    .A(_04539_),
    .Y(_04543_),
    .D(_04542_));
 sg13g2_a22oi_1 _22096_ (.Y(_04544_),
    .B1(_04186_),
    .B2(_03742_),
    .A2(_04177_),
    .A1(net165));
 sg13g2_nand2_1 _22097_ (.Y(_04545_),
    .A(_03642_),
    .B(_04202_));
 sg13g2_nand2_1 _22098_ (.Y(_04546_),
    .A(_03668_),
    .B(_04207_));
 sg13g2_nand3_1 _22099_ (.B(_04545_),
    .C(_04546_),
    .A(_04544_),
    .Y(_04547_));
 sg13g2_nor2_1 _22100_ (.A(_04543_),
    .B(_04547_),
    .Y(_04548_));
 sg13g2_nand3_1 _22101_ (.B(_04538_),
    .C(_04548_),
    .A(_04520_),
    .Y(_04549_));
 sg13g2_nand2b_1 _22102_ (.Y(_04550_),
    .B(net1116),
    .A_N(_04548_));
 sg13g2_nand2b_1 _22103_ (.Y(_04551_),
    .B(_04550_),
    .A_N(net1073));
 sg13g2_nand3_1 _22104_ (.B(_04549_),
    .C(_04551_),
    .A(_04537_),
    .Y(_04552_));
 sg13g2_nand2_1 _22105_ (.Y(_04553_),
    .A(_11122_),
    .B(net167));
 sg13g2_mux2_1 _22106_ (.A0(net1047),
    .A1(net1046),
    .S(_04553_),
    .X(_04554_));
 sg13g2_nand3_1 _22107_ (.B(_03678_),
    .C(_03680_),
    .A(net237),
    .Y(_04555_));
 sg13g2_o21ai_1 _22108_ (.B1(_04555_),
    .Y(_04556_),
    .A1(net1033),
    .A2(_04554_));
 sg13g2_a221oi_1 _22109_ (.B2(_04228_),
    .C1(net122),
    .B1(net126),
    .A1(net225),
    .Y(_04557_),
    .A2(net162));
 sg13g2_nor2b_1 _22110_ (.A(_04557_),
    .B_N(_09889_),
    .Y(_04558_));
 sg13g2_a221oi_1 _22111_ (.B2(_04558_),
    .C1(net331),
    .B1(_04215_),
    .A1(net1048),
    .Y(_04559_),
    .A2(_11411_));
 sg13g2_nand2_1 _22112_ (.Y(_04560_),
    .A(net279),
    .B(_04505_));
 sg13g2_nor2_1 _22113_ (.A(_03915_),
    .B(_04505_),
    .Y(_04561_));
 sg13g2_a21o_1 _22114_ (.A2(_04560_),
    .A1(net127),
    .B1(_04561_),
    .X(_04562_));
 sg13g2_and2_1 _22115_ (.A(_04553_),
    .B(_04555_),
    .X(_04563_));
 sg13g2_xnor2_1 _22116_ (.Y(_04564_),
    .A(_04562_),
    .B(_04563_));
 sg13g2_o21ai_1 _22117_ (.B1(net241),
    .Y(_04565_),
    .A1(_11563_),
    .A2(_03696_));
 sg13g2_o21ai_1 _22118_ (.B1(_04565_),
    .Y(_04566_),
    .A1(_03915_),
    .A2(_04524_));
 sg13g2_buf_1 _22119_ (.A(_04566_),
    .X(_04567_));
 sg13g2_xnor2_1 _22120_ (.Y(_04568_),
    .A(_04563_),
    .B(_04567_));
 sg13g2_a22oi_1 _22121_ (.Y(_04569_),
    .B1(_04568_),
    .B2(_04237_),
    .A2(_04564_),
    .A1(_09180_));
 sg13g2_nand4_1 _22122_ (.B(_04556_),
    .C(_04559_),
    .A(_04552_),
    .Y(_04570_),
    .D(_04569_));
 sg13g2_o21ai_1 _22123_ (.B1(_04570_),
    .Y(_04571_),
    .A1(_04143_),
    .A2(\cpu.ex.c_mult[3] ));
 sg13g2_nand2_1 _22124_ (.Y(_04572_),
    .A(net701),
    .B(net794));
 sg13g2_a21o_1 _22125_ (.A2(_04572_),
    .A1(net96),
    .B1(_04267_),
    .X(_04573_));
 sg13g2_nor2_1 _22126_ (.A(net702),
    .B(_04572_),
    .Y(_04574_));
 sg13g2_o21ai_1 _22127_ (.B1(_04263_),
    .Y(_04575_),
    .A1(_00272_),
    .A2(_04501_));
 sg13g2_a221oi_1 _22128_ (.B2(net96),
    .C1(_04575_),
    .B1(_04574_),
    .A1(net702),
    .Y(_04576_),
    .A2(_04573_));
 sg13g2_o21ai_1 _22129_ (.B1(_04576_),
    .Y(_00987_),
    .A1(net82),
    .A2(_04571_));
 sg13g2_nand2b_1 _22130_ (.Y(_04577_),
    .B(_03703_),
    .A_N(_03688_));
 sg13g2_a21oi_1 _22131_ (.A1(_03678_),
    .A2(_03680_),
    .Y(_04578_),
    .B1(_11122_));
 sg13g2_o21ai_1 _22132_ (.B1(_03795_),
    .Y(_04579_),
    .A1(_04578_),
    .A2(_04562_));
 sg13g2_xnor2_1 _22133_ (.Y(_04580_),
    .A(_04577_),
    .B(_04579_));
 sg13g2_nor2_1 _22134_ (.A(net237),
    .B(_04567_),
    .Y(_04581_));
 sg13g2_nand2_1 _22135_ (.Y(_04582_),
    .A(net237),
    .B(_04567_));
 sg13g2_o21ai_1 _22136_ (.B1(_04582_),
    .Y(_04583_),
    .A1(net125),
    .A2(_04581_));
 sg13g2_xor2_1 _22137_ (.B(_04583_),
    .A(_04577_),
    .X(_04584_));
 sg13g2_nand2_1 _22138_ (.Y(_04585_),
    .A(net127),
    .B(net126));
 sg13g2_a221oi_1 _22139_ (.B2(net225),
    .C1(net129),
    .B1(net155),
    .A1(net124),
    .Y(_04586_),
    .A2(net162));
 sg13g2_nand2_1 _22140_ (.Y(_04587_),
    .A(_09889_),
    .B(_04508_));
 sg13g2_a21o_1 _22141_ (.A2(_04586_),
    .A1(_04585_),
    .B1(_04587_),
    .X(_04588_));
 sg13g2_a21oi_1 _22142_ (.A1(net1048),
    .A2(_10383_),
    .Y(_04589_),
    .B1(net331));
 sg13g2_mux2_1 _22143_ (.A0(net1046),
    .A1(net1047),
    .S(_03688_),
    .X(_04590_));
 sg13g2_o21ai_1 _22144_ (.B1(_03703_),
    .Y(_04591_),
    .A1(net1115),
    .A2(_04590_));
 sg13g2_a22oi_1 _22145_ (.Y(_04592_),
    .B1(_04177_),
    .B2(net136),
    .A2(net180),
    .A1(_04180_));
 sg13g2_a22oi_1 _22146_ (.Y(_04593_),
    .B1(net157),
    .B2(net138),
    .A2(net199),
    .A1(net130));
 sg13g2_a22oi_1 _22147_ (.Y(_04594_),
    .B1(net158),
    .B2(net137),
    .A2(net154),
    .A1(net128));
 sg13g2_nand4_1 _22148_ (.B(_04592_),
    .C(_04593_),
    .A(_04356_),
    .Y(_04595_),
    .D(_04594_));
 sg13g2_nand2_1 _22149_ (.Y(_04596_),
    .A(net132),
    .B(net160));
 sg13g2_o21ai_1 _22150_ (.B1(_04145_),
    .Y(_04597_),
    .A1(_11487_),
    .A2(_11599_));
 sg13g2_a21oi_1 _22151_ (.A1(net134),
    .A2(net156),
    .Y(_04598_),
    .B1(net161));
 sg13g2_nand2_1 _22152_ (.Y(_04599_),
    .A(net163),
    .B(_04148_));
 sg13g2_nand4_1 _22153_ (.B(_04597_),
    .C(_04598_),
    .A(_04596_),
    .Y(_04600_),
    .D(_04599_));
 sg13g2_nand2b_1 _22154_ (.Y(_04601_),
    .B(net161),
    .A_N(net131));
 sg13g2_and2_1 _22155_ (.A(_04213_),
    .B(_04601_),
    .X(_04602_));
 sg13g2_o21ai_1 _22156_ (.B1(_04602_),
    .Y(_04603_),
    .A1(_04595_),
    .A2(_04600_));
 sg13g2_nand4_1 _22157_ (.B(_04589_),
    .C(_04591_),
    .A(_04588_),
    .Y(_04604_),
    .D(_04603_));
 sg13g2_a221oi_1 _22158_ (.B2(_04237_),
    .C1(_04604_),
    .B1(_04584_),
    .A1(net1045),
    .Y(_04605_),
    .A2(_04580_));
 sg13g2_a21o_1 _22159_ (.A2(_11609_),
    .A1(net331),
    .B1(_04605_),
    .X(_04606_));
 sg13g2_nor2_1 _22160_ (.A(_08264_),
    .B(_04339_),
    .Y(_04607_));
 sg13g2_nor3_1 _22161_ (.A(_08579_),
    .B(net781),
    .C(_04260_),
    .Y(_04608_));
 sg13g2_a21oi_1 _22162_ (.A1(net96),
    .A2(_04339_),
    .Y(_04609_),
    .B1(_04267_));
 sg13g2_nor2_1 _22163_ (.A(_08817_),
    .B(_04609_),
    .Y(_04610_));
 sg13g2_a221oi_1 _22164_ (.B2(_08616_),
    .C1(_04610_),
    .B1(_04608_),
    .A1(net96),
    .Y(_04611_),
    .A2(_04607_));
 sg13g2_o21ai_1 _22165_ (.B1(_04611_),
    .Y(_00988_),
    .A1(net82),
    .A2(_04606_));
 sg13g2_and2_1 _22166_ (.A(net163),
    .B(net156),
    .X(_04612_));
 sg13g2_and2_1 _22167_ (.A(net138),
    .B(net158),
    .X(_04613_));
 sg13g2_nand2_1 _22168_ (.Y(_04614_),
    .A(net132),
    .B(net179));
 sg13g2_nand2_1 _22169_ (.Y(_04615_),
    .A(net133),
    .B(net181));
 sg13g2_a22oi_1 _22170_ (.Y(_04616_),
    .B1(_04186_),
    .B2(net164),
    .A2(net199),
    .A1(net165));
 sg13g2_a22oi_1 _22171_ (.Y(_04617_),
    .B1(_04359_),
    .B2(net166),
    .A2(net180),
    .A1(_03742_));
 sg13g2_nand4_1 _22172_ (.B(_04615_),
    .C(_04616_),
    .A(_04614_),
    .Y(_04618_),
    .D(_04617_));
 sg13g2_nor4_1 _22173_ (.A(_04317_),
    .B(_04612_),
    .C(_04613_),
    .D(_04618_),
    .Y(_04619_));
 sg13g2_or3_1 _22174_ (.A(_11487_),
    .B(_11599_),
    .C(net157),
    .X(_04620_));
 sg13g2_nand2_1 _22175_ (.Y(_04621_),
    .A(_04145_),
    .B(_04620_));
 sg13g2_o21ai_1 _22176_ (.B1(_04621_),
    .Y(_04622_),
    .A1(_04218_),
    .A2(_04619_));
 sg13g2_o21ai_1 _22177_ (.B1(_04622_),
    .Y(_04623_),
    .A1(net134),
    .A2(_04303_));
 sg13g2_nand2_1 _22178_ (.Y(_04624_),
    .A(net125),
    .B(net126));
 sg13g2_a21oi_1 _22179_ (.A1(net225),
    .A2(net160),
    .Y(_04625_),
    .B1(net122));
 sg13g2_a22oi_1 _22180_ (.Y(_04626_),
    .B1(net155),
    .B2(net124),
    .A2(net162),
    .A1(net127));
 sg13g2_nand3_1 _22181_ (.B(_04625_),
    .C(_04626_),
    .A(_04624_),
    .Y(_04627_));
 sg13g2_and2_1 _22182_ (.A(_09889_),
    .B(_04537_),
    .X(_04628_));
 sg13g2_inv_1 _22183_ (.Y(_04629_),
    .A(_09001_));
 sg13g2_o21ai_1 _22184_ (.B1(_04143_),
    .Y(_04630_),
    .A1(_04629_),
    .A2(net141));
 sg13g2_a21oi_1 _22185_ (.A1(_04627_),
    .A2(_04628_),
    .Y(_04631_),
    .B1(_04630_));
 sg13g2_nand2_1 _22186_ (.Y(_04632_),
    .A(_11614_),
    .B(_03668_));
 sg13g2_mux2_1 _22187_ (.A0(_09101_),
    .A1(net1046),
    .S(_04632_),
    .X(_04633_));
 sg13g2_nand2b_1 _22188_ (.Y(_04634_),
    .B(_11675_),
    .A_N(_03668_));
 sg13g2_o21ai_1 _22189_ (.B1(_04634_),
    .Y(_04635_),
    .A1(net1033),
    .A2(_04633_));
 sg13g2_a22oi_1 _22190_ (.Y(_04636_),
    .B1(_03799_),
    .B2(_03802_),
    .A2(_03793_),
    .A1(_03788_));
 sg13g2_buf_1 _22191_ (.A(_04636_),
    .X(_04637_));
 sg13g2_and2_1 _22192_ (.A(_04634_),
    .B(_04632_),
    .X(_04638_));
 sg13g2_xnor2_1 _22193_ (.Y(_04639_),
    .A(_04637_),
    .B(_04638_));
 sg13g2_xor2_1 _22194_ (.B(_04638_),
    .A(_03706_),
    .X(_04640_));
 sg13g2_a22oi_1 _22195_ (.Y(_04641_),
    .B1(_04640_),
    .B2(_04237_),
    .A2(_04639_),
    .A1(_09180_));
 sg13g2_nand4_1 _22196_ (.B(_04631_),
    .C(_04635_),
    .A(_04623_),
    .Y(_04642_),
    .D(_04641_));
 sg13g2_o21ai_1 _22197_ (.B1(_04642_),
    .Y(_04643_),
    .A1(_04143_),
    .A2(\cpu.ex.c_mult[5] ));
 sg13g2_buf_1 _22198_ (.A(_08829_),
    .X(_04644_));
 sg13g2_xnor2_1 _22199_ (.Y(_04645_),
    .A(_10981_),
    .B(_04340_));
 sg13g2_a22oi_1 _22200_ (.Y(_04646_),
    .B1(_04645_),
    .B2(_04345_),
    .A2(net61),
    .A1(net964));
 sg13g2_o21ai_1 _22201_ (.B1(_04646_),
    .Y(_00989_),
    .A1(_04141_),
    .A2(_04643_));
 sg13g2_nand2_1 _22202_ (.Y(_04647_),
    .A(_03671_),
    .B(_03658_));
 sg13g2_o21ai_1 _22203_ (.B1(_03807_),
    .Y(_04648_),
    .A1(_03813_),
    .A2(_04637_));
 sg13g2_xor2_1 _22204_ (.B(_04648_),
    .A(_04647_),
    .X(_04649_));
 sg13g2_nand2_1 _22205_ (.Y(_04650_),
    .A(_04289_),
    .B(_04290_));
 sg13g2_xnor2_1 _22206_ (.Y(_04651_),
    .A(_04650_),
    .B(_04647_));
 sg13g2_nand2_1 _22207_ (.Y(_04652_),
    .A(_03659_),
    .B(net129));
 sg13g2_a22oi_1 _22208_ (.Y(_04653_),
    .B1(_04186_),
    .B2(net166),
    .A2(_04177_),
    .A1(net138));
 sg13g2_nand2_1 _22209_ (.Y(_04654_),
    .A(net165),
    .B(_04174_));
 sg13g2_nand2_1 _22210_ (.Y(_04655_),
    .A(_03826_),
    .B(net156));
 sg13g2_a21oi_1 _22211_ (.A1(net130),
    .A2(net181),
    .Y(_04656_),
    .B1(_04152_));
 sg13g2_nand4_1 _22212_ (.B(_04654_),
    .C(_04655_),
    .A(_04653_),
    .Y(_04657_),
    .D(_04656_));
 sg13g2_nand2_1 _22213_ (.Y(_04658_),
    .A(net136),
    .B(_04158_));
 sg13g2_nand3_1 _22214_ (.B(_04454_),
    .C(_04658_),
    .A(_04357_),
    .Y(_04659_));
 sg13g2_o21ai_1 _22215_ (.B1(_04213_),
    .Y(_04660_),
    .A1(_04657_),
    .A2(_04659_));
 sg13g2_o21ai_1 _22216_ (.B1(_04145_),
    .Y(_04661_),
    .A1(net158),
    .A2(_04620_));
 sg13g2_nand2_1 _22217_ (.Y(_04662_),
    .A(_04660_),
    .B(_04661_));
 sg13g2_mux2_1 _22218_ (.A0(net1124),
    .A1(_09166_),
    .S(_03671_),
    .X(_04663_));
 sg13g2_o21ai_1 _22219_ (.B1(_03658_),
    .Y(_04664_),
    .A1(net1115),
    .A2(_04663_));
 sg13g2_a21oi_1 _22220_ (.A1(_09001_),
    .A2(_11470_),
    .Y(_04665_),
    .B1(_11534_));
 sg13g2_a22oi_1 _22221_ (.Y(_04666_),
    .B1(net156),
    .B2(net123),
    .A2(net180),
    .A1(net225));
 sg13g2_a22oi_1 _22222_ (.Y(_04667_),
    .B1(net179),
    .B2(_03699_),
    .A2(net181),
    .A1(_04228_));
 sg13g2_a21oi_1 _22223_ (.A1(net167),
    .A2(net162),
    .Y(_04668_),
    .B1(net161));
 sg13g2_nand3_1 _22224_ (.B(_04667_),
    .C(_04668_),
    .A(_04666_),
    .Y(_04669_));
 sg13g2_nand3_1 _22225_ (.B(_04601_),
    .C(_04669_),
    .A(_09889_),
    .Y(_04670_));
 sg13g2_nand3_1 _22226_ (.B(_04665_),
    .C(_04670_),
    .A(_04664_),
    .Y(_04671_));
 sg13g2_a221oi_1 _22227_ (.B2(_04662_),
    .C1(_04671_),
    .B1(_04652_),
    .A1(_04237_),
    .Y(_04672_),
    .A2(_04651_));
 sg13g2_o21ai_1 _22228_ (.B1(_04672_),
    .Y(_04673_),
    .A1(net832),
    .A2(_04649_));
 sg13g2_o21ai_1 _22229_ (.B1(_04673_),
    .Y(_04674_),
    .A1(net278),
    .A2(\cpu.ex.c_mult[6] ));
 sg13g2_buf_1 _22230_ (.A(_08777_),
    .X(_04675_));
 sg13g2_nand2_1 _22231_ (.Y(_04676_),
    .A(_08829_),
    .B(_04340_));
 sg13g2_xnor2_1 _22232_ (.Y(_04677_),
    .A(_03651_),
    .B(_04676_));
 sg13g2_a22oi_1 _22233_ (.Y(_04678_),
    .B1(_04677_),
    .B2(_04345_),
    .A2(_04268_),
    .A1(net963));
 sg13g2_o21ai_1 _22234_ (.B1(_04678_),
    .Y(_00990_),
    .A1(_04141_),
    .A2(_04674_));
 sg13g2_nand2_1 _22235_ (.Y(_04679_),
    .A(_03671_),
    .B(_04293_));
 sg13g2_xnor2_1 _22236_ (.Y(_04680_),
    .A(_04679_),
    .B(_04295_));
 sg13g2_and3_1 _22237_ (.X(_04681_),
    .A(_03805_),
    .B(_04637_),
    .C(_03807_));
 sg13g2_nor2b_1 _22238_ (.A(_04681_),
    .B_N(_03815_),
    .Y(_04682_));
 sg13g2_xor2_1 _22239_ (.B(_04295_),
    .A(_04682_),
    .X(_04683_));
 sg13g2_nor2_1 _22240_ (.A(_08256_),
    .B(net154),
    .Y(_04684_));
 sg13g2_nor3_1 _22241_ (.A(_03773_),
    .B(_04310_),
    .C(_04684_),
    .Y(_04685_));
 sg13g2_a221oi_1 _22242_ (.B2(net132),
    .C1(_04685_),
    .B1(net126),
    .A1(net136),
    .Y(_04686_),
    .A2(net159));
 sg13g2_a221oi_1 _22243_ (.B2(_04301_),
    .C1(_04476_),
    .B1(net160),
    .A1(net137),
    .Y(_04687_),
    .A2(_04159_));
 sg13g2_nand3_1 _22244_ (.B(_04686_),
    .C(_04687_),
    .A(_04401_),
    .Y(_04688_));
 sg13g2_nand2_1 _22245_ (.Y(_04689_),
    .A(_03714_),
    .B(net122));
 sg13g2_nand3_1 _22246_ (.B(_04688_),
    .C(_04689_),
    .A(_04213_),
    .Y(_04690_));
 sg13g2_o21ai_1 _22247_ (.B1(net1032),
    .Y(_04691_),
    .A1(_04163_),
    .A2(_04303_));
 sg13g2_a22oi_1 _22248_ (.Y(_04692_),
    .B1(net155),
    .B2(_04322_),
    .A2(net159),
    .A1(_04324_));
 sg13g2_nand2_1 _22249_ (.Y(_04693_),
    .A(net198),
    .B(net182));
 sg13g2_a21oi_1 _22250_ (.A1(_04316_),
    .A2(net160),
    .Y(_04694_),
    .B1(_04153_));
 sg13g2_nand4_1 _22251_ (.B(_04692_),
    .C(_04693_),
    .A(_04546_),
    .Y(_04695_),
    .D(_04694_));
 sg13g2_nand2b_1 _22252_ (.Y(_04696_),
    .B(_04695_),
    .A_N(_04691_));
 sg13g2_mux2_1 _22253_ (.A0(_09101_),
    .A1(_09167_),
    .S(_03650_),
    .X(_04697_));
 sg13g2_o21ai_1 _22254_ (.B1(_03660_),
    .Y(_04698_),
    .A1(net1033),
    .A2(_04697_));
 sg13g2_a21oi_1 _22255_ (.A1(net1048),
    .A2(_11442_),
    .Y(_04699_),
    .B1(_04246_));
 sg13g2_nand4_1 _22256_ (.B(_04696_),
    .C(_04698_),
    .A(_04690_),
    .Y(_04700_),
    .D(_04699_));
 sg13g2_a21oi_1 _22257_ (.A1(net1045),
    .A2(_04683_),
    .Y(_04701_),
    .B1(_04700_));
 sg13g2_o21ai_1 _22258_ (.B1(_04701_),
    .Y(_04702_),
    .A1(_04224_),
    .A2(_04680_));
 sg13g2_o21ai_1 _22259_ (.B1(_04702_),
    .Y(_04703_),
    .A1(net278),
    .A2(\cpu.ex.c_mult[7] ));
 sg13g2_buf_1 _22260_ (.A(_08797_),
    .X(_04704_));
 sg13g2_nand3_1 _22261_ (.B(_08777_),
    .C(_04340_),
    .A(_08829_),
    .Y(_04705_));
 sg13g2_xnor2_1 _22262_ (.Y(_04706_),
    .A(_03645_),
    .B(_04705_));
 sg13g2_a22oi_1 _22263_ (.Y(_04707_),
    .B1(_04706_),
    .B2(net81),
    .A2(net61),
    .A1(net962));
 sg13g2_o21ai_1 _22264_ (.B1(_04707_),
    .Y(_00991_),
    .A1(_04140_),
    .A2(_04703_));
 sg13g2_nor3_1 _22265_ (.A(_04288_),
    .B(_04297_),
    .C(_04299_),
    .Y(_04708_));
 sg13g2_nand2_1 _22266_ (.Y(_04709_),
    .A(_11719_),
    .B(net135));
 sg13g2_and2_1 _22267_ (.A(_03719_),
    .B(_04709_),
    .X(_04710_));
 sg13g2_xor2_1 _22268_ (.B(_04710_),
    .A(_03818_),
    .X(_04711_));
 sg13g2_a22oi_1 _22269_ (.Y(_04712_),
    .B1(net154),
    .B2(_04230_),
    .A2(net199),
    .A1(_04228_));
 sg13g2_a22oi_1 _22270_ (.Y(_04713_),
    .B1(net155),
    .B2(net123),
    .A2(net160),
    .A1(net167));
 sg13g2_a22oi_1 _22271_ (.Y(_04714_),
    .B1(net162),
    .B2(net131),
    .A2(net180),
    .A1(net127));
 sg13g2_nand4_1 _22272_ (.B(_04712_),
    .C(_04713_),
    .A(_04598_),
    .Y(_04715_),
    .D(_04714_));
 sg13g2_nand3_1 _22273_ (.B(_04652_),
    .C(_04715_),
    .A(net1032),
    .Y(_04716_));
 sg13g2_nand2_1 _22274_ (.Y(_04717_),
    .A(net1073),
    .B(_04311_));
 sg13g2_a22oi_1 _22275_ (.Y(_04718_),
    .B1(_04162_),
    .B2(net136),
    .A2(_04175_),
    .A1(net137));
 sg13g2_a22oi_1 _22276_ (.Y(_04719_),
    .B1(_04207_),
    .B2(net133),
    .A2(_04158_),
    .A1(net138));
 sg13g2_nand2_1 _22277_ (.Y(_04720_),
    .A(_04449_),
    .B(_04719_));
 sg13g2_a21oi_1 _22278_ (.A1(net128),
    .A2(net155),
    .Y(_04721_),
    .B1(_04720_));
 sg13g2_nand3_1 _22279_ (.B(_04718_),
    .C(_04721_),
    .A(_04717_),
    .Y(_04722_));
 sg13g2_nand2_1 _22280_ (.Y(_04723_),
    .A(_03720_),
    .B(net122));
 sg13g2_nand3_1 _22281_ (.B(_04722_),
    .C(_04723_),
    .A(_04213_),
    .Y(_04724_));
 sg13g2_nand2_1 _22282_ (.Y(_04725_),
    .A(net1048),
    .B(_03784_));
 sg13g2_mux2_1 _22283_ (.A0(net1124),
    .A1(_09166_),
    .S(_04709_),
    .X(_04726_));
 sg13g2_o21ai_1 _22284_ (.B1(_03719_),
    .Y(_04727_),
    .A1(_09886_),
    .A2(_04726_));
 sg13g2_nand4_1 _22285_ (.B(_04724_),
    .C(_04725_),
    .A(_04716_),
    .Y(_04728_),
    .D(_04727_));
 sg13g2_a21oi_1 _22286_ (.A1(_09181_),
    .A2(_04711_),
    .Y(_04729_),
    .B1(_04728_));
 sg13g2_nand2_1 _22287_ (.Y(_04730_),
    .A(_03674_),
    .B(_03708_));
 sg13g2_xor2_1 _22288_ (.B(_04710_),
    .A(_04730_),
    .X(_04731_));
 sg13g2_a22oi_1 _22289_ (.Y(_04732_),
    .B1(_04731_),
    .B2(_04288_),
    .A2(_04729_),
    .A1(_04708_));
 sg13g2_mux2_1 _22290_ (.A0(\cpu.ex.c_mult[8] ),
    .A1(_04732_),
    .S(net278),
    .X(_04733_));
 sg13g2_nand2b_1 _22291_ (.Y(_04734_),
    .B(_04733_),
    .A_N(_04140_));
 sg13g2_xnor2_1 _22292_ (.Y(_04735_),
    .A(_10737_),
    .B(_04341_));
 sg13g2_a22oi_1 _22293_ (.Y(_04736_),
    .B1(_04735_),
    .B2(net81),
    .A2(_04268_),
    .A1(\cpu.ex.pc[8] ));
 sg13g2_nand2_1 _22294_ (.Y(_00992_),
    .A(_04734_),
    .B(_04736_));
 sg13g2_a221oi_1 _22295_ (.B2(_11714_),
    .C1(_04270_),
    .B1(_11727_),
    .A1(\cpu.ex.r_mult[9] ),
    .Y(_04737_),
    .A2(net411));
 sg13g2_and2_1 _22296_ (.A(_03721_),
    .B(_03712_),
    .X(_04738_));
 sg13g2_nor2_1 _22297_ (.A(net190),
    .B(net135),
    .Y(_04739_));
 sg13g2_a21oi_1 _22298_ (.A1(_03818_),
    .A2(_03828_),
    .Y(_04740_),
    .B1(_04739_));
 sg13g2_xnor2_1 _22299_ (.Y(_04741_),
    .A(_04738_),
    .B(_04740_));
 sg13g2_nand2_1 _22300_ (.Y(_04742_),
    .A(net1045),
    .B(_04741_));
 sg13g2_nand3_1 _22301_ (.B(_03674_),
    .C(_03708_),
    .A(net135),
    .Y(_04743_));
 sg13g2_a21oi_1 _22302_ (.A1(_03674_),
    .A2(_03708_),
    .Y(_04744_),
    .B1(net135));
 sg13g2_a21oi_1 _22303_ (.A1(_11667_),
    .A2(_04743_),
    .Y(_04745_),
    .B1(_04744_));
 sg13g2_xnor2_1 _22304_ (.Y(_04746_),
    .A(_04745_),
    .B(_04738_));
 sg13g2_nand2b_1 _22305_ (.Y(_04747_),
    .B(_04288_),
    .A_N(_04746_));
 sg13g2_a22oi_1 _22306_ (.Y(_04748_),
    .B1(_04207_),
    .B2(_04196_),
    .A2(_04148_),
    .A1(_03753_));
 sg13g2_a22oi_1 _22307_ (.Y(_04749_),
    .B1(_04191_),
    .B2(net164),
    .A2(_04174_),
    .A1(_03642_));
 sg13g2_a21oi_1 _22308_ (.A1(net166),
    .A2(net181),
    .Y(_04750_),
    .B1(_04151_));
 sg13g2_nand3_1 _22309_ (.B(_04749_),
    .C(_04750_),
    .A(_04748_),
    .Y(_04751_));
 sg13g2_and2_1 _22310_ (.A(_03643_),
    .B(net199),
    .X(_04752_));
 sg13g2_or3_1 _22311_ (.A(_04311_),
    .B(_04752_),
    .C(_04751_),
    .X(_04753_));
 sg13g2_a22oi_1 _22312_ (.Y(_04754_),
    .B1(_04753_),
    .B2(net1073),
    .A2(_04751_),
    .A1(_09880_));
 sg13g2_inv_1 _22313_ (.Y(_04755_),
    .A(_04754_));
 sg13g2_a22oi_1 _22314_ (.Y(_04756_),
    .B1(_04186_),
    .B2(_04228_),
    .A2(net180),
    .A1(net167));
 sg13g2_a22oi_1 _22315_ (.Y(_04757_),
    .B1(_04359_),
    .B2(_04230_),
    .A2(net181),
    .A1(_03801_));
 sg13g2_nand3_1 _22316_ (.B(_04756_),
    .C(_04757_),
    .A(_04541_),
    .Y(_04758_));
 sg13g2_a221oi_1 _22317_ (.B2(net131),
    .C1(_04612_),
    .B1(net179),
    .A1(_03699_),
    .Y(_04759_),
    .A2(net199));
 sg13g2_nand2b_1 _22318_ (.Y(_04760_),
    .B(_04759_),
    .A_N(_04758_));
 sg13g2_nand3_1 _22319_ (.B(_04689_),
    .C(_04760_),
    .A(_09889_),
    .Y(_04761_));
 sg13g2_mux2_1 _22320_ (.A0(net1124),
    .A1(_09166_),
    .S(_03712_),
    .X(_04762_));
 sg13g2_o21ai_1 _22321_ (.B1(_03721_),
    .Y(_04763_),
    .A1(net1115),
    .A2(_04762_));
 sg13g2_nand2_1 _22322_ (.Y(_04764_),
    .A(_09002_),
    .B(net238));
 sg13g2_nand3_1 _22323_ (.B(_04763_),
    .C(_04764_),
    .A(_04761_),
    .Y(_04765_));
 sg13g2_a21oi_1 _22324_ (.A1(_04330_),
    .A2(_04755_),
    .Y(_04766_),
    .B1(_04765_));
 sg13g2_and4_1 _22325_ (.A(_04300_),
    .B(_04742_),
    .C(_04747_),
    .D(_04766_),
    .X(_04767_));
 sg13g2_a21o_1 _22326_ (.A2(_04737_),
    .A1(_11726_),
    .B1(_04767_),
    .X(_04768_));
 sg13g2_xnor2_1 _22327_ (.Y(_04769_),
    .A(_11109_),
    .B(_04342_));
 sg13g2_a22oi_1 _22328_ (.Y(_04770_),
    .B1(_04769_),
    .B2(net81),
    .A2(_04267_),
    .A1(_08786_));
 sg13g2_o21ai_1 _22329_ (.B1(_04770_),
    .Y(_00993_),
    .A1(_04140_),
    .A2(_04768_));
 sg13g2_nand3_1 _22330_ (.B(_03818_),
    .C(_03828_),
    .A(_03824_),
    .Y(_04771_));
 sg13g2_nand2_1 _22331_ (.Y(_04772_),
    .A(_04279_),
    .B(_04771_));
 sg13g2_nand2_1 _22332_ (.Y(_04773_),
    .A(_11731_),
    .B(_04180_));
 sg13g2_nand2_1 _22333_ (.Y(_04774_),
    .A(_04773_),
    .B(_03734_));
 sg13g2_xnor2_1 _22334_ (.Y(_04775_),
    .A(_04772_),
    .B(_04774_));
 sg13g2_and2_1 _22335_ (.A(_09181_),
    .B(_04775_),
    .X(_04776_));
 sg13g2_a221oi_1 _22336_ (.B2(net134),
    .C1(_04214_),
    .B1(_04307_),
    .A1(net127),
    .Y(_04777_),
    .A2(net154));
 sg13g2_a22oi_1 _22337_ (.Y(_04778_),
    .B1(_04177_),
    .B2(net124),
    .A2(net182),
    .A1(net125));
 sg13g2_nand2_1 _22338_ (.Y(_04779_),
    .A(net131),
    .B(net181));
 sg13g2_nand2_1 _22339_ (.Y(_04780_),
    .A(_04599_),
    .B(_04779_));
 sg13g2_a221oi_1 _22340_ (.B2(net198),
    .C1(_04780_),
    .B1(net158),
    .A1(net123),
    .Y(_04781_),
    .A2(net159));
 sg13g2_nand4_1 _22341_ (.B(_04777_),
    .C(_04778_),
    .A(_04655_),
    .Y(_04782_),
    .D(_04781_));
 sg13g2_and2_1 _22342_ (.A(_09890_),
    .B(_04723_),
    .X(_04783_));
 sg13g2_nand2_1 _22343_ (.Y(_04784_),
    .A(_04301_),
    .B(_04208_));
 sg13g2_a21oi_1 _22344_ (.A1(_03643_),
    .A2(_04161_),
    .Y(_04785_),
    .B1(_04152_));
 sg13g2_a22oi_1 _22345_ (.Y(_04786_),
    .B1(_04192_),
    .B2(net166),
    .A2(net162),
    .A1(net136));
 sg13g2_nand3_1 _22346_ (.B(_04785_),
    .C(_04786_),
    .A(_04784_),
    .Y(_04787_));
 sg13g2_nand2_1 _22347_ (.Y(_04788_),
    .A(_04213_),
    .B(_04787_));
 sg13g2_o21ai_1 _22348_ (.B1(_04145_),
    .Y(_04789_),
    .A1(net159),
    .A2(_04159_));
 sg13g2_nand3_1 _22349_ (.B(_04788_),
    .C(_04789_),
    .A(_04717_),
    .Y(_04790_));
 sg13g2_mux2_1 _22350_ (.A0(_09100_),
    .A1(_09166_),
    .S(_04773_),
    .X(_04791_));
 sg13g2_o21ai_1 _22351_ (.B1(_03734_),
    .Y(_04792_),
    .A1(net1115),
    .A2(_04791_));
 sg13g2_o21ai_1 _22352_ (.B1(_04792_),
    .Y(_04793_),
    .A1(_04629_),
    .A2(_11563_));
 sg13g2_a221oi_1 _22353_ (.B2(_04370_),
    .C1(_04793_),
    .B1(_04790_),
    .A1(_04782_),
    .Y(_04794_),
    .A2(_04783_));
 sg13g2_nand2_1 _22354_ (.Y(_04795_),
    .A(_04708_),
    .B(_04794_));
 sg13g2_xor2_1 _22355_ (.B(_04774_),
    .A(_04284_),
    .X(_04796_));
 sg13g2_nand2_1 _22356_ (.Y(_04797_),
    .A(_04288_),
    .B(_04796_));
 sg13g2_o21ai_1 _22357_ (.B1(_04797_),
    .Y(_04798_),
    .A1(_04776_),
    .A2(_04795_));
 sg13g2_nand2_1 _22358_ (.Y(_04799_),
    .A(_04270_),
    .B(_04798_));
 sg13g2_o21ai_1 _22359_ (.B1(_04799_),
    .Y(_04800_),
    .A1(net278),
    .A2(\cpu.ex.c_mult[10] ));
 sg13g2_buf_1 _22360_ (.A(_08807_),
    .X(_04801_));
 sg13g2_nand2_1 _22361_ (.Y(_04802_),
    .A(_08786_),
    .B(_04342_));
 sg13g2_xor2_1 _22362_ (.B(_04802_),
    .A(_10738_),
    .X(_04803_));
 sg13g2_a22oi_1 _22363_ (.Y(_04804_),
    .B1(_04803_),
    .B2(net96),
    .A2(_04267_),
    .A1(net961));
 sg13g2_o21ai_1 _22364_ (.B1(_04804_),
    .Y(_00994_),
    .A1(_04140_),
    .A2(_04800_));
 sg13g2_mux2_1 _22365_ (.A0(\cpu.dec.r_set_cc ),
    .A1(_10223_),
    .S(_03635_),
    .X(_00997_));
 sg13g2_buf_1 _22366_ (.A(_00254_),
    .X(_04805_));
 sg13g2_nor4_1 _22367_ (.A(net1111),
    .B(net1110),
    .C(_04805_),
    .D(_03575_),
    .Y(_04806_));
 sg13g2_buf_2 _22368_ (.A(_04806_),
    .X(_04807_));
 sg13g2_buf_1 _22369_ (.A(_04807_),
    .X(_04808_));
 sg13g2_mux2_1 _22370_ (.A0(_10539_),
    .A1(_03589_),
    .S(_04808_),
    .X(_00998_));
 sg13g2_buf_1 _22371_ (.A(net967),
    .X(_04809_));
 sg13g2_mux2_1 _22372_ (.A0(_10395_),
    .A1(_04809_),
    .S(_04808_),
    .X(_00999_));
 sg13g2_mux2_1 _22373_ (.A0(_10373_),
    .A1(net455),
    .S(net511),
    .X(_01000_));
 sg13g2_mux2_1 _22374_ (.A0(\cpu.ex.r_sp[13] ),
    .A1(net454),
    .S(net511),
    .X(_01001_));
 sg13g2_buf_1 _22375_ (.A(net520),
    .X(_04810_));
 sg13g2_mux2_1 _22376_ (.A0(_10825_),
    .A1(_04810_),
    .S(net511),
    .X(_01002_));
 sg13g2_mux2_1 _22377_ (.A0(_10937_),
    .A1(net720),
    .S(net511),
    .X(_01003_));
 sg13g2_mux2_1 _22378_ (.A0(_10482_),
    .A1(_03591_),
    .S(net511),
    .X(_01004_));
 sg13g2_mux2_1 _22379_ (.A0(_10436_),
    .A1(net518),
    .S(net511),
    .X(_01005_));
 sg13g2_mux2_1 _22380_ (.A0(_10871_),
    .A1(net517),
    .S(net511),
    .X(_01006_));
 sg13g2_mux2_1 _22381_ (.A0(_10898_),
    .A1(net593),
    .S(_04807_),
    .X(_01007_));
 sg13g2_mux2_1 _22382_ (.A0(_10788_),
    .A1(net723),
    .S(_04807_),
    .X(_01008_));
 sg13g2_nand2_1 _22383_ (.Y(_04811_),
    .A(net841),
    .B(_04807_));
 sg13g2_o21ai_1 _22384_ (.B1(_04811_),
    .Y(_01009_),
    .A1(_10953_),
    .A2(net511));
 sg13g2_buf_1 _22385_ (.A(net845),
    .X(_04812_));
 sg13g2_mux2_1 _22386_ (.A0(_10682_),
    .A1(_04812_),
    .S(_04807_),
    .X(_01010_));
 sg13g2_mux2_1 _22387_ (.A0(_11101_),
    .A1(net837),
    .S(_04807_),
    .X(_01011_));
 sg13g2_mux2_1 _22388_ (.A0(_10716_),
    .A1(net836),
    .S(_04807_),
    .X(_01012_));
 sg13g2_or2_1 _22389_ (.X(_04813_),
    .B(_03575_),
    .A(_10228_));
 sg13g2_buf_1 _22390_ (.A(_04813_),
    .X(_04814_));
 sg13g2_buf_1 _22391_ (.A(_04814_),
    .X(_04815_));
 sg13g2_nor2b_1 _22392_ (.A(_04805_),
    .B_N(net920),
    .Y(_04816_));
 sg13g2_nand2_1 _22393_ (.Y(_04817_),
    .A(_03573_),
    .B(_04816_));
 sg13g2_and2_1 _22394_ (.A(_08621_),
    .B(net1110),
    .X(_04818_));
 sg13g2_a21oi_1 _22395_ (.A1(_03576_),
    .A2(\cpu.ex.r_wb_swapsp ),
    .Y(_04819_),
    .B1(_04818_));
 sg13g2_or4_1 _22396_ (.A(net1111),
    .B(_04805_),
    .C(_03575_),
    .D(_04819_),
    .X(_04820_));
 sg13g2_buf_1 _22397_ (.A(_04820_),
    .X(_04821_));
 sg13g2_buf_1 _22398_ (.A(_04821_),
    .X(_04822_));
 sg13g2_nand2_1 _22399_ (.Y(_04823_),
    .A(\cpu.ex.r_stmp[0] ),
    .B(net449));
 sg13g2_o21ai_1 _22400_ (.B1(_04823_),
    .Y(_01013_),
    .A1(net510),
    .A2(_04817_));
 sg13g2_mux2_1 _22401_ (.A0(net1104),
    .A1(_10716_),
    .S(net510),
    .X(_04824_));
 sg13g2_buf_1 _22402_ (.A(_04821_),
    .X(_04825_));
 sg13g2_mux2_1 _22403_ (.A0(_04824_),
    .A1(\cpu.ex.r_stmp[10] ),
    .S(net448),
    .X(_01014_));
 sg13g2_mux2_1 _22404_ (.A0(net1107),
    .A1(_10395_),
    .S(_04815_),
    .X(_04826_));
 sg13g2_mux2_1 _22405_ (.A0(_04826_),
    .A1(\cpu.ex.r_stmp[11] ),
    .S(net448),
    .X(_01015_));
 sg13g2_buf_1 _22406_ (.A(_04814_),
    .X(_04827_));
 sg13g2_mux2_1 _22407_ (.A0(net620),
    .A1(_10373_),
    .S(net509),
    .X(_04828_));
 sg13g2_mux2_1 _22408_ (.A0(_04828_),
    .A1(\cpu.ex.r_stmp[12] ),
    .S(net448),
    .X(_01016_));
 sg13g2_mux2_1 _22409_ (.A0(net614),
    .A1(\cpu.ex.r_sp[13] ),
    .S(net509),
    .X(_04829_));
 sg13g2_mux2_1 _22410_ (.A0(_04829_),
    .A1(\cpu.ex.r_stmp[13] ),
    .S(net449),
    .X(_01017_));
 sg13g2_mux2_1 _22411_ (.A0(net605),
    .A1(_10825_),
    .S(net509),
    .X(_04830_));
 sg13g2_mux2_1 _22412_ (.A0(_04830_),
    .A1(\cpu.ex.r_stmp[14] ),
    .S(net449),
    .X(_01018_));
 sg13g2_nor2_1 _22413_ (.A(net676),
    .B(net509),
    .Y(_04831_));
 sg13g2_a21oi_1 _22414_ (.A1(_10937_),
    .A2(net510),
    .Y(_04832_),
    .B1(_04831_));
 sg13g2_nand2_1 _22415_ (.Y(_04833_),
    .A(\cpu.ex.r_stmp[15] ),
    .B(_04822_));
 sg13g2_o21ai_1 _22416_ (.B1(_04833_),
    .Y(_01019_),
    .A1(net448),
    .A2(_04832_));
 sg13g2_nor2_1 _22417_ (.A(_10180_),
    .B(net509),
    .Y(_04834_));
 sg13g2_a21oi_1 _22418_ (.A1(_10539_),
    .A2(_04815_),
    .Y(_04835_),
    .B1(_04834_));
 sg13g2_nand2_1 _22419_ (.Y(_04836_),
    .A(\cpu.ex.r_stmp[1] ),
    .B(net449));
 sg13g2_o21ai_1 _22420_ (.B1(_04836_),
    .Y(_01020_),
    .A1(net448),
    .A2(_04835_));
 sg13g2_nor2_1 _22421_ (.A(_09524_),
    .B(net509),
    .Y(_04837_));
 sg13g2_a21oi_1 _22422_ (.A1(_10482_),
    .A2(net510),
    .Y(_04838_),
    .B1(_04837_));
 sg13g2_nand2_1 _22423_ (.Y(_04839_),
    .A(\cpu.ex.r_stmp[2] ),
    .B(net449));
 sg13g2_o21ai_1 _22424_ (.B1(_04839_),
    .Y(_01021_),
    .A1(_04825_),
    .A2(_04838_));
 sg13g2_nor2_1 _22425_ (.A(_09342_),
    .B(net509),
    .Y(_04840_));
 sg13g2_a21oi_1 _22426_ (.A1(_10436_),
    .A2(net510),
    .Y(_04841_),
    .B1(_04840_));
 sg13g2_nand2_1 _22427_ (.Y(_04842_),
    .A(\cpu.ex.r_stmp[3] ),
    .B(net449));
 sg13g2_o21ai_1 _22428_ (.B1(_04842_),
    .Y(_01022_),
    .A1(_04825_),
    .A2(_04841_));
 sg13g2_nor2_1 _22429_ (.A(net650),
    .B(_04814_),
    .Y(_04843_));
 sg13g2_a21oi_1 _22430_ (.A1(_10871_),
    .A2(net510),
    .Y(_04844_),
    .B1(_04843_));
 sg13g2_nand2_1 _22431_ (.Y(_04845_),
    .A(\cpu.ex.r_stmp[4] ),
    .B(_04821_));
 sg13g2_o21ai_1 _22432_ (.B1(_04845_),
    .Y(_01023_),
    .A1(net448),
    .A2(_04844_));
 sg13g2_nor2_1 _22433_ (.A(net730),
    .B(_04814_),
    .Y(_04846_));
 sg13g2_a21oi_1 _22434_ (.A1(_10898_),
    .A2(net510),
    .Y(_04847_),
    .B1(_04846_));
 sg13g2_nand2_1 _22435_ (.Y(_04848_),
    .A(\cpu.ex.r_stmp[5] ),
    .B(_04821_));
 sg13g2_o21ai_1 _22436_ (.B1(_04848_),
    .Y(_01024_),
    .A1(net448),
    .A2(_04847_));
 sg13g2_mux2_1 _22437_ (.A0(net1028),
    .A1(_10788_),
    .S(net509),
    .X(_04849_));
 sg13g2_mux2_1 _22438_ (.A0(_04849_),
    .A1(\cpu.ex.r_stmp[6] ),
    .S(net449),
    .X(_01025_));
 sg13g2_nor2_1 _22439_ (.A(_02979_),
    .B(_04814_),
    .Y(_04850_));
 sg13g2_a21oi_1 _22440_ (.A1(\cpu.ex.r_sp[7] ),
    .A2(net510),
    .Y(_04851_),
    .B1(_04850_));
 sg13g2_nand2_1 _22441_ (.Y(_04852_),
    .A(\cpu.ex.r_stmp[7] ),
    .B(_04821_));
 sg13g2_o21ai_1 _22442_ (.B1(_04852_),
    .Y(_01026_),
    .A1(net448),
    .A2(_04851_));
 sg13g2_mux2_1 _22443_ (.A0(net1043),
    .A1(_10682_),
    .S(_04827_),
    .X(_04853_));
 sg13g2_mux2_1 _22444_ (.A0(_04853_),
    .A1(\cpu.ex.r_stmp[8] ),
    .S(net449),
    .X(_01027_));
 sg13g2_mux2_1 _22445_ (.A0(_11085_),
    .A1(_11101_),
    .S(_04827_),
    .X(_04854_));
 sg13g2_mux2_1 _22446_ (.A0(_04854_),
    .A1(\cpu.ex.r_stmp[9] ),
    .S(_04822_),
    .X(_01028_));
 sg13g2_nand2_1 _22447_ (.Y(_04855_),
    .A(_11520_),
    .B(net331));
 sg13g2_a221oi_1 _22448_ (.B2(net58),
    .C1(_04855_),
    .B1(_11480_),
    .A1(_11515_),
    .Y(_04856_),
    .A2(_11511_));
 sg13g2_buf_1 _22449_ (.A(_04856_),
    .X(_04857_));
 sg13g2_buf_1 _22450_ (.A(_11528_),
    .X(_04858_));
 sg13g2_buf_1 _22451_ (.A(net584),
    .X(_04859_));
 sg13g2_buf_1 _22452_ (.A(_04251_),
    .X(_04860_));
 sg13g2_inv_1 _22453_ (.Y(_04861_),
    .A(net124));
 sg13g2_a22oi_1 _22454_ (.Y(_04862_),
    .B1(net137),
    .B2(_04171_),
    .A2(net114),
    .A1(_11019_));
 sg13g2_nand2_1 _22455_ (.Y(_04863_),
    .A(net123),
    .B(net179));
 sg13g2_a22oi_1 _22456_ (.Y(_04864_),
    .B1(_04359_),
    .B2(net132),
    .A2(_04194_),
    .A1(net133));
 sg13g2_a22oi_1 _22457_ (.Y(_04865_),
    .B1(_04202_),
    .B2(_03753_),
    .A2(_04148_),
    .A1(_03682_));
 sg13g2_nand4_1 _22458_ (.B(_04779_),
    .C(_04864_),
    .A(_04863_),
    .Y(_04866_),
    .D(_04865_));
 sg13g2_a221oi_1 _22459_ (.B2(net136),
    .C1(_04866_),
    .B1(_04205_),
    .A1(_04155_),
    .Y(_04867_),
    .A2(net154));
 sg13g2_o21ai_1 _22460_ (.B1(_04867_),
    .Y(_04868_),
    .A1(_04518_),
    .A2(_04862_));
 sg13g2_nand2_1 _22461_ (.Y(_04869_),
    .A(_04196_),
    .B(net157));
 sg13g2_nand4_1 _22462_ (.B(_04455_),
    .C(_04585_),
    .A(_04365_),
    .Y(_04870_),
    .D(_04869_));
 sg13g2_o21ai_1 _22463_ (.B1(_04213_),
    .Y(_04871_),
    .A1(_04868_),
    .A2(_04870_));
 sg13g2_nand2_1 _22464_ (.Y(_04872_),
    .A(_11487_),
    .B(_04145_));
 sg13g2_a22oi_1 _22465_ (.Y(_04873_),
    .B1(_04871_),
    .B2(_04872_),
    .A2(net129),
    .A1(_04861_));
 sg13g2_nand2_1 _22466_ (.Y(_04874_),
    .A(_04220_),
    .B(_04224_));
 sg13g2_o21ai_1 _22467_ (.B1(net198),
    .Y(_04875_),
    .A1(net1033),
    .A2(_04874_));
 sg13g2_nand2b_1 _22468_ (.Y(_04876_),
    .B(_03693_),
    .A_N(net1047));
 sg13g2_or2_1 _22469_ (.X(_04877_),
    .B(_04874_),
    .A(net198));
 sg13g2_a21oi_1 _22470_ (.A1(_04876_),
    .A2(_04877_),
    .Y(_04878_),
    .B1(net1033));
 sg13g2_a21oi_1 _22471_ (.A1(_11510_),
    .A2(_04875_),
    .Y(_04879_),
    .B1(_04878_));
 sg13g2_o21ai_1 _22472_ (.B1(_04143_),
    .Y(_04880_),
    .A1(_04629_),
    .A2(_11667_));
 sg13g2_nor3_2 _22473_ (.A(_04873_),
    .B(_04879_),
    .C(_04880_),
    .Y(_04881_));
 sg13g2_or4_1 _22474_ (.A(net508),
    .B(_11540_),
    .C(net197),
    .D(_04881_),
    .X(_04882_));
 sg13g2_nand2_1 _22475_ (.Y(_04883_),
    .A(net1060),
    .B(_11544_));
 sg13g2_buf_1 _22476_ (.A(_04883_),
    .X(_04884_));
 sg13g2_buf_2 _22477_ (.A(_04884_),
    .X(_04885_));
 sg13g2_nand2b_1 _22478_ (.Y(_04886_),
    .B(net1042),
    .A_N(net1043));
 sg13g2_nor2_1 _22479_ (.A(net1028),
    .B(_04886_),
    .Y(_04887_));
 sg13g2_buf_2 _22480_ (.A(_04887_),
    .X(_04888_));
 sg13g2_a21oi_1 _22481_ (.A1(_10050_),
    .A2(net893),
    .Y(_04889_),
    .B1(net1034));
 sg13g2_nor3_1 _22482_ (.A(net1030),
    .B(net784),
    .C(_04889_),
    .Y(_04890_));
 sg13g2_nor2_1 _22483_ (.A(_10889_),
    .B(net780),
    .Y(_04891_));
 sg13g2_o21ai_1 _22484_ (.B1(net767),
    .Y(_04892_),
    .A1(_04890_),
    .A2(_04891_));
 sg13g2_nor3_1 _22485_ (.A(net1030),
    .B(net696),
    .C(_09567_),
    .Y(_04893_));
 sg13g2_o21ai_1 _22486_ (.B1(net1039),
    .Y(_04894_),
    .A1(_09394_),
    .A2(_04893_));
 sg13g2_nand2_1 _22487_ (.Y(_04895_),
    .A(net894),
    .B(net1034));
 sg13g2_o21ai_1 _22488_ (.B1(_04895_),
    .Y(_04896_),
    .A1(net780),
    .A2(net1034));
 sg13g2_nand2_1 _22489_ (.Y(_04897_),
    .A(net783),
    .B(_10050_));
 sg13g2_buf_1 _22490_ (.A(_04897_),
    .X(_04898_));
 sg13g2_nand2_1 _22491_ (.Y(_04899_),
    .A(net893),
    .B(_09567_));
 sg13g2_o21ai_1 _22492_ (.B1(_04895_),
    .Y(_04900_),
    .A1(_04898_),
    .A2(_04899_));
 sg13g2_a22oi_1 _22493_ (.Y(_04901_),
    .B1(_04900_),
    .B2(net1030),
    .A2(_04896_),
    .A1(net783));
 sg13g2_nand3_1 _22494_ (.B(_04894_),
    .C(_04901_),
    .A(_04892_),
    .Y(_04902_));
 sg13g2_buf_2 _22495_ (.A(_04902_),
    .X(_04903_));
 sg13g2_nand3_1 _22496_ (.B(_09220_),
    .C(_04903_),
    .A(_09219_),
    .Y(_04904_));
 sg13g2_nand2_1 _22497_ (.Y(_04905_),
    .A(net893),
    .B(net784));
 sg13g2_buf_2 _22498_ (.A(_04905_),
    .X(_04906_));
 sg13g2_nor3_1 _22499_ (.A(net783),
    .B(net1039),
    .C(_04906_),
    .Y(_04907_));
 sg13g2_buf_1 _22500_ (.A(_04907_),
    .X(_04908_));
 sg13g2_and2_1 _22501_ (.A(net862),
    .B(_04908_),
    .X(_04909_));
 sg13g2_buf_1 _22502_ (.A(_04909_),
    .X(_04910_));
 sg13g2_buf_1 _22503_ (.A(_09567_),
    .X(_04911_));
 sg13g2_nand2_1 _22504_ (.Y(_04912_),
    .A(net893),
    .B(_09341_));
 sg13g2_buf_1 _22505_ (.A(_04912_),
    .X(_04913_));
 sg13g2_nor3_2 _22506_ (.A(net960),
    .B(net648),
    .C(net583),
    .Y(_04914_));
 sg13g2_buf_2 _22507_ (.A(\cpu.gpio.r_src_o[4][0] ),
    .X(_04915_));
 sg13g2_a22oi_1 _22508_ (.Y(_04916_),
    .B1(_04914_),
    .B2(_04915_),
    .A2(_04910_),
    .A1(_09219_));
 sg13g2_nor3_1 _22509_ (.A(net1030),
    .B(net648),
    .C(net583),
    .Y(_04917_));
 sg13g2_buf_2 _22510_ (.A(_04917_),
    .X(_04918_));
 sg13g2_nand2_1 _22511_ (.Y(_04919_),
    .A(net783),
    .B(_09271_));
 sg13g2_buf_1 _22512_ (.A(_04919_),
    .X(_04920_));
 sg13g2_nor3_1 _22513_ (.A(_09567_),
    .B(_04906_),
    .C(_04920_),
    .Y(_04921_));
 sg13g2_buf_1 _22514_ (.A(_04921_),
    .X(_04922_));
 sg13g2_buf_2 _22515_ (.A(\cpu.gpio.r_src_io[6][0] ),
    .X(_04923_));
 sg13g2_a22oi_1 _22516_ (.Y(_04924_),
    .B1(net446),
    .B2(_04923_),
    .A2(_04918_),
    .A1(_09220_));
 sg13g2_buf_2 _22517_ (.A(\cpu.gpio.r_uart_rx_src[0] ),
    .X(_04925_));
 sg13g2_nor3_1 _22518_ (.A(_09998_),
    .B(net1039),
    .C(_02739_),
    .Y(_04926_));
 sg13g2_buf_1 _22519_ (.A(_04926_),
    .X(_04927_));
 sg13g2_buf_1 _22520_ (.A(net541),
    .X(_04928_));
 sg13g2_nand2_1 _22521_ (.Y(_04929_),
    .A(net900),
    .B(net444));
 sg13g2_nor2_1 _22522_ (.A(net1034),
    .B(_04929_),
    .Y(_04930_));
 sg13g2_buf_1 _22523_ (.A(_04930_),
    .X(_04931_));
 sg13g2_buf_2 _22524_ (.A(\cpu.gpio.r_spi_miso_src[0][0] ),
    .X(_04932_));
 sg13g2_buf_2 _22525_ (.A(\cpu.gpio.r_src_o[6][0] ),
    .X(_04933_));
 sg13g2_nor3_2 _22526_ (.A(net862),
    .B(net648),
    .C(_04920_),
    .Y(_04934_));
 sg13g2_nor3_1 _22527_ (.A(_09567_),
    .B(net583),
    .C(_04906_),
    .Y(_04935_));
 sg13g2_buf_1 _22528_ (.A(_04935_),
    .X(_04936_));
 sg13g2_buf_2 _22529_ (.A(\cpu.gpio.r_src_io[4][0] ),
    .X(_04937_));
 sg13g2_a22oi_1 _22530_ (.Y(_04938_),
    .B1(net443),
    .B2(_04937_),
    .A2(_04934_),
    .A1(_04933_));
 sg13g2_inv_1 _22531_ (.Y(_04939_),
    .A(_04938_));
 sg13g2_a221oi_1 _22532_ (.B2(_04932_),
    .C1(_04939_),
    .B1(_04931_),
    .A1(_04925_),
    .Y(_04940_),
    .A2(net445));
 sg13g2_nand4_1 _22533_ (.B(_04916_),
    .C(_04924_),
    .A(_04904_),
    .Y(_04941_),
    .D(_04940_));
 sg13g2_nand2_1 _22534_ (.Y(_04942_),
    .A(net784),
    .B(_04895_));
 sg13g2_buf_2 _22535_ (.A(_00226_),
    .X(_04943_));
 sg13g2_or2_1 _22536_ (.X(_04944_),
    .B(_04943_),
    .A(net784));
 sg13g2_o21ai_1 _22537_ (.B1(_04944_),
    .Y(_04945_),
    .A1(net783),
    .A2(_04899_));
 sg13g2_nor2_1 _22538_ (.A(_09521_),
    .B(_09416_),
    .Y(_04946_));
 sg13g2_nor2_1 _22539_ (.A(net1039),
    .B(_04946_),
    .Y(_04947_));
 sg13g2_a221oi_1 _22540_ (.B2(net1039),
    .C1(_04947_),
    .B1(_04945_),
    .A1(net767),
    .Y(_04948_),
    .A2(_04942_));
 sg13g2_nand2_1 _22541_ (.Y(_04949_),
    .A(net767),
    .B(net1039));
 sg13g2_buf_2 _22542_ (.A(_04949_),
    .X(_04950_));
 sg13g2_nor3_1 _22543_ (.A(net1030),
    .B(_04950_),
    .C(_04906_),
    .Y(_04951_));
 sg13g2_buf_2 _22544_ (.A(_04951_),
    .X(_04952_));
 sg13g2_nor3_1 _22545_ (.A(_04948_),
    .B(net445),
    .C(_04952_),
    .Y(_04953_));
 sg13g2_buf_2 _22546_ (.A(_04953_),
    .X(_04954_));
 sg13g2_inv_1 _22547_ (.Y(_04955_),
    .A(_00312_));
 sg13g2_nor2_1 _22548_ (.A(_04950_),
    .B(_04906_),
    .Y(_04956_));
 sg13g2_buf_1 _22549_ (.A(_04956_),
    .X(_04957_));
 sg13g2_a221oi_1 _22550_ (.B2(_11982_),
    .C1(net858),
    .B1(net447),
    .A1(_04955_),
    .Y(_04958_),
    .A2(_04957_));
 sg13g2_a21oi_1 _22551_ (.A1(\cpu.spi.r_mode[2][0] ),
    .A2(net447),
    .Y(_04959_),
    .B1(net862));
 sg13g2_a22oi_1 _22552_ (.Y(_04960_),
    .B1(\cpu.spi.r_timeout[0] ),
    .B2(net632),
    .A2(_04943_),
    .A1(_09252_));
 sg13g2_nand3_1 _22553_ (.B(net780),
    .C(\cpu.spi.r_ready ),
    .A(net889),
    .Y(_04961_));
 sg13g2_o21ai_1 _22554_ (.B1(_04961_),
    .Y(_04962_),
    .A1(net763),
    .A2(_04960_));
 sg13g2_nor3_1 _22555_ (.A(_09567_),
    .B(_04950_),
    .C(_04906_),
    .Y(_04963_));
 sg13g2_buf_2 _22556_ (.A(_04963_),
    .X(_04964_));
 sg13g2_buf_1 _22557_ (.A(\cpu.spi.r_clk_count[2][0] ),
    .X(_04965_));
 sg13g2_nand3_1 _22558_ (.B(_09567_),
    .C(net623),
    .A(_09272_),
    .Y(_04966_));
 sg13g2_buf_2 _22559_ (.A(_04966_),
    .X(_04967_));
 sg13g2_nor2_1 _22560_ (.A(_00311_),
    .B(_04967_),
    .Y(_04968_));
 sg13g2_a221oi_1 _22561_ (.B2(_04965_),
    .C1(_04968_),
    .B1(_04964_),
    .A1(net695),
    .Y(_04969_),
    .A2(_04962_));
 sg13g2_o21ai_1 _22562_ (.B1(_04969_),
    .Y(_04970_),
    .A1(_04958_),
    .A2(_04959_));
 sg13g2_a221oi_1 _22563_ (.B2(_09320_),
    .C1(_04970_),
    .B1(_04954_),
    .A1(\cpu.spi.r_mode[1][0] ),
    .Y(_04971_),
    .A2(net445));
 sg13g2_buf_1 _22564_ (.A(\cpu.intr.r_clock_count[16] ),
    .X(_04972_));
 sg13g2_nand2_1 _22565_ (.Y(_04973_),
    .A(net782),
    .B(_09965_));
 sg13g2_o21ai_1 _22566_ (.B1(_04973_),
    .Y(_04974_),
    .A1(net782),
    .A2(_00283_));
 sg13g2_buf_1 _22567_ (.A(_09419_),
    .X(_04975_));
 sg13g2_buf_1 _22568_ (.A(net507),
    .X(_04976_));
 sg13g2_buf_1 _22569_ (.A(net442),
    .X(_04977_));
 sg13g2_buf_1 _22570_ (.A(net399),
    .X(_04978_));
 sg13g2_and2_1 _22571_ (.A(net900),
    .B(\cpu.intr.r_clock_cmp[16] ),
    .X(_04979_));
 sg13g2_a21oi_1 _22572_ (.A1(net889),
    .A2(\cpu.intr.r_clock_cmp[0] ),
    .Y(_04980_),
    .B1(_04979_));
 sg13g2_nor2_1 _22573_ (.A(net648),
    .B(_04950_),
    .Y(_04981_));
 sg13g2_buf_1 _22574_ (.A(_04981_),
    .X(_04982_));
 sg13g2_o21ai_1 _22575_ (.B1(_04982_),
    .Y(_04983_),
    .A1(_09248_),
    .A2(_09249_));
 sg13g2_o21ai_1 _22576_ (.B1(_04983_),
    .Y(_04984_),
    .A1(net653),
    .A2(_04980_));
 sg13g2_a221oi_1 _22577_ (.B2(net361),
    .C1(_04984_),
    .B1(_04974_),
    .A1(_04972_),
    .Y(_04985_),
    .A2(net412));
 sg13g2_nand3_1 _22578_ (.B(\cpu.intr.r_timer_reload[16] ),
    .C(net374),
    .A(net674),
    .Y(_04986_));
 sg13g2_buf_1 _22579_ (.A(net621),
    .X(_04987_));
 sg13g2_buf_1 _22580_ (.A(net506),
    .X(_04988_));
 sg13g2_buf_1 _22581_ (.A(_04988_),
    .X(_04989_));
 sg13g2_a22oi_1 _22582_ (.Y(_04990_),
    .B1(net398),
    .B2(_10128_),
    .A2(net374),
    .A1(\cpu.intr.r_timer_reload[0] ));
 sg13g2_or2_1 _22583_ (.X(_04991_),
    .B(_04990_),
    .A(net674));
 sg13g2_nor2_1 _22584_ (.A(net648),
    .B(_04898_),
    .Y(_04992_));
 sg13g2_buf_1 _22585_ (.A(_04992_),
    .X(_04993_));
 sg13g2_buf_1 _22586_ (.A(_04993_),
    .X(_04994_));
 sg13g2_a21oi_1 _22587_ (.A1(_04950_),
    .A2(net583),
    .Y(_04995_),
    .B1(net696));
 sg13g2_nor2_1 _22588_ (.A(net894),
    .B(_04995_),
    .Y(_04996_));
 sg13g2_buf_1 _22589_ (.A(_04996_),
    .X(_04997_));
 sg13g2_o21ai_1 _22590_ (.B1(net396),
    .Y(_04998_),
    .A1(_09248_),
    .A2(_09249_));
 sg13g2_inv_1 _22591_ (.Y(_04999_),
    .A(_04998_));
 sg13g2_o21ai_1 _22592_ (.B1(\cpu.intr.r_enable[0] ),
    .Y(_05000_),
    .A1(net397),
    .A2(_04999_));
 sg13g2_nand4_1 _22593_ (.B(_04986_),
    .C(_04991_),
    .A(_04985_),
    .Y(_05001_),
    .D(_05000_));
 sg13g2_nand2_1 _22594_ (.Y(_05002_),
    .A(_04886_),
    .B(_10001_));
 sg13g2_buf_1 _22595_ (.A(_05002_),
    .X(_05003_));
 sg13g2_o21ai_1 _22596_ (.B1(net733),
    .Y(_05004_),
    .A1(_09421_),
    .A2(_09732_));
 sg13g2_buf_2 _22597_ (.A(_05004_),
    .X(_05005_));
 sg13g2_a22oi_1 _22598_ (.Y(_05006_),
    .B1(net447),
    .B2(\cpu.uart.r_div_value[0] ),
    .A2(_04957_),
    .A1(\cpu.uart.r_div_value[8] ));
 sg13g2_nor2_1 _22599_ (.A(net648),
    .B(_04920_),
    .Y(_05007_));
 sg13g2_buf_1 _22600_ (.A(_05007_),
    .X(_05008_));
 sg13g2_a22oi_1 _22601_ (.Y(_05009_),
    .B1(net440),
    .B2(\cpu.uart.r_x_invert ),
    .A2(_04993_),
    .A1(_09248_));
 sg13g2_nand2_1 _22602_ (.Y(_05010_),
    .A(_05006_),
    .B(_05009_));
 sg13g2_a21oi_1 _22603_ (.A1(\cpu.uart.r_in[0] ),
    .A2(_05005_),
    .Y(_05011_),
    .B1(_05010_));
 sg13g2_o21ai_1 _22604_ (.B1(net1041),
    .Y(_05012_),
    .A1(net582),
    .A2(_05011_));
 sg13g2_a21oi_1 _22605_ (.A1(_10059_),
    .A2(_05001_),
    .Y(_05013_),
    .B1(_05012_));
 sg13g2_o21ai_1 _22606_ (.B1(_05013_),
    .Y(_05014_),
    .A1(_09208_),
    .A2(_04971_));
 sg13g2_a21oi_1 _22607_ (.A1(_04888_),
    .A2(_04941_),
    .Y(_05015_),
    .B1(_05014_));
 sg13g2_buf_1 _22608_ (.A(net626),
    .X(_05016_));
 sg13g2_buf_1 _22609_ (.A(net505),
    .X(_05017_));
 sg13g2_a22oi_1 _22610_ (.Y(_05018_),
    .B1(net624),
    .B2(\cpu.dcache.r_data[3][0] ),
    .A2(net625),
    .A1(\cpu.dcache.r_data[2][0] ));
 sg13g2_a22oi_1 _22611_ (.Y(_05019_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[4][0] ),
    .A2(net541),
    .A1(\cpu.dcache.r_data[5][0] ));
 sg13g2_nand2_1 _22612_ (.Y(_05020_),
    .A(_05018_),
    .B(_05019_));
 sg13g2_a221oi_1 _22613_ (.B2(\cpu.dcache.r_data[6][0] ),
    .C1(_05020_),
    .B1(net507),
    .A1(\cpu.dcache.r_data[7][0] ),
    .Y(_05021_),
    .A2(net540));
 sg13g2_nor2_1 _22614_ (.A(\cpu.dcache.r_data[0][0] ),
    .B(_04913_),
    .Y(_05022_));
 sg13g2_a21oi_1 _22615_ (.A1(_04913_),
    .A2(_05021_),
    .Y(_05023_),
    .B1(_05022_));
 sg13g2_nand3b_1 _22616_ (.B(net439),
    .C(_05021_),
    .Y(_05024_),
    .A_N(\cpu.dcache.r_data[1][0] ));
 sg13g2_o21ai_1 _22617_ (.B1(_05024_),
    .Y(_05025_),
    .A1(net439),
    .A2(_05023_));
 sg13g2_buf_1 _22618_ (.A(net624),
    .X(_05026_));
 sg13g2_buf_1 _22619_ (.A(net504),
    .X(_05027_));
 sg13g2_buf_1 _22620_ (.A(net444),
    .X(_05028_));
 sg13g2_a22oi_1 _22621_ (.Y(_05029_),
    .B1(net395),
    .B2(\cpu.dcache.r_data[5][16] ),
    .A2(net438),
    .A1(\cpu.dcache.r_data[3][16] ));
 sg13g2_buf_1 _22622_ (.A(net625),
    .X(_05030_));
 sg13g2_buf_1 _22623_ (.A(net503),
    .X(_05031_));
 sg13g2_a22oi_1 _22624_ (.Y(_05032_),
    .B1(net437),
    .B2(\cpu.dcache.r_data[2][16] ),
    .A2(net505),
    .A1(\cpu.dcache.r_data[1][16] ));
 sg13g2_mux2_1 _22625_ (.A0(\cpu.dcache.r_data[4][16] ),
    .A1(\cpu.dcache.r_data[6][16] ),
    .S(net696),
    .X(_05033_));
 sg13g2_a22oi_1 _22626_ (.Y(_05034_),
    .B1(_05033_),
    .B2(net767),
    .A2(_09521_),
    .A1(\cpu.dcache.r_data[7][16] ));
 sg13g2_nand2b_1 _22627_ (.Y(_05035_),
    .B(net894),
    .A_N(_05034_));
 sg13g2_nand3_1 _22628_ (.B(_05032_),
    .C(_05035_),
    .A(_05029_),
    .Y(_05036_));
 sg13g2_mux2_1 _22629_ (.A0(\cpu.dcache.r_data[0][16] ),
    .A1(_05036_),
    .S(_09517_),
    .X(_05037_));
 sg13g2_a21oi_2 _22630_ (.B1(_08580_),
    .Y(_05038_),
    .A2(net1125),
    .A1(net1126));
 sg13g2_nor3_2 _22631_ (.A(_08576_),
    .B(_09209_),
    .C(_08584_),
    .Y(_05039_));
 sg13g2_nand2_1 _22632_ (.Y(_05040_),
    .A(_05038_),
    .B(_05039_));
 sg13g2_buf_2 _22633_ (.A(_05040_),
    .X(_05041_));
 sg13g2_a21oi_1 _22634_ (.A1(net615),
    .A2(_05037_),
    .Y(_05042_),
    .B1(_05041_));
 sg13g2_o21ai_1 _22635_ (.B1(_05042_),
    .Y(_05043_),
    .A1(net537),
    .A2(_05025_));
 sg13g2_buf_1 _22636_ (.A(net619),
    .X(_05044_));
 sg13g2_buf_1 _22637_ (.A(_05044_),
    .X(_05045_));
 sg13g2_a22oi_1 _22638_ (.Y(_05046_),
    .B1(_05028_),
    .B2(\cpu.dcache.r_data[5][24] ),
    .A2(net505),
    .A1(\cpu.dcache.r_data[1][24] ));
 sg13g2_a22oi_1 _22639_ (.Y(_05047_),
    .B1(net438),
    .B2(\cpu.dcache.r_data[3][24] ),
    .A2(net437),
    .A1(\cpu.dcache.r_data[2][24] ));
 sg13g2_mux2_1 _22640_ (.A0(\cpu.dcache.r_data[4][24] ),
    .A1(\cpu.dcache.r_data[6][24] ),
    .S(net696),
    .X(_05048_));
 sg13g2_a22oi_1 _22641_ (.Y(_05049_),
    .B1(_05048_),
    .B2(net767),
    .A2(_09521_),
    .A1(\cpu.dcache.r_data[7][24] ));
 sg13g2_nand2b_1 _22642_ (.Y(_05050_),
    .B(_09555_),
    .A_N(_05049_));
 sg13g2_and4_1 _22643_ (.A(_09517_),
    .B(_05046_),
    .C(_05047_),
    .D(_05050_),
    .X(_05051_));
 sg13g2_a21oi_1 _22644_ (.A1(_00309_),
    .A2(_05045_),
    .Y(_05052_),
    .B1(_05051_));
 sg13g2_a22oi_1 _22645_ (.Y(_05053_),
    .B1(_05027_),
    .B2(\cpu.dcache.r_data[3][8] ),
    .A2(net437),
    .A1(\cpu.dcache.r_data[2][8] ));
 sg13g2_a22oi_1 _22646_ (.Y(_05054_),
    .B1(net395),
    .B2(\cpu.dcache.r_data[5][8] ),
    .A2(net505),
    .A1(\cpu.dcache.r_data[1][8] ));
 sg13g2_inv_1 _22647_ (.Y(_05055_),
    .A(_00310_));
 sg13g2_a22oi_1 _22648_ (.Y(_05056_),
    .B1(net502),
    .B2(_05055_),
    .A2(net472),
    .A1(\cpu.dcache.r_data[7][8] ));
 sg13g2_a22oi_1 _22649_ (.Y(_05057_),
    .B1(net441),
    .B2(\cpu.dcache.r_data[4][8] ),
    .A2(net442),
    .A1(\cpu.dcache.r_data[6][8] ));
 sg13g2_nand4_1 _22650_ (.B(_05054_),
    .C(_05056_),
    .A(_05053_),
    .Y(_05058_),
    .D(_05057_));
 sg13g2_and2_1 _22651_ (.A(_10052_),
    .B(_05058_),
    .X(_05059_));
 sg13g2_a21oi_1 _22652_ (.A1(net997),
    .A2(_05052_),
    .Y(_05060_),
    .B1(_05059_));
 sg13g2_a21oi_1 _22653_ (.A1(_09992_),
    .A2(_05037_),
    .Y(_05061_),
    .B1(_12016_));
 sg13g2_nand3b_1 _22654_ (.B(net1060),
    .C(_08610_),
    .Y(_05062_),
    .A_N(_08584_));
 sg13g2_buf_2 _22655_ (.A(_05062_),
    .X(_05063_));
 sg13g2_mux2_1 _22656_ (.A0(_05060_),
    .A1(_05061_),
    .S(_05063_),
    .X(_05064_));
 sg13g2_buf_1 _22657_ (.A(_05039_),
    .X(_05065_));
 sg13g2_nor2_1 _22658_ (.A(net997),
    .B(net717),
    .Y(_05066_));
 sg13g2_a22oi_1 _22659_ (.Y(_05067_),
    .B1(_05025_),
    .B2(_05066_),
    .A2(_05064_),
    .A1(_05041_));
 sg13g2_a21oi_1 _22660_ (.A1(_05043_),
    .A2(_05067_),
    .Y(_05068_),
    .B1(net848));
 sg13g2_nor3_1 _22661_ (.A(_04884_),
    .B(_05015_),
    .C(_05068_),
    .Y(_05069_));
 sg13g2_a21oi_1 _22662_ (.A1(net833),
    .A2(net78),
    .Y(_05070_),
    .B1(_05069_));
 sg13g2_o21ai_1 _22663_ (.B1(net721),
    .Y(_05071_),
    .A1(net584),
    .A2(net197));
 sg13g2_mux2_1 _22664_ (.A0(_05070_),
    .A1(_05071_),
    .S(net191),
    .X(_05072_));
 sg13g2_o21ai_1 _22665_ (.B1(_05072_),
    .Y(_01029_),
    .A1(_04857_),
    .A2(_04882_));
 sg13g2_nand2_1 _22666_ (.Y(_05073_),
    .A(net191),
    .B(net226));
 sg13g2_nor2_2 _22667_ (.A(net508),
    .B(_05073_),
    .Y(_05074_));
 sg13g2_nand3b_1 _22668_ (.B(net226),
    .C(_04858_),
    .Y(_05075_),
    .A_N(_04803_));
 sg13g2_o21ai_1 _22669_ (.B1(_05075_),
    .Y(_05076_),
    .A1(net961),
    .A2(net226));
 sg13g2_inv_1 _22670_ (.Y(_05077_),
    .A(_09208_));
 sg13g2_inv_1 _22671_ (.Y(_05078_),
    .A(_00157_));
 sg13g2_buf_1 _22672_ (.A(\cpu.spi.r_clk_count[2][7] ),
    .X(_05079_));
 sg13g2_a22oi_1 _22673_ (.Y(_05080_),
    .B1(_04964_),
    .B2(_05079_),
    .A2(_04952_),
    .A1(_05078_));
 sg13g2_nor2_1 _22674_ (.A(net780),
    .B(_04920_),
    .Y(_05081_));
 sg13g2_buf_2 _22675_ (.A(_05081_),
    .X(_05082_));
 sg13g2_nor2_1 _22676_ (.A(_00156_),
    .B(_04967_),
    .Y(_05083_));
 sg13g2_a21oi_1 _22677_ (.A1(\cpu.spi.r_timeout[7] ),
    .A2(_05082_),
    .Y(_05084_),
    .B1(_05083_));
 sg13g2_nand2b_1 _22678_ (.Y(_05085_),
    .B(_04954_),
    .A_N(_00220_));
 sg13g2_nand3_1 _22679_ (.B(_05084_),
    .C(_05085_),
    .A(_05080_),
    .Y(_05086_));
 sg13g2_and3_1 _22680_ (.X(_05087_),
    .A(_09227_),
    .B(net960),
    .C(_04982_));
 sg13g2_o21ai_1 _22681_ (.B1(\cpu.gpio.r_enable_io[7] ),
    .Y(_05088_),
    .A1(_04952_),
    .A2(_05087_));
 sg13g2_nand2_1 _22682_ (.Y(_05089_),
    .A(net895),
    .B(_10120_));
 sg13g2_nand2b_1 _22683_ (.Y(_05090_),
    .B(_05007_),
    .A_N(_00159_));
 sg13g2_o21ai_1 _22684_ (.B1(_05090_),
    .Y(_05091_),
    .A1(_00161_),
    .A2(_05089_));
 sg13g2_nor2b_1 _22685_ (.A(_00158_),
    .B_N(net446),
    .Y(_05092_));
 sg13g2_a221oi_1 _22686_ (.B2(_09999_),
    .C1(_05092_),
    .B1(_05091_),
    .A1(_09217_),
    .Y(_05093_),
    .A2(_04918_));
 sg13g2_buf_1 _22687_ (.A(\cpu.gpio.r_src_io[5][3] ),
    .X(_05094_));
 sg13g2_nand2_2 _22688_ (.Y(_05095_),
    .A(net1034),
    .B(_04993_));
 sg13g2_nor2_1 _22689_ (.A(_00160_),
    .B(_05095_),
    .Y(_05096_));
 sg13g2_a221oi_1 _22690_ (.B2(_05094_),
    .C1(_05096_),
    .B1(net443),
    .A1(\cpu.gpio.r_enable_in[7] ),
    .Y(_05097_),
    .A2(net362));
 sg13g2_nand2_1 _22691_ (.Y(_05098_),
    .A(_05093_),
    .B(_05097_));
 sg13g2_nor2_1 _22692_ (.A(net1039),
    .B(_10110_),
    .Y(_05099_));
 sg13g2_buf_1 _22693_ (.A(_05099_),
    .X(_05100_));
 sg13g2_a22oi_1 _22694_ (.Y(_05101_),
    .B1(net501),
    .B2(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .A2(_10122_),
    .A1(\cpu.gpio.genblk2[7].srcs_io[0] ));
 sg13g2_nand2_1 _22695_ (.Y(_05102_),
    .A(net889),
    .B(net10));
 sg13g2_o21ai_1 _22696_ (.B1(_05102_),
    .Y(_05103_),
    .A1(net889),
    .A2(_00162_));
 sg13g2_a22oi_1 _22697_ (.Y(_05104_),
    .B1(_05103_),
    .B2(net444),
    .A2(_05007_),
    .A1(_09227_));
 sg13g2_a21oi_1 _22698_ (.A1(_05101_),
    .A2(_05104_),
    .Y(_05105_),
    .B1(net1034));
 sg13g2_nor2_1 _22699_ (.A(_05098_),
    .B(_05105_),
    .Y(_05106_));
 sg13g2_nand2b_1 _22700_ (.Y(_05107_),
    .B(_04903_),
    .A_N(_09218_));
 sg13g2_nand3_1 _22701_ (.B(_05106_),
    .C(_05107_),
    .A(_05088_),
    .Y(_05108_));
 sg13g2_a22oi_1 _22702_ (.Y(_05109_),
    .B1(_05005_),
    .B2(\cpu.uart.r_in[7] ),
    .A2(net447),
    .A1(\cpu.uart.r_div_value[7] ));
 sg13g2_nor2_1 _22703_ (.A(_10001_),
    .B(net396),
    .Y(_05110_));
 sg13g2_buf_2 _22704_ (.A(\cpu.intr.r_clock_count[23] ),
    .X(_05111_));
 sg13g2_mux2_1 _22705_ (.A0(_09967_),
    .A1(_09987_),
    .S(net900),
    .X(_05112_));
 sg13g2_a22oi_1 _22706_ (.Y(_05113_),
    .B1(_05112_),
    .B2(net442),
    .A2(_10122_),
    .A1(_05111_));
 sg13g2_mux2_1 _22707_ (.A0(\cpu.intr.r_clock_cmp[7] ),
    .A1(\cpu.intr.r_clock_cmp[23] ),
    .S(net1039),
    .X(_05114_));
 sg13g2_mux2_1 _22708_ (.A0(\cpu.intr.r_timer_reload[7] ),
    .A1(\cpu.intr.r_timer_reload[23] ),
    .S(net900),
    .X(_05115_));
 sg13g2_a22oi_1 _22709_ (.Y(_05116_),
    .B1(_05115_),
    .B2(net472),
    .A2(_05114_),
    .A1(net444));
 sg13g2_nand2_1 _22710_ (.Y(_05117_),
    .A(_10171_),
    .B(net501));
 sg13g2_nand3_1 _22711_ (.B(_05116_),
    .C(_05117_),
    .A(_05113_),
    .Y(_05118_));
 sg13g2_nand2_1 _22712_ (.Y(_05119_),
    .A(_05110_),
    .B(_05118_));
 sg13g2_o21ai_1 _22713_ (.B1(_05119_),
    .Y(_05120_),
    .A1(net582),
    .A2(_05109_));
 sg13g2_a221oi_1 _22714_ (.B2(_04888_),
    .C1(_05120_),
    .B1(_05108_),
    .A1(_05077_),
    .Y(_05121_),
    .A2(_05086_));
 sg13g2_nor2_1 _22715_ (.A(_08581_),
    .B(_05063_),
    .Y(_05122_));
 sg13g2_buf_1 _22716_ (.A(_05122_),
    .X(_05123_));
 sg13g2_a22oi_1 _22717_ (.Y(_05124_),
    .B1(net623),
    .B2(\cpu.dcache.r_data[6][7] ),
    .A2(net626),
    .A1(\cpu.dcache.r_data[1][7] ));
 sg13g2_a22oi_1 _22718_ (.Y(_05125_),
    .B1(net504),
    .B2(\cpu.dcache.r_data[3][7] ),
    .A2(net625),
    .A1(\cpu.dcache.r_data[2][7] ));
 sg13g2_a22oi_1 _22719_ (.Y(_05126_),
    .B1(net541),
    .B2(\cpu.dcache.r_data[5][7] ),
    .A2(net540),
    .A1(\cpu.dcache.r_data[7][7] ));
 sg13g2_inv_1 _22720_ (.Y(_05127_),
    .A(_00152_));
 sg13g2_a22oi_1 _22721_ (.Y(_05128_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[4][7] ),
    .A2(net619),
    .A1(_05127_));
 sg13g2_nand4_1 _22722_ (.B(_05125_),
    .C(_05126_),
    .A(_05124_),
    .Y(_05129_),
    .D(_05128_));
 sg13g2_buf_1 _22723_ (.A(_05129_),
    .X(_05130_));
 sg13g2_a22oi_1 _22724_ (.Y(_05131_),
    .B1(net626),
    .B2(\cpu.dcache.r_data[1][23] ),
    .A2(net540),
    .A1(\cpu.dcache.r_data[7][23] ));
 sg13g2_a22oi_1 _22725_ (.Y(_05132_),
    .B1(net623),
    .B2(\cpu.dcache.r_data[6][23] ),
    .A2(net503),
    .A1(\cpu.dcache.r_data[2][23] ));
 sg13g2_inv_1 _22726_ (.Y(_05133_),
    .A(_00153_));
 sg13g2_a22oi_1 _22727_ (.Y(_05134_),
    .B1(net619),
    .B2(_05133_),
    .A2(net541),
    .A1(\cpu.dcache.r_data[5][23] ));
 sg13g2_a22oi_1 _22728_ (.Y(_05135_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[4][23] ),
    .A2(net504),
    .A1(\cpu.dcache.r_data[3][23] ));
 sg13g2_nand4_1 _22729_ (.B(_05132_),
    .C(_05134_),
    .A(_05131_),
    .Y(_05136_),
    .D(_05135_));
 sg13g2_buf_1 _22730_ (.A(_05136_),
    .X(_05137_));
 sg13g2_nor2_1 _22731_ (.A(_10051_),
    .B(_12016_),
    .Y(_05138_));
 sg13g2_a221oi_1 _22732_ (.B2(_05138_),
    .C1(_05039_),
    .B1(_05137_),
    .A1(_12016_),
    .Y(_05139_),
    .A2(_05130_));
 sg13g2_a22oi_1 _22733_ (.Y(_05140_),
    .B1(net507),
    .B2(\cpu.dcache.r_data[6][15] ),
    .A2(net626),
    .A1(\cpu.dcache.r_data[1][15] ));
 sg13g2_a22oi_1 _22734_ (.Y(_05141_),
    .B1(net504),
    .B2(\cpu.dcache.r_data[3][15] ),
    .A2(net503),
    .A1(\cpu.dcache.r_data[2][15] ));
 sg13g2_a22oi_1 _22735_ (.Y(_05142_),
    .B1(net541),
    .B2(\cpu.dcache.r_data[5][15] ),
    .A2(net540),
    .A1(\cpu.dcache.r_data[7][15] ));
 sg13g2_inv_1 _22736_ (.Y(_05143_),
    .A(_00155_));
 sg13g2_a22oi_1 _22737_ (.Y(_05144_),
    .B1(_04987_),
    .B2(\cpu.dcache.r_data[4][15] ),
    .A2(net619),
    .A1(_05143_));
 sg13g2_nand4_1 _22738_ (.B(_05141_),
    .C(_05142_),
    .A(_05140_),
    .Y(_05145_),
    .D(_05144_));
 sg13g2_a22oi_1 _22739_ (.Y(_05146_),
    .B1(_04975_),
    .B2(\cpu.dcache.r_data[6][31] ),
    .A2(net626),
    .A1(\cpu.dcache.r_data[1][31] ));
 sg13g2_a22oi_1 _22740_ (.Y(_05147_),
    .B1(net541),
    .B2(\cpu.dcache.r_data[5][31] ),
    .A2(_05030_),
    .A1(\cpu.dcache.r_data[2][31] ));
 sg13g2_inv_1 _22741_ (.Y(_05148_),
    .A(_00154_));
 sg13g2_a22oi_1 _22742_ (.Y(_05149_),
    .B1(_04987_),
    .B2(\cpu.dcache.r_data[4][31] ),
    .A2(_09641_),
    .A1(_05148_));
 sg13g2_a22oi_1 _22743_ (.Y(_05150_),
    .B1(net504),
    .B2(\cpu.dcache.r_data[3][31] ),
    .A2(net540),
    .A1(\cpu.dcache.r_data[7][31] ));
 sg13g2_nand4_1 _22744_ (.B(_05147_),
    .C(_05149_),
    .A(_05146_),
    .Y(_05151_),
    .D(_05150_));
 sg13g2_a221oi_1 _22745_ (.B2(net997),
    .C1(_05063_),
    .B1(_05151_),
    .A1(net889),
    .Y(_05152_),
    .A2(_05145_));
 sg13g2_nor3_1 _22746_ (.A(_05123_),
    .B(_05139_),
    .C(_05152_),
    .Y(_05153_));
 sg13g2_nand2_1 _22747_ (.Y(_05154_),
    .A(_09273_),
    .B(_05137_));
 sg13g2_nand2_1 _22748_ (.Y(_05155_),
    .A(_10051_),
    .B(_05130_));
 sg13g2_a21oi_1 _22749_ (.A1(_05154_),
    .A2(_05155_),
    .Y(_05156_),
    .B1(_05041_));
 sg13g2_nor3_1 _22750_ (.A(net1041),
    .B(_05153_),
    .C(_05156_),
    .Y(_05157_));
 sg13g2_a21oi_2 _22751_ (.B1(_05157_),
    .Y(_05158_),
    .A2(_05121_),
    .A1(net1041));
 sg13g2_nor2_1 _22752_ (.A(_11527_),
    .B(_05158_),
    .Y(_05159_));
 sg13g2_buf_1 _22753_ (.A(_05123_),
    .X(_05160_));
 sg13g2_a22oi_1 _22754_ (.Y(_05161_),
    .B1(net507),
    .B2(\cpu.dcache.r_data[6][10] ),
    .A2(net503),
    .A1(\cpu.dcache.r_data[2][10] ));
 sg13g2_a22oi_1 _22755_ (.Y(_05162_),
    .B1(net504),
    .B2(\cpu.dcache.r_data[3][10] ),
    .A2(net472),
    .A1(\cpu.dcache.r_data[7][10] ));
 sg13g2_inv_1 _22756_ (.Y(_05163_),
    .A(_00103_));
 sg13g2_a22oi_1 _22757_ (.Y(_05164_),
    .B1(net619),
    .B2(_05163_),
    .A2(net444),
    .A1(\cpu.dcache.r_data[5][10] ));
 sg13g2_a22oi_1 _22758_ (.Y(_05165_),
    .B1(net506),
    .B2(\cpu.dcache.r_data[4][10] ),
    .A2(net505),
    .A1(\cpu.dcache.r_data[1][10] ));
 sg13g2_nand4_1 _22759_ (.B(_05162_),
    .C(_05164_),
    .A(_05161_),
    .Y(_05166_),
    .D(_05165_));
 sg13g2_a22oi_1 _22760_ (.Y(_05167_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[4][26] ),
    .A2(net624),
    .A1(\cpu.dcache.r_data[3][26] ));
 sg13g2_a22oi_1 _22761_ (.Y(_05168_),
    .B1(_09533_),
    .B2(\cpu.dcache.r_data[5][26] ),
    .A2(net623),
    .A1(\cpu.dcache.r_data[6][26] ));
 sg13g2_nand2_1 _22762_ (.Y(_05169_),
    .A(_05167_),
    .B(_05168_));
 sg13g2_a221oi_1 _22763_ (.B2(\cpu.dcache.r_data[2][26] ),
    .C1(_05169_),
    .B1(net503),
    .A1(\cpu.dcache.r_data[7][26] ),
    .Y(_05170_),
    .A2(_09757_));
 sg13g2_mux2_1 _22764_ (.A0(_00102_),
    .A1(_05170_),
    .S(net648),
    .X(_05171_));
 sg13g2_nor2_1 _22765_ (.A(\cpu.dcache.r_data[1][26] ),
    .B(_12211_),
    .Y(_05172_));
 sg13g2_a22oi_1 _22766_ (.Y(_05173_),
    .B1(_05172_),
    .B2(_05170_),
    .A2(_05171_),
    .A1(_12211_));
 sg13g2_mux2_1 _22767_ (.A0(_05166_),
    .A1(_05173_),
    .S(net615),
    .X(_05174_));
 sg13g2_nor3_1 _22768_ (.A(net1058),
    .B(_10001_),
    .C(_04997_),
    .Y(_05175_));
 sg13g2_buf_2 _22769_ (.A(_05175_),
    .X(_05176_));
 sg13g2_buf_1 _22770_ (.A(\cpu.intr.r_clock_count[26] ),
    .X(_05177_));
 sg13g2_buf_1 _22771_ (.A(net501),
    .X(_05178_));
 sg13g2_a22oi_1 _22772_ (.Y(_05179_),
    .B1(net435),
    .B2(_10188_),
    .A2(net373),
    .A1(_05177_));
 sg13g2_buf_1 _22773_ (.A(_05028_),
    .X(_05180_));
 sg13g2_buf_1 _22774_ (.A(net360),
    .X(_05181_));
 sg13g2_a22oi_1 _22775_ (.Y(_05182_),
    .B1(net329),
    .B2(\cpu.intr.r_clock_cmp[10] ),
    .A2(net335),
    .A1(\cpu.intr.r_timer_reload[10] ));
 sg13g2_or2_1 _22776_ (.X(_05183_),
    .B(_05182_),
    .A(net617));
 sg13g2_nor2_1 _22777_ (.A(net900),
    .B(_02739_),
    .Y(_05184_));
 sg13g2_buf_2 _22778_ (.A(_05184_),
    .X(_05185_));
 sg13g2_nor2_1 _22779_ (.A(net889),
    .B(net653),
    .Y(_05186_));
 sg13g2_buf_2 _22780_ (.A(_05186_),
    .X(_05187_));
 sg13g2_a22oi_1 _22781_ (.Y(_05188_),
    .B1(_05187_),
    .B2(\cpu.intr.r_clock_cmp[26] ),
    .A2(_05185_),
    .A1(_09966_));
 sg13g2_nand3_1 _22782_ (.B(_05183_),
    .C(_05188_),
    .A(_05179_),
    .Y(_05189_));
 sg13g2_a221oi_1 _22783_ (.B2(_05189_),
    .C1(net1125),
    .B1(_05176_),
    .A1(_05160_),
    .Y(_05190_),
    .A2(_05174_));
 sg13g2_nor3_1 _22784_ (.A(_04884_),
    .B(_05159_),
    .C(_05190_),
    .Y(_05191_));
 sg13g2_a21oi_1 _22785_ (.A1(net1104),
    .A2(net78),
    .Y(_05192_),
    .B1(_05191_));
 sg13g2_mux2_1 _22786_ (.A0(_05076_),
    .A1(_05192_),
    .S(_11540_),
    .X(_05193_));
 sg13g2_a21oi_1 _22787_ (.A1(_04800_),
    .A2(_05074_),
    .Y(_01030_),
    .B1(_05193_));
 sg13g2_a21o_1 _22788_ (.A2(_11526_),
    .A1(_11524_),
    .B1(_11527_),
    .X(_05194_));
 sg13g2_buf_1 _22789_ (.A(_05194_),
    .X(_05195_));
 sg13g2_nor2_1 _22790_ (.A(net581),
    .B(_04344_),
    .Y(_05196_));
 sg13g2_nor2_1 _22791_ (.A(_11540_),
    .B(net197),
    .Y(_05197_));
 sg13g2_nand2_1 _22792_ (.Y(_05198_),
    .A(net191),
    .B(_04251_));
 sg13g2_inv_1 _22793_ (.Y(_05199_),
    .A(net1119));
 sg13g2_mux2_1 _22794_ (.A0(\cpu.dcache.r_data[1][27] ),
    .A1(\cpu.dcache.r_data[3][27] ),
    .S(_09201_),
    .X(_05200_));
 sg13g2_a22oi_1 _22795_ (.Y(_05201_),
    .B1(_05200_),
    .B2(_09286_),
    .A2(_09732_),
    .A1(\cpu.dcache.r_data[2][27] ));
 sg13g2_inv_1 _22796_ (.Y(_05202_),
    .A(_00112_));
 sg13g2_mux2_1 _22797_ (.A0(\cpu.dcache.r_data[5][27] ),
    .A1(\cpu.dcache.r_data[7][27] ),
    .S(net696),
    .X(_05203_));
 sg13g2_a22oi_1 _22798_ (.Y(_05204_),
    .B1(_05203_),
    .B2(_09270_),
    .A2(_09557_),
    .A1(\cpu.dcache.r_data[4][27] ));
 sg13g2_nor2_1 _22799_ (.A(_11931_),
    .B(_05204_),
    .Y(_05205_));
 sg13g2_a221oi_1 _22800_ (.B2(_05202_),
    .C1(_05205_),
    .B1(_05045_),
    .A1(\cpu.dcache.r_data[6][27] ),
    .Y(_05206_),
    .A2(net399));
 sg13g2_o21ai_1 _22801_ (.B1(_05206_),
    .Y(_05207_),
    .A1(_05199_),
    .A2(_05201_));
 sg13g2_a22oi_1 _22802_ (.Y(_05208_),
    .B1(net360),
    .B2(\cpu.dcache.r_data[5][11] ),
    .A2(net439),
    .A1(\cpu.dcache.r_data[1][11] ));
 sg13g2_buf_1 _22803_ (.A(_05031_),
    .X(_05209_));
 sg13g2_a22oi_1 _22804_ (.Y(_05210_),
    .B1(net394),
    .B2(\cpu.dcache.r_data[2][11] ),
    .A2(net413),
    .A1(\cpu.dcache.r_data[7][11] ));
 sg13g2_inv_1 _22805_ (.Y(_05211_),
    .A(_00113_));
 sg13g2_a22oi_1 _22806_ (.Y(_05212_),
    .B1(net436),
    .B2(_05211_),
    .A2(net399),
    .A1(\cpu.dcache.r_data[6][11] ));
 sg13g2_buf_1 _22807_ (.A(net438),
    .X(_05213_));
 sg13g2_a22oi_1 _22808_ (.Y(_05214_),
    .B1(net441),
    .B2(\cpu.dcache.r_data[4][11] ),
    .A2(_05213_),
    .A1(\cpu.dcache.r_data[3][11] ));
 sg13g2_nand4_1 _22809_ (.B(_05210_),
    .C(_05212_),
    .A(_05208_),
    .Y(_05215_),
    .D(_05214_));
 sg13g2_and2_1 _22810_ (.A(net673),
    .B(_05215_),
    .X(_05216_));
 sg13g2_a21o_1 _22811_ (.A2(_05207_),
    .A1(net615),
    .B1(_05216_),
    .X(_05217_));
 sg13g2_buf_1 _22812_ (.A(\cpu.intr.r_clock_count[27] ),
    .X(_05218_));
 sg13g2_a22oi_1 _22813_ (.Y(_05219_),
    .B1(net435),
    .B2(_10193_),
    .A2(net412),
    .A1(_05218_));
 sg13g2_a22oi_1 _22814_ (.Y(_05220_),
    .B1(net329),
    .B2(\cpu.intr.r_clock_cmp[11] ),
    .A2(net374),
    .A1(\cpu.intr.r_timer_reload[11] ));
 sg13g2_or2_1 _22815_ (.X(_05221_),
    .B(_05220_),
    .A(net617));
 sg13g2_a22oi_1 _22816_ (.Y(_05222_),
    .B1(_05187_),
    .B2(\cpu.intr.r_clock_cmp[27] ),
    .A2(_05185_),
    .A1(\cpu.intr.r_timer_count[11] ));
 sg13g2_nand3_1 _22817_ (.B(_05221_),
    .C(_05222_),
    .A(_05219_),
    .Y(_05223_));
 sg13g2_a221oi_1 _22818_ (.B2(_05176_),
    .C1(net1125),
    .B1(_05223_),
    .A1(_05123_),
    .Y(_05224_),
    .A2(_05217_));
 sg13g2_nor3_1 _22819_ (.A(_04884_),
    .B(_05159_),
    .C(_05224_),
    .Y(_05225_));
 sg13g2_a21oi_1 _22820_ (.A1(net1107),
    .A2(net78),
    .Y(_05226_),
    .B1(_05225_));
 sg13g2_nand2_1 _22821_ (.Y(_05227_),
    .A(_11540_),
    .B(_05226_));
 sg13g2_o21ai_1 _22822_ (.B1(_05227_),
    .Y(_05228_),
    .A1(\cpu.ex.pc[11] ),
    .A2(_05198_));
 sg13g2_a221oi_1 _22823_ (.B2(_05197_),
    .C1(_05228_),
    .B1(_05196_),
    .A1(_04337_),
    .Y(_01031_),
    .A2(_05074_));
 sg13g2_buf_1 _22824_ (.A(_04138_),
    .X(_05229_));
 sg13g2_nand3b_1 _22825_ (.B(net226),
    .C(net508),
    .Y(_05230_),
    .A_N(_04386_));
 sg13g2_o21ai_1 _22826_ (.B1(_05230_),
    .Y(_05231_),
    .A1(_08618_),
    .A2(net196));
 sg13g2_buf_1 _22827_ (.A(net191),
    .X(_05232_));
 sg13g2_buf_1 _22828_ (.A(\cpu.intr.r_clock_count[28] ),
    .X(_05233_));
 sg13g2_a22oi_1 _22829_ (.Y(_05234_),
    .B1(net435),
    .B2(_10200_),
    .A2(net373),
    .A1(_05233_));
 sg13g2_a22oi_1 _22830_ (.Y(_05235_),
    .B1(net329),
    .B2(\cpu.intr.r_clock_cmp[12] ),
    .A2(net335),
    .A1(\cpu.intr.r_timer_reload[12] ));
 sg13g2_or2_1 _22831_ (.X(_05236_),
    .B(_05235_),
    .A(net537));
 sg13g2_a22oi_1 _22832_ (.Y(_05237_),
    .B1(_05187_),
    .B2(\cpu.intr.r_clock_cmp[28] ),
    .A2(_05185_),
    .A1(\cpu.intr.r_timer_count[12] ));
 sg13g2_nand3_1 _22833_ (.B(_05236_),
    .C(_05237_),
    .A(_05234_),
    .Y(_05238_));
 sg13g2_a22oi_1 _22834_ (.Y(_05239_),
    .B1(net505),
    .B2(\cpu.dcache.r_data[1][28] ),
    .A2(net540),
    .A1(\cpu.dcache.r_data[7][28] ));
 sg13g2_a22oi_1 _22835_ (.Y(_05240_),
    .B1(net444),
    .B2(\cpu.dcache.r_data[5][28] ),
    .A2(_05026_),
    .A1(\cpu.dcache.r_data[3][28] ));
 sg13g2_inv_1 _22836_ (.Y(_05241_),
    .A(_00123_));
 sg13g2_a22oi_1 _22837_ (.Y(_05242_),
    .B1(_09641_),
    .B2(_05241_),
    .A2(_04975_),
    .A1(\cpu.dcache.r_data[6][28] ));
 sg13g2_a22oi_1 _22838_ (.Y(_05243_),
    .B1(net506),
    .B2(\cpu.dcache.r_data[4][28] ),
    .A2(_05030_),
    .A1(\cpu.dcache.r_data[2][28] ));
 sg13g2_nand4_1 _22839_ (.B(_05240_),
    .C(_05242_),
    .A(_05239_),
    .Y(_05244_),
    .D(_05243_));
 sg13g2_buf_1 _22840_ (.A(_05244_),
    .X(_05245_));
 sg13g2_a22oi_1 _22841_ (.Y(_05246_),
    .B1(net438),
    .B2(\cpu.dcache.r_data[3][12] ),
    .A2(net437),
    .A1(\cpu.dcache.r_data[2][12] ));
 sg13g2_a22oi_1 _22842_ (.Y(_05247_),
    .B1(_04928_),
    .B2(\cpu.dcache.r_data[5][12] ),
    .A2(net505),
    .A1(\cpu.dcache.r_data[1][12] ));
 sg13g2_inv_1 _22843_ (.Y(_05248_),
    .A(_00124_));
 sg13g2_a22oi_1 _22844_ (.Y(_05249_),
    .B1(net502),
    .B2(_05248_),
    .A2(net472),
    .A1(\cpu.dcache.r_data[7][12] ));
 sg13g2_a22oi_1 _22845_ (.Y(_05250_),
    .B1(net506),
    .B2(\cpu.dcache.r_data[4][12] ),
    .A2(net442),
    .A1(\cpu.dcache.r_data[6][12] ));
 sg13g2_nand4_1 _22846_ (.B(_05247_),
    .C(_05249_),
    .A(_05246_),
    .Y(_05251_),
    .D(_05250_));
 sg13g2_and2_1 _22847_ (.A(net673),
    .B(_05251_),
    .X(_05252_));
 sg13g2_a21o_1 _22848_ (.A2(_05245_),
    .A1(net538),
    .B1(_05252_),
    .X(_05253_));
 sg13g2_a22oi_1 _22849_ (.Y(_05254_),
    .B1(_05253_),
    .B2(_05160_),
    .A2(_05238_),
    .A1(_05176_));
 sg13g2_a21oi_1 _22850_ (.A1(_08583_),
    .A2(_05158_),
    .Y(_05255_),
    .B1(_11536_));
 sg13g2_buf_1 _22851_ (.A(_05255_),
    .X(_05256_));
 sg13g2_o21ai_1 _22852_ (.B1(_05256_),
    .Y(_05257_),
    .A1(net966),
    .A2(_05254_));
 sg13g2_nand2b_1 _22853_ (.Y(_05258_),
    .B(net83),
    .A_N(net620));
 sg13g2_o21ai_1 _22854_ (.B1(_05258_),
    .Y(_05259_),
    .A1(net83),
    .A2(_05257_));
 sg13g2_a221oi_1 _22855_ (.B2(net153),
    .C1(_05259_),
    .B1(_05231_),
    .A1(_04384_),
    .Y(_01032_),
    .A2(_05074_));
 sg13g2_a22oi_1 _22856_ (.Y(_05260_),
    .B1(_05209_),
    .B2(\cpu.dcache.r_data[2][29] ),
    .A2(_09995_),
    .A1(\cpu.dcache.r_data[7][29] ));
 sg13g2_a22oi_1 _22857_ (.Y(_05261_),
    .B1(net395),
    .B2(\cpu.dcache.r_data[5][29] ),
    .A2(net438),
    .A1(\cpu.dcache.r_data[3][29] ));
 sg13g2_a22oi_1 _22858_ (.Y(_05262_),
    .B1(net441),
    .B2(\cpu.dcache.r_data[4][29] ),
    .A2(_05017_),
    .A1(\cpu.dcache.r_data[1][29] ));
 sg13g2_inv_1 _22859_ (.Y(_05263_),
    .A(_00130_));
 sg13g2_a22oi_1 _22860_ (.Y(_05264_),
    .B1(net502),
    .B2(_05263_),
    .A2(net442),
    .A1(\cpu.dcache.r_data[6][29] ));
 sg13g2_nand4_1 _22861_ (.B(_05261_),
    .C(_05262_),
    .A(_05260_),
    .Y(_05265_),
    .D(_05264_));
 sg13g2_a22oi_1 _22862_ (.Y(_05266_),
    .B1(_04977_),
    .B2(\cpu.dcache.r_data[6][13] ),
    .A2(_05213_),
    .A1(\cpu.dcache.r_data[3][13] ));
 sg13g2_a22oi_1 _22863_ (.Y(_05267_),
    .B1(net360),
    .B2(\cpu.dcache.r_data[5][13] ),
    .A2(_05017_),
    .A1(\cpu.dcache.r_data[1][13] ));
 sg13g2_a22oi_1 _22864_ (.Y(_05268_),
    .B1(net441),
    .B2(\cpu.dcache.r_data[4][13] ),
    .A2(net394),
    .A1(\cpu.dcache.r_data[2][13] ));
 sg13g2_inv_1 _22865_ (.Y(_05269_),
    .A(_00131_));
 sg13g2_a22oi_1 _22866_ (.Y(_05270_),
    .B1(net436),
    .B2(_05269_),
    .A2(_09995_),
    .A1(\cpu.dcache.r_data[7][13] ));
 sg13g2_nand4_1 _22867_ (.B(_05267_),
    .C(_05268_),
    .A(_05266_),
    .Y(_05271_),
    .D(_05270_));
 sg13g2_mux2_1 _22868_ (.A0(_05265_),
    .A1(_05271_),
    .S(net616),
    .X(_05272_));
 sg13g2_and2_1 _22869_ (.A(_10206_),
    .B(net398),
    .X(_05273_));
 sg13g2_a221oi_1 _22870_ (.B2(\cpu.intr.r_clock_cmp[13] ),
    .C1(_05273_),
    .B1(net329),
    .A1(\cpu.intr.r_timer_reload[13] ),
    .Y(_05274_),
    .A2(net335));
 sg13g2_buf_1 _22871_ (.A(\cpu.intr.r_clock_count[29] ),
    .X(_05275_));
 sg13g2_and2_1 _22872_ (.A(\cpu.intr.r_timer_count[13] ),
    .B(_05185_),
    .X(_05276_));
 sg13g2_a221oi_1 _22873_ (.B2(\cpu.intr.r_clock_cmp[29] ),
    .C1(_05276_),
    .B1(_05187_),
    .A1(_05275_),
    .Y(_05277_),
    .A2(net373));
 sg13g2_o21ai_1 _22874_ (.B1(_05277_),
    .Y(_05278_),
    .A1(net537),
    .A2(_05274_));
 sg13g2_a22oi_1 _22875_ (.Y(_05279_),
    .B1(_05278_),
    .B2(_05176_),
    .A2(_05272_),
    .A1(net500));
 sg13g2_o21ai_1 _22876_ (.B1(_05256_),
    .Y(_05280_),
    .A1(net966),
    .A2(_05279_));
 sg13g2_mux2_1 _22877_ (.A0(_05280_),
    .A1(net614),
    .S(net83),
    .X(_05281_));
 sg13g2_o21ai_1 _22878_ (.B1(_05281_),
    .Y(_05282_),
    .A1(_08666_),
    .A2(_05198_));
 sg13g2_a21oi_1 _22879_ (.A1(net508),
    .A2(_04429_),
    .Y(_05283_),
    .B1(_05073_));
 sg13g2_o21ai_1 _22880_ (.B1(_05283_),
    .Y(_05284_),
    .A1(net508),
    .A2(_04427_));
 sg13g2_nor2b_1 _22881_ (.A(_05282_),
    .B_N(_05284_),
    .Y(_01033_));
 sg13g2_a22oi_1 _22882_ (.Y(_05285_),
    .B1(net398),
    .B2(_10210_),
    .A2(net335),
    .A1(\cpu.intr.r_timer_reload[14] ));
 sg13g2_buf_1 _22883_ (.A(\cpu.intr.r_clock_count[30] ),
    .X(_05286_));
 sg13g2_and2_1 _22884_ (.A(net900),
    .B(\cpu.intr.r_clock_cmp[30] ),
    .X(_05287_));
 sg13g2_a21oi_1 _22885_ (.A1(net763),
    .A2(\cpu.intr.r_clock_cmp[14] ),
    .Y(_05288_),
    .B1(_05287_));
 sg13g2_nor2_1 _22886_ (.A(net653),
    .B(_05288_),
    .Y(_05289_));
 sg13g2_a221oi_1 _22887_ (.B2(\cpu.intr.r_timer_count[14] ),
    .C1(_05289_),
    .B1(_05185_),
    .A1(_05286_),
    .Y(_05290_),
    .A2(net412));
 sg13g2_o21ai_1 _22888_ (.B1(_05290_),
    .Y(_05291_),
    .A1(net615),
    .A2(_05285_));
 sg13g2_a22oi_1 _22889_ (.Y(_05292_),
    .B1(_05016_),
    .B2(\cpu.dcache.r_data[1][30] ),
    .A2(net472),
    .A1(\cpu.dcache.r_data[7][30] ));
 sg13g2_a22oi_1 _22890_ (.Y(_05293_),
    .B1(net395),
    .B2(\cpu.dcache.r_data[5][30] ),
    .A2(net438),
    .A1(\cpu.dcache.r_data[3][30] ));
 sg13g2_inv_1 _22891_ (.Y(_05294_),
    .A(_00142_));
 sg13g2_a22oi_1 _22892_ (.Y(_05295_),
    .B1(net502),
    .B2(_05294_),
    .A2(_04976_),
    .A1(\cpu.dcache.r_data[6][30] ));
 sg13g2_a22oi_1 _22893_ (.Y(_05296_),
    .B1(net441),
    .B2(\cpu.dcache.r_data[4][30] ),
    .A2(net437),
    .A1(\cpu.dcache.r_data[2][30] ));
 sg13g2_nand4_1 _22894_ (.B(_05293_),
    .C(_05295_),
    .A(_05292_),
    .Y(_05297_),
    .D(_05296_));
 sg13g2_a22oi_1 _22895_ (.Y(_05298_),
    .B1(net506),
    .B2(\cpu.dcache.r_data[4][14] ),
    .A2(_05016_),
    .A1(\cpu.dcache.r_data[1][14] ));
 sg13g2_a22oi_1 _22896_ (.Y(_05299_),
    .B1(_05026_),
    .B2(\cpu.dcache.r_data[3][14] ),
    .A2(net503),
    .A1(\cpu.dcache.r_data[2][14] ));
 sg13g2_a22oi_1 _22897_ (.Y(_05300_),
    .B1(net444),
    .B2(\cpu.dcache.r_data[5][14] ),
    .A2(net507),
    .A1(\cpu.dcache.r_data[6][14] ));
 sg13g2_inv_1 _22898_ (.Y(_05301_),
    .A(_00143_));
 sg13g2_a22oi_1 _22899_ (.Y(_05302_),
    .B1(net619),
    .B2(_05301_),
    .A2(net472),
    .A1(\cpu.dcache.r_data[7][14] ));
 sg13g2_nand4_1 _22900_ (.B(_05299_),
    .C(_05300_),
    .A(_05298_),
    .Y(_05303_),
    .D(_05302_));
 sg13g2_mux2_1 _22901_ (.A0(_05297_),
    .A1(_05303_),
    .S(net673),
    .X(_05304_));
 sg13g2_a22oi_1 _22902_ (.Y(_05305_),
    .B1(_05304_),
    .B2(_05123_),
    .A2(_05291_),
    .A1(_05176_));
 sg13g2_nor2_1 _22903_ (.A(net1125),
    .B(_05305_),
    .Y(_05306_));
 sg13g2_nor2b_1 _22904_ (.A(_05306_),
    .B_N(_05256_),
    .Y(_05307_));
 sg13g2_or4_1 _22905_ (.A(net508),
    .B(net83),
    .C(net197),
    .D(_05307_),
    .X(_05308_));
 sg13g2_buf_1 _22906_ (.A(_11540_),
    .X(_05309_));
 sg13g2_buf_1 _22907_ (.A(_04884_),
    .X(_05310_));
 sg13g2_nand2_1 _22908_ (.Y(_05311_),
    .A(net605),
    .B(net78));
 sg13g2_o21ai_1 _22909_ (.B1(_05311_),
    .Y(_05312_),
    .A1(_05310_),
    .A2(_05307_));
 sg13g2_nor2_1 _22910_ (.A(net581),
    .B(_04251_),
    .Y(_05313_));
 sg13g2_a22oi_1 _22911_ (.Y(_05314_),
    .B1(_04466_),
    .B2(_05313_),
    .A2(net197),
    .A1(net915));
 sg13g2_nor2_1 _22912_ (.A(_11540_),
    .B(_05314_),
    .Y(_05315_));
 sg13g2_a21oi_1 _22913_ (.A1(_05309_),
    .A2(_05312_),
    .Y(_05316_),
    .B1(_05315_));
 sg13g2_o21ai_1 _22914_ (.B1(_05316_),
    .Y(_01034_),
    .A1(_04464_),
    .A2(_05308_));
 sg13g2_nor2_1 _22915_ (.A(net581),
    .B(_04499_),
    .Y(_05317_));
 sg13g2_buf_1 _22916_ (.A(\cpu.intr.r_clock_count[31] ),
    .X(_05318_));
 sg13g2_a22oi_1 _22917_ (.Y(_05319_),
    .B1(net435),
    .B2(_10217_),
    .A2(net373),
    .A1(_05318_));
 sg13g2_a22oi_1 _22918_ (.Y(_05320_),
    .B1(net329),
    .B2(\cpu.intr.r_clock_cmp[15] ),
    .A2(net374),
    .A1(\cpu.intr.r_timer_reload[15] ));
 sg13g2_or2_1 _22919_ (.X(_05321_),
    .B(_05320_),
    .A(net617));
 sg13g2_a22oi_1 _22920_ (.Y(_05322_),
    .B1(_05187_),
    .B2(\cpu.intr.r_clock_cmp[31] ),
    .A2(_05185_),
    .A1(\cpu.intr.r_timer_count[15] ));
 sg13g2_nand3_1 _22921_ (.B(_05321_),
    .C(_05322_),
    .A(_05319_),
    .Y(_05323_));
 sg13g2_mux2_1 _22922_ (.A0(_05145_),
    .A1(_05151_),
    .S(net615),
    .X(_05324_));
 sg13g2_a22oi_1 _22923_ (.Y(_05325_),
    .B1(_05324_),
    .B2(net500),
    .A2(_05323_),
    .A1(_05176_));
 sg13g2_o21ai_1 _22924_ (.B1(_05256_),
    .Y(_05326_),
    .A1(_08583_),
    .A2(_05325_));
 sg13g2_nor2_1 _22925_ (.A(_03634_),
    .B(_05326_),
    .Y(_05327_));
 sg13g2_a21oi_1 _22926_ (.A1(net676),
    .A2(net83),
    .Y(_05328_),
    .B1(_05327_));
 sg13g2_o21ai_1 _22927_ (.B1(_05328_),
    .Y(_05329_),
    .A1(_08538_),
    .A2(_05198_));
 sg13g2_a221oi_1 _22928_ (.B2(_05197_),
    .C1(_05329_),
    .B1(_05317_),
    .A1(_04497_),
    .Y(_01035_),
    .A2(_05074_));
 sg13g2_nand2_1 _22929_ (.Y(_05330_),
    .A(_11110_),
    .B(_11528_));
 sg13g2_o21ai_1 _22930_ (.B1(_05330_),
    .Y(_05331_),
    .A1(net584),
    .A2(_04249_));
 sg13g2_nand2_1 _22931_ (.Y(_05332_),
    .A(net196),
    .B(_05331_));
 sg13g2_o21ai_1 _22932_ (.B1(_05332_),
    .Y(_05333_),
    .A1(net923),
    .A2(net196));
 sg13g2_buf_1 _22933_ (.A(net191),
    .X(_05334_));
 sg13g2_inv_1 _22934_ (.Y(_05335_),
    .A(_00095_));
 sg13g2_buf_1 _22935_ (.A(_04952_),
    .X(_05336_));
 sg13g2_buf_1 _22936_ (.A(\cpu.spi.r_clk_count[2][1] ),
    .X(_05337_));
 sg13g2_a22oi_1 _22937_ (.Y(_05338_),
    .B1(_04964_),
    .B2(_05337_),
    .A2(net392),
    .A1(_05335_));
 sg13g2_mux2_1 _22938_ (.A0(_11939_),
    .A1(_11938_),
    .S(net858),
    .X(_05339_));
 sg13g2_a22oi_1 _22939_ (.Y(_05340_),
    .B1(_05339_),
    .B2(net447),
    .A2(_05082_),
    .A1(\cpu.spi.r_timeout[1] ));
 sg13g2_or2_1 _22940_ (.X(_05341_),
    .B(_04967_),
    .A(_00094_));
 sg13g2_nand3_1 _22941_ (.B(_05340_),
    .C(_05341_),
    .A(_05338_),
    .Y(_05342_));
 sg13g2_a221oi_1 _22942_ (.B2(_09319_),
    .C1(_05342_),
    .B1(_04954_),
    .A1(_11942_),
    .Y(_05343_),
    .A2(net445));
 sg13g2_nand2b_1 _22943_ (.Y(_05344_),
    .B(_05077_),
    .A_N(_05343_));
 sg13g2_inv_1 _22944_ (.Y(_05345_),
    .A(\cpu.intr.r_clock ));
 sg13g2_buf_1 _22945_ (.A(_04982_),
    .X(_05346_));
 sg13g2_a21oi_1 _22946_ (.A1(_09251_),
    .A2(net396),
    .Y(_05347_),
    .B1(_05346_));
 sg13g2_a22oi_1 _22947_ (.Y(_05348_),
    .B1(net329),
    .B2(\cpu.intr.r_clock_cmp[1] ),
    .A2(net361),
    .A1(_09968_));
 sg13g2_a221oi_1 _22948_ (.B2(\cpu.intr.r_clock_cmp[17] ),
    .C1(net763),
    .B1(net360),
    .A1(\cpu.intr.r_timer_reload[17] ),
    .Y(_05349_),
    .A2(net374));
 sg13g2_a21oi_1 _22949_ (.A1(net673),
    .A2(_05348_),
    .Y(_05350_),
    .B1(_05349_));
 sg13g2_nand2_1 _22950_ (.Y(_05351_),
    .A(_10129_),
    .B(net501));
 sg13g2_buf_2 _22951_ (.A(\cpu.intr.r_clock_count[17] ),
    .X(_05352_));
 sg13g2_a22oi_1 _22952_ (.Y(_05353_),
    .B1(_04993_),
    .B2(_09251_),
    .A2(net412),
    .A1(_05352_));
 sg13g2_nand3_1 _22953_ (.B(\cpu.intr.r_timer_reload[1] ),
    .C(net374),
    .A(net763),
    .Y(_05354_));
 sg13g2_nand3_1 _22954_ (.B(_09964_),
    .C(_04978_),
    .A(net674),
    .Y(_05355_));
 sg13g2_nand4_1 _22955_ (.B(_05353_),
    .C(_05354_),
    .A(_05351_),
    .Y(_05356_),
    .D(_05355_));
 sg13g2_nor2_1 _22956_ (.A(_05350_),
    .B(_05356_),
    .Y(_05357_));
 sg13g2_o21ai_1 _22957_ (.B1(_05357_),
    .Y(_05358_),
    .A1(_05345_),
    .A2(_05347_));
 sg13g2_nand3_1 _22958_ (.B(_09226_),
    .C(_04903_),
    .A(_09225_),
    .Y(_05359_));
 sg13g2_nand2b_1 _22959_ (.Y(_05360_),
    .B(_04931_),
    .A_N(_00100_));
 sg13g2_buf_2 _22960_ (.A(\cpu.gpio.r_src_io[4][1] ),
    .X(_05361_));
 sg13g2_nand2_1 _22961_ (.Y(_05362_),
    .A(net858),
    .B(net440));
 sg13g2_nand2b_1 _22962_ (.Y(_05363_),
    .B(net446),
    .A_N(_00096_));
 sg13g2_o21ai_1 _22963_ (.B1(_05363_),
    .Y(_05364_),
    .A1(_00097_),
    .A2(_05362_));
 sg13g2_a221oi_1 _22964_ (.B2(_05361_),
    .C1(_05364_),
    .B1(net443),
    .A1(_09226_),
    .Y(_05365_),
    .A2(_04918_));
 sg13g2_inv_1 _22965_ (.Y(_05366_),
    .A(_00099_));
 sg13g2_nor2_1 _22966_ (.A(_00098_),
    .B(_05095_),
    .Y(_05367_));
 sg13g2_a221oi_1 _22967_ (.B2(_09225_),
    .C1(_05367_),
    .B1(net362),
    .A1(_05366_),
    .Y(_05368_),
    .A2(net445));
 sg13g2_nand4_1 _22968_ (.B(_05360_),
    .C(_05365_),
    .A(_05359_),
    .Y(_05369_),
    .D(_05368_));
 sg13g2_a22oi_1 _22969_ (.Y(_05370_),
    .B1(net440),
    .B2(\cpu.uart.r_r_invert ),
    .A2(net397),
    .A1(_09249_));
 sg13g2_a22oi_1 _22970_ (.Y(_05371_),
    .B1(net447),
    .B2(\cpu.uart.r_div_value[1] ),
    .A2(_04957_),
    .A1(\cpu.uart.r_div_value[9] ));
 sg13g2_nand2_1 _22971_ (.Y(_05372_),
    .A(_05370_),
    .B(_05371_));
 sg13g2_a21oi_1 _22972_ (.A1(\cpu.uart.r_in[1] ),
    .A2(_05005_),
    .Y(_05373_),
    .B1(_05372_));
 sg13g2_o21ai_1 _22973_ (.B1(net1041),
    .Y(_05374_),
    .A1(net582),
    .A2(_05373_));
 sg13g2_a221oi_1 _22974_ (.B2(_04888_),
    .C1(_05374_),
    .B1(_05369_),
    .A1(_10059_),
    .Y(_05375_),
    .A2(_05358_));
 sg13g2_a22oi_1 _22975_ (.Y(_05376_),
    .B1(_04976_),
    .B2(\cpu.dcache.r_data[6][25] ),
    .A2(net439),
    .A1(\cpu.dcache.r_data[1][25] ));
 sg13g2_a22oi_1 _22976_ (.Y(_05377_),
    .B1(_05031_),
    .B2(\cpu.dcache.r_data[2][25] ),
    .A2(net413),
    .A1(\cpu.dcache.r_data[7][25] ));
 sg13g2_inv_1 _22977_ (.Y(_05378_),
    .A(_00092_));
 sg13g2_a22oi_1 _22978_ (.Y(_05379_),
    .B1(_05044_),
    .B2(_05378_),
    .A2(net395),
    .A1(\cpu.dcache.r_data[5][25] ));
 sg13g2_a22oi_1 _22979_ (.Y(_05380_),
    .B1(_04988_),
    .B2(\cpu.dcache.r_data[4][25] ),
    .A2(_05027_),
    .A1(\cpu.dcache.r_data[3][25] ));
 sg13g2_nand4_1 _22980_ (.B(_05377_),
    .C(_05379_),
    .A(_05376_),
    .Y(_05381_),
    .D(_05380_));
 sg13g2_buf_1 _22981_ (.A(net439),
    .X(_05382_));
 sg13g2_a22oi_1 _22982_ (.Y(_05383_),
    .B1(_04977_),
    .B2(\cpu.dcache.r_data[6][9] ),
    .A2(net390),
    .A1(\cpu.dcache.r_data[1][9] ));
 sg13g2_a22oi_1 _22983_ (.Y(_05384_),
    .B1(net360),
    .B2(\cpu.dcache.r_data[5][9] ),
    .A2(_05209_),
    .A1(\cpu.dcache.r_data[2][9] ));
 sg13g2_inv_1 _22984_ (.Y(_05385_),
    .A(_00093_));
 sg13g2_a22oi_1 _22985_ (.Y(_05386_),
    .B1(net398),
    .B2(\cpu.dcache.r_data[4][9] ),
    .A2(net436),
    .A1(_05385_));
 sg13g2_a22oi_1 _22986_ (.Y(_05387_),
    .B1(net393),
    .B2(\cpu.dcache.r_data[3][9] ),
    .A2(net413),
    .A1(\cpu.dcache.r_data[7][9] ));
 sg13g2_nand4_1 _22987_ (.B(_05384_),
    .C(_05386_),
    .A(_05383_),
    .Y(_05388_),
    .D(_05387_));
 sg13g2_and2_1 _22988_ (.A(_10053_),
    .B(_05388_),
    .X(_05389_));
 sg13g2_a21oi_1 _22989_ (.A1(net997),
    .A2(_05381_),
    .Y(_05390_),
    .B1(_05389_));
 sg13g2_a22oi_1 _22990_ (.Y(_05391_),
    .B1(net399),
    .B2(\cpu.dcache.r_data[6][17] ),
    .A2(net393),
    .A1(\cpu.dcache.r_data[3][17] ));
 sg13g2_a22oi_1 _22991_ (.Y(_05392_),
    .B1(net360),
    .B2(\cpu.dcache.r_data[5][17] ),
    .A2(_05382_),
    .A1(\cpu.dcache.r_data[1][17] ));
 sg13g2_a22oi_1 _22992_ (.Y(_05393_),
    .B1(net398),
    .B2(\cpu.dcache.r_data[4][17] ),
    .A2(net394),
    .A1(\cpu.dcache.r_data[2][17] ));
 sg13g2_inv_1 _22993_ (.Y(_05394_),
    .A(_00091_));
 sg13g2_a22oi_1 _22994_ (.Y(_05395_),
    .B1(net436),
    .B2(_05394_),
    .A2(net413),
    .A1(\cpu.dcache.r_data[7][17] ));
 sg13g2_nand4_1 _22995_ (.B(_05392_),
    .C(_05393_),
    .A(_05391_),
    .Y(_05396_),
    .D(_05395_));
 sg13g2_buf_1 _22996_ (.A(_05396_),
    .X(_05397_));
 sg13g2_a22oi_1 _22997_ (.Y(_05398_),
    .B1(net438),
    .B2(\cpu.dcache.r_data[3][1] ),
    .A2(_09994_),
    .A1(\cpu.dcache.r_data[7][1] ));
 sg13g2_a22oi_1 _22998_ (.Y(_05399_),
    .B1(net506),
    .B2(\cpu.dcache.r_data[4][1] ),
    .A2(net437),
    .A1(\cpu.dcache.r_data[2][1] ));
 sg13g2_a22oi_1 _22999_ (.Y(_05400_),
    .B1(_04928_),
    .B2(\cpu.dcache.r_data[5][1] ),
    .A2(net507),
    .A1(\cpu.dcache.r_data[6][1] ));
 sg13g2_nand3_1 _23000_ (.B(_05399_),
    .C(_05400_),
    .A(_05398_),
    .Y(_05401_));
 sg13g2_nand2b_1 _23001_ (.Y(_05402_),
    .B(net895),
    .A_N(\cpu.dcache.r_data[0][1] ));
 sg13g2_o21ai_1 _23002_ (.B1(_05402_),
    .Y(_05403_),
    .A1(net895),
    .A2(_05401_));
 sg13g2_o21ai_1 _23003_ (.B1(net390),
    .Y(_05404_),
    .A1(\cpu.dcache.r_data[1][1] ),
    .A2(_05401_));
 sg13g2_o21ai_1 _23004_ (.B1(_05404_),
    .Y(_05405_),
    .A1(net390),
    .A2(_05403_));
 sg13g2_buf_1 _23005_ (.A(_12016_),
    .X(_05406_));
 sg13g2_a221oi_1 _23006_ (.B2(net959),
    .C1(net717),
    .B1(_05405_),
    .A1(_05138_),
    .Y(_05407_),
    .A2(_05397_));
 sg13g2_a21oi_1 _23007_ (.A1(net717),
    .A2(_05390_),
    .Y(_05408_),
    .B1(_05407_));
 sg13g2_nand2_1 _23008_ (.Y(_05409_),
    .A(_10106_),
    .B(_05397_));
 sg13g2_nand2_1 _23009_ (.Y(_05410_),
    .A(net616),
    .B(_05405_));
 sg13g2_a21oi_1 _23010_ (.A1(_05409_),
    .A2(_05410_),
    .Y(_05411_),
    .B1(_05041_));
 sg13g2_a21oi_1 _23011_ (.A1(_05041_),
    .A2(_05408_),
    .Y(_05412_),
    .B1(_05411_));
 sg13g2_a221oi_1 _23012_ (.B2(net1058),
    .C1(net78),
    .B1(_05412_),
    .A1(_05344_),
    .Y(_05413_),
    .A2(_05375_));
 sg13g2_a21oi_1 _23013_ (.A1(net538),
    .A2(net77),
    .Y(_05414_),
    .B1(_05413_));
 sg13g2_nor2_1 _23014_ (.A(net151),
    .B(_05414_),
    .Y(_05415_));
 sg13g2_a21o_1 _23015_ (.A2(_05333_),
    .A1(net153),
    .B1(_05415_),
    .X(_01036_));
 sg13g2_buf_1 _23016_ (.A(net152),
    .X(_05416_));
 sg13g2_a22oi_1 _23017_ (.Y(_05417_),
    .B1(net441),
    .B2(\cpu.dcache.r_data[4][2] ),
    .A2(net438),
    .A1(\cpu.dcache.r_data[3][2] ));
 sg13g2_a22oi_1 _23018_ (.Y(_05418_),
    .B1(net437),
    .B2(\cpu.dcache.r_data[2][2] ),
    .A2(net439),
    .A1(\cpu.dcache.r_data[1][2] ));
 sg13g2_a22oi_1 _23019_ (.Y(_05419_),
    .B1(net395),
    .B2(\cpu.dcache.r_data[5][2] ),
    .A2(net442),
    .A1(\cpu.dcache.r_data[6][2] ));
 sg13g2_a22oi_1 _23020_ (.Y(_05420_),
    .B1(net502),
    .B2(\cpu.dcache.r_data[0][2] ),
    .A2(_09994_),
    .A1(\cpu.dcache.r_data[7][2] ));
 sg13g2_nand4_1 _23021_ (.B(_05418_),
    .C(_05419_),
    .A(_05417_),
    .Y(_05421_),
    .D(_05420_));
 sg13g2_a22oi_1 _23022_ (.Y(_05422_),
    .B1(net394),
    .B2(\cpu.dcache.r_data[2][18] ),
    .A2(net413),
    .A1(\cpu.dcache.r_data[7][18] ));
 sg13g2_a22oi_1 _23023_ (.Y(_05423_),
    .B1(net399),
    .B2(\cpu.dcache.r_data[6][18] ),
    .A2(net393),
    .A1(\cpu.dcache.r_data[3][18] ));
 sg13g2_inv_1 _23024_ (.Y(_05424_),
    .A(_00101_));
 sg13g2_a22oi_1 _23025_ (.Y(_05425_),
    .B1(net502),
    .B2(_05424_),
    .A2(net395),
    .A1(\cpu.dcache.r_data[5][18] ));
 sg13g2_a22oi_1 _23026_ (.Y(_05426_),
    .B1(net441),
    .B2(\cpu.dcache.r_data[4][18] ),
    .A2(net439),
    .A1(\cpu.dcache.r_data[1][18] ));
 sg13g2_nand4_1 _23027_ (.B(_05423_),
    .C(_05425_),
    .A(_05422_),
    .Y(_05427_),
    .D(_05426_));
 sg13g2_mux2_1 _23028_ (.A0(_05421_),
    .A1(_05427_),
    .S(net538),
    .X(_05428_));
 sg13g2_a221oi_1 _23029_ (.B2(_05138_),
    .C1(net717),
    .B1(_05427_),
    .A1(net959),
    .Y(_05429_),
    .A2(_05421_));
 sg13g2_a221oi_1 _23030_ (.B2(_12039_),
    .C1(_05063_),
    .B1(_05173_),
    .A1(net616),
    .Y(_05430_),
    .A2(_05166_));
 sg13g2_o21ai_1 _23031_ (.B1(_05041_),
    .Y(_05431_),
    .A1(_05429_),
    .A2(_05430_));
 sg13g2_o21ai_1 _23032_ (.B1(_05431_),
    .Y(_05432_),
    .A1(_05041_),
    .A2(_05428_));
 sg13g2_and2_1 _23033_ (.A(_09323_),
    .B(_04954_),
    .X(_05433_));
 sg13g2_inv_1 _23034_ (.Y(_05434_),
    .A(_00105_));
 sg13g2_buf_1 _23035_ (.A(_04957_),
    .X(_05435_));
 sg13g2_buf_1 _23036_ (.A(net447),
    .X(_05436_));
 sg13g2_nor3_1 _23037_ (.A(net617),
    .B(_00281_),
    .C(_02739_),
    .Y(_05437_));
 sg13g2_a221oi_1 _23038_ (.B2(_11928_),
    .C1(_05437_),
    .B1(_05436_),
    .A1(_05434_),
    .Y(_05438_),
    .A2(_05435_));
 sg13g2_buf_1 _23039_ (.A(\cpu.spi.r_clk_count[2][2] ),
    .X(_05439_));
 sg13g2_and2_1 _23040_ (.A(net858),
    .B(_11932_),
    .X(_05440_));
 sg13g2_a22oi_1 _23041_ (.Y(_05441_),
    .B1(_05440_),
    .B2(net447),
    .A2(_05082_),
    .A1(\cpu.spi.r_timeout[2] ));
 sg13g2_o21ai_1 _23042_ (.B1(_05441_),
    .Y(_05442_),
    .A1(_00104_),
    .A2(_04967_));
 sg13g2_a21oi_1 _23043_ (.A1(_05439_),
    .A2(_04964_),
    .Y(_05443_),
    .B1(_05442_));
 sg13g2_o21ai_1 _23044_ (.B1(_05443_),
    .Y(_05444_),
    .A1(net735),
    .A2(_05438_));
 sg13g2_o21ai_1 _23045_ (.B1(_05077_),
    .Y(_05445_),
    .A1(_05433_),
    .A2(_05444_));
 sg13g2_nand2b_1 _23046_ (.Y(_05446_),
    .B(_04903_),
    .A_N(_09216_));
 sg13g2_inv_1 _23047_ (.Y(_05447_),
    .A(_00108_));
 sg13g2_buf_1 _23048_ (.A(\cpu.gpio.r_src_io[4][2] ),
    .X(_05448_));
 sg13g2_a22oi_1 _23049_ (.Y(_05449_),
    .B1(net443),
    .B2(_05448_),
    .A2(_04914_),
    .A1(_05447_));
 sg13g2_a22oi_1 _23050_ (.Y(_05450_),
    .B1(_04918_),
    .B2(_09215_),
    .A2(net362),
    .A1(\cpu.gpio.r_enable_in[2] ));
 sg13g2_inv_1 _23051_ (.Y(_05451_),
    .A(_00109_));
 sg13g2_inv_1 _23052_ (.Y(_05452_),
    .A(_00110_));
 sg13g2_nand2b_1 _23053_ (.Y(_05453_),
    .B(net446),
    .A_N(_00106_));
 sg13g2_o21ai_1 _23054_ (.B1(_05453_),
    .Y(_05454_),
    .A1(_00107_),
    .A2(_05362_));
 sg13g2_a221oi_1 _23055_ (.B2(_05452_),
    .C1(_05454_),
    .B1(_04931_),
    .A1(_05451_),
    .Y(_05455_),
    .A2(net445));
 sg13g2_nand4_1 _23056_ (.B(_05449_),
    .C(_05450_),
    .A(_05446_),
    .Y(_05456_),
    .D(_05455_));
 sg13g2_mux2_1 _23057_ (.A0(\cpu.intr.r_timer_count[2] ),
    .A1(_09963_),
    .S(net617),
    .X(_05457_));
 sg13g2_nand2_1 _23058_ (.Y(_05458_),
    .A(net361),
    .B(_05457_));
 sg13g2_mux2_1 _23059_ (.A0(\cpu.intr.r_clock_cmp[2] ),
    .A1(\cpu.intr.r_clock_cmp[18] ),
    .S(net617),
    .X(_05459_));
 sg13g2_a22oi_1 _23060_ (.Y(_05460_),
    .B1(_05459_),
    .B2(net329),
    .A2(net391),
    .A1(_09245_));
 sg13g2_buf_2 _23061_ (.A(\cpu.intr.r_clock_count[18] ),
    .X(_05461_));
 sg13g2_nand2_1 _23062_ (.Y(_05462_),
    .A(net674),
    .B(\cpu.intr.r_timer_reload[18] ));
 sg13g2_nand2_1 _23063_ (.Y(_05463_),
    .A(net673),
    .B(\cpu.intr.r_timer_reload[2] ));
 sg13g2_a21oi_1 _23064_ (.A1(_05462_),
    .A2(_05463_),
    .Y(_05464_),
    .B1(net539));
 sg13g2_a221oi_1 _23065_ (.B2(_10142_),
    .C1(_05464_),
    .B1(net435),
    .A1(_05461_),
    .Y(_05465_),
    .A2(net373));
 sg13g2_a21oi_1 _23066_ (.A1(_09245_),
    .A2(net396),
    .Y(_05466_),
    .B1(net397));
 sg13g2_nand2b_1 _23067_ (.Y(_05467_),
    .B(\cpu.intr.r_enable[2] ),
    .A_N(_05466_));
 sg13g2_nand4_1 _23068_ (.B(_05460_),
    .C(_05465_),
    .A(_05458_),
    .Y(_05468_),
    .D(_05467_));
 sg13g2_and2_1 _23069_ (.A(\cpu.uart.r_in[2] ),
    .B(_05005_),
    .X(_05469_));
 sg13g2_a221oi_1 _23070_ (.B2(\cpu.uart.r_div_value[2] ),
    .C1(_05469_),
    .B1(net388),
    .A1(_09952_),
    .Y(_05470_),
    .A2(net389));
 sg13g2_o21ai_1 _23071_ (.B1(net848),
    .Y(_05471_),
    .A1(net582),
    .A2(_05470_));
 sg13g2_a221oi_1 _23072_ (.B2(_10059_),
    .C1(_05471_),
    .B1(_05468_),
    .A1(_04888_),
    .Y(_05472_),
    .A2(_05456_));
 sg13g2_a221oi_1 _23073_ (.B2(_05472_),
    .C1(net77),
    .B1(_05445_),
    .A1(net1058),
    .Y(_05473_),
    .A2(_05432_));
 sg13g2_a21oi_1 _23074_ (.A1(net596),
    .A2(net77),
    .Y(_05474_),
    .B1(_05473_));
 sg13g2_o21ai_1 _23075_ (.B1(net226),
    .Y(_05475_),
    .A1(net794),
    .A2(_05195_));
 sg13g2_nor3_1 _23076_ (.A(net701),
    .B(net923),
    .C(net581),
    .Y(_05476_));
 sg13g2_a21o_1 _23077_ (.A2(_04535_),
    .A1(net581),
    .B1(_05476_),
    .X(_05477_));
 sg13g2_a221oi_1 _23078_ (.B2(net196),
    .C1(_05309_),
    .B1(_05477_),
    .A1(net701),
    .Y(_05478_),
    .A2(_05475_));
 sg13g2_a21oi_1 _23079_ (.A1(net121),
    .A2(_05474_),
    .Y(_01037_),
    .B1(_05478_));
 sg13g2_and2_1 _23080_ (.A(net794),
    .B(net704),
    .X(_05479_));
 sg13g2_mux2_1 _23081_ (.A0(_05479_),
    .A1(_04571_),
    .S(net581),
    .X(_05480_));
 sg13g2_nand2_1 _23082_ (.Y(_05481_),
    .A(net584),
    .B(_04572_));
 sg13g2_a21oi_1 _23083_ (.A1(net196),
    .A2(_05481_),
    .Y(_05482_),
    .B1(net702));
 sg13g2_a21oi_1 _23084_ (.A1(_05229_),
    .A2(_05480_),
    .Y(_05483_),
    .B1(_05482_));
 sg13g2_nand2_1 _23085_ (.Y(_05484_),
    .A(net997),
    .B(_05207_));
 sg13g2_nor2_1 _23086_ (.A(_05063_),
    .B(_05216_),
    .Y(_05485_));
 sg13g2_mux2_1 _23087_ (.A0(\cpu.dcache.r_data[1][3] ),
    .A1(\cpu.dcache.r_data[3][3] ),
    .S(net696),
    .X(_05486_));
 sg13g2_a22oi_1 _23088_ (.Y(_05487_),
    .B1(_05486_),
    .B2(net695),
    .A2(_09732_),
    .A1(\cpu.dcache.r_data[2][3] ));
 sg13g2_nor2_1 _23089_ (.A(_05199_),
    .B(_05487_),
    .Y(_05488_));
 sg13g2_mux2_1 _23090_ (.A0(\cpu.dcache.r_data[5][3] ),
    .A1(\cpu.dcache.r_data[7][3] ),
    .S(net696),
    .X(_05489_));
 sg13g2_a22oi_1 _23091_ (.Y(_05490_),
    .B1(_05489_),
    .B2(net695),
    .A2(_09557_),
    .A1(\cpu.dcache.r_data[4][3] ));
 sg13g2_a22oi_1 _23092_ (.Y(_05491_),
    .B1(net502),
    .B2(\cpu.dcache.r_data[0][3] ),
    .A2(net442),
    .A1(\cpu.dcache.r_data[6][3] ));
 sg13g2_o21ai_1 _23093_ (.B1(_05491_),
    .Y(_05492_),
    .A1(net733),
    .A2(_05490_));
 sg13g2_nor2_1 _23094_ (.A(_05488_),
    .B(_05492_),
    .Y(_05493_));
 sg13g2_a22oi_1 _23095_ (.Y(_05494_),
    .B1(net507),
    .B2(\cpu.dcache.r_data[6][19] ),
    .A2(net503),
    .A1(\cpu.dcache.r_data[2][19] ));
 sg13g2_a22oi_1 _23096_ (.Y(_05495_),
    .B1(net506),
    .B2(\cpu.dcache.r_data[4][19] ),
    .A2(net504),
    .A1(\cpu.dcache.r_data[3][19] ));
 sg13g2_a22oi_1 _23097_ (.Y(_05496_),
    .B1(net444),
    .B2(\cpu.dcache.r_data[5][19] ),
    .A2(net472),
    .A1(\cpu.dcache.r_data[7][19] ));
 sg13g2_nand3_1 _23098_ (.B(_05495_),
    .C(_05496_),
    .A(_05494_),
    .Y(_05497_));
 sg13g2_nand2_1 _23099_ (.Y(_05498_),
    .A(_00111_),
    .B(net895));
 sg13g2_o21ai_1 _23100_ (.B1(_05498_),
    .Y(_05499_),
    .A1(net895),
    .A2(_05497_));
 sg13g2_o21ai_1 _23101_ (.B1(net390),
    .Y(_05500_),
    .A1(\cpu.dcache.r_data[1][19] ),
    .A2(_05497_));
 sg13g2_o21ai_1 _23102_ (.B1(_05500_),
    .Y(_05501_),
    .A1(net390),
    .A2(_05499_));
 sg13g2_nand2_1 _23103_ (.Y(_05502_),
    .A(net997),
    .B(_05063_));
 sg13g2_a22oi_1 _23104_ (.Y(_05503_),
    .B1(_05502_),
    .B2(_05041_),
    .A2(_05501_),
    .A1(_09993_));
 sg13g2_a221oi_1 _23105_ (.B2(_05066_),
    .C1(_05503_),
    .B1(_05493_),
    .A1(_05484_),
    .Y(_05504_),
    .A2(_05485_));
 sg13g2_o21ai_1 _23106_ (.B1(_05503_),
    .Y(_05505_),
    .A1(net537),
    .A2(_05493_));
 sg13g2_o21ai_1 _23107_ (.B1(_05505_),
    .Y(_05506_),
    .A1(net500),
    .A2(_05504_));
 sg13g2_inv_1 _23108_ (.Y(_05507_),
    .A(_00115_));
 sg13g2_buf_1 _23109_ (.A(\cpu.spi.r_clk_count[2][3] ),
    .X(_05508_));
 sg13g2_a22oi_1 _23110_ (.Y(_05509_),
    .B1(_04964_),
    .B2(_05508_),
    .A2(net392),
    .A1(_05507_));
 sg13g2_nor2_1 _23111_ (.A(_00114_),
    .B(_04967_),
    .Y(_05510_));
 sg13g2_a21oi_1 _23112_ (.A1(\cpu.spi.r_timeout[3] ),
    .A2(_05082_),
    .Y(_05511_),
    .B1(_05510_));
 sg13g2_nand2_1 _23113_ (.Y(_05512_),
    .A(_09317_),
    .B(_04954_));
 sg13g2_nand3_1 _23114_ (.B(_05511_),
    .C(_05512_),
    .A(_05509_),
    .Y(_05513_));
 sg13g2_nand2_1 _23115_ (.Y(_05514_),
    .A(_05077_),
    .B(_05513_));
 sg13g2_nand2b_1 _23116_ (.Y(_05515_),
    .B(net446),
    .A_N(_00116_));
 sg13g2_nor2_1 _23117_ (.A(net858),
    .B(net782),
    .Y(_05516_));
 sg13g2_nor3_1 _23118_ (.A(net862),
    .B(net763),
    .C(_00117_),
    .Y(_05517_));
 sg13g2_a21oi_1 _23119_ (.A1(_09230_),
    .A2(_05516_),
    .Y(_05518_),
    .B1(_05517_));
 sg13g2_nand3b_1 _23120_ (.B(net895),
    .C(net695),
    .Y(_05519_),
    .A_N(_05518_));
 sg13g2_nand2_1 _23121_ (.Y(_05520_),
    .A(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .B(net501));
 sg13g2_o21ai_1 _23122_ (.B1(_05520_),
    .Y(_05521_),
    .A1(_00119_),
    .A2(_04929_));
 sg13g2_buf_1 _23123_ (.A(\cpu.gpio.r_src_io[4][3] ),
    .X(_05522_));
 sg13g2_a22oi_1 _23124_ (.Y(_05523_),
    .B1(net443),
    .B2(_05522_),
    .A2(net362),
    .A1(_09229_));
 sg13g2_o21ai_1 _23125_ (.B1(_05523_),
    .Y(_05524_),
    .A1(_00118_),
    .A2(_05095_));
 sg13g2_a21oi_1 _23126_ (.A1(net960),
    .A2(_05521_),
    .Y(_05525_),
    .B1(_05524_));
 sg13g2_nand3_1 _23127_ (.B(_09230_),
    .C(_04903_),
    .A(_09229_),
    .Y(_05526_));
 sg13g2_nand4_1 _23128_ (.B(_05519_),
    .C(_05525_),
    .A(_05515_),
    .Y(_05527_),
    .D(_05526_));
 sg13g2_a21o_1 _23129_ (.A2(net361),
    .A1(_09962_),
    .B1(net673),
    .X(_05528_));
 sg13g2_a221oi_1 _23130_ (.B2(\cpu.intr.r_clock_cmp[19] ),
    .C1(_05528_),
    .B1(_05181_),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .Y(_05529_),
    .A2(_09997_));
 sg13g2_a21oi_1 _23131_ (.A1(\cpu.intr.r_timer_reload[3] ),
    .A2(net335),
    .Y(_05530_),
    .B1(net615));
 sg13g2_buf_1 _23132_ (.A(\cpu.intr.r_clock_count[19] ),
    .X(_05531_));
 sg13g2_nand2_1 _23133_ (.Y(_05532_),
    .A(_10147_),
    .B(net501));
 sg13g2_nor2_1 _23134_ (.A(net900),
    .B(net653),
    .Y(_05533_));
 sg13g2_buf_1 _23135_ (.A(_05533_),
    .X(_05534_));
 sg13g2_a22oi_1 _23136_ (.Y(_05535_),
    .B1(net499),
    .B2(\cpu.intr.r_clock_cmp[3] ),
    .A2(_05185_),
    .A1(\cpu.intr.r_timer_count[3] ));
 sg13g2_a21oi_1 _23137_ (.A1(_09246_),
    .A2(net396),
    .Y(_05536_),
    .B1(net391));
 sg13g2_nand2b_1 _23138_ (.Y(_05537_),
    .B(\cpu.intr.r_swi ),
    .A_N(_05536_));
 sg13g2_nand3_1 _23139_ (.B(_05535_),
    .C(_05537_),
    .A(_05532_),
    .Y(_05538_));
 sg13g2_a221oi_1 _23140_ (.B2(_09246_),
    .C1(_05538_),
    .B1(net397),
    .A1(_05531_),
    .Y(_05539_),
    .A2(_10124_));
 sg13g2_o21ai_1 _23141_ (.B1(_05539_),
    .Y(_05540_),
    .A1(_05529_),
    .A2(_05530_));
 sg13g2_and2_1 _23142_ (.A(\cpu.uart.r_in[3] ),
    .B(_05005_),
    .X(_05541_));
 sg13g2_a221oi_1 _23143_ (.B2(\cpu.uart.r_div_value[3] ),
    .C1(_05541_),
    .B1(net388),
    .A1(\cpu.uart.r_div_value[11] ),
    .Y(_05542_),
    .A2(net389));
 sg13g2_o21ai_1 _23144_ (.B1(net1041),
    .Y(_05543_),
    .A1(net582),
    .A2(_05542_));
 sg13g2_a221oi_1 _23145_ (.B2(_10059_),
    .C1(_05543_),
    .B1(_05540_),
    .A1(_04888_),
    .Y(_05544_),
    .A2(_05527_));
 sg13g2_a221oi_1 _23146_ (.B2(_05544_),
    .C1(net78),
    .B1(_05514_),
    .A1(net1058),
    .Y(_05545_),
    .A2(_05506_));
 sg13g2_a21oi_1 _23147_ (.A1(net632),
    .A2(_05310_),
    .Y(_05546_),
    .B1(_05545_));
 sg13g2_nor2_1 _23148_ (.A(net191),
    .B(_05546_),
    .Y(_05547_));
 sg13g2_a21o_1 _23149_ (.A2(_05483_),
    .A1(_05232_),
    .B1(_05547_),
    .X(_01038_));
 sg13g2_o21ai_1 _23150_ (.B1(net196),
    .Y(_05548_),
    .A1(net581),
    .A2(_05479_));
 sg13g2_nand2_1 _23151_ (.Y(_05549_),
    .A(net584),
    .B(_04607_));
 sg13g2_o21ai_1 _23152_ (.B1(_05549_),
    .Y(_05550_),
    .A1(net508),
    .A2(_04606_));
 sg13g2_a22oi_1 _23153_ (.Y(_05551_),
    .B1(_05550_),
    .B2(_05229_),
    .A2(_05548_),
    .A1(_08264_));
 sg13g2_a21oi_1 _23154_ (.A1(net1060),
    .A2(_11544_),
    .Y(_05552_),
    .B1(net650));
 sg13g2_mux2_1 _23155_ (.A0(\cpu.intr.r_timer_count[4] ),
    .A1(_09986_),
    .S(net782),
    .X(_05553_));
 sg13g2_mux2_1 _23156_ (.A0(\cpu.intr.r_clock_cmp[4] ),
    .A1(\cpu.intr.r_clock_cmp[20] ),
    .S(net782),
    .X(_05554_));
 sg13g2_a22oi_1 _23157_ (.Y(_05555_),
    .B1(_05554_),
    .B2(net329),
    .A2(_05553_),
    .A1(net361));
 sg13g2_mux2_1 _23158_ (.A0(\cpu.intr.r_timer_reload[4] ),
    .A1(\cpu.intr.r_timer_reload[20] ),
    .S(_09287_),
    .X(_05556_));
 sg13g2_a22oi_1 _23159_ (.Y(_05557_),
    .B1(_05556_),
    .B2(net335),
    .A2(net397),
    .A1(_09214_));
 sg13g2_buf_1 _23160_ (.A(\cpu.intr.r_clock_count[20] ),
    .X(_05558_));
 sg13g2_a22oi_1 _23161_ (.Y(_05559_),
    .B1(net435),
    .B2(_10153_),
    .A2(net412),
    .A1(_05558_));
 sg13g2_o21ai_1 _23162_ (.B1(_09244_),
    .Y(_05560_),
    .A1(_05346_),
    .A2(net396));
 sg13g2_nand4_1 _23163_ (.B(_05557_),
    .C(_05559_),
    .A(_05555_),
    .Y(_05561_),
    .D(_05560_));
 sg13g2_inv_1 _23164_ (.Y(_05562_),
    .A(_09214_));
 sg13g2_a21oi_1 _23165_ (.A1(_05562_),
    .A2(net396),
    .Y(_05563_),
    .B1(_10001_));
 sg13g2_nand2_1 _23166_ (.Y(_05564_),
    .A(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .B(net501));
 sg13g2_a22oi_1 _23167_ (.Y(_05565_),
    .B1(net499),
    .B2(net7),
    .A2(_10122_),
    .A1(\cpu.gpio.genblk2[4].srcs_io[0] ));
 sg13g2_a21oi_1 _23168_ (.A1(_09238_),
    .A2(_04982_),
    .Y(_05566_),
    .B1(net440));
 sg13g2_nand2b_1 _23169_ (.Y(_05567_),
    .B(_09239_),
    .A_N(_05566_));
 sg13g2_nand3_1 _23170_ (.B(_05565_),
    .C(_05567_),
    .A(_05564_),
    .Y(_05568_));
 sg13g2_nand3_1 _23171_ (.B(_09234_),
    .C(_04903_),
    .A(_09233_),
    .Y(_05569_));
 sg13g2_buf_2 _23172_ (.A(\cpu.gpio.r_src_o[3][0] ),
    .X(_05570_));
 sg13g2_nand3_1 _23173_ (.B(_05570_),
    .C(_04982_),
    .A(_09999_),
    .Y(_05571_));
 sg13g2_nand3_1 _23174_ (.B(net862),
    .C(_04957_),
    .A(_09238_),
    .Y(_05572_));
 sg13g2_buf_2 _23175_ (.A(\cpu.gpio.r_spi_miso_src[1][0] ),
    .X(_05573_));
 sg13g2_nand2_1 _23176_ (.Y(_05574_),
    .A(_05573_),
    .B(_04931_));
 sg13g2_buf_2 _23177_ (.A(\cpu.gpio.r_src_o[7][0] ),
    .X(_05575_));
 sg13g2_buf_2 _23178_ (.A(\cpu.gpio.r_src_io[5][0] ),
    .X(_05576_));
 sg13g2_a22oi_1 _23179_ (.Y(_05577_),
    .B1(net443),
    .B2(_05576_),
    .A2(_04934_),
    .A1(_05575_));
 sg13g2_and4_1 _23180_ (.A(_05571_),
    .B(_05572_),
    .C(_05574_),
    .D(_05577_),
    .X(_05578_));
 sg13g2_a22oi_1 _23181_ (.Y(_05579_),
    .B1(_04918_),
    .B2(_09234_),
    .A2(net362),
    .A1(_09233_));
 sg13g2_buf_2 _23182_ (.A(\cpu.gpio.r_src_o[5][0] ),
    .X(_05580_));
 sg13g2_buf_2 _23183_ (.A(\cpu.gpio.r_src_io[7][0] ),
    .X(_05581_));
 sg13g2_a22oi_1 _23184_ (.Y(_05582_),
    .B1(net446),
    .B2(_05581_),
    .A2(_04914_),
    .A1(_05580_));
 sg13g2_nand4_1 _23185_ (.B(_05578_),
    .C(_05579_),
    .A(_05569_),
    .Y(_05583_),
    .D(_05582_));
 sg13g2_a21o_1 _23186_ (.A2(_05568_),
    .A1(net960),
    .B1(_05583_),
    .X(_05584_));
 sg13g2_inv_1 _23187_ (.Y(_05585_),
    .A(_00126_));
 sg13g2_buf_1 _23188_ (.A(\cpu.spi.r_clk_count[2][4] ),
    .X(_05586_));
 sg13g2_nand2_1 _23189_ (.Y(_05587_),
    .A(\cpu.spi.r_timeout[4] ),
    .B(_05082_));
 sg13g2_o21ai_1 _23190_ (.B1(_05587_),
    .Y(_05588_),
    .A1(_00125_),
    .A2(_04967_));
 sg13g2_a221oi_1 _23191_ (.B2(_05586_),
    .C1(_05588_),
    .B1(_04964_),
    .A1(_05585_),
    .Y(_05589_),
    .A2(net392));
 sg13g2_nand2_1 _23192_ (.Y(_05590_),
    .A(_09325_),
    .B(_04954_));
 sg13g2_a21oi_1 _23193_ (.A1(_05589_),
    .A2(_05590_),
    .Y(_05591_),
    .B1(_09208_));
 sg13g2_a221oi_1 _23194_ (.B2(_04888_),
    .C1(_05591_),
    .B1(_05584_),
    .A1(_05561_),
    .Y(_05592_),
    .A2(_05563_));
 sg13g2_a221oi_1 _23195_ (.B2(\cpu.uart.r_in[4] ),
    .C1(net582),
    .B1(_05005_),
    .A1(\cpu.uart.r_div_value[4] ),
    .Y(_05593_),
    .A2(net388));
 sg13g2_a21oi_1 _23196_ (.A1(_05003_),
    .A2(_05592_),
    .Y(_05594_),
    .B1(_05593_));
 sg13g2_o21ai_1 _23197_ (.B1(_05065_),
    .Y(_05595_),
    .A1(_05038_),
    .A2(_05252_));
 sg13g2_a22oi_1 _23198_ (.Y(_05596_),
    .B1(net393),
    .B2(\cpu.dcache.r_data[3][4] ),
    .A2(net394),
    .A1(\cpu.dcache.r_data[2][4] ));
 sg13g2_a22oi_1 _23199_ (.Y(_05597_),
    .B1(_05180_),
    .B2(\cpu.dcache.r_data[5][4] ),
    .A2(net390),
    .A1(\cpu.dcache.r_data[1][4] ));
 sg13g2_inv_1 _23200_ (.Y(_05598_),
    .A(_00121_));
 sg13g2_a22oi_1 _23201_ (.Y(_05599_),
    .B1(net436),
    .B2(_05598_),
    .A2(net399),
    .A1(\cpu.dcache.r_data[6][4] ));
 sg13g2_a22oi_1 _23202_ (.Y(_05600_),
    .B1(net398),
    .B2(\cpu.dcache.r_data[4][4] ),
    .A2(net374),
    .A1(\cpu.dcache.r_data[7][4] ));
 sg13g2_nand4_1 _23203_ (.B(_05597_),
    .C(_05599_),
    .A(_05596_),
    .Y(_05601_),
    .D(_05600_));
 sg13g2_buf_1 _23204_ (.A(_05601_),
    .X(_05602_));
 sg13g2_a22oi_1 _23205_ (.Y(_05603_),
    .B1(net507),
    .B2(\cpu.dcache.r_data[6][20] ),
    .A2(net504),
    .A1(\cpu.dcache.r_data[3][20] ));
 sg13g2_a22oi_1 _23206_ (.Y(_05604_),
    .B1(net541),
    .B2(\cpu.dcache.r_data[5][20] ),
    .A2(net505),
    .A1(\cpu.dcache.r_data[1][20] ));
 sg13g2_a22oi_1 _23207_ (.Y(_05605_),
    .B1(net506),
    .B2(\cpu.dcache.r_data[4][20] ),
    .A2(net503),
    .A1(\cpu.dcache.r_data[2][20] ));
 sg13g2_inv_1 _23208_ (.Y(_05606_),
    .A(_00122_));
 sg13g2_a22oi_1 _23209_ (.Y(_05607_),
    .B1(net619),
    .B2(_05606_),
    .A2(net540),
    .A1(\cpu.dcache.r_data[7][20] ));
 sg13g2_and4_1 _23210_ (.A(_05603_),
    .B(_05604_),
    .C(_05605_),
    .D(_05607_),
    .X(_05608_));
 sg13g2_buf_1 _23211_ (.A(_05608_),
    .X(_05609_));
 sg13g2_inv_1 _23212_ (.Y(_05610_),
    .A(_05609_));
 sg13g2_nor2_1 _23213_ (.A(_10052_),
    .B(net717),
    .Y(_05611_));
 sg13g2_a22oi_1 _23214_ (.Y(_05612_),
    .B1(_05610_),
    .B2(_05611_),
    .A2(_05245_),
    .A1(_05065_));
 sg13g2_nor2_1 _23215_ (.A(net959),
    .B(_05612_),
    .Y(_05613_));
 sg13g2_a21oi_1 _23216_ (.A1(_05066_),
    .A2(_05602_),
    .Y(_05614_),
    .B1(_05613_));
 sg13g2_nand2_1 _23217_ (.Y(_05615_),
    .A(net537),
    .B(_05609_));
 sg13g2_o21ai_1 _23218_ (.B1(_05615_),
    .Y(_05616_),
    .A1(net537),
    .A2(_05602_));
 sg13g2_a221oi_1 _23219_ (.B2(net500),
    .C1(net848),
    .B1(_05616_),
    .A1(_05595_),
    .Y(_05617_),
    .A2(_05614_));
 sg13g2_a21oi_1 _23220_ (.A1(net848),
    .A2(_05594_),
    .Y(_05618_),
    .B1(_05617_));
 sg13g2_nor2_1 _23221_ (.A(net77),
    .B(_05618_),
    .Y(_05619_));
 sg13g2_o21ai_1 _23222_ (.B1(net152),
    .Y(_05620_),
    .A1(_05552_),
    .A2(_05619_));
 sg13g2_o21ai_1 _23223_ (.B1(_05620_),
    .Y(_01039_),
    .A1(_05416_),
    .A2(_05551_));
 sg13g2_buf_2 _23224_ (.A(\cpu.intr.r_clock_count[21] ),
    .X(_05621_));
 sg13g2_inv_1 _23225_ (.Y(_05622_),
    .A(\cpu.intr.r_timer_reload[21] ));
 sg13g2_nor2_1 _23226_ (.A(net889),
    .B(_05622_),
    .Y(_05623_));
 sg13g2_a21oi_1 _23227_ (.A1(net763),
    .A2(\cpu.intr.r_timer_reload[5] ),
    .Y(_05624_),
    .B1(_05623_));
 sg13g2_nor2_1 _23228_ (.A(net539),
    .B(_05624_),
    .Y(_05625_));
 sg13g2_a221oi_1 _23229_ (.B2(_10159_),
    .C1(_05625_),
    .B1(net501),
    .A1(_05621_),
    .Y(_05626_),
    .A2(net412));
 sg13g2_mux2_1 _23230_ (.A0(\cpu.intr.r_timer_count[5] ),
    .A1(_09985_),
    .S(_09287_),
    .X(_05627_));
 sg13g2_a22oi_1 _23231_ (.Y(_05628_),
    .B1(_05627_),
    .B2(net361),
    .A2(_04994_),
    .A1(_09253_));
 sg13g2_mux2_1 _23232_ (.A0(\cpu.intr.r_clock_cmp[5] ),
    .A1(\cpu.intr.r_clock_cmp[21] ),
    .S(net782),
    .X(_05629_));
 sg13g2_a22oi_1 _23233_ (.Y(_05630_),
    .B1(_05629_),
    .B2(_05181_),
    .A2(net391),
    .A1(_09252_));
 sg13g2_nand3_1 _23234_ (.B(_09253_),
    .C(net396),
    .A(_09252_),
    .Y(_05631_));
 sg13g2_nand4_1 _23235_ (.B(_05628_),
    .C(_05630_),
    .A(_05626_),
    .Y(_05632_),
    .D(_05631_));
 sg13g2_nand3_1 _23236_ (.B(_09236_),
    .C(_04903_),
    .A(_09235_),
    .Y(_05633_));
 sg13g2_nand2_1 _23237_ (.Y(_05634_),
    .A(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .B(_05100_));
 sg13g2_a22oi_1 _23238_ (.Y(_05635_),
    .B1(net499),
    .B2(net8),
    .A2(_10122_),
    .A1(\cpu.gpio.genblk2[5].srcs_io[0] ));
 sg13g2_a21oi_1 _23239_ (.A1(_09240_),
    .A2(_04982_),
    .Y(_05636_),
    .B1(net440));
 sg13g2_nand2b_1 _23240_ (.Y(_05637_),
    .B(_09241_),
    .A_N(_05636_));
 sg13g2_nand3_1 _23241_ (.B(_05635_),
    .C(_05637_),
    .A(_05634_),
    .Y(_05638_));
 sg13g2_nand2b_1 _23242_ (.Y(_05639_),
    .B(_04931_),
    .A_N(_00138_));
 sg13g2_inv_1 _23243_ (.Y(_05640_),
    .A(_00134_));
 sg13g2_a22oi_1 _23244_ (.Y(_05641_),
    .B1(net446),
    .B2(_05640_),
    .A2(net362),
    .A1(_09235_));
 sg13g2_nand2b_1 _23245_ (.Y(_05642_),
    .B(_05007_),
    .A_N(_00135_));
 sg13g2_o21ai_1 _23246_ (.B1(_05642_),
    .Y(_05643_),
    .A1(_00137_),
    .A2(_05089_));
 sg13g2_nor2_1 _23247_ (.A(_00136_),
    .B(_05095_),
    .Y(_05644_));
 sg13g2_a221oi_1 _23248_ (.B2(_11925_),
    .C1(_05644_),
    .B1(_05643_),
    .A1(_09236_),
    .Y(_05645_),
    .A2(_04918_));
 sg13g2_buf_2 _23249_ (.A(\cpu.gpio.r_src_io[5][1] ),
    .X(_05646_));
 sg13g2_a22oi_1 _23250_ (.Y(_05647_),
    .B1(_04936_),
    .B2(_05646_),
    .A2(_04952_),
    .A1(_09240_));
 sg13g2_nand4_1 _23251_ (.B(_05641_),
    .C(_05645_),
    .A(_05639_),
    .Y(_05648_),
    .D(_05647_));
 sg13g2_a21oi_1 _23252_ (.A1(_04911_),
    .A2(_05638_),
    .Y(_05649_),
    .B1(_05648_));
 sg13g2_nand2_1 _23253_ (.Y(_05650_),
    .A(_05633_),
    .B(_05649_));
 sg13g2_inv_1 _23254_ (.Y(_05651_),
    .A(_00133_));
 sg13g2_buf_1 _23255_ (.A(\cpu.spi.r_clk_count[2][5] ),
    .X(_05652_));
 sg13g2_nand2_1 _23256_ (.Y(_05653_),
    .A(\cpu.spi.r_timeout[5] ),
    .B(_05082_));
 sg13g2_o21ai_1 _23257_ (.B1(_05653_),
    .Y(_05654_),
    .A1(_00132_),
    .A2(_04967_));
 sg13g2_a221oi_1 _23258_ (.B2(_05652_),
    .C1(_05654_),
    .B1(_04964_),
    .A1(_05651_),
    .Y(_05655_),
    .A2(_04952_));
 sg13g2_nand2_1 _23259_ (.Y(_05656_),
    .A(_09324_),
    .B(_04954_));
 sg13g2_a21oi_1 _23260_ (.A1(_05655_),
    .A2(_05656_),
    .Y(_05657_),
    .B1(_09208_));
 sg13g2_a221oi_1 _23261_ (.B2(_04888_),
    .C1(_05657_),
    .B1(_05650_),
    .A1(_10059_),
    .Y(_05658_),
    .A2(_05632_));
 sg13g2_a221oi_1 _23262_ (.B2(\cpu.uart.r_in[5] ),
    .C1(net582),
    .B1(_05005_),
    .A1(\cpu.uart.r_div_value[5] ),
    .Y(_05659_),
    .A2(net388));
 sg13g2_a21oi_1 _23263_ (.A1(_05003_),
    .A2(_05658_),
    .Y(_05660_),
    .B1(_05659_));
 sg13g2_a21oi_1 _23264_ (.A1(net616),
    .A2(_05271_),
    .Y(_05661_),
    .B1(_05038_));
 sg13g2_nand2b_1 _23265_ (.Y(_05662_),
    .B(net717),
    .A_N(_05661_));
 sg13g2_a22oi_1 _23266_ (.Y(_05663_),
    .B1(net390),
    .B2(\cpu.dcache.r_data[1][5] ),
    .A2(_09996_),
    .A1(\cpu.dcache.r_data[7][5] ));
 sg13g2_a22oi_1 _23267_ (.Y(_05664_),
    .B1(_04978_),
    .B2(\cpu.dcache.r_data[6][5] ),
    .A2(net394),
    .A1(\cpu.dcache.r_data[2][5] ));
 sg13g2_inv_1 _23268_ (.Y(_05665_),
    .A(_00128_));
 sg13g2_a22oi_1 _23269_ (.Y(_05666_),
    .B1(net436),
    .B2(_05665_),
    .A2(net360),
    .A1(\cpu.dcache.r_data[5][5] ));
 sg13g2_a22oi_1 _23270_ (.Y(_05667_),
    .B1(net398),
    .B2(\cpu.dcache.r_data[4][5] ),
    .A2(net393),
    .A1(\cpu.dcache.r_data[3][5] ));
 sg13g2_nand4_1 _23271_ (.B(_05664_),
    .C(_05666_),
    .A(_05663_),
    .Y(_05668_),
    .D(_05667_));
 sg13g2_buf_1 _23272_ (.A(_05668_),
    .X(_05669_));
 sg13g2_a22oi_1 _23273_ (.Y(_05670_),
    .B1(net399),
    .B2(\cpu.dcache.r_data[6][21] ),
    .A2(net393),
    .A1(\cpu.dcache.r_data[3][21] ));
 sg13g2_a22oi_1 _23274_ (.Y(_05671_),
    .B1(_05180_),
    .B2(\cpu.dcache.r_data[5][21] ),
    .A2(_05382_),
    .A1(\cpu.dcache.r_data[1][21] ));
 sg13g2_a22oi_1 _23275_ (.Y(_05672_),
    .B1(_04989_),
    .B2(\cpu.dcache.r_data[4][21] ),
    .A2(net394),
    .A1(\cpu.dcache.r_data[2][21] ));
 sg13g2_inv_1 _23276_ (.Y(_05673_),
    .A(_00129_));
 sg13g2_a22oi_1 _23277_ (.Y(_05674_),
    .B1(net436),
    .B2(_05673_),
    .A2(net413),
    .A1(\cpu.dcache.r_data[7][21] ));
 sg13g2_nand4_1 _23278_ (.B(_05671_),
    .C(_05672_),
    .A(_05670_),
    .Y(_05675_),
    .D(_05674_));
 sg13g2_buf_1 _23279_ (.A(_05675_),
    .X(_05676_));
 sg13g2_a22oi_1 _23280_ (.Y(_05677_),
    .B1(_05611_),
    .B2(_05676_),
    .A2(_05265_),
    .A1(net717));
 sg13g2_nor2_1 _23281_ (.A(net959),
    .B(_05677_),
    .Y(_05678_));
 sg13g2_a21oi_1 _23282_ (.A1(_05066_),
    .A2(_05669_),
    .Y(_05679_),
    .B1(_05678_));
 sg13g2_or2_1 _23283_ (.X(_05680_),
    .B(_05676_),
    .A(net616));
 sg13g2_o21ai_1 _23284_ (.B1(_05680_),
    .Y(_05681_),
    .A1(net537),
    .A2(_05669_));
 sg13g2_a221oi_1 _23285_ (.B2(net500),
    .C1(net848),
    .B1(_05681_),
    .A1(_05662_),
    .Y(_05682_),
    .A2(_05679_));
 sg13g2_a21oi_1 _23286_ (.A1(net848),
    .A2(_05660_),
    .Y(_05683_),
    .B1(_05682_));
 sg13g2_nor2_1 _23287_ (.A(net77),
    .B(_05683_),
    .Y(_05684_));
 sg13g2_a21oi_1 _23288_ (.A1(net598),
    .A2(net77),
    .Y(_05685_),
    .B1(_05684_));
 sg13g2_nand2_1 _23289_ (.Y(_05686_),
    .A(net584),
    .B(_04645_));
 sg13g2_o21ai_1 _23290_ (.B1(_05686_),
    .Y(_05687_),
    .A1(net584),
    .A2(_04643_));
 sg13g2_mux2_1 _23291_ (.A0(net964),
    .A1(_05687_),
    .S(net226),
    .X(_05688_));
 sg13g2_nand2_1 _23292_ (.Y(_05689_),
    .A(net151),
    .B(_05688_));
 sg13g2_o21ai_1 _23293_ (.B1(_05689_),
    .Y(_01040_),
    .A1(net153),
    .A2(_05685_));
 sg13g2_nand2_1 _23294_ (.Y(_05690_),
    .A(net584),
    .B(_04677_));
 sg13g2_o21ai_1 _23295_ (.B1(_05690_),
    .Y(_05691_),
    .A1(_04858_),
    .A2(_04674_));
 sg13g2_and2_1 _23296_ (.A(net963),
    .B(_04860_),
    .X(_05692_));
 sg13g2_a21oi_1 _23297_ (.A1(net196),
    .A2(_05691_),
    .Y(_05693_),
    .B1(_05692_));
 sg13g2_buf_1 _23298_ (.A(_11540_),
    .X(_05694_));
 sg13g2_a22oi_1 _23299_ (.Y(_05695_),
    .B1(net360),
    .B2(\cpu.dcache.r_data[5][6] ),
    .A2(net393),
    .A1(\cpu.dcache.r_data[3][6] ));
 sg13g2_a22oi_1 _23300_ (.Y(_05696_),
    .B1(net399),
    .B2(\cpu.dcache.r_data[6][6] ),
    .A2(net394),
    .A1(\cpu.dcache.r_data[2][6] ));
 sg13g2_a22oi_1 _23301_ (.Y(_05697_),
    .B1(net398),
    .B2(\cpu.dcache.r_data[4][6] ),
    .A2(net390),
    .A1(\cpu.dcache.r_data[1][6] ));
 sg13g2_inv_1 _23302_ (.Y(_05698_),
    .A(_00140_));
 sg13g2_a22oi_1 _23303_ (.Y(_05699_),
    .B1(net436),
    .B2(_05698_),
    .A2(_09996_),
    .A1(\cpu.dcache.r_data[7][6] ));
 sg13g2_nand4_1 _23304_ (.B(_05696_),
    .C(_05697_),
    .A(_05695_),
    .Y(_05700_),
    .D(_05699_));
 sg13g2_a22oi_1 _23305_ (.Y(_05701_),
    .B1(net442),
    .B2(\cpu.dcache.r_data[6][22] ),
    .A2(net393),
    .A1(\cpu.dcache.r_data[3][22] ));
 sg13g2_a22oi_1 _23306_ (.Y(_05702_),
    .B1(net395),
    .B2(\cpu.dcache.r_data[5][22] ),
    .A2(net439),
    .A1(\cpu.dcache.r_data[1][22] ));
 sg13g2_a22oi_1 _23307_ (.Y(_05703_),
    .B1(net441),
    .B2(\cpu.dcache.r_data[4][22] ),
    .A2(net437),
    .A1(\cpu.dcache.r_data[2][22] ));
 sg13g2_inv_1 _23308_ (.Y(_05704_),
    .A(_00141_));
 sg13g2_a22oi_1 _23309_ (.Y(_05705_),
    .B1(net502),
    .B2(_05704_),
    .A2(net413),
    .A1(\cpu.dcache.r_data[7][22] ));
 sg13g2_nand4_1 _23310_ (.B(_05702_),
    .C(_05703_),
    .A(_05701_),
    .Y(_05706_),
    .D(_05705_));
 sg13g2_mux2_1 _23311_ (.A0(_05700_),
    .A1(_05706_),
    .S(_10106_),
    .X(_05707_));
 sg13g2_a221oi_1 _23312_ (.B2(_05138_),
    .C1(net717),
    .B1(_05706_),
    .A1(_12016_),
    .Y(_05708_),
    .A2(_05700_));
 sg13g2_a221oi_1 _23313_ (.B2(_10053_),
    .C1(_05063_),
    .B1(_05303_),
    .A1(net997),
    .Y(_05709_),
    .A2(_05297_));
 sg13g2_nor3_1 _23314_ (.A(_05123_),
    .B(_05708_),
    .C(_05709_),
    .Y(_05710_));
 sg13g2_a21o_1 _23315_ (.A2(_05707_),
    .A1(net500),
    .B1(_05710_),
    .X(_05711_));
 sg13g2_inv_1 _23316_ (.Y(_05712_),
    .A(_00150_));
 sg13g2_a22oi_1 _23317_ (.Y(_05713_),
    .B1(_05178_),
    .B2(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .A2(_05187_),
    .A1(_05712_));
 sg13g2_a22oi_1 _23318_ (.Y(_05714_),
    .B1(_05534_),
    .B2(net9),
    .A2(_10123_),
    .A1(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_a21oi_1 _23319_ (.A1(_05713_),
    .A2(_05714_),
    .Y(_05715_),
    .B1(net1034));
 sg13g2_nand3_1 _23320_ (.B(_09222_),
    .C(_04903_),
    .A(_09221_),
    .Y(_05716_));
 sg13g2_and3_1 _23321_ (.X(_05717_),
    .A(_09231_),
    .B(net960),
    .C(net391));
 sg13g2_o21ai_1 _23322_ (.B1(\cpu.gpio.r_enable_io[6] ),
    .Y(_05718_),
    .A1(net392),
    .A2(_05717_));
 sg13g2_inv_1 _23323_ (.Y(_05719_),
    .A(_00146_));
 sg13g2_buf_1 _23324_ (.A(\cpu.gpio.r_src_io[5][2] ),
    .X(_05720_));
 sg13g2_nand2_1 _23325_ (.Y(_05721_),
    .A(_05720_),
    .B(net443));
 sg13g2_o21ai_1 _23326_ (.B1(_05721_),
    .Y(_05722_),
    .A1(_00148_),
    .A2(_05095_));
 sg13g2_a221oi_1 _23327_ (.B2(_05719_),
    .C1(_05722_),
    .B1(_04922_),
    .A1(_09221_),
    .Y(_05723_),
    .A2(_04910_));
 sg13g2_nand2b_1 _23328_ (.Y(_05724_),
    .B(_05008_),
    .A_N(_00147_));
 sg13g2_o21ai_1 _23329_ (.B1(_05724_),
    .Y(_05725_),
    .A1(_00149_),
    .A2(_05089_));
 sg13g2_and3_1 _23330_ (.X(_05726_),
    .A(_09231_),
    .B(_04911_),
    .C(_05008_));
 sg13g2_a221oi_1 _23331_ (.B2(_11925_),
    .C1(_05726_),
    .B1(_05725_),
    .A1(_09222_),
    .Y(_05727_),
    .A2(_04918_));
 sg13g2_nand4_1 _23332_ (.B(_05718_),
    .C(_05723_),
    .A(_05716_),
    .Y(_05728_),
    .D(_05727_));
 sg13g2_o21ai_1 _23333_ (.B1(_04888_),
    .Y(_05729_),
    .A1(_05715_),
    .A2(_05728_));
 sg13g2_a22oi_1 _23334_ (.Y(_05730_),
    .B1(_05005_),
    .B2(\cpu.uart.r_in[6] ),
    .A2(net388),
    .A1(\cpu.uart.r_div_value[6] ));
 sg13g2_or2_1 _23335_ (.X(_05731_),
    .B(_05730_),
    .A(net582));
 sg13g2_mux2_1 _23336_ (.A0(_10165_),
    .A1(\cpu.intr.r_timer_count[6] ),
    .S(net632),
    .X(_05732_));
 sg13g2_a22oi_1 _23337_ (.Y(_05733_),
    .B1(_05732_),
    .B2(net767),
    .A2(_09521_),
    .A1(\cpu.intr.r_timer_reload[6] ));
 sg13g2_mux2_1 _23338_ (.A0(\cpu.intr.r_clock_cmp[22] ),
    .A1(\cpu.intr.r_timer_reload[22] ),
    .S(net632),
    .X(_05734_));
 sg13g2_a221oi_1 _23339_ (.B2(net695),
    .C1(net763),
    .B1(_05734_),
    .A1(_09988_),
    .Y(_05735_),
    .A2(_09732_));
 sg13g2_a21o_1 _23340_ (.A2(_05733_),
    .A1(net673),
    .B1(_05735_),
    .X(_05736_));
 sg13g2_buf_1 _23341_ (.A(\cpu.intr.r_clock_count[22] ),
    .X(_05737_));
 sg13g2_a22oi_1 _23342_ (.Y(_05738_),
    .B1(net499),
    .B2(\cpu.intr.r_clock_cmp[6] ),
    .A2(net412),
    .A1(_05737_));
 sg13g2_o21ai_1 _23343_ (.B1(_05738_),
    .Y(_05739_),
    .A1(net733),
    .A2(_05736_));
 sg13g2_inv_1 _23344_ (.Y(_05740_),
    .A(_00145_));
 sg13g2_buf_1 _23345_ (.A(\cpu.spi.r_clk_count[2][6] ),
    .X(_05741_));
 sg13g2_a22oi_1 _23346_ (.Y(_05742_),
    .B1(_04964_),
    .B2(_05741_),
    .A2(net392),
    .A1(_05740_));
 sg13g2_nor2_1 _23347_ (.A(_00144_),
    .B(_04967_),
    .Y(_05743_));
 sg13g2_a21oi_1 _23348_ (.A1(\cpu.spi.r_timeout[6] ),
    .A2(_05082_),
    .Y(_05744_),
    .B1(_05743_));
 sg13g2_nand2_1 _23349_ (.Y(_05745_),
    .A(_09318_),
    .B(_04954_));
 sg13g2_nand3_1 _23350_ (.B(_05744_),
    .C(_05745_),
    .A(_05742_),
    .Y(_05746_));
 sg13g2_a22oi_1 _23351_ (.Y(_05747_),
    .B1(_05746_),
    .B2(_05077_),
    .A2(_05739_),
    .A1(_05110_));
 sg13g2_nand4_1 _23352_ (.B(_05729_),
    .C(_05731_),
    .A(net848),
    .Y(_05748_),
    .D(_05747_));
 sg13g2_o21ai_1 _23353_ (.B1(_05748_),
    .Y(_05749_),
    .A1(net848),
    .A2(_05711_));
 sg13g2_nand2_1 _23354_ (.Y(_05750_),
    .A(net1028),
    .B(net78));
 sg13g2_o21ai_1 _23355_ (.B1(_05750_),
    .Y(_05751_),
    .A1(net77),
    .A2(_05749_));
 sg13g2_nand2_1 _23356_ (.Y(_05752_),
    .A(net150),
    .B(_05751_));
 sg13g2_o21ai_1 _23357_ (.B1(_05752_),
    .Y(_01041_),
    .A1(net121),
    .A2(_05693_));
 sg13g2_nor2_1 _23358_ (.A(net581),
    .B(_04706_),
    .Y(_05753_));
 sg13g2_nor2_1 _23359_ (.A(net78),
    .B(_05158_),
    .Y(_05754_));
 sg13g2_a21oi_1 _23360_ (.A1(_10974_),
    .A2(_04885_),
    .Y(_05755_),
    .B1(_05754_));
 sg13g2_nand3b_1 _23361_ (.B(_11537_),
    .C(_04860_),
    .Y(_05756_),
    .A_N(net962));
 sg13g2_o21ai_1 _23362_ (.B1(_05756_),
    .Y(_05757_),
    .A1(net191),
    .A2(_05755_));
 sg13g2_a221oi_1 _23363_ (.B2(_05197_),
    .C1(_05757_),
    .B1(_05753_),
    .A1(_04703_),
    .Y(_01042_),
    .A2(_05074_));
 sg13g2_and2_1 _23364_ (.A(net508),
    .B(_04735_),
    .X(_05758_));
 sg13g2_a21oi_1 _23365_ (.A1(_05195_),
    .A2(_04733_),
    .Y(_05759_),
    .B1(_05758_));
 sg13g2_o21ai_1 _23366_ (.B1(_05334_),
    .Y(_05760_),
    .A1(\cpu.ex.pc[8] ),
    .A2(net196));
 sg13g2_buf_2 _23367_ (.A(\cpu.intr.r_clock_count[24] ),
    .X(_05761_));
 sg13g2_a22oi_1 _23368_ (.Y(_05762_),
    .B1(net499),
    .B2(\cpu.intr.r_clock_cmp[8] ),
    .A2(net373),
    .A1(_05761_));
 sg13g2_a22oi_1 _23369_ (.Y(_05763_),
    .B1(net361),
    .B2(\cpu.intr.r_timer_count[8] ),
    .A2(net335),
    .A1(\cpu.intr.r_timer_reload[8] ));
 sg13g2_or2_1 _23370_ (.X(_05764_),
    .B(_05763_),
    .A(net617));
 sg13g2_a22oi_1 _23371_ (.Y(_05765_),
    .B1(net435),
    .B2(_10175_),
    .A2(_05187_),
    .A1(\cpu.intr.r_clock_cmp[24] ));
 sg13g2_nand3_1 _23372_ (.B(_05764_),
    .C(_05765_),
    .A(_05762_),
    .Y(_05766_));
 sg13g2_a21o_1 _23373_ (.A2(_05052_),
    .A1(_10134_),
    .B1(_05059_),
    .X(_05767_));
 sg13g2_a22oi_1 _23374_ (.Y(_05768_),
    .B1(_05767_),
    .B2(net500),
    .A2(_05766_),
    .A1(_05176_));
 sg13g2_o21ai_1 _23375_ (.B1(_05256_),
    .Y(_05769_),
    .A1(net966),
    .A2(_05768_));
 sg13g2_mux2_1 _23376_ (.A0(_05769_),
    .A1(_09203_),
    .S(_04885_),
    .X(_05770_));
 sg13g2_nand2_1 _23377_ (.Y(_05771_),
    .A(net150),
    .B(_05770_));
 sg13g2_a22oi_1 _23378_ (.Y(_01043_),
    .B1(_05760_),
    .B2(_05771_),
    .A2(_05759_),
    .A1(_05197_));
 sg13g2_a21oi_1 _23379_ (.A1(_04859_),
    .A2(_04769_),
    .Y(_05772_),
    .B1(_05073_));
 sg13g2_o21ai_1 _23380_ (.B1(_05772_),
    .Y(_05773_),
    .A1(_04859_),
    .A2(_04768_));
 sg13g2_a21o_1 _23381_ (.A2(_05381_),
    .A1(_10134_),
    .B1(_05389_),
    .X(_05774_));
 sg13g2_buf_1 _23382_ (.A(\cpu.intr.r_clock_count[25] ),
    .X(_05775_));
 sg13g2_a22oi_1 _23383_ (.Y(_05776_),
    .B1(net499),
    .B2(\cpu.intr.r_clock_cmp[9] ),
    .A2(net373),
    .A1(_05775_));
 sg13g2_a22oi_1 _23384_ (.Y(_05777_),
    .B1(net361),
    .B2(\cpu.intr.r_timer_count[9] ),
    .A2(net335),
    .A1(\cpu.intr.r_timer_reload[9] ));
 sg13g2_or2_1 _23385_ (.X(_05778_),
    .B(_05777_),
    .A(net615));
 sg13g2_a22oi_1 _23386_ (.Y(_05779_),
    .B1(net435),
    .B2(_10183_),
    .A2(_05187_),
    .A1(\cpu.intr.r_clock_cmp[25] ));
 sg13g2_nand3_1 _23387_ (.B(_05778_),
    .C(_05779_),
    .A(_05776_),
    .Y(_05780_));
 sg13g2_a22oi_1 _23388_ (.Y(_05781_),
    .B1(_05780_),
    .B2(_05176_),
    .A2(_05774_),
    .A1(net500));
 sg13g2_o21ai_1 _23389_ (.B1(_05256_),
    .Y(_05782_),
    .A1(_03034_),
    .A2(_05781_));
 sg13g2_o21ai_1 _23390_ (.B1(_05782_),
    .Y(_05783_),
    .A1(_08786_),
    .A2(_05198_));
 sg13g2_nor2_1 _23391_ (.A(net83),
    .B(_05783_),
    .Y(_05784_));
 sg13g2_and2_1 _23392_ (.A(_02984_),
    .B(net83),
    .X(_05785_));
 sg13g2_a21o_1 _23393_ (.A2(_05784_),
    .A1(_05773_),
    .B1(_05785_),
    .X(_01044_));
 sg13g2_a21oi_1 _23394_ (.A1(_03531_),
    .A2(\cpu.dec.r_rd[0] ),
    .Y(_05786_),
    .B1(net197));
 sg13g2_nand2_1 _23395_ (.Y(_05787_),
    .A(net1018),
    .B(net150));
 sg13g2_o21ai_1 _23396_ (.B1(_05787_),
    .Y(_01045_),
    .A1(_05416_),
    .A2(_05786_));
 sg13g2_a21oi_1 _23397_ (.A1(_03531_),
    .A2(\cpu.dec.r_rd[1] ),
    .Y(_05788_),
    .B1(net197));
 sg13g2_nand2_1 _23398_ (.Y(_05789_),
    .A(net1019),
    .B(_05694_));
 sg13g2_o21ai_1 _23399_ (.B1(_05789_),
    .Y(_01046_),
    .A1(net121),
    .A2(_05788_));
 sg13g2_nor3_1 _23400_ (.A(\cpu.dec.r_store ),
    .B(_09294_),
    .C(net197),
    .Y(_05790_));
 sg13g2_nand3_1 _23401_ (.B(net151),
    .C(_05790_),
    .A(\cpu.dec.r_rd[2] ),
    .Y(_05791_));
 sg13g2_o21ai_1 _23402_ (.B1(_05791_),
    .Y(_01047_),
    .A1(_03576_),
    .A2(net153));
 sg13g2_nand3_1 _23403_ (.B(net151),
    .C(_05790_),
    .A(\cpu.dec.r_rd[3] ),
    .Y(_05792_));
 sg13g2_o21ai_1 _23404_ (.B1(_05792_),
    .Y(_01048_),
    .A1(_10226_),
    .A2(_05232_));
 sg13g2_mux2_1 _23405_ (.A0(\cpu.dec.r_swapsp ),
    .A1(\cpu.ex.r_wb_swapsp ),
    .S(net150),
    .X(_01049_));
 sg13g2_and2_1 _23406_ (.A(_10988_),
    .B(_11004_),
    .X(_05793_));
 sg13g2_nand2_1 _23407_ (.Y(_05794_),
    .A(net850),
    .B(net150));
 sg13g2_o21ai_1 _23408_ (.B1(_05794_),
    .Y(_01050_),
    .A1(_05793_),
    .A2(net121));
 sg13g2_a22oi_1 _23409_ (.Y(_05795_),
    .B1(net533),
    .B2(_10496_),
    .A2(_10253_),
    .A1(_03590_));
 sg13g2_a221oi_1 _23410_ (.B2(_11185_),
    .C1(net966),
    .B1(net533),
    .A1(net1104),
    .Y(_05796_),
    .A2(net534));
 sg13g2_a21oi_1 _23411_ (.A1(net834),
    .A2(_05795_),
    .Y(_05797_),
    .B1(_05796_));
 sg13g2_mux2_1 _23412_ (.A0(_10191_),
    .A1(_05797_),
    .S(net153),
    .X(_01051_));
 sg13g2_and2_1 _23413_ (.A(_10461_),
    .B(_10462_),
    .X(_05798_));
 sg13g2_a221oi_1 _23414_ (.B2(_10407_),
    .C1(net966),
    .B1(net533),
    .A1(net1107),
    .Y(_05799_),
    .A2(net534));
 sg13g2_a21oi_1 _23415_ (.A1(net834),
    .A2(_05798_),
    .Y(_05800_),
    .B1(_05799_));
 sg13g2_mux2_1 _23416_ (.A0(_10198_),
    .A1(_05800_),
    .S(net153),
    .X(_01052_));
 sg13g2_or3_1 _23417_ (.A(_11305_),
    .B(_11317_),
    .C(_11321_),
    .X(_05801_));
 sg13g2_nand2_1 _23418_ (.Y(_05802_),
    .A(net834),
    .B(_05801_));
 sg13g2_o21ai_1 _23419_ (.B1(_05802_),
    .Y(_05803_),
    .A1(net834),
    .A2(_10377_));
 sg13g2_mux2_1 _23420_ (.A0(_10203_),
    .A1(_05803_),
    .S(net153),
    .X(_01053_));
 sg13g2_nand3_1 _23421_ (.B(_11354_),
    .C(_11355_),
    .A(net966),
    .Y(_05804_));
 sg13g2_o21ai_1 _23422_ (.B1(_05804_),
    .Y(_05805_),
    .A1(net834),
    .A2(_10317_));
 sg13g2_nand2_1 _23423_ (.Y(_05806_),
    .A(_10205_),
    .B(_05694_));
 sg13g2_o21ai_1 _23424_ (.B1(_05806_),
    .Y(_01054_),
    .A1(net121),
    .A2(_05805_));
 sg13g2_nor2_2 _23425_ (.A(_11255_),
    .B(_11256_),
    .Y(_05807_));
 sg13g2_mux2_1 _23426_ (.A0(_05807_),
    .A1(_11466_),
    .S(_11527_),
    .X(_05808_));
 sg13g2_nand2_1 _23427_ (.Y(_05809_),
    .A(_10215_),
    .B(net152));
 sg13g2_o21ai_1 _23428_ (.B1(_05809_),
    .Y(_01055_),
    .A1(net150),
    .A2(_05808_));
 sg13g2_nor2_1 _23429_ (.A(net834),
    .B(_11438_),
    .Y(_05810_));
 sg13g2_a21oi_1 _23430_ (.A1(net834),
    .A2(_11284_),
    .Y(_05811_),
    .B1(_05810_));
 sg13g2_nand2_1 _23431_ (.Y(_05812_),
    .A(_10220_),
    .B(net152));
 sg13g2_o21ai_1 _23432_ (.B1(_05812_),
    .Y(_01056_),
    .A1(net150),
    .A2(_05811_));
 sg13g2_a21oi_1 _23433_ (.A1(_10537_),
    .A2(_10545_),
    .Y(_05813_),
    .B1(_10315_));
 sg13g2_a21o_1 _23434_ (.A2(_10253_),
    .A1(_10107_),
    .B1(_05813_),
    .X(_05814_));
 sg13g2_nand2_1 _23435_ (.Y(_05815_),
    .A(_05814_),
    .B(_05334_));
 sg13g2_o21ai_1 _23436_ (.B1(_05815_),
    .Y(_01057_),
    .A1(net762),
    .A2(net153));
 sg13g2_nand2_1 _23437_ (.Y(_05816_),
    .A(_02709_),
    .B(net152));
 sg13g2_o21ai_1 _23438_ (.B1(_05816_),
    .Y(_01058_),
    .A1(_05795_),
    .A2(net121));
 sg13g2_nand2_1 _23439_ (.Y(_05817_),
    .A(net974),
    .B(net152));
 sg13g2_o21ai_1 _23440_ (.B1(_05817_),
    .Y(_01059_),
    .A1(_05798_),
    .A2(net121));
 sg13g2_mux2_1 _23441_ (.A0(_10152_),
    .A1(_05801_),
    .S(net151),
    .X(_01060_));
 sg13g2_nand2_1 _23442_ (.Y(_05818_),
    .A(_11354_),
    .B(_11355_));
 sg13g2_mux2_1 _23443_ (.A0(_10158_),
    .A1(_05818_),
    .S(net151),
    .X(_01061_));
 sg13g2_nand2_1 _23444_ (.Y(_05819_),
    .A(net982),
    .B(net152));
 sg13g2_o21ai_1 _23445_ (.B1(_05819_),
    .Y(_01062_),
    .A1(_05807_),
    .A2(net121));
 sg13g2_mux2_1 _23446_ (.A0(_10105_),
    .A1(_11284_),
    .S(net151),
    .X(_01063_));
 sg13g2_nor3_1 _23447_ (.A(_03034_),
    .B(_11151_),
    .C(_11152_),
    .Y(_05820_));
 sg13g2_a21oi_1 _23448_ (.A1(_03035_),
    .A2(_05793_),
    .Y(_05821_),
    .B1(_05820_));
 sg13g2_mux2_1 _23449_ (.A0(_10181_),
    .A1(_05821_),
    .S(net151),
    .X(_01064_));
 sg13g2_nor2_1 _23450_ (.A(_11219_),
    .B(_11221_),
    .Y(_05822_));
 sg13g2_nor2_1 _23451_ (.A(net966),
    .B(_05822_),
    .Y(_05823_));
 sg13g2_a21oi_1 _23452_ (.A1(net834),
    .A2(_05814_),
    .Y(_05824_),
    .B1(_05823_));
 sg13g2_nand2_1 _23453_ (.Y(_05825_),
    .A(_10186_),
    .B(net152));
 sg13g2_o21ai_1 _23454_ (.B1(_05825_),
    .Y(_01065_),
    .A1(net150),
    .A2(_05824_));
 sg13g2_or3_1 _23455_ (.A(_11008_),
    .B(_10500_),
    .C(_10465_),
    .X(_05826_));
 sg13g2_buf_1 _23456_ (.A(_05826_),
    .X(_05827_));
 sg13g2_o21ai_1 _23457_ (.B1(_03384_),
    .Y(_05828_),
    .A1(_10520_),
    .A2(_05827_));
 sg13g2_buf_1 _23458_ (.A(_05828_),
    .X(_05829_));
 sg13g2_nor4_2 _23459_ (.A(_08476_),
    .B(_04805_),
    .C(_10228_),
    .Y(_05830_),
    .D(_03610_));
 sg13g2_and2_1 _23460_ (.A(_05829_),
    .B(_05830_),
    .X(_05831_));
 sg13g2_buf_1 _23461_ (.A(_05831_),
    .X(_05832_));
 sg13g2_o21ai_1 _23462_ (.B1(_09877_),
    .Y(_05833_),
    .A1(net294),
    .A2(_05832_));
 sg13g2_buf_1 _23463_ (.A(_05833_),
    .X(_05834_));
 sg13g2_buf_1 _23464_ (.A(_00286_),
    .X(_05835_));
 sg13g2_nand2b_1 _23465_ (.Y(_05836_),
    .B(net965),
    .A_N(_05835_));
 sg13g2_o21ai_1 _23466_ (.B1(_05836_),
    .Y(_05837_),
    .A1(net965),
    .A2(net620));
 sg13g2_nand2_1 _23467_ (.Y(_05838_),
    .A(_05832_),
    .B(_05837_));
 sg13g2_mux2_1 _23468_ (.A0(net620),
    .A1(_08618_),
    .S(_08574_),
    .X(_05839_));
 sg13g2_mux2_1 _23469_ (.A0(_05838_),
    .A1(_05839_),
    .S(net294),
    .X(_05840_));
 sg13g2_nor2_1 _23470_ (.A(net618),
    .B(_05840_),
    .Y(_05841_));
 sg13g2_a21oi_1 _23471_ (.A1(_10844_),
    .A2(_05834_),
    .Y(_01068_),
    .B1(_05841_));
 sg13g2_buf_1 _23472_ (.A(_10304_),
    .X(_05842_));
 sg13g2_inv_2 _23473_ (.Y(_05843_),
    .A(net958));
 sg13g2_nor2_1 _23474_ (.A(net1108),
    .B(_05843_),
    .Y(_05844_));
 sg13g2_buf_2 _23475_ (.A(_05844_),
    .X(_05845_));
 sg13g2_nand2_1 _23476_ (.Y(_05846_),
    .A(net1108),
    .B(_05843_));
 sg13g2_buf_2 _23477_ (.A(_05846_),
    .X(_05847_));
 sg13g2_nand3b_1 _23478_ (.B(_05847_),
    .C(net965),
    .Y(_05848_),
    .A_N(_05845_));
 sg13g2_o21ai_1 _23479_ (.B1(_05848_),
    .Y(_05849_),
    .A1(net965),
    .A2(net614));
 sg13g2_nand2_1 _23480_ (.Y(_05850_),
    .A(_05832_),
    .B(_05849_));
 sg13g2_mux2_1 _23481_ (.A0(net614),
    .A1(_08666_),
    .S(_08574_),
    .X(_05851_));
 sg13g2_mux2_1 _23482_ (.A0(_05850_),
    .A1(_05851_),
    .S(net294),
    .X(_05852_));
 sg13g2_nor2_1 _23483_ (.A(net618),
    .B(_05852_),
    .Y(_05853_));
 sg13g2_a21oi_1 _23484_ (.A1(_05843_),
    .A2(_05834_),
    .Y(_01069_),
    .B1(_05853_));
 sg13g2_inv_2 _23485_ (.Y(_05854_),
    .A(net1103));
 sg13g2_nand2_1 _23486_ (.Y(_05855_),
    .A(net1108),
    .B(net958));
 sg13g2_buf_2 _23487_ (.A(_05855_),
    .X(_05856_));
 sg13g2_nor2_1 _23488_ (.A(net1103),
    .B(_05856_),
    .Y(_05857_));
 sg13g2_buf_1 _23489_ (.A(net1103),
    .X(_05858_));
 sg13g2_nand2_1 _23490_ (.Y(_05859_),
    .A(net957),
    .B(_05856_));
 sg13g2_nand3b_1 _23491_ (.B(_05859_),
    .C(net965),
    .Y(_05860_),
    .A_N(_05857_));
 sg13g2_o21ai_1 _23492_ (.B1(_05860_),
    .Y(_05861_),
    .A1(net965),
    .A2(net605));
 sg13g2_nand3_1 _23493_ (.B(_05832_),
    .C(_05861_),
    .A(net330),
    .Y(_05862_));
 sg13g2_nor2_1 _23494_ (.A(net605),
    .B(_08574_),
    .Y(_05863_));
 sg13g2_a21oi_1 _23495_ (.A1(_08871_),
    .A2(_08574_),
    .Y(_05864_),
    .B1(_05863_));
 sg13g2_or2_1 _23496_ (.X(_05865_),
    .B(_05864_),
    .A(net330));
 sg13g2_a21oi_1 _23497_ (.A1(_05862_),
    .A2(_05865_),
    .Y(_05866_),
    .B1(net618));
 sg13g2_a21oi_1 _23498_ (.A1(_05854_),
    .A2(_05834_),
    .Y(_01070_),
    .B1(_05866_));
 sg13g2_inv_1 _23499_ (.Y(_05867_),
    .A(_10947_));
 sg13g2_nand3_1 _23500_ (.B(net958),
    .C(net1103),
    .A(net1108),
    .Y(_05868_));
 sg13g2_buf_1 _23501_ (.A(_05868_),
    .X(_05869_));
 sg13g2_xnor2_1 _23502_ (.Y(_05870_),
    .A(net956),
    .B(_05869_));
 sg13g2_nand2_1 _23503_ (.Y(_05871_),
    .A(net965),
    .B(_05870_));
 sg13g2_o21ai_1 _23504_ (.B1(_05871_),
    .Y(_05872_),
    .A1(net965),
    .A2(net860));
 sg13g2_nand3_1 _23505_ (.B(_05832_),
    .C(_05872_),
    .A(net330),
    .Y(_05873_));
 sg13g2_nand2_1 _23506_ (.Y(_05874_),
    .A(_08551_),
    .B(_08558_));
 sg13g2_nor2_1 _23507_ (.A(net860),
    .B(_08574_),
    .Y(_05875_));
 sg13g2_o21ai_1 _23508_ (.B1(net294),
    .Y(_05876_),
    .A1(_05874_),
    .A2(_05875_));
 sg13g2_a21oi_1 _23509_ (.A1(_05873_),
    .A2(_05876_),
    .Y(_05877_),
    .B1(_09296_));
 sg13g2_a21oi_1 _23510_ (.A1(_05867_),
    .A2(_05834_),
    .Y(_01071_),
    .B1(_05877_));
 sg13g2_buf_1 _23511_ (.A(net595),
    .X(_05878_));
 sg13g2_buf_2 _23512_ (.A(_00188_),
    .X(_05879_));
 sg13g2_buf_1 _23513_ (.A(_10472_),
    .X(_05880_));
 sg13g2_buf_1 _23514_ (.A(_10947_),
    .X(_05881_));
 sg13g2_nor2_2 _23515_ (.A(net955),
    .B(net954),
    .Y(_05882_));
 sg13g2_nand2_1 _23516_ (.Y(_05883_),
    .A(_05879_),
    .B(_05882_));
 sg13g2_nand2_1 _23517_ (.Y(_05884_),
    .A(net1126),
    .B(_05830_));
 sg13g2_nor2_1 _23518_ (.A(_10444_),
    .B(_05884_),
    .Y(_05885_));
 sg13g2_nand3_1 _23519_ (.B(_05843_),
    .C(_05885_),
    .A(_10844_),
    .Y(_05886_));
 sg13g2_buf_1 _23520_ (.A(_05886_),
    .X(_05887_));
 sg13g2_nor2_1 _23521_ (.A(_05883_),
    .B(_05887_),
    .Y(_05888_));
 sg13g2_buf_1 _23522_ (.A(_05888_),
    .X(_05889_));
 sg13g2_buf_1 _23523_ (.A(_05889_),
    .X(_05890_));
 sg13g2_mux2_1 _23524_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(_05878_),
    .S(net277),
    .X(_01139_));
 sg13g2_mux2_1 _23525_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(net450),
    .S(net277),
    .X(_01140_));
 sg13g2_mux2_1 _23526_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(_03588_),
    .S(_05890_),
    .X(_01141_));
 sg13g2_mux2_1 _23527_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(net593),
    .S(net277),
    .X(_01142_));
 sg13g2_mux2_1 _23528_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(_03016_),
    .S(net277),
    .X(_01143_));
 sg13g2_mux2_1 _23529_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(net719),
    .S(net277),
    .X(_01144_));
 sg13g2_mux2_1 _23530_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(net718),
    .S(net277),
    .X(_01145_));
 sg13g2_mux2_1 _23531_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(_03019_),
    .S(net277),
    .X(_01146_));
 sg13g2_buf_1 _23532_ (.A(net968),
    .X(_05891_));
 sg13g2_mux2_1 _23533_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(net830),
    .S(net277),
    .X(_01147_));
 sg13g2_mux2_1 _23534_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(net831),
    .S(_05890_),
    .X(_01148_));
 sg13g2_mux2_1 _23535_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(net455),
    .S(_05889_),
    .X(_01149_));
 sg13g2_mux2_1 _23536_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(net454),
    .S(_05889_),
    .X(_01150_));
 sg13g2_buf_1 _23537_ (.A(_05885_),
    .X(_05892_));
 sg13g2_nand2_1 _23538_ (.Y(_05893_),
    .A(_05854_),
    .B(_05845_));
 sg13g2_buf_2 _23539_ (.A(_05893_),
    .X(_05894_));
 sg13g2_nand2_2 _23540_ (.Y(_05895_),
    .A(net864),
    .B(net954));
 sg13g2_nor2_2 _23541_ (.A(_05894_),
    .B(_05895_),
    .Y(_05896_));
 sg13g2_and2_1 _23542_ (.A(net434),
    .B(_05896_),
    .X(_05897_));
 sg13g2_buf_1 _23543_ (.A(_05897_),
    .X(_05898_));
 sg13g2_buf_1 _23544_ (.A(_05898_),
    .X(_05899_));
 sg13g2_mux2_1 _23545_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A1(net498),
    .S(net328),
    .X(_01151_));
 sg13g2_mux2_1 _23546_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A1(net450),
    .S(net328),
    .X(_01152_));
 sg13g2_mux2_1 _23547_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A1(_03588_),
    .S(net328),
    .X(_01153_));
 sg13g2_mux2_1 _23548_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A1(net593),
    .S(net328),
    .X(_01154_));
 sg13g2_buf_1 _23549_ (.A(net847),
    .X(_05900_));
 sg13g2_mux2_1 _23550_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A1(net716),
    .S(net328),
    .X(_01155_));
 sg13g2_mux2_1 _23551_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A1(net719),
    .S(net328),
    .X(_01156_));
 sg13g2_mux2_1 _23552_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A1(net718),
    .S(_05899_),
    .X(_01157_));
 sg13g2_buf_1 _23553_ (.A(_11085_),
    .X(_05901_));
 sg13g2_mux2_1 _23554_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A1(_05901_),
    .S(_05899_),
    .X(_01158_));
 sg13g2_mux2_1 _23555_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A1(net830),
    .S(net328),
    .X(_01159_));
 sg13g2_mux2_1 _23556_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A1(_04809_),
    .S(net328),
    .X(_01160_));
 sg13g2_mux2_1 _23557_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A1(net455),
    .S(_05898_),
    .X(_01161_));
 sg13g2_mux2_1 _23558_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A1(net454),
    .S(_05898_),
    .X(_01162_));
 sg13g2_buf_1 _23559_ (.A(net1108),
    .X(_05902_));
 sg13g2_nand2_1 _23560_ (.Y(_05903_),
    .A(net864),
    .B(_05902_));
 sg13g2_nand3_1 _23561_ (.B(_05854_),
    .C(_05881_),
    .A(_05842_),
    .Y(_05904_));
 sg13g2_nor2_1 _23562_ (.A(_05903_),
    .B(_05904_),
    .Y(_05905_));
 sg13g2_buf_2 _23563_ (.A(_05905_),
    .X(_05906_));
 sg13g2_and2_1 _23564_ (.A(net434),
    .B(_05906_),
    .X(_05907_));
 sg13g2_buf_1 _23565_ (.A(_05907_),
    .X(_05908_));
 sg13g2_buf_1 _23566_ (.A(_05908_),
    .X(_05909_));
 sg13g2_mux2_1 _23567_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .A1(net498),
    .S(net327),
    .X(_01163_));
 sg13g2_mux2_1 _23568_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .A1(net450),
    .S(net327),
    .X(_01164_));
 sg13g2_buf_1 _23569_ (.A(net860),
    .X(_05910_));
 sg13g2_mux2_1 _23570_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .A1(net715),
    .S(net327),
    .X(_01165_));
 sg13g2_mux2_1 _23571_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .A1(_03617_),
    .S(net327),
    .X(_01166_));
 sg13g2_mux2_1 _23572_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .A1(net716),
    .S(net327),
    .X(_01167_));
 sg13g2_mux2_1 _23573_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .A1(net719),
    .S(net327),
    .X(_01168_));
 sg13g2_mux2_1 _23574_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .A1(net718),
    .S(net327),
    .X(_01169_));
 sg13g2_mux2_1 _23575_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .A1(_05901_),
    .S(_05909_),
    .X(_01170_));
 sg13g2_mux2_1 _23576_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .A1(net830),
    .S(net327),
    .X(_01171_));
 sg13g2_mux2_1 _23577_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .A1(net831),
    .S(_05909_),
    .X(_01172_));
 sg13g2_mux2_1 _23578_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .A1(net455),
    .S(_05908_),
    .X(_01173_));
 sg13g2_mux2_1 _23579_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .A1(net454),
    .S(_05908_),
    .X(_01174_));
 sg13g2_nor2_2 _23580_ (.A(net955),
    .B(net956),
    .Y(_05911_));
 sg13g2_nand2b_1 _23581_ (.Y(_05912_),
    .B(_05911_),
    .A_N(_05879_));
 sg13g2_buf_1 _23582_ (.A(_05912_),
    .X(_05913_));
 sg13g2_nor2_1 _23583_ (.A(_05887_),
    .B(_05913_),
    .Y(_05914_));
 sg13g2_buf_1 _23584_ (.A(_05914_),
    .X(_05915_));
 sg13g2_buf_1 _23585_ (.A(_05915_),
    .X(_05916_));
 sg13g2_mux2_1 _23586_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(_05878_),
    .S(net276),
    .X(_01175_));
 sg13g2_mux2_1 _23587_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(net450),
    .S(net276),
    .X(_01176_));
 sg13g2_mux2_1 _23588_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(net715),
    .S(net276),
    .X(_01177_));
 sg13g2_mux2_1 _23589_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(_03617_),
    .S(net276),
    .X(_01178_));
 sg13g2_mux2_1 _23590_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(net716),
    .S(net276),
    .X(_01179_));
 sg13g2_mux2_1 _23591_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(_03618_),
    .S(net276),
    .X(_01180_));
 sg13g2_mux2_1 _23592_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(net718),
    .S(_05916_),
    .X(_01181_));
 sg13g2_mux2_1 _23593_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(net953),
    .S(net276),
    .X(_01182_));
 sg13g2_mux2_1 _23594_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(_05891_),
    .S(net276),
    .X(_01183_));
 sg13g2_mux2_1 _23595_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(net831),
    .S(_05916_),
    .X(_01184_));
 sg13g2_mux2_1 _23596_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(net455),
    .S(_05915_),
    .X(_01185_));
 sg13g2_mux2_1 _23597_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(net454),
    .S(_05915_),
    .X(_01186_));
 sg13g2_nand2b_1 _23598_ (.Y(_05917_),
    .B(_05885_),
    .A_N(_05847_));
 sg13g2_buf_2 _23599_ (.A(_05917_),
    .X(_05918_));
 sg13g2_nor2_1 _23600_ (.A(_05913_),
    .B(_05918_),
    .Y(_05919_));
 sg13g2_buf_1 _23601_ (.A(_05919_),
    .X(_05920_));
 sg13g2_buf_1 _23602_ (.A(_05920_),
    .X(_05921_));
 sg13g2_mux2_1 _23603_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A1(net498),
    .S(net275),
    .X(_01187_));
 sg13g2_mux2_1 _23604_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A1(net450),
    .S(net275),
    .X(_01188_));
 sg13g2_mux2_1 _23605_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A1(_05910_),
    .S(net275),
    .X(_01189_));
 sg13g2_buf_1 _23606_ (.A(_02990_),
    .X(_05922_));
 sg13g2_mux2_1 _23607_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A1(net580),
    .S(net275),
    .X(_01190_));
 sg13g2_mux2_1 _23608_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A1(net716),
    .S(net275),
    .X(_01191_));
 sg13g2_mux2_1 _23609_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A1(_03618_),
    .S(net275),
    .X(_01192_));
 sg13g2_mux2_1 _23610_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A1(net718),
    .S(_05921_),
    .X(_01193_));
 sg13g2_mux2_1 _23611_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A1(net953),
    .S(net275),
    .X(_01194_));
 sg13g2_mux2_1 _23612_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A1(_05891_),
    .S(net275),
    .X(_01195_));
 sg13g2_mux2_1 _23613_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A1(net831),
    .S(_05921_),
    .X(_01196_));
 sg13g2_mux2_1 _23614_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A1(net455),
    .S(_05920_),
    .X(_01197_));
 sg13g2_mux2_1 _23615_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A1(net454),
    .S(_05920_),
    .X(_01198_));
 sg13g2_nand2_1 _23616_ (.Y(_05923_),
    .A(_05845_),
    .B(net434));
 sg13g2_nor2_1 _23617_ (.A(_05913_),
    .B(_05923_),
    .Y(_05924_));
 sg13g2_buf_1 _23618_ (.A(_05924_),
    .X(_05925_));
 sg13g2_buf_1 _23619_ (.A(_05925_),
    .X(_05926_));
 sg13g2_mux2_1 _23620_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A1(net498),
    .S(net274),
    .X(_01199_));
 sg13g2_mux2_1 _23621_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A1(net450),
    .S(net274),
    .X(_01200_));
 sg13g2_mux2_1 _23622_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A1(_05910_),
    .S(net274),
    .X(_01201_));
 sg13g2_mux2_1 _23623_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A1(net580),
    .S(net274),
    .X(_01202_));
 sg13g2_mux2_1 _23624_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A1(_05900_),
    .S(net274),
    .X(_01203_));
 sg13g2_buf_1 _23625_ (.A(_09205_),
    .X(_05927_));
 sg13g2_mux2_1 _23626_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A1(_05927_),
    .S(net274),
    .X(_01204_));
 sg13g2_mux2_1 _23627_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A1(net718),
    .S(_05926_),
    .X(_01205_));
 sg13g2_mux2_1 _23628_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A1(net953),
    .S(net274),
    .X(_01206_));
 sg13g2_mux2_1 _23629_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A1(net830),
    .S(net274),
    .X(_01207_));
 sg13g2_mux2_1 _23630_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A1(net831),
    .S(_05926_),
    .X(_01208_));
 sg13g2_mux2_1 _23631_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A1(_03629_),
    .S(_05925_),
    .X(_01209_));
 sg13g2_mux2_1 _23632_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A1(_03630_),
    .S(_05925_),
    .X(_01210_));
 sg13g2_or2_1 _23633_ (.X(_05928_),
    .B(_05884_),
    .A(_10444_));
 sg13g2_buf_2 _23634_ (.A(_05928_),
    .X(_05929_));
 sg13g2_nor3_1 _23635_ (.A(_05856_),
    .B(_05929_),
    .C(_05913_),
    .Y(_05930_));
 sg13g2_buf_1 _23636_ (.A(_05930_),
    .X(_05931_));
 sg13g2_buf_1 _23637_ (.A(_05931_),
    .X(_05932_));
 sg13g2_mux2_1 _23638_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .A1(net498),
    .S(net326),
    .X(_01211_));
 sg13g2_mux2_1 _23639_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .A1(_04810_),
    .S(net326),
    .X(_01212_));
 sg13g2_mux2_1 _23640_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .A1(net715),
    .S(net326),
    .X(_01213_));
 sg13g2_mux2_1 _23641_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .A1(_05922_),
    .S(net326),
    .X(_01214_));
 sg13g2_mux2_1 _23642_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .A1(_05900_),
    .S(net326),
    .X(_01215_));
 sg13g2_mux2_1 _23643_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .A1(_05927_),
    .S(net326),
    .X(_01216_));
 sg13g2_mux2_1 _23644_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .A1(net718),
    .S(_05932_),
    .X(_01217_));
 sg13g2_mux2_1 _23645_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .A1(net953),
    .S(net326),
    .X(_01218_));
 sg13g2_mux2_1 _23646_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .A1(net830),
    .S(net326),
    .X(_01219_));
 sg13g2_mux2_1 _23647_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .A1(net831),
    .S(_05932_),
    .X(_01220_));
 sg13g2_mux2_1 _23648_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .A1(_03629_),
    .S(_05931_),
    .X(_01221_));
 sg13g2_mux2_1 _23649_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .A1(_03630_),
    .S(_05931_),
    .X(_01222_));
 sg13g2_nand2_2 _23650_ (.Y(_05933_),
    .A(net955),
    .B(net956));
 sg13g2_nor2_1 _23651_ (.A(net958),
    .B(net1103),
    .Y(_05934_));
 sg13g2_buf_1 _23652_ (.A(_05934_),
    .X(_05935_));
 sg13g2_nand2_1 _23653_ (.Y(_05936_),
    .A(_10844_),
    .B(_05935_));
 sg13g2_nor3_1 _23654_ (.A(_05929_),
    .B(_05933_),
    .C(_05936_),
    .Y(_05937_));
 sg13g2_buf_1 _23655_ (.A(_05937_),
    .X(_05938_));
 sg13g2_buf_1 _23656_ (.A(_05938_),
    .X(_05939_));
 sg13g2_mux2_1 _23657_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(net498),
    .S(net325),
    .X(_01223_));
 sg13g2_mux2_1 _23658_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(net450),
    .S(net325),
    .X(_01224_));
 sg13g2_mux2_1 _23659_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(net715),
    .S(net325),
    .X(_01225_));
 sg13g2_mux2_1 _23660_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(net580),
    .S(net325),
    .X(_01226_));
 sg13g2_mux2_1 _23661_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(net716),
    .S(net325),
    .X(_01227_));
 sg13g2_mux2_1 _23662_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(net829),
    .S(_05939_),
    .X(_01228_));
 sg13g2_mux2_1 _23663_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(net718),
    .S(net325),
    .X(_01229_));
 sg13g2_mux2_1 _23664_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(net953),
    .S(net325),
    .X(_01230_));
 sg13g2_mux2_1 _23665_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(net830),
    .S(net325),
    .X(_01231_));
 sg13g2_mux2_1 _23666_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(net831),
    .S(_05939_),
    .X(_01232_));
 sg13g2_buf_1 _23667_ (.A(_09461_),
    .X(_05940_));
 sg13g2_mux2_1 _23668_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(_05940_),
    .S(_05938_),
    .X(_01233_));
 sg13g2_buf_1 _23669_ (.A(_10238_),
    .X(_05941_));
 sg13g2_mux2_1 _23670_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(net496),
    .S(_05938_),
    .X(_01234_));
 sg13g2_nor4_1 _23671_ (.A(net864),
    .B(net957),
    .C(net954),
    .D(_05918_),
    .Y(_05942_));
 sg13g2_buf_1 _23672_ (.A(_05942_),
    .X(_05943_));
 sg13g2_buf_1 _23673_ (.A(_05943_),
    .X(_05944_));
 sg13g2_mux2_1 _23674_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A1(net498),
    .S(net273),
    .X(_01235_));
 sg13g2_mux2_1 _23675_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A1(net450),
    .S(net273),
    .X(_01236_));
 sg13g2_mux2_1 _23676_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A1(net715),
    .S(net273),
    .X(_01237_));
 sg13g2_mux2_1 _23677_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A1(net580),
    .S(net273),
    .X(_01238_));
 sg13g2_mux2_1 _23678_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A1(net716),
    .S(_05944_),
    .X(_01239_));
 sg13g2_mux2_1 _23679_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A1(net829),
    .S(net273),
    .X(_01240_));
 sg13g2_mux2_1 _23680_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A1(_04812_),
    .S(net273),
    .X(_01241_));
 sg13g2_mux2_1 _23681_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A1(net953),
    .S(net273),
    .X(_01242_));
 sg13g2_mux2_1 _23682_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A1(net830),
    .S(net273),
    .X(_01243_));
 sg13g2_mux2_1 _23683_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A1(net831),
    .S(_05944_),
    .X(_01244_));
 sg13g2_mux2_1 _23684_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A1(_05940_),
    .S(_05943_),
    .X(_01245_));
 sg13g2_mux2_1 _23685_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A1(net496),
    .S(_05943_),
    .X(_01246_));
 sg13g2_nor2_2 _23686_ (.A(_05894_),
    .B(_05933_),
    .Y(_05945_));
 sg13g2_and2_1 _23687_ (.A(_05892_),
    .B(_05945_),
    .X(_05946_));
 sg13g2_buf_1 _23688_ (.A(_05946_),
    .X(_05947_));
 sg13g2_buf_1 _23689_ (.A(_05947_),
    .X(_05948_));
 sg13g2_mux2_1 _23690_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A1(net498),
    .S(net324),
    .X(_01247_));
 sg13g2_buf_1 _23691_ (.A(_11895_),
    .X(_05949_));
 sg13g2_mux2_1 _23692_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A1(_05949_),
    .S(net324),
    .X(_01248_));
 sg13g2_mux2_1 _23693_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A1(net715),
    .S(net324),
    .X(_01249_));
 sg13g2_mux2_1 _23694_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A1(net580),
    .S(net324),
    .X(_01250_));
 sg13g2_mux2_1 _23695_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A1(net716),
    .S(_05948_),
    .X(_01251_));
 sg13g2_mux2_1 _23696_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A1(net829),
    .S(net324),
    .X(_01252_));
 sg13g2_buf_1 _23697_ (.A(_09203_),
    .X(_05950_));
 sg13g2_mux2_1 _23698_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A1(net828),
    .S(net324),
    .X(_01253_));
 sg13g2_mux2_1 _23699_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A1(net953),
    .S(net324),
    .X(_01254_));
 sg13g2_mux2_1 _23700_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A1(net830),
    .S(net324),
    .X(_01255_));
 sg13g2_buf_1 _23701_ (.A(net1107),
    .X(_05951_));
 sg13g2_mux2_1 _23702_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A1(_05951_),
    .S(_05948_),
    .X(_01256_));
 sg13g2_mux2_1 _23703_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A1(net497),
    .S(_05947_),
    .X(_01257_));
 sg13g2_mux2_1 _23704_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A1(_05941_),
    .S(_05947_),
    .X(_01258_));
 sg13g2_buf_1 _23705_ (.A(net595),
    .X(_05952_));
 sg13g2_nand2_1 _23706_ (.Y(_05953_),
    .A(_05880_),
    .B(_05902_));
 sg13g2_nor4_1 _23707_ (.A(_05843_),
    .B(net1103),
    .C(_05881_),
    .D(_05953_),
    .Y(_05954_));
 sg13g2_buf_2 _23708_ (.A(_05954_),
    .X(_05955_));
 sg13g2_and2_1 _23709_ (.A(net434),
    .B(_05955_),
    .X(_05956_));
 sg13g2_buf_1 _23710_ (.A(_05956_),
    .X(_05957_));
 sg13g2_buf_1 _23711_ (.A(_05957_),
    .X(_05958_));
 sg13g2_mux2_1 _23712_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .A1(_05952_),
    .S(net323),
    .X(_01259_));
 sg13g2_mux2_1 _23713_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .A1(_05949_),
    .S(net323),
    .X(_01260_));
 sg13g2_mux2_1 _23714_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .A1(net715),
    .S(net323),
    .X(_01261_));
 sg13g2_mux2_1 _23715_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .A1(net580),
    .S(net323),
    .X(_01262_));
 sg13g2_mux2_1 _23716_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .A1(net716),
    .S(_05958_),
    .X(_01263_));
 sg13g2_mux2_1 _23717_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .A1(net829),
    .S(net323),
    .X(_01264_));
 sg13g2_mux2_1 _23718_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .A1(_05950_),
    .S(net323),
    .X(_01265_));
 sg13g2_mux2_1 _23719_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .A1(net953),
    .S(net323),
    .X(_01266_));
 sg13g2_buf_1 _23720_ (.A(net1104),
    .X(_05959_));
 sg13g2_mux2_1 _23721_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .A1(net950),
    .S(net323),
    .X(_01267_));
 sg13g2_mux2_1 _23722_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .A1(_05951_),
    .S(_05958_),
    .X(_01268_));
 sg13g2_mux2_1 _23723_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .A1(net497),
    .S(_05957_),
    .X(_01269_));
 sg13g2_mux2_1 _23724_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .A1(_05941_),
    .S(_05957_),
    .X(_01270_));
 sg13g2_nor2_1 _23725_ (.A(_05883_),
    .B(_05918_),
    .Y(_05960_));
 sg13g2_buf_1 _23726_ (.A(_05960_),
    .X(_05961_));
 sg13g2_buf_1 _23727_ (.A(_05961_),
    .X(_05962_));
 sg13g2_mux2_1 _23728_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A1(_05952_),
    .S(net272),
    .X(_01271_));
 sg13g2_mux2_1 _23729_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A1(net495),
    .S(net272),
    .X(_01272_));
 sg13g2_mux2_1 _23730_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A1(net715),
    .S(_05962_),
    .X(_01273_));
 sg13g2_mux2_1 _23731_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A1(_05922_),
    .S(_05962_),
    .X(_01274_));
 sg13g2_buf_1 _23732_ (.A(_10057_),
    .X(_05963_));
 sg13g2_mux2_1 _23733_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A1(net827),
    .S(net272),
    .X(_01275_));
 sg13g2_mux2_1 _23734_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A1(net829),
    .S(net272),
    .X(_01276_));
 sg13g2_mux2_1 _23735_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A1(_05950_),
    .S(net272),
    .X(_01277_));
 sg13g2_buf_1 _23736_ (.A(_11085_),
    .X(_05964_));
 sg13g2_mux2_1 _23737_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A1(_05964_),
    .S(net272),
    .X(_01278_));
 sg13g2_mux2_1 _23738_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A1(net950),
    .S(net272),
    .X(_01279_));
 sg13g2_mux2_1 _23739_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A1(net951),
    .S(net272),
    .X(_01280_));
 sg13g2_mux2_1 _23740_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A1(net497),
    .S(_05961_),
    .X(_01281_));
 sg13g2_mux2_1 _23741_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A1(net496),
    .S(_05961_),
    .X(_01282_));
 sg13g2_or2_1 _23742_ (.X(_05965_),
    .B(_05933_),
    .A(_05879_));
 sg13g2_buf_1 _23743_ (.A(_05965_),
    .X(_05966_));
 sg13g2_nor2_1 _23744_ (.A(_05887_),
    .B(_05966_),
    .Y(_05967_));
 sg13g2_buf_1 _23745_ (.A(_05967_),
    .X(_05968_));
 sg13g2_buf_1 _23746_ (.A(_05968_),
    .X(_05969_));
 sg13g2_mux2_1 _23747_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(net494),
    .S(_05969_),
    .X(_01283_));
 sg13g2_mux2_1 _23748_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(net495),
    .S(net271),
    .X(_01284_));
 sg13g2_buf_1 _23749_ (.A(_11905_),
    .X(_05970_));
 sg13g2_mux2_1 _23750_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(net714),
    .S(net271),
    .X(_01285_));
 sg13g2_mux2_1 _23751_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(net580),
    .S(net271),
    .X(_01286_));
 sg13g2_mux2_1 _23752_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(net827),
    .S(net271),
    .X(_01287_));
 sg13g2_mux2_1 _23753_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(net829),
    .S(net271),
    .X(_01288_));
 sg13g2_mux2_1 _23754_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(net828),
    .S(net271),
    .X(_01289_));
 sg13g2_mux2_1 _23755_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(net949),
    .S(net271),
    .X(_01290_));
 sg13g2_mux2_1 _23756_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(net950),
    .S(net271),
    .X(_01291_));
 sg13g2_mux2_1 _23757_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(net951),
    .S(_05969_),
    .X(_01292_));
 sg13g2_mux2_1 _23758_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(net497),
    .S(_05968_),
    .X(_01293_));
 sg13g2_mux2_1 _23759_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(net496),
    .S(_05968_),
    .X(_01294_));
 sg13g2_nor2_1 _23760_ (.A(_05918_),
    .B(_05966_),
    .Y(_05971_));
 sg13g2_buf_1 _23761_ (.A(_05971_),
    .X(_05972_));
 sg13g2_buf_1 _23762_ (.A(_05972_),
    .X(_05973_));
 sg13g2_mux2_1 _23763_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A1(net494),
    .S(_05973_),
    .X(_01295_));
 sg13g2_mux2_1 _23764_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A1(net495),
    .S(net270),
    .X(_01296_));
 sg13g2_mux2_1 _23765_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A1(net714),
    .S(net270),
    .X(_01297_));
 sg13g2_mux2_1 _23766_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A1(net580),
    .S(net270),
    .X(_01298_));
 sg13g2_mux2_1 _23767_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A1(net827),
    .S(net270),
    .X(_01299_));
 sg13g2_mux2_1 _23768_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A1(net829),
    .S(net270),
    .X(_01300_));
 sg13g2_mux2_1 _23769_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A1(net828),
    .S(net270),
    .X(_01301_));
 sg13g2_mux2_1 _23770_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A1(net949),
    .S(net270),
    .X(_01302_));
 sg13g2_mux2_1 _23771_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A1(net950),
    .S(net270),
    .X(_01303_));
 sg13g2_mux2_1 _23772_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A1(net951),
    .S(_05973_),
    .X(_01304_));
 sg13g2_mux2_1 _23773_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A1(net497),
    .S(_05972_),
    .X(_01305_));
 sg13g2_mux2_1 _23774_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A1(net496),
    .S(_05972_),
    .X(_01306_));
 sg13g2_nor2_1 _23775_ (.A(_05923_),
    .B(_05966_),
    .Y(_05974_));
 sg13g2_buf_1 _23776_ (.A(_05974_),
    .X(_05975_));
 sg13g2_buf_1 _23777_ (.A(_05975_),
    .X(_05976_));
 sg13g2_mux2_1 _23778_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A1(net494),
    .S(_05976_),
    .X(_01307_));
 sg13g2_mux2_1 _23779_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A1(net495),
    .S(net269),
    .X(_01308_));
 sg13g2_mux2_1 _23780_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A1(net714),
    .S(net269),
    .X(_01309_));
 sg13g2_buf_1 _23781_ (.A(_02990_),
    .X(_05977_));
 sg13g2_mux2_1 _23782_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A1(net579),
    .S(net269),
    .X(_01310_));
 sg13g2_mux2_1 _23783_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A1(net827),
    .S(net269),
    .X(_01311_));
 sg13g2_mux2_1 _23784_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A1(net829),
    .S(net269),
    .X(_01312_));
 sg13g2_mux2_1 _23785_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A1(net828),
    .S(net269),
    .X(_01313_));
 sg13g2_mux2_1 _23786_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A1(net949),
    .S(net269),
    .X(_01314_));
 sg13g2_mux2_1 _23787_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A1(net950),
    .S(net269),
    .X(_01315_));
 sg13g2_mux2_1 _23788_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A1(net951),
    .S(_05976_),
    .X(_01316_));
 sg13g2_mux2_1 _23789_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A1(net497),
    .S(_05975_),
    .X(_01317_));
 sg13g2_mux2_1 _23790_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A1(net496),
    .S(_05975_),
    .X(_01318_));
 sg13g2_nor3_1 _23791_ (.A(_05856_),
    .B(_05929_),
    .C(_05966_),
    .Y(_05978_));
 sg13g2_buf_1 _23792_ (.A(_05978_),
    .X(_05979_));
 sg13g2_buf_1 _23793_ (.A(_05979_),
    .X(_05980_));
 sg13g2_mux2_1 _23794_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .A1(net494),
    .S(_05980_),
    .X(_01319_));
 sg13g2_mux2_1 _23795_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .A1(net495),
    .S(net322),
    .X(_01320_));
 sg13g2_mux2_1 _23796_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .A1(net714),
    .S(net322),
    .X(_01321_));
 sg13g2_mux2_1 _23797_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .A1(net579),
    .S(net322),
    .X(_01322_));
 sg13g2_mux2_1 _23798_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .A1(net827),
    .S(net322),
    .X(_01323_));
 sg13g2_buf_1 _23799_ (.A(_09205_),
    .X(_05981_));
 sg13g2_mux2_1 _23800_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .A1(_05981_),
    .S(net322),
    .X(_01324_));
 sg13g2_mux2_1 _23801_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .A1(net828),
    .S(net322),
    .X(_01325_));
 sg13g2_mux2_1 _23802_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .A1(net949),
    .S(net322),
    .X(_01326_));
 sg13g2_mux2_1 _23803_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .A1(net950),
    .S(net322),
    .X(_01327_));
 sg13g2_mux2_1 _23804_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .A1(net951),
    .S(_05980_),
    .X(_01328_));
 sg13g2_mux2_1 _23805_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .A1(net497),
    .S(_05979_),
    .X(_01329_));
 sg13g2_mux2_1 _23806_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .A1(net496),
    .S(_05979_),
    .X(_01330_));
 sg13g2_nand2_2 _23807_ (.Y(_05982_),
    .A(net955),
    .B(net954));
 sg13g2_nor3_1 _23808_ (.A(_05929_),
    .B(_05936_),
    .C(_05982_),
    .Y(_05983_));
 sg13g2_buf_1 _23809_ (.A(_05983_),
    .X(_05984_));
 sg13g2_buf_1 _23810_ (.A(_05984_),
    .X(_05985_));
 sg13g2_mux2_1 _23811_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(net494),
    .S(net321),
    .X(_01331_));
 sg13g2_mux2_1 _23812_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(net495),
    .S(net321),
    .X(_01332_));
 sg13g2_mux2_1 _23813_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(net714),
    .S(net321),
    .X(_01333_));
 sg13g2_mux2_1 _23814_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(net579),
    .S(net321),
    .X(_01334_));
 sg13g2_mux2_1 _23815_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(net827),
    .S(net321),
    .X(_01335_));
 sg13g2_mux2_1 _23816_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(net826),
    .S(net321),
    .X(_01336_));
 sg13g2_mux2_1 _23817_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(net828),
    .S(_05985_),
    .X(_01337_));
 sg13g2_mux2_1 _23818_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(net949),
    .S(net321),
    .X(_01338_));
 sg13g2_mux2_1 _23819_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(net950),
    .S(net321),
    .X(_01339_));
 sg13g2_mux2_1 _23820_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(net951),
    .S(_05985_),
    .X(_01340_));
 sg13g2_mux2_1 _23821_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(net497),
    .S(_05984_),
    .X(_01341_));
 sg13g2_mux2_1 _23822_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(net496),
    .S(_05984_),
    .X(_01342_));
 sg13g2_nor2_1 _23823_ (.A(net864),
    .B(net1103),
    .Y(_05986_));
 sg13g2_nand2_1 _23824_ (.Y(_05987_),
    .A(net954),
    .B(_05986_));
 sg13g2_nor2_1 _23825_ (.A(_05918_),
    .B(_05987_),
    .Y(_05988_));
 sg13g2_buf_2 _23826_ (.A(_05988_),
    .X(_05989_));
 sg13g2_buf_1 _23827_ (.A(_05989_),
    .X(_05990_));
 sg13g2_mux2_1 _23828_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A1(net494),
    .S(net268),
    .X(_01343_));
 sg13g2_mux2_1 _23829_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A1(net495),
    .S(net268),
    .X(_01344_));
 sg13g2_mux2_1 _23830_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A1(net714),
    .S(net268),
    .X(_01345_));
 sg13g2_mux2_1 _23831_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A1(net579),
    .S(net268),
    .X(_01346_));
 sg13g2_mux2_1 _23832_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A1(_05963_),
    .S(net268),
    .X(_01347_));
 sg13g2_mux2_1 _23833_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A1(net826),
    .S(net268),
    .X(_01348_));
 sg13g2_mux2_1 _23834_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A1(net828),
    .S(_05990_),
    .X(_01349_));
 sg13g2_mux2_1 _23835_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A1(net949),
    .S(net268),
    .X(_01350_));
 sg13g2_mux2_1 _23836_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A1(net950),
    .S(net268),
    .X(_01351_));
 sg13g2_mux2_1 _23837_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A1(net951),
    .S(_05990_),
    .X(_01352_));
 sg13g2_buf_1 _23838_ (.A(net620),
    .X(_05991_));
 sg13g2_mux2_1 _23839_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A1(net493),
    .S(_05989_),
    .X(_01353_));
 sg13g2_buf_1 _23840_ (.A(_10238_),
    .X(_05992_));
 sg13g2_mux2_1 _23841_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A1(net492),
    .S(_05989_),
    .X(_01354_));
 sg13g2_nor2_1 _23842_ (.A(_05894_),
    .B(_05982_),
    .Y(_05993_));
 sg13g2_and2_1 _23843_ (.A(_05892_),
    .B(_05993_),
    .X(_05994_));
 sg13g2_buf_1 _23844_ (.A(_05994_),
    .X(_05995_));
 sg13g2_buf_1 _23845_ (.A(_05995_),
    .X(_05996_));
 sg13g2_mux2_1 _23846_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A1(net494),
    .S(net320),
    .X(_01355_));
 sg13g2_mux2_1 _23847_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A1(net495),
    .S(net320),
    .X(_01356_));
 sg13g2_mux2_1 _23848_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A1(_05970_),
    .S(net320),
    .X(_01357_));
 sg13g2_mux2_1 _23849_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A1(net579),
    .S(net320),
    .X(_01358_));
 sg13g2_mux2_1 _23850_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A1(net827),
    .S(net320),
    .X(_01359_));
 sg13g2_mux2_1 _23851_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A1(_05981_),
    .S(net320),
    .X(_01360_));
 sg13g2_mux2_1 _23852_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A1(net828),
    .S(_05996_),
    .X(_01361_));
 sg13g2_mux2_1 _23853_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A1(net949),
    .S(net320),
    .X(_01362_));
 sg13g2_mux2_1 _23854_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A1(_05959_),
    .S(net320),
    .X(_01363_));
 sg13g2_mux2_1 _23855_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A1(net951),
    .S(_05996_),
    .X(_01364_));
 sg13g2_mux2_1 _23856_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A1(net493),
    .S(_05995_),
    .X(_01365_));
 sg13g2_mux2_1 _23857_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A1(net492),
    .S(_05995_),
    .X(_01366_));
 sg13g2_nor2_2 _23858_ (.A(_05904_),
    .B(_05953_),
    .Y(_05997_));
 sg13g2_and2_1 _23859_ (.A(net434),
    .B(_05997_),
    .X(_05998_));
 sg13g2_buf_1 _23860_ (.A(_05998_),
    .X(_05999_));
 sg13g2_buf_1 _23861_ (.A(_05999_),
    .X(_06000_));
 sg13g2_mux2_1 _23862_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .A1(net494),
    .S(net319),
    .X(_01367_));
 sg13g2_buf_1 _23863_ (.A(net605),
    .X(_06001_));
 sg13g2_mux2_1 _23864_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .A1(net491),
    .S(net319),
    .X(_01368_));
 sg13g2_mux2_1 _23865_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .A1(_05970_),
    .S(net319),
    .X(_01369_));
 sg13g2_mux2_1 _23866_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .A1(net579),
    .S(net319),
    .X(_01370_));
 sg13g2_mux2_1 _23867_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .A1(_05963_),
    .S(_06000_),
    .X(_01371_));
 sg13g2_mux2_1 _23868_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .A1(net826),
    .S(net319),
    .X(_01372_));
 sg13g2_buf_1 _23869_ (.A(net1043),
    .X(_06002_));
 sg13g2_mux2_1 _23870_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .A1(net825),
    .S(net319),
    .X(_01373_));
 sg13g2_mux2_1 _23871_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .A1(net949),
    .S(net319),
    .X(_01374_));
 sg13g2_mux2_1 _23872_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .A1(_05959_),
    .S(net319),
    .X(_01375_));
 sg13g2_buf_1 _23873_ (.A(_10386_),
    .X(_06003_));
 sg13g2_mux2_1 _23874_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .A1(net948),
    .S(_06000_),
    .X(_01376_));
 sg13g2_mux2_1 _23875_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .A1(net493),
    .S(_05999_),
    .X(_01377_));
 sg13g2_mux2_1 _23876_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .A1(net492),
    .S(_05999_),
    .X(_01378_));
 sg13g2_buf_1 _23877_ (.A(net595),
    .X(_06004_));
 sg13g2_or2_1 _23878_ (.X(_06005_),
    .B(_05982_),
    .A(_05879_));
 sg13g2_buf_1 _23879_ (.A(_06005_),
    .X(_06006_));
 sg13g2_nor2_1 _23880_ (.A(_05887_),
    .B(_06006_),
    .Y(_06007_));
 sg13g2_buf_1 _23881_ (.A(_06007_),
    .X(_06008_));
 sg13g2_buf_1 _23882_ (.A(_06008_),
    .X(_06009_));
 sg13g2_mux2_1 _23883_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(net490),
    .S(net267),
    .X(_01379_));
 sg13g2_mux2_1 _23884_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(net491),
    .S(net267),
    .X(_01380_));
 sg13g2_mux2_1 _23885_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(net714),
    .S(net267),
    .X(_01381_));
 sg13g2_mux2_1 _23886_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(net579),
    .S(net267),
    .X(_01382_));
 sg13g2_mux2_1 _23887_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(net827),
    .S(net267),
    .X(_01383_));
 sg13g2_mux2_1 _23888_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(net826),
    .S(_06009_),
    .X(_01384_));
 sg13g2_mux2_1 _23889_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(net825),
    .S(net267),
    .X(_01385_));
 sg13g2_mux2_1 _23890_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(_05964_),
    .S(_06009_),
    .X(_01386_));
 sg13g2_buf_1 _23891_ (.A(_10703_),
    .X(_06010_));
 sg13g2_mux2_1 _23892_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(net947),
    .S(net267),
    .X(_01387_));
 sg13g2_mux2_1 _23893_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(net948),
    .S(net267),
    .X(_01388_));
 sg13g2_mux2_1 _23894_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(net493),
    .S(_06008_),
    .X(_01389_));
 sg13g2_mux2_1 _23895_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(net492),
    .S(_06008_),
    .X(_01390_));
 sg13g2_nor2_1 _23896_ (.A(_05918_),
    .B(_06006_),
    .Y(_06011_));
 sg13g2_buf_1 _23897_ (.A(_06011_),
    .X(_06012_));
 sg13g2_buf_1 _23898_ (.A(_06012_),
    .X(_06013_));
 sg13g2_mux2_1 _23899_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A1(net490),
    .S(net266),
    .X(_01391_));
 sg13g2_mux2_1 _23900_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A1(net491),
    .S(net266),
    .X(_01392_));
 sg13g2_mux2_1 _23901_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A1(net714),
    .S(net266),
    .X(_01393_));
 sg13g2_mux2_1 _23902_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A1(net579),
    .S(net266),
    .X(_01394_));
 sg13g2_buf_1 _23903_ (.A(_10057_),
    .X(_06014_));
 sg13g2_mux2_1 _23904_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A1(net824),
    .S(net266),
    .X(_01395_));
 sg13g2_mux2_1 _23905_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A1(net826),
    .S(_06013_),
    .X(_01396_));
 sg13g2_mux2_1 _23906_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A1(net825),
    .S(net266),
    .X(_01397_));
 sg13g2_buf_1 _23907_ (.A(_11085_),
    .X(_06015_));
 sg13g2_mux2_1 _23908_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A1(net946),
    .S(_06013_),
    .X(_01398_));
 sg13g2_mux2_1 _23909_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A1(net947),
    .S(net266),
    .X(_01399_));
 sg13g2_mux2_1 _23910_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A1(net948),
    .S(net266),
    .X(_01400_));
 sg13g2_mux2_1 _23911_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A1(net493),
    .S(_06012_),
    .X(_01401_));
 sg13g2_mux2_1 _23912_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A1(net492),
    .S(_06012_),
    .X(_01402_));
 sg13g2_nor2_1 _23913_ (.A(_05883_),
    .B(_05923_),
    .Y(_06016_));
 sg13g2_buf_1 _23914_ (.A(_06016_),
    .X(_06017_));
 sg13g2_buf_1 _23915_ (.A(_06017_),
    .X(_06018_));
 sg13g2_mux2_1 _23916_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A1(net490),
    .S(net265),
    .X(_01403_));
 sg13g2_mux2_1 _23917_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A1(net491),
    .S(net265),
    .X(_01404_));
 sg13g2_buf_1 _23918_ (.A(net860),
    .X(_06019_));
 sg13g2_mux2_1 _23919_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A1(_06019_),
    .S(net265),
    .X(_01405_));
 sg13g2_mux2_1 _23920_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A1(_05977_),
    .S(net265),
    .X(_01406_));
 sg13g2_mux2_1 _23921_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A1(net824),
    .S(_06018_),
    .X(_01407_));
 sg13g2_mux2_1 _23922_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A1(net826),
    .S(net265),
    .X(_01408_));
 sg13g2_mux2_1 _23923_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A1(net825),
    .S(net265),
    .X(_01409_));
 sg13g2_mux2_1 _23924_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A1(net946),
    .S(_06018_),
    .X(_01410_));
 sg13g2_mux2_1 _23925_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A1(_06010_),
    .S(net265),
    .X(_01411_));
 sg13g2_mux2_1 _23926_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A1(net948),
    .S(net265),
    .X(_01412_));
 sg13g2_mux2_1 _23927_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A1(_05991_),
    .S(_06017_),
    .X(_01413_));
 sg13g2_mux2_1 _23928_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A1(_05992_),
    .S(_06017_),
    .X(_01414_));
 sg13g2_nor2_1 _23929_ (.A(_05923_),
    .B(_06006_),
    .Y(_06020_));
 sg13g2_buf_1 _23930_ (.A(_06020_),
    .X(_06021_));
 sg13g2_buf_1 _23931_ (.A(_06021_),
    .X(_06022_));
 sg13g2_mux2_1 _23932_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A1(net490),
    .S(net264),
    .X(_01415_));
 sg13g2_mux2_1 _23933_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A1(net491),
    .S(net264),
    .X(_01416_));
 sg13g2_mux2_1 _23934_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A1(net713),
    .S(net264),
    .X(_01417_));
 sg13g2_mux2_1 _23935_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A1(_05977_),
    .S(net264),
    .X(_01418_));
 sg13g2_mux2_1 _23936_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A1(net824),
    .S(net264),
    .X(_01419_));
 sg13g2_mux2_1 _23937_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A1(net826),
    .S(_06022_),
    .X(_01420_));
 sg13g2_mux2_1 _23938_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A1(net825),
    .S(net264),
    .X(_01421_));
 sg13g2_mux2_1 _23939_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A1(net946),
    .S(_06022_),
    .X(_01422_));
 sg13g2_mux2_1 _23940_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A1(net947),
    .S(net264),
    .X(_01423_));
 sg13g2_mux2_1 _23941_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A1(net948),
    .S(net264),
    .X(_01424_));
 sg13g2_mux2_1 _23942_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A1(_05991_),
    .S(_06021_),
    .X(_01425_));
 sg13g2_mux2_1 _23943_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A1(net492),
    .S(_06021_),
    .X(_01426_));
 sg13g2_nor3_1 _23944_ (.A(_05856_),
    .B(_05929_),
    .C(_06006_),
    .Y(_06023_));
 sg13g2_buf_1 _23945_ (.A(_06023_),
    .X(_06024_));
 sg13g2_buf_1 _23946_ (.A(_06024_),
    .X(_06025_));
 sg13g2_mux2_1 _23947_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .A1(net490),
    .S(net318),
    .X(_01427_));
 sg13g2_mux2_1 _23948_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .A1(net491),
    .S(net318),
    .X(_01428_));
 sg13g2_mux2_1 _23949_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .A1(net713),
    .S(net318),
    .X(_01429_));
 sg13g2_mux2_1 _23950_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .A1(net598),
    .S(net318),
    .X(_01430_));
 sg13g2_mux2_1 _23951_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .A1(net824),
    .S(net318),
    .X(_01431_));
 sg13g2_mux2_1 _23952_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .A1(net826),
    .S(_06025_),
    .X(_01432_));
 sg13g2_mux2_1 _23953_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .A1(net825),
    .S(net318),
    .X(_01433_));
 sg13g2_mux2_1 _23954_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .A1(net946),
    .S(_06025_),
    .X(_01434_));
 sg13g2_mux2_1 _23955_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .A1(net947),
    .S(net318),
    .X(_01435_));
 sg13g2_mux2_1 _23956_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .A1(net948),
    .S(net318),
    .X(_01436_));
 sg13g2_mux2_1 _23957_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .A1(net493),
    .S(_06024_),
    .X(_01437_));
 sg13g2_mux2_1 _23958_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .A1(net492),
    .S(_06024_),
    .X(_01438_));
 sg13g2_nor3_1 _23959_ (.A(_05856_),
    .B(_05883_),
    .C(_05929_),
    .Y(_06026_));
 sg13g2_buf_1 _23960_ (.A(_06026_),
    .X(_06027_));
 sg13g2_buf_1 _23961_ (.A(_06027_),
    .X(_06028_));
 sg13g2_mux2_1 _23962_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .A1(net490),
    .S(net317),
    .X(_01439_));
 sg13g2_mux2_1 _23963_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .A1(net491),
    .S(net317),
    .X(_01440_));
 sg13g2_mux2_1 _23964_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .A1(_06019_),
    .S(net317),
    .X(_01441_));
 sg13g2_mux2_1 _23965_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .A1(net598),
    .S(net317),
    .X(_01442_));
 sg13g2_mux2_1 _23966_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .A1(net824),
    .S(_06028_),
    .X(_01443_));
 sg13g2_mux2_1 _23967_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .A1(net841),
    .S(net317),
    .X(_01444_));
 sg13g2_mux2_1 _23968_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .A1(net825),
    .S(net317),
    .X(_01445_));
 sg13g2_mux2_1 _23969_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .A1(net946),
    .S(_06028_),
    .X(_01446_));
 sg13g2_mux2_1 _23970_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .A1(_06010_),
    .S(net317),
    .X(_01447_));
 sg13g2_mux2_1 _23971_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .A1(net948),
    .S(net317),
    .X(_01448_));
 sg13g2_mux2_1 _23972_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .A1(net493),
    .S(_06027_),
    .X(_01449_));
 sg13g2_mux2_1 _23973_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .A1(_05992_),
    .S(_06027_),
    .X(_01450_));
 sg13g2_nand2_1 _23974_ (.Y(_06029_),
    .A(net1103),
    .B(net956));
 sg13g2_nor3_1 _23975_ (.A(net955),
    .B(_05887_),
    .C(_06029_),
    .Y(_06030_));
 sg13g2_buf_1 _23976_ (.A(_06030_),
    .X(_06031_));
 sg13g2_buf_1 _23977_ (.A(_06031_),
    .X(_06032_));
 sg13g2_mux2_1 _23978_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(net490),
    .S(net263),
    .X(_01451_));
 sg13g2_mux2_1 _23979_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(net491),
    .S(net263),
    .X(_01452_));
 sg13g2_mux2_1 _23980_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(net713),
    .S(net263),
    .X(_01453_));
 sg13g2_mux2_1 _23981_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(net598),
    .S(_06032_),
    .X(_01454_));
 sg13g2_mux2_1 _23982_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(net824),
    .S(net263),
    .X(_01455_));
 sg13g2_mux2_1 _23983_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(net841),
    .S(net263),
    .X(_01456_));
 sg13g2_mux2_1 _23984_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(net825),
    .S(net263),
    .X(_01457_));
 sg13g2_mux2_1 _23985_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(net946),
    .S(net263),
    .X(_01458_));
 sg13g2_mux2_1 _23986_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(net947),
    .S(net263),
    .X(_01459_));
 sg13g2_mux2_1 _23987_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(net948),
    .S(_06032_),
    .X(_01460_));
 sg13g2_mux2_1 _23988_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(net493),
    .S(_06031_),
    .X(_01461_));
 sg13g2_mux2_1 _23989_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(net492),
    .S(_06031_),
    .X(_01462_));
 sg13g2_nor3_1 _23990_ (.A(_05842_),
    .B(_05903_),
    .C(_06029_),
    .Y(_06033_));
 sg13g2_buf_2 _23991_ (.A(_06033_),
    .X(_06034_));
 sg13g2_and2_1 _23992_ (.A(net434),
    .B(_06034_),
    .X(_06035_));
 sg13g2_buf_1 _23993_ (.A(_06035_),
    .X(_06036_));
 sg13g2_buf_1 _23994_ (.A(_06036_),
    .X(_06037_));
 sg13g2_mux2_1 _23995_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A1(net490),
    .S(net316),
    .X(_01463_));
 sg13g2_mux2_1 _23996_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A1(_06001_),
    .S(net316),
    .X(_01464_));
 sg13g2_mux2_1 _23997_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A1(net713),
    .S(net316),
    .X(_01465_));
 sg13g2_mux2_1 _23998_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A1(net598),
    .S(_06037_),
    .X(_01466_));
 sg13g2_mux2_1 _23999_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A1(net824),
    .S(net316),
    .X(_01467_));
 sg13g2_mux2_1 _24000_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A1(net841),
    .S(_06037_),
    .X(_01468_));
 sg13g2_mux2_1 _24001_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A1(_06002_),
    .S(net316),
    .X(_01469_));
 sg13g2_mux2_1 _24002_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A1(net946),
    .S(net316),
    .X(_01470_));
 sg13g2_mux2_1 _24003_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A1(net947),
    .S(net316),
    .X(_01471_));
 sg13g2_mux2_1 _24004_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A1(_06003_),
    .S(net316),
    .X(_01472_));
 sg13g2_mux2_1 _24005_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A1(net522),
    .S(_06036_),
    .X(_01473_));
 sg13g2_mux2_1 _24006_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A1(net521),
    .S(_06036_),
    .X(_01474_));
 sg13g2_nor2_1 _24007_ (.A(_05854_),
    .B(net954),
    .Y(_06038_));
 sg13g2_nand2_1 _24008_ (.Y(_06039_),
    .A(net958),
    .B(_06038_));
 sg13g2_nor3_2 _24009_ (.A(_05880_),
    .B(net952),
    .C(_06039_),
    .Y(_06040_));
 sg13g2_and2_1 _24010_ (.A(net434),
    .B(_06040_),
    .X(_06041_));
 sg13g2_buf_1 _24011_ (.A(_06041_),
    .X(_06042_));
 sg13g2_buf_1 _24012_ (.A(_06042_),
    .X(_06043_));
 sg13g2_mux2_1 _24013_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A1(_06004_),
    .S(net315),
    .X(_01475_));
 sg13g2_mux2_1 _24014_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A1(_06001_),
    .S(net315),
    .X(_01476_));
 sg13g2_mux2_1 _24015_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A1(net713),
    .S(net315),
    .X(_01477_));
 sg13g2_mux2_1 _24016_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A1(net598),
    .S(_06043_),
    .X(_01478_));
 sg13g2_mux2_1 _24017_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A1(_06014_),
    .S(net315),
    .X(_01479_));
 sg13g2_mux2_1 _24018_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A1(net841),
    .S(net315),
    .X(_01480_));
 sg13g2_mux2_1 _24019_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A1(_06002_),
    .S(net315),
    .X(_01481_));
 sg13g2_mux2_1 _24020_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A1(_06015_),
    .S(net315),
    .X(_01482_));
 sg13g2_mux2_1 _24021_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A1(net947),
    .S(net315),
    .X(_01483_));
 sg13g2_mux2_1 _24022_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A1(_06003_),
    .S(_06043_),
    .X(_01484_));
 sg13g2_mux2_1 _24023_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A1(net522),
    .S(_06042_),
    .X(_01485_));
 sg13g2_mux2_1 _24024_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A1(net521),
    .S(_06042_),
    .X(_01486_));
 sg13g2_nor2_1 _24025_ (.A(_05903_),
    .B(_06039_),
    .Y(_06044_));
 sg13g2_buf_2 _24026_ (.A(_06044_),
    .X(_06045_));
 sg13g2_and2_1 _24027_ (.A(net434),
    .B(_06045_),
    .X(_06046_));
 sg13g2_buf_1 _24028_ (.A(_06046_),
    .X(_06047_));
 sg13g2_buf_1 _24029_ (.A(_06047_),
    .X(_06048_));
 sg13g2_mux2_1 _24030_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .A1(_06004_),
    .S(net314),
    .X(_01487_));
 sg13g2_mux2_1 _24031_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .A1(net520),
    .S(net314),
    .X(_01488_));
 sg13g2_mux2_1 _24032_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .A1(net713),
    .S(net314),
    .X(_01489_));
 sg13g2_mux2_1 _24033_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .A1(net598),
    .S(_06048_),
    .X(_01490_));
 sg13g2_mux2_1 _24034_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .A1(_06014_),
    .S(net314),
    .X(_01491_));
 sg13g2_mux2_1 _24035_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .A1(net841),
    .S(net314),
    .X(_01492_));
 sg13g2_mux2_1 _24036_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .A1(net845),
    .S(net314),
    .X(_01493_));
 sg13g2_mux2_1 _24037_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .A1(net946),
    .S(net314),
    .X(_01494_));
 sg13g2_mux2_1 _24038_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .A1(net947),
    .S(net314),
    .X(_01495_));
 sg13g2_mux2_1 _24039_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .A1(net967),
    .S(_06048_),
    .X(_01496_));
 sg13g2_mux2_1 _24040_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .A1(net522),
    .S(_06047_),
    .X(_01497_));
 sg13g2_mux2_1 _24041_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .A1(net521),
    .S(_06047_),
    .X(_01498_));
 sg13g2_nor3_1 _24042_ (.A(_05929_),
    .B(_05895_),
    .C(_05936_),
    .Y(_06049_));
 sg13g2_buf_1 _24043_ (.A(_06049_),
    .X(_06050_));
 sg13g2_buf_1 _24044_ (.A(_06050_),
    .X(_06051_));
 sg13g2_mux2_1 _24045_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(_03593_),
    .S(net313),
    .X(_01499_));
 sg13g2_mux2_1 _24046_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(_03586_),
    .S(net313),
    .X(_01500_));
 sg13g2_mux2_1 _24047_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(net713),
    .S(net313),
    .X(_01501_));
 sg13g2_mux2_1 _24048_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(_02991_),
    .S(net313),
    .X(_01502_));
 sg13g2_mux2_1 _24049_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(net824),
    .S(_06051_),
    .X(_01503_));
 sg13g2_mux2_1 _24050_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(_02996_),
    .S(net313),
    .X(_01504_));
 sg13g2_mux2_1 _24051_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(net845),
    .S(_06051_),
    .X(_01505_));
 sg13g2_mux2_1 _24052_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(_06015_),
    .S(net313),
    .X(_01506_));
 sg13g2_mux2_1 _24053_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(net968),
    .S(net313),
    .X(_01507_));
 sg13g2_mux2_1 _24054_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(net967),
    .S(net313),
    .X(_01508_));
 sg13g2_mux2_1 _24055_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(_03582_),
    .S(_06050_),
    .X(_01509_));
 sg13g2_mux2_1 _24056_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(_03584_),
    .S(_06050_),
    .X(_01510_));
 sg13g2_nor3_1 _24057_ (.A(_05858_),
    .B(_05895_),
    .C(_05918_),
    .Y(_06052_));
 sg13g2_buf_1 _24058_ (.A(_06052_),
    .X(_06053_));
 sg13g2_buf_1 _24059_ (.A(_06053_),
    .X(_06054_));
 sg13g2_mux2_1 _24060_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A1(_03593_),
    .S(net262),
    .X(_01511_));
 sg13g2_mux2_1 _24061_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A1(_03586_),
    .S(net262),
    .X(_01512_));
 sg13g2_mux2_1 _24062_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A1(net713),
    .S(net262),
    .X(_01513_));
 sg13g2_mux2_1 _24063_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A1(_02991_),
    .S(_06054_),
    .X(_01514_));
 sg13g2_mux2_1 _24064_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A1(net847),
    .S(_06054_),
    .X(_01515_));
 sg13g2_mux2_1 _24065_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A1(_02996_),
    .S(net262),
    .X(_01516_));
 sg13g2_mux2_1 _24066_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A1(_02982_),
    .S(net262),
    .X(_01517_));
 sg13g2_mux2_1 _24067_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A1(net969),
    .S(net262),
    .X(_01518_));
 sg13g2_mux2_1 _24068_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A1(_02986_),
    .S(net262),
    .X(_01519_));
 sg13g2_mux2_1 _24069_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A1(_02988_),
    .S(net262),
    .X(_01520_));
 sg13g2_mux2_1 _24070_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A1(_03582_),
    .S(_06053_),
    .X(_01521_));
 sg13g2_mux2_1 _24071_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A1(_03584_),
    .S(_06053_),
    .X(_01522_));
 sg13g2_and2_1 _24072_ (.A(_05879_),
    .B(_05882_),
    .X(_06055_));
 sg13g2_buf_1 _24073_ (.A(_06055_),
    .X(_06056_));
 sg13g2_and3_1 _24074_ (.X(_06057_),
    .A(_08582_),
    .B(_10444_),
    .C(_05830_));
 sg13g2_buf_1 _24075_ (.A(_06057_),
    .X(_06058_));
 sg13g2_and3_1 _24076_ (.X(_06059_),
    .A(_10844_),
    .B(_05843_),
    .C(_06058_));
 sg13g2_buf_1 _24077_ (.A(_06059_),
    .X(_06060_));
 sg13g2_nand2_1 _24078_ (.Y(_06061_),
    .A(_06056_),
    .B(_06060_));
 sg13g2_buf_2 _24079_ (.A(_06061_),
    .X(_06062_));
 sg13g2_buf_1 _24080_ (.A(_06062_),
    .X(_06063_));
 sg13g2_nand2_1 _24081_ (.Y(_06064_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .B(_06062_));
 sg13g2_o21ai_1 _24082_ (.B1(_06064_),
    .Y(_01523_),
    .A1(net586),
    .A2(net261));
 sg13g2_mux2_1 _24083_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .S(net261),
    .X(_01524_));
 sg13g2_nand2_1 _24084_ (.Y(_06065_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .B(_06062_));
 sg13g2_o21ai_1 _24085_ (.B1(_06065_),
    .Y(_01525_),
    .A1(net587),
    .A2(net261));
 sg13g2_nand2_1 _24086_ (.Y(_06066_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .B(_06062_));
 sg13g2_o21ai_1 _24087_ (.B1(_06066_),
    .Y(_01526_),
    .A1(net652),
    .A2(_06063_));
 sg13g2_mux2_1 _24088_ (.A0(net729),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .S(net261),
    .X(_01527_));
 sg13g2_nand2_1 _24089_ (.Y(_06067_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .B(_06062_));
 sg13g2_o21ai_1 _24090_ (.B1(_06067_),
    .Y(_01528_),
    .A1(net728),
    .A2(_06063_));
 sg13g2_mux2_1 _24091_ (.A0(net727),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .S(net261),
    .X(_01529_));
 sg13g2_mux2_1 _24092_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .S(net261),
    .X(_01530_));
 sg13g2_mux2_1 _24093_ (.A0(net843),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .S(net261),
    .X(_01531_));
 sg13g2_mux2_1 _24094_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .S(net261),
    .X(_01532_));
 sg13g2_mux2_1 _24095_ (.A0(net453),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .S(_06062_),
    .X(_01533_));
 sg13g2_mux2_1 _24096_ (.A0(net452),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .S(_06062_),
    .X(_01534_));
 sg13g2_buf_1 _24097_ (.A(_06058_),
    .X(_06068_));
 sg13g2_nand2_1 _24098_ (.Y(_06069_),
    .A(_05896_),
    .B(_06068_));
 sg13g2_buf_2 _24099_ (.A(_06069_),
    .X(_06070_));
 sg13g2_buf_1 _24100_ (.A(_06070_),
    .X(_06071_));
 sg13g2_nand2_1 _24101_ (.Y(_06072_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .B(_06070_));
 sg13g2_o21ai_1 _24102_ (.B1(_06072_),
    .Y(_01535_),
    .A1(_03866_),
    .A2(net312));
 sg13g2_mux2_1 _24103_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .S(net312),
    .X(_01536_));
 sg13g2_nand2_1 _24104_ (.Y(_06073_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .B(_06070_));
 sg13g2_o21ai_1 _24105_ (.B1(_06073_),
    .Y(_01537_),
    .A1(net587),
    .A2(net312));
 sg13g2_nand2_1 _24106_ (.Y(_06074_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .B(_06070_));
 sg13g2_o21ai_1 _24107_ (.B1(_06074_),
    .Y(_01538_),
    .A1(net652),
    .A2(_06071_));
 sg13g2_mux2_1 _24108_ (.A0(net729),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .S(net312),
    .X(_01539_));
 sg13g2_nand2_1 _24109_ (.Y(_06075_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .B(_06070_));
 sg13g2_o21ai_1 _24110_ (.B1(_06075_),
    .Y(_01540_),
    .A1(net728),
    .A2(_06071_));
 sg13g2_mux2_1 _24111_ (.A0(net727),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .S(net312),
    .X(_01541_));
 sg13g2_mux2_1 _24112_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .S(net312),
    .X(_01542_));
 sg13g2_mux2_1 _24113_ (.A0(net843),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .S(net312),
    .X(_01543_));
 sg13g2_mux2_1 _24114_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .S(net312),
    .X(_01544_));
 sg13g2_mux2_1 _24115_ (.A0(net453),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .S(_06070_),
    .X(_01545_));
 sg13g2_mux2_1 _24116_ (.A0(_03859_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .S(_06070_),
    .X(_01546_));
 sg13g2_nand2_1 _24117_ (.Y(_06076_),
    .A(_05906_),
    .B(net433));
 sg13g2_buf_2 _24118_ (.A(_06076_),
    .X(_06077_));
 sg13g2_buf_1 _24119_ (.A(_06077_),
    .X(_06078_));
 sg13g2_nand2_1 _24120_ (.Y(_06079_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .B(_06077_));
 sg13g2_o21ai_1 _24121_ (.B1(_06079_),
    .Y(_01547_),
    .A1(net586),
    .A2(net311));
 sg13g2_mux2_1 _24122_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S(net311),
    .X(_01548_));
 sg13g2_nand2_1 _24123_ (.Y(_06080_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .B(_06077_));
 sg13g2_o21ai_1 _24124_ (.B1(_06080_),
    .Y(_01549_),
    .A1(net587),
    .A2(net311));
 sg13g2_nand2_1 _24125_ (.Y(_06081_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .B(_06077_));
 sg13g2_o21ai_1 _24126_ (.B1(_06081_),
    .Y(_01550_),
    .A1(net652),
    .A2(_06078_));
 sg13g2_mux2_1 _24127_ (.A0(net729),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S(net311),
    .X(_01551_));
 sg13g2_nand2_1 _24128_ (.Y(_06082_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .B(_06077_));
 sg13g2_o21ai_1 _24129_ (.B1(_06082_),
    .Y(_01552_),
    .A1(net728),
    .A2(_06078_));
 sg13g2_mux2_1 _24130_ (.A0(net727),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S(net311),
    .X(_01553_));
 sg13g2_mux2_1 _24131_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S(net311),
    .X(_01554_));
 sg13g2_mux2_1 _24132_ (.A0(net843),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S(net311),
    .X(_01555_));
 sg13g2_mux2_1 _24133_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S(net311),
    .X(_01556_));
 sg13g2_mux2_1 _24134_ (.A0(_03858_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S(_06077_),
    .X(_01557_));
 sg13g2_mux2_1 _24135_ (.A0(_03859_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S(_06077_),
    .X(_01558_));
 sg13g2_nor2_1 _24136_ (.A(_05879_),
    .B(_05895_),
    .Y(_06083_));
 sg13g2_nand2_1 _24137_ (.Y(_06084_),
    .A(_06083_),
    .B(_06060_));
 sg13g2_buf_2 _24138_ (.A(_06084_),
    .X(_06085_));
 sg13g2_buf_1 _24139_ (.A(_06085_),
    .X(_06086_));
 sg13g2_nand2_1 _24140_ (.Y(_06087_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .B(_06085_));
 sg13g2_o21ai_1 _24141_ (.B1(_06087_),
    .Y(_01559_),
    .A1(net586),
    .A2(net260));
 sg13g2_mux2_1 _24142_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .S(net260),
    .X(_01560_));
 sg13g2_nand2_1 _24143_ (.Y(_06088_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .B(_06085_));
 sg13g2_o21ai_1 _24144_ (.B1(_06088_),
    .Y(_01561_),
    .A1(net587),
    .A2(net260));
 sg13g2_nand2_1 _24145_ (.Y(_06089_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .B(_06085_));
 sg13g2_o21ai_1 _24146_ (.B1(_06089_),
    .Y(_01562_),
    .A1(net652),
    .A2(_06086_));
 sg13g2_mux2_1 _24147_ (.A0(net729),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .S(net260),
    .X(_01563_));
 sg13g2_nand2_1 _24148_ (.Y(_06090_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .B(_06085_));
 sg13g2_o21ai_1 _24149_ (.B1(_06090_),
    .Y(_01564_),
    .A1(net728),
    .A2(_06086_));
 sg13g2_mux2_1 _24150_ (.A0(net727),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .S(net260),
    .X(_01565_));
 sg13g2_mux2_1 _24151_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .S(net260),
    .X(_01566_));
 sg13g2_mux2_1 _24152_ (.A0(net843),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .S(net260),
    .X(_01567_));
 sg13g2_mux2_1 _24153_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .S(net260),
    .X(_01568_));
 sg13g2_mux2_1 _24154_ (.A0(net453),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .S(_06085_),
    .X(_01569_));
 sg13g2_mux2_1 _24155_ (.A0(net452),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .S(_06085_),
    .X(_01570_));
 sg13g2_nor2b_1 _24156_ (.A(_05847_),
    .B_N(net489),
    .Y(_06091_));
 sg13g2_buf_2 _24157_ (.A(_06091_),
    .X(_06092_));
 sg13g2_nand2_1 _24158_ (.Y(_06093_),
    .A(_06083_),
    .B(_06092_));
 sg13g2_buf_2 _24159_ (.A(_06093_),
    .X(_06094_));
 sg13g2_buf_1 _24160_ (.A(_06094_),
    .X(_06095_));
 sg13g2_nand2_1 _24161_ (.Y(_06096_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .B(_06094_));
 sg13g2_o21ai_1 _24162_ (.B1(_06096_),
    .Y(_01571_),
    .A1(net586),
    .A2(net259));
 sg13g2_mux2_1 _24163_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .S(net259),
    .X(_01572_));
 sg13g2_nand2_1 _24164_ (.Y(_06097_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .B(_06094_));
 sg13g2_o21ai_1 _24165_ (.B1(_06097_),
    .Y(_01573_),
    .A1(net587),
    .A2(net259));
 sg13g2_nand2_1 _24166_ (.Y(_06098_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .B(_06094_));
 sg13g2_o21ai_1 _24167_ (.B1(_06098_),
    .Y(_01574_),
    .A1(net652),
    .A2(_06095_));
 sg13g2_mux2_1 _24168_ (.A0(net729),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .S(net259),
    .X(_01575_));
 sg13g2_nand2_1 _24169_ (.Y(_06099_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .B(_06094_));
 sg13g2_o21ai_1 _24170_ (.B1(_06099_),
    .Y(_01576_),
    .A1(net728),
    .A2(_06095_));
 sg13g2_mux2_1 _24171_ (.A0(net727),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .S(net259),
    .X(_01577_));
 sg13g2_mux2_1 _24172_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .S(net259),
    .X(_01578_));
 sg13g2_mux2_1 _24173_ (.A0(net843),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .S(net259),
    .X(_01579_));
 sg13g2_mux2_1 _24174_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .S(net259),
    .X(_01580_));
 sg13g2_mux2_1 _24175_ (.A0(net453),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .S(_06094_),
    .X(_01581_));
 sg13g2_mux2_1 _24176_ (.A0(net452),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .S(_06094_),
    .X(_01582_));
 sg13g2_nand3_1 _24177_ (.B(_06083_),
    .C(net433),
    .A(_05845_),
    .Y(_06100_));
 sg13g2_buf_2 _24178_ (.A(_06100_),
    .X(_06101_));
 sg13g2_buf_1 _24179_ (.A(_06101_),
    .X(_06102_));
 sg13g2_nand2_1 _24180_ (.Y(_06103_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .B(_06101_));
 sg13g2_o21ai_1 _24181_ (.B1(_06103_),
    .Y(_01583_),
    .A1(net586),
    .A2(net310));
 sg13g2_mux2_1 _24182_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .S(net310),
    .X(_01584_));
 sg13g2_nand2_1 _24183_ (.Y(_06104_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .B(_06101_));
 sg13g2_o21ai_1 _24184_ (.B1(_06104_),
    .Y(_01585_),
    .A1(_03861_),
    .A2(net310));
 sg13g2_nand2_1 _24185_ (.Y(_06105_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .B(_06101_));
 sg13g2_o21ai_1 _24186_ (.B1(_06105_),
    .Y(_01586_),
    .A1(net652),
    .A2(_06102_));
 sg13g2_mux2_1 _24187_ (.A0(net729),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .S(net310),
    .X(_01587_));
 sg13g2_nand2_1 _24188_ (.Y(_06106_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .B(_06101_));
 sg13g2_o21ai_1 _24189_ (.B1(_06106_),
    .Y(_01588_),
    .A1(net728),
    .A2(_06102_));
 sg13g2_mux2_1 _24190_ (.A0(net727),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .S(net310),
    .X(_01589_));
 sg13g2_mux2_1 _24191_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .S(net310),
    .X(_01590_));
 sg13g2_mux2_1 _24192_ (.A0(net843),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .S(net310),
    .X(_01591_));
 sg13g2_mux2_1 _24193_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .S(net310),
    .X(_01592_));
 sg13g2_mux2_1 _24194_ (.A0(net453),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .S(_06101_),
    .X(_01593_));
 sg13g2_mux2_1 _24195_ (.A0(net452),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .S(_06101_),
    .X(_01594_));
 sg13g2_nor2b_1 _24196_ (.A(_05856_),
    .B_N(net489),
    .Y(_06107_));
 sg13g2_nand2_1 _24197_ (.Y(_06108_),
    .A(_06083_),
    .B(_06107_));
 sg13g2_buf_2 _24198_ (.A(_06108_),
    .X(_06109_));
 sg13g2_buf_1 _24199_ (.A(_06109_),
    .X(_06110_));
 sg13g2_nand2_1 _24200_ (.Y(_06111_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .B(_06109_));
 sg13g2_o21ai_1 _24201_ (.B1(_06111_),
    .Y(_01595_),
    .A1(_03866_),
    .A2(net309));
 sg13g2_mux2_1 _24202_ (.A0(_03860_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S(net309),
    .X(_01596_));
 sg13g2_nand2_1 _24203_ (.Y(_06112_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .B(_06109_));
 sg13g2_o21ai_1 _24204_ (.B1(_06112_),
    .Y(_01597_),
    .A1(_03861_),
    .A2(net309));
 sg13g2_nand2_1 _24205_ (.Y(_06113_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .B(_06109_));
 sg13g2_o21ai_1 _24206_ (.B1(_06113_),
    .Y(_01598_),
    .A1(net652),
    .A2(_06110_));
 sg13g2_mux2_1 _24207_ (.A0(net729),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S(net309),
    .X(_01599_));
 sg13g2_nand2_1 _24208_ (.Y(_06114_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .B(_06109_));
 sg13g2_o21ai_1 _24209_ (.B1(_06114_),
    .Y(_01600_),
    .A1(net728),
    .A2(_06110_));
 sg13g2_mux2_1 _24210_ (.A0(net727),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S(net309),
    .X(_01601_));
 sg13g2_mux2_1 _24211_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S(net309),
    .X(_01602_));
 sg13g2_mux2_1 _24212_ (.A0(net843),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S(net309),
    .X(_01603_));
 sg13g2_mux2_1 _24213_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S(net309),
    .X(_01604_));
 sg13g2_mux2_1 _24214_ (.A0(net453),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S(_06109_),
    .X(_01605_));
 sg13g2_mux2_1 _24215_ (.A0(net452),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S(_06109_),
    .X(_01606_));
 sg13g2_nor3_2 _24216_ (.A(net952),
    .B(net958),
    .C(net957),
    .Y(_06115_));
 sg13g2_nand4_1 _24217_ (.B(net956),
    .C(_06115_),
    .A(net955),
    .Y(_06116_),
    .D(net489));
 sg13g2_buf_2 _24218_ (.A(_06116_),
    .X(_06117_));
 sg13g2_buf_1 _24219_ (.A(_06117_),
    .X(_06118_));
 sg13g2_nand2_1 _24220_ (.Y(_06119_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .B(_06117_));
 sg13g2_o21ai_1 _24221_ (.B1(_06119_),
    .Y(_01607_),
    .A1(net586),
    .A2(net359));
 sg13g2_mux2_1 _24222_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .S(net359),
    .X(_01608_));
 sg13g2_nand2_1 _24223_ (.Y(_06120_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .B(_06117_));
 sg13g2_o21ai_1 _24224_ (.B1(_06120_),
    .Y(_01609_),
    .A1(net587),
    .A2(net359));
 sg13g2_buf_1 _24225_ (.A(net730),
    .X(_06121_));
 sg13g2_nand2_1 _24226_ (.Y(_06122_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .B(_06117_));
 sg13g2_o21ai_1 _24227_ (.B1(_06122_),
    .Y(_01610_),
    .A1(net647),
    .A2(_06118_));
 sg13g2_buf_1 _24228_ (.A(net847),
    .X(_06123_));
 sg13g2_mux2_1 _24229_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .S(_06118_),
    .X(_01611_));
 sg13g2_buf_1 _24230_ (.A(net846),
    .X(_06124_));
 sg13g2_nand2_1 _24231_ (.Y(_06125_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .B(_06117_));
 sg13g2_o21ai_1 _24232_ (.B1(_06125_),
    .Y(_01612_),
    .A1(net711),
    .A2(net359));
 sg13g2_buf_1 _24233_ (.A(net845),
    .X(_06126_));
 sg13g2_mux2_1 _24234_ (.A0(net710),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .S(net359),
    .X(_01613_));
 sg13g2_buf_1 _24235_ (.A(net969),
    .X(_06127_));
 sg13g2_mux2_1 _24236_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .S(net359),
    .X(_01614_));
 sg13g2_buf_1 _24237_ (.A(net968),
    .X(_06128_));
 sg13g2_mux2_1 _24238_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .S(net359),
    .X(_01615_));
 sg13g2_buf_1 _24239_ (.A(net967),
    .X(_06129_));
 sg13g2_mux2_1 _24240_ (.A0(net821),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .S(net359),
    .X(_01616_));
 sg13g2_mux2_1 _24241_ (.A0(net453),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .S(_06117_),
    .X(_01617_));
 sg13g2_mux2_1 _24242_ (.A0(net452),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .S(_06117_),
    .X(_01618_));
 sg13g2_nand3_1 _24243_ (.B(_05986_),
    .C(_06092_),
    .A(net956),
    .Y(_06130_));
 sg13g2_buf_2 _24244_ (.A(_06130_),
    .X(_06131_));
 sg13g2_buf_1 _24245_ (.A(_06131_),
    .X(_06132_));
 sg13g2_nand2_1 _24246_ (.Y(_06133_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .B(_06131_));
 sg13g2_o21ai_1 _24247_ (.B1(_06133_),
    .Y(_01619_),
    .A1(net586),
    .A2(net258));
 sg13g2_mux2_1 _24248_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .S(net258),
    .X(_01620_));
 sg13g2_nand2_1 _24249_ (.Y(_06134_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .B(_06131_));
 sg13g2_o21ai_1 _24250_ (.B1(_06134_),
    .Y(_01621_),
    .A1(net587),
    .A2(net258));
 sg13g2_nand2_1 _24251_ (.Y(_06135_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .B(_06131_));
 sg13g2_o21ai_1 _24252_ (.B1(_06135_),
    .Y(_01622_),
    .A1(net647),
    .A2(_06132_));
 sg13g2_mux2_1 _24253_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .S(_06132_),
    .X(_01623_));
 sg13g2_nand2_1 _24254_ (.Y(_06136_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .B(_06131_));
 sg13g2_o21ai_1 _24255_ (.B1(_06136_),
    .Y(_01624_),
    .A1(net711),
    .A2(net258));
 sg13g2_mux2_1 _24256_ (.A0(net710),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .S(net258),
    .X(_01625_));
 sg13g2_mux2_1 _24257_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .S(net258),
    .X(_01626_));
 sg13g2_mux2_1 _24258_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .S(net258),
    .X(_01627_));
 sg13g2_mux2_1 _24259_ (.A0(net821),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .S(net258),
    .X(_01628_));
 sg13g2_mux2_1 _24260_ (.A0(net453),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .S(_06131_),
    .X(_01629_));
 sg13g2_mux2_1 _24261_ (.A0(net452),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .S(_06131_),
    .X(_01630_));
 sg13g2_buf_1 _24262_ (.A(net650),
    .X(_06137_));
 sg13g2_nand2_1 _24263_ (.Y(_06138_),
    .A(_05945_),
    .B(net433));
 sg13g2_buf_2 _24264_ (.A(_06138_),
    .X(_06139_));
 sg13g2_buf_1 _24265_ (.A(_06139_),
    .X(_06140_));
 sg13g2_nand2_1 _24266_ (.Y(_06141_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .B(_06139_));
 sg13g2_o21ai_1 _24267_ (.B1(_06141_),
    .Y(_01631_),
    .A1(_06137_),
    .A2(net308));
 sg13g2_buf_1 _24268_ (.A(net520),
    .X(_06142_));
 sg13g2_mux2_1 _24269_ (.A0(net432),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .S(net308),
    .X(_01632_));
 sg13g2_buf_1 _24270_ (.A(net676),
    .X(_06143_));
 sg13g2_nand2_1 _24271_ (.Y(_06144_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .B(_06139_));
 sg13g2_o21ai_1 _24272_ (.B1(_06144_),
    .Y(_01633_),
    .A1(net577),
    .A2(net308));
 sg13g2_nand2_1 _24273_ (.Y(_06145_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .B(_06139_));
 sg13g2_o21ai_1 _24274_ (.B1(_06145_),
    .Y(_01634_),
    .A1(net647),
    .A2(_06140_));
 sg13g2_mux2_1 _24275_ (.A0(_06123_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .S(net308),
    .X(_01635_));
 sg13g2_nand2_1 _24276_ (.Y(_06146_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .B(_06139_));
 sg13g2_o21ai_1 _24277_ (.B1(_06146_),
    .Y(_01636_),
    .A1(_06124_),
    .A2(_06140_));
 sg13g2_mux2_1 _24278_ (.A0(_06126_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .S(net308),
    .X(_01637_));
 sg13g2_mux2_1 _24279_ (.A0(_06127_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .S(net308),
    .X(_01638_));
 sg13g2_mux2_1 _24280_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .S(net308),
    .X(_01639_));
 sg13g2_mux2_1 _24281_ (.A0(net821),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .S(net308),
    .X(_01640_));
 sg13g2_buf_1 _24282_ (.A(net522),
    .X(_06147_));
 sg13g2_mux2_1 _24283_ (.A0(_06147_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .S(_06139_),
    .X(_01641_));
 sg13g2_buf_1 _24284_ (.A(net521),
    .X(_06148_));
 sg13g2_mux2_1 _24285_ (.A0(_06148_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .S(_06139_),
    .X(_01642_));
 sg13g2_nand2_1 _24286_ (.Y(_06149_),
    .A(_05955_),
    .B(net433));
 sg13g2_buf_2 _24287_ (.A(_06149_),
    .X(_06150_));
 sg13g2_buf_1 _24288_ (.A(_06150_),
    .X(_06151_));
 sg13g2_nand2_1 _24289_ (.Y(_06152_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .B(_06150_));
 sg13g2_o21ai_1 _24290_ (.B1(_06152_),
    .Y(_01643_),
    .A1(net578),
    .A2(net307));
 sg13g2_mux2_1 _24291_ (.A0(_06142_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S(net307),
    .X(_01644_));
 sg13g2_nand2_1 _24292_ (.Y(_06153_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .B(_06150_));
 sg13g2_o21ai_1 _24293_ (.B1(_06153_),
    .Y(_01645_),
    .A1(net577),
    .A2(net307));
 sg13g2_nand2_1 _24294_ (.Y(_06154_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .B(_06150_));
 sg13g2_o21ai_1 _24295_ (.B1(_06154_),
    .Y(_01646_),
    .A1(net647),
    .A2(_06151_));
 sg13g2_mux2_1 _24296_ (.A0(_06123_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S(_06151_),
    .X(_01647_));
 sg13g2_nand2_1 _24297_ (.Y(_06155_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .B(_06150_));
 sg13g2_o21ai_1 _24298_ (.B1(_06155_),
    .Y(_01648_),
    .A1(_06124_),
    .A2(net307));
 sg13g2_mux2_1 _24299_ (.A0(_06126_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S(net307),
    .X(_01649_));
 sg13g2_mux2_1 _24300_ (.A0(_06127_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S(net307),
    .X(_01650_));
 sg13g2_mux2_1 _24301_ (.A0(_06128_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S(net307),
    .X(_01651_));
 sg13g2_mux2_1 _24302_ (.A0(_06129_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S(net307),
    .X(_01652_));
 sg13g2_mux2_1 _24303_ (.A0(net431),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S(_06150_),
    .X(_01653_));
 sg13g2_mux2_1 _24304_ (.A0(_06148_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S(_06150_),
    .X(_01654_));
 sg13g2_nand2_1 _24305_ (.Y(_06156_),
    .A(_06056_),
    .B(_06092_));
 sg13g2_buf_2 _24306_ (.A(_06156_),
    .X(_06157_));
 sg13g2_buf_1 _24307_ (.A(_06157_),
    .X(_06158_));
 sg13g2_nand2_1 _24308_ (.Y(_06159_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .B(_06157_));
 sg13g2_o21ai_1 _24309_ (.B1(_06159_),
    .Y(_01655_),
    .A1(_06137_),
    .A2(net257));
 sg13g2_mux2_1 _24310_ (.A0(net432),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .S(net257),
    .X(_01656_));
 sg13g2_nand2_1 _24311_ (.Y(_06160_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .B(_06157_));
 sg13g2_o21ai_1 _24312_ (.B1(_06160_),
    .Y(_01657_),
    .A1(net577),
    .A2(net257));
 sg13g2_nand2_1 _24313_ (.Y(_06161_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .B(_06157_));
 sg13g2_o21ai_1 _24314_ (.B1(_06161_),
    .Y(_01658_),
    .A1(net647),
    .A2(_06158_));
 sg13g2_mux2_1 _24315_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .S(net257),
    .X(_01659_));
 sg13g2_nand2_1 _24316_ (.Y(_06162_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .B(_06157_));
 sg13g2_o21ai_1 _24317_ (.B1(_06162_),
    .Y(_01660_),
    .A1(net711),
    .A2(_06158_));
 sg13g2_mux2_1 _24318_ (.A0(net710),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .S(net257),
    .X(_01661_));
 sg13g2_mux2_1 _24319_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .S(net257),
    .X(_01662_));
 sg13g2_mux2_1 _24320_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .S(net257),
    .X(_01663_));
 sg13g2_mux2_1 _24321_ (.A0(_06129_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .S(net257),
    .X(_01664_));
 sg13g2_mux2_1 _24322_ (.A0(_06147_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .S(_06157_),
    .X(_01665_));
 sg13g2_mux2_1 _24323_ (.A0(net430),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .S(_06157_),
    .X(_01666_));
 sg13g2_nor2_1 _24324_ (.A(_05879_),
    .B(_05933_),
    .Y(_06163_));
 sg13g2_nand2_1 _24325_ (.Y(_06164_),
    .A(_06163_),
    .B(_06060_));
 sg13g2_buf_2 _24326_ (.A(_06164_),
    .X(_06165_));
 sg13g2_buf_1 _24327_ (.A(_06165_),
    .X(_06166_));
 sg13g2_nand2_1 _24328_ (.Y(_06167_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .B(_06165_));
 sg13g2_o21ai_1 _24329_ (.B1(_06167_),
    .Y(_01667_),
    .A1(net578),
    .A2(net256));
 sg13g2_mux2_1 _24330_ (.A0(net432),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .S(net256),
    .X(_01668_));
 sg13g2_nand2_1 _24331_ (.Y(_06168_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .B(_06165_));
 sg13g2_o21ai_1 _24332_ (.B1(_06168_),
    .Y(_01669_),
    .A1(net577),
    .A2(net256));
 sg13g2_nand2_1 _24333_ (.Y(_06169_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .B(_06165_));
 sg13g2_o21ai_1 _24334_ (.B1(_06169_),
    .Y(_01670_),
    .A1(net647),
    .A2(net256));
 sg13g2_mux2_1 _24335_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .S(_06166_),
    .X(_01671_));
 sg13g2_nand2_1 _24336_ (.Y(_06170_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .B(_06165_));
 sg13g2_o21ai_1 _24337_ (.B1(_06170_),
    .Y(_01672_),
    .A1(net711),
    .A2(_06166_));
 sg13g2_mux2_1 _24338_ (.A0(net710),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .S(net256),
    .X(_01673_));
 sg13g2_mux2_1 _24339_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .S(net256),
    .X(_01674_));
 sg13g2_mux2_1 _24340_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .S(net256),
    .X(_01675_));
 sg13g2_mux2_1 _24341_ (.A0(net821),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .S(net256),
    .X(_01676_));
 sg13g2_mux2_1 _24342_ (.A0(net431),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .S(_06165_),
    .X(_01677_));
 sg13g2_mux2_1 _24343_ (.A0(net430),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .S(_06165_),
    .X(_01678_));
 sg13g2_nand2_1 _24344_ (.Y(_06171_),
    .A(_06163_),
    .B(_06092_));
 sg13g2_buf_2 _24345_ (.A(_06171_),
    .X(_06172_));
 sg13g2_buf_1 _24346_ (.A(_06172_),
    .X(_06173_));
 sg13g2_nand2_1 _24347_ (.Y(_06174_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .B(_06172_));
 sg13g2_o21ai_1 _24348_ (.B1(_06174_),
    .Y(_01679_),
    .A1(net578),
    .A2(net255));
 sg13g2_mux2_1 _24349_ (.A0(net432),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .S(net255),
    .X(_01680_));
 sg13g2_nand2_1 _24350_ (.Y(_06175_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .B(_06172_));
 sg13g2_o21ai_1 _24351_ (.B1(_06175_),
    .Y(_01681_),
    .A1(net577),
    .A2(net255));
 sg13g2_nand2_1 _24352_ (.Y(_06176_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .B(_06172_));
 sg13g2_o21ai_1 _24353_ (.B1(_06176_),
    .Y(_01682_),
    .A1(net647),
    .A2(net255));
 sg13g2_mux2_1 _24354_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .S(_06173_),
    .X(_01683_));
 sg13g2_nand2_1 _24355_ (.Y(_06177_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .B(_06172_));
 sg13g2_o21ai_1 _24356_ (.B1(_06177_),
    .Y(_01684_),
    .A1(net711),
    .A2(_06173_));
 sg13g2_mux2_1 _24357_ (.A0(net710),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .S(net255),
    .X(_01685_));
 sg13g2_mux2_1 _24358_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .S(net255),
    .X(_01686_));
 sg13g2_mux2_1 _24359_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .S(net255),
    .X(_01687_));
 sg13g2_mux2_1 _24360_ (.A0(net821),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .S(net255),
    .X(_01688_));
 sg13g2_mux2_1 _24361_ (.A0(net431),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .S(_06172_),
    .X(_01689_));
 sg13g2_mux2_1 _24362_ (.A0(net430),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .S(_06172_),
    .X(_01690_));
 sg13g2_nand3_1 _24363_ (.B(_06163_),
    .C(net489),
    .A(_05845_),
    .Y(_06178_));
 sg13g2_buf_2 _24364_ (.A(_06178_),
    .X(_06179_));
 sg13g2_buf_1 _24365_ (.A(_06179_),
    .X(_06180_));
 sg13g2_nand2_1 _24366_ (.Y(_06181_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .B(_06179_));
 sg13g2_o21ai_1 _24367_ (.B1(_06181_),
    .Y(_01691_),
    .A1(net578),
    .A2(net358));
 sg13g2_mux2_1 _24368_ (.A0(net432),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .S(net358),
    .X(_01692_));
 sg13g2_nand2_1 _24369_ (.Y(_06182_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .B(_06179_));
 sg13g2_o21ai_1 _24370_ (.B1(_06182_),
    .Y(_01693_),
    .A1(_06143_),
    .A2(net358));
 sg13g2_nand2_1 _24371_ (.Y(_06183_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .B(_06179_));
 sg13g2_o21ai_1 _24372_ (.B1(_06183_),
    .Y(_01694_),
    .A1(_06121_),
    .A2(net358));
 sg13g2_mux2_1 _24373_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .S(_06180_),
    .X(_01695_));
 sg13g2_nand2_1 _24374_ (.Y(_06184_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .B(_06179_));
 sg13g2_o21ai_1 _24375_ (.B1(_06184_),
    .Y(_01696_),
    .A1(net711),
    .A2(_06180_));
 sg13g2_mux2_1 _24376_ (.A0(net710),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .S(net358),
    .X(_01697_));
 sg13g2_mux2_1 _24377_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .S(net358),
    .X(_01698_));
 sg13g2_mux2_1 _24378_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .S(net358),
    .X(_01699_));
 sg13g2_mux2_1 _24379_ (.A0(net821),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .S(net358),
    .X(_01700_));
 sg13g2_mux2_1 _24380_ (.A0(net431),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .S(_06179_),
    .X(_01701_));
 sg13g2_mux2_1 _24381_ (.A0(net430),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .S(_06179_),
    .X(_01702_));
 sg13g2_nand2_1 _24382_ (.Y(_06185_),
    .A(_06163_),
    .B(_06107_));
 sg13g2_buf_2 _24383_ (.A(_06185_),
    .X(_06186_));
 sg13g2_buf_1 _24384_ (.A(_06186_),
    .X(_06187_));
 sg13g2_nand2_1 _24385_ (.Y(_06188_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .B(_06186_));
 sg13g2_o21ai_1 _24386_ (.B1(_06188_),
    .Y(_01703_),
    .A1(net578),
    .A2(net306));
 sg13g2_mux2_1 _24387_ (.A0(net432),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S(net306),
    .X(_01704_));
 sg13g2_nand2_1 _24388_ (.Y(_06189_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .B(_06186_));
 sg13g2_o21ai_1 _24389_ (.B1(_06189_),
    .Y(_01705_),
    .A1(_06143_),
    .A2(net306));
 sg13g2_nand2_1 _24390_ (.Y(_06190_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .B(_06186_));
 sg13g2_o21ai_1 _24391_ (.B1(_06190_),
    .Y(_01706_),
    .A1(_06121_),
    .A2(net306));
 sg13g2_mux2_1 _24392_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S(_06187_),
    .X(_01707_));
 sg13g2_nand2_1 _24393_ (.Y(_06191_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .B(_06186_));
 sg13g2_o21ai_1 _24394_ (.B1(_06191_),
    .Y(_01708_),
    .A1(net711),
    .A2(_06187_));
 sg13g2_mux2_1 _24395_ (.A0(net710),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S(net306),
    .X(_01709_));
 sg13g2_mux2_1 _24396_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S(net306),
    .X(_01710_));
 sg13g2_mux2_1 _24397_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S(net306),
    .X(_01711_));
 sg13g2_mux2_1 _24398_ (.A0(net821),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S(net306),
    .X(_01712_));
 sg13g2_mux2_1 _24399_ (.A0(net431),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S(_06186_),
    .X(_01713_));
 sg13g2_mux2_1 _24400_ (.A0(net430),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S(_06186_),
    .X(_01714_));
 sg13g2_inv_1 _24401_ (.Y(_06192_),
    .A(_05982_));
 sg13g2_nand3_1 _24402_ (.B(_06192_),
    .C(net489),
    .A(_06115_),
    .Y(_06193_));
 sg13g2_buf_2 _24403_ (.A(_06193_),
    .X(_06194_));
 sg13g2_buf_1 _24404_ (.A(_06194_),
    .X(_06195_));
 sg13g2_nand2_1 _24405_ (.Y(_06196_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .B(_06194_));
 sg13g2_o21ai_1 _24406_ (.B1(_06196_),
    .Y(_01715_),
    .A1(net578),
    .A2(net357));
 sg13g2_mux2_1 _24407_ (.A0(net432),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .S(net357),
    .X(_01716_));
 sg13g2_nand2_1 _24408_ (.Y(_06197_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .B(_06194_));
 sg13g2_o21ai_1 _24409_ (.B1(_06197_),
    .Y(_01717_),
    .A1(net577),
    .A2(net357));
 sg13g2_nand2_1 _24410_ (.Y(_06198_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .B(_06194_));
 sg13g2_o21ai_1 _24411_ (.B1(_06198_),
    .Y(_01718_),
    .A1(net647),
    .A2(net357));
 sg13g2_mux2_1 _24412_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .S(_06195_),
    .X(_01719_));
 sg13g2_nand2_1 _24413_ (.Y(_06199_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .B(_06194_));
 sg13g2_o21ai_1 _24414_ (.B1(_06199_),
    .Y(_01720_),
    .A1(net711),
    .A2(_06195_));
 sg13g2_mux2_1 _24415_ (.A0(net710),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .S(net357),
    .X(_01721_));
 sg13g2_mux2_1 _24416_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .S(net357),
    .X(_01722_));
 sg13g2_mux2_1 _24417_ (.A0(_06128_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .S(net357),
    .X(_01723_));
 sg13g2_mux2_1 _24418_ (.A0(net821),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .S(net357),
    .X(_01724_));
 sg13g2_mux2_1 _24419_ (.A0(net431),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .S(_06194_),
    .X(_01725_));
 sg13g2_mux2_1 _24420_ (.A0(net430),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .S(_06194_),
    .X(_01726_));
 sg13g2_nand2b_1 _24421_ (.Y(_06200_),
    .B(_06092_),
    .A_N(_05987_));
 sg13g2_buf_2 _24422_ (.A(_06200_),
    .X(_06201_));
 sg13g2_buf_1 _24423_ (.A(_06201_),
    .X(_06202_));
 sg13g2_nand2_1 _24424_ (.Y(_06203_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .B(_06201_));
 sg13g2_o21ai_1 _24425_ (.B1(_06203_),
    .Y(_01727_),
    .A1(net578),
    .A2(net254));
 sg13g2_mux2_1 _24426_ (.A0(net432),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .S(net254),
    .X(_01728_));
 sg13g2_nand2_1 _24427_ (.Y(_06204_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .B(_06201_));
 sg13g2_o21ai_1 _24428_ (.B1(_06204_),
    .Y(_01729_),
    .A1(net577),
    .A2(net254));
 sg13g2_buf_1 _24429_ (.A(net730),
    .X(_06205_));
 sg13g2_nand2_1 _24430_ (.Y(_06206_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .B(_06201_));
 sg13g2_o21ai_1 _24431_ (.B1(_06206_),
    .Y(_01730_),
    .A1(net646),
    .A2(net254));
 sg13g2_buf_1 _24432_ (.A(net847),
    .X(_06207_));
 sg13g2_mux2_1 _24433_ (.A0(net709),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .S(_06202_),
    .X(_01731_));
 sg13g2_buf_1 _24434_ (.A(net846),
    .X(_06208_));
 sg13g2_nand2_1 _24435_ (.Y(_06209_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .B(_06201_));
 sg13g2_o21ai_1 _24436_ (.B1(_06209_),
    .Y(_01732_),
    .A1(net708),
    .A2(_06202_));
 sg13g2_buf_1 _24437_ (.A(net845),
    .X(_06210_));
 sg13g2_mux2_1 _24438_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .S(net254),
    .X(_01733_));
 sg13g2_buf_1 _24439_ (.A(net969),
    .X(_06211_));
 sg13g2_mux2_1 _24440_ (.A0(net820),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .S(net254),
    .X(_01734_));
 sg13g2_buf_1 _24441_ (.A(net968),
    .X(_06212_));
 sg13g2_mux2_1 _24442_ (.A0(net819),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .S(net254),
    .X(_01735_));
 sg13g2_buf_1 _24443_ (.A(net967),
    .X(_06213_));
 sg13g2_mux2_1 _24444_ (.A0(net818),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .S(net254),
    .X(_01736_));
 sg13g2_mux2_1 _24445_ (.A0(net431),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .S(_06201_),
    .X(_01737_));
 sg13g2_mux2_1 _24446_ (.A0(net430),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .S(_06201_),
    .X(_01738_));
 sg13g2_nand2_1 _24447_ (.Y(_06214_),
    .A(_05993_),
    .B(net433));
 sg13g2_buf_2 _24448_ (.A(_06214_),
    .X(_06215_));
 sg13g2_buf_1 _24449_ (.A(_06215_),
    .X(_06216_));
 sg13g2_nand2_1 _24450_ (.Y(_06217_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .B(_06215_));
 sg13g2_o21ai_1 _24451_ (.B1(_06217_),
    .Y(_01739_),
    .A1(net578),
    .A2(net305));
 sg13g2_mux2_1 _24452_ (.A0(_06142_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .S(net305),
    .X(_01740_));
 sg13g2_nand2_1 _24453_ (.Y(_06218_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .B(_06215_));
 sg13g2_o21ai_1 _24454_ (.B1(_06218_),
    .Y(_01741_),
    .A1(net577),
    .A2(net305));
 sg13g2_nand2_1 _24455_ (.Y(_06219_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .B(_06215_));
 sg13g2_o21ai_1 _24456_ (.B1(_06219_),
    .Y(_01742_),
    .A1(net646),
    .A2(net305));
 sg13g2_mux2_1 _24457_ (.A0(net709),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .S(_06216_),
    .X(_01743_));
 sg13g2_nand2_1 _24458_ (.Y(_06220_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .B(_06215_));
 sg13g2_o21ai_1 _24459_ (.B1(_06220_),
    .Y(_01744_),
    .A1(net708),
    .A2(net305));
 sg13g2_mux2_1 _24460_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .S(net305),
    .X(_01745_));
 sg13g2_mux2_1 _24461_ (.A0(net820),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .S(net305),
    .X(_01746_));
 sg13g2_mux2_1 _24462_ (.A0(net819),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .S(net305),
    .X(_01747_));
 sg13g2_mux2_1 _24463_ (.A0(net818),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .S(_06216_),
    .X(_01748_));
 sg13g2_mux2_1 _24464_ (.A0(net431),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .S(_06215_),
    .X(_01749_));
 sg13g2_mux2_1 _24465_ (.A0(net430),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .S(_06215_),
    .X(_01750_));
 sg13g2_buf_1 _24466_ (.A(net650),
    .X(_06221_));
 sg13g2_nand2_1 _24467_ (.Y(_06222_),
    .A(_05997_),
    .B(net433));
 sg13g2_buf_2 _24468_ (.A(_06222_),
    .X(_06223_));
 sg13g2_buf_1 _24469_ (.A(_06223_),
    .X(_06224_));
 sg13g2_nand2_1 _24470_ (.Y(_06225_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .B(_06223_));
 sg13g2_o21ai_1 _24471_ (.B1(_06225_),
    .Y(_01751_),
    .A1(net576),
    .A2(net304));
 sg13g2_buf_1 _24472_ (.A(net520),
    .X(_06226_));
 sg13g2_mux2_1 _24473_ (.A0(net429),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S(net304),
    .X(_01752_));
 sg13g2_buf_1 _24474_ (.A(net676),
    .X(_06227_));
 sg13g2_nand2_1 _24475_ (.Y(_06228_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .B(_06223_));
 sg13g2_o21ai_1 _24476_ (.B1(_06228_),
    .Y(_01753_),
    .A1(_06227_),
    .A2(net304));
 sg13g2_nand2_1 _24477_ (.Y(_06229_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .B(_06223_));
 sg13g2_o21ai_1 _24478_ (.B1(_06229_),
    .Y(_01754_),
    .A1(net646),
    .A2(net304));
 sg13g2_mux2_1 _24479_ (.A0(net709),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S(_06224_),
    .X(_01755_));
 sg13g2_nand2_1 _24480_ (.Y(_06230_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .B(_06223_));
 sg13g2_o21ai_1 _24481_ (.B1(_06230_),
    .Y(_01756_),
    .A1(net708),
    .A2(_06224_));
 sg13g2_mux2_1 _24482_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S(net304),
    .X(_01757_));
 sg13g2_mux2_1 _24483_ (.A0(net820),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S(net304),
    .X(_01758_));
 sg13g2_mux2_1 _24484_ (.A0(net819),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S(net304),
    .X(_01759_));
 sg13g2_mux2_1 _24485_ (.A0(net818),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S(net304),
    .X(_01760_));
 sg13g2_buf_1 _24486_ (.A(net522),
    .X(_06231_));
 sg13g2_mux2_1 _24487_ (.A0(net428),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S(_06223_),
    .X(_01761_));
 sg13g2_buf_1 _24488_ (.A(net521),
    .X(_06232_));
 sg13g2_mux2_1 _24489_ (.A0(net427),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S(_06223_),
    .X(_01762_));
 sg13g2_nor2_1 _24490_ (.A(_05879_),
    .B(_05982_),
    .Y(_06233_));
 sg13g2_nand2_1 _24491_ (.Y(_06234_),
    .A(_06233_),
    .B(_06060_));
 sg13g2_buf_2 _24492_ (.A(_06234_),
    .X(_06235_));
 sg13g2_buf_1 _24493_ (.A(_06235_),
    .X(_06236_));
 sg13g2_nand2_1 _24494_ (.Y(_06237_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .B(_06235_));
 sg13g2_o21ai_1 _24495_ (.B1(_06237_),
    .Y(_01763_),
    .A1(net576),
    .A2(net253));
 sg13g2_mux2_1 _24496_ (.A0(net429),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .S(net253),
    .X(_01764_));
 sg13g2_nand2_1 _24497_ (.Y(_06238_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .B(_06235_));
 sg13g2_o21ai_1 _24498_ (.B1(_06238_),
    .Y(_01765_),
    .A1(net575),
    .A2(net253));
 sg13g2_nand2_1 _24499_ (.Y(_06239_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .B(_06235_));
 sg13g2_o21ai_1 _24500_ (.B1(_06239_),
    .Y(_01766_),
    .A1(net646),
    .A2(net253));
 sg13g2_mux2_1 _24501_ (.A0(net709),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .S(_06236_),
    .X(_01767_));
 sg13g2_nand2_1 _24502_ (.Y(_06240_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .B(_06235_));
 sg13g2_o21ai_1 _24503_ (.B1(_06240_),
    .Y(_01768_),
    .A1(net708),
    .A2(net253));
 sg13g2_mux2_1 _24504_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .S(net253),
    .X(_01769_));
 sg13g2_mux2_1 _24505_ (.A0(net820),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .S(net253),
    .X(_01770_));
 sg13g2_mux2_1 _24506_ (.A0(net819),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .S(net253),
    .X(_01771_));
 sg13g2_mux2_1 _24507_ (.A0(net818),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .S(_06236_),
    .X(_01772_));
 sg13g2_mux2_1 _24508_ (.A0(net428),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .S(_06235_),
    .X(_01773_));
 sg13g2_mux2_1 _24509_ (.A0(net427),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .S(_06235_),
    .X(_01774_));
 sg13g2_nand2_1 _24510_ (.Y(_06241_),
    .A(_06233_),
    .B(_06092_));
 sg13g2_buf_2 _24511_ (.A(_06241_),
    .X(_06242_));
 sg13g2_buf_1 _24512_ (.A(_06242_),
    .X(_06243_));
 sg13g2_nand2_1 _24513_ (.Y(_06244_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .B(_06242_));
 sg13g2_o21ai_1 _24514_ (.B1(_06244_),
    .Y(_01775_),
    .A1(net576),
    .A2(net252));
 sg13g2_mux2_1 _24515_ (.A0(net429),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .S(net252),
    .X(_01776_));
 sg13g2_nand2_1 _24516_ (.Y(_06245_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .B(_06242_));
 sg13g2_o21ai_1 _24517_ (.B1(_06245_),
    .Y(_01777_),
    .A1(net575),
    .A2(net252));
 sg13g2_nand2_1 _24518_ (.Y(_06246_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .B(_06242_));
 sg13g2_o21ai_1 _24519_ (.B1(_06246_),
    .Y(_01778_),
    .A1(net646),
    .A2(net252));
 sg13g2_mux2_1 _24520_ (.A0(net709),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .S(_06243_),
    .X(_01779_));
 sg13g2_nand2_1 _24521_ (.Y(_06247_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .B(_06242_));
 sg13g2_o21ai_1 _24522_ (.B1(_06247_),
    .Y(_01780_),
    .A1(net708),
    .A2(net252));
 sg13g2_mux2_1 _24523_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .S(net252),
    .X(_01781_));
 sg13g2_mux2_1 _24524_ (.A0(net820),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .S(net252),
    .X(_01782_));
 sg13g2_mux2_1 _24525_ (.A0(net819),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .S(net252),
    .X(_01783_));
 sg13g2_mux2_1 _24526_ (.A0(net818),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .S(_06243_),
    .X(_01784_));
 sg13g2_mux2_1 _24527_ (.A0(net428),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .S(_06242_),
    .X(_01785_));
 sg13g2_mux2_1 _24528_ (.A0(net427),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .S(_06242_),
    .X(_01786_));
 sg13g2_nand3_1 _24529_ (.B(_06056_),
    .C(net489),
    .A(_05845_),
    .Y(_06248_));
 sg13g2_buf_2 _24530_ (.A(_06248_),
    .X(_06249_));
 sg13g2_buf_1 _24531_ (.A(_06249_),
    .X(_06250_));
 sg13g2_nand2_1 _24532_ (.Y(_06251_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .B(_06249_));
 sg13g2_o21ai_1 _24533_ (.B1(_06251_),
    .Y(_01787_),
    .A1(net576),
    .A2(net356));
 sg13g2_mux2_1 _24534_ (.A0(net429),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .S(net356),
    .X(_01788_));
 sg13g2_nand2_1 _24535_ (.Y(_06252_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .B(_06249_));
 sg13g2_o21ai_1 _24536_ (.B1(_06252_),
    .Y(_01789_),
    .A1(_06227_),
    .A2(net356));
 sg13g2_nand2_1 _24537_ (.Y(_06253_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .B(_06249_));
 sg13g2_o21ai_1 _24538_ (.B1(_06253_),
    .Y(_01790_),
    .A1(net646),
    .A2(_06250_));
 sg13g2_mux2_1 _24539_ (.A0(net709),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .S(net356),
    .X(_01791_));
 sg13g2_nand2_1 _24540_ (.Y(_06254_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .B(_06249_));
 sg13g2_o21ai_1 _24541_ (.B1(_06254_),
    .Y(_01792_),
    .A1(_06208_),
    .A2(_06250_));
 sg13g2_mux2_1 _24542_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .S(net356),
    .X(_01793_));
 sg13g2_mux2_1 _24543_ (.A0(_06211_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .S(net356),
    .X(_01794_));
 sg13g2_mux2_1 _24544_ (.A0(net819),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .S(net356),
    .X(_01795_));
 sg13g2_mux2_1 _24545_ (.A0(net818),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .S(net356),
    .X(_01796_));
 sg13g2_mux2_1 _24546_ (.A0(net428),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .S(_06249_),
    .X(_01797_));
 sg13g2_mux2_1 _24547_ (.A0(net427),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .S(_06249_),
    .X(_01798_));
 sg13g2_nand3_1 _24548_ (.B(_06233_),
    .C(net489),
    .A(_05845_),
    .Y(_06255_));
 sg13g2_buf_2 _24549_ (.A(_06255_),
    .X(_06256_));
 sg13g2_buf_1 _24550_ (.A(_06256_),
    .X(_06257_));
 sg13g2_nand2_1 _24551_ (.Y(_06258_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .B(_06256_));
 sg13g2_o21ai_1 _24552_ (.B1(_06258_),
    .Y(_01799_),
    .A1(net576),
    .A2(net355));
 sg13g2_mux2_1 _24553_ (.A0(net429),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .S(net355),
    .X(_01800_));
 sg13g2_nand2_1 _24554_ (.Y(_06259_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .B(_06256_));
 sg13g2_o21ai_1 _24555_ (.B1(_06259_),
    .Y(_01801_),
    .A1(net575),
    .A2(net355));
 sg13g2_nand2_1 _24556_ (.Y(_06260_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .B(_06256_));
 sg13g2_o21ai_1 _24557_ (.B1(_06260_),
    .Y(_01802_),
    .A1(net646),
    .A2(net355));
 sg13g2_mux2_1 _24558_ (.A0(net709),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .S(_06257_),
    .X(_01803_));
 sg13g2_nand2_1 _24559_ (.Y(_06261_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .B(_06256_));
 sg13g2_o21ai_1 _24560_ (.B1(_06261_),
    .Y(_01804_),
    .A1(net708),
    .A2(net355));
 sg13g2_mux2_1 _24561_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .S(net355),
    .X(_01805_));
 sg13g2_mux2_1 _24562_ (.A0(net820),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .S(net355),
    .X(_01806_));
 sg13g2_mux2_1 _24563_ (.A0(net819),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .S(net355),
    .X(_01807_));
 sg13g2_mux2_1 _24564_ (.A0(net818),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .S(_06257_),
    .X(_01808_));
 sg13g2_mux2_1 _24565_ (.A0(net428),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .S(_06256_),
    .X(_01809_));
 sg13g2_mux2_1 _24566_ (.A0(net427),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .S(_06256_),
    .X(_01810_));
 sg13g2_nand2_1 _24567_ (.Y(_06262_),
    .A(_06233_),
    .B(_06107_));
 sg13g2_buf_2 _24568_ (.A(_06262_),
    .X(_06263_));
 sg13g2_buf_1 _24569_ (.A(_06263_),
    .X(_06264_));
 sg13g2_nand2_1 _24570_ (.Y(_06265_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .B(_06263_));
 sg13g2_o21ai_1 _24571_ (.B1(_06265_),
    .Y(_01811_),
    .A1(net576),
    .A2(net303));
 sg13g2_mux2_1 _24572_ (.A0(net429),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S(net303),
    .X(_01812_));
 sg13g2_nand2_1 _24573_ (.Y(_06266_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .B(_06263_));
 sg13g2_o21ai_1 _24574_ (.B1(_06266_),
    .Y(_01813_),
    .A1(net575),
    .A2(net303));
 sg13g2_nand2_1 _24575_ (.Y(_06267_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .B(_06263_));
 sg13g2_o21ai_1 _24576_ (.B1(_06267_),
    .Y(_01814_),
    .A1(net646),
    .A2(net303));
 sg13g2_mux2_1 _24577_ (.A0(net709),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S(_06264_),
    .X(_01815_));
 sg13g2_nand2_1 _24578_ (.Y(_06268_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .B(_06263_));
 sg13g2_o21ai_1 _24579_ (.B1(_06268_),
    .Y(_01816_),
    .A1(net708),
    .A2(net303));
 sg13g2_mux2_1 _24580_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S(net303),
    .X(_01817_));
 sg13g2_mux2_1 _24581_ (.A0(net820),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S(net303),
    .X(_01818_));
 sg13g2_mux2_1 _24582_ (.A0(net819),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S(net303),
    .X(_01819_));
 sg13g2_mux2_1 _24583_ (.A0(net818),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S(_06264_),
    .X(_01820_));
 sg13g2_mux2_1 _24584_ (.A0(net428),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S(_06263_),
    .X(_01821_));
 sg13g2_mux2_1 _24585_ (.A0(net427),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S(_06263_),
    .X(_01822_));
 sg13g2_nand2_1 _24586_ (.Y(_06269_),
    .A(_06056_),
    .B(_06107_));
 sg13g2_buf_2 _24587_ (.A(_06269_),
    .X(_06270_));
 sg13g2_buf_1 _24588_ (.A(_06270_),
    .X(_06271_));
 sg13g2_nand2_1 _24589_ (.Y(_06272_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .B(_06270_));
 sg13g2_o21ai_1 _24590_ (.B1(_06272_),
    .Y(_01823_),
    .A1(net576),
    .A2(net302));
 sg13g2_mux2_1 _24591_ (.A0(net429),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S(net302),
    .X(_01824_));
 sg13g2_nand2_1 _24592_ (.Y(_06273_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .B(_06270_));
 sg13g2_o21ai_1 _24593_ (.B1(_06273_),
    .Y(_01825_),
    .A1(net575),
    .A2(net302));
 sg13g2_nand2_1 _24594_ (.Y(_06274_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .B(_06270_));
 sg13g2_o21ai_1 _24595_ (.B1(_06274_),
    .Y(_01826_),
    .A1(_06205_),
    .A2(_06271_));
 sg13g2_mux2_1 _24596_ (.A0(_06207_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S(net302),
    .X(_01827_));
 sg13g2_nand2_1 _24597_ (.Y(_06275_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .B(_06270_));
 sg13g2_o21ai_1 _24598_ (.B1(_06275_),
    .Y(_01828_),
    .A1(_06208_),
    .A2(_06271_));
 sg13g2_mux2_1 _24599_ (.A0(_06210_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S(net302),
    .X(_01829_));
 sg13g2_mux2_1 _24600_ (.A0(_06211_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S(net302),
    .X(_01830_));
 sg13g2_mux2_1 _24601_ (.A0(_06212_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S(net302),
    .X(_01831_));
 sg13g2_mux2_1 _24602_ (.A0(_06213_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S(net302),
    .X(_01832_));
 sg13g2_mux2_1 _24603_ (.A0(net428),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S(_06270_),
    .X(_01833_));
 sg13g2_mux2_1 _24604_ (.A0(net427),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S(_06270_),
    .X(_01834_));
 sg13g2_nand3_1 _24605_ (.B(_06038_),
    .C(_06060_),
    .A(net864),
    .Y(_06276_));
 sg13g2_buf_2 _24606_ (.A(_06276_),
    .X(_06277_));
 sg13g2_buf_1 _24607_ (.A(_06277_),
    .X(_06278_));
 sg13g2_nand2_1 _24608_ (.Y(_06279_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .B(_06277_));
 sg13g2_o21ai_1 _24609_ (.B1(_06279_),
    .Y(_01835_),
    .A1(net576),
    .A2(net251));
 sg13g2_mux2_1 _24610_ (.A0(_06226_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .S(net251),
    .X(_01836_));
 sg13g2_nand2_1 _24611_ (.Y(_06280_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .B(_06277_));
 sg13g2_o21ai_1 _24612_ (.B1(_06280_),
    .Y(_01837_),
    .A1(net575),
    .A2(net251));
 sg13g2_nand2_1 _24613_ (.Y(_06281_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .B(_06277_));
 sg13g2_o21ai_1 _24614_ (.B1(_06281_),
    .Y(_01838_),
    .A1(_06205_),
    .A2(_06278_));
 sg13g2_mux2_1 _24615_ (.A0(_06207_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .S(_06278_),
    .X(_01839_));
 sg13g2_nand2_1 _24616_ (.Y(_06282_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .B(_06277_));
 sg13g2_o21ai_1 _24617_ (.B1(_06282_),
    .Y(_01840_),
    .A1(net708),
    .A2(net251));
 sg13g2_mux2_1 _24618_ (.A0(_06210_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .S(net251),
    .X(_01841_));
 sg13g2_mux2_1 _24619_ (.A0(net820),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .S(net251),
    .X(_01842_));
 sg13g2_mux2_1 _24620_ (.A0(_06212_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .S(net251),
    .X(_01843_));
 sg13g2_mux2_1 _24621_ (.A0(_06213_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .S(net251),
    .X(_01844_));
 sg13g2_mux2_1 _24622_ (.A0(net428),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .S(_06277_),
    .X(_01845_));
 sg13g2_mux2_1 _24623_ (.A0(net427),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .S(_06277_),
    .X(_01846_));
 sg13g2_nand2_1 _24624_ (.Y(_06283_),
    .A(_06034_),
    .B(_06068_));
 sg13g2_buf_2 _24625_ (.A(_06283_),
    .X(_06284_));
 sg13g2_buf_1 _24626_ (.A(_06284_),
    .X(_06285_));
 sg13g2_nand2_1 _24627_ (.Y(_06286_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .B(_06284_));
 sg13g2_o21ai_1 _24628_ (.B1(_06286_),
    .Y(_01847_),
    .A1(_06221_),
    .A2(net301));
 sg13g2_mux2_1 _24629_ (.A0(net429),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .S(net301),
    .X(_01848_));
 sg13g2_nand2_1 _24630_ (.Y(_06287_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .B(_06284_));
 sg13g2_o21ai_1 _24631_ (.B1(_06287_),
    .Y(_01849_),
    .A1(net575),
    .A2(net301));
 sg13g2_nand2_1 _24632_ (.Y(_06288_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .B(_06284_));
 sg13g2_o21ai_1 _24633_ (.B1(_06288_),
    .Y(_01850_),
    .A1(net730),
    .A2(_06285_));
 sg13g2_mux2_1 _24634_ (.A0(net726),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .S(net301),
    .X(_01851_));
 sg13g2_nand2_1 _24635_ (.Y(_06289_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .B(_06284_));
 sg13g2_o21ai_1 _24636_ (.B1(_06289_),
    .Y(_01852_),
    .A1(net846),
    .A2(_06285_));
 sg13g2_mux2_1 _24637_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .S(net301),
    .X(_01853_));
 sg13g2_mux2_1 _24638_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .S(net301),
    .X(_01854_));
 sg13g2_mux2_1 _24639_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .S(net301),
    .X(_01855_));
 sg13g2_mux2_1 _24640_ (.A0(net838),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .S(net301),
    .X(_01856_));
 sg13g2_mux2_1 _24641_ (.A0(_06231_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .S(_06284_),
    .X(_01857_));
 sg13g2_mux2_1 _24642_ (.A0(_06232_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .S(_06284_),
    .X(_01858_));
 sg13g2_nand2_1 _24643_ (.Y(_06290_),
    .A(_06040_),
    .B(net433));
 sg13g2_buf_2 _24644_ (.A(_06290_),
    .X(_06291_));
 sg13g2_buf_1 _24645_ (.A(_06291_),
    .X(_06292_));
 sg13g2_nand2_1 _24646_ (.Y(_06293_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .B(_06291_));
 sg13g2_o21ai_1 _24647_ (.B1(_06293_),
    .Y(_01859_),
    .A1(_06221_),
    .A2(net300));
 sg13g2_mux2_1 _24648_ (.A0(_06226_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .S(net300),
    .X(_01860_));
 sg13g2_nand2_1 _24649_ (.Y(_06294_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .B(_06291_));
 sg13g2_o21ai_1 _24650_ (.B1(_06294_),
    .Y(_01861_),
    .A1(net575),
    .A2(net300));
 sg13g2_nand2_1 _24651_ (.Y(_06295_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .B(_06291_));
 sg13g2_o21ai_1 _24652_ (.B1(_06295_),
    .Y(_01862_),
    .A1(net730),
    .A2(_06292_));
 sg13g2_mux2_1 _24653_ (.A0(net726),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .S(net300),
    .X(_01863_));
 sg13g2_nand2_1 _24654_ (.Y(_06296_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .B(_06291_));
 sg13g2_o21ai_1 _24655_ (.B1(_06296_),
    .Y(_01864_),
    .A1(net846),
    .A2(_06292_));
 sg13g2_mux2_1 _24656_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .S(net300),
    .X(_01865_));
 sg13g2_mux2_1 _24657_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .S(net300),
    .X(_01866_));
 sg13g2_mux2_1 _24658_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .S(net300),
    .X(_01867_));
 sg13g2_mux2_1 _24659_ (.A0(net838),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .S(net300),
    .X(_01868_));
 sg13g2_mux2_1 _24660_ (.A0(_06231_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .S(_06291_),
    .X(_01869_));
 sg13g2_mux2_1 _24661_ (.A0(_06232_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .S(_06291_),
    .X(_01870_));
 sg13g2_nand2_1 _24662_ (.Y(_06297_),
    .A(_06045_),
    .B(net433));
 sg13g2_buf_2 _24663_ (.A(_06297_),
    .X(_06298_));
 sg13g2_buf_1 _24664_ (.A(_06298_),
    .X(_06299_));
 sg13g2_nand2_1 _24665_ (.Y(_06300_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .B(_06298_));
 sg13g2_o21ai_1 _24666_ (.B1(_06300_),
    .Y(_01871_),
    .A1(net650),
    .A2(net299));
 sg13g2_mux2_1 _24667_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S(net299),
    .X(_01872_));
 sg13g2_nand2_1 _24668_ (.Y(_06301_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .B(_06298_));
 sg13g2_o21ai_1 _24669_ (.B1(_06301_),
    .Y(_01873_),
    .A1(net676),
    .A2(_06299_));
 sg13g2_nand2_1 _24670_ (.Y(_06302_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .B(_06298_));
 sg13g2_o21ai_1 _24671_ (.B1(_06302_),
    .Y(_01874_),
    .A1(net730),
    .A2(net299));
 sg13g2_mux2_1 _24672_ (.A0(net726),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S(net299),
    .X(_01875_));
 sg13g2_nand2_1 _24673_ (.Y(_06303_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .B(_06298_));
 sg13g2_o21ai_1 _24674_ (.B1(_06303_),
    .Y(_01876_),
    .A1(net846),
    .A2(_06299_));
 sg13g2_mux2_1 _24675_ (.A0(_02998_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S(net299),
    .X(_01877_));
 sg13g2_mux2_1 _24676_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S(net299),
    .X(_01878_));
 sg13g2_mux2_1 _24677_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S(net299),
    .X(_01879_));
 sg13g2_mux2_1 _24678_ (.A0(net838),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S(net299),
    .X(_01880_));
 sg13g2_mux2_1 _24679_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S(_06298_),
    .X(_01881_));
 sg13g2_mux2_1 _24680_ (.A0(_03585_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S(_06298_),
    .X(_01882_));
 sg13g2_nand3_1 _24681_ (.B(_06115_),
    .C(net489),
    .A(_05911_),
    .Y(_06304_));
 sg13g2_buf_2 _24682_ (.A(_06304_),
    .X(_06305_));
 sg13g2_buf_1 _24683_ (.A(_06305_),
    .X(_06306_));
 sg13g2_nand2_1 _24684_ (.Y(_06307_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .B(_06305_));
 sg13g2_o21ai_1 _24685_ (.B1(_06307_),
    .Y(_01883_),
    .A1(net650),
    .A2(net354));
 sg13g2_mux2_1 _24686_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .S(net354),
    .X(_01884_));
 sg13g2_nand2_1 _24687_ (.Y(_06308_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .B(_06305_));
 sg13g2_o21ai_1 _24688_ (.B1(_06308_),
    .Y(_01885_),
    .A1(net676),
    .A2(_06306_));
 sg13g2_nand2_1 _24689_ (.Y(_06309_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .B(_06305_));
 sg13g2_o21ai_1 _24690_ (.B1(_06309_),
    .Y(_01886_),
    .A1(net730),
    .A2(net354));
 sg13g2_mux2_1 _24691_ (.A0(net726),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .S(net354),
    .X(_01887_));
 sg13g2_nand2_1 _24692_ (.Y(_06310_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .B(_06305_));
 sg13g2_o21ai_1 _24693_ (.B1(_06310_),
    .Y(_01888_),
    .A1(net846),
    .A2(_06306_));
 sg13g2_mux2_1 _24694_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .S(net354),
    .X(_01889_));
 sg13g2_mux2_1 _24695_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .S(net354),
    .X(_01890_));
 sg13g2_mux2_1 _24696_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .S(net354),
    .X(_01891_));
 sg13g2_mux2_1 _24697_ (.A0(net838),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .S(net354),
    .X(_01892_));
 sg13g2_mux2_1 _24698_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .S(_06305_),
    .X(_01893_));
 sg13g2_mux2_1 _24699_ (.A0(net458),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .S(_06305_),
    .X(_01894_));
 sg13g2_nand3_1 _24700_ (.B(_05911_),
    .C(_06092_),
    .A(_05854_),
    .Y(_06311_));
 sg13g2_buf_2 _24701_ (.A(_06311_),
    .X(_06312_));
 sg13g2_buf_1 _24702_ (.A(_06312_),
    .X(_06313_));
 sg13g2_nand2_1 _24703_ (.Y(_06314_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .B(_06312_));
 sg13g2_o21ai_1 _24704_ (.B1(_06314_),
    .Y(_01895_),
    .A1(_03865_),
    .A2(net250));
 sg13g2_mux2_1 _24705_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .S(net250),
    .X(_01896_));
 sg13g2_nand2_1 _24706_ (.Y(_06315_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .B(_06312_));
 sg13g2_o21ai_1 _24707_ (.B1(_06315_),
    .Y(_01897_),
    .A1(net676),
    .A2(_06313_));
 sg13g2_nand2_1 _24708_ (.Y(_06316_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .B(_06312_));
 sg13g2_o21ai_1 _24709_ (.B1(_06316_),
    .Y(_01898_),
    .A1(_02970_),
    .A2(net250));
 sg13g2_mux2_1 _24710_ (.A0(net726),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .S(net250),
    .X(_01899_));
 sg13g2_nand2_1 _24711_ (.Y(_06317_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .B(_06312_));
 sg13g2_o21ai_1 _24712_ (.B1(_06317_),
    .Y(_01900_),
    .A1(net846),
    .A2(_06313_));
 sg13g2_mux2_1 _24713_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .S(net250),
    .X(_01901_));
 sg13g2_mux2_1 _24714_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .S(net250),
    .X(_01902_));
 sg13g2_mux2_1 _24715_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .S(net250),
    .X(_01903_));
 sg13g2_mux2_1 _24716_ (.A0(net838),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .S(net250),
    .X(_01904_));
 sg13g2_mux2_1 _24717_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .S(_06312_),
    .X(_01905_));
 sg13g2_mux2_1 _24718_ (.A0(_03585_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .S(_06312_),
    .X(_01906_));
 sg13g2_buf_1 _24719_ (.A(net596),
    .X(_06318_));
 sg13g2_mux2_1 _24720_ (.A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(net488),
    .S(_05889_),
    .X(_01907_));
 sg13g2_mux2_1 _24721_ (.A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(net488),
    .S(_05898_),
    .X(_01908_));
 sg13g2_mux2_1 _24722_ (.A0(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A1(net488),
    .S(_05908_),
    .X(_01909_));
 sg13g2_mux2_1 _24723_ (.A0(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A1(net488),
    .S(_05915_),
    .X(_01910_));
 sg13g2_mux2_1 _24724_ (.A0(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .A1(net488),
    .S(_05920_),
    .X(_01911_));
 sg13g2_mux2_1 _24725_ (.A0(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A1(net488),
    .S(_05925_),
    .X(_01912_));
 sg13g2_mux2_1 _24726_ (.A0(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .A1(net488),
    .S(_05931_),
    .X(_01913_));
 sg13g2_mux2_1 _24727_ (.A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(_06318_),
    .S(_05938_),
    .X(_01914_));
 sg13g2_mux2_1 _24728_ (.A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(_06318_),
    .S(_05943_),
    .X(_01915_));
 sg13g2_mux2_1 _24729_ (.A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(net488),
    .S(_05947_),
    .X(_01916_));
 sg13g2_buf_1 _24730_ (.A(net596),
    .X(_06319_));
 sg13g2_mux2_1 _24731_ (.A0(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A1(net487),
    .S(_05957_),
    .X(_01917_));
 sg13g2_mux2_1 _24732_ (.A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(net487),
    .S(_05961_),
    .X(_01918_));
 sg13g2_mux2_1 _24733_ (.A0(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .A1(net487),
    .S(_05968_),
    .X(_01919_));
 sg13g2_mux2_1 _24734_ (.A0(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .A1(_06319_),
    .S(_05972_),
    .X(_01920_));
 sg13g2_mux2_1 _24735_ (.A0(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .A1(net487),
    .S(_05975_),
    .X(_01921_));
 sg13g2_mux2_1 _24736_ (.A0(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .A1(net487),
    .S(_05979_),
    .X(_01922_));
 sg13g2_mux2_1 _24737_ (.A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(net487),
    .S(_05984_),
    .X(_01923_));
 sg13g2_mux2_1 _24738_ (.A0(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A1(net487),
    .S(_05989_),
    .X(_01924_));
 sg13g2_mux2_1 _24739_ (.A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(_06319_),
    .S(_05995_),
    .X(_01925_));
 sg13g2_mux2_1 _24740_ (.A0(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A1(net487),
    .S(_05999_),
    .X(_01926_));
 sg13g2_buf_1 _24741_ (.A(net596),
    .X(_06320_));
 sg13g2_mux2_1 _24742_ (.A0(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A1(net486),
    .S(_06008_),
    .X(_01927_));
 sg13g2_mux2_1 _24743_ (.A0(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .A1(net486),
    .S(_06012_),
    .X(_01928_));
 sg13g2_mux2_1 _24744_ (.A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(_06320_),
    .S(_06017_),
    .X(_01929_));
 sg13g2_mux2_1 _24745_ (.A0(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A1(_06320_),
    .S(_06021_),
    .X(_01930_));
 sg13g2_mux2_1 _24746_ (.A0(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .A1(net486),
    .S(_06024_),
    .X(_01931_));
 sg13g2_mux2_1 _24747_ (.A0(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A1(net486),
    .S(_06027_),
    .X(_01932_));
 sg13g2_mux2_1 _24748_ (.A0(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .A1(net486),
    .S(_06031_),
    .X(_01933_));
 sg13g2_mux2_1 _24749_ (.A0(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .A1(net486),
    .S(_06036_),
    .X(_01934_));
 sg13g2_mux2_1 _24750_ (.A0(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .A1(net486),
    .S(_06042_),
    .X(_01935_));
 sg13g2_mux2_1 _24751_ (.A0(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .A1(net486),
    .S(_06047_),
    .X(_01936_));
 sg13g2_mux2_1 _24752_ (.A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(_03590_),
    .S(_06050_),
    .X(_01937_));
 sg13g2_mux2_1 _24753_ (.A0(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A1(net596),
    .S(_06053_),
    .X(_01938_));
 sg13g2_nor2_1 _24754_ (.A(net1028),
    .B(_09261_),
    .Y(_06321_));
 sg13g2_and3_1 _24755_ (.X(_06322_),
    .A(net1042),
    .B(_00233_),
    .C(_06321_));
 sg13g2_buf_1 _24756_ (.A(_06322_),
    .X(_06323_));
 sg13g2_and2_1 _24757_ (.A(net891),
    .B(_06323_),
    .X(_06324_));
 sg13g2_buf_2 _24758_ (.A(_06324_),
    .X(_06325_));
 sg13g2_nand3_1 _24759_ (.B(_10124_),
    .C(_06325_),
    .A(net960),
    .Y(_06326_));
 sg13g2_buf_1 _24760_ (.A(_06326_),
    .X(_06327_));
 sg13g2_mux2_1 _24761_ (.A0(net884),
    .A1(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .S(_06327_),
    .X(_01955_));
 sg13g2_mux2_1 _24762_ (.A0(net883),
    .A1(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .S(_06327_),
    .X(_01956_));
 sg13g2_mux2_1 _24763_ (.A0(net882),
    .A1(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .S(_06327_),
    .X(_01957_));
 sg13g2_mux2_1 _24764_ (.A0(net888),
    .A1(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .S(_06327_),
    .X(_01958_));
 sg13g2_nand3_1 _24765_ (.B(_05178_),
    .C(_06325_),
    .A(net960),
    .Y(_06328_));
 sg13g2_buf_2 _24766_ (.A(_06328_),
    .X(_06329_));
 sg13g2_mux2_1 _24767_ (.A0(net885),
    .A1(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .S(_06329_),
    .X(_01959_));
 sg13g2_mux2_1 _24768_ (.A0(net884),
    .A1(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .S(_06329_),
    .X(_01960_));
 sg13g2_mux2_1 _24769_ (.A0(net883),
    .A1(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .S(_06329_),
    .X(_01961_));
 sg13g2_mux2_1 _24770_ (.A0(net882),
    .A1(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .S(_06329_),
    .X(_01962_));
 sg13g2_mux2_1 _24771_ (.A0(net888),
    .A1(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .S(_06329_),
    .X(_01963_));
 sg13g2_nand2_1 _24772_ (.Y(_06330_),
    .A(_04931_),
    .B(_06325_));
 sg13g2_buf_1 _24773_ (.A(_06330_),
    .X(_06331_));
 sg13g2_mux2_1 _24774_ (.A0(net890),
    .A1(_04932_),
    .S(net76),
    .X(_01964_));
 sg13g2_buf_1 _24775_ (.A(\cpu.gpio.r_spi_miso_src[0][1] ),
    .X(_06332_));
 sg13g2_nand2_1 _24776_ (.Y(_06333_),
    .A(_06332_),
    .B(net76));
 sg13g2_o21ai_1 _24777_ (.B1(_06333_),
    .Y(_01965_),
    .A1(net762),
    .A2(net76));
 sg13g2_mux2_1 _24778_ (.A0(net886),
    .A1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .S(net76),
    .X(_01966_));
 sg13g2_mux2_1 _24779_ (.A0(net885),
    .A1(\cpu.gpio.r_spi_miso_src[0][3] ),
    .S(net76),
    .X(_01967_));
 sg13g2_mux2_1 _24780_ (.A0(net884),
    .A1(_05573_),
    .S(net76),
    .X(_01968_));
 sg13g2_buf_1 _24781_ (.A(\cpu.gpio.r_spi_miso_src[1][1] ),
    .X(_06334_));
 sg13g2_mux2_1 _24782_ (.A0(net883),
    .A1(_06334_),
    .S(net76),
    .X(_01969_));
 sg13g2_mux2_1 _24783_ (.A0(net882),
    .A1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .S(_06331_),
    .X(_01970_));
 sg13g2_mux2_1 _24784_ (.A0(_10105_),
    .A1(\cpu.gpio.r_spi_miso_src[1][3] ),
    .S(net76),
    .X(_01971_));
 sg13g2_nand2_1 _24785_ (.Y(_06335_),
    .A(net443),
    .B(_06325_));
 sg13g2_buf_1 _24786_ (.A(_06335_),
    .X(_06336_));
 sg13g2_mux2_1 _24787_ (.A0(net890),
    .A1(_04937_),
    .S(net75),
    .X(_01972_));
 sg13g2_nand2_1 _24788_ (.Y(_06337_),
    .A(_05361_),
    .B(net75));
 sg13g2_o21ai_1 _24789_ (.B1(_06337_),
    .Y(_01973_),
    .A1(net762),
    .A2(net75));
 sg13g2_mux2_1 _24790_ (.A0(net886),
    .A1(_05448_),
    .S(net75),
    .X(_01974_));
 sg13g2_mux2_1 _24791_ (.A0(net885),
    .A1(_05522_),
    .S(net75),
    .X(_01975_));
 sg13g2_mux2_1 _24792_ (.A0(net884),
    .A1(_05576_),
    .S(net75),
    .X(_01976_));
 sg13g2_mux2_1 _24793_ (.A0(net883),
    .A1(_05646_),
    .S(net75),
    .X(_01977_));
 sg13g2_mux2_1 _24794_ (.A0(net882),
    .A1(_05720_),
    .S(_06336_),
    .X(_01978_));
 sg13g2_mux2_1 _24795_ (.A0(net888),
    .A1(_05094_),
    .S(net75),
    .X(_01979_));
 sg13g2_nand2_1 _24796_ (.Y(_06338_),
    .A(net446),
    .B(_06325_));
 sg13g2_buf_1 _24797_ (.A(_06338_),
    .X(_06339_));
 sg13g2_mux2_1 _24798_ (.A0(net890),
    .A1(_04923_),
    .S(net74),
    .X(_01980_));
 sg13g2_buf_1 _24799_ (.A(\cpu.gpio.r_src_io[6][1] ),
    .X(_06340_));
 sg13g2_nand2_1 _24800_ (.Y(_06341_),
    .A(_06340_),
    .B(net74));
 sg13g2_o21ai_1 _24801_ (.B1(_06341_),
    .Y(_01981_),
    .A1(net887),
    .A2(net74));
 sg13g2_mux2_1 _24802_ (.A0(net886),
    .A1(\cpu.gpio.r_src_io[6][2] ),
    .S(_06339_),
    .X(_01982_));
 sg13g2_mux2_1 _24803_ (.A0(net885),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .S(net74),
    .X(_01983_));
 sg13g2_mux2_1 _24804_ (.A0(net884),
    .A1(_05581_),
    .S(net74),
    .X(_01984_));
 sg13g2_buf_1 _24805_ (.A(\cpu.gpio.r_src_io[7][1] ),
    .X(_06342_));
 sg13g2_mux2_1 _24806_ (.A0(net883),
    .A1(_06342_),
    .S(net74),
    .X(_01985_));
 sg13g2_mux2_1 _24807_ (.A0(net882),
    .A1(\cpu.gpio.r_src_io[7][2] ),
    .S(net74),
    .X(_01986_));
 sg13g2_mux2_1 _24808_ (.A0(net888),
    .A1(\cpu.gpio.r_src_io[7][3] ),
    .S(net74),
    .X(_01987_));
 sg13g2_and3_1 _24809_ (.X(_06343_),
    .A(net651),
    .B(net391),
    .C(_06325_));
 sg13g2_buf_1 _24810_ (.A(_06343_),
    .X(_06344_));
 sg13g2_mux2_1 _24811_ (.A0(_05570_),
    .A1(net992),
    .S(_06344_),
    .X(_01988_));
 sg13g2_buf_1 _24812_ (.A(\cpu.gpio.r_src_o[3][1] ),
    .X(_06345_));
 sg13g2_mux2_1 _24813_ (.A0(_06345_),
    .A1(_12136_),
    .S(_06344_),
    .X(_01989_));
 sg13g2_mux2_1 _24814_ (.A0(\cpu.gpio.r_src_o[3][2] ),
    .A1(net989),
    .S(_06344_),
    .X(_01990_));
 sg13g2_mux2_1 _24815_ (.A0(\cpu.gpio.r_src_o[3][3] ),
    .A1(net851),
    .S(_06344_),
    .X(_01991_));
 sg13g2_nand2_1 _24816_ (.Y(_06346_),
    .A(_04914_),
    .B(_06325_));
 sg13g2_buf_1 _24817_ (.A(_06346_),
    .X(_06347_));
 sg13g2_mux2_1 _24818_ (.A0(_10049_),
    .A1(_04915_),
    .S(_06347_),
    .X(_01992_));
 sg13g2_buf_1 _24819_ (.A(\cpu.gpio.r_src_o[4][1] ),
    .X(_06348_));
 sg13g2_nand2_1 _24820_ (.Y(_06349_),
    .A(_06348_),
    .B(net73));
 sg13g2_o21ai_1 _24821_ (.B1(_06349_),
    .Y(_01993_),
    .A1(net887),
    .A2(net73));
 sg13g2_mux2_1 _24822_ (.A0(net886),
    .A1(\cpu.gpio.r_src_o[4][2] ),
    .S(net73),
    .X(_01994_));
 sg13g2_mux2_1 _24823_ (.A0(_10146_),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .S(net73),
    .X(_01995_));
 sg13g2_mux2_1 _24824_ (.A0(net884),
    .A1(_05580_),
    .S(net73),
    .X(_01996_));
 sg13g2_buf_1 _24825_ (.A(\cpu.gpio.r_src_o[5][1] ),
    .X(_06350_));
 sg13g2_mux2_1 _24826_ (.A0(net883),
    .A1(_06350_),
    .S(net73),
    .X(_01997_));
 sg13g2_mux2_1 _24827_ (.A0(net882),
    .A1(\cpu.gpio.r_src_o[5][2] ),
    .S(net73),
    .X(_01998_));
 sg13g2_mux2_1 _24828_ (.A0(net888),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .S(net73),
    .X(_01999_));
 sg13g2_nand2_2 _24829_ (.Y(_06351_),
    .A(_04934_),
    .B(_06325_));
 sg13g2_mux2_1 _24830_ (.A0(net884),
    .A1(_05575_),
    .S(_06351_),
    .X(_02004_));
 sg13g2_buf_1 _24831_ (.A(\cpu.gpio.r_src_o[7][1] ),
    .X(_06352_));
 sg13g2_mux2_1 _24832_ (.A0(net883),
    .A1(_06352_),
    .S(_06351_),
    .X(_02005_));
 sg13g2_mux2_1 _24833_ (.A0(_10164_),
    .A1(\cpu.gpio.r_src_o[7][2] ),
    .S(_06351_),
    .X(_02006_));
 sg13g2_mux2_1 _24834_ (.A0(net888),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .S(_06351_),
    .X(_02007_));
 sg13g2_buf_1 _24835_ (.A(net970),
    .X(_06353_));
 sg13g2_and2_1 _24836_ (.A(net786),
    .B(_08359_),
    .X(_06354_));
 sg13g2_buf_4 _24837_ (.X(_06355_),
    .A(_06354_));
 sg13g2_buf_1 _24838_ (.A(\cpu.icache.r_offset[2] ),
    .X(_06356_));
 sg13g2_buf_2 _24839_ (.A(_00251_),
    .X(_06357_));
 sg13g2_buf_1 _24840_ (.A(\cpu.icache.r_offset[1] ),
    .X(_06358_));
 sg13g2_buf_1 _24841_ (.A(\cpu.icache.r_offset[0] ),
    .X(_06359_));
 sg13g2_nand2b_1 _24842_ (.Y(_06360_),
    .B(_06359_),
    .A_N(_06358_));
 sg13g2_nor3_1 _24843_ (.A(_06356_),
    .B(_06357_),
    .C(_06360_),
    .Y(_06361_));
 sg13g2_buf_2 _24844_ (.A(_06361_),
    .X(_06362_));
 sg13g2_nand2_2 _24845_ (.Y(_06363_),
    .A(_06355_),
    .B(_06362_));
 sg13g2_mux2_1 _24846_ (.A0(net817),
    .A1(\cpu.icache.r_data[0][0] ),
    .S(_06363_),
    .X(_02011_));
 sg13g2_buf_1 _24847_ (.A(net972),
    .X(_06364_));
 sg13g2_buf_1 _24848_ (.A(_00252_),
    .X(_06365_));
 sg13g2_inv_1 _24849_ (.Y(_06366_),
    .A(_06365_));
 sg13g2_nand2_1 _24850_ (.Y(_06367_),
    .A(_06358_),
    .B(_06359_));
 sg13g2_nor3_1 _24851_ (.A(_06357_),
    .B(_06366_),
    .C(_06367_),
    .Y(_06368_));
 sg13g2_buf_2 _24852_ (.A(_06368_),
    .X(_06369_));
 sg13g2_nand2_2 _24853_ (.Y(_06370_),
    .A(_06355_),
    .B(_06369_));
 sg13g2_mux2_1 _24854_ (.A0(net816),
    .A1(\cpu.icache.r_data[0][10] ),
    .S(_06370_),
    .X(_02012_));
 sg13g2_buf_1 _24855_ (.A(net971),
    .X(_06371_));
 sg13g2_mux2_1 _24856_ (.A0(net815),
    .A1(\cpu.icache.r_data[0][11] ),
    .S(_06370_),
    .X(_02013_));
 sg13g2_nand2b_1 _24857_ (.Y(_06372_),
    .B(_06358_),
    .A_N(_06359_));
 sg13g2_nor3_1 _24858_ (.A(_06356_),
    .B(_06357_),
    .C(_06372_),
    .Y(_06373_));
 sg13g2_buf_2 _24859_ (.A(_06373_),
    .X(_06374_));
 sg13g2_nand2_2 _24860_ (.Y(_06375_),
    .A(_06355_),
    .B(_06374_));
 sg13g2_mux2_1 _24861_ (.A0(net817),
    .A1(\cpu.icache.r_data[0][12] ),
    .S(_06375_),
    .X(_02014_));
 sg13g2_buf_1 _24862_ (.A(_12156_),
    .X(_06376_));
 sg13g2_mux2_1 _24863_ (.A0(net814),
    .A1(\cpu.icache.r_data[0][13] ),
    .S(_06375_),
    .X(_02015_));
 sg13g2_mux2_1 _24864_ (.A0(net816),
    .A1(\cpu.icache.r_data[0][14] ),
    .S(_06375_),
    .X(_02016_));
 sg13g2_mux2_1 _24865_ (.A0(net815),
    .A1(\cpu.icache.r_data[0][15] ),
    .S(_06375_),
    .X(_02017_));
 sg13g2_nor3_1 _24866_ (.A(_06357_),
    .B(_06365_),
    .C(_06360_),
    .Y(_06377_));
 sg13g2_buf_2 _24867_ (.A(_06377_),
    .X(_06378_));
 sg13g2_nand2_2 _24868_ (.Y(_06379_),
    .A(_06355_),
    .B(_06378_));
 sg13g2_mux2_1 _24869_ (.A0(net817),
    .A1(\cpu.icache.r_data[0][16] ),
    .S(_06379_),
    .X(_02018_));
 sg13g2_mux2_1 _24870_ (.A0(net814),
    .A1(\cpu.icache.r_data[0][17] ),
    .S(_06379_),
    .X(_02019_));
 sg13g2_mux2_1 _24871_ (.A0(net816),
    .A1(\cpu.icache.r_data[0][18] ),
    .S(_06379_),
    .X(_02020_));
 sg13g2_mux2_1 _24872_ (.A0(net815),
    .A1(\cpu.icache.r_data[0][19] ),
    .S(_06379_),
    .X(_02021_));
 sg13g2_mux2_1 _24873_ (.A0(net814),
    .A1(\cpu.icache.r_data[0][1] ),
    .S(_06363_),
    .X(_02022_));
 sg13g2_nor4_1 _24874_ (.A(_06358_),
    .B(_06359_),
    .C(_06357_),
    .D(_06365_),
    .Y(_06380_));
 sg13g2_buf_2 _24875_ (.A(_06380_),
    .X(_06381_));
 sg13g2_nand2_2 _24876_ (.Y(_06382_),
    .A(_06355_),
    .B(_06381_));
 sg13g2_mux2_1 _24877_ (.A0(net817),
    .A1(\cpu.icache.r_data[0][20] ),
    .S(_06382_),
    .X(_02023_));
 sg13g2_mux2_1 _24878_ (.A0(net814),
    .A1(\cpu.icache.r_data[0][21] ),
    .S(_06382_),
    .X(_02024_));
 sg13g2_mux2_1 _24879_ (.A0(net816),
    .A1(\cpu.icache.r_data[0][22] ),
    .S(_06382_),
    .X(_02025_));
 sg13g2_mux2_1 _24880_ (.A0(net815),
    .A1(\cpu.icache.r_data[0][23] ),
    .S(_06382_),
    .X(_02026_));
 sg13g2_inv_1 _24881_ (.Y(_06383_),
    .A(\cpu.i_wstrobe_d ));
 sg13g2_nor3_1 _24882_ (.A(_06365_),
    .B(_06383_),
    .C(_06367_),
    .Y(_06384_));
 sg13g2_buf_2 _24883_ (.A(_06384_),
    .X(_06385_));
 sg13g2_nand2_1 _24884_ (.Y(_06386_),
    .A(_06355_),
    .B(_06385_));
 sg13g2_buf_1 _24885_ (.A(_06386_),
    .X(_06387_));
 sg13g2_buf_1 _24886_ (.A(_06387_),
    .X(_06388_));
 sg13g2_mux2_1 _24887_ (.A0(net817),
    .A1(\cpu.icache.r_data[0][24] ),
    .S(net387),
    .X(_02027_));
 sg13g2_mux2_1 _24888_ (.A0(net814),
    .A1(\cpu.icache.r_data[0][25] ),
    .S(net387),
    .X(_02028_));
 sg13g2_mux2_1 _24889_ (.A0(net816),
    .A1(\cpu.icache.r_data[0][26] ),
    .S(net387),
    .X(_02029_));
 sg13g2_mux2_1 _24890_ (.A0(net815),
    .A1(\cpu.icache.r_data[0][27] ),
    .S(net387),
    .X(_02030_));
 sg13g2_nor3_1 _24891_ (.A(_06357_),
    .B(_06365_),
    .C(_06372_),
    .Y(_06389_));
 sg13g2_buf_4 _24892_ (.X(_06390_),
    .A(_06389_));
 sg13g2_nand2_2 _24893_ (.Y(_06391_),
    .A(_06355_),
    .B(_06390_));
 sg13g2_mux2_1 _24894_ (.A0(_06353_),
    .A1(\cpu.icache.r_data[0][28] ),
    .S(_06391_),
    .X(_02031_));
 sg13g2_mux2_1 _24895_ (.A0(net814),
    .A1(\cpu.icache.r_data[0][29] ),
    .S(_06391_),
    .X(_02032_));
 sg13g2_mux2_1 _24896_ (.A0(net816),
    .A1(\cpu.icache.r_data[0][2] ),
    .S(_06363_),
    .X(_02033_));
 sg13g2_mux2_1 _24897_ (.A0(net816),
    .A1(\cpu.icache.r_data[0][30] ),
    .S(_06391_),
    .X(_02034_));
 sg13g2_mux2_1 _24898_ (.A0(net815),
    .A1(\cpu.icache.r_data[0][31] ),
    .S(_06391_),
    .X(_02035_));
 sg13g2_mux2_1 _24899_ (.A0(net815),
    .A1(\cpu.icache.r_data[0][3] ),
    .S(_06363_),
    .X(_02036_));
 sg13g2_nor4_1 _24900_ (.A(_06358_),
    .B(_06359_),
    .C(_06356_),
    .D(_06357_),
    .Y(_06392_));
 sg13g2_buf_2 _24901_ (.A(_06392_),
    .X(_06393_));
 sg13g2_nand2_2 _24902_ (.Y(_06394_),
    .A(_06355_),
    .B(_06393_));
 sg13g2_mux2_1 _24903_ (.A0(net817),
    .A1(\cpu.icache.r_data[0][4] ),
    .S(_06394_),
    .X(_02037_));
 sg13g2_mux2_1 _24904_ (.A0(net814),
    .A1(\cpu.icache.r_data[0][5] ),
    .S(_06394_),
    .X(_02038_));
 sg13g2_mux2_1 _24905_ (.A0(net816),
    .A1(\cpu.icache.r_data[0][6] ),
    .S(_06394_),
    .X(_02039_));
 sg13g2_mux2_1 _24906_ (.A0(net815),
    .A1(\cpu.icache.r_data[0][7] ),
    .S(_06394_),
    .X(_02040_));
 sg13g2_mux2_1 _24907_ (.A0(_06353_),
    .A1(\cpu.icache.r_data[0][8] ),
    .S(_06370_),
    .X(_02041_));
 sg13g2_mux2_1 _24908_ (.A0(net814),
    .A1(\cpu.icache.r_data[0][9] ),
    .S(_06370_),
    .X(_02042_));
 sg13g2_buf_1 _24909_ (.A(net970),
    .X(_06395_));
 sg13g2_and2_1 _24910_ (.A(net546),
    .B(_06362_),
    .X(_06396_));
 sg13g2_buf_1 _24911_ (.A(_06396_),
    .X(_06397_));
 sg13g2_mux2_1 _24912_ (.A0(\cpu.icache.r_data[1][0] ),
    .A1(net813),
    .S(_06397_),
    .X(_02043_));
 sg13g2_buf_1 _24913_ (.A(net972),
    .X(_06398_));
 sg13g2_and2_1 _24914_ (.A(_08682_),
    .B(_06369_),
    .X(_06399_));
 sg13g2_buf_1 _24915_ (.A(_06399_),
    .X(_06400_));
 sg13g2_mux2_1 _24916_ (.A0(\cpu.icache.r_data[1][10] ),
    .A1(net812),
    .S(_06400_),
    .X(_02044_));
 sg13g2_buf_1 _24917_ (.A(net971),
    .X(_06401_));
 sg13g2_mux2_1 _24918_ (.A0(\cpu.icache.r_data[1][11] ),
    .A1(net811),
    .S(_06400_),
    .X(_02045_));
 sg13g2_and2_1 _24919_ (.A(net546),
    .B(_06374_),
    .X(_06402_));
 sg13g2_buf_1 _24920_ (.A(_06402_),
    .X(_06403_));
 sg13g2_mux2_1 _24921_ (.A0(\cpu.icache.r_data[1][12] ),
    .A1(net813),
    .S(_06403_),
    .X(_02046_));
 sg13g2_buf_1 _24922_ (.A(_12156_),
    .X(_06404_));
 sg13g2_mux2_1 _24923_ (.A0(\cpu.icache.r_data[1][13] ),
    .A1(net810),
    .S(_06403_),
    .X(_02047_));
 sg13g2_mux2_1 _24924_ (.A0(\cpu.icache.r_data[1][14] ),
    .A1(net812),
    .S(_06403_),
    .X(_02048_));
 sg13g2_mux2_1 _24925_ (.A0(\cpu.icache.r_data[1][15] ),
    .A1(_06401_),
    .S(_06403_),
    .X(_02049_));
 sg13g2_and2_1 _24926_ (.A(net546),
    .B(_06378_),
    .X(_06405_));
 sg13g2_buf_2 _24927_ (.A(_06405_),
    .X(_06406_));
 sg13g2_mux2_1 _24928_ (.A0(\cpu.icache.r_data[1][16] ),
    .A1(net813),
    .S(_06406_),
    .X(_02050_));
 sg13g2_mux2_1 _24929_ (.A0(\cpu.icache.r_data[1][17] ),
    .A1(net810),
    .S(_06406_),
    .X(_02051_));
 sg13g2_mux2_1 _24930_ (.A0(\cpu.icache.r_data[1][18] ),
    .A1(net812),
    .S(_06406_),
    .X(_02052_));
 sg13g2_mux2_1 _24931_ (.A0(\cpu.icache.r_data[1][19] ),
    .A1(net811),
    .S(_06406_),
    .X(_02053_));
 sg13g2_mux2_1 _24932_ (.A0(\cpu.icache.r_data[1][1] ),
    .A1(net810),
    .S(_06397_),
    .X(_02054_));
 sg13g2_buf_1 _24933_ (.A(_12073_),
    .X(_06407_));
 sg13g2_and2_1 _24934_ (.A(net546),
    .B(_06381_),
    .X(_06408_));
 sg13g2_buf_1 _24935_ (.A(_06408_),
    .X(_06409_));
 sg13g2_mux2_1 _24936_ (.A0(\cpu.icache.r_data[1][20] ),
    .A1(net945),
    .S(_06409_),
    .X(_02055_));
 sg13g2_buf_1 _24937_ (.A(_12156_),
    .X(_06410_));
 sg13g2_mux2_1 _24938_ (.A0(\cpu.icache.r_data[1][21] ),
    .A1(net809),
    .S(_06409_),
    .X(_02056_));
 sg13g2_buf_1 _24939_ (.A(_12090_),
    .X(_06411_));
 sg13g2_mux2_1 _24940_ (.A0(\cpu.icache.r_data[1][22] ),
    .A1(net944),
    .S(_06409_),
    .X(_02057_));
 sg13g2_buf_1 _24941_ (.A(_12096_),
    .X(_06412_));
 sg13g2_mux2_1 _24942_ (.A0(\cpu.icache.r_data[1][23] ),
    .A1(net943),
    .S(_06409_),
    .X(_02058_));
 sg13g2_and2_1 _24943_ (.A(net546),
    .B(_06385_),
    .X(_06413_));
 sg13g2_buf_2 _24944_ (.A(_06413_),
    .X(_06414_));
 sg13g2_mux2_1 _24945_ (.A0(\cpu.icache.r_data[1][24] ),
    .A1(net945),
    .S(_06414_),
    .X(_02059_));
 sg13g2_mux2_1 _24946_ (.A0(\cpu.icache.r_data[1][25] ),
    .A1(net809),
    .S(_06414_),
    .X(_02060_));
 sg13g2_mux2_1 _24947_ (.A0(\cpu.icache.r_data[1][26] ),
    .A1(net944),
    .S(_06414_),
    .X(_02061_));
 sg13g2_mux2_1 _24948_ (.A0(\cpu.icache.r_data[1][27] ),
    .A1(net943),
    .S(_06414_),
    .X(_02062_));
 sg13g2_and2_1 _24949_ (.A(net546),
    .B(_06390_),
    .X(_06415_));
 sg13g2_buf_1 _24950_ (.A(_06415_),
    .X(_06416_));
 sg13g2_mux2_1 _24951_ (.A0(\cpu.icache.r_data[1][28] ),
    .A1(net945),
    .S(_06416_),
    .X(_02063_));
 sg13g2_mux2_1 _24952_ (.A0(\cpu.icache.r_data[1][29] ),
    .A1(_06410_),
    .S(_06416_),
    .X(_02064_));
 sg13g2_mux2_1 _24953_ (.A0(\cpu.icache.r_data[1][2] ),
    .A1(net944),
    .S(_06397_),
    .X(_02065_));
 sg13g2_mux2_1 _24954_ (.A0(\cpu.icache.r_data[1][30] ),
    .A1(net944),
    .S(_06416_),
    .X(_02066_));
 sg13g2_mux2_1 _24955_ (.A0(\cpu.icache.r_data[1][31] ),
    .A1(net943),
    .S(_06416_),
    .X(_02067_));
 sg13g2_mux2_1 _24956_ (.A0(\cpu.icache.r_data[1][3] ),
    .A1(net943),
    .S(_06397_),
    .X(_02068_));
 sg13g2_and2_1 _24957_ (.A(net546),
    .B(_06393_),
    .X(_06417_));
 sg13g2_buf_1 _24958_ (.A(_06417_),
    .X(_06418_));
 sg13g2_mux2_1 _24959_ (.A0(\cpu.icache.r_data[1][4] ),
    .A1(net945),
    .S(_06418_),
    .X(_02069_));
 sg13g2_mux2_1 _24960_ (.A0(\cpu.icache.r_data[1][5] ),
    .A1(net809),
    .S(_06418_),
    .X(_02070_));
 sg13g2_mux2_1 _24961_ (.A0(\cpu.icache.r_data[1][6] ),
    .A1(_06411_),
    .S(_06418_),
    .X(_02071_));
 sg13g2_mux2_1 _24962_ (.A0(\cpu.icache.r_data[1][7] ),
    .A1(net943),
    .S(_06418_),
    .X(_02072_));
 sg13g2_mux2_1 _24963_ (.A0(\cpu.icache.r_data[1][8] ),
    .A1(_06407_),
    .S(_06400_),
    .X(_02073_));
 sg13g2_mux2_1 _24964_ (.A0(\cpu.icache.r_data[1][9] ),
    .A1(_06410_),
    .S(_06400_),
    .X(_02074_));
 sg13g2_and2_1 _24965_ (.A(net480),
    .B(_06362_),
    .X(_06419_));
 sg13g2_buf_1 _24966_ (.A(_06419_),
    .X(_06420_));
 sg13g2_mux2_1 _24967_ (.A0(\cpu.icache.r_data[2][0] ),
    .A1(net945),
    .S(_06420_),
    .X(_02075_));
 sg13g2_and2_1 _24968_ (.A(_08685_),
    .B(_06369_),
    .X(_06421_));
 sg13g2_buf_1 _24969_ (.A(_06421_),
    .X(_06422_));
 sg13g2_mux2_1 _24970_ (.A0(\cpu.icache.r_data[2][10] ),
    .A1(_06411_),
    .S(_06422_),
    .X(_02076_));
 sg13g2_mux2_1 _24971_ (.A0(\cpu.icache.r_data[2][11] ),
    .A1(_06412_),
    .S(_06422_),
    .X(_02077_));
 sg13g2_and2_1 _24972_ (.A(net480),
    .B(_06374_),
    .X(_06423_));
 sg13g2_buf_1 _24973_ (.A(_06423_),
    .X(_06424_));
 sg13g2_mux2_1 _24974_ (.A0(\cpu.icache.r_data[2][12] ),
    .A1(_06407_),
    .S(_06424_),
    .X(_02078_));
 sg13g2_mux2_1 _24975_ (.A0(\cpu.icache.r_data[2][13] ),
    .A1(net809),
    .S(_06424_),
    .X(_02079_));
 sg13g2_mux2_1 _24976_ (.A0(\cpu.icache.r_data[2][14] ),
    .A1(net944),
    .S(_06424_),
    .X(_02080_));
 sg13g2_mux2_1 _24977_ (.A0(\cpu.icache.r_data[2][15] ),
    .A1(net943),
    .S(_06424_),
    .X(_02081_));
 sg13g2_and2_1 _24978_ (.A(net480),
    .B(_06378_),
    .X(_06425_));
 sg13g2_buf_1 _24979_ (.A(_06425_),
    .X(_06426_));
 sg13g2_mux2_1 _24980_ (.A0(\cpu.icache.r_data[2][16] ),
    .A1(net945),
    .S(_06426_),
    .X(_02082_));
 sg13g2_mux2_1 _24981_ (.A0(\cpu.icache.r_data[2][17] ),
    .A1(net809),
    .S(_06426_),
    .X(_02083_));
 sg13g2_mux2_1 _24982_ (.A0(\cpu.icache.r_data[2][18] ),
    .A1(net944),
    .S(_06426_),
    .X(_02084_));
 sg13g2_mux2_1 _24983_ (.A0(\cpu.icache.r_data[2][19] ),
    .A1(net943),
    .S(_06426_),
    .X(_02085_));
 sg13g2_mux2_1 _24984_ (.A0(\cpu.icache.r_data[2][1] ),
    .A1(net809),
    .S(_06420_),
    .X(_02086_));
 sg13g2_and2_1 _24985_ (.A(net480),
    .B(_06381_),
    .X(_06427_));
 sg13g2_buf_1 _24986_ (.A(_06427_),
    .X(_06428_));
 sg13g2_mux2_1 _24987_ (.A0(\cpu.icache.r_data[2][20] ),
    .A1(net945),
    .S(_06428_),
    .X(_02087_));
 sg13g2_mux2_1 _24988_ (.A0(\cpu.icache.r_data[2][21] ),
    .A1(net809),
    .S(_06428_),
    .X(_02088_));
 sg13g2_mux2_1 _24989_ (.A0(\cpu.icache.r_data[2][22] ),
    .A1(net944),
    .S(_06428_),
    .X(_02089_));
 sg13g2_mux2_1 _24990_ (.A0(\cpu.icache.r_data[2][23] ),
    .A1(net943),
    .S(_06428_),
    .X(_02090_));
 sg13g2_and2_1 _24991_ (.A(net480),
    .B(_06385_),
    .X(_06429_));
 sg13g2_buf_2 _24992_ (.A(_06429_),
    .X(_06430_));
 sg13g2_mux2_1 _24993_ (.A0(\cpu.icache.r_data[2][24] ),
    .A1(net945),
    .S(_06430_),
    .X(_02091_));
 sg13g2_mux2_1 _24994_ (.A0(\cpu.icache.r_data[2][25] ),
    .A1(net809),
    .S(_06430_),
    .X(_02092_));
 sg13g2_mux2_1 _24995_ (.A0(\cpu.icache.r_data[2][26] ),
    .A1(net944),
    .S(_06430_),
    .X(_02093_));
 sg13g2_mux2_1 _24996_ (.A0(\cpu.icache.r_data[2][27] ),
    .A1(_06412_),
    .S(_06430_),
    .X(_02094_));
 sg13g2_buf_1 _24997_ (.A(_12073_),
    .X(_06431_));
 sg13g2_and2_1 _24998_ (.A(net480),
    .B(_06390_),
    .X(_06432_));
 sg13g2_buf_1 _24999_ (.A(_06432_),
    .X(_06433_));
 sg13g2_mux2_1 _25000_ (.A0(\cpu.icache.r_data[2][28] ),
    .A1(net942),
    .S(_06433_),
    .X(_02095_));
 sg13g2_buf_1 _25001_ (.A(_12156_),
    .X(_06434_));
 sg13g2_mux2_1 _25002_ (.A0(\cpu.icache.r_data[2][29] ),
    .A1(net808),
    .S(_06433_),
    .X(_02096_));
 sg13g2_buf_1 _25003_ (.A(_12090_),
    .X(_06435_));
 sg13g2_mux2_1 _25004_ (.A0(\cpu.icache.r_data[2][2] ),
    .A1(net941),
    .S(_06420_),
    .X(_02097_));
 sg13g2_mux2_1 _25005_ (.A0(\cpu.icache.r_data[2][30] ),
    .A1(net941),
    .S(_06433_),
    .X(_02098_));
 sg13g2_buf_1 _25006_ (.A(_12096_),
    .X(_06436_));
 sg13g2_mux2_1 _25007_ (.A0(\cpu.icache.r_data[2][31] ),
    .A1(net940),
    .S(_06433_),
    .X(_02099_));
 sg13g2_mux2_1 _25008_ (.A0(\cpu.icache.r_data[2][3] ),
    .A1(net940),
    .S(_06420_),
    .X(_02100_));
 sg13g2_and2_1 _25009_ (.A(net480),
    .B(_06393_),
    .X(_06437_));
 sg13g2_buf_1 _25010_ (.A(_06437_),
    .X(_06438_));
 sg13g2_mux2_1 _25011_ (.A0(\cpu.icache.r_data[2][4] ),
    .A1(net942),
    .S(_06438_),
    .X(_02101_));
 sg13g2_mux2_1 _25012_ (.A0(\cpu.icache.r_data[2][5] ),
    .A1(net808),
    .S(_06438_),
    .X(_02102_));
 sg13g2_mux2_1 _25013_ (.A0(\cpu.icache.r_data[2][6] ),
    .A1(net941),
    .S(_06438_),
    .X(_02103_));
 sg13g2_mux2_1 _25014_ (.A0(\cpu.icache.r_data[2][7] ),
    .A1(net940),
    .S(_06438_),
    .X(_02104_));
 sg13g2_mux2_1 _25015_ (.A0(\cpu.icache.r_data[2][8] ),
    .A1(net942),
    .S(_06422_),
    .X(_02105_));
 sg13g2_mux2_1 _25016_ (.A0(\cpu.icache.r_data[2][9] ),
    .A1(net808),
    .S(_06422_),
    .X(_02106_));
 sg13g2_nand2_2 _25017_ (.Y(_06439_),
    .A(net425),
    .B(_06362_));
 sg13g2_mux2_1 _25018_ (.A0(net817),
    .A1(\cpu.icache.r_data[3][0] ),
    .S(_06439_),
    .X(_02107_));
 sg13g2_and2_1 _25019_ (.A(net425),
    .B(_06369_),
    .X(_06440_));
 sg13g2_buf_1 _25020_ (.A(_06440_),
    .X(_06441_));
 sg13g2_mux2_1 _25021_ (.A0(\cpu.icache.r_data[3][10] ),
    .A1(net941),
    .S(_06441_),
    .X(_02108_));
 sg13g2_mux2_1 _25022_ (.A0(\cpu.icache.r_data[3][11] ),
    .A1(_06436_),
    .S(_06441_),
    .X(_02109_));
 sg13g2_nand2_2 _25023_ (.Y(_06442_),
    .A(net425),
    .B(_06374_));
 sg13g2_mux2_1 _25024_ (.A0(net817),
    .A1(\cpu.icache.r_data[3][12] ),
    .S(_06442_),
    .X(_02110_));
 sg13g2_mux2_1 _25025_ (.A0(_06376_),
    .A1(\cpu.icache.r_data[3][13] ),
    .S(_06442_),
    .X(_02111_));
 sg13g2_mux2_1 _25026_ (.A0(_06364_),
    .A1(\cpu.icache.r_data[3][14] ),
    .S(_06442_),
    .X(_02112_));
 sg13g2_mux2_1 _25027_ (.A0(_06371_),
    .A1(\cpu.icache.r_data[3][15] ),
    .S(_06442_),
    .X(_02113_));
 sg13g2_buf_1 _25028_ (.A(_02835_),
    .X(_06443_));
 sg13g2_nand2_2 _25029_ (.Y(_06444_),
    .A(net425),
    .B(_06378_));
 sg13g2_mux2_1 _25030_ (.A0(net807),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(_06444_),
    .X(_02114_));
 sg13g2_mux2_1 _25031_ (.A0(_06376_),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(_06444_),
    .X(_02115_));
 sg13g2_mux2_1 _25032_ (.A0(_06364_),
    .A1(\cpu.icache.r_data[3][18] ),
    .S(_06444_),
    .X(_02116_));
 sg13g2_mux2_1 _25033_ (.A0(_06371_),
    .A1(\cpu.icache.r_data[3][19] ),
    .S(_06444_),
    .X(_02117_));
 sg13g2_buf_1 _25034_ (.A(_12156_),
    .X(_06445_));
 sg13g2_mux2_1 _25035_ (.A0(net806),
    .A1(\cpu.icache.r_data[3][1] ),
    .S(_06439_),
    .X(_02118_));
 sg13g2_nand2_2 _25036_ (.Y(_06446_),
    .A(net425),
    .B(_06381_));
 sg13g2_mux2_1 _25037_ (.A0(net807),
    .A1(\cpu.icache.r_data[3][20] ),
    .S(_06446_),
    .X(_02119_));
 sg13g2_mux2_1 _25038_ (.A0(net806),
    .A1(\cpu.icache.r_data[3][21] ),
    .S(_06446_),
    .X(_02120_));
 sg13g2_buf_1 _25039_ (.A(_02823_),
    .X(_06447_));
 sg13g2_mux2_1 _25040_ (.A0(net805),
    .A1(\cpu.icache.r_data[3][22] ),
    .S(_06446_),
    .X(_02121_));
 sg13g2_buf_1 _25041_ (.A(_02831_),
    .X(_06448_));
 sg13g2_mux2_1 _25042_ (.A0(net804),
    .A1(\cpu.icache.r_data[3][23] ),
    .S(_06446_),
    .X(_02122_));
 sg13g2_nand2_1 _25043_ (.Y(_06449_),
    .A(_08655_),
    .B(_06385_));
 sg13g2_buf_1 _25044_ (.A(_06449_),
    .X(_06450_));
 sg13g2_buf_1 _25045_ (.A(_06450_),
    .X(_06451_));
 sg13g2_mux2_1 _25046_ (.A0(net807),
    .A1(\cpu.icache.r_data[3][24] ),
    .S(net249),
    .X(_02123_));
 sg13g2_mux2_1 _25047_ (.A0(_06445_),
    .A1(\cpu.icache.r_data[3][25] ),
    .S(net249),
    .X(_02124_));
 sg13g2_mux2_1 _25048_ (.A0(net805),
    .A1(\cpu.icache.r_data[3][26] ),
    .S(net249),
    .X(_02125_));
 sg13g2_mux2_1 _25049_ (.A0(net804),
    .A1(\cpu.icache.r_data[3][27] ),
    .S(net249),
    .X(_02126_));
 sg13g2_nand2_2 _25050_ (.Y(_06452_),
    .A(net425),
    .B(_06390_));
 sg13g2_mux2_1 _25051_ (.A0(_06443_),
    .A1(\cpu.icache.r_data[3][28] ),
    .S(_06452_),
    .X(_02127_));
 sg13g2_mux2_1 _25052_ (.A0(net806),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(_06452_),
    .X(_02128_));
 sg13g2_mux2_1 _25053_ (.A0(net805),
    .A1(\cpu.icache.r_data[3][2] ),
    .S(_06439_),
    .X(_02129_));
 sg13g2_mux2_1 _25054_ (.A0(net805),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(_06452_),
    .X(_02130_));
 sg13g2_mux2_1 _25055_ (.A0(_06448_),
    .A1(\cpu.icache.r_data[3][31] ),
    .S(_06452_),
    .X(_02131_));
 sg13g2_mux2_1 _25056_ (.A0(net804),
    .A1(\cpu.icache.r_data[3][3] ),
    .S(_06439_),
    .X(_02132_));
 sg13g2_nand2_2 _25057_ (.Y(_06453_),
    .A(net425),
    .B(_06393_));
 sg13g2_mux2_1 _25058_ (.A0(_06443_),
    .A1(\cpu.icache.r_data[3][4] ),
    .S(_06453_),
    .X(_02133_));
 sg13g2_mux2_1 _25059_ (.A0(net806),
    .A1(\cpu.icache.r_data[3][5] ),
    .S(_06453_),
    .X(_02134_));
 sg13g2_mux2_1 _25060_ (.A0(_06447_),
    .A1(\cpu.icache.r_data[3][6] ),
    .S(_06453_),
    .X(_02135_));
 sg13g2_mux2_1 _25061_ (.A0(net804),
    .A1(\cpu.icache.r_data[3][7] ),
    .S(_06453_),
    .X(_02136_));
 sg13g2_mux2_1 _25062_ (.A0(\cpu.icache.r_data[3][8] ),
    .A1(net942),
    .S(_06441_),
    .X(_02137_));
 sg13g2_mux2_1 _25063_ (.A0(\cpu.icache.r_data[3][9] ),
    .A1(net808),
    .S(_06441_),
    .X(_02138_));
 sg13g2_nand2_2 _25064_ (.Y(_06454_),
    .A(net545),
    .B(_06362_));
 sg13g2_mux2_1 _25065_ (.A0(net807),
    .A1(\cpu.icache.r_data[4][0] ),
    .S(_06454_),
    .X(_02139_));
 sg13g2_and2_1 _25066_ (.A(net545),
    .B(_06369_),
    .X(_06455_));
 sg13g2_buf_1 _25067_ (.A(_06455_),
    .X(_06456_));
 sg13g2_mux2_1 _25068_ (.A0(\cpu.icache.r_data[4][10] ),
    .A1(_06435_),
    .S(_06456_),
    .X(_02140_));
 sg13g2_mux2_1 _25069_ (.A0(\cpu.icache.r_data[4][11] ),
    .A1(net940),
    .S(_06456_),
    .X(_02141_));
 sg13g2_nand2_2 _25070_ (.Y(_06457_),
    .A(net545),
    .B(_06374_));
 sg13g2_mux2_1 _25071_ (.A0(net807),
    .A1(\cpu.icache.r_data[4][12] ),
    .S(_06457_),
    .X(_02142_));
 sg13g2_mux2_1 _25072_ (.A0(net806),
    .A1(\cpu.icache.r_data[4][13] ),
    .S(_06457_),
    .X(_02143_));
 sg13g2_mux2_1 _25073_ (.A0(net805),
    .A1(\cpu.icache.r_data[4][14] ),
    .S(_06457_),
    .X(_02144_));
 sg13g2_mux2_1 _25074_ (.A0(net804),
    .A1(\cpu.icache.r_data[4][15] ),
    .S(_06457_),
    .X(_02145_));
 sg13g2_nand2_2 _25075_ (.Y(_06458_),
    .A(net545),
    .B(_06378_));
 sg13g2_mux2_1 _25076_ (.A0(net807),
    .A1(\cpu.icache.r_data[4][16] ),
    .S(_06458_),
    .X(_02146_));
 sg13g2_mux2_1 _25077_ (.A0(net806),
    .A1(\cpu.icache.r_data[4][17] ),
    .S(_06458_),
    .X(_02147_));
 sg13g2_mux2_1 _25078_ (.A0(net805),
    .A1(\cpu.icache.r_data[4][18] ),
    .S(_06458_),
    .X(_02148_));
 sg13g2_mux2_1 _25079_ (.A0(net804),
    .A1(\cpu.icache.r_data[4][19] ),
    .S(_06458_),
    .X(_02149_));
 sg13g2_mux2_1 _25080_ (.A0(net806),
    .A1(\cpu.icache.r_data[4][1] ),
    .S(_06454_),
    .X(_02150_));
 sg13g2_nand2_2 _25081_ (.Y(_06459_),
    .A(net545),
    .B(_06381_));
 sg13g2_mux2_1 _25082_ (.A0(net807),
    .A1(\cpu.icache.r_data[4][20] ),
    .S(_06459_),
    .X(_02151_));
 sg13g2_mux2_1 _25083_ (.A0(net806),
    .A1(\cpu.icache.r_data[4][21] ),
    .S(_06459_),
    .X(_02152_));
 sg13g2_mux2_1 _25084_ (.A0(net805),
    .A1(\cpu.icache.r_data[4][22] ),
    .S(_06459_),
    .X(_02153_));
 sg13g2_mux2_1 _25085_ (.A0(net804),
    .A1(\cpu.icache.r_data[4][23] ),
    .S(_06459_),
    .X(_02154_));
 sg13g2_and2_1 _25086_ (.A(net545),
    .B(_06385_),
    .X(_06460_));
 sg13g2_buf_2 _25087_ (.A(_06460_),
    .X(_06461_));
 sg13g2_mux2_1 _25088_ (.A0(\cpu.icache.r_data[4][24] ),
    .A1(net942),
    .S(_06461_),
    .X(_02155_));
 sg13g2_mux2_1 _25089_ (.A0(\cpu.icache.r_data[4][25] ),
    .A1(net808),
    .S(_06461_),
    .X(_02156_));
 sg13g2_mux2_1 _25090_ (.A0(\cpu.icache.r_data[4][26] ),
    .A1(net941),
    .S(_06461_),
    .X(_02157_));
 sg13g2_mux2_1 _25091_ (.A0(\cpu.icache.r_data[4][27] ),
    .A1(net940),
    .S(_06461_),
    .X(_02158_));
 sg13g2_nand2_2 _25092_ (.Y(_06462_),
    .A(_08683_),
    .B(_06390_));
 sg13g2_mux2_1 _25093_ (.A0(net807),
    .A1(\cpu.icache.r_data[4][28] ),
    .S(_06462_),
    .X(_02159_));
 sg13g2_mux2_1 _25094_ (.A0(_06445_),
    .A1(\cpu.icache.r_data[4][29] ),
    .S(_06462_),
    .X(_02160_));
 sg13g2_mux2_1 _25095_ (.A0(net805),
    .A1(\cpu.icache.r_data[4][2] ),
    .S(_06454_),
    .X(_02161_));
 sg13g2_mux2_1 _25096_ (.A0(_06447_),
    .A1(\cpu.icache.r_data[4][30] ),
    .S(_06462_),
    .X(_02162_));
 sg13g2_mux2_1 _25097_ (.A0(_06448_),
    .A1(\cpu.icache.r_data[4][31] ),
    .S(_06462_),
    .X(_02163_));
 sg13g2_mux2_1 _25098_ (.A0(net804),
    .A1(\cpu.icache.r_data[4][3] ),
    .S(_06454_),
    .X(_02164_));
 sg13g2_buf_1 _25099_ (.A(_02835_),
    .X(_06463_));
 sg13g2_nand2_2 _25100_ (.Y(_06464_),
    .A(net545),
    .B(_06393_));
 sg13g2_mux2_1 _25101_ (.A0(net803),
    .A1(\cpu.icache.r_data[4][4] ),
    .S(_06464_),
    .X(_02165_));
 sg13g2_buf_1 _25102_ (.A(_12156_),
    .X(_06465_));
 sg13g2_mux2_1 _25103_ (.A0(net802),
    .A1(\cpu.icache.r_data[4][5] ),
    .S(_06464_),
    .X(_02166_));
 sg13g2_buf_1 _25104_ (.A(_02823_),
    .X(_06466_));
 sg13g2_mux2_1 _25105_ (.A0(net801),
    .A1(\cpu.icache.r_data[4][6] ),
    .S(_06464_),
    .X(_02167_));
 sg13g2_buf_1 _25106_ (.A(_02831_),
    .X(_06467_));
 sg13g2_mux2_1 _25107_ (.A0(net800),
    .A1(\cpu.icache.r_data[4][7] ),
    .S(_06464_),
    .X(_02168_));
 sg13g2_mux2_1 _25108_ (.A0(\cpu.icache.r_data[4][8] ),
    .A1(net942),
    .S(_06456_),
    .X(_02169_));
 sg13g2_mux2_1 _25109_ (.A0(\cpu.icache.r_data[4][9] ),
    .A1(net808),
    .S(_06456_),
    .X(_02170_));
 sg13g2_nand2_2 _25110_ (.Y(_06468_),
    .A(net542),
    .B(_06362_));
 sg13g2_mux2_1 _25111_ (.A0(net803),
    .A1(\cpu.icache.r_data[5][0] ),
    .S(_06468_),
    .X(_02171_));
 sg13g2_nand2_2 _25112_ (.Y(_06469_),
    .A(net542),
    .B(_06369_));
 sg13g2_mux2_1 _25113_ (.A0(_06466_),
    .A1(\cpu.icache.r_data[5][10] ),
    .S(_06469_),
    .X(_02172_));
 sg13g2_mux2_1 _25114_ (.A0(_06467_),
    .A1(\cpu.icache.r_data[5][11] ),
    .S(_06469_),
    .X(_02173_));
 sg13g2_nand2_2 _25115_ (.Y(_06470_),
    .A(net542),
    .B(_06374_));
 sg13g2_mux2_1 _25116_ (.A0(net803),
    .A1(\cpu.icache.r_data[5][12] ),
    .S(_06470_),
    .X(_02174_));
 sg13g2_mux2_1 _25117_ (.A0(_06465_),
    .A1(\cpu.icache.r_data[5][13] ),
    .S(_06470_),
    .X(_02175_));
 sg13g2_mux2_1 _25118_ (.A0(net801),
    .A1(\cpu.icache.r_data[5][14] ),
    .S(_06470_),
    .X(_02176_));
 sg13g2_mux2_1 _25119_ (.A0(net800),
    .A1(\cpu.icache.r_data[5][15] ),
    .S(_06470_),
    .X(_02177_));
 sg13g2_nand2_2 _25120_ (.Y(_06471_),
    .A(net542),
    .B(_06378_));
 sg13g2_mux2_1 _25121_ (.A0(net803),
    .A1(\cpu.icache.r_data[5][16] ),
    .S(_06471_),
    .X(_02178_));
 sg13g2_mux2_1 _25122_ (.A0(net802),
    .A1(\cpu.icache.r_data[5][17] ),
    .S(_06471_),
    .X(_02179_));
 sg13g2_mux2_1 _25123_ (.A0(net801),
    .A1(\cpu.icache.r_data[5][18] ),
    .S(_06471_),
    .X(_02180_));
 sg13g2_mux2_1 _25124_ (.A0(net800),
    .A1(\cpu.icache.r_data[5][19] ),
    .S(_06471_),
    .X(_02181_));
 sg13g2_mux2_1 _25125_ (.A0(_06465_),
    .A1(\cpu.icache.r_data[5][1] ),
    .S(_06468_),
    .X(_02182_));
 sg13g2_nand2_2 _25126_ (.Y(_06472_),
    .A(net542),
    .B(_06381_));
 sg13g2_mux2_1 _25127_ (.A0(net803),
    .A1(\cpu.icache.r_data[5][20] ),
    .S(_06472_),
    .X(_02183_));
 sg13g2_mux2_1 _25128_ (.A0(net802),
    .A1(\cpu.icache.r_data[5][21] ),
    .S(_06472_),
    .X(_02184_));
 sg13g2_mux2_1 _25129_ (.A0(net801),
    .A1(\cpu.icache.r_data[5][22] ),
    .S(_06472_),
    .X(_02185_));
 sg13g2_mux2_1 _25130_ (.A0(net800),
    .A1(\cpu.icache.r_data[5][23] ),
    .S(_06472_),
    .X(_02186_));
 sg13g2_nand2_1 _25131_ (.Y(_06473_),
    .A(net542),
    .B(_06385_));
 sg13g2_buf_2 _25132_ (.A(_06473_),
    .X(_06474_));
 sg13g2_mux2_1 _25133_ (.A0(_06463_),
    .A1(\cpu.icache.r_data[5][24] ),
    .S(_06474_),
    .X(_02187_));
 sg13g2_mux2_1 _25134_ (.A0(net802),
    .A1(\cpu.icache.r_data[5][25] ),
    .S(_06474_),
    .X(_02188_));
 sg13g2_mux2_1 _25135_ (.A0(net801),
    .A1(\cpu.icache.r_data[5][26] ),
    .S(_06474_),
    .X(_02189_));
 sg13g2_mux2_1 _25136_ (.A0(net800),
    .A1(\cpu.icache.r_data[5][27] ),
    .S(_06474_),
    .X(_02190_));
 sg13g2_nand2_2 _25137_ (.Y(_06475_),
    .A(net542),
    .B(_06390_));
 sg13g2_mux2_1 _25138_ (.A0(_06463_),
    .A1(\cpu.icache.r_data[5][28] ),
    .S(_06475_),
    .X(_02191_));
 sg13g2_mux2_1 _25139_ (.A0(net802),
    .A1(\cpu.icache.r_data[5][29] ),
    .S(_06475_),
    .X(_02192_));
 sg13g2_mux2_1 _25140_ (.A0(net801),
    .A1(\cpu.icache.r_data[5][2] ),
    .S(_06468_),
    .X(_02193_));
 sg13g2_mux2_1 _25141_ (.A0(_06466_),
    .A1(\cpu.icache.r_data[5][30] ),
    .S(_06475_),
    .X(_02194_));
 sg13g2_mux2_1 _25142_ (.A0(net800),
    .A1(\cpu.icache.r_data[5][31] ),
    .S(_06475_),
    .X(_02195_));
 sg13g2_mux2_1 _25143_ (.A0(net800),
    .A1(\cpu.icache.r_data[5][3] ),
    .S(_06468_),
    .X(_02196_));
 sg13g2_nand2_2 _25144_ (.Y(_06476_),
    .A(_09078_),
    .B(_06393_));
 sg13g2_mux2_1 _25145_ (.A0(net803),
    .A1(\cpu.icache.r_data[5][4] ),
    .S(_06476_),
    .X(_02197_));
 sg13g2_mux2_1 _25146_ (.A0(net802),
    .A1(\cpu.icache.r_data[5][5] ),
    .S(_06476_),
    .X(_02198_));
 sg13g2_mux2_1 _25147_ (.A0(net801),
    .A1(\cpu.icache.r_data[5][6] ),
    .S(_06476_),
    .X(_02199_));
 sg13g2_mux2_1 _25148_ (.A0(net800),
    .A1(\cpu.icache.r_data[5][7] ),
    .S(_06476_),
    .X(_02200_));
 sg13g2_mux2_1 _25149_ (.A0(net803),
    .A1(\cpu.icache.r_data[5][8] ),
    .S(_06469_),
    .X(_02201_));
 sg13g2_mux2_1 _25150_ (.A0(net802),
    .A1(\cpu.icache.r_data[5][9] ),
    .S(_06469_),
    .X(_02202_));
 sg13g2_nand2_2 _25151_ (.Y(_06477_),
    .A(net544),
    .B(_06362_));
 sg13g2_mux2_1 _25152_ (.A0(net803),
    .A1(\cpu.icache.r_data[6][0] ),
    .S(_06477_),
    .X(_02203_));
 sg13g2_nand2_2 _25153_ (.Y(_06478_),
    .A(net544),
    .B(_06369_));
 sg13g2_mux2_1 _25154_ (.A0(net801),
    .A1(\cpu.icache.r_data[6][10] ),
    .S(_06478_),
    .X(_02204_));
 sg13g2_mux2_1 _25155_ (.A0(_06467_),
    .A1(\cpu.icache.r_data[6][11] ),
    .S(_06478_),
    .X(_02205_));
 sg13g2_nand2_2 _25156_ (.Y(_06479_),
    .A(net544),
    .B(_06374_));
 sg13g2_mux2_1 _25157_ (.A0(net813),
    .A1(\cpu.icache.r_data[6][12] ),
    .S(_06479_),
    .X(_02206_));
 sg13g2_mux2_1 _25158_ (.A0(net802),
    .A1(\cpu.icache.r_data[6][13] ),
    .S(_06479_),
    .X(_02207_));
 sg13g2_mux2_1 _25159_ (.A0(net812),
    .A1(\cpu.icache.r_data[6][14] ),
    .S(_06479_),
    .X(_02208_));
 sg13g2_mux2_1 _25160_ (.A0(net811),
    .A1(\cpu.icache.r_data[6][15] ),
    .S(_06479_),
    .X(_02209_));
 sg13g2_nand2_2 _25161_ (.Y(_06480_),
    .A(net544),
    .B(_06378_));
 sg13g2_mux2_1 _25162_ (.A0(net813),
    .A1(\cpu.icache.r_data[6][16] ),
    .S(_06480_),
    .X(_02210_));
 sg13g2_mux2_1 _25163_ (.A0(net810),
    .A1(\cpu.icache.r_data[6][17] ),
    .S(_06480_),
    .X(_02211_));
 sg13g2_mux2_1 _25164_ (.A0(net812),
    .A1(\cpu.icache.r_data[6][18] ),
    .S(_06480_),
    .X(_02212_));
 sg13g2_mux2_1 _25165_ (.A0(net811),
    .A1(\cpu.icache.r_data[6][19] ),
    .S(_06480_),
    .X(_02213_));
 sg13g2_mux2_1 _25166_ (.A0(net810),
    .A1(\cpu.icache.r_data[6][1] ),
    .S(_06477_),
    .X(_02214_));
 sg13g2_nand2_2 _25167_ (.Y(_06481_),
    .A(net544),
    .B(_06381_));
 sg13g2_mux2_1 _25168_ (.A0(net813),
    .A1(\cpu.icache.r_data[6][20] ),
    .S(_06481_),
    .X(_02215_));
 sg13g2_mux2_1 _25169_ (.A0(net810),
    .A1(\cpu.icache.r_data[6][21] ),
    .S(_06481_),
    .X(_02216_));
 sg13g2_mux2_1 _25170_ (.A0(net812),
    .A1(\cpu.icache.r_data[6][22] ),
    .S(_06481_),
    .X(_02217_));
 sg13g2_mux2_1 _25171_ (.A0(net811),
    .A1(\cpu.icache.r_data[6][23] ),
    .S(_06481_),
    .X(_02218_));
 sg13g2_nand2_1 _25172_ (.Y(_06482_),
    .A(_08922_),
    .B(_06385_));
 sg13g2_buf_2 _25173_ (.A(_06482_),
    .X(_06483_));
 sg13g2_mux2_1 _25174_ (.A0(net813),
    .A1(\cpu.icache.r_data[6][24] ),
    .S(_06483_),
    .X(_02219_));
 sg13g2_mux2_1 _25175_ (.A0(_06404_),
    .A1(\cpu.icache.r_data[6][25] ),
    .S(_06483_),
    .X(_02220_));
 sg13g2_mux2_1 _25176_ (.A0(net812),
    .A1(\cpu.icache.r_data[6][26] ),
    .S(_06483_),
    .X(_02221_));
 sg13g2_mux2_1 _25177_ (.A0(net811),
    .A1(\cpu.icache.r_data[6][27] ),
    .S(_06483_),
    .X(_02222_));
 sg13g2_nand2_2 _25178_ (.Y(_06484_),
    .A(net544),
    .B(_06390_));
 sg13g2_mux2_1 _25179_ (.A0(net813),
    .A1(\cpu.icache.r_data[6][28] ),
    .S(_06484_),
    .X(_02223_));
 sg13g2_mux2_1 _25180_ (.A0(net810),
    .A1(\cpu.icache.r_data[6][29] ),
    .S(_06484_),
    .X(_02224_));
 sg13g2_mux2_1 _25181_ (.A0(net812),
    .A1(\cpu.icache.r_data[6][2] ),
    .S(_06477_),
    .X(_02225_));
 sg13g2_mux2_1 _25182_ (.A0(_06398_),
    .A1(\cpu.icache.r_data[6][30] ),
    .S(_06484_),
    .X(_02226_));
 sg13g2_mux2_1 _25183_ (.A0(net811),
    .A1(\cpu.icache.r_data[6][31] ),
    .S(_06484_),
    .X(_02227_));
 sg13g2_mux2_1 _25184_ (.A0(net811),
    .A1(\cpu.icache.r_data[6][3] ),
    .S(_06477_),
    .X(_02228_));
 sg13g2_nand2_2 _25185_ (.Y(_06485_),
    .A(_08922_),
    .B(_06393_));
 sg13g2_mux2_1 _25186_ (.A0(_06395_),
    .A1(\cpu.icache.r_data[6][4] ),
    .S(_06485_),
    .X(_02229_));
 sg13g2_mux2_1 _25187_ (.A0(net810),
    .A1(\cpu.icache.r_data[6][5] ),
    .S(_06485_),
    .X(_02230_));
 sg13g2_mux2_1 _25188_ (.A0(_06398_),
    .A1(\cpu.icache.r_data[6][6] ),
    .S(_06485_),
    .X(_02231_));
 sg13g2_mux2_1 _25189_ (.A0(_06401_),
    .A1(\cpu.icache.r_data[6][7] ),
    .S(_06485_),
    .X(_02232_));
 sg13g2_mux2_1 _25190_ (.A0(_06395_),
    .A1(\cpu.icache.r_data[6][8] ),
    .S(_06478_),
    .X(_02233_));
 sg13g2_mux2_1 _25191_ (.A0(_06404_),
    .A1(\cpu.icache.r_data[6][9] ),
    .S(_06478_),
    .X(_02234_));
 sg13g2_and2_1 _25192_ (.A(net543),
    .B(_06362_),
    .X(_06486_));
 sg13g2_buf_1 _25193_ (.A(_06486_),
    .X(_06487_));
 sg13g2_mux2_1 _25194_ (.A0(\cpu.icache.r_data[7][0] ),
    .A1(net942),
    .S(_06487_),
    .X(_02235_));
 sg13g2_and2_1 _25195_ (.A(net543),
    .B(_06369_),
    .X(_06488_));
 sg13g2_buf_1 _25196_ (.A(_06488_),
    .X(_06489_));
 sg13g2_mux2_1 _25197_ (.A0(\cpu.icache.r_data[7][10] ),
    .A1(net941),
    .S(_06489_),
    .X(_02236_));
 sg13g2_mux2_1 _25198_ (.A0(\cpu.icache.r_data[7][11] ),
    .A1(_06436_),
    .S(_06489_),
    .X(_02237_));
 sg13g2_and2_1 _25199_ (.A(net543),
    .B(_06374_),
    .X(_06490_));
 sg13g2_buf_1 _25200_ (.A(_06490_),
    .X(_06491_));
 sg13g2_mux2_1 _25201_ (.A0(\cpu.icache.r_data[7][12] ),
    .A1(_06431_),
    .S(_06491_),
    .X(_02238_));
 sg13g2_mux2_1 _25202_ (.A0(\cpu.icache.r_data[7][13] ),
    .A1(net808),
    .S(_06491_),
    .X(_02239_));
 sg13g2_mux2_1 _25203_ (.A0(\cpu.icache.r_data[7][14] ),
    .A1(net941),
    .S(_06491_),
    .X(_02240_));
 sg13g2_mux2_1 _25204_ (.A0(\cpu.icache.r_data[7][15] ),
    .A1(net940),
    .S(_06491_),
    .X(_02241_));
 sg13g2_and2_1 _25205_ (.A(net543),
    .B(_06378_),
    .X(_06492_));
 sg13g2_buf_1 _25206_ (.A(_06492_),
    .X(_06493_));
 sg13g2_mux2_1 _25207_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(_06431_),
    .S(_06493_),
    .X(_02242_));
 sg13g2_mux2_1 _25208_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(_06434_),
    .S(_06493_),
    .X(_02243_));
 sg13g2_mux2_1 _25209_ (.A0(\cpu.icache.r_data[7][18] ),
    .A1(_06435_),
    .S(_06493_),
    .X(_02244_));
 sg13g2_mux2_1 _25210_ (.A0(\cpu.icache.r_data[7][19] ),
    .A1(net940),
    .S(_06493_),
    .X(_02245_));
 sg13g2_mux2_1 _25211_ (.A0(\cpu.icache.r_data[7][1] ),
    .A1(_06434_),
    .S(_06487_),
    .X(_02246_));
 sg13g2_and2_1 _25212_ (.A(net543),
    .B(_06381_),
    .X(_06494_));
 sg13g2_buf_1 _25213_ (.A(_06494_),
    .X(_06495_));
 sg13g2_mux2_1 _25214_ (.A0(\cpu.icache.r_data[7][20] ),
    .A1(net942),
    .S(_06495_),
    .X(_02247_));
 sg13g2_mux2_1 _25215_ (.A0(\cpu.icache.r_data[7][21] ),
    .A1(net808),
    .S(_06495_),
    .X(_02248_));
 sg13g2_mux2_1 _25216_ (.A0(\cpu.icache.r_data[7][22] ),
    .A1(net941),
    .S(_06495_),
    .X(_02249_));
 sg13g2_mux2_1 _25217_ (.A0(\cpu.icache.r_data[7][23] ),
    .A1(net940),
    .S(_06495_),
    .X(_02250_));
 sg13g2_and2_1 _25218_ (.A(net543),
    .B(_06385_),
    .X(_06496_));
 sg13g2_buf_2 _25219_ (.A(_06496_),
    .X(_06497_));
 sg13g2_mux2_1 _25220_ (.A0(\cpu.icache.r_data[7][24] ),
    .A1(net1000),
    .S(_06497_),
    .X(_02251_));
 sg13g2_mux2_1 _25221_ (.A0(\cpu.icache.r_data[7][25] ),
    .A1(net991),
    .S(_06497_),
    .X(_02252_));
 sg13g2_mux2_1 _25222_ (.A0(\cpu.icache.r_data[7][26] ),
    .A1(net996),
    .S(_06497_),
    .X(_02253_));
 sg13g2_mux2_1 _25223_ (.A0(\cpu.icache.r_data[7][27] ),
    .A1(net995),
    .S(_06497_),
    .X(_02254_));
 sg13g2_and2_1 _25224_ (.A(_08947_),
    .B(_06390_),
    .X(_06498_));
 sg13g2_buf_1 _25225_ (.A(_06498_),
    .X(_06499_));
 sg13g2_mux2_1 _25226_ (.A0(\cpu.icache.r_data[7][28] ),
    .A1(net1000),
    .S(_06499_),
    .X(_02255_));
 sg13g2_mux2_1 _25227_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(net991),
    .S(_06499_),
    .X(_02256_));
 sg13g2_mux2_1 _25228_ (.A0(\cpu.icache.r_data[7][2] ),
    .A1(net996),
    .S(_06487_),
    .X(_02257_));
 sg13g2_mux2_1 _25229_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(_12046_),
    .S(_06499_),
    .X(_02258_));
 sg13g2_mux2_1 _25230_ (.A0(\cpu.icache.r_data[7][31] ),
    .A1(net995),
    .S(_06499_),
    .X(_02259_));
 sg13g2_mux2_1 _25231_ (.A0(\cpu.icache.r_data[7][3] ),
    .A1(_12063_),
    .S(_06487_),
    .X(_02260_));
 sg13g2_and2_1 _25232_ (.A(net543),
    .B(_06393_),
    .X(_06500_));
 sg13g2_buf_2 _25233_ (.A(_06500_),
    .X(_06501_));
 sg13g2_mux2_1 _25234_ (.A0(\cpu.icache.r_data[7][4] ),
    .A1(_12023_),
    .S(_06501_),
    .X(_02261_));
 sg13g2_mux2_1 _25235_ (.A0(\cpu.icache.r_data[7][5] ),
    .A1(_12133_),
    .S(_06501_),
    .X(_02262_));
 sg13g2_mux2_1 _25236_ (.A0(\cpu.icache.r_data[7][6] ),
    .A1(_12046_),
    .S(_06501_),
    .X(_02263_));
 sg13g2_mux2_1 _25237_ (.A0(\cpu.icache.r_data[7][7] ),
    .A1(_12063_),
    .S(_06501_),
    .X(_02264_));
 sg13g2_mux2_1 _25238_ (.A0(\cpu.icache.r_data[7][8] ),
    .A1(_12023_),
    .S(_06489_),
    .X(_02265_));
 sg13g2_mux2_1 _25239_ (.A0(\cpu.icache.r_data[7][9] ),
    .A1(_12133_),
    .S(_06489_),
    .X(_02266_));
 sg13g2_buf_1 _25240_ (.A(_06387_),
    .X(_06502_));
 sg13g2_mux2_1 _25241_ (.A0(net964),
    .A1(\cpu.icache.r_tag[0][5] ),
    .S(net386),
    .X(_02270_));
 sg13g2_buf_1 _25242_ (.A(_06387_),
    .X(_06503_));
 sg13g2_buf_1 _25243_ (.A(net385),
    .X(_06504_));
 sg13g2_nand2_1 _25244_ (.Y(_06505_),
    .A(\cpu.icache.r_tag[0][15] ),
    .B(net386));
 sg13g2_o21ai_1 _25245_ (.B1(_06505_),
    .Y(_02271_),
    .A1(net474),
    .A2(net353));
 sg13g2_nand2_1 _25246_ (.Y(_06506_),
    .A(\cpu.icache.r_tag[0][16] ),
    .B(net386));
 sg13g2_o21ai_1 _25247_ (.B1(_06506_),
    .Y(_02272_),
    .A1(net421),
    .A2(net353));
 sg13g2_nand2_1 _25248_ (.Y(_06507_),
    .A(\cpu.icache.r_tag[0][17] ),
    .B(_06502_));
 sg13g2_o21ai_1 _25249_ (.B1(_06507_),
    .Y(_02273_),
    .A1(net475),
    .A2(_06504_));
 sg13g2_nand2_1 _25250_ (.Y(_06508_),
    .A(\cpu.icache.r_tag[0][18] ),
    .B(net386));
 sg13g2_o21ai_1 _25251_ (.B1(_06508_),
    .Y(_02274_),
    .A1(net423),
    .A2(net353));
 sg13g2_nand2_1 _25252_ (.Y(_06509_),
    .A(\cpu.icache.r_tag[0][19] ),
    .B(net386));
 sg13g2_o21ai_1 _25253_ (.B1(_06509_),
    .Y(_02275_),
    .A1(net424),
    .A2(net353));
 sg13g2_nand2_1 _25254_ (.Y(_06510_),
    .A(\cpu.icache.r_tag[0][20] ),
    .B(_06502_));
 sg13g2_o21ai_1 _25255_ (.B1(_06510_),
    .Y(_02276_),
    .A1(net479),
    .A2(net353));
 sg13g2_nand2_1 _25256_ (.Y(_06511_),
    .A(\cpu.icache.r_tag[0][21] ),
    .B(net385));
 sg13g2_o21ai_1 _25257_ (.B1(_06511_),
    .Y(_02277_),
    .A1(net422),
    .A2(net353));
 sg13g2_nand2_1 _25258_ (.Y(_06512_),
    .A(\cpu.icache.r_tag[0][22] ),
    .B(net385));
 sg13g2_o21ai_1 _25259_ (.B1(_06512_),
    .Y(_02278_),
    .A1(net420),
    .A2(_06504_));
 sg13g2_nand2_1 _25260_ (.Y(_06513_),
    .A(\cpu.icache.r_tag[0][23] ),
    .B(net385));
 sg13g2_o21ai_1 _25261_ (.B1(_06513_),
    .Y(_02279_),
    .A1(net477),
    .A2(net353));
 sg13g2_mux2_1 _25262_ (.A0(net963),
    .A1(\cpu.icache.r_tag[0][6] ),
    .S(net386),
    .X(_02280_));
 sg13g2_mux2_1 _25263_ (.A0(net962),
    .A1(\cpu.icache.r_tag[0][7] ),
    .S(net386),
    .X(_02281_));
 sg13g2_nand2_1 _25264_ (.Y(_06514_),
    .A(\cpu.icache.r_tag[0][8] ),
    .B(_06503_));
 sg13g2_o21ai_1 _25265_ (.B1(_06514_),
    .Y(_02282_),
    .A1(net1050),
    .A2(net387));
 sg13g2_nand2_1 _25266_ (.Y(_06515_),
    .A(\cpu.icache.r_tag[0][9] ),
    .B(_06503_));
 sg13g2_o21ai_1 _25267_ (.B1(_06515_),
    .Y(_02283_),
    .A1(net906),
    .A2(net387));
 sg13g2_mux2_1 _25268_ (.A0(net961),
    .A1(\cpu.icache.r_tag[0][10] ),
    .S(net386),
    .X(_02284_));
 sg13g2_nand2_1 _25269_ (.Y(_06516_),
    .A(\cpu.icache.r_tag[0][11] ),
    .B(net385));
 sg13g2_o21ai_1 _25270_ (.B1(_06516_),
    .Y(_02285_),
    .A1(net1051),
    .A2(net387));
 sg13g2_nand2_1 _25271_ (.Y(_06517_),
    .A(\cpu.icache.r_tag[0][12] ),
    .B(net385));
 sg13g2_o21ai_1 _25272_ (.B1(_06517_),
    .Y(_02286_),
    .A1(net384),
    .A2(net387));
 sg13g2_nand2_1 _25273_ (.Y(_06518_),
    .A(\cpu.icache.r_tag[0][13] ),
    .B(net385));
 sg13g2_o21ai_1 _25274_ (.B1(_06518_),
    .Y(_02287_),
    .A1(net383),
    .A2(_06388_));
 sg13g2_nand2_1 _25275_ (.Y(_06519_),
    .A(\cpu.icache.r_tag[0][14] ),
    .B(net385));
 sg13g2_o21ai_1 _25276_ (.B1(_06519_),
    .Y(_02288_),
    .A1(net476),
    .A2(_06388_));
 sg13g2_nor3_1 _25277_ (.A(_06357_),
    .B(_06365_),
    .C(_06367_),
    .Y(_06520_));
 sg13g2_buf_1 _25278_ (.A(_06520_),
    .X(_06521_));
 sg13g2_nand2_1 _25279_ (.Y(_06522_),
    .A(net546),
    .B(_06521_));
 sg13g2_buf_1 _25280_ (.A(_06522_),
    .X(_06523_));
 sg13g2_buf_1 _25281_ (.A(_06523_),
    .X(_06524_));
 sg13g2_mux2_1 _25282_ (.A0(net964),
    .A1(\cpu.icache.r_tag[1][5] ),
    .S(net352),
    .X(_02289_));
 sg13g2_buf_1 _25283_ (.A(_06523_),
    .X(_06525_));
 sg13g2_nand2_1 _25284_ (.Y(_06526_),
    .A(\cpu.icache.r_tag[1][15] ),
    .B(net352));
 sg13g2_o21ai_1 _25285_ (.B1(_06526_),
    .Y(_02290_),
    .A1(net474),
    .A2(_06525_));
 sg13g2_buf_1 _25286_ (.A(_06523_),
    .X(_06527_));
 sg13g2_nand2_1 _25287_ (.Y(_06528_),
    .A(\cpu.icache.r_tag[1][16] ),
    .B(net350));
 sg13g2_o21ai_1 _25288_ (.B1(_06528_),
    .Y(_02291_),
    .A1(net421),
    .A2(net351));
 sg13g2_nand2_1 _25289_ (.Y(_06529_),
    .A(\cpu.icache.r_tag[1][17] ),
    .B(net350));
 sg13g2_o21ai_1 _25290_ (.B1(_06529_),
    .Y(_02292_),
    .A1(net475),
    .A2(net351));
 sg13g2_nand2_1 _25291_ (.Y(_06530_),
    .A(\cpu.icache.r_tag[1][18] ),
    .B(net350));
 sg13g2_o21ai_1 _25292_ (.B1(_06530_),
    .Y(_02293_),
    .A1(net423),
    .A2(net351));
 sg13g2_nand2_1 _25293_ (.Y(_06531_),
    .A(\cpu.icache.r_tag[1][19] ),
    .B(net350));
 sg13g2_o21ai_1 _25294_ (.B1(_06531_),
    .Y(_02294_),
    .A1(net424),
    .A2(net351));
 sg13g2_nand2_1 _25295_ (.Y(_06532_),
    .A(\cpu.icache.r_tag[1][20] ),
    .B(net350));
 sg13g2_o21ai_1 _25296_ (.B1(_06532_),
    .Y(_02295_),
    .A1(net479),
    .A2(net351));
 sg13g2_nand2_1 _25297_ (.Y(_06533_),
    .A(\cpu.icache.r_tag[1][21] ),
    .B(net350));
 sg13g2_o21ai_1 _25298_ (.B1(_06533_),
    .Y(_02296_),
    .A1(net422),
    .A2(net351));
 sg13g2_nand2_1 _25299_ (.Y(_06534_),
    .A(\cpu.icache.r_tag[1][22] ),
    .B(net350));
 sg13g2_o21ai_1 _25300_ (.B1(_06534_),
    .Y(_02297_),
    .A1(net420),
    .A2(net351));
 sg13g2_nand2_1 _25301_ (.Y(_06535_),
    .A(\cpu.icache.r_tag[1][23] ),
    .B(_06527_));
 sg13g2_o21ai_1 _25302_ (.B1(_06535_),
    .Y(_02298_),
    .A1(_08758_),
    .A2(net351));
 sg13g2_mux2_1 _25303_ (.A0(net963),
    .A1(\cpu.icache.r_tag[1][6] ),
    .S(net352),
    .X(_02299_));
 sg13g2_mux2_1 _25304_ (.A0(net962),
    .A1(\cpu.icache.r_tag[1][7] ),
    .S(_06524_),
    .X(_02300_));
 sg13g2_nand2_1 _25305_ (.Y(_06536_),
    .A(\cpu.icache.r_tag[1][8] ),
    .B(net350));
 sg13g2_o21ai_1 _25306_ (.B1(_06536_),
    .Y(_02301_),
    .A1(net1050),
    .A2(_06525_));
 sg13g2_nand2_1 _25307_ (.Y(_06537_),
    .A(\cpu.icache.r_tag[1][9] ),
    .B(_06527_));
 sg13g2_o21ai_1 _25308_ (.B1(_06537_),
    .Y(_02302_),
    .A1(net906),
    .A2(net352));
 sg13g2_mux2_1 _25309_ (.A0(net961),
    .A1(\cpu.icache.r_tag[1][10] ),
    .S(_06524_),
    .X(_02303_));
 sg13g2_nand2_1 _25310_ (.Y(_06538_),
    .A(\cpu.icache.r_tag[1][11] ),
    .B(_06523_));
 sg13g2_o21ai_1 _25311_ (.B1(_06538_),
    .Y(_02304_),
    .A1(net1051),
    .A2(net352));
 sg13g2_nand2_1 _25312_ (.Y(_06539_),
    .A(\cpu.icache.r_tag[1][12] ),
    .B(_06523_));
 sg13g2_o21ai_1 _25313_ (.B1(_06539_),
    .Y(_02305_),
    .A1(net384),
    .A2(net352));
 sg13g2_nand2_1 _25314_ (.Y(_06540_),
    .A(\cpu.icache.r_tag[1][13] ),
    .B(_06523_));
 sg13g2_o21ai_1 _25315_ (.B1(_06540_),
    .Y(_02306_),
    .A1(net383),
    .A2(net352));
 sg13g2_nand2_1 _25316_ (.Y(_06541_),
    .A(\cpu.icache.r_tag[1][14] ),
    .B(_06523_));
 sg13g2_o21ai_1 _25317_ (.B1(_06541_),
    .Y(_02307_),
    .A1(net476),
    .A2(net352));
 sg13g2_nand2_1 _25318_ (.Y(_06542_),
    .A(net480),
    .B(_06521_));
 sg13g2_buf_1 _25319_ (.A(_06542_),
    .X(_06543_));
 sg13g2_buf_1 _25320_ (.A(_06543_),
    .X(_06544_));
 sg13g2_mux2_1 _25321_ (.A0(net964),
    .A1(\cpu.icache.r_tag[2][5] ),
    .S(net298),
    .X(_02308_));
 sg13g2_buf_1 _25322_ (.A(_06543_),
    .X(_06545_));
 sg13g2_nand2_1 _25323_ (.Y(_06546_),
    .A(\cpu.icache.r_tag[2][15] ),
    .B(net298));
 sg13g2_o21ai_1 _25324_ (.B1(_06546_),
    .Y(_02309_),
    .A1(net474),
    .A2(net297));
 sg13g2_buf_1 _25325_ (.A(_06543_),
    .X(_06547_));
 sg13g2_nand2_1 _25326_ (.Y(_06548_),
    .A(\cpu.icache.r_tag[2][16] ),
    .B(net296));
 sg13g2_o21ai_1 _25327_ (.B1(_06548_),
    .Y(_02310_),
    .A1(_08944_),
    .A2(net297));
 sg13g2_nand2_1 _25328_ (.Y(_06549_),
    .A(\cpu.icache.r_tag[2][17] ),
    .B(net296));
 sg13g2_o21ai_1 _25329_ (.B1(_06549_),
    .Y(_02311_),
    .A1(net475),
    .A2(net297));
 sg13g2_nand2_1 _25330_ (.Y(_06550_),
    .A(\cpu.icache.r_tag[2][18] ),
    .B(net296));
 sg13g2_o21ai_1 _25331_ (.B1(_06550_),
    .Y(_02312_),
    .A1(net423),
    .A2(net297));
 sg13g2_nand2_1 _25332_ (.Y(_06551_),
    .A(\cpu.icache.r_tag[2][19] ),
    .B(net296));
 sg13g2_o21ai_1 _25333_ (.B1(_06551_),
    .Y(_02313_),
    .A1(net424),
    .A2(net297));
 sg13g2_nand2_1 _25334_ (.Y(_06552_),
    .A(\cpu.icache.r_tag[2][20] ),
    .B(net296));
 sg13g2_o21ai_1 _25335_ (.B1(_06552_),
    .Y(_02314_),
    .A1(net479),
    .A2(_06545_));
 sg13g2_nand2_1 _25336_ (.Y(_06553_),
    .A(\cpu.icache.r_tag[2][21] ),
    .B(net296));
 sg13g2_o21ai_1 _25337_ (.B1(_06553_),
    .Y(_02315_),
    .A1(net422),
    .A2(net297));
 sg13g2_nand2_1 _25338_ (.Y(_06554_),
    .A(\cpu.icache.r_tag[2][22] ),
    .B(net296));
 sg13g2_o21ai_1 _25339_ (.B1(_06554_),
    .Y(_02316_),
    .A1(net420),
    .A2(_06545_));
 sg13g2_nand2_1 _25340_ (.Y(_06555_),
    .A(\cpu.icache.r_tag[2][23] ),
    .B(net296));
 sg13g2_o21ai_1 _25341_ (.B1(_06555_),
    .Y(_02317_),
    .A1(net477),
    .A2(net297));
 sg13g2_mux2_1 _25342_ (.A0(net963),
    .A1(\cpu.icache.r_tag[2][6] ),
    .S(net298),
    .X(_02318_));
 sg13g2_mux2_1 _25343_ (.A0(net962),
    .A1(\cpu.icache.r_tag[2][7] ),
    .S(_06544_),
    .X(_02319_));
 sg13g2_nand2_1 _25344_ (.Y(_06556_),
    .A(\cpu.icache.r_tag[2][8] ),
    .B(_06547_));
 sg13g2_o21ai_1 _25345_ (.B1(_06556_),
    .Y(_02320_),
    .A1(net1050),
    .A2(net297));
 sg13g2_nand2_1 _25346_ (.Y(_06557_),
    .A(\cpu.icache.r_tag[2][9] ),
    .B(_06547_));
 sg13g2_o21ai_1 _25347_ (.B1(_06557_),
    .Y(_02321_),
    .A1(net906),
    .A2(net298));
 sg13g2_mux2_1 _25348_ (.A0(net961),
    .A1(\cpu.icache.r_tag[2][10] ),
    .S(_06544_),
    .X(_02322_));
 sg13g2_nand2_1 _25349_ (.Y(_06558_),
    .A(\cpu.icache.r_tag[2][11] ),
    .B(_06543_));
 sg13g2_o21ai_1 _25350_ (.B1(_06558_),
    .Y(_02323_),
    .A1(net1051),
    .A2(net298));
 sg13g2_nand2_1 _25351_ (.Y(_06559_),
    .A(\cpu.icache.r_tag[2][12] ),
    .B(_06543_));
 sg13g2_o21ai_1 _25352_ (.B1(_06559_),
    .Y(_02324_),
    .A1(net384),
    .A2(net298));
 sg13g2_nand2_1 _25353_ (.Y(_06560_),
    .A(\cpu.icache.r_tag[2][13] ),
    .B(_06543_));
 sg13g2_o21ai_1 _25354_ (.B1(_06560_),
    .Y(_02325_),
    .A1(net383),
    .A2(net298));
 sg13g2_nand2_1 _25355_ (.Y(_06561_),
    .A(\cpu.icache.r_tag[2][14] ),
    .B(_06543_));
 sg13g2_o21ai_1 _25356_ (.B1(_06561_),
    .Y(_02326_),
    .A1(net476),
    .A2(net298));
 sg13g2_buf_1 _25357_ (.A(_06450_),
    .X(_06562_));
 sg13g2_mux2_1 _25358_ (.A0(net964),
    .A1(\cpu.icache.r_tag[3][5] ),
    .S(net248),
    .X(_02327_));
 sg13g2_buf_1 _25359_ (.A(_06450_),
    .X(_06563_));
 sg13g2_buf_1 _25360_ (.A(net247),
    .X(_06564_));
 sg13g2_nand2_1 _25361_ (.Y(_06565_),
    .A(\cpu.icache.r_tag[3][15] ),
    .B(net248));
 sg13g2_o21ai_1 _25362_ (.B1(_06565_),
    .Y(_02328_),
    .A1(net474),
    .A2(_06564_));
 sg13g2_nand2_1 _25363_ (.Y(_06566_),
    .A(\cpu.icache.r_tag[3][16] ),
    .B(net248));
 sg13g2_o21ai_1 _25364_ (.B1(_06566_),
    .Y(_02329_),
    .A1(net421),
    .A2(net224));
 sg13g2_nand2_1 _25365_ (.Y(_06567_),
    .A(\cpu.icache.r_tag[3][17] ),
    .B(net248));
 sg13g2_o21ai_1 _25366_ (.B1(_06567_),
    .Y(_02330_),
    .A1(net475),
    .A2(net224));
 sg13g2_nand2_1 _25367_ (.Y(_06568_),
    .A(\cpu.icache.r_tag[3][18] ),
    .B(net248));
 sg13g2_o21ai_1 _25368_ (.B1(_06568_),
    .Y(_02331_),
    .A1(net423),
    .A2(net224));
 sg13g2_nand2_1 _25369_ (.Y(_06569_),
    .A(\cpu.icache.r_tag[3][19] ),
    .B(net248));
 sg13g2_o21ai_1 _25370_ (.B1(_06569_),
    .Y(_02332_),
    .A1(net424),
    .A2(_06564_));
 sg13g2_nand2_1 _25371_ (.Y(_06570_),
    .A(\cpu.icache.r_tag[3][20] ),
    .B(net248));
 sg13g2_o21ai_1 _25372_ (.B1(_06570_),
    .Y(_02333_),
    .A1(net479),
    .A2(net224));
 sg13g2_nand2_1 _25373_ (.Y(_06571_),
    .A(\cpu.icache.r_tag[3][21] ),
    .B(net247));
 sg13g2_o21ai_1 _25374_ (.B1(_06571_),
    .Y(_02334_),
    .A1(net422),
    .A2(net224));
 sg13g2_nand2_1 _25375_ (.Y(_06572_),
    .A(\cpu.icache.r_tag[3][22] ),
    .B(net247));
 sg13g2_o21ai_1 _25376_ (.B1(_06572_),
    .Y(_02335_),
    .A1(net420),
    .A2(net224));
 sg13g2_nand2_1 _25377_ (.Y(_06573_),
    .A(\cpu.icache.r_tag[3][23] ),
    .B(net247));
 sg13g2_o21ai_1 _25378_ (.B1(_06573_),
    .Y(_02336_),
    .A1(net477),
    .A2(net224));
 sg13g2_mux2_1 _25379_ (.A0(net963),
    .A1(\cpu.icache.r_tag[3][6] ),
    .S(net248),
    .X(_02337_));
 sg13g2_mux2_1 _25380_ (.A0(net962),
    .A1(\cpu.icache.r_tag[3][7] ),
    .S(_06562_),
    .X(_02338_));
 sg13g2_nand2_1 _25381_ (.Y(_06574_),
    .A(\cpu.icache.r_tag[3][8] ),
    .B(_06563_));
 sg13g2_o21ai_1 _25382_ (.B1(_06574_),
    .Y(_02339_),
    .A1(net1050),
    .A2(_06451_));
 sg13g2_nand2_1 _25383_ (.Y(_06575_),
    .A(\cpu.icache.r_tag[3][9] ),
    .B(_06563_));
 sg13g2_o21ai_1 _25384_ (.B1(_06575_),
    .Y(_02340_),
    .A1(net906),
    .A2(_06451_));
 sg13g2_mux2_1 _25385_ (.A0(net961),
    .A1(\cpu.icache.r_tag[3][10] ),
    .S(_06562_),
    .X(_02341_));
 sg13g2_nand2_1 _25386_ (.Y(_06576_),
    .A(\cpu.icache.r_tag[3][11] ),
    .B(net247));
 sg13g2_o21ai_1 _25387_ (.B1(_06576_),
    .Y(_02342_),
    .A1(net1051),
    .A2(net249));
 sg13g2_nand2_1 _25388_ (.Y(_06577_),
    .A(\cpu.icache.r_tag[3][12] ),
    .B(net247));
 sg13g2_o21ai_1 _25389_ (.B1(_06577_),
    .Y(_02343_),
    .A1(net384),
    .A2(net249));
 sg13g2_nand2_1 _25390_ (.Y(_06578_),
    .A(\cpu.icache.r_tag[3][13] ),
    .B(net247));
 sg13g2_o21ai_1 _25391_ (.B1(_06578_),
    .Y(_02344_),
    .A1(net383),
    .A2(net249));
 sg13g2_nand2_1 _25392_ (.Y(_06579_),
    .A(\cpu.icache.r_tag[3][14] ),
    .B(net247));
 sg13g2_o21ai_1 _25393_ (.B1(_06579_),
    .Y(_02345_),
    .A1(net476),
    .A2(net249));
 sg13g2_nand2_1 _25394_ (.Y(_06580_),
    .A(net545),
    .B(_06521_));
 sg13g2_buf_1 _25395_ (.A(_06580_),
    .X(_06581_));
 sg13g2_buf_1 _25396_ (.A(_06581_),
    .X(_06582_));
 sg13g2_mux2_1 _25397_ (.A0(net964),
    .A1(\cpu.icache.r_tag[4][5] ),
    .S(net349),
    .X(_02346_));
 sg13g2_buf_1 _25398_ (.A(_06581_),
    .X(_06583_));
 sg13g2_nand2_1 _25399_ (.Y(_06584_),
    .A(\cpu.icache.r_tag[4][15] ),
    .B(net349));
 sg13g2_o21ai_1 _25400_ (.B1(_06584_),
    .Y(_02347_),
    .A1(net474),
    .A2(net348));
 sg13g2_buf_1 _25401_ (.A(_06581_),
    .X(_06585_));
 sg13g2_nand2_1 _25402_ (.Y(_06586_),
    .A(\cpu.icache.r_tag[4][16] ),
    .B(net347));
 sg13g2_o21ai_1 _25403_ (.B1(_06586_),
    .Y(_02348_),
    .A1(net421),
    .A2(net348));
 sg13g2_nand2_1 _25404_ (.Y(_06587_),
    .A(\cpu.icache.r_tag[4][17] ),
    .B(net347));
 sg13g2_o21ai_1 _25405_ (.B1(_06587_),
    .Y(_02349_),
    .A1(net475),
    .A2(net348));
 sg13g2_nand2_1 _25406_ (.Y(_06588_),
    .A(\cpu.icache.r_tag[4][18] ),
    .B(net347));
 sg13g2_o21ai_1 _25407_ (.B1(_06588_),
    .Y(_02350_),
    .A1(net423),
    .A2(net348));
 sg13g2_nand2_1 _25408_ (.Y(_06589_),
    .A(\cpu.icache.r_tag[4][19] ),
    .B(net347));
 sg13g2_o21ai_1 _25409_ (.B1(_06589_),
    .Y(_02351_),
    .A1(_08735_),
    .A2(net348));
 sg13g2_nand2_1 _25410_ (.Y(_06590_),
    .A(\cpu.icache.r_tag[4][20] ),
    .B(net347));
 sg13g2_o21ai_1 _25411_ (.B1(_06590_),
    .Y(_02352_),
    .A1(net479),
    .A2(net348));
 sg13g2_nand2_1 _25412_ (.Y(_06591_),
    .A(\cpu.icache.r_tag[4][21] ),
    .B(net347));
 sg13g2_o21ai_1 _25413_ (.B1(_06591_),
    .Y(_02353_),
    .A1(net422),
    .A2(net348));
 sg13g2_nand2_1 _25414_ (.Y(_06592_),
    .A(\cpu.icache.r_tag[4][22] ),
    .B(net347));
 sg13g2_o21ai_1 _25415_ (.B1(_06592_),
    .Y(_02354_),
    .A1(net420),
    .A2(net348));
 sg13g2_nand2_1 _25416_ (.Y(_06593_),
    .A(\cpu.icache.r_tag[4][23] ),
    .B(_06585_));
 sg13g2_o21ai_1 _25417_ (.B1(_06593_),
    .Y(_02355_),
    .A1(net477),
    .A2(_06583_));
 sg13g2_mux2_1 _25418_ (.A0(net963),
    .A1(\cpu.icache.r_tag[4][6] ),
    .S(net349),
    .X(_02356_));
 sg13g2_mux2_1 _25419_ (.A0(net962),
    .A1(\cpu.icache.r_tag[4][7] ),
    .S(net349),
    .X(_02357_));
 sg13g2_nand2_1 _25420_ (.Y(_06594_),
    .A(\cpu.icache.r_tag[4][8] ),
    .B(_06585_));
 sg13g2_o21ai_1 _25421_ (.B1(_06594_),
    .Y(_02358_),
    .A1(net1050),
    .A2(_06583_));
 sg13g2_nand2_1 _25422_ (.Y(_06595_),
    .A(\cpu.icache.r_tag[4][9] ),
    .B(net347));
 sg13g2_o21ai_1 _25423_ (.B1(_06595_),
    .Y(_02359_),
    .A1(net906),
    .A2(net349));
 sg13g2_mux2_1 _25424_ (.A0(net961),
    .A1(\cpu.icache.r_tag[4][10] ),
    .S(_06582_),
    .X(_02360_));
 sg13g2_nand2_1 _25425_ (.Y(_06596_),
    .A(\cpu.icache.r_tag[4][11] ),
    .B(_06581_));
 sg13g2_o21ai_1 _25426_ (.B1(_06596_),
    .Y(_02361_),
    .A1(net1051),
    .A2(_06582_));
 sg13g2_nand2_1 _25427_ (.Y(_06597_),
    .A(\cpu.icache.r_tag[4][12] ),
    .B(_06581_));
 sg13g2_o21ai_1 _25428_ (.B1(_06597_),
    .Y(_02362_),
    .A1(net384),
    .A2(net349));
 sg13g2_nand2_1 _25429_ (.Y(_06598_),
    .A(\cpu.icache.r_tag[4][13] ),
    .B(_06581_));
 sg13g2_o21ai_1 _25430_ (.B1(_06598_),
    .Y(_02363_),
    .A1(net383),
    .A2(net349));
 sg13g2_nand2_1 _25431_ (.Y(_06599_),
    .A(\cpu.icache.r_tag[4][14] ),
    .B(_06581_));
 sg13g2_o21ai_1 _25432_ (.B1(_06599_),
    .Y(_02364_),
    .A1(net476),
    .A2(net349));
 sg13g2_nand2_1 _25433_ (.Y(_06600_),
    .A(_09078_),
    .B(_06521_));
 sg13g2_buf_1 _25434_ (.A(_06600_),
    .X(_06601_));
 sg13g2_buf_1 _25435_ (.A(_06601_),
    .X(_06602_));
 sg13g2_mux2_1 _25436_ (.A0(net964),
    .A1(\cpu.icache.r_tag[5][5] ),
    .S(net346),
    .X(_02365_));
 sg13g2_buf_1 _25437_ (.A(_06601_),
    .X(_06603_));
 sg13g2_nand2_1 _25438_ (.Y(_06604_),
    .A(\cpu.icache.r_tag[5][15] ),
    .B(net346));
 sg13g2_o21ai_1 _25439_ (.B1(_06604_),
    .Y(_02366_),
    .A1(net474),
    .A2(net345));
 sg13g2_buf_1 _25440_ (.A(_06601_),
    .X(_06605_));
 sg13g2_nand2_1 _25441_ (.Y(_06606_),
    .A(\cpu.icache.r_tag[5][16] ),
    .B(net344));
 sg13g2_o21ai_1 _25442_ (.B1(_06606_),
    .Y(_02367_),
    .A1(net421),
    .A2(net345));
 sg13g2_nand2_1 _25443_ (.Y(_06607_),
    .A(\cpu.icache.r_tag[5][17] ),
    .B(net344));
 sg13g2_o21ai_1 _25444_ (.B1(_06607_),
    .Y(_02368_),
    .A1(net475),
    .A2(net345));
 sg13g2_nand2_1 _25445_ (.Y(_06608_),
    .A(\cpu.icache.r_tag[5][18] ),
    .B(net344));
 sg13g2_o21ai_1 _25446_ (.B1(_06608_),
    .Y(_02369_),
    .A1(net423),
    .A2(net345));
 sg13g2_nand2_1 _25447_ (.Y(_06609_),
    .A(\cpu.icache.r_tag[5][19] ),
    .B(net344));
 sg13g2_o21ai_1 _25448_ (.B1(_06609_),
    .Y(_02370_),
    .A1(net424),
    .A2(net345));
 sg13g2_nand2_1 _25449_ (.Y(_06610_),
    .A(\cpu.icache.r_tag[5][20] ),
    .B(_06605_));
 sg13g2_o21ai_1 _25450_ (.B1(_06610_),
    .Y(_02371_),
    .A1(net479),
    .A2(_06603_));
 sg13g2_nand2_1 _25451_ (.Y(_06611_),
    .A(\cpu.icache.r_tag[5][21] ),
    .B(net344));
 sg13g2_o21ai_1 _25452_ (.B1(_06611_),
    .Y(_02372_),
    .A1(net422),
    .A2(net345));
 sg13g2_nand2_1 _25453_ (.Y(_06612_),
    .A(\cpu.icache.r_tag[5][22] ),
    .B(_06605_));
 sg13g2_o21ai_1 _25454_ (.B1(_06612_),
    .Y(_02373_),
    .A1(net420),
    .A2(_06603_));
 sg13g2_nand2_1 _25455_ (.Y(_06613_),
    .A(\cpu.icache.r_tag[5][23] ),
    .B(net344));
 sg13g2_o21ai_1 _25456_ (.B1(_06613_),
    .Y(_02374_),
    .A1(net477),
    .A2(net345));
 sg13g2_mux2_1 _25457_ (.A0(net963),
    .A1(\cpu.icache.r_tag[5][6] ),
    .S(net346),
    .X(_02375_));
 sg13g2_mux2_1 _25458_ (.A0(net962),
    .A1(\cpu.icache.r_tag[5][7] ),
    .S(_06602_),
    .X(_02376_));
 sg13g2_nand2_1 _25459_ (.Y(_06614_),
    .A(\cpu.icache.r_tag[5][8] ),
    .B(net344));
 sg13g2_o21ai_1 _25460_ (.B1(_06614_),
    .Y(_02377_),
    .A1(net1050),
    .A2(net345));
 sg13g2_nand2_1 _25461_ (.Y(_06615_),
    .A(\cpu.icache.r_tag[5][9] ),
    .B(net344));
 sg13g2_o21ai_1 _25462_ (.B1(_06615_),
    .Y(_02378_),
    .A1(net906),
    .A2(net346));
 sg13g2_mux2_1 _25463_ (.A0(net961),
    .A1(\cpu.icache.r_tag[5][10] ),
    .S(_06602_),
    .X(_02379_));
 sg13g2_nand2_1 _25464_ (.Y(_06616_),
    .A(\cpu.icache.r_tag[5][11] ),
    .B(_06601_));
 sg13g2_o21ai_1 _25465_ (.B1(_06616_),
    .Y(_02380_),
    .A1(net1051),
    .A2(net346));
 sg13g2_nand2_1 _25466_ (.Y(_06617_),
    .A(\cpu.icache.r_tag[5][12] ),
    .B(_06601_));
 sg13g2_o21ai_1 _25467_ (.B1(_06617_),
    .Y(_02381_),
    .A1(net384),
    .A2(net346));
 sg13g2_nand2_1 _25468_ (.Y(_06618_),
    .A(\cpu.icache.r_tag[5][13] ),
    .B(_06601_));
 sg13g2_o21ai_1 _25469_ (.B1(_06618_),
    .Y(_02382_),
    .A1(net383),
    .A2(net346));
 sg13g2_nand2_1 _25470_ (.Y(_06619_),
    .A(\cpu.icache.r_tag[5][14] ),
    .B(_06601_));
 sg13g2_o21ai_1 _25471_ (.B1(_06619_),
    .Y(_02383_),
    .A1(net476),
    .A2(net346));
 sg13g2_nand2_1 _25472_ (.Y(_06620_),
    .A(net544),
    .B(_06521_));
 sg13g2_buf_1 _25473_ (.A(_06620_),
    .X(_06621_));
 sg13g2_buf_1 _25474_ (.A(_06621_),
    .X(_06622_));
 sg13g2_mux2_1 _25475_ (.A0(_04644_),
    .A1(\cpu.icache.r_tag[6][5] ),
    .S(_06622_),
    .X(_02384_));
 sg13g2_buf_1 _25476_ (.A(_06621_),
    .X(_06623_));
 sg13g2_nand2_1 _25477_ (.Y(_06624_),
    .A(\cpu.icache.r_tag[6][15] ),
    .B(net343));
 sg13g2_o21ai_1 _25478_ (.B1(_06624_),
    .Y(_02385_),
    .A1(net474),
    .A2(net342));
 sg13g2_buf_1 _25479_ (.A(_06621_),
    .X(_06625_));
 sg13g2_nand2_1 _25480_ (.Y(_06626_),
    .A(\cpu.icache.r_tag[6][16] ),
    .B(net341));
 sg13g2_o21ai_1 _25481_ (.B1(_06626_),
    .Y(_02386_),
    .A1(net421),
    .A2(net342));
 sg13g2_nand2_1 _25482_ (.Y(_06627_),
    .A(\cpu.icache.r_tag[6][17] ),
    .B(net341));
 sg13g2_o21ai_1 _25483_ (.B1(_06627_),
    .Y(_02387_),
    .A1(net475),
    .A2(net342));
 sg13g2_nand2_1 _25484_ (.Y(_06628_),
    .A(\cpu.icache.r_tag[6][18] ),
    .B(net341));
 sg13g2_o21ai_1 _25485_ (.B1(_06628_),
    .Y(_02388_),
    .A1(net423),
    .A2(net342));
 sg13g2_nand2_1 _25486_ (.Y(_06629_),
    .A(\cpu.icache.r_tag[6][19] ),
    .B(_06625_));
 sg13g2_o21ai_1 _25487_ (.B1(_06629_),
    .Y(_02389_),
    .A1(net424),
    .A2(_06623_));
 sg13g2_nand2_1 _25488_ (.Y(_06630_),
    .A(\cpu.icache.r_tag[6][20] ),
    .B(_06625_));
 sg13g2_o21ai_1 _25489_ (.B1(_06630_),
    .Y(_02390_),
    .A1(net479),
    .A2(_06623_));
 sg13g2_nand2_1 _25490_ (.Y(_06631_),
    .A(\cpu.icache.r_tag[6][21] ),
    .B(net341));
 sg13g2_o21ai_1 _25491_ (.B1(_06631_),
    .Y(_02391_),
    .A1(net422),
    .A2(net342));
 sg13g2_nand2_1 _25492_ (.Y(_06632_),
    .A(\cpu.icache.r_tag[6][22] ),
    .B(net341));
 sg13g2_o21ai_1 _25493_ (.B1(_06632_),
    .Y(_02392_),
    .A1(net420),
    .A2(net342));
 sg13g2_nand2_1 _25494_ (.Y(_06633_),
    .A(\cpu.icache.r_tag[6][23] ),
    .B(net341));
 sg13g2_o21ai_1 _25495_ (.B1(_06633_),
    .Y(_02393_),
    .A1(net477),
    .A2(net342));
 sg13g2_mux2_1 _25496_ (.A0(_04675_),
    .A1(\cpu.icache.r_tag[6][6] ),
    .S(net343),
    .X(_02394_));
 sg13g2_mux2_1 _25497_ (.A0(_04704_),
    .A1(\cpu.icache.r_tag[6][7] ),
    .S(net343),
    .X(_02395_));
 sg13g2_nand2_1 _25498_ (.Y(_06634_),
    .A(\cpu.icache.r_tag[6][8] ),
    .B(net341));
 sg13g2_o21ai_1 _25499_ (.B1(_06634_),
    .Y(_02396_),
    .A1(net1050),
    .A2(net342));
 sg13g2_nand2_1 _25500_ (.Y(_06635_),
    .A(\cpu.icache.r_tag[6][9] ),
    .B(net341));
 sg13g2_o21ai_1 _25501_ (.B1(_06635_),
    .Y(_02397_),
    .A1(net906),
    .A2(net343));
 sg13g2_mux2_1 _25502_ (.A0(_04801_),
    .A1(\cpu.icache.r_tag[6][10] ),
    .S(net343),
    .X(_02398_));
 sg13g2_nand2_1 _25503_ (.Y(_06636_),
    .A(\cpu.icache.r_tag[6][11] ),
    .B(_06621_));
 sg13g2_o21ai_1 _25504_ (.B1(_06636_),
    .Y(_02399_),
    .A1(net1051),
    .A2(net343));
 sg13g2_nand2_1 _25505_ (.Y(_06637_),
    .A(\cpu.icache.r_tag[6][12] ),
    .B(_06621_));
 sg13g2_o21ai_1 _25506_ (.B1(_06637_),
    .Y(_02400_),
    .A1(net384),
    .A2(net343));
 sg13g2_nand2_1 _25507_ (.Y(_06638_),
    .A(\cpu.icache.r_tag[6][13] ),
    .B(_06621_));
 sg13g2_o21ai_1 _25508_ (.B1(_06638_),
    .Y(_02401_),
    .A1(net383),
    .A2(net343));
 sg13g2_nand2_1 _25509_ (.Y(_06639_),
    .A(\cpu.icache.r_tag[6][14] ),
    .B(_06621_));
 sg13g2_o21ai_1 _25510_ (.B1(_06639_),
    .Y(_02402_),
    .A1(net476),
    .A2(_06622_));
 sg13g2_nand2_1 _25511_ (.Y(_06640_),
    .A(net543),
    .B(_06521_));
 sg13g2_buf_1 _25512_ (.A(_06640_),
    .X(_06641_));
 sg13g2_buf_1 _25513_ (.A(_06641_),
    .X(_06642_));
 sg13g2_mux2_1 _25514_ (.A0(_04644_),
    .A1(\cpu.icache.r_tag[7][5] ),
    .S(net340),
    .X(_02403_));
 sg13g2_buf_1 _25515_ (.A(_06641_),
    .X(_06643_));
 sg13g2_nand2_1 _25516_ (.Y(_06644_),
    .A(\cpu.icache.r_tag[7][15] ),
    .B(net340));
 sg13g2_o21ai_1 _25517_ (.B1(_06644_),
    .Y(_02404_),
    .A1(_08988_),
    .A2(net339));
 sg13g2_buf_1 _25518_ (.A(_06641_),
    .X(_06645_));
 sg13g2_nand2_1 _25519_ (.Y(_06646_),
    .A(\cpu.icache.r_tag[7][16] ),
    .B(net338));
 sg13g2_o21ai_1 _25520_ (.B1(_06646_),
    .Y(_02405_),
    .A1(net421),
    .A2(net339));
 sg13g2_nand2_1 _25521_ (.Y(_06647_),
    .A(\cpu.icache.r_tag[7][17] ),
    .B(net338));
 sg13g2_o21ai_1 _25522_ (.B1(_06647_),
    .Y(_02406_),
    .A1(net475),
    .A2(net339));
 sg13g2_nand2_1 _25523_ (.Y(_06648_),
    .A(\cpu.icache.r_tag[7][18] ),
    .B(net338));
 sg13g2_o21ai_1 _25524_ (.B1(_06648_),
    .Y(_02407_),
    .A1(net423),
    .A2(net339));
 sg13g2_nand2_1 _25525_ (.Y(_06649_),
    .A(\cpu.icache.r_tag[7][19] ),
    .B(net338));
 sg13g2_o21ai_1 _25526_ (.B1(_06649_),
    .Y(_02408_),
    .A1(net424),
    .A2(net339));
 sg13g2_nand2_1 _25527_ (.Y(_06650_),
    .A(\cpu.icache.r_tag[7][20] ),
    .B(_06645_));
 sg13g2_o21ai_1 _25528_ (.B1(_06650_),
    .Y(_02409_),
    .A1(_08713_),
    .A2(_06643_));
 sg13g2_nand2_1 _25529_ (.Y(_06651_),
    .A(\cpu.icache.r_tag[7][21] ),
    .B(net338));
 sg13g2_o21ai_1 _25530_ (.B1(_06651_),
    .Y(_02410_),
    .A1(_08920_),
    .A2(net339));
 sg13g2_nand2_1 _25531_ (.Y(_06652_),
    .A(\cpu.icache.r_tag[7][22] ),
    .B(_06645_));
 sg13g2_o21ai_1 _25532_ (.B1(_06652_),
    .Y(_02411_),
    .A1(_08966_),
    .A2(net339));
 sg13g2_nand2_1 _25533_ (.Y(_06653_),
    .A(\cpu.icache.r_tag[7][23] ),
    .B(net338));
 sg13g2_o21ai_1 _25534_ (.B1(_06653_),
    .Y(_02412_),
    .A1(net477),
    .A2(net339));
 sg13g2_mux2_1 _25535_ (.A0(_04675_),
    .A1(\cpu.icache.r_tag[7][6] ),
    .S(net340),
    .X(_02413_));
 sg13g2_mux2_1 _25536_ (.A0(_04704_),
    .A1(\cpu.icache.r_tag[7][7] ),
    .S(net340),
    .X(_02414_));
 sg13g2_nand2_1 _25537_ (.Y(_06654_),
    .A(\cpu.icache.r_tag[7][8] ),
    .B(net338));
 sg13g2_o21ai_1 _25538_ (.B1(_06654_),
    .Y(_02415_),
    .A1(_08820_),
    .A2(_06643_));
 sg13g2_nand2_1 _25539_ (.Y(_06655_),
    .A(\cpu.icache.r_tag[7][9] ),
    .B(net338));
 sg13g2_o21ai_1 _25540_ (.B1(_06655_),
    .Y(_02416_),
    .A1(_08788_),
    .A2(net340));
 sg13g2_mux2_1 _25541_ (.A0(_04801_),
    .A1(\cpu.icache.r_tag[7][10] ),
    .S(net340),
    .X(_02417_));
 sg13g2_nand2_1 _25542_ (.Y(_06656_),
    .A(\cpu.icache.r_tag[7][11] ),
    .B(_06641_));
 sg13g2_o21ai_1 _25543_ (.B1(_06656_),
    .Y(_02418_),
    .A1(_08769_),
    .A2(_06642_));
 sg13g2_nand2_1 _25544_ (.Y(_06657_),
    .A(\cpu.icache.r_tag[7][12] ),
    .B(_06641_));
 sg13g2_o21ai_1 _25545_ (.B1(_06657_),
    .Y(_02419_),
    .A1(_08648_),
    .A2(net340));
 sg13g2_nand2_1 _25546_ (.Y(_06658_),
    .A(\cpu.icache.r_tag[7][13] ),
    .B(_06641_));
 sg13g2_o21ai_1 _25547_ (.B1(_06658_),
    .Y(_02420_),
    .A1(_08681_),
    .A2(net340));
 sg13g2_nand2_1 _25548_ (.Y(_06659_),
    .A(\cpu.icache.r_tag[7][14] ),
    .B(_06641_));
 sg13g2_o21ai_1 _25549_ (.B1(_06659_),
    .Y(_02421_),
    .A1(_08879_),
    .A2(_06642_));
 sg13g2_and2_1 _25550_ (.A(net171),
    .B(net499),
    .X(_06660_));
 sg13g2_buf_2 _25551_ (.A(_06660_),
    .X(_06661_));
 sg13g2_buf_1 _25552_ (.A(_06661_),
    .X(_06662_));
 sg13g2_mux2_1 _25553_ (.A0(\cpu.intr.r_clock_cmp[0] ),
    .A1(net890),
    .S(_06662_),
    .X(_02431_));
 sg13g2_mux2_1 _25554_ (.A0(\cpu.intr.r_clock_cmp[10] ),
    .A1(_10191_),
    .S(net95),
    .X(_02432_));
 sg13g2_mux2_1 _25555_ (.A0(\cpu.intr.r_clock_cmp[11] ),
    .A1(_10198_),
    .S(net95),
    .X(_02433_));
 sg13g2_mux2_1 _25556_ (.A0(\cpu.intr.r_clock_cmp[12] ),
    .A1(_10203_),
    .S(net95),
    .X(_02434_));
 sg13g2_mux2_1 _25557_ (.A0(\cpu.intr.r_clock_cmp[13] ),
    .A1(_10205_),
    .S(net95),
    .X(_02435_));
 sg13g2_mux2_1 _25558_ (.A0(\cpu.intr.r_clock_cmp[14] ),
    .A1(_10215_),
    .S(_06662_),
    .X(_02436_));
 sg13g2_mux2_1 _25559_ (.A0(\cpu.intr.r_clock_cmp[15] ),
    .A1(_10220_),
    .S(net95),
    .X(_02437_));
 sg13g2_nor2_1 _25560_ (.A(_10061_),
    .B(_04929_),
    .Y(_06663_));
 sg13g2_buf_2 _25561_ (.A(_06663_),
    .X(_06664_));
 sg13g2_buf_1 _25562_ (.A(_06664_),
    .X(_06665_));
 sg13g2_mux2_1 _25563_ (.A0(\cpu.intr.r_clock_cmp[16] ),
    .A1(net890),
    .S(net94),
    .X(_02438_));
 sg13g2_buf_1 _25564_ (.A(_10069_),
    .X(_06666_));
 sg13g2_mux2_1 _25565_ (.A0(\cpu.intr.r_clock_cmp[17] ),
    .A1(net939),
    .S(net94),
    .X(_02439_));
 sg13g2_mux2_1 _25566_ (.A0(\cpu.intr.r_clock_cmp[18] ),
    .A1(net886),
    .S(net94),
    .X(_02440_));
 sg13g2_mux2_1 _25567_ (.A0(\cpu.intr.r_clock_cmp[19] ),
    .A1(net885),
    .S(net94),
    .X(_02441_));
 sg13g2_mux2_1 _25568_ (.A0(\cpu.intr.r_clock_cmp[1] ),
    .A1(net939),
    .S(net95),
    .X(_02442_));
 sg13g2_mux2_1 _25569_ (.A0(\cpu.intr.r_clock_cmp[20] ),
    .A1(net992),
    .S(net94),
    .X(_02443_));
 sg13g2_mux2_1 _25570_ (.A0(\cpu.intr.r_clock_cmp[21] ),
    .A1(net990),
    .S(_06665_),
    .X(_02444_));
 sg13g2_mux2_1 _25571_ (.A0(\cpu.intr.r_clock_cmp[22] ),
    .A1(net989),
    .S(net94),
    .X(_02445_));
 sg13g2_mux2_1 _25572_ (.A0(\cpu.intr.r_clock_cmp[23] ),
    .A1(net851),
    .S(_06665_),
    .X(_02446_));
 sg13g2_mux2_1 _25573_ (.A0(\cpu.intr.r_clock_cmp[24] ),
    .A1(_10181_),
    .S(net94),
    .X(_02447_));
 sg13g2_mux2_1 _25574_ (.A0(\cpu.intr.r_clock_cmp[25] ),
    .A1(_10186_),
    .S(net94),
    .X(_02448_));
 sg13g2_mux2_1 _25575_ (.A0(\cpu.intr.r_clock_cmp[26] ),
    .A1(_10191_),
    .S(_06664_),
    .X(_02449_));
 sg13g2_mux2_1 _25576_ (.A0(\cpu.intr.r_clock_cmp[27] ),
    .A1(_10198_),
    .S(_06664_),
    .X(_02450_));
 sg13g2_mux2_1 _25577_ (.A0(\cpu.intr.r_clock_cmp[28] ),
    .A1(_10203_),
    .S(_06664_),
    .X(_02451_));
 sg13g2_mux2_1 _25578_ (.A0(\cpu.intr.r_clock_cmp[29] ),
    .A1(_10205_),
    .S(_06664_),
    .X(_02452_));
 sg13g2_mux2_1 _25579_ (.A0(\cpu.intr.r_clock_cmp[2] ),
    .A1(net886),
    .S(net95),
    .X(_02453_));
 sg13g2_mux2_1 _25580_ (.A0(\cpu.intr.r_clock_cmp[30] ),
    .A1(_10215_),
    .S(_06664_),
    .X(_02454_));
 sg13g2_mux2_1 _25581_ (.A0(\cpu.intr.r_clock_cmp[31] ),
    .A1(_10220_),
    .S(_06664_),
    .X(_02455_));
 sg13g2_mux2_1 _25582_ (.A0(\cpu.intr.r_clock_cmp[3] ),
    .A1(net885),
    .S(net95),
    .X(_02456_));
 sg13g2_mux2_1 _25583_ (.A0(\cpu.intr.r_clock_cmp[4] ),
    .A1(net992),
    .S(_06661_),
    .X(_02457_));
 sg13g2_mux2_1 _25584_ (.A0(\cpu.intr.r_clock_cmp[5] ),
    .A1(net990),
    .S(_06661_),
    .X(_02458_));
 sg13g2_mux2_1 _25585_ (.A0(\cpu.intr.r_clock_cmp[6] ),
    .A1(net989),
    .S(_06661_),
    .X(_02459_));
 sg13g2_mux2_1 _25586_ (.A0(\cpu.intr.r_clock_cmp[7] ),
    .A1(net851),
    .S(_06661_),
    .X(_02460_));
 sg13g2_mux2_1 _25587_ (.A0(\cpu.intr.r_clock_cmp[8] ),
    .A1(_10181_),
    .S(_06661_),
    .X(_02461_));
 sg13g2_mux2_1 _25588_ (.A0(\cpu.intr.r_clock_cmp[9] ),
    .A1(_10186_),
    .S(_06661_),
    .X(_02462_));
 sg13g2_nor3_1 _25589_ (.A(net538),
    .B(net539),
    .C(_10061_),
    .Y(_06667_));
 sg13g2_buf_2 _25590_ (.A(_06667_),
    .X(_06668_));
 sg13g2_buf_1 _25591_ (.A(_06668_),
    .X(_06669_));
 sg13g2_mux2_1 _25592_ (.A0(\cpu.intr.r_timer_reload[0] ),
    .A1(net890),
    .S(net93),
    .X(_02486_));
 sg13g2_mux2_1 _25593_ (.A0(\cpu.intr.r_timer_reload[10] ),
    .A1(_10191_),
    .S(net93),
    .X(_02487_));
 sg13g2_mux2_1 _25594_ (.A0(\cpu.intr.r_timer_reload[11] ),
    .A1(_10198_),
    .S(net93),
    .X(_02488_));
 sg13g2_mux2_1 _25595_ (.A0(\cpu.intr.r_timer_reload[12] ),
    .A1(_10203_),
    .S(net93),
    .X(_02489_));
 sg13g2_mux2_1 _25596_ (.A0(\cpu.intr.r_timer_reload[13] ),
    .A1(_10205_),
    .S(net93),
    .X(_02490_));
 sg13g2_mux2_1 _25597_ (.A0(\cpu.intr.r_timer_reload[14] ),
    .A1(_10215_),
    .S(net93),
    .X(_02491_));
 sg13g2_mux2_1 _25598_ (.A0(\cpu.intr.r_timer_reload[15] ),
    .A1(_10220_),
    .S(net93),
    .X(_02492_));
 sg13g2_mux2_1 _25599_ (.A0(\cpu.intr.r_timer_reload[16] ),
    .A1(net890),
    .S(net104),
    .X(_02493_));
 sg13g2_inv_1 _25600_ (.Y(_06670_),
    .A(\cpu.intr.r_timer_reload[17] ));
 sg13g2_o21ai_1 _25601_ (.B1(_10071_),
    .Y(_02494_),
    .A1(_06670_),
    .A2(net104));
 sg13g2_inv_1 _25602_ (.Y(_06671_),
    .A(\cpu.intr.r_timer_reload[18] ));
 sg13g2_o21ai_1 _25603_ (.B1(_10076_),
    .Y(_02495_),
    .A1(_06671_),
    .A2(net104));
 sg13g2_inv_1 _25604_ (.Y(_06672_),
    .A(\cpu.intr.r_timer_reload[19] ));
 sg13g2_o21ai_1 _25605_ (.B1(_10081_),
    .Y(_02496_),
    .A1(_06672_),
    .A2(net104));
 sg13g2_mux2_1 _25606_ (.A0(\cpu.intr.r_timer_reload[1] ),
    .A1(net939),
    .S(_06669_),
    .X(_02497_));
 sg13g2_mux2_1 _25607_ (.A0(\cpu.intr.r_timer_reload[20] ),
    .A1(net992),
    .S(net104),
    .X(_02498_));
 sg13g2_o21ai_1 _25608_ (.B1(_10093_),
    .Y(_02499_),
    .A1(_05622_),
    .A2(_10064_));
 sg13g2_inv_1 _25609_ (.Y(_06673_),
    .A(\cpu.intr.r_timer_reload[22] ));
 sg13g2_o21ai_1 _25610_ (.B1(_10099_),
    .Y(_02500_),
    .A1(_06673_),
    .A2(net104));
 sg13g2_mux2_1 _25611_ (.A0(\cpu.intr.r_timer_reload[23] ),
    .A1(net851),
    .S(_10063_),
    .X(_02501_));
 sg13g2_mux2_1 _25612_ (.A0(\cpu.intr.r_timer_reload[2] ),
    .A1(_10133_),
    .S(net93),
    .X(_02502_));
 sg13g2_mux2_1 _25613_ (.A0(\cpu.intr.r_timer_reload[3] ),
    .A1(_10146_),
    .S(_06669_),
    .X(_02503_));
 sg13g2_mux2_1 _25614_ (.A0(\cpu.intr.r_timer_reload[4] ),
    .A1(net992),
    .S(_06668_),
    .X(_02504_));
 sg13g2_mux2_1 _25615_ (.A0(\cpu.intr.r_timer_reload[5] ),
    .A1(_12136_),
    .S(_06668_),
    .X(_02505_));
 sg13g2_mux2_1 _25616_ (.A0(\cpu.intr.r_timer_reload[6] ),
    .A1(net989),
    .S(_06668_),
    .X(_02506_));
 sg13g2_mux2_1 _25617_ (.A0(\cpu.intr.r_timer_reload[7] ),
    .A1(net851),
    .S(_06668_),
    .X(_02507_));
 sg13g2_mux2_1 _25618_ (.A0(\cpu.intr.r_timer_reload[8] ),
    .A1(_10181_),
    .S(_06668_),
    .X(_02508_));
 sg13g2_mux2_1 _25619_ (.A0(\cpu.intr.r_timer_reload[9] ),
    .A1(_10186_),
    .S(_06668_),
    .X(_02509_));
 sg13g2_nand2b_1 _25620_ (.Y(_06674_),
    .B(_09869_),
    .A_N(_09830_));
 sg13g2_nor4_2 _25621_ (.A(_11914_),
    .B(_11916_),
    .C(_11917_),
    .Y(_06675_),
    .D(_11884_));
 sg13g2_nor2_1 _25622_ (.A(_09844_),
    .B(_09832_),
    .Y(_06676_));
 sg13g2_nor2_1 _25623_ (.A(_11882_),
    .B(_09854_),
    .Y(_06677_));
 sg13g2_nand4_1 _25624_ (.B(_06675_),
    .C(_06676_),
    .A(_11880_),
    .Y(_06678_),
    .D(_06677_));
 sg13g2_a21oi_1 _25625_ (.A1(_09390_),
    .A2(_06674_),
    .Y(_06679_),
    .B1(_06678_));
 sg13g2_buf_1 _25626_ (.A(_06679_),
    .X(_06680_));
 sg13g2_mux2_1 _25627_ (.A0(\cpu.qspi.r_read_delay[0][0] ),
    .A1(\cpu.qspi.r_read_delay[1][0] ),
    .S(_09863_),
    .X(_06681_));
 sg13g2_mux2_1 _25628_ (.A0(_06681_),
    .A1(\cpu.qspi.r_read_delay[2][0] ),
    .S(net245),
    .X(_06682_));
 sg13g2_or4_1 _25629_ (.A(_09843_),
    .B(_09853_),
    .C(net1031),
    .D(net1118),
    .X(_06683_));
 sg13g2_buf_1 _25630_ (.A(_06683_),
    .X(_06684_));
 sg13g2_inv_1 _25631_ (.Y(_06685_),
    .A(_09835_));
 sg13g2_a21o_1 _25632_ (.A2(_06685_),
    .A1(net1117),
    .B1(_09851_),
    .X(_06686_));
 sg13g2_a221oi_1 _25633_ (.B2(_00178_),
    .C1(_06686_),
    .B1(_06684_),
    .A1(net1114),
    .Y(_06687_),
    .A2(_06682_));
 sg13g2_nor2_1 _25634_ (.A(_09835_),
    .B(net29),
    .Y(_06688_));
 sg13g2_a21oi_1 _25635_ (.A1(net29),
    .A2(_06687_),
    .Y(_02510_),
    .B1(_06688_));
 sg13g2_nor2_1 _25636_ (.A(\cpu.qspi.r_read_delay[1][1] ),
    .B(net245),
    .Y(_06689_));
 sg13g2_mux2_1 _25637_ (.A0(\cpu.qspi.r_read_delay[0][1] ),
    .A1(\cpu.qspi.r_read_delay[2][1] ),
    .S(net245),
    .X(_06690_));
 sg13g2_nor2_1 _25638_ (.A(net88),
    .B(_06690_),
    .Y(_06691_));
 sg13g2_a21oi_1 _25639_ (.A1(net88),
    .A2(_06689_),
    .Y(_06692_),
    .B1(_06691_));
 sg13g2_xnor2_1 _25640_ (.Y(_06693_),
    .A(_09835_),
    .B(_09836_));
 sg13g2_nor2_1 _25641_ (.A(net1117),
    .B(_06684_),
    .Y(_06694_));
 sg13g2_mux2_1 _25642_ (.A0(_06693_),
    .A1(_09911_),
    .S(_06694_),
    .X(_06695_));
 sg13g2_a21oi_1 _25643_ (.A1(net1114),
    .A2(_06692_),
    .Y(_06696_),
    .B1(_06695_));
 sg13g2_nand2_1 _25644_ (.Y(_06697_),
    .A(_11881_),
    .B(_06696_));
 sg13g2_mux2_1 _25645_ (.A0(_09836_),
    .A1(_06697_),
    .S(net29),
    .X(_02511_));
 sg13g2_mux2_1 _25646_ (.A0(\cpu.qspi.r_read_delay[0][2] ),
    .A1(\cpu.qspi.r_read_delay[1][2] ),
    .S(net88),
    .X(_06698_));
 sg13g2_mux2_1 _25647_ (.A0(_06698_),
    .A1(\cpu.qspi.r_read_delay[2][2] ),
    .S(net245),
    .X(_06699_));
 sg13g2_nor2_1 _25648_ (.A(_09835_),
    .B(_09836_),
    .Y(_06700_));
 sg13g2_xor2_1 _25649_ (.B(_06700_),
    .A(_00179_),
    .X(_06701_));
 sg13g2_nor4_2 _25650_ (.A(_09843_),
    .B(_09853_),
    .C(net1031),
    .Y(_06702_),
    .D(net1118));
 sg13g2_o21ai_1 _25651_ (.B1(_09912_),
    .Y(_06703_),
    .A1(net1117),
    .A2(_06702_));
 sg13g2_a22oi_1 _25652_ (.Y(_06704_),
    .B1(_06701_),
    .B2(_06703_),
    .A2(_06694_),
    .A1(net1114));
 sg13g2_or2_1 _25653_ (.X(_06705_),
    .B(_06704_),
    .A(_09851_));
 sg13g2_a21oi_1 _25654_ (.A1(net1114),
    .A2(_06699_),
    .Y(_06706_),
    .B1(_06705_));
 sg13g2_nor2_1 _25655_ (.A(_09837_),
    .B(net29),
    .Y(_06707_));
 sg13g2_a21oi_1 _25656_ (.A1(_06680_),
    .A2(_06706_),
    .Y(_02512_),
    .B1(_06707_));
 sg13g2_a21oi_1 _25657_ (.A1(_09912_),
    .A2(_06702_),
    .Y(_06708_),
    .B1(_09838_));
 sg13g2_nand2b_1 _25658_ (.Y(_06709_),
    .B(net29),
    .A_N(_06708_));
 sg13g2_mux2_1 _25659_ (.A0(\cpu.qspi.r_read_delay[0][3] ),
    .A1(\cpu.qspi.r_read_delay[1][3] ),
    .S(net88),
    .X(_06710_));
 sg13g2_mux2_1 _25660_ (.A0(_06710_),
    .A1(\cpu.qspi.r_read_delay[2][3] ),
    .S(net245),
    .X(_06711_));
 sg13g2_nand2_1 _25661_ (.Y(_06712_),
    .A(_09912_),
    .B(_06702_));
 sg13g2_a22oi_1 _25662_ (.Y(_06713_),
    .B1(_06712_),
    .B2(_09840_),
    .A2(_06711_),
    .A1(net1114));
 sg13g2_nor2b_1 _25663_ (.A(_06713_),
    .B_N(net29),
    .Y(_06714_));
 sg13g2_a21o_1 _25664_ (.A2(_06709_),
    .A1(\cpu.qspi.r_count[3] ),
    .B1(_06714_),
    .X(_02513_));
 sg13g2_and2_1 _25665_ (.A(_09840_),
    .B(_06684_),
    .X(_06715_));
 sg13g2_nor3_1 _25666_ (.A(_09834_),
    .B(_09840_),
    .C(_06694_),
    .Y(_06716_));
 sg13g2_a21oi_1 _25667_ (.A1(_09834_),
    .A2(_06715_),
    .Y(_06717_),
    .B1(_06716_));
 sg13g2_nor2_1 _25668_ (.A(\cpu.qspi.r_count[4] ),
    .B(net29),
    .Y(_06718_));
 sg13g2_a21oi_1 _25669_ (.A1(net29),
    .A2(_06717_),
    .Y(_02514_),
    .B1(_06718_));
 sg13g2_and2_1 _25670_ (.A(_10000_),
    .B(_06321_),
    .X(_06719_));
 sg13g2_buf_2 _25671_ (.A(_06719_),
    .X(_06720_));
 sg13g2_and2_1 _25672_ (.A(_09289_),
    .B(_06720_),
    .X(_06721_));
 sg13g2_buf_1 _25673_ (.A(_06721_),
    .X(_06722_));
 sg13g2_nand2_1 _25674_ (.Y(_06723_),
    .A(net850),
    .B(_06722_));
 sg13g2_nand2_1 _25675_ (.Y(_06724_),
    .A(_09289_),
    .B(_06720_));
 sg13g2_buf_1 _25676_ (.A(_06724_),
    .X(_06725_));
 sg13g2_nand2_1 _25677_ (.Y(_06726_),
    .A(\cpu.qspi.r_read_delay[0][0] ),
    .B(_06725_));
 sg13g2_a21oi_1 _25678_ (.A1(_06723_),
    .A2(_06726_),
    .Y(_02525_),
    .B1(net630));
 sg13g2_nand2_1 _25679_ (.Y(_06727_),
    .A(_06666_),
    .B(_06722_));
 sg13g2_nand2_1 _25680_ (.Y(_06728_),
    .A(\cpu.qspi.r_read_delay[0][1] ),
    .B(_06725_));
 sg13g2_a21oi_1 _25681_ (.A1(_06727_),
    .A2(_06728_),
    .Y(_02526_),
    .B1(net630));
 sg13g2_buf_1 _25682_ (.A(net764),
    .X(_06729_));
 sg13g2_nand2_1 _25683_ (.Y(_06730_),
    .A(net849),
    .B(_06722_));
 sg13g2_nand2_1 _25684_ (.Y(_06731_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_06725_));
 sg13g2_nand3_1 _25685_ (.B(_06730_),
    .C(_06731_),
    .A(net645),
    .Y(_02527_));
 sg13g2_nand2_1 _25686_ (.Y(_06732_),
    .A(net974),
    .B(_06722_));
 sg13g2_nand2_1 _25687_ (.Y(_06733_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_06725_));
 sg13g2_buf_2 _25688_ (.A(net781),
    .X(_06734_));
 sg13g2_buf_1 _25689_ (.A(_06734_),
    .X(_06735_));
 sg13g2_a21oi_1 _25690_ (.A1(_06732_),
    .A2(_06733_),
    .Y(_02528_),
    .B1(net574));
 sg13g2_and2_1 _25691_ (.A(_10120_),
    .B(_06720_),
    .X(_06736_));
 sg13g2_buf_1 _25692_ (.A(_06736_),
    .X(_06737_));
 sg13g2_nand2_1 _25693_ (.Y(_06738_),
    .A(net850),
    .B(_06737_));
 sg13g2_nand2_1 _25694_ (.Y(_06739_),
    .A(_10120_),
    .B(_06720_));
 sg13g2_buf_1 _25695_ (.A(_06739_),
    .X(_06740_));
 sg13g2_nand2_1 _25696_ (.Y(_06741_),
    .A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_06740_));
 sg13g2_a21oi_1 _25697_ (.A1(_06738_),
    .A2(_06741_),
    .Y(_02529_),
    .B1(net574));
 sg13g2_nand2_1 _25698_ (.Y(_06742_),
    .A(_06666_),
    .B(_06737_));
 sg13g2_nand2_1 _25699_ (.Y(_06743_),
    .A(\cpu.qspi.r_read_delay[1][1] ),
    .B(_06740_));
 sg13g2_a21oi_1 _25700_ (.A1(_06742_),
    .A2(_06743_),
    .Y(_02530_),
    .B1(net574));
 sg13g2_nand2_1 _25701_ (.Y(_06744_),
    .A(net849),
    .B(_06737_));
 sg13g2_nand2_1 _25702_ (.Y(_06745_),
    .A(\cpu.qspi.r_read_delay[1][2] ),
    .B(_06740_));
 sg13g2_nand3_1 _25703_ (.B(_06744_),
    .C(_06745_),
    .A(net645),
    .Y(_02531_));
 sg13g2_nand2_1 _25704_ (.Y(_06746_),
    .A(net974),
    .B(_06737_));
 sg13g2_nand2_1 _25705_ (.Y(_06747_),
    .A(\cpu.qspi.r_read_delay[1][3] ),
    .B(_06740_));
 sg13g2_a21oi_1 _25706_ (.A1(_06746_),
    .A2(_06747_),
    .Y(_02532_),
    .B1(net574));
 sg13g2_buf_1 _25707_ (.A(net1029),
    .X(_06748_));
 sg13g2_nor2b_1 _25708_ (.A(net583),
    .B_N(_06720_),
    .Y(_06749_));
 sg13g2_buf_1 _25709_ (.A(_06749_),
    .X(_06750_));
 sg13g2_nand2_1 _25710_ (.Y(_06751_),
    .A(net799),
    .B(_06750_));
 sg13g2_nand2b_1 _25711_ (.Y(_06752_),
    .B(_06720_),
    .A_N(net583));
 sg13g2_buf_1 _25712_ (.A(_06752_),
    .X(_06753_));
 sg13g2_nand2_1 _25713_ (.Y(_06754_),
    .A(\cpu.qspi.r_read_delay[2][0] ),
    .B(_06753_));
 sg13g2_a21oi_1 _25714_ (.A1(_06751_),
    .A2(_06754_),
    .Y(_02533_),
    .B1(net574));
 sg13g2_nand2_1 _25715_ (.Y(_06755_),
    .A(net939),
    .B(_06750_));
 sg13g2_nand2_1 _25716_ (.Y(_06756_),
    .A(\cpu.qspi.r_read_delay[2][1] ),
    .B(_06753_));
 sg13g2_a21oi_1 _25717_ (.A1(_06755_),
    .A2(_06756_),
    .Y(_02534_),
    .B1(net574));
 sg13g2_nand2_1 _25718_ (.Y(_06757_),
    .A(net849),
    .B(_06750_));
 sg13g2_nand2_1 _25719_ (.Y(_06758_),
    .A(\cpu.qspi.r_read_delay[2][2] ),
    .B(_06753_));
 sg13g2_nand3_1 _25720_ (.B(_06757_),
    .C(_06758_),
    .A(net645),
    .Y(_02535_));
 sg13g2_nand2_1 _25721_ (.Y(_06759_),
    .A(net974),
    .B(_06750_));
 sg13g2_nand2_1 _25722_ (.Y(_06760_),
    .A(\cpu.qspi.r_read_delay[2][3] ),
    .B(_06753_));
 sg13g2_a21oi_1 _25723_ (.A1(_06759_),
    .A2(_06760_),
    .Y(_02536_),
    .B1(net574));
 sg13g2_a22oi_1 _25724_ (.Y(_06761_),
    .B1(net88),
    .B2(\cpu.qspi.r_mask[1] ),
    .A2(_09865_),
    .A1(\cpu.qspi.r_mask[2] ));
 sg13g2_nand2_1 _25725_ (.Y(_06762_),
    .A(\cpu.qspi.r_mask[0] ),
    .B(_09866_));
 sg13g2_nand3_1 _25726_ (.B(_06761_),
    .C(_06762_),
    .A(_11882_),
    .Y(_06763_));
 sg13g2_nor3_2 _25727_ (.A(_09843_),
    .B(_09844_),
    .C(_09832_),
    .Y(_06764_));
 sg13g2_nor2_1 _25728_ (.A(net1114),
    .B(net1117),
    .Y(_06765_));
 sg13g2_nand4_1 _25729_ (.B(_06763_),
    .C(_06764_),
    .A(_09831_),
    .Y(_06766_),
    .D(_06765_));
 sg13g2_buf_2 _25730_ (.A(_06766_),
    .X(_06767_));
 sg13g2_buf_1 _25731_ (.A(net892),
    .X(_06768_));
 sg13g2_nor2_1 _25732_ (.A(_09820_),
    .B(_09825_),
    .Y(_06769_));
 sg13g2_buf_1 _25733_ (.A(_06769_),
    .X(_06770_));
 sg13g2_mux2_1 _25734_ (.A0(_09435_),
    .A1(net382),
    .S(net113),
    .X(_06771_));
 sg13g2_nand2_1 _25735_ (.Y(_06772_),
    .A(_09856_),
    .B(_06771_));
 sg13g2_o21ai_1 _25736_ (.B1(_06772_),
    .Y(_06773_),
    .A1(net706),
    .A2(_08648_));
 sg13g2_buf_1 _25737_ (.A(_06770_),
    .X(_06774_));
 sg13g2_mux2_1 _25738_ (.A0(_09692_),
    .A1(_09686_),
    .S(net92),
    .X(_06775_));
 sg13g2_nand2_1 _25739_ (.Y(_06776_),
    .A(_06768_),
    .B(_06775_));
 sg13g2_o21ai_1 _25740_ (.B1(_06776_),
    .Y(_06777_),
    .A1(net706),
    .A2(_08944_));
 sg13g2_buf_1 _25741_ (.A(net1128),
    .X(_06778_));
 sg13g2_buf_1 _25742_ (.A(net938),
    .X(_06779_));
 sg13g2_nor2_1 _25743_ (.A(_09391_),
    .B(_11542_),
    .Y(_06780_));
 sg13g2_nand3_1 _25744_ (.B(_09821_),
    .C(_06780_),
    .A(_00233_),
    .Y(_06781_));
 sg13g2_o21ai_1 _25745_ (.B1(_06781_),
    .Y(_06782_),
    .A1(_09592_),
    .A2(net113));
 sg13g2_nor2_1 _25746_ (.A(net938),
    .B(_06782_),
    .Y(_06783_));
 sg13g2_a21oi_1 _25747_ (.A1(net798),
    .A2(_10737_),
    .Y(_06784_),
    .B1(_06783_));
 sg13g2_inv_1 _25748_ (.Y(_06785_),
    .A(_09854_));
 sg13g2_nor2_1 _25749_ (.A(_09853_),
    .B(net1118),
    .Y(_06786_));
 sg13g2_nand2_1 _25750_ (.Y(_06787_),
    .A(_06675_),
    .B(_06786_));
 sg13g2_nor4_1 _25751_ (.A(_11882_),
    .B(_09900_),
    .C(_09854_),
    .D(\cpu.qspi.r_state[11] ),
    .Y(_06788_));
 sg13g2_nand2_1 _25752_ (.Y(_06789_),
    .A(_09899_),
    .B(_06788_));
 sg13g2_nor3_2 _25753_ (.A(_09851_),
    .B(_06787_),
    .C(_06789_),
    .Y(_06790_));
 sg13g2_nor2_1 _25754_ (.A(_11882_),
    .B(_06790_),
    .Y(_06791_));
 sg13g2_o21ai_1 _25755_ (.B1(_06791_),
    .Y(_06792_),
    .A1(_06785_),
    .A2(net142));
 sg13g2_mux2_1 _25756_ (.A0(_05058_),
    .A1(_05251_),
    .S(_12006_),
    .X(_06793_));
 sg13g2_nor2b_1 _25757_ (.A(_05025_),
    .B_N(_12030_),
    .Y(_06794_));
 sg13g2_a21o_1 _25758_ (.A2(_06793_),
    .A1(net998),
    .B1(_06794_),
    .X(_06795_));
 sg13g2_mux2_1 _25759_ (.A0(_05052_),
    .A1(_05037_),
    .S(_12004_),
    .X(_06796_));
 sg13g2_and2_1 _25760_ (.A(net1096),
    .B(net994),
    .X(_06797_));
 sg13g2_a21oi_1 _25761_ (.A1(_12002_),
    .A2(_05609_),
    .Y(_06798_),
    .B1(net998));
 sg13g2_and3_1 _25762_ (.X(_06799_),
    .A(net998),
    .B(_12002_),
    .C(_05245_));
 sg13g2_o21ai_1 _25763_ (.B1(_12006_),
    .Y(_06800_),
    .A1(_06798_),
    .A2(_06799_));
 sg13g2_o21ai_1 _25764_ (.B1(_06800_),
    .Y(_06801_),
    .A1(_12103_),
    .A2(_12027_));
 sg13g2_a221oi_1 _25765_ (.B2(_06797_),
    .C1(_06801_),
    .B1(_06796_),
    .A1(net999),
    .Y(_06802_),
    .A2(_06795_));
 sg13g2_nor2b_1 _25766_ (.A(_12123_),
    .B_N(_12026_),
    .Y(_06803_));
 sg13g2_nor2_1 _25767_ (.A(net994),
    .B(_06803_),
    .Y(_06804_));
 sg13g2_inv_1 _25768_ (.Y(_06805_),
    .A(_06804_));
 sg13g2_o21ai_1 _25769_ (.B1(net1118),
    .Y(_06806_),
    .A1(_05602_),
    .A2(_06805_));
 sg13g2_inv_1 _25770_ (.Y(_06807_),
    .A(_09833_));
 sg13g2_nand2_1 _25771_ (.Y(_06808_),
    .A(_08264_),
    .B(net1128));
 sg13g2_o21ai_1 _25772_ (.B1(_06808_),
    .Y(_06809_),
    .A1(net1128),
    .A2(_11931_));
 sg13g2_a22oi_1 _25773_ (.Y(_06810_),
    .B1(_06809_),
    .B2(_11917_),
    .A2(\cpu.qspi.r_state[0] ),
    .A1(_06807_));
 sg13g2_o21ai_1 _25774_ (.B1(_06810_),
    .Y(_06811_),
    .A1(_06802_),
    .A2(_06806_));
 sg13g2_nor2_1 _25775_ (.A(_06792_),
    .B(_06811_),
    .Y(_06812_));
 sg13g2_o21ai_1 _25776_ (.B1(_06812_),
    .Y(_06813_),
    .A1(_11915_),
    .A2(_06784_));
 sg13g2_a221oi_1 _25777_ (.B2(_11916_),
    .C1(_06813_),
    .B1(_06777_),
    .A1(_11884_),
    .Y(_06814_),
    .A2(_06773_));
 sg13g2_nand2_1 _25778_ (.Y(_06815_),
    .A(_09900_),
    .B(_09833_));
 sg13g2_nand3_1 _25779_ (.B(_09836_),
    .C(_06815_),
    .A(_06685_),
    .Y(_06816_));
 sg13g2_o21ai_1 _25780_ (.B1(_06816_),
    .Y(_06817_),
    .A1(_06685_),
    .A2(_06815_));
 sg13g2_nor2_1 _25781_ (.A(_09837_),
    .B(_06817_),
    .Y(_06818_));
 sg13g2_nand3b_1 _25782_ (.B(_00178_),
    .C(_06815_),
    .Y(_06819_),
    .A_N(_09836_));
 sg13g2_nor2b_1 _25783_ (.A(net1031),
    .B_N(net142),
    .Y(_06820_));
 sg13g2_o21ai_1 _25784_ (.B1(_09837_),
    .Y(_06821_),
    .A1(_06819_),
    .A2(_06820_));
 sg13g2_nor3_1 _25785_ (.A(net1031),
    .B(_09835_),
    .C(_06821_),
    .Y(_06822_));
 sg13g2_nor2_1 _25786_ (.A(_06818_),
    .B(_06822_),
    .Y(_06823_));
 sg13g2_o21ai_1 _25787_ (.B1(_06818_),
    .Y(_06824_),
    .A1(net1031),
    .A2(_09836_));
 sg13g2_o21ai_1 _25788_ (.B1(_06824_),
    .Y(_06825_),
    .A1(_09836_),
    .A2(_06821_));
 sg13g2_inv_1 _25789_ (.Y(_06826_),
    .A(_06825_));
 sg13g2_o21ai_1 _25790_ (.B1(_06826_),
    .Y(_06827_),
    .A1(net142),
    .A2(_06823_));
 sg13g2_o21ai_1 _25791_ (.B1(_06827_),
    .Y(_06828_),
    .A1(_09853_),
    .A2(net1031));
 sg13g2_xnor2_1 _25792_ (.Y(_06829_),
    .A(net142),
    .B(_09869_));
 sg13g2_a221oi_1 _25793_ (.B2(_06790_),
    .C1(_06767_),
    .B1(_06829_),
    .A1(_06814_),
    .Y(_06830_),
    .A2(_06828_));
 sg13g2_a21o_1 _25794_ (.A2(_06767_),
    .A1(net11),
    .B1(_06830_),
    .X(_02541_));
 sg13g2_nor2_1 _25795_ (.A(_09574_),
    .B(net92),
    .Y(_06831_));
 sg13g2_a21oi_1 _25796_ (.A1(_09568_),
    .A2(net92),
    .Y(_06832_),
    .B1(_06831_));
 sg13g2_nand2b_1 _25797_ (.Y(_06833_),
    .B(net798),
    .A_N(_10981_));
 sg13g2_o21ai_1 _25798_ (.B1(_06833_),
    .Y(_06834_),
    .A1(net798),
    .A2(_06832_));
 sg13g2_and2_1 _25799_ (.A(net1096),
    .B(_12026_),
    .X(_06835_));
 sg13g2_a221oi_1 _25800_ (.B2(_05405_),
    .C1(net998),
    .B1(_06835_),
    .A1(_12006_),
    .Y(_06836_),
    .A2(_05676_));
 sg13g2_mux2_1 _25801_ (.A0(_05271_),
    .A1(_05388_),
    .S(net1096),
    .X(_06837_));
 sg13g2_a21oi_1 _25802_ (.A1(net999),
    .A2(_06837_),
    .Y(_06838_),
    .B1(_12004_));
 sg13g2_mux2_1 _25803_ (.A0(_05265_),
    .A1(_05381_),
    .S(net1096),
    .X(_06839_));
 sg13g2_a22oi_1 _25804_ (.Y(_06840_),
    .B1(_06839_),
    .B2(net998),
    .A2(_05397_),
    .A1(_12030_));
 sg13g2_nand2b_1 _25805_ (.Y(_06841_),
    .B(net994),
    .A_N(_06840_));
 sg13g2_o21ai_1 _25806_ (.B1(_06841_),
    .Y(_06842_),
    .A1(_06836_),
    .A2(_06838_));
 sg13g2_mux2_1 _25807_ (.A0(_05669_),
    .A1(_06842_),
    .S(_06805_),
    .X(_06843_));
 sg13g2_a221oi_1 _25808_ (.B2(_09846_),
    .C1(_06792_),
    .B1(_06843_),
    .A1(_11917_),
    .Y(_06844_),
    .A2(_06834_));
 sg13g2_nand2_1 _25809_ (.Y(_06845_),
    .A(net380),
    .B(net113));
 sg13g2_o21ai_1 _25810_ (.B1(_06845_),
    .Y(_06846_),
    .A1(_09529_),
    .A2(net92));
 sg13g2_nand2_1 _25811_ (.Y(_06847_),
    .A(net706),
    .B(_06846_));
 sg13g2_o21ai_1 _25812_ (.B1(_06847_),
    .Y(_06848_),
    .A1(net706),
    .A2(_08900_));
 sg13g2_mux2_1 _25813_ (.A0(_09605_),
    .A1(_00235_),
    .S(net92),
    .X(_06849_));
 sg13g2_and2_1 _25814_ (.A(net798),
    .B(_11109_),
    .X(_06850_));
 sg13g2_a21oi_1 _25815_ (.A1(net706),
    .A2(_06849_),
    .Y(_06851_),
    .B1(_06850_));
 sg13g2_mux2_1 _25816_ (.A0(_09471_),
    .A1(net381),
    .S(net92),
    .X(_06852_));
 sg13g2_nor2_1 _25817_ (.A(net892),
    .B(_08681_),
    .Y(_06853_));
 sg13g2_a21oi_1 _25818_ (.A1(net706),
    .A2(_06852_),
    .Y(_06854_),
    .B1(_06853_));
 sg13g2_nor2b_1 _25819_ (.A(_06854_),
    .B_N(_11884_),
    .Y(_06855_));
 sg13g2_a221oi_1 _25820_ (.B2(_11914_),
    .C1(_06855_),
    .B1(_06851_),
    .A1(_11916_),
    .Y(_06856_),
    .A2(_06848_));
 sg13g2_a221oi_1 _25821_ (.B2(_06856_),
    .C1(_06767_),
    .B1(_06844_),
    .A1(_09869_),
    .Y(_06857_),
    .A2(_06790_));
 sg13g2_a21o_1 _25822_ (.A2(_06767_),
    .A1(net12),
    .B1(_06857_),
    .X(_02542_));
 sg13g2_mux2_1 _25823_ (.A0(_09761_),
    .A1(_09754_),
    .S(net92),
    .X(_06858_));
 sg13g2_nor2_1 _25824_ (.A(net892),
    .B(_08855_),
    .Y(_06859_));
 sg13g2_a21oi_1 _25825_ (.A1(net706),
    .A2(_06858_),
    .Y(_06860_),
    .B1(_06859_));
 sg13g2_nor2b_1 _25826_ (.A(_06860_),
    .B_N(_11916_),
    .Y(_06861_));
 sg13g2_a221oi_1 _25827_ (.B2(_05427_),
    .C1(net998),
    .B1(_06797_),
    .A1(_12006_),
    .Y(_06862_),
    .A2(_05706_));
 sg13g2_mux2_1 _25828_ (.A0(_05173_),
    .A1(_05297_),
    .S(_12006_),
    .X(_06863_));
 sg13g2_a21oi_1 _25829_ (.A1(_12103_),
    .A2(_06863_),
    .Y(_06864_),
    .B1(_12004_));
 sg13g2_mux2_1 _25830_ (.A0(_05166_),
    .A1(_05303_),
    .S(_12006_),
    .X(_06865_));
 sg13g2_a22oi_1 _25831_ (.Y(_06866_),
    .B1(_06865_),
    .B2(_12028_),
    .A2(_05421_),
    .A1(_12030_));
 sg13g2_nand2b_1 _25832_ (.Y(_06867_),
    .B(net999),
    .A_N(_06866_));
 sg13g2_o21ai_1 _25833_ (.B1(_06867_),
    .Y(_06868_),
    .A1(_06862_),
    .A2(_06864_));
 sg13g2_mux2_1 _25834_ (.A0(_05700_),
    .A1(_06868_),
    .S(_06805_),
    .X(_06869_));
 sg13g2_nand3_1 _25835_ (.B(_09821_),
    .C(_06780_),
    .A(_00229_),
    .Y(_06870_));
 sg13g2_o21ai_1 _25836_ (.B1(_06870_),
    .Y(_06871_),
    .A1(_09581_),
    .A2(net113));
 sg13g2_nand2_1 _25837_ (.Y(_06872_),
    .A(net938),
    .B(_03651_));
 sg13g2_o21ai_1 _25838_ (.B1(_06872_),
    .Y(_06873_),
    .A1(net938),
    .A2(_06871_));
 sg13g2_mux2_1 _25839_ (.A0(_08279_),
    .A1(net767),
    .S(net892),
    .X(_06874_));
 sg13g2_o21ai_1 _25840_ (.B1(_06791_),
    .Y(_06875_),
    .A1(_00180_),
    .A2(_06874_));
 sg13g2_a221oi_1 _25841_ (.B2(_11917_),
    .C1(_06875_),
    .B1(_06873_),
    .A1(net1118),
    .Y(_06876_),
    .A2(_06869_));
 sg13g2_inv_1 _25842_ (.Y(_06877_),
    .A(_09623_));
 sg13g2_mux2_1 _25843_ (.A0(_06877_),
    .A1(_00237_),
    .S(net113),
    .X(_06878_));
 sg13g2_nand2b_1 _25844_ (.Y(_06879_),
    .B(_06778_),
    .A_N(_10738_));
 sg13g2_o21ai_1 _25845_ (.B1(_06879_),
    .Y(_06880_),
    .A1(net938),
    .A2(_06878_));
 sg13g2_mux2_1 _25846_ (.A0(_09537_),
    .A1(net379),
    .S(net113),
    .X(_06881_));
 sg13g2_nor2_1 _25847_ (.A(net892),
    .B(_08879_),
    .Y(_06882_));
 sg13g2_a21o_1 _25848_ (.A2(_06881_),
    .A1(net892),
    .B1(_06882_),
    .X(_06883_));
 sg13g2_a22oi_1 _25849_ (.Y(_06884_),
    .B1(_06883_),
    .B2(_11884_),
    .A2(_06880_),
    .A1(_11914_));
 sg13g2_nand2_1 _25850_ (.Y(_06885_),
    .A(_06876_),
    .B(_06884_));
 sg13g2_nor2_1 _25851_ (.A(_06861_),
    .B(_06885_),
    .Y(_06886_));
 sg13g2_nor2_1 _25852_ (.A(net142),
    .B(_09869_),
    .Y(_06887_));
 sg13g2_nor2b_1 _25853_ (.A(_06887_),
    .B_N(_06790_),
    .Y(_06888_));
 sg13g2_nor3_1 _25854_ (.A(_06767_),
    .B(_06886_),
    .C(_06888_),
    .Y(_06889_));
 sg13g2_a21o_1 _25855_ (.A2(_06767_),
    .A1(net13),
    .B1(_06889_),
    .X(_02543_));
 sg13g2_mux2_1 _25856_ (.A0(_09699_),
    .A1(_09713_),
    .S(net113),
    .X(_06890_));
 sg13g2_nand2_1 _25857_ (.Y(_06891_),
    .A(net1128),
    .B(_08988_));
 sg13g2_o21ai_1 _25858_ (.B1(_06891_),
    .Y(_06892_),
    .A1(net938),
    .A2(_06890_));
 sg13g2_nor2b_1 _25859_ (.A(_06892_),
    .B_N(_11884_),
    .Y(_06893_));
 sg13g2_and2_1 _25860_ (.A(net702),
    .B(net1128),
    .X(_06894_));
 sg13g2_a21oi_1 _25861_ (.A1(net892),
    .A2(_09266_),
    .Y(_06895_),
    .B1(_06894_));
 sg13g2_o21ai_1 _25862_ (.B1(_06677_),
    .Y(_06896_),
    .A1(_00180_),
    .A2(_06895_));
 sg13g2_mux4_1 _25863_ (.S0(_12004_),
    .A0(_05151_),
    .A1(_05137_),
    .A2(_05207_),
    .A3(_05501_),
    .S1(net1096),
    .X(_06897_));
 sg13g2_inv_1 _25864_ (.Y(_06898_),
    .A(_05493_));
 sg13g2_mux2_1 _25865_ (.A0(_05145_),
    .A1(_05215_),
    .S(net1096),
    .X(_06899_));
 sg13g2_a22oi_1 _25866_ (.Y(_06900_),
    .B1(_06899_),
    .B2(net998),
    .A2(_06898_),
    .A1(_12030_));
 sg13g2_nor2b_1 _25867_ (.A(_06900_),
    .B_N(net999),
    .Y(_06901_));
 sg13g2_a221oi_1 _25868_ (.B2(net994),
    .C1(_06901_),
    .B1(_06897_),
    .A1(_05130_),
    .Y(_06902_),
    .A2(_06804_));
 sg13g2_nor2b_1 _25869_ (.A(_06902_),
    .B_N(_09846_),
    .Y(_06903_));
 sg13g2_nor4_1 _25870_ (.A(_06790_),
    .B(_06893_),
    .C(_06896_),
    .D(_06903_),
    .Y(_06904_));
 sg13g2_mux2_1 _25871_ (.A0(_09648_),
    .A1(net378),
    .S(net113),
    .X(_06905_));
 sg13g2_nor2_1 _25872_ (.A(net938),
    .B(_06905_),
    .Y(_06906_));
 sg13g2_a21oi_1 _25873_ (.A1(net798),
    .A2(_08758_),
    .Y(_06907_),
    .B1(_06906_));
 sg13g2_nor3_1 _25874_ (.A(_09859_),
    .B(_09861_),
    .C(_11880_),
    .Y(_06908_));
 sg13g2_mux2_1 _25875_ (.A0(_09565_),
    .A1(_00239_),
    .S(net92),
    .X(_06909_));
 sg13g2_nand2_1 _25876_ (.Y(_06910_),
    .A(net938),
    .B(_04338_));
 sg13g2_o21ai_1 _25877_ (.B1(_06910_),
    .Y(_06911_),
    .A1(net798),
    .A2(_06909_));
 sg13g2_a22oi_1 _25878_ (.Y(_06912_),
    .B1(_06911_),
    .B2(_11914_),
    .A2(_06908_),
    .A1(_06907_));
 sg13g2_nand2_1 _25879_ (.Y(_06913_),
    .A(_00231_),
    .B(_06774_));
 sg13g2_o21ai_1 _25880_ (.B1(_06913_),
    .Y(_06914_),
    .A1(_09616_),
    .A2(_06774_));
 sg13g2_nand2_1 _25881_ (.Y(_06915_),
    .A(_06778_),
    .B(_03645_));
 sg13g2_o21ai_1 _25882_ (.B1(_06915_),
    .Y(_06916_),
    .A1(net798),
    .A2(_06914_));
 sg13g2_mux2_1 _25883_ (.A0(_09671_),
    .A1(_09665_),
    .S(_06770_),
    .X(_06917_));
 sg13g2_nand2_1 _25884_ (.Y(_06918_),
    .A(_09856_),
    .B(_06917_));
 sg13g2_o21ai_1 _25885_ (.B1(_06918_),
    .Y(_06919_),
    .A1(net706),
    .A2(_08735_));
 sg13g2_a22oi_1 _25886_ (.Y(_06920_),
    .B1(_06919_),
    .B2(_11916_),
    .A2(_06916_),
    .A1(_11917_));
 sg13g2_and3_1 _25887_ (.X(_06921_),
    .A(_06904_),
    .B(_06912_),
    .C(_06920_));
 sg13g2_nor3_1 _25888_ (.A(_06767_),
    .B(_06888_),
    .C(_06921_),
    .Y(_06922_));
 sg13g2_a21o_1 _25889_ (.A2(_06767_),
    .A1(net14),
    .B1(_06922_),
    .X(_02544_));
 sg13g2_mux4_1 _25890_ (.S0(_05573_),
    .A0(_09234_),
    .A1(_09236_),
    .A2(_09222_),
    .A3(_09217_),
    .S1(_06334_),
    .X(_06923_));
 sg13g2_mux4_1 _25891_ (.S0(_05573_),
    .A0(_09220_),
    .A1(_09226_),
    .A2(_09215_),
    .A3(_09230_),
    .S1(_06334_),
    .X(_06924_));
 sg13g2_nor2b_1 _25892_ (.A(\cpu.gpio.r_spi_miso_src[1][2] ),
    .B_N(_06924_),
    .Y(_06925_));
 sg13g2_a21oi_1 _25893_ (.A1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .A2(_06923_),
    .Y(_06926_),
    .B1(_06925_));
 sg13g2_mux4_1 _25894_ (.S0(_05573_),
    .A0(_09239_),
    .A1(_09241_),
    .A2(_09231_),
    .A3(_09227_),
    .S1(_06334_),
    .X(_06927_));
 sg13g2_nand3_1 _25895_ (.B(\cpu.gpio.r_spi_miso_src[1][3] ),
    .C(_06927_),
    .A(_05712_),
    .Y(_06928_));
 sg13g2_o21ai_1 _25896_ (.B1(_06928_),
    .Y(_06929_),
    .A1(\cpu.gpio.r_spi_miso_src[1][3] ),
    .A2(_06926_));
 sg13g2_mux4_1 _25897_ (.S0(_04932_),
    .A0(_09234_),
    .A1(_09236_),
    .A2(_09222_),
    .A3(_09217_),
    .S1(_06332_),
    .X(_06930_));
 sg13g2_mux4_1 _25898_ (.S0(_04932_),
    .A0(_09220_),
    .A1(_09226_),
    .A2(_09215_),
    .A3(_09230_),
    .S1(_06332_),
    .X(_06931_));
 sg13g2_nor2b_1 _25899_ (.A(\cpu.gpio.r_spi_miso_src[0][2] ),
    .B_N(_06931_),
    .Y(_06932_));
 sg13g2_a21oi_1 _25900_ (.A1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .A2(_06930_),
    .Y(_06933_),
    .B1(_06932_));
 sg13g2_mux4_1 _25901_ (.S0(_04932_),
    .A0(_09239_),
    .A1(_09241_),
    .A2(_09231_),
    .A3(_09227_),
    .S1(_06332_),
    .X(_06934_));
 sg13g2_nand3_1 _25902_ (.B(\cpu.gpio.r_spi_miso_src[0][3] ),
    .C(_06934_),
    .A(_05452_),
    .Y(_06935_));
 sg13g2_o21ai_1 _25903_ (.B1(_06935_),
    .Y(_06936_),
    .A1(\cpu.gpio.r_spi_miso_src[0][3] ),
    .A2(_06933_));
 sg13g2_mux2_1 _25904_ (.A0(_06929_),
    .A1(_06936_),
    .S(_11959_),
    .X(_06937_));
 sg13g2_nor2_1 _25905_ (.A(net1122),
    .B(_11985_),
    .Y(_06938_));
 sg13g2_nor2b_1 _25906_ (.A(net1038),
    .B_N(net1122),
    .Y(_06939_));
 sg13g2_a22oi_1 _25907_ (.Y(_06940_),
    .B1(_06939_),
    .B2(net604),
    .A2(_06938_),
    .A1(net1038));
 sg13g2_nor3_1 _25908_ (.A(net781),
    .B(net419),
    .C(_06940_),
    .Y(_06941_));
 sg13g2_buf_4 _25909_ (.X(_06942_),
    .A(_06941_));
 sg13g2_mux2_1 _25910_ (.A0(_09320_),
    .A1(_06937_),
    .S(_06942_),
    .X(_02584_));
 sg13g2_mux2_1 _25911_ (.A0(_09319_),
    .A1(_09320_),
    .S(_06942_),
    .X(_02585_));
 sg13g2_mux2_1 _25912_ (.A0(_09323_),
    .A1(_09319_),
    .S(_06942_),
    .X(_02586_));
 sg13g2_mux2_1 _25913_ (.A0(_09317_),
    .A1(_09323_),
    .S(_06942_),
    .X(_02587_));
 sg13g2_mux2_1 _25914_ (.A0(_09325_),
    .A1(_09317_),
    .S(_06942_),
    .X(_02588_));
 sg13g2_mux2_1 _25915_ (.A0(_09324_),
    .A1(_09325_),
    .S(_06942_),
    .X(_02589_));
 sg13g2_mux2_1 _25916_ (.A0(_09318_),
    .A1(_09324_),
    .S(_06942_),
    .X(_02590_));
 sg13g2_mux2_1 _25917_ (.A0(\cpu.spi.r_in[7] ),
    .A1(_09318_),
    .S(_06942_),
    .X(_02591_));
 sg13g2_nand2_1 _25918_ (.Y(_06943_),
    .A(_09285_),
    .B(_09290_));
 sg13g2_nor2_1 _25919_ (.A(_09285_),
    .B(_09195_),
    .Y(_06944_));
 sg13g2_a22oi_1 _25920_ (.Y(_06945_),
    .B1(_06944_),
    .B2(_11924_),
    .A2(_11986_),
    .A1(net1121));
 sg13g2_nand4_1 _25921_ (.B(_11981_),
    .C(_11991_),
    .A(_06943_),
    .Y(_06946_),
    .D(_06945_));
 sg13g2_buf_1 _25922_ (.A(_06946_),
    .X(_06947_));
 sg13g2_buf_1 _25923_ (.A(_00223_),
    .X(_06948_));
 sg13g2_nor2b_1 _25924_ (.A(net604),
    .B_N(_00221_),
    .Y(_06949_));
 sg13g2_o21ai_1 _25925_ (.B1(_09357_),
    .Y(_06950_),
    .A1(_06948_),
    .A2(_06949_));
 sg13g2_o21ai_1 _25926_ (.B1(_06950_),
    .Y(_06951_),
    .A1(_09357_),
    .A2(_10047_));
 sg13g2_a21oi_1 _25927_ (.A1(_11924_),
    .A2(_06951_),
    .Y(_06952_),
    .B1(net72));
 sg13g2_a21o_1 _25928_ (.A2(net72),
    .A1(\cpu.spi.r_out[0] ),
    .B1(_06952_),
    .X(_02599_));
 sg13g2_mux2_1 _25929_ (.A0(_00181_),
    .A1(_00221_),
    .S(net604),
    .X(_06953_));
 sg13g2_nor2_1 _25930_ (.A(_09195_),
    .B(net854),
    .Y(_06954_));
 sg13g2_buf_2 _25931_ (.A(_06954_),
    .X(_06955_));
 sg13g2_a22oi_1 _25932_ (.Y(_06956_),
    .B1(_06955_),
    .B2(_10069_),
    .A2(net854),
    .A1(\cpu.spi.r_out[0] ));
 sg13g2_o21ai_1 _25933_ (.B1(_06956_),
    .Y(_06957_),
    .A1(net898),
    .A2(_06953_));
 sg13g2_mux2_1 _25934_ (.A0(_06957_),
    .A1(\cpu.spi.r_out[1] ),
    .S(_06947_),
    .X(_02600_));
 sg13g2_mux2_1 _25935_ (.A0(_00182_),
    .A1(_00181_),
    .S(net604),
    .X(_06958_));
 sg13g2_a22oi_1 _25936_ (.Y(_06959_),
    .B1(_06955_),
    .B2(net1020),
    .A2(net854),
    .A1(\cpu.spi.r_out[1] ));
 sg13g2_o21ai_1 _25937_ (.B1(_06959_),
    .Y(_06960_),
    .A1(net898),
    .A2(_06958_));
 sg13g2_mux2_1 _25938_ (.A0(_06960_),
    .A1(\cpu.spi.r_out[2] ),
    .S(net72),
    .X(_02601_));
 sg13g2_mux2_1 _25939_ (.A0(_00285_),
    .A1(_00182_),
    .S(net604),
    .X(_06961_));
 sg13g2_a22oi_1 _25940_ (.Y(_06962_),
    .B1(_06955_),
    .B2(_10079_),
    .A2(net854),
    .A1(\cpu.spi.r_out[2] ));
 sg13g2_o21ai_1 _25941_ (.B1(_06962_),
    .Y(_06963_),
    .A1(net898),
    .A2(_06961_));
 sg13g2_mux2_1 _25942_ (.A0(_06963_),
    .A1(\cpu.spi.r_out[3] ),
    .S(net72),
    .X(_02602_));
 sg13g2_mux2_1 _25943_ (.A0(_00183_),
    .A1(_00285_),
    .S(net604),
    .X(_06964_));
 sg13g2_a22oi_1 _25944_ (.Y(_06965_),
    .B1(_06955_),
    .B2(_10085_),
    .A2(net854),
    .A1(\cpu.spi.r_out[3] ));
 sg13g2_o21ai_1 _25945_ (.B1(_06965_),
    .Y(_06966_),
    .A1(net898),
    .A2(_06964_));
 sg13g2_mux2_1 _25946_ (.A0(_06966_),
    .A1(\cpu.spi.r_out[4] ),
    .S(net72),
    .X(_02603_));
 sg13g2_mux2_1 _25947_ (.A0(_00184_),
    .A1(_00183_),
    .S(net604),
    .X(_06967_));
 sg13g2_a22oi_1 _25948_ (.Y(_06968_),
    .B1(_06955_),
    .B2(_10091_),
    .A2(net854),
    .A1(\cpu.spi.r_out[4] ));
 sg13g2_o21ai_1 _25949_ (.B1(_06968_),
    .Y(_06969_),
    .A1(net898),
    .A2(_06967_));
 sg13g2_mux2_1 _25950_ (.A0(_06969_),
    .A1(\cpu.spi.r_out[5] ),
    .S(net72),
    .X(_02604_));
 sg13g2_buf_1 _25951_ (.A(_00185_),
    .X(_06970_));
 sg13g2_mux2_1 _25952_ (.A0(_06970_),
    .A1(_00184_),
    .S(_11993_),
    .X(_06971_));
 sg13g2_a22oi_1 _25953_ (.Y(_06972_),
    .B1(_06955_),
    .B2(_10097_),
    .A2(net854),
    .A1(\cpu.spi.r_out[5] ));
 sg13g2_o21ai_1 _25954_ (.B1(_06972_),
    .Y(_06973_),
    .A1(_09340_),
    .A2(_06971_));
 sg13g2_mux2_1 _25955_ (.A0(_06973_),
    .A1(\cpu.spi.r_out[6] ),
    .S(net72),
    .X(_02605_));
 sg13g2_buf_1 _25956_ (.A(_00279_),
    .X(_06974_));
 sg13g2_mux2_1 _25957_ (.A0(_06974_),
    .A1(_06970_),
    .S(_11993_),
    .X(_06975_));
 sg13g2_a22oi_1 _25958_ (.Y(_06976_),
    .B1(_06955_),
    .B2(_10103_),
    .A2(net854),
    .A1(\cpu.spi.r_out[6] ));
 sg13g2_o21ai_1 _25959_ (.B1(_06976_),
    .Y(_06977_),
    .A1(_09340_),
    .A2(_06975_));
 sg13g2_mux2_1 _25960_ (.A0(_06977_),
    .A1(\cpu.spi.r_out[7] ),
    .S(net72),
    .X(_02606_));
 sg13g2_or2_1 _25961_ (.X(_06978_),
    .B(_09355_),
    .A(net781));
 sg13g2_buf_1 _25962_ (.A(_06978_),
    .X(_06979_));
 sg13g2_nand2_1 _25963_ (.Y(_06980_),
    .A(net732),
    .B(_06979_));
 sg13g2_o21ai_1 _25964_ (.B1(_06980_),
    .Y(_02609_),
    .A1(_03865_),
    .A2(_06979_));
 sg13g2_nand2_1 _25965_ (.Y(_06981_),
    .A(net857),
    .B(_06979_));
 sg13g2_o21ai_1 _25966_ (.B1(_06981_),
    .Y(_02610_),
    .A1(_02970_),
    .A2(_06979_));
 sg13g2_and2_1 _25967_ (.A(_09344_),
    .B(_05082_),
    .X(_06982_));
 sg13g2_buf_4 _25968_ (.X(_06983_),
    .A(_06982_));
 sg13g2_mux2_1 _25969_ (.A0(\cpu.spi.r_timeout[0] ),
    .A1(net890),
    .S(_06983_),
    .X(_02614_));
 sg13g2_mux2_1 _25970_ (.A0(\cpu.spi.r_timeout[1] ),
    .A1(net939),
    .S(_06983_),
    .X(_02615_));
 sg13g2_mux2_1 _25971_ (.A0(\cpu.spi.r_timeout[2] ),
    .A1(net886),
    .S(_06983_),
    .X(_02616_));
 sg13g2_mux2_1 _25972_ (.A0(\cpu.spi.r_timeout[3] ),
    .A1(net885),
    .S(_06983_),
    .X(_02617_));
 sg13g2_mux2_1 _25973_ (.A0(\cpu.spi.r_timeout[4] ),
    .A1(_12130_),
    .S(_06983_),
    .X(_02618_));
 sg13g2_mux2_1 _25974_ (.A0(\cpu.spi.r_timeout[5] ),
    .A1(net990),
    .S(_06983_),
    .X(_02619_));
 sg13g2_mux2_1 _25975_ (.A0(\cpu.spi.r_timeout[6] ),
    .A1(net989),
    .S(_06983_),
    .X(_02620_));
 sg13g2_mux2_1 _25976_ (.A0(\cpu.spi.r_timeout[7] ),
    .A1(net851),
    .S(_06983_),
    .X(_02621_));
 sg13g2_nand2_1 _25977_ (.Y(_06984_),
    .A(_09196_),
    .B(_11988_));
 sg13g2_nand2_1 _25978_ (.Y(_06985_),
    .A(_09316_),
    .B(_09329_));
 sg13g2_or4_1 _25979_ (.A(_00224_),
    .B(_09193_),
    .C(_09301_),
    .D(_06985_),
    .X(_06986_));
 sg13g2_o21ai_1 _25980_ (.B1(net1038),
    .Y(_06987_),
    .A1(_09193_),
    .A2(_06985_));
 sg13g2_nand4_1 _25981_ (.B(_06984_),
    .C(_06986_),
    .A(_11981_),
    .Y(_06988_),
    .D(_06987_));
 sg13g2_buf_2 _25982_ (.A(_06988_),
    .X(_06989_));
 sg13g2_buf_1 _25983_ (.A(_06989_),
    .X(_06990_));
 sg13g2_and2_1 _25984_ (.A(net897),
    .B(\cpu.spi.r_timeout[0] ),
    .X(_06991_));
 sg13g2_a21oi_1 _25985_ (.A1(net898),
    .A2(_00282_),
    .Y(_06992_),
    .B1(_06991_));
 sg13g2_nand2_1 _25986_ (.Y(_06993_),
    .A(_09303_),
    .B(net60));
 sg13g2_o21ai_1 _25987_ (.B1(_06993_),
    .Y(_02622_),
    .A1(net60),
    .A2(_06992_));
 sg13g2_nor3_1 _25988_ (.A(_09303_),
    .B(_09304_),
    .C(_06989_),
    .Y(_06994_));
 sg13g2_a21oi_1 _25989_ (.A1(_09303_),
    .A2(_09304_),
    .Y(_06995_),
    .B1(_06994_));
 sg13g2_nor2_1 _25990_ (.A(_09196_),
    .B(_06989_),
    .Y(_06996_));
 sg13g2_buf_2 _25991_ (.A(_06996_),
    .X(_06997_));
 sg13g2_a22oi_1 _25992_ (.Y(_06998_),
    .B1(_06997_),
    .B2(\cpu.spi.r_timeout[1] ),
    .A2(net60),
    .A1(_09304_));
 sg13g2_o21ai_1 _25993_ (.B1(_06998_),
    .Y(_02623_),
    .A1(_09358_),
    .A2(_06995_));
 sg13g2_a22oi_1 _25994_ (.Y(_06999_),
    .B1(_06997_),
    .B2(\cpu.spi.r_timeout[2] ),
    .A2(_06990_),
    .A1(\cpu.spi.r_timeout_count[2] ));
 sg13g2_o21ai_1 _25995_ (.B1(\cpu.spi.r_timeout_count[2] ),
    .Y(_07000_),
    .A1(_09303_),
    .A2(_09304_));
 sg13g2_o21ai_1 _25996_ (.B1(_07000_),
    .Y(_07001_),
    .A1(_09306_),
    .A2(_06990_));
 sg13g2_nand2_1 _25997_ (.Y(_07002_),
    .A(net898),
    .B(_07001_));
 sg13g2_nand2_1 _25998_ (.Y(_02624_),
    .A(_06999_),
    .B(_07002_));
 sg13g2_nor2_1 _25999_ (.A(_09308_),
    .B(_06989_),
    .Y(_07003_));
 sg13g2_a21oi_1 _26000_ (.A1(\cpu.spi.r_timeout_count[3] ),
    .A2(_09306_),
    .Y(_07004_),
    .B1(_07003_));
 sg13g2_a22oi_1 _26001_ (.Y(_07005_),
    .B1(_06997_),
    .B2(\cpu.spi.r_timeout[3] ),
    .A2(net60),
    .A1(\cpu.spi.r_timeout_count[3] ));
 sg13g2_o21ai_1 _26002_ (.B1(_07005_),
    .Y(_02625_),
    .A1(net897),
    .A2(_07004_));
 sg13g2_nor2_1 _26003_ (.A(_09310_),
    .B(_06989_),
    .Y(_07006_));
 sg13g2_a21oi_1 _26004_ (.A1(\cpu.spi.r_timeout_count[4] ),
    .A2(_09308_),
    .Y(_07007_),
    .B1(_07006_));
 sg13g2_a22oi_1 _26005_ (.Y(_07008_),
    .B1(_06997_),
    .B2(\cpu.spi.r_timeout[4] ),
    .A2(net60),
    .A1(\cpu.spi.r_timeout_count[4] ));
 sg13g2_o21ai_1 _26006_ (.B1(_07008_),
    .Y(_02626_),
    .A1(net897),
    .A2(_07007_));
 sg13g2_nor2_1 _26007_ (.A(_09312_),
    .B(_06989_),
    .Y(_07009_));
 sg13g2_a21oi_1 _26008_ (.A1(\cpu.spi.r_timeout_count[5] ),
    .A2(_09310_),
    .Y(_07010_),
    .B1(_07009_));
 sg13g2_a22oi_1 _26009_ (.Y(_07011_),
    .B1(_06997_),
    .B2(\cpu.spi.r_timeout[5] ),
    .A2(net60),
    .A1(\cpu.spi.r_timeout_count[5] ));
 sg13g2_o21ai_1 _26010_ (.B1(_07011_),
    .Y(_02627_),
    .A1(net897),
    .A2(_07010_));
 sg13g2_nor2_1 _26011_ (.A(_09314_),
    .B(_06989_),
    .Y(_07012_));
 sg13g2_a21oi_1 _26012_ (.A1(\cpu.spi.r_timeout_count[6] ),
    .A2(_09312_),
    .Y(_07013_),
    .B1(_07012_));
 sg13g2_a22oi_1 _26013_ (.Y(_07014_),
    .B1(_06997_),
    .B2(\cpu.spi.r_timeout[6] ),
    .A2(net60),
    .A1(\cpu.spi.r_timeout_count[6] ));
 sg13g2_o21ai_1 _26014_ (.B1(_07014_),
    .Y(_02628_),
    .A1(net897),
    .A2(_07013_));
 sg13g2_nor3_1 _26015_ (.A(_09302_),
    .B(_09314_),
    .C(_06989_),
    .Y(_07015_));
 sg13g2_a21oi_1 _26016_ (.A1(_09302_),
    .A2(_09314_),
    .Y(_07016_),
    .B1(_07015_));
 sg13g2_a22oi_1 _26017_ (.Y(_07017_),
    .B1(_06997_),
    .B2(\cpu.spi.r_timeout[7] ),
    .A2(net60),
    .A1(_09302_));
 sg13g2_o21ai_1 _26018_ (.B1(_07017_),
    .Y(_02629_),
    .A1(net897),
    .A2(_07016_));
 sg13g2_buf_1 _26019_ (.A(\cpu.uart.r_rcnt[0] ),
    .X(_07018_));
 sg13g2_nor2_1 _26020_ (.A(_07018_),
    .B(\cpu.uart.r_rcnt[1] ),
    .Y(_07019_));
 sg13g2_nand2_1 _26021_ (.Y(_07020_),
    .A(_09930_),
    .B(_07019_));
 sg13g2_nor2_1 _26022_ (.A(net899),
    .B(_07020_),
    .Y(_07021_));
 sg13g2_buf_1 _26023_ (.A(\cpu.uart.r_rstate[3] ),
    .X(_07022_));
 sg13g2_buf_1 _26024_ (.A(net1080),
    .X(_07023_));
 sg13g2_buf_1 _26025_ (.A(\cpu.uart.r_rstate[1] ),
    .X(_07024_));
 sg13g2_buf_1 _26026_ (.A(\cpu.uart.r_rstate[2] ),
    .X(_07025_));
 sg13g2_nor2_2 _26027_ (.A(net1079),
    .B(_07025_),
    .Y(_07026_));
 sg13g2_buf_2 _26028_ (.A(\cpu.uart.r_rstate[0] ),
    .X(_07027_));
 sg13g2_inv_1 _26029_ (.Y(_07028_),
    .A(_07027_));
 sg13g2_nand3_1 _26030_ (.B(_07023_),
    .C(_07026_),
    .A(_07028_),
    .Y(_07029_));
 sg13g2_o21ai_1 _26031_ (.B1(_07029_),
    .Y(_07030_),
    .A1(_07023_),
    .A2(_07026_));
 sg13g2_and2_1 _26032_ (.A(_07021_),
    .B(_07030_),
    .X(_07031_));
 sg13g2_buf_2 _26033_ (.A(_07031_),
    .X(_07032_));
 sg13g2_mux2_1 _26034_ (.A0(\cpu.uart.r_ib[0] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(_07032_),
    .X(_02642_));
 sg13g2_mux2_1 _26035_ (.A0(\cpu.uart.r_ib[1] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(_07032_),
    .X(_02643_));
 sg13g2_mux2_1 _26036_ (.A0(\cpu.uart.r_ib[2] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(_07032_),
    .X(_02644_));
 sg13g2_mux2_1 _26037_ (.A0(\cpu.uart.r_ib[3] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(_07032_),
    .X(_02645_));
 sg13g2_mux2_1 _26038_ (.A0(\cpu.uart.r_ib[4] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(_07032_),
    .X(_02646_));
 sg13g2_mux2_1 _26039_ (.A0(\cpu.uart.r_ib[5] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(_07032_),
    .X(_02647_));
 sg13g2_xor2_1 _26040_ (.B(\cpu.uart.r_r ),
    .A(\cpu.uart.r_r_invert ),
    .X(_07033_));
 sg13g2_mux2_1 _26041_ (.A0(\cpu.uart.r_ib[6] ),
    .A1(_07033_),
    .S(_07032_),
    .X(_02648_));
 sg13g2_and4_1 _26042_ (.A(_07027_),
    .B(net937),
    .C(_07021_),
    .D(_07026_),
    .X(_07034_));
 sg13g2_buf_1 _26043_ (.A(_07034_),
    .X(_07035_));
 sg13g2_mux2_1 _26044_ (.A0(\cpu.uart.r_in[0] ),
    .A1(\cpu.uart.r_ib[0] ),
    .S(net178),
    .X(_02649_));
 sg13g2_mux2_1 _26045_ (.A0(\cpu.uart.r_in[1] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(net178),
    .X(_02650_));
 sg13g2_mux2_1 _26046_ (.A0(\cpu.uart.r_in[2] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(net178),
    .X(_02651_));
 sg13g2_mux2_1 _26047_ (.A0(\cpu.uart.r_in[3] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(net178),
    .X(_02652_));
 sg13g2_mux2_1 _26048_ (.A0(\cpu.uart.r_in[4] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(net178),
    .X(_02653_));
 sg13g2_mux2_1 _26049_ (.A0(\cpu.uart.r_in[5] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(net178),
    .X(_02654_));
 sg13g2_mux2_1 _26050_ (.A0(\cpu.uart.r_in[6] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(net178),
    .X(_02655_));
 sg13g2_mux2_1 _26051_ (.A0(\cpu.uart.r_in[7] ),
    .A1(_07033_),
    .S(_07035_),
    .X(_02656_));
 sg13g2_buf_1 _26052_ (.A(\cpu.uart.r_xstate[1] ),
    .X(_07036_));
 sg13g2_buf_1 _26053_ (.A(_07036_),
    .X(_07037_));
 sg13g2_buf_1 _26054_ (.A(\cpu.uart.r_xstate[0] ),
    .X(_07038_));
 sg13g2_buf_1 _26055_ (.A(_07038_),
    .X(_07039_));
 sg13g2_nor2_1 _26056_ (.A(net1043),
    .B(net1042),
    .Y(_07040_));
 sg13g2_and3_1 _26057_ (.X(_07041_),
    .A(net1030),
    .B(_07040_),
    .C(_06321_));
 sg13g2_buf_2 _26058_ (.A(_07041_),
    .X(_07042_));
 sg13g2_nand2_1 _26059_ (.Y(_07043_),
    .A(net391),
    .B(_07042_));
 sg13g2_buf_1 _26060_ (.A(\cpu.uart.r_xstate[3] ),
    .X(_07044_));
 sg13g2_buf_1 _26061_ (.A(_07044_),
    .X(_07045_));
 sg13g2_buf_1 _26062_ (.A(\cpu.uart.r_xstate[2] ),
    .X(_07046_));
 sg13g2_nor2_1 _26063_ (.A(net934),
    .B(_07046_),
    .Y(_07047_));
 sg13g2_o21ai_1 _26064_ (.B1(_07047_),
    .Y(_07048_),
    .A1(net935),
    .A2(_07043_));
 sg13g2_nand3_1 _26065_ (.B(net391),
    .C(_07042_),
    .A(_07039_),
    .Y(_07049_));
 sg13g2_nand3_1 _26066_ (.B(_07045_),
    .C(_07049_),
    .A(net936),
    .Y(_07050_));
 sg13g2_o21ai_1 _26067_ (.B1(_07050_),
    .Y(_07051_),
    .A1(net936),
    .A2(_07048_));
 sg13g2_buf_1 _26068_ (.A(_07046_),
    .X(_07052_));
 sg13g2_nor2_1 _26069_ (.A(_07037_),
    .B(_07046_),
    .Y(_07053_));
 sg13g2_xnor2_1 _26070_ (.Y(_07054_),
    .A(net934),
    .B(_07053_));
 sg13g2_buf_2 _26071_ (.A(_07054_),
    .X(_07055_));
 sg13g2_buf_1 _26072_ (.A(\cpu.uart.r_xcnt[0] ),
    .X(_07056_));
 sg13g2_nor2_1 _26073_ (.A(_07056_),
    .B(\cpu.uart.r_xcnt[1] ),
    .Y(_07057_));
 sg13g2_nand2_1 _26074_ (.Y(_07058_),
    .A(_09930_),
    .B(_07057_));
 sg13g2_buf_1 _26075_ (.A(_07058_),
    .X(_07059_));
 sg13g2_a221oi_1 _26076_ (.B2(_07059_),
    .C1(net899),
    .B1(_07055_),
    .A1(net934),
    .Y(_07060_),
    .A2(net933));
 sg13g2_nand2b_1 _26077_ (.Y(_07061_),
    .B(_07060_),
    .A_N(_07051_));
 sg13g2_buf_1 _26078_ (.A(_07061_),
    .X(_07062_));
 sg13g2_buf_1 _26079_ (.A(_07062_),
    .X(_07063_));
 sg13g2_buf_1 _26080_ (.A(_07055_),
    .X(_07064_));
 sg13g2_nor2b_1 _26081_ (.A(_07064_),
    .B_N(_10047_),
    .Y(_07065_));
 sg13g2_a21oi_1 _26082_ (.A1(\cpu.uart.r_out[1] ),
    .A2(net573),
    .Y(_07066_),
    .B1(_07065_));
 sg13g2_nand2_1 _26083_ (.Y(_07067_),
    .A(\cpu.uart.r_out[0] ),
    .B(net30));
 sg13g2_o21ai_1 _26084_ (.B1(_07067_),
    .Y(_02657_),
    .A1(_07063_),
    .A2(_07066_));
 sg13g2_nor2_1 _26085_ (.A(net887),
    .B(_07064_),
    .Y(_07068_));
 sg13g2_a21oi_1 _26086_ (.A1(\cpu.uart.r_out[2] ),
    .A2(net573),
    .Y(_07069_),
    .B1(_07068_));
 sg13g2_nand2_1 _26087_ (.Y(_07070_),
    .A(\cpu.uart.r_out[1] ),
    .B(_07063_));
 sg13g2_o21ai_1 _26088_ (.B1(_07070_),
    .Y(_02658_),
    .A1(net30),
    .A2(_07069_));
 sg13g2_nor2b_1 _26089_ (.A(_07055_),
    .B_N(net1020),
    .Y(_07071_));
 sg13g2_a21oi_1 _26090_ (.A1(\cpu.uart.r_out[3] ),
    .A2(net573),
    .Y(_07072_),
    .B1(_07071_));
 sg13g2_nand2_1 _26091_ (.Y(_07073_),
    .A(\cpu.uart.r_out[2] ),
    .B(_07062_));
 sg13g2_o21ai_1 _26092_ (.B1(_07073_),
    .Y(_02659_),
    .A1(net30),
    .A2(_07072_));
 sg13g2_nor2b_1 _26093_ (.A(_07055_),
    .B_N(net1113),
    .Y(_07074_));
 sg13g2_a21oi_1 _26094_ (.A1(\cpu.uart.r_out[4] ),
    .A2(net573),
    .Y(_07075_),
    .B1(_07074_));
 sg13g2_nand2_1 _26095_ (.Y(_07076_),
    .A(\cpu.uart.r_out[3] ),
    .B(_07062_));
 sg13g2_o21ai_1 _26096_ (.B1(_07076_),
    .Y(_02660_),
    .A1(net30),
    .A2(_07075_));
 sg13g2_nor2b_1 _26097_ (.A(_07055_),
    .B_N(_10085_),
    .Y(_07077_));
 sg13g2_a21oi_1 _26098_ (.A1(\cpu.uart.r_out[5] ),
    .A2(net573),
    .Y(_07078_),
    .B1(_07077_));
 sg13g2_nand2_1 _26099_ (.Y(_07079_),
    .A(\cpu.uart.r_out[4] ),
    .B(_07062_));
 sg13g2_o21ai_1 _26100_ (.B1(_07079_),
    .Y(_02661_),
    .A1(net30),
    .A2(_07078_));
 sg13g2_nor2b_1 _26101_ (.A(_07055_),
    .B_N(_10091_),
    .Y(_07080_));
 sg13g2_a21oi_1 _26102_ (.A1(\cpu.uart.r_out[6] ),
    .A2(net573),
    .Y(_07081_),
    .B1(_07080_));
 sg13g2_nand2_1 _26103_ (.Y(_07082_),
    .A(\cpu.uart.r_out[5] ),
    .B(_07062_));
 sg13g2_o21ai_1 _26104_ (.B1(_07082_),
    .Y(_02662_),
    .A1(net30),
    .A2(_07081_));
 sg13g2_nor2b_1 _26105_ (.A(_07055_),
    .B_N(_10097_),
    .Y(_07083_));
 sg13g2_a21oi_1 _26106_ (.A1(\cpu.uart.r_out[7] ),
    .A2(net573),
    .Y(_07084_),
    .B1(_07083_));
 sg13g2_nand2_1 _26107_ (.Y(_07085_),
    .A(\cpu.uart.r_out[6] ),
    .B(_07062_));
 sg13g2_o21ai_1 _26108_ (.B1(_07085_),
    .Y(_02663_),
    .A1(net30),
    .A2(_07084_));
 sg13g2_nor3_1 _26109_ (.A(_06974_),
    .B(net573),
    .C(_07062_),
    .Y(_07086_));
 sg13g2_a21o_1 _26110_ (.A2(net30),
    .A1(\cpu.uart.r_out[7] ),
    .B1(_07086_),
    .X(_02664_));
 sg13g2_nand2b_1 _26111_ (.Y(_07087_),
    .B(_09959_),
    .A_N(_09919_));
 sg13g2_buf_1 _26112_ (.A(_07087_),
    .X(_07088_));
 sg13g2_nor3_1 _26113_ (.A(net1079),
    .B(_07025_),
    .C(net1080),
    .Y(_07089_));
 sg13g2_a22oi_1 _26114_ (.Y(_07090_),
    .B1(_07088_),
    .B2(_07089_),
    .A2(net1080),
    .A1(net1079));
 sg13g2_nor4_1 _26115_ (.A(_07027_),
    .B(\cpu.uart.r_rstate[1] ),
    .C(_07025_),
    .D(net1080),
    .Y(_07091_));
 sg13g2_buf_1 _26116_ (.A(_07025_),
    .X(_07092_));
 sg13g2_a21o_1 _26117_ (.A2(_07088_),
    .A1(_07024_),
    .B1(net932),
    .X(_07093_));
 sg13g2_a22oi_1 _26118_ (.Y(_07094_),
    .B1(_07093_),
    .B2(net1080),
    .A2(_07091_),
    .A1(_07033_));
 sg13g2_o21ai_1 _26119_ (.B1(_07094_),
    .Y(_07095_),
    .A1(_07028_),
    .A2(_07090_));
 sg13g2_nor2_1 _26120_ (.A(_07028_),
    .B(net1079),
    .Y(_07096_));
 sg13g2_nor2b_1 _26121_ (.A(_07022_),
    .B_N(_07033_),
    .Y(_07097_));
 sg13g2_nand2_1 _26122_ (.Y(_07098_),
    .A(net1079),
    .B(net1080));
 sg13g2_nor2_1 _26123_ (.A(_07027_),
    .B(_07098_),
    .Y(_07099_));
 sg13g2_a21oi_1 _26124_ (.A1(_07096_),
    .A2(_07097_),
    .Y(_07100_),
    .B1(_07099_));
 sg13g2_nor3_1 _26125_ (.A(_07092_),
    .B(_07020_),
    .C(_07100_),
    .Y(_07101_));
 sg13g2_xor2_1 _26126_ (.B(_07026_),
    .A(net1080),
    .X(_07102_));
 sg13g2_o21ai_1 _26127_ (.B1(net891),
    .Y(_07103_),
    .A1(_09930_),
    .A2(_07102_));
 sg13g2_nor3_1 _26128_ (.A(_07095_),
    .B(_07101_),
    .C(_07103_),
    .Y(_07104_));
 sg13g2_and2_1 _26129_ (.A(_07027_),
    .B(net1079),
    .X(_07105_));
 sg13g2_buf_1 _26130_ (.A(_07105_),
    .X(_07106_));
 sg13g2_o21ai_1 _26131_ (.B1(net937),
    .Y(_07107_),
    .A1(net932),
    .A2(_07106_));
 sg13g2_nor2b_1 _26132_ (.A(_07091_),
    .B_N(_07107_),
    .Y(_07108_));
 sg13g2_and2_1 _26133_ (.A(_07104_),
    .B(_07108_),
    .X(_07109_));
 sg13g2_nor2_1 _26134_ (.A(_07018_),
    .B(_07104_),
    .Y(_07110_));
 sg13g2_a21oi_1 _26135_ (.A1(_07018_),
    .A2(_07109_),
    .Y(_02667_),
    .B1(_07110_));
 sg13g2_nand2_1 _26136_ (.Y(_07111_),
    .A(_07018_),
    .B(_07108_));
 sg13g2_nand2_1 _26137_ (.Y(_07112_),
    .A(_07104_),
    .B(_07111_));
 sg13g2_a22oi_1 _26138_ (.Y(_07113_),
    .B1(_07112_),
    .B2(\cpu.uart.r_rcnt[1] ),
    .A2(_07109_),
    .A1(_07019_));
 sg13g2_inv_1 _26139_ (.Y(_02668_),
    .A(_07113_));
 sg13g2_buf_1 _26140_ (.A(\cpu.gpio.genblk1[3].srcs_o[1] ),
    .X(_07114_));
 sg13g2_and2_1 _26141_ (.A(_07045_),
    .B(_07052_),
    .X(_07115_));
 sg13g2_buf_1 _26142_ (.A(_07115_),
    .X(_07116_));
 sg13g2_nor2_2 _26143_ (.A(_07036_),
    .B(_07038_),
    .Y(_07117_));
 sg13g2_o21ai_1 _26144_ (.B1(_07117_),
    .Y(_07118_),
    .A1(_07047_),
    .A2(_07116_));
 sg13g2_nand3b_1 _26145_ (.B(net934),
    .C(net936),
    .Y(_07119_),
    .A_N(_07052_));
 sg13g2_buf_1 _26146_ (.A(_07119_),
    .X(_07120_));
 sg13g2_nand3_1 _26147_ (.B(_07118_),
    .C(_07120_),
    .A(net891),
    .Y(_07121_));
 sg13g2_nand2_1 _26148_ (.Y(_07122_),
    .A(\cpu.uart.r_out[0] ),
    .B(_07055_));
 sg13g2_xor2_1 _26149_ (.B(_07122_),
    .A(\cpu.uart.r_x_invert ),
    .X(_07123_));
 sg13g2_nand2_1 _26150_ (.Y(_07124_),
    .A(_00278_),
    .B(_07121_));
 sg13g2_o21ai_1 _26151_ (.B1(_07124_),
    .Y(_07125_),
    .A1(_07121_),
    .A2(_07123_));
 sg13g2_inv_1 _26152_ (.Y(_07126_),
    .A(_07044_));
 sg13g2_nand2_1 _26153_ (.Y(_07127_),
    .A(net936),
    .B(net935));
 sg13g2_nor4_2 _26154_ (.A(_07126_),
    .B(net933),
    .C(_07043_),
    .Y(_07128_),
    .D(_07127_));
 sg13g2_nand2_1 _26155_ (.Y(_07129_),
    .A(_07038_),
    .B(net934));
 sg13g2_nand3_1 _26156_ (.B(_07059_),
    .C(_07129_),
    .A(_07037_),
    .Y(_07130_));
 sg13g2_nor2_1 _26157_ (.A(_07044_),
    .B(_07059_),
    .Y(_07131_));
 sg13g2_a21oi_1 _26158_ (.A1(net934),
    .A2(_07117_),
    .Y(_07132_),
    .B1(_07131_));
 sg13g2_nor2b_1 _26159_ (.A(_07044_),
    .B_N(_07038_),
    .Y(_07133_));
 sg13g2_a21oi_1 _26160_ (.A1(_09930_),
    .A2(_07057_),
    .Y(_07134_),
    .B1(_07126_));
 sg13g2_a21oi_1 _26161_ (.A1(_07088_),
    .A2(_07133_),
    .Y(_07135_),
    .B1(_07134_));
 sg13g2_nor2b_1 _26162_ (.A(_07135_),
    .B_N(_07053_),
    .Y(_07136_));
 sg13g2_a21oi_1 _26163_ (.A1(_07046_),
    .A2(_07132_),
    .Y(_07137_),
    .B1(_07136_));
 sg13g2_nand2_1 _26164_ (.Y(_07138_),
    .A(_07130_),
    .B(_07137_));
 sg13g2_o21ai_1 _26165_ (.B1(net891),
    .Y(_07139_),
    .A1(_07128_),
    .A2(_07138_));
 sg13g2_mux2_1 _26166_ (.A0(_07114_),
    .A1(_07125_),
    .S(_07139_),
    .X(_02673_));
 sg13g2_a21o_1 _26167_ (.A2(_07057_),
    .A1(net935),
    .B1(net933),
    .X(_07140_));
 sg13g2_or2_1 _26168_ (.X(_07141_),
    .B(_07057_),
    .A(net935));
 sg13g2_a22oi_1 _26169_ (.Y(_07142_),
    .B1(_07141_),
    .B2(net933),
    .A2(_07140_),
    .A1(net936));
 sg13g2_and2_1 _26170_ (.A(_07047_),
    .B(_07117_),
    .X(_07143_));
 sg13g2_buf_1 _26171_ (.A(_07143_),
    .X(_07144_));
 sg13g2_nor2_1 _26172_ (.A(net899),
    .B(_07144_),
    .Y(_07145_));
 sg13g2_o21ai_1 _26173_ (.B1(_07145_),
    .Y(_07146_),
    .A1(_07126_),
    .A2(_07142_));
 sg13g2_nor3_1 _26174_ (.A(_07088_),
    .B(_07128_),
    .C(_07146_),
    .Y(_07147_));
 sg13g2_inv_1 _26175_ (.Y(_07148_),
    .A(_07117_));
 sg13g2_a22oi_1 _26176_ (.Y(_07149_),
    .B1(_07148_),
    .B2(_07116_),
    .A2(_07053_),
    .A1(_07126_));
 sg13g2_nand2_1 _26177_ (.Y(_07150_),
    .A(_07147_),
    .B(_07149_));
 sg13g2_nor2b_1 _26178_ (.A(_07056_),
    .B_N(_07147_),
    .Y(_07151_));
 sg13g2_a21oi_1 _26179_ (.A1(_07056_),
    .A2(_07150_),
    .Y(_07152_),
    .B1(_07151_));
 sg13g2_inv_1 _26180_ (.Y(_02676_),
    .A(_07152_));
 sg13g2_nand2_1 _26181_ (.Y(_07153_),
    .A(_07056_),
    .B(_07149_));
 sg13g2_nand2_1 _26182_ (.Y(_07154_),
    .A(_07147_),
    .B(_07153_));
 sg13g2_o21ai_1 _26183_ (.B1(\cpu.uart.r_xcnt[1] ),
    .Y(_07155_),
    .A1(_07056_),
    .A2(_07150_));
 sg13g2_o21ai_1 _26184_ (.B1(_07155_),
    .Y(_02677_),
    .A1(\cpu.uart.r_xcnt[1] ),
    .A2(_07154_));
 sg13g2_buf_1 _26185_ (.A(_10117_),
    .X(_07156_));
 sg13g2_buf_1 _26186_ (.A(net80),
    .X(_07157_));
 sg13g2_buf_1 _26187_ (.A(_10126_),
    .X(_07158_));
 sg13g2_inv_1 _26188_ (.Y(_07159_),
    .A(_04972_));
 sg13g2_nand2_1 _26189_ (.Y(_07160_),
    .A(_10210_),
    .B(_10212_));
 sg13g2_nand2_1 _26190_ (.Y(_07161_),
    .A(_10217_),
    .B(_10167_));
 sg13g2_nor3_2 _26191_ (.A(_07159_),
    .B(_07160_),
    .C(_07161_),
    .Y(_07162_));
 sg13g2_nand2_1 _26192_ (.Y(_07163_),
    .A(net91),
    .B(_07162_));
 sg13g2_o21ai_1 _26193_ (.B1(_07163_),
    .Y(_07164_),
    .A1(net1029),
    .A2(net102));
 sg13g2_nor2_1 _26194_ (.A(_07160_),
    .B(_07161_),
    .Y(_07165_));
 sg13g2_o21ai_1 _26195_ (.B1(net87),
    .Y(_07166_),
    .A1(_10141_),
    .A2(_07165_));
 sg13g2_a22oi_1 _26196_ (.Y(_02463_),
    .B1(_07166_),
    .B2(_07159_),
    .A2(_07164_),
    .A1(net71));
 sg13g2_and2_1 _26197_ (.A(_05352_),
    .B(_07162_),
    .X(_07167_));
 sg13g2_buf_1 _26198_ (.A(_07167_),
    .X(_07168_));
 sg13g2_nand2_1 _26199_ (.Y(_07169_),
    .A(net91),
    .B(_07168_));
 sg13g2_o21ai_1 _26200_ (.B1(_07169_),
    .Y(_07170_),
    .A1(net1027),
    .A2(_10127_));
 sg13g2_o21ai_1 _26201_ (.B1(net87),
    .Y(_07171_),
    .A1(net86),
    .A2(_07162_));
 sg13g2_inv_1 _26202_ (.Y(_07172_),
    .A(_05352_));
 sg13g2_a22oi_1 _26203_ (.Y(_02464_),
    .B1(_07171_),
    .B2(_07172_),
    .A2(_07170_),
    .A1(net71));
 sg13g2_nand3_1 _26204_ (.B(_07158_),
    .C(_07168_),
    .A(_05461_),
    .Y(_07173_));
 sg13g2_o21ai_1 _26205_ (.B1(_07173_),
    .Y(_07174_),
    .A1(net1026),
    .A2(_10127_));
 sg13g2_o21ai_1 _26206_ (.B1(_07156_),
    .Y(_07175_),
    .A1(_10141_),
    .A2(_07168_));
 sg13g2_inv_1 _26207_ (.Y(_07176_),
    .A(_05461_));
 sg13g2_a22oi_1 _26208_ (.Y(_02465_),
    .B1(_07175_),
    .B2(_07176_),
    .A2(_07174_),
    .A1(_07157_));
 sg13g2_buf_1 _26209_ (.A(_10126_),
    .X(_07177_));
 sg13g2_nand4_1 _26210_ (.B(_04972_),
    .C(_05352_),
    .A(_10217_),
    .Y(_07178_),
    .D(_05461_));
 sg13g2_nor2_2 _26211_ (.A(_10218_),
    .B(_07178_),
    .Y(_07179_));
 sg13g2_nand3_1 _26212_ (.B(_07158_),
    .C(_07179_),
    .A(_05531_),
    .Y(_07180_));
 sg13g2_o21ai_1 _26213_ (.B1(_07180_),
    .Y(_07181_),
    .A1(net1025),
    .A2(_07177_));
 sg13g2_o21ai_1 _26214_ (.B1(_07156_),
    .Y(_07182_),
    .A1(net86),
    .A2(_07179_));
 sg13g2_inv_1 _26215_ (.Y(_07183_),
    .A(_05531_));
 sg13g2_a22oi_1 _26216_ (.Y(_02466_),
    .B1(_07182_),
    .B2(_07183_),
    .A2(_07181_),
    .A1(net71));
 sg13g2_nand3_1 _26217_ (.B(_05531_),
    .C(_07168_),
    .A(_05461_),
    .Y(_07184_));
 sg13g2_nor3_1 _26218_ (.A(_05558_),
    .B(_10140_),
    .C(_07184_),
    .Y(_07185_));
 sg13g2_a21oi_1 _26219_ (.A1(net1024),
    .A2(net100),
    .Y(_07186_),
    .B1(_07185_));
 sg13g2_a21oi_1 _26220_ (.A1(net91),
    .A2(_07184_),
    .Y(_07187_),
    .B1(_10136_));
 sg13g2_nand2b_1 _26221_ (.Y(_07188_),
    .B(_05558_),
    .A_N(_07187_));
 sg13g2_o21ai_1 _26222_ (.B1(_07188_),
    .Y(_02467_),
    .A1(net101),
    .A2(_07186_));
 sg13g2_and2_1 _26223_ (.A(_05531_),
    .B(_05558_),
    .X(_07189_));
 sg13g2_buf_1 _26224_ (.A(_07189_),
    .X(_07190_));
 sg13g2_nand4_1 _26225_ (.B(_10126_),
    .C(_07179_),
    .A(_05621_),
    .Y(_07191_),
    .D(_07190_));
 sg13g2_o21ai_1 _26226_ (.B1(_07191_),
    .Y(_07192_),
    .A1(net1023),
    .A2(net102));
 sg13g2_nand2_1 _26227_ (.Y(_07193_),
    .A(_07179_),
    .B(_07190_));
 sg13g2_a21oi_1 _26228_ (.A1(_07177_),
    .A2(_07193_),
    .Y(_07194_),
    .B1(net116));
 sg13g2_nor2_1 _26229_ (.A(_05621_),
    .B(_07194_),
    .Y(_07195_));
 sg13g2_a21oi_1 _26230_ (.A1(_07157_),
    .A2(_07192_),
    .Y(_02468_),
    .B1(_07195_));
 sg13g2_inv_1 _26231_ (.Y(_07196_),
    .A(_05737_));
 sg13g2_nand3_1 _26232_ (.B(_05461_),
    .C(_07162_),
    .A(_05352_),
    .Y(_07197_));
 sg13g2_nand2_1 _26233_ (.Y(_07198_),
    .A(_05621_),
    .B(_07190_));
 sg13g2_nor3_2 _26234_ (.A(_07196_),
    .B(_07197_),
    .C(_07198_),
    .Y(_07199_));
 sg13g2_nand2_1 _26235_ (.Y(_07200_),
    .A(net91),
    .B(_07199_));
 sg13g2_o21ai_1 _26236_ (.B1(_07200_),
    .Y(_07201_),
    .A1(net1022),
    .A2(net90));
 sg13g2_nor2_1 _26237_ (.A(_07197_),
    .B(_07198_),
    .Y(_07202_));
 sg13g2_o21ai_1 _26238_ (.B1(net80),
    .Y(_07203_),
    .A1(net86),
    .A2(_07202_));
 sg13g2_a22oi_1 _26239_ (.Y(_02469_),
    .B1(_07203_),
    .B2(_07196_),
    .A2(_07201_),
    .A1(net87));
 sg13g2_nand4_1 _26240_ (.B(_05737_),
    .C(_07179_),
    .A(_05621_),
    .Y(_07204_),
    .D(_07190_));
 sg13g2_buf_1 _26241_ (.A(_07204_),
    .X(_07205_));
 sg13g2_nor2_1 _26242_ (.A(net100),
    .B(_07205_),
    .Y(_07206_));
 sg13g2_nand2_1 _26243_ (.Y(_07207_),
    .A(_05111_),
    .B(_07206_));
 sg13g2_o21ai_1 _26244_ (.B1(_07207_),
    .Y(_07208_),
    .A1(net1021),
    .A2(net102));
 sg13g2_a21oi_1 _26245_ (.A1(net90),
    .A2(_07205_),
    .Y(_07209_),
    .B1(net116));
 sg13g2_nor2_1 _26246_ (.A(_05111_),
    .B(_07209_),
    .Y(_07210_));
 sg13g2_a21oi_1 _26247_ (.A1(net71),
    .A2(_07208_),
    .Y(_02470_),
    .B1(_07210_));
 sg13g2_nand3_1 _26248_ (.B(_05761_),
    .C(_07199_),
    .A(_05111_),
    .Y(_07211_));
 sg13g2_buf_1 _26249_ (.A(_07211_),
    .X(_07212_));
 sg13g2_nor2_1 _26250_ (.A(_10139_),
    .B(_07212_),
    .Y(_07213_));
 sg13g2_inv_1 _26251_ (.Y(_07214_),
    .A(_07213_));
 sg13g2_o21ai_1 _26252_ (.B1(_07214_),
    .Y(_07215_),
    .A1(_10181_),
    .A2(net102));
 sg13g2_a21o_1 _26253_ (.A2(_07199_),
    .A1(_05111_),
    .B1(net100),
    .X(_07216_));
 sg13g2_a21oi_1 _26254_ (.A1(net80),
    .A2(_07216_),
    .Y(_07217_),
    .B1(_05761_));
 sg13g2_a21oi_1 _26255_ (.A1(net71),
    .A2(_07215_),
    .Y(_02471_),
    .B1(_07217_));
 sg13g2_nand2_1 _26256_ (.Y(_07218_),
    .A(_05775_),
    .B(_07213_));
 sg13g2_o21ai_1 _26257_ (.B1(_07218_),
    .Y(_07219_),
    .A1(_10186_),
    .A2(net90));
 sg13g2_a21o_1 _26258_ (.A2(_07212_),
    .A1(net90),
    .B1(net101),
    .X(_07220_));
 sg13g2_inv_1 _26259_ (.Y(_07221_),
    .A(_05775_));
 sg13g2_a22oi_1 _26260_ (.Y(_02472_),
    .B1(_07220_),
    .B2(_07221_),
    .A2(_07219_),
    .A1(net87));
 sg13g2_and2_1 _26261_ (.A(_05775_),
    .B(_05177_),
    .X(_07222_));
 sg13g2_buf_1 _26262_ (.A(_07222_),
    .X(_07223_));
 sg13g2_nand2_1 _26263_ (.Y(_07224_),
    .A(_07213_),
    .B(_07223_));
 sg13g2_o21ai_1 _26264_ (.B1(_07224_),
    .Y(_07225_),
    .A1(_10191_),
    .A2(net102));
 sg13g2_o21ai_1 _26265_ (.B1(net91),
    .Y(_07226_),
    .A1(_07221_),
    .A2(_07212_));
 sg13g2_a21oi_1 _26266_ (.A1(net80),
    .A2(_07226_),
    .Y(_07227_),
    .B1(_05177_));
 sg13g2_a21oi_1 _26267_ (.A1(net71),
    .A2(_07225_),
    .Y(_02473_),
    .B1(_07227_));
 sg13g2_inv_1 _26268_ (.Y(_07228_),
    .A(_05218_));
 sg13g2_nand3_1 _26269_ (.B(_05761_),
    .C(_07223_),
    .A(_05111_),
    .Y(_07229_));
 sg13g2_nor2_1 _26270_ (.A(_07228_),
    .B(_07229_),
    .Y(_07230_));
 sg13g2_nand2_1 _26271_ (.Y(_07231_),
    .A(_07206_),
    .B(_07230_));
 sg13g2_o21ai_1 _26272_ (.B1(_07231_),
    .Y(_07232_),
    .A1(_10198_),
    .A2(net90));
 sg13g2_o21ai_1 _26273_ (.B1(net90),
    .Y(_07233_),
    .A1(_07205_),
    .A2(_07229_));
 sg13g2_nand2_1 _26274_ (.Y(_07234_),
    .A(net87),
    .B(_07233_));
 sg13g2_a22oi_1 _26275_ (.Y(_02474_),
    .B1(_07234_),
    .B2(_07228_),
    .A2(_07232_),
    .A1(net87));
 sg13g2_nand4_1 _26276_ (.B(_10126_),
    .C(_07199_),
    .A(_05233_),
    .Y(_07235_),
    .D(_07230_));
 sg13g2_o21ai_1 _26277_ (.B1(_07235_),
    .Y(_07236_),
    .A1(_10203_),
    .A2(net102));
 sg13g2_a21o_1 _26278_ (.A2(_07230_),
    .A1(_07199_),
    .B1(net100),
    .X(_07237_));
 sg13g2_a21oi_1 _26279_ (.A1(net80),
    .A2(_07237_),
    .Y(_07238_),
    .B1(_05233_));
 sg13g2_a21oi_1 _26280_ (.A1(net71),
    .A2(_07236_),
    .Y(_02475_),
    .B1(_07238_));
 sg13g2_nand2_1 _26281_ (.Y(_07239_),
    .A(_05233_),
    .B(_07230_));
 sg13g2_nor2_1 _26282_ (.A(_07205_),
    .B(_07239_),
    .Y(_07240_));
 sg13g2_nand3_1 _26283_ (.B(net91),
    .C(_07240_),
    .A(_05275_),
    .Y(_07241_));
 sg13g2_o21ai_1 _26284_ (.B1(_07241_),
    .Y(_07242_),
    .A1(_10205_),
    .A2(net90));
 sg13g2_o21ai_1 _26285_ (.B1(net80),
    .Y(_07243_),
    .A1(net86),
    .A2(_07240_));
 sg13g2_inv_1 _26286_ (.Y(_07244_),
    .A(_05275_));
 sg13g2_a22oi_1 _26287_ (.Y(_02476_),
    .B1(_07243_),
    .B2(_07244_),
    .A2(_07242_),
    .A1(net87));
 sg13g2_inv_1 _26288_ (.Y(_07245_),
    .A(_05286_));
 sg13g2_nand4_1 _26289_ (.B(_05233_),
    .C(_05275_),
    .A(_05218_),
    .Y(_07246_),
    .D(_07223_));
 sg13g2_buf_1 _26290_ (.A(_07246_),
    .X(_07247_));
 sg13g2_or3_1 _26291_ (.A(_07245_),
    .B(_07214_),
    .C(_07247_),
    .X(_07248_));
 sg13g2_o21ai_1 _26292_ (.B1(_07248_),
    .Y(_07249_),
    .A1(_10215_),
    .A2(net102));
 sg13g2_o21ai_1 _26293_ (.B1(net91),
    .Y(_07250_),
    .A1(_07212_),
    .A2(_07247_));
 sg13g2_a21oi_1 _26294_ (.A1(net80),
    .A2(_07250_),
    .Y(_07251_),
    .B1(_05286_));
 sg13g2_a21oi_1 _26295_ (.A1(net71),
    .A2(_07249_),
    .Y(_02477_),
    .B1(_07251_));
 sg13g2_nand3_1 _26296_ (.B(_05761_),
    .C(_05286_),
    .A(_05111_),
    .Y(_07252_));
 sg13g2_nor3_1 _26297_ (.A(_07205_),
    .B(_07247_),
    .C(_07252_),
    .Y(_07253_));
 sg13g2_nand3_1 _26298_ (.B(net91),
    .C(_07253_),
    .A(_05318_),
    .Y(_07254_));
 sg13g2_o21ai_1 _26299_ (.B1(_07254_),
    .Y(_07255_),
    .A1(_10220_),
    .A2(net90));
 sg13g2_o21ai_1 _26300_ (.B1(net80),
    .Y(_07256_),
    .A1(net86),
    .A2(_07253_));
 sg13g2_inv_1 _26301_ (.Y(_07257_),
    .A(_05318_));
 sg13g2_a22oi_1 _26302_ (.Y(_02478_),
    .B1(_07256_),
    .B2(_07257_),
    .A2(_07255_),
    .A1(net87));
 sg13g2_nor2_1 _26303_ (.A(\cpu.r_clk_invert ),
    .B(net618),
    .Y(_07258_));
 sg13g2_a21oi_1 _26304_ (.A1(_09217_),
    .A2(net629),
    .Y(_02545_),
    .B1(_07258_));
 sg13g2_nand2b_1 _26305_ (.Y(_07259_),
    .B(net891),
    .A_N(\cpu.d_flush_all ));
 sg13g2_buf_2 _26306_ (.A(_07259_),
    .X(_07260_));
 sg13g2_nor2b_1 _26307_ (.A(\cpu.dcache.r_valid[0] ),
    .B_N(net469),
    .Y(_07261_));
 sg13g2_nand3_1 _26308_ (.B(_02953_),
    .C(_02958_),
    .A(_09391_),
    .Y(_07262_));
 sg13g2_buf_2 _26309_ (.A(_07262_),
    .X(_07263_));
 sg13g2_nor2_1 _26310_ (.A(net603),
    .B(_07263_),
    .Y(_07264_));
 sg13g2_nor3_1 _26311_ (.A(_07260_),
    .B(_07261_),
    .C(_07264_),
    .Y(_00739_));
 sg13g2_nor2_1 _26312_ (.A(\cpu.dcache.r_valid[1] ),
    .B(net464),
    .Y(_07265_));
 sg13g2_nor2_1 _26313_ (.A(net601),
    .B(_07263_),
    .Y(_07266_));
 sg13g2_nor3_1 _26314_ (.A(_07260_),
    .B(_07265_),
    .C(_07266_),
    .Y(_00740_));
 sg13g2_nor2_1 _26315_ (.A(\cpu.dcache.r_valid[2] ),
    .B(net333),
    .Y(_07267_));
 sg13g2_nor2_1 _26316_ (.A(net407),
    .B(_07263_),
    .Y(_07268_));
 sg13g2_nor3_1 _26317_ (.A(_07260_),
    .B(_07267_),
    .C(_07268_),
    .Y(_00741_));
 sg13g2_nor2_1 _26318_ (.A(\cpu.dcache.r_valid[3] ),
    .B(net402),
    .Y(_07269_));
 sg13g2_nor2_1 _26319_ (.A(net528),
    .B(_07263_),
    .Y(_07270_));
 sg13g2_nor3_1 _26320_ (.A(_07260_),
    .B(_07269_),
    .C(_07270_),
    .Y(_00742_));
 sg13g2_inv_1 _26321_ (.Y(_07271_),
    .A(\cpu.dcache.r_valid[4] ));
 sg13g2_inv_1 _26322_ (.Y(_07272_),
    .A(_07263_));
 sg13g2_a221oi_1 _26323_ (.B2(_04989_),
    .C1(_07260_),
    .B1(_07272_),
    .A1(_07271_),
    .Y(_00743_),
    .A2(net463));
 sg13g2_nor2_1 _26324_ (.A(\cpu.dcache.r_valid[5] ),
    .B(net460),
    .Y(_07273_));
 sg13g2_nor2_1 _26325_ (.A(net599),
    .B(_07263_),
    .Y(_07274_));
 sg13g2_nor3_1 _26326_ (.A(_07260_),
    .B(_07273_),
    .C(_07274_),
    .Y(_00744_));
 sg13g2_nor2_1 _26327_ (.A(\cpu.dcache.r_valid[6] ),
    .B(net400),
    .Y(_07275_));
 sg13g2_nor2_1 _26328_ (.A(net525),
    .B(_07263_),
    .Y(_07276_));
 sg13g2_nor3_1 _26329_ (.A(_07260_),
    .B(_07275_),
    .C(_07276_),
    .Y(_00745_));
 sg13g2_nor2_1 _26330_ (.A(\cpu.dcache.r_valid[7] ),
    .B(net365),
    .Y(_07277_));
 sg13g2_nor2_1 _26331_ (.A(net466),
    .B(_07263_),
    .Y(_07278_));
 sg13g2_nor3_1 _26332_ (.A(_07260_),
    .B(_07277_),
    .C(_07278_),
    .Y(_00746_));
 sg13g2_nor3_1 _26333_ (.A(net1019),
    .B(net1018),
    .C(_10228_),
    .Y(_07279_));
 sg13g2_nand2_1 _26334_ (.Y(_07280_),
    .A(_04816_),
    .B(_07279_));
 sg13g2_buf_1 _26335_ (.A(_07280_),
    .X(_07281_));
 sg13g2_nor2_1 _26336_ (.A(net650),
    .B(_07281_),
    .Y(_07282_));
 sg13g2_a21oi_1 _26337_ (.A1(_08475_),
    .A2(_07281_),
    .Y(_07283_),
    .B1(_07282_));
 sg13g2_nor3_1 _26338_ (.A(net294),
    .B(_09353_),
    .C(_07283_),
    .Y(_00795_));
 sg13g2_and4_1 _26339_ (.A(net721),
    .B(_11008_),
    .C(\cpu.dec.do_flush_all ),
    .D(net658),
    .X(_00928_));
 sg13g2_and4_1 _26340_ (.A(net721),
    .B(_10520_),
    .C(\cpu.dec.do_flush_all ),
    .D(net658),
    .X(_00946_));
 sg13g2_nand2_1 _26341_ (.Y(_07284_),
    .A(_04260_),
    .B(_10743_));
 sg13g2_a22oi_1 _26342_ (.Y(_07285_),
    .B1(_07284_),
    .B2(net330),
    .A2(_09365_),
    .A1(_06768_));
 sg13g2_nor2b_1 _26343_ (.A(_11524_),
    .B_N(_10628_),
    .Y(_07286_));
 sg13g2_nand3_1 _26344_ (.B(net658),
    .C(_07286_),
    .A(net721),
    .Y(_07287_));
 sg13g2_mux2_1 _26345_ (.A0(_10526_),
    .A1(_09257_),
    .S(_07287_),
    .X(_07288_));
 sg13g2_nor2_1 _26346_ (.A(_10749_),
    .B(net572),
    .Y(_07289_));
 sg13g2_a21oi_1 _26347_ (.A1(net572),
    .A2(_07288_),
    .Y(_07290_),
    .B1(_07289_));
 sg13g2_nor3_1 _26348_ (.A(net618),
    .B(_07285_),
    .C(_07290_),
    .Y(_00947_));
 sg13g2_nor4_1 _26349_ (.A(_09210_),
    .B(_00296_),
    .C(_04857_),
    .D(_04881_),
    .Y(_07291_));
 sg13g2_nand2_1 _26350_ (.Y(_07292_),
    .A(_08468_),
    .B(net658));
 sg13g2_nor2_1 _26351_ (.A(_00308_),
    .B(_07292_),
    .Y(_07293_));
 sg13g2_nand3b_1 _26352_ (.B(net1058),
    .C(net891),
    .Y(_07294_),
    .A_N(_12009_));
 sg13g2_a21oi_1 _26353_ (.A1(_09827_),
    .A2(_07294_),
    .Y(_07295_),
    .B1(_08468_));
 sg13g2_nor2_1 _26354_ (.A(_09294_),
    .B(_07295_),
    .Y(_07296_));
 sg13g2_o21ai_1 _26355_ (.B1(_07296_),
    .Y(_07297_),
    .A1(_09210_),
    .A2(_07293_));
 sg13g2_nor2_1 _26356_ (.A(_07291_),
    .B(_07297_),
    .Y(_01066_));
 sg13g2_nand2b_1 _26357_ (.Y(_07298_),
    .B(_07293_),
    .A_N(_04881_));
 sg13g2_a22oi_1 _26358_ (.Y(_07299_),
    .B1(_07293_),
    .B2(_11527_),
    .A2(_07296_),
    .A1(_08466_));
 sg13g2_o21ai_1 _26359_ (.B1(_07299_),
    .Y(_01067_),
    .A1(_04857_),
    .A2(_07298_));
 sg13g2_inv_1 _26360_ (.Y(_07300_),
    .A(\cpu.icache.r_valid[0] ));
 sg13g2_nand2b_1 _26361_ (.Y(_07301_),
    .B(_09877_),
    .A_N(\cpu.ex.i_flush_all ));
 sg13g2_buf_2 _26362_ (.A(_07301_),
    .X(_07302_));
 sg13g2_a21oi_1 _26363_ (.A1(_07300_),
    .A2(net353),
    .Y(_02422_),
    .B1(_07302_));
 sg13g2_nor2_1 _26364_ (.A(\cpu.icache.r_valid[1] ),
    .B(_06414_),
    .Y(_07303_));
 sg13g2_nor2_1 _26365_ (.A(_07302_),
    .B(_07303_),
    .Y(_02423_));
 sg13g2_nor2_1 _26366_ (.A(\cpu.icache.r_valid[2] ),
    .B(_06430_),
    .Y(_07304_));
 sg13g2_nor2_1 _26367_ (.A(_07302_),
    .B(_07304_),
    .Y(_02424_));
 sg13g2_inv_1 _26368_ (.Y(_07305_),
    .A(\cpu.icache.r_valid[3] ));
 sg13g2_a21oi_1 _26369_ (.A1(_07305_),
    .A2(net224),
    .Y(_02425_),
    .B1(_07302_));
 sg13g2_nor2_1 _26370_ (.A(\cpu.icache.r_valid[4] ),
    .B(_06461_),
    .Y(_07306_));
 sg13g2_nor2_1 _26371_ (.A(_07302_),
    .B(_07306_),
    .Y(_02426_));
 sg13g2_inv_1 _26372_ (.Y(_07307_),
    .A(\cpu.icache.r_valid[5] ));
 sg13g2_a21oi_1 _26373_ (.A1(_07307_),
    .A2(_06474_),
    .Y(_02427_),
    .B1(_07302_));
 sg13g2_inv_1 _26374_ (.Y(_07308_),
    .A(\cpu.icache.r_valid[6] ));
 sg13g2_a21oi_1 _26375_ (.A1(_07308_),
    .A2(_06483_),
    .Y(_02428_),
    .B1(_07302_));
 sg13g2_nor2_1 _26376_ (.A(\cpu.icache.r_valid[7] ),
    .B(_06497_),
    .Y(_07309_));
 sg13g2_nor2_1 _26377_ (.A(_07302_),
    .B(_07309_),
    .Y(_02429_));
 sg13g2_nand3_1 _26378_ (.B(net171),
    .C(_05435_),
    .A(net1113),
    .Y(_07310_));
 sg13g2_nand2_1 _26379_ (.Y(_07311_),
    .A(\cpu.intr.r_swi ),
    .B(_07310_));
 sg13g2_nand3_1 _26380_ (.B(net171),
    .C(_05436_),
    .A(net1025),
    .Y(_07312_));
 sg13g2_a21oi_1 _26381_ (.A1(_07311_),
    .A2(_07312_),
    .Y(_00315_),
    .B1(net574));
 sg13g2_nor2_1 _26382_ (.A(_02953_),
    .B(net1094),
    .Y(_07313_));
 sg13g2_nor2b_1 _26383_ (.A(_07313_),
    .B_N(_00313_),
    .Y(_00584_));
 sg13g2_nor2_1 _26384_ (.A(_12030_),
    .B(_12074_),
    .Y(_07314_));
 sg13g2_nor2_1 _26385_ (.A(_07313_),
    .B(_07314_),
    .Y(_00585_));
 sg13g2_xnor2_1 _26386_ (.Y(_07315_),
    .A(net999),
    .B(_12007_));
 sg13g2_nor2b_1 _26387_ (.A(_07313_),
    .B_N(_07315_),
    .Y(_00586_));
 sg13g2_nor2_1 _26388_ (.A(_09342_),
    .B(net572),
    .Y(_07316_));
 sg13g2_a21oi_1 _26389_ (.A1(net1057),
    .A2(net572),
    .Y(_07317_),
    .B1(_07316_));
 sg13g2_nor2_1 _26390_ (.A(net631),
    .B(_07317_),
    .Y(_00796_));
 sg13g2_a21oi_2 _26391_ (.B1(net226),
    .Y(_07318_),
    .A2(_04252_),
    .A1(_11522_));
 sg13g2_nor2b_1 _26392_ (.A(net721),
    .B_N(_07318_),
    .Y(_07319_));
 sg13g2_nand3b_1 _26393_ (.B(_04260_),
    .C(_07286_),
    .Y(_07320_),
    .A_N(_10762_));
 sg13g2_a21oi_1 _26394_ (.A1(net721),
    .A2(_07320_),
    .Y(_07321_),
    .B1(_09293_));
 sg13g2_nor2_1 _26395_ (.A(_03848_),
    .B(_07321_),
    .Y(_07322_));
 sg13g2_nor2_1 _26396_ (.A(_10762_),
    .B(_07322_),
    .Y(_07323_));
 sg13g2_a21oi_1 _26397_ (.A1(_10749_),
    .A2(_07322_),
    .Y(_07324_),
    .B1(_07323_));
 sg13g2_nor2_1 _26398_ (.A(_07318_),
    .B(_07324_),
    .Y(_07325_));
 sg13g2_o21ai_1 _26399_ (.B1(_09879_),
    .Y(_00797_),
    .A1(_07319_),
    .A2(_07325_));
 sg13g2_nand2_1 _26400_ (.Y(_07326_),
    .A(_10969_),
    .B(net572));
 sg13g2_o21ai_1 _26401_ (.B1(_07326_),
    .Y(_07327_),
    .A1(_02979_),
    .A2(net572));
 sg13g2_and2_1 _26402_ (.A(_06729_),
    .B(_07327_),
    .X(_00798_));
 sg13g2_nor4_1 _26403_ (.A(\cpu.ex.r_branch_stall ),
    .B(_11521_),
    .C(\cpu.dec.r_store ),
    .D(_07292_),
    .Y(_07328_));
 sg13g2_nor3_1 _26404_ (.A(_11517_),
    .B(_07295_),
    .C(_07328_),
    .Y(_07329_));
 sg13g2_nand2_1 _26405_ (.Y(_07330_),
    .A(_08580_),
    .B(_11523_));
 sg13g2_o21ai_1 _26406_ (.B1(net77),
    .Y(_07331_),
    .A1(_07329_),
    .A2(_07330_));
 sg13g2_nand2_1 _26407_ (.Y(_07332_),
    .A(_06779_),
    .B(_09014_));
 sg13g2_o21ai_1 _26408_ (.B1(_07332_),
    .Y(_07333_),
    .A1(_06779_),
    .A2(_07331_));
 sg13g2_nand2_1 _26409_ (.Y(_00944_),
    .A(_09879_),
    .B(_07333_));
 sg13g2_nand2_1 _26410_ (.Y(_07334_),
    .A(_09391_),
    .B(net1036));
 sg13g2_nand3_1 _26411_ (.B(\cpu.dec.do_flush_write ),
    .C(_04260_),
    .A(net721),
    .Y(_07335_));
 sg13g2_a21oi_1 _26412_ (.A1(_07334_),
    .A2(_07335_),
    .Y(_00945_),
    .B1(_06735_));
 sg13g2_nand2_1 _26413_ (.Y(_07336_),
    .A(\cpu.dec.io ),
    .B(_04260_));
 sg13g2_nand2_1 _26414_ (.Y(_07337_),
    .A(_02952_),
    .B(net1036));
 sg13g2_a21oi_1 _26415_ (.A1(_07336_),
    .A2(_07337_),
    .Y(_00948_),
    .B1(_06735_));
 sg13g2_nor2b_1 _26416_ (.A(_09257_),
    .B_N(_07318_),
    .Y(_07338_));
 sg13g2_nand2_1 _26417_ (.Y(_07339_),
    .A(_10526_),
    .B(net572));
 sg13g2_o21ai_1 _26418_ (.B1(_07339_),
    .Y(_07340_),
    .A1(_10180_),
    .A2(net572));
 sg13g2_nor2_1 _26419_ (.A(_07318_),
    .B(_07340_),
    .Y(_07341_));
 sg13g2_nor3_1 _26420_ (.A(_09954_),
    .B(_07338_),
    .C(_07341_),
    .Y(_00995_));
 sg13g2_inv_1 _26421_ (.Y(_07342_),
    .A(_11544_));
 sg13g2_a22oi_1 _26422_ (.Y(_07343_),
    .B1(_07342_),
    .B2(net1060),
    .A2(_04260_),
    .A1(_11521_));
 sg13g2_nor2_1 _26423_ (.A(_09297_),
    .B(_07343_),
    .Y(_00996_));
 sg13g2_and2_1 _26424_ (.A(_10749_),
    .B(_05832_),
    .X(_07344_));
 sg13g2_buf_1 _26425_ (.A(_07344_),
    .X(_07345_));
 sg13g2_mux2_1 _26426_ (.A0(_10444_),
    .A1(_09266_),
    .S(_07345_),
    .X(_07346_));
 sg13g2_nand2_1 _26427_ (.Y(_07347_),
    .A(_04257_),
    .B(_07346_));
 sg13g2_buf_1 _26428_ (.A(_06734_),
    .X(_07348_));
 sg13g2_a21oi_1 _26429_ (.A1(_11522_),
    .A2(_07347_),
    .Y(_01072_),
    .B1(net571));
 sg13g2_nor2_1 _26430_ (.A(_09449_),
    .B(_04257_),
    .Y(_07349_));
 sg13g2_nand2_1 _26431_ (.Y(_07350_),
    .A(net596),
    .B(_07345_));
 sg13g2_o21ai_1 _26432_ (.B1(_07350_),
    .Y(_07351_),
    .A1(_10637_),
    .A2(_07345_));
 sg13g2_nor2_1 _26433_ (.A(net294),
    .B(_07351_),
    .Y(_07352_));
 sg13g2_nor3_1 _26434_ (.A(_09954_),
    .B(_07349_),
    .C(_07352_),
    .Y(_01073_));
 sg13g2_mux2_1 _26435_ (.A0(\cpu.ex.mmu_read[1] ),
    .A1(_10107_),
    .S(_07345_),
    .X(_07353_));
 sg13g2_a21oi_1 _26436_ (.A1(_08537_),
    .A2(_07353_),
    .Y(_07354_),
    .B1(_10734_));
 sg13g2_nor2_1 _26437_ (.A(_09297_),
    .B(_07354_),
    .Y(_01074_));
 sg13g2_buf_1 _26438_ (.A(_09296_),
    .X(_07355_));
 sg13g2_nor2_1 _26439_ (.A(_10472_),
    .B(net1108),
    .Y(_07356_));
 sg13g2_and3_1 _26440_ (.X(_07357_),
    .A(net956),
    .B(net1081),
    .C(_05935_));
 sg13g2_buf_1 _26441_ (.A(_07357_),
    .X(_07358_));
 sg13g2_and2_1 _26442_ (.A(_07356_),
    .B(_07358_),
    .X(_07359_));
 sg13g2_buf_1 _26443_ (.A(_07359_),
    .X(_07360_));
 sg13g2_nor2b_1 _26444_ (.A(_00255_),
    .B_N(_05830_),
    .Y(_07361_));
 sg13g2_o21ai_1 _26445_ (.B1(_07361_),
    .Y(_07362_),
    .A1(_10749_),
    .A2(_00253_));
 sg13g2_a21o_1 _26446_ (.A2(_07362_),
    .A1(_05829_),
    .B1(_08615_),
    .X(_07363_));
 sg13g2_buf_1 _26447_ (.A(_07363_),
    .X(_07364_));
 sg13g2_buf_1 _26448_ (.A(_05829_),
    .X(_07365_));
 sg13g2_nand2b_1 _26449_ (.Y(_07366_),
    .B(net569),
    .A_N(_07364_));
 sg13g2_buf_1 _26450_ (.A(_07366_),
    .X(_07367_));
 sg13g2_a21oi_1 _26451_ (.A1(_03384_),
    .A2(_11008_),
    .Y(_07368_),
    .B1(_07365_));
 sg13g2_nor2_1 _26452_ (.A(_07364_),
    .B(_07368_),
    .Y(_07369_));
 sg13g2_buf_2 _26453_ (.A(_07369_),
    .X(_07370_));
 sg13g2_o21ai_1 _26454_ (.B1(_07370_),
    .Y(_07371_),
    .A1(_07360_),
    .A2(net177));
 sg13g2_nor2_1 _26455_ (.A(_10054_),
    .B(_07366_),
    .Y(_07372_));
 sg13g2_buf_2 _26456_ (.A(_07372_),
    .X(_07373_));
 sg13g2_buf_1 _26457_ (.A(_07373_),
    .X(_07374_));
 sg13g2_a22oi_1 _26458_ (.Y(_07375_),
    .B1(net120),
    .B2(_07360_),
    .A2(_07371_),
    .A1(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_nor2_1 _26459_ (.A(net570),
    .B(_07375_),
    .Y(_01075_));
 sg13g2_nor2_2 _26460_ (.A(net959),
    .B(_05894_),
    .Y(_07376_));
 sg13g2_nor2_1 _26461_ (.A(net864),
    .B(net1108),
    .Y(_07377_));
 sg13g2_a21oi_1 _26462_ (.A1(net1081),
    .A2(_05935_),
    .Y(_07378_),
    .B1(net956));
 sg13g2_a21o_1 _26463_ (.A2(_07358_),
    .A1(net952),
    .B1(_07378_),
    .X(_07379_));
 sg13g2_and2_1 _26464_ (.A(net864),
    .B(_07379_),
    .X(_07380_));
 sg13g2_a21oi_1 _26465_ (.A1(_07358_),
    .A2(_07377_),
    .Y(_07381_),
    .B1(_07380_));
 sg13g2_buf_2 _26466_ (.A(_07381_),
    .X(_07382_));
 sg13g2_nor2_1 _26467_ (.A(_07367_),
    .B(_07382_),
    .Y(_07383_));
 sg13g2_buf_1 _26468_ (.A(net177),
    .X(_07384_));
 sg13g2_buf_1 _26469_ (.A(_07370_),
    .X(_07385_));
 sg13g2_o21ai_1 _26470_ (.B1(net148),
    .Y(_07386_),
    .A1(_05896_),
    .A2(net149));
 sg13g2_a22oi_1 _26471_ (.Y(_07387_),
    .B1(_07386_),
    .B2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A2(_07383_),
    .A1(_07376_));
 sg13g2_nor2_1 _26472_ (.A(net570),
    .B(_07387_),
    .Y(_01076_));
 sg13g2_o21ai_1 _26473_ (.B1(_07385_),
    .Y(_07388_),
    .A1(_05906_),
    .A2(_07384_));
 sg13g2_a22oi_1 _26474_ (.Y(_07389_),
    .B1(_07388_),
    .B2(\cpu.genblk1.mmu.r_valid_d[11] ),
    .A2(_07373_),
    .A1(_05906_));
 sg13g2_nor2_1 _26475_ (.A(net570),
    .B(_07389_),
    .Y(_01077_));
 sg13g2_nor4_1 _26476_ (.A(net952),
    .B(net958),
    .C(_05854_),
    .D(net959),
    .Y(_07390_));
 sg13g2_buf_1 _26477_ (.A(_07390_),
    .X(_07391_));
 sg13g2_nor3_1 _26478_ (.A(net952),
    .B(net958),
    .C(_05854_),
    .Y(_07392_));
 sg13g2_o21ai_1 _26479_ (.B1(_05835_),
    .Y(_07393_),
    .A1(_05857_),
    .A2(_07392_));
 sg13g2_nor2_1 _26480_ (.A(_07382_),
    .B(_07393_),
    .Y(_07394_));
 sg13g2_o21ai_1 _26481_ (.B1(net148),
    .Y(_07395_),
    .A1(net149),
    .A2(_07394_));
 sg13g2_a22oi_1 _26482_ (.Y(_07396_),
    .B1(_07395_),
    .B2(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A2(_07391_),
    .A1(_07383_));
 sg13g2_nor2_1 _26483_ (.A(net570),
    .B(_07396_),
    .Y(_01078_));
 sg13g2_nand3_1 _26484_ (.B(_05843_),
    .C(net957),
    .A(net952),
    .Y(_07397_));
 sg13g2_buf_1 _26485_ (.A(_07397_),
    .X(_07398_));
 sg13g2_nor2_2 _26486_ (.A(_07382_),
    .B(_07398_),
    .Y(_07399_));
 sg13g2_o21ai_1 _26487_ (.B1(net148),
    .Y(_07400_),
    .A1(net149),
    .A2(_07399_));
 sg13g2_a22oi_1 _26488_ (.Y(_07401_),
    .B1(_07400_),
    .B2(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(_07399_),
    .A1(net120));
 sg13g2_nor2_1 _26489_ (.A(net570),
    .B(_07401_),
    .Y(_01079_));
 sg13g2_nor4_1 _26490_ (.A(net952),
    .B(_05843_),
    .C(_05854_),
    .D(net959),
    .Y(_07402_));
 sg13g2_buf_2 _26491_ (.A(_07402_),
    .X(_07403_));
 sg13g2_nand2_1 _26492_ (.Y(_07404_),
    .A(_05858_),
    .B(_05845_));
 sg13g2_nor2_1 _26493_ (.A(_07382_),
    .B(_07404_),
    .Y(_07405_));
 sg13g2_o21ai_1 _26494_ (.B1(net148),
    .Y(_07406_),
    .A1(net149),
    .A2(_07405_));
 sg13g2_a22oi_1 _26495_ (.Y(_07407_),
    .B1(_07406_),
    .B2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A2(_07403_),
    .A1(_07383_));
 sg13g2_nor2_1 _26496_ (.A(net570),
    .B(_07407_),
    .Y(_01080_));
 sg13g2_nor2_2 _26497_ (.A(_05869_),
    .B(_07382_),
    .Y(_07408_));
 sg13g2_o21ai_1 _26498_ (.B1(_07385_),
    .Y(_07409_),
    .A1(_07384_),
    .A2(_07408_));
 sg13g2_a22oi_1 _26499_ (.Y(_07410_),
    .B1(_07409_),
    .B2(\cpu.genblk1.mmu.r_valid_d[15] ),
    .A2(_07408_),
    .A1(net120));
 sg13g2_nor2_1 _26500_ (.A(net570),
    .B(_07410_),
    .Y(_01081_));
 sg13g2_a21oi_1 _26501_ (.A1(_03384_),
    .A2(_10500_),
    .Y(_07411_),
    .B1(_07365_));
 sg13g2_or2_1 _26502_ (.X(_07412_),
    .B(_07411_),
    .A(_07364_));
 sg13g2_buf_1 _26503_ (.A(_07412_),
    .X(_07413_));
 sg13g2_a21o_1 _26504_ (.A2(_07377_),
    .A1(_07358_),
    .B1(_07380_),
    .X(_07414_));
 sg13g2_buf_1 _26505_ (.A(_07414_),
    .X(_07415_));
 sg13g2_o21ai_1 _26506_ (.B1(_05869_),
    .Y(_07416_),
    .A1(_05882_),
    .A2(_05936_));
 sg13g2_and2_1 _26507_ (.A(net1081),
    .B(_07416_),
    .X(_07417_));
 sg13g2_buf_1 _26508_ (.A(_07417_),
    .X(_07418_));
 sg13g2_nor2_1 _26509_ (.A(_10520_),
    .B(_05827_),
    .Y(_07419_));
 sg13g2_nor2b_1 _26510_ (.A(_07419_),
    .B_N(_03384_),
    .Y(_07420_));
 sg13g2_buf_1 _26511_ (.A(_07420_),
    .X(_07421_));
 sg13g2_buf_1 _26512_ (.A(net568),
    .X(_07422_));
 sg13g2_a21oi_1 _26513_ (.A1(_07415_),
    .A2(_07418_),
    .Y(_07423_),
    .B1(net485));
 sg13g2_o21ai_1 _26514_ (.B1(\cpu.genblk1.mmu.r_valid_d[16] ),
    .Y(_07424_),
    .A1(net176),
    .A2(_07423_));
 sg13g2_nor2_1 _26515_ (.A(_07364_),
    .B(_07411_),
    .Y(_07425_));
 sg13g2_buf_1 _26516_ (.A(_07425_),
    .X(_07426_));
 sg13g2_a21oi_1 _26517_ (.A1(net1081),
    .A2(_05882_),
    .Y(_07427_),
    .B1(_05406_));
 sg13g2_and2_1 _26518_ (.A(_06115_),
    .B(_07427_),
    .X(_07428_));
 sg13g2_buf_1 _26519_ (.A(_07428_),
    .X(_07429_));
 sg13g2_nand4_1 _26520_ (.B(_07415_),
    .C(net175),
    .A(net569),
    .Y(_07430_),
    .D(_07429_));
 sg13g2_a21oi_1 _26521_ (.A1(_07424_),
    .A2(_07430_),
    .Y(_01082_),
    .B1(_07348_));
 sg13g2_nor2_1 _26522_ (.A(net954),
    .B(net1081),
    .Y(_07431_));
 sg13g2_a22oi_1 _26523_ (.Y(_07432_),
    .B1(_07356_),
    .B2(_07431_),
    .A2(_06192_),
    .A1(net1081));
 sg13g2_inv_1 _26524_ (.Y(_07433_),
    .A(_07432_));
 sg13g2_nand2b_1 _26525_ (.Y(_07434_),
    .B(net952),
    .A_N(net1081));
 sg13g2_a21oi_1 _26526_ (.A1(_05935_),
    .A2(_07434_),
    .Y(_07435_),
    .B1(net954));
 sg13g2_a22oi_1 _26527_ (.Y(_07436_),
    .B1(_07435_),
    .B2(net955),
    .A2(_07433_),
    .A1(_05935_));
 sg13g2_buf_2 _26528_ (.A(_07436_),
    .X(_07437_));
 sg13g2_nor3_1 _26529_ (.A(net957),
    .B(_05847_),
    .C(_07437_),
    .Y(_07438_));
 sg13g2_nand2_1 _26530_ (.Y(_07439_),
    .A(net120),
    .B(_07438_));
 sg13g2_nor2_1 _26531_ (.A(_07421_),
    .B(_07438_),
    .Y(_07440_));
 sg13g2_o21ai_1 _26532_ (.B1(\cpu.genblk1.mmu.r_valid_d[17] ),
    .Y(_07441_),
    .A1(net176),
    .A2(_07440_));
 sg13g2_a21oi_1 _26533_ (.A1(_07439_),
    .A2(_07441_),
    .Y(_01083_),
    .B1(net571));
 sg13g2_nor2_1 _26534_ (.A(_07367_),
    .B(_07437_),
    .Y(_07442_));
 sg13g2_o21ai_1 _26535_ (.B1(net175),
    .Y(_07443_),
    .A1(net485),
    .A2(_05945_));
 sg13g2_a22oi_1 _26536_ (.Y(_07444_),
    .B1(_07443_),
    .B2(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A2(_07442_),
    .A1(_07376_));
 sg13g2_nor2_1 _26537_ (.A(_07355_),
    .B(_07444_),
    .Y(_01084_));
 sg13g2_o21ai_1 _26538_ (.B1(net175),
    .Y(_07445_),
    .A1(net485),
    .A2(_05955_));
 sg13g2_a22oi_1 _26539_ (.Y(_07446_),
    .B1(_07445_),
    .B2(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(_07373_),
    .A1(_05955_));
 sg13g2_nor2_1 _26540_ (.A(_07355_),
    .B(_07446_),
    .Y(_01085_));
 sg13g2_a22oi_1 _26541_ (.Y(_07447_),
    .B1(_07377_),
    .B2(_07431_),
    .A2(_05911_),
    .A1(net1081));
 sg13g2_inv_1 _26542_ (.Y(_07448_),
    .A(_07447_));
 sg13g2_a22oi_1 _26543_ (.Y(_07449_),
    .B1(_07448_),
    .B2(_05935_),
    .A2(_07435_),
    .A1(net864));
 sg13g2_buf_1 _26544_ (.A(_07449_),
    .X(_07450_));
 sg13g2_nor3_2 _26545_ (.A(net957),
    .B(_05847_),
    .C(net426),
    .Y(_07451_));
 sg13g2_o21ai_1 _26546_ (.B1(net148),
    .Y(_07452_),
    .A1(net149),
    .A2(_07451_));
 sg13g2_a22oi_1 _26547_ (.Y(_07453_),
    .B1(_07452_),
    .B2(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(_07451_),
    .A1(net120));
 sg13g2_nor2_1 _26548_ (.A(net570),
    .B(_07453_),
    .Y(_01086_));
 sg13g2_nand2_1 _26549_ (.Y(_07454_),
    .A(_07391_),
    .B(_07442_));
 sg13g2_inv_1 _26550_ (.Y(_07455_),
    .A(_07393_));
 sg13g2_inv_1 _26551_ (.Y(_07456_),
    .A(_07437_));
 sg13g2_a21oi_1 _26552_ (.A1(_07455_),
    .A2(_07456_),
    .Y(_07457_),
    .B1(net568));
 sg13g2_o21ai_1 _26553_ (.B1(\cpu.genblk1.mmu.r_valid_d[20] ),
    .Y(_07458_),
    .A1(net176),
    .A2(_07457_));
 sg13g2_a21oi_1 _26554_ (.A1(_07454_),
    .A2(_07458_),
    .Y(_01087_),
    .B1(net571));
 sg13g2_buf_1 _26555_ (.A(_09296_),
    .X(_07459_));
 sg13g2_nor2_2 _26556_ (.A(_07398_),
    .B(_07437_),
    .Y(_07460_));
 sg13g2_o21ai_1 _26557_ (.B1(net175),
    .Y(_07461_),
    .A1(net485),
    .A2(_07460_));
 sg13g2_a22oi_1 _26558_ (.Y(_07462_),
    .B1(_07461_),
    .B2(\cpu.genblk1.mmu.r_valid_d[21] ),
    .A2(_07460_),
    .A1(net120));
 sg13g2_nor2_1 _26559_ (.A(_07459_),
    .B(_07462_),
    .Y(_01088_));
 sg13g2_nor2_1 _26560_ (.A(_07404_),
    .B(_07437_),
    .Y(_07463_));
 sg13g2_nor2_1 _26561_ (.A(net485),
    .B(_07463_),
    .Y(_07464_));
 sg13g2_o21ai_1 _26562_ (.B1(\cpu.genblk1.mmu.r_valid_d[22] ),
    .Y(_07465_),
    .A1(net176),
    .A2(_07464_));
 sg13g2_nand4_1 _26563_ (.B(_07403_),
    .C(net175),
    .A(net569),
    .Y(_07466_),
    .D(_07456_));
 sg13g2_a21oi_1 _26564_ (.A1(_07465_),
    .A2(_07466_),
    .Y(_01089_),
    .B1(net571));
 sg13g2_nor2_1 _26565_ (.A(_05953_),
    .B(_06039_),
    .Y(_07467_));
 sg13g2_nand2_1 _26566_ (.Y(_07468_),
    .A(net120),
    .B(_07467_));
 sg13g2_nor2_1 _26567_ (.A(net568),
    .B(_07467_),
    .Y(_07469_));
 sg13g2_o21ai_1 _26568_ (.B1(\cpu.genblk1.mmu.r_valid_d[23] ),
    .Y(_07470_),
    .A1(net176),
    .A2(_07469_));
 sg13g2_a21oi_1 _26569_ (.A1(_07468_),
    .A2(_07470_),
    .Y(_01090_),
    .B1(net571));
 sg13g2_nand2_1 _26570_ (.Y(_07471_),
    .A(_07429_),
    .B(_07442_));
 sg13g2_a21oi_1 _26571_ (.A1(_07418_),
    .A2(_07456_),
    .Y(_07472_),
    .B1(net568));
 sg13g2_o21ai_1 _26572_ (.B1(\cpu.genblk1.mmu.r_valid_d[24] ),
    .Y(_07473_),
    .A1(_07413_),
    .A2(_07472_));
 sg13g2_a21oi_1 _26573_ (.A1(_07471_),
    .A2(_07473_),
    .Y(_01091_),
    .B1(_07348_));
 sg13g2_a21o_1 _26574_ (.A2(_07379_),
    .A1(net955),
    .B1(_07360_),
    .X(_07474_));
 sg13g2_buf_1 _26575_ (.A(_07474_),
    .X(_07475_));
 sg13g2_inv_1 _26576_ (.Y(_07476_),
    .A(net337));
 sg13g2_nor3_2 _26577_ (.A(net957),
    .B(_05847_),
    .C(_07476_),
    .Y(_07477_));
 sg13g2_o21ai_1 _26578_ (.B1(_07426_),
    .Y(_07478_),
    .A1(net485),
    .A2(_07477_));
 sg13g2_a22oi_1 _26579_ (.Y(_07479_),
    .B1(_07478_),
    .B2(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(_07477_),
    .A1(_07374_));
 sg13g2_nor2_1 _26580_ (.A(net567),
    .B(_07479_),
    .Y(_01092_));
 sg13g2_nor2_1 _26581_ (.A(net485),
    .B(_07364_),
    .Y(_07480_));
 sg13g2_nand3_1 _26582_ (.B(_07376_),
    .C(net337),
    .A(_07480_),
    .Y(_07481_));
 sg13g2_nor2_1 _26583_ (.A(net568),
    .B(_05993_),
    .Y(_07482_));
 sg13g2_o21ai_1 _26584_ (.B1(\cpu.genblk1.mmu.r_valid_d[26] ),
    .Y(_07483_),
    .A1(net176),
    .A2(_07482_));
 sg13g2_a21oi_1 _26585_ (.A1(_07481_),
    .A2(_07483_),
    .Y(_01093_),
    .B1(net571));
 sg13g2_nand2_1 _26586_ (.Y(_07484_),
    .A(_05997_),
    .B(_07374_));
 sg13g2_nor2_1 _26587_ (.A(net568),
    .B(_05997_),
    .Y(_07485_));
 sg13g2_o21ai_1 _26588_ (.B1(\cpu.genblk1.mmu.r_valid_d[27] ),
    .Y(_07486_),
    .A1(net176),
    .A2(_07485_));
 sg13g2_a21oi_1 _26589_ (.A1(_07484_),
    .A2(_07486_),
    .Y(_01094_),
    .B1(net571));
 sg13g2_nand3_1 _26590_ (.B(_07391_),
    .C(net337),
    .A(_07480_),
    .Y(_07487_));
 sg13g2_a21oi_1 _26591_ (.A1(_07455_),
    .A2(net337),
    .Y(_07488_),
    .B1(net568));
 sg13g2_o21ai_1 _26592_ (.B1(\cpu.genblk1.mmu.r_valid_d[28] ),
    .Y(_07489_),
    .A1(_07413_),
    .A2(_07488_));
 sg13g2_a21oi_1 _26593_ (.A1(_07487_),
    .A2(_07489_),
    .Y(_01095_),
    .B1(net571));
 sg13g2_nor2_2 _26594_ (.A(_07398_),
    .B(_07476_),
    .Y(_07490_));
 sg13g2_o21ai_1 _26595_ (.B1(net175),
    .Y(_07491_),
    .A1(_07422_),
    .A2(_07490_));
 sg13g2_a22oi_1 _26596_ (.Y(_07492_),
    .B1(_07491_),
    .B2(\cpu.genblk1.mmu.r_valid_d[29] ),
    .A2(_07490_),
    .A1(net120));
 sg13g2_nor2_1 _26597_ (.A(net567),
    .B(_07492_),
    .Y(_01096_));
 sg13g2_nor2_1 _26598_ (.A(_05894_),
    .B(net426),
    .Y(_07493_));
 sg13g2_o21ai_1 _26599_ (.B1(_07370_),
    .Y(_07494_),
    .A1(net177),
    .A2(_07493_));
 sg13g2_nor3_1 _26600_ (.A(_05406_),
    .B(_05894_),
    .C(net426),
    .Y(_07495_));
 sg13g2_a22oi_1 _26601_ (.Y(_07496_),
    .B1(_07495_),
    .B2(_07480_),
    .A2(_07494_),
    .A1(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_nor2_1 _26602_ (.A(net567),
    .B(_07496_),
    .Y(_01097_));
 sg13g2_inv_1 _26603_ (.Y(_07497_),
    .A(_07404_));
 sg13g2_a21oi_1 _26604_ (.A1(_07497_),
    .A2(net337),
    .Y(_07498_),
    .B1(net485));
 sg13g2_o21ai_1 _26605_ (.B1(\cpu.genblk1.mmu.r_valid_d[30] ),
    .Y(_07499_),
    .A1(net176),
    .A2(_07498_));
 sg13g2_nand4_1 _26606_ (.B(_07403_),
    .C(net175),
    .A(net569),
    .Y(_07500_),
    .D(_07475_));
 sg13g2_buf_1 _26607_ (.A(_06734_),
    .X(_07501_));
 sg13g2_a21oi_1 _26608_ (.A1(_07499_),
    .A2(_07500_),
    .Y(_01098_),
    .B1(net566));
 sg13g2_nor2_2 _26609_ (.A(_05869_),
    .B(_07476_),
    .Y(_07502_));
 sg13g2_o21ai_1 _26610_ (.B1(net175),
    .Y(_07503_),
    .A1(_07422_),
    .A2(_07502_));
 sg13g2_a22oi_1 _26611_ (.Y(_07504_),
    .B1(_07503_),
    .B2(\cpu.genblk1.mmu.r_valid_d[31] ),
    .A2(_07502_),
    .A1(_07373_));
 sg13g2_nor2_1 _26612_ (.A(_07459_),
    .B(_07504_),
    .Y(_01099_));
 sg13g2_nor2b_2 _26613_ (.A(net426),
    .B_N(_05857_),
    .Y(_07505_));
 sg13g2_o21ai_1 _26614_ (.B1(net148),
    .Y(_07506_),
    .A1(net177),
    .A2(_07505_));
 sg13g2_a22oi_1 _26615_ (.Y(_07507_),
    .B1(_07506_),
    .B2(\cpu.genblk1.mmu.r_valid_d[3] ),
    .A2(_07505_),
    .A1(_07373_));
 sg13g2_nor2_1 _26616_ (.A(net567),
    .B(_07507_),
    .Y(_01100_));
 sg13g2_nor2_1 _26617_ (.A(net177),
    .B(net426),
    .Y(_07508_));
 sg13g2_nor2_1 _26618_ (.A(_07393_),
    .B(net426),
    .Y(_07509_));
 sg13g2_o21ai_1 _26619_ (.B1(net148),
    .Y(_07510_),
    .A1(net177),
    .A2(_07509_));
 sg13g2_a22oi_1 _26620_ (.Y(_07511_),
    .B1(_07510_),
    .B2(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A2(_07508_),
    .A1(_07391_));
 sg13g2_nor2_1 _26621_ (.A(net567),
    .B(_07511_),
    .Y(_01101_));
 sg13g2_o21ai_1 _26622_ (.B1(net148),
    .Y(_07512_),
    .A1(_06034_),
    .A2(net149));
 sg13g2_a22oi_1 _26623_ (.Y(_07513_),
    .B1(_07512_),
    .B2(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(_07373_),
    .A1(_06034_));
 sg13g2_nor2_1 _26624_ (.A(net567),
    .B(_07513_),
    .Y(_01102_));
 sg13g2_o21ai_1 _26625_ (.B1(_07370_),
    .Y(_07514_),
    .A1(_06040_),
    .A2(net149));
 sg13g2_a22oi_1 _26626_ (.Y(_07515_),
    .B1(_07514_),
    .B2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A2(_07508_),
    .A1(_07403_));
 sg13g2_nor2_1 _26627_ (.A(net567),
    .B(_07515_),
    .Y(_01103_));
 sg13g2_o21ai_1 _26628_ (.B1(_07370_),
    .Y(_07516_),
    .A1(_06045_),
    .A2(net149));
 sg13g2_a22oi_1 _26629_ (.Y(_07517_),
    .B1(_07516_),
    .B2(\cpu.genblk1.mmu.r_valid_d[7] ),
    .A2(_07373_),
    .A1(_06045_));
 sg13g2_nor2_1 _26630_ (.A(net567),
    .B(_07517_),
    .Y(_01104_));
 sg13g2_buf_1 _26631_ (.A(_09296_),
    .X(_07518_));
 sg13g2_nor2b_1 _26632_ (.A(_07450_),
    .B_N(_07418_),
    .Y(_07519_));
 sg13g2_o21ai_1 _26633_ (.B1(_07370_),
    .Y(_07520_),
    .A1(net177),
    .A2(_07519_));
 sg13g2_a22oi_1 _26634_ (.Y(_07521_),
    .B1(_07520_),
    .B2(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A2(_07508_),
    .A1(_07429_));
 sg13g2_nor2_1 _26635_ (.A(net565),
    .B(_07521_),
    .Y(_01105_));
 sg13g2_nor3_2 _26636_ (.A(net957),
    .B(_05847_),
    .C(_07382_),
    .Y(_07522_));
 sg13g2_o21ai_1 _26637_ (.B1(_07370_),
    .Y(_07523_),
    .A1(net177),
    .A2(_07522_));
 sg13g2_a22oi_1 _26638_ (.Y(_07524_),
    .B1(_07523_),
    .B2(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(_07522_),
    .A1(_07373_));
 sg13g2_nor2_1 _26639_ (.A(_07518_),
    .B(_07524_),
    .Y(_01106_));
 sg13g2_nand2_1 _26640_ (.Y(_07525_),
    .A(_08582_),
    .B(_00253_));
 sg13g2_a21oi_1 _26641_ (.A1(_07361_),
    .A2(_07525_),
    .Y(_07526_),
    .B1(_07421_));
 sg13g2_nand2b_1 _26642_ (.Y(_07527_),
    .B(net330),
    .A_N(_07526_));
 sg13g2_buf_1 _26643_ (.A(_07527_),
    .X(_07528_));
 sg13g2_nand2b_1 _26644_ (.Y(_07529_),
    .B(net569),
    .A_N(_07528_));
 sg13g2_buf_2 _26645_ (.A(_07529_),
    .X(_07530_));
 sg13g2_nor2b_1 _26646_ (.A(_10520_),
    .B_N(_03384_),
    .Y(_07531_));
 sg13g2_a21oi_1 _26647_ (.A1(_05827_),
    .A2(_07531_),
    .Y(_07532_),
    .B1(_07528_));
 sg13g2_buf_2 _26648_ (.A(_07532_),
    .X(_07533_));
 sg13g2_o21ai_1 _26649_ (.B1(_07533_),
    .Y(_07534_),
    .A1(_07360_),
    .A2(_07530_));
 sg13g2_nor2_1 _26650_ (.A(_10054_),
    .B(_07530_),
    .Y(_07535_));
 sg13g2_buf_2 _26651_ (.A(_07535_),
    .X(_07536_));
 sg13g2_buf_1 _26652_ (.A(_07536_),
    .X(_07537_));
 sg13g2_a22oi_1 _26653_ (.Y(_07538_),
    .B1(net112),
    .B2(_07360_),
    .A2(_07534_),
    .A1(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_nor2_1 _26654_ (.A(net565),
    .B(_07538_),
    .Y(_01107_));
 sg13g2_nor2_1 _26655_ (.A(net568),
    .B(_07528_),
    .Y(_07539_));
 sg13g2_and2_1 _26656_ (.A(_07376_),
    .B(_07539_),
    .X(_07540_));
 sg13g2_buf_1 _26657_ (.A(_07540_),
    .X(_07541_));
 sg13g2_buf_1 _26658_ (.A(_07530_),
    .X(_07542_));
 sg13g2_buf_1 _26659_ (.A(_07533_),
    .X(_07543_));
 sg13g2_o21ai_1 _26660_ (.B1(net146),
    .Y(_07544_),
    .A1(_05896_),
    .A2(net147));
 sg13g2_a22oi_1 _26661_ (.Y(_07545_),
    .B1(_07544_),
    .B2(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A2(_07541_),
    .A1(_07415_));
 sg13g2_nor2_1 _26662_ (.A(net565),
    .B(_07545_),
    .Y(_01108_));
 sg13g2_o21ai_1 _26663_ (.B1(net146),
    .Y(_07546_),
    .A1(_05906_),
    .A2(net147));
 sg13g2_a22oi_1 _26664_ (.Y(_07547_),
    .B1(_07546_),
    .B2(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A2(net112),
    .A1(_05906_));
 sg13g2_nor2_1 _26665_ (.A(net565),
    .B(_07547_),
    .Y(_01109_));
 sg13g2_and2_1 _26666_ (.A(_07391_),
    .B(_07539_),
    .X(_07548_));
 sg13g2_buf_1 _26667_ (.A(_07548_),
    .X(_07549_));
 sg13g2_o21ai_1 _26668_ (.B1(_07543_),
    .Y(_07550_),
    .A1(_07394_),
    .A2(net147));
 sg13g2_a22oi_1 _26669_ (.Y(_07551_),
    .B1(_07550_),
    .B2(\cpu.genblk1.mmu.r_valid_i[12] ),
    .A2(_07549_),
    .A1(_07415_));
 sg13g2_nor2_1 _26670_ (.A(net565),
    .B(_07551_),
    .Y(_01110_));
 sg13g2_o21ai_1 _26671_ (.B1(net146),
    .Y(_07552_),
    .A1(_07399_),
    .A2(net147));
 sg13g2_a22oi_1 _26672_ (.Y(_07553_),
    .B1(_07552_),
    .B2(\cpu.genblk1.mmu.r_valid_i[13] ),
    .A2(net112),
    .A1(_07399_));
 sg13g2_nor2_1 _26673_ (.A(net565),
    .B(_07553_),
    .Y(_01111_));
 sg13g2_o21ai_1 _26674_ (.B1(_07533_),
    .Y(_07554_),
    .A1(_07405_),
    .A2(_07530_));
 sg13g2_nand2_1 _26675_ (.Y(_07555_),
    .A(\cpu.genblk1.mmu.r_valid_i[14] ),
    .B(_07554_));
 sg13g2_nand3_1 _26676_ (.B(_07403_),
    .C(_07539_),
    .A(_07415_),
    .Y(_07556_));
 sg13g2_a21oi_1 _26677_ (.A1(_07555_),
    .A2(_07556_),
    .Y(_01112_),
    .B1(net566));
 sg13g2_o21ai_1 _26678_ (.B1(net146),
    .Y(_07557_),
    .A1(_07408_),
    .A2(net147));
 sg13g2_a22oi_1 _26679_ (.Y(_07558_),
    .B1(_07557_),
    .B2(\cpu.genblk1.mmu.r_valid_i[15] ),
    .A2(net112),
    .A1(_07408_));
 sg13g2_nor2_1 _26680_ (.A(net565),
    .B(_07558_),
    .Y(_01113_));
 sg13g2_a21oi_1 _26681_ (.A1(_03384_),
    .A2(_10465_),
    .Y(_07559_),
    .B1(net569));
 sg13g2_or2_1 _26682_ (.X(_07560_),
    .B(_07559_),
    .A(_07528_));
 sg13g2_buf_1 _26683_ (.A(_07560_),
    .X(_07561_));
 sg13g2_o21ai_1 _26684_ (.B1(\cpu.genblk1.mmu.r_valid_i[16] ),
    .Y(_07562_),
    .A1(_07423_),
    .A2(net174));
 sg13g2_nor2_1 _26685_ (.A(_07528_),
    .B(_07559_),
    .Y(_07563_));
 sg13g2_buf_1 _26686_ (.A(_07563_),
    .X(_07564_));
 sg13g2_nand4_1 _26687_ (.B(_07415_),
    .C(_07429_),
    .A(net569),
    .Y(_07565_),
    .D(net173));
 sg13g2_a21oi_1 _26688_ (.A1(_07562_),
    .A2(_07565_),
    .Y(_01114_),
    .B1(net566));
 sg13g2_nand2_1 _26689_ (.Y(_07566_),
    .A(_07438_),
    .B(net112));
 sg13g2_o21ai_1 _26690_ (.B1(\cpu.genblk1.mmu.r_valid_i[17] ),
    .Y(_07567_),
    .A1(_07440_),
    .A2(net174));
 sg13g2_a21oi_1 _26691_ (.A1(_07566_),
    .A2(_07567_),
    .Y(_01115_),
    .B1(net566));
 sg13g2_o21ai_1 _26692_ (.B1(net173),
    .Y(_07568_),
    .A1(_05945_),
    .A2(net147));
 sg13g2_a22oi_1 _26693_ (.Y(_07569_),
    .B1(_07568_),
    .B2(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A2(_07541_),
    .A1(_07456_));
 sg13g2_nor2_1 _26694_ (.A(_07518_),
    .B(_07569_),
    .Y(_01116_));
 sg13g2_o21ai_1 _26695_ (.B1(net173),
    .Y(_07570_),
    .A1(_05955_),
    .A2(_07542_));
 sg13g2_a22oi_1 _26696_ (.Y(_07571_),
    .B1(_07570_),
    .B2(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A2(_07537_),
    .A1(_05955_));
 sg13g2_nor2_1 _26697_ (.A(net565),
    .B(_07571_),
    .Y(_01117_));
 sg13g2_buf_1 _26698_ (.A(_09296_),
    .X(_07572_));
 sg13g2_o21ai_1 _26699_ (.B1(net146),
    .Y(_07573_),
    .A1(_07451_),
    .A2(net147));
 sg13g2_a22oi_1 _26700_ (.Y(_07574_),
    .B1(_07573_),
    .B2(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A2(net112),
    .A1(_07451_));
 sg13g2_nor2_1 _26701_ (.A(net564),
    .B(_07574_),
    .Y(_01118_));
 sg13g2_nor2_1 _26702_ (.A(_07437_),
    .B(_07530_),
    .Y(_07575_));
 sg13g2_nand2_1 _26703_ (.Y(_07576_),
    .A(_07391_),
    .B(_07575_));
 sg13g2_o21ai_1 _26704_ (.B1(\cpu.genblk1.mmu.r_valid_i[20] ),
    .Y(_07577_),
    .A1(_07457_),
    .A2(net174));
 sg13g2_a21oi_1 _26705_ (.A1(_07576_),
    .A2(_07577_),
    .Y(_01119_),
    .B1(net566));
 sg13g2_o21ai_1 _26706_ (.B1(net173),
    .Y(_07578_),
    .A1(_07460_),
    .A2(net147));
 sg13g2_a22oi_1 _26707_ (.Y(_07579_),
    .B1(_07578_),
    .B2(\cpu.genblk1.mmu.r_valid_i[21] ),
    .A2(net112),
    .A1(_07460_));
 sg13g2_nor2_1 _26708_ (.A(_07572_),
    .B(_07579_),
    .Y(_01120_));
 sg13g2_o21ai_1 _26709_ (.B1(_07564_),
    .Y(_07580_),
    .A1(_07463_),
    .A2(_07542_));
 sg13g2_a22oi_1 _26710_ (.Y(_07581_),
    .B1(_07580_),
    .B2(\cpu.genblk1.mmu.r_valid_i[22] ),
    .A2(_07575_),
    .A1(_07403_));
 sg13g2_nor2_1 _26711_ (.A(_07572_),
    .B(_07581_),
    .Y(_01121_));
 sg13g2_nand2_1 _26712_ (.Y(_07582_),
    .A(_07467_),
    .B(_07537_));
 sg13g2_o21ai_1 _26713_ (.B1(\cpu.genblk1.mmu.r_valid_i[23] ),
    .Y(_07583_),
    .A1(_07469_),
    .A2(net174));
 sg13g2_a21oi_1 _26714_ (.A1(_07582_),
    .A2(_07583_),
    .Y(_01122_),
    .B1(net566));
 sg13g2_nand2_1 _26715_ (.Y(_07584_),
    .A(_07429_),
    .B(_07575_));
 sg13g2_o21ai_1 _26716_ (.B1(\cpu.genblk1.mmu.r_valid_i[24] ),
    .Y(_07585_),
    .A1(_07472_),
    .A2(net174));
 sg13g2_a21oi_1 _26717_ (.A1(_07584_),
    .A2(_07585_),
    .Y(_01123_),
    .B1(_07501_));
 sg13g2_buf_1 _26718_ (.A(_07530_),
    .X(_07586_));
 sg13g2_o21ai_1 _26719_ (.B1(net173),
    .Y(_07587_),
    .A1(_07477_),
    .A2(_07586_));
 sg13g2_a22oi_1 _26720_ (.Y(_07588_),
    .B1(_07587_),
    .B2(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A2(_07536_),
    .A1(_07477_));
 sg13g2_nor2_1 _26721_ (.A(net564),
    .B(_07588_),
    .Y(_01124_));
 sg13g2_nand2_1 _26722_ (.Y(_07589_),
    .A(net337),
    .B(_07541_));
 sg13g2_o21ai_1 _26723_ (.B1(\cpu.genblk1.mmu.r_valid_i[26] ),
    .Y(_07590_),
    .A1(_07482_),
    .A2(net174));
 sg13g2_a21oi_1 _26724_ (.A1(_07589_),
    .A2(_07590_),
    .Y(_01125_),
    .B1(net566));
 sg13g2_nand2_1 _26725_ (.Y(_07591_),
    .A(_05997_),
    .B(net112));
 sg13g2_o21ai_1 _26726_ (.B1(\cpu.genblk1.mmu.r_valid_i[27] ),
    .Y(_07592_),
    .A1(_07485_),
    .A2(net174));
 sg13g2_a21oi_1 _26727_ (.A1(_07591_),
    .A2(_07592_),
    .Y(_01126_),
    .B1(net566));
 sg13g2_nand2_1 _26728_ (.Y(_07593_),
    .A(net337),
    .B(_07549_));
 sg13g2_o21ai_1 _26729_ (.B1(\cpu.genblk1.mmu.r_valid_i[28] ),
    .Y(_07594_),
    .A1(_07488_),
    .A2(net174));
 sg13g2_a21oi_1 _26730_ (.A1(_07593_),
    .A2(_07594_),
    .Y(_01127_),
    .B1(_07501_));
 sg13g2_o21ai_1 _26731_ (.B1(net173),
    .Y(_07595_),
    .A1(_07490_),
    .A2(_07586_));
 sg13g2_a22oi_1 _26732_ (.Y(_07596_),
    .B1(_07595_),
    .B2(\cpu.genblk1.mmu.r_valid_i[29] ),
    .A2(_07536_),
    .A1(_07490_));
 sg13g2_nor2_1 _26733_ (.A(net564),
    .B(_07596_),
    .Y(_01128_));
 sg13g2_o21ai_1 _26734_ (.B1(_07543_),
    .Y(_07597_),
    .A1(_07493_),
    .A2(net145));
 sg13g2_a22oi_1 _26735_ (.Y(_07598_),
    .B1(_07597_),
    .B2(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(_07539_),
    .A1(_07495_));
 sg13g2_nor2_1 _26736_ (.A(net564),
    .B(_07598_),
    .Y(_01129_));
 sg13g2_o21ai_1 _26737_ (.B1(\cpu.genblk1.mmu.r_valid_i[30] ),
    .Y(_07599_),
    .A1(_07498_),
    .A2(_07561_));
 sg13g2_nand4_1 _26738_ (.B(_07403_),
    .C(net337),
    .A(net569),
    .Y(_07600_),
    .D(net173));
 sg13g2_buf_2 _26739_ (.A(_06734_),
    .X(_07601_));
 sg13g2_a21oi_1 _26740_ (.A1(_07599_),
    .A2(_07600_),
    .Y(_01130_),
    .B1(_07601_));
 sg13g2_o21ai_1 _26741_ (.B1(net173),
    .Y(_07602_),
    .A1(_07502_),
    .A2(net145));
 sg13g2_a22oi_1 _26742_ (.Y(_07603_),
    .B1(_07602_),
    .B2(\cpu.genblk1.mmu.r_valid_i[31] ),
    .A2(_07536_),
    .A1(_07502_));
 sg13g2_nor2_1 _26743_ (.A(net564),
    .B(_07603_),
    .Y(_01131_));
 sg13g2_o21ai_1 _26744_ (.B1(net146),
    .Y(_07604_),
    .A1(_07505_),
    .A2(net145));
 sg13g2_a22oi_1 _26745_ (.Y(_07605_),
    .B1(_07604_),
    .B2(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(_07536_),
    .A1(_07505_));
 sg13g2_nor2_1 _26746_ (.A(net564),
    .B(_07605_),
    .Y(_01132_));
 sg13g2_inv_1 _26747_ (.Y(_07606_),
    .A(net426));
 sg13g2_o21ai_1 _26748_ (.B1(net146),
    .Y(_07607_),
    .A1(_07509_),
    .A2(net145));
 sg13g2_a22oi_1 _26749_ (.Y(_07608_),
    .B1(_07607_),
    .B2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A2(_07549_),
    .A1(_07606_));
 sg13g2_nor2_1 _26750_ (.A(net564),
    .B(_07608_),
    .Y(_01133_));
 sg13g2_o21ai_1 _26751_ (.B1(net146),
    .Y(_07609_),
    .A1(_06034_),
    .A2(net145));
 sg13g2_a22oi_1 _26752_ (.Y(_07610_),
    .B1(_07609_),
    .B2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A2(_07536_),
    .A1(_06034_));
 sg13g2_nor2_1 _26753_ (.A(net564),
    .B(_07610_),
    .Y(_01134_));
 sg13g2_buf_1 _26754_ (.A(_09296_),
    .X(_07611_));
 sg13g2_o21ai_1 _26755_ (.B1(_07533_),
    .Y(_07612_),
    .A1(_06040_),
    .A2(_07530_));
 sg13g2_nor2_1 _26756_ (.A(net426),
    .B(_07530_),
    .Y(_07613_));
 sg13g2_a22oi_1 _26757_ (.Y(_07614_),
    .B1(_07613_),
    .B2(_07403_),
    .A2(_07612_),
    .A1(\cpu.genblk1.mmu.r_valid_i[6] ));
 sg13g2_nor2_1 _26758_ (.A(net562),
    .B(_07614_),
    .Y(_01135_));
 sg13g2_o21ai_1 _26759_ (.B1(_07533_),
    .Y(_07615_),
    .A1(_06045_),
    .A2(net145));
 sg13g2_a22oi_1 _26760_ (.Y(_07616_),
    .B1(_07615_),
    .B2(\cpu.genblk1.mmu.r_valid_i[7] ),
    .A2(_07536_),
    .A1(_06045_));
 sg13g2_nor2_1 _26761_ (.A(net562),
    .B(_07616_),
    .Y(_01136_));
 sg13g2_o21ai_1 _26762_ (.B1(_07533_),
    .Y(_07617_),
    .A1(_07519_),
    .A2(net145));
 sg13g2_a22oi_1 _26763_ (.Y(_07618_),
    .B1(_07617_),
    .B2(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A2(_07613_),
    .A1(_07429_));
 sg13g2_nor2_1 _26764_ (.A(_07611_),
    .B(_07618_),
    .Y(_01137_));
 sg13g2_o21ai_1 _26765_ (.B1(_07533_),
    .Y(_07619_),
    .A1(_07522_),
    .A2(net145));
 sg13g2_a22oi_1 _26766_ (.Y(_07620_),
    .B1(_07619_),
    .B2(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A2(_07536_),
    .A1(_07522_));
 sg13g2_nor2_1 _26767_ (.A(_07611_),
    .B(_07620_),
    .Y(_01138_));
 sg13g2_and2_1 _26768_ (.A(net362),
    .B(_06323_),
    .X(_07621_));
 sg13g2_buf_2 _26769_ (.A(_07621_),
    .X(_07622_));
 sg13g2_nand2_1 _26770_ (.Y(_07623_),
    .A(net799),
    .B(_07622_));
 sg13g2_nand2_1 _26771_ (.Y(_07624_),
    .A(net362),
    .B(_06323_));
 sg13g2_buf_2 _26772_ (.A(_07624_),
    .X(_07625_));
 sg13g2_nand2_1 _26773_ (.Y(_07626_),
    .A(_09219_),
    .B(_07625_));
 sg13g2_a21oi_1 _26774_ (.A1(_07623_),
    .A2(_07626_),
    .Y(_01939_),
    .B1(net563));
 sg13g2_nand2_1 _26775_ (.Y(_07627_),
    .A(net939),
    .B(_07622_));
 sg13g2_nand2_1 _26776_ (.Y(_07628_),
    .A(_09225_),
    .B(_07625_));
 sg13g2_a21oi_1 _26777_ (.A1(_07627_),
    .A2(_07628_),
    .Y(_01940_),
    .B1(net563));
 sg13g2_nand2_1 _26778_ (.Y(_07629_),
    .A(net849),
    .B(_07622_));
 sg13g2_nand2_1 _26779_ (.Y(_07630_),
    .A(\cpu.gpio.r_enable_in[2] ),
    .B(_07625_));
 sg13g2_a21oi_1 _26780_ (.A1(_07629_),
    .A2(_07630_),
    .Y(_01941_),
    .B1(net563));
 sg13g2_nand2_1 _26781_ (.Y(_07631_),
    .A(_10080_),
    .B(_07622_));
 sg13g2_nand2_1 _26782_ (.Y(_07632_),
    .A(_09229_),
    .B(_07625_));
 sg13g2_a21oi_1 _26783_ (.A1(_07631_),
    .A2(_07632_),
    .Y(_01942_),
    .B1(_07601_));
 sg13g2_nand2_1 _26784_ (.Y(_07633_),
    .A(net1024),
    .B(_07622_));
 sg13g2_nand2_1 _26785_ (.Y(_07634_),
    .A(_09233_),
    .B(_07625_));
 sg13g2_a21oi_1 _26786_ (.A1(_07633_),
    .A2(_07634_),
    .Y(_01943_),
    .B1(net563));
 sg13g2_nand2_1 _26787_ (.Y(_07635_),
    .A(net1023),
    .B(_07622_));
 sg13g2_nand2_1 _26788_ (.Y(_07636_),
    .A(_09235_),
    .B(_07625_));
 sg13g2_a21oi_1 _26789_ (.A1(_07635_),
    .A2(_07636_),
    .Y(_01944_),
    .B1(net563));
 sg13g2_nand2_1 _26790_ (.Y(_07637_),
    .A(net1022),
    .B(_07622_));
 sg13g2_nand2_1 _26791_ (.Y(_07638_),
    .A(_09221_),
    .B(_07625_));
 sg13g2_a21oi_1 _26792_ (.A1(_07637_),
    .A2(_07638_),
    .Y(_01945_),
    .B1(net563));
 sg13g2_nand2_1 _26793_ (.Y(_07639_),
    .A(net1021),
    .B(_07622_));
 sg13g2_nand2_1 _26794_ (.Y(_07640_),
    .A(\cpu.gpio.r_enable_in[7] ),
    .B(_07625_));
 sg13g2_a21oi_1 _26795_ (.A1(_07639_),
    .A2(_07640_),
    .Y(_01946_),
    .B1(net563));
 sg13g2_buf_1 _26796_ (.A(_06323_),
    .X(_07641_));
 sg13g2_nand3_1 _26797_ (.B(net392),
    .C(net111),
    .A(_10086_),
    .Y(_07642_));
 sg13g2_nand2_1 _26798_ (.Y(_07643_),
    .A(net392),
    .B(net111));
 sg13g2_nand2_1 _26799_ (.Y(_07644_),
    .A(_09238_),
    .B(_07643_));
 sg13g2_a21oi_1 _26800_ (.A1(_07642_),
    .A2(_07644_),
    .Y(_01947_),
    .B1(net563));
 sg13g2_nand3_1 _26801_ (.B(net392),
    .C(net111),
    .A(net1023),
    .Y(_07645_));
 sg13g2_nand2_1 _26802_ (.Y(_07646_),
    .A(_09240_),
    .B(_07643_));
 sg13g2_buf_1 _26803_ (.A(_06734_),
    .X(_07647_));
 sg13g2_a21oi_1 _26804_ (.A1(_07645_),
    .A2(_07646_),
    .Y(_01948_),
    .B1(net561));
 sg13g2_nand3_1 _26805_ (.B(_05336_),
    .C(_07641_),
    .A(net1022),
    .Y(_07648_));
 sg13g2_nand2_1 _26806_ (.Y(_07649_),
    .A(\cpu.gpio.r_enable_io[6] ),
    .B(_07643_));
 sg13g2_a21oi_1 _26807_ (.A1(_07648_),
    .A2(_07649_),
    .Y(_01949_),
    .B1(net561));
 sg13g2_nand3_1 _26808_ (.B(_05336_),
    .C(_07641_),
    .A(net1021),
    .Y(_07650_));
 sg13g2_nand2_1 _26809_ (.Y(_07651_),
    .A(\cpu.gpio.r_enable_io[7] ),
    .B(_07643_));
 sg13g2_a21oi_1 _26810_ (.A1(_07650_),
    .A2(_07651_),
    .Y(_01950_),
    .B1(net561));
 sg13g2_nand3_1 _26811_ (.B(net499),
    .C(_06323_),
    .A(net960),
    .Y(_07652_));
 sg13g2_buf_1 _26812_ (.A(_07652_),
    .X(_07653_));
 sg13g2_mux2_1 _26813_ (.A0(net1024),
    .A1(net7),
    .S(_07653_),
    .X(_07654_));
 sg13g2_and2_1 _26814_ (.A(net645),
    .B(_07654_),
    .X(_01951_));
 sg13g2_mux2_1 _26815_ (.A0(net1023),
    .A1(net8),
    .S(_07653_),
    .X(_07655_));
 sg13g2_and2_1 _26816_ (.A(net645),
    .B(_07655_),
    .X(_01952_));
 sg13g2_buf_1 _26817_ (.A(net764),
    .X(_07656_));
 sg13g2_mux2_1 _26818_ (.A0(net1022),
    .A1(net9),
    .S(_07653_),
    .X(_07657_));
 sg13g2_and2_1 _26819_ (.A(net644),
    .B(_07657_),
    .X(_01953_));
 sg13g2_mux2_1 _26820_ (.A0(_10103_),
    .A1(net10),
    .S(_07653_),
    .X(_07658_));
 sg13g2_and2_1 _26821_ (.A(net644),
    .B(_07658_),
    .X(_01954_));
 sg13g2_nand2_1 _26822_ (.Y(_07659_),
    .A(_04934_),
    .B(_06323_));
 sg13g2_buf_1 _26823_ (.A(_07659_),
    .X(_07660_));
 sg13g2_nor2_1 _26824_ (.A(net799),
    .B(_07660_),
    .Y(_07661_));
 sg13g2_a21oi_1 _26825_ (.A1(_04934_),
    .A2(net111),
    .Y(_07662_),
    .B1(_04933_));
 sg13g2_o21ai_1 _26826_ (.B1(net675),
    .Y(_02000_),
    .A1(_07661_),
    .A2(_07662_));
 sg13g2_buf_1 _26827_ (.A(\cpu.gpio.r_src_o[6][1] ),
    .X(_07663_));
 sg13g2_nand2_1 _26828_ (.Y(_07664_),
    .A(_07663_),
    .B(_07660_));
 sg13g2_o21ai_1 _26829_ (.B1(_07664_),
    .Y(_07665_),
    .A1(net887),
    .A2(_07660_));
 sg13g2_and2_1 _26830_ (.A(net644),
    .B(_07665_),
    .X(_02001_));
 sg13g2_mux2_1 _26831_ (.A0(_10075_),
    .A1(\cpu.gpio.r_src_o[6][2] ),
    .S(_07660_),
    .X(_07666_));
 sg13g2_and2_1 _26832_ (.A(net644),
    .B(_07666_),
    .X(_02002_));
 sg13g2_mux2_1 _26833_ (.A0(net1025),
    .A1(\cpu.gpio.r_src_o[6][3] ),
    .S(_07660_),
    .X(_07667_));
 sg13g2_and2_1 _26834_ (.A(net644),
    .B(_07667_),
    .X(_02003_));
 sg13g2_nand3_1 _26835_ (.B(net445),
    .C(net111),
    .A(_06748_),
    .Y(_07668_));
 sg13g2_nand2_1 _26836_ (.Y(_07669_),
    .A(net445),
    .B(net111));
 sg13g2_nand2_1 _26837_ (.Y(_07670_),
    .A(_04925_),
    .B(_07669_));
 sg13g2_a21oi_1 _26838_ (.A1(_07668_),
    .A2(_07670_),
    .Y(_02008_),
    .B1(net561));
 sg13g2_nand3_1 _26839_ (.B(_04927_),
    .C(net111),
    .A(net1027),
    .Y(_07671_));
 sg13g2_nand2_1 _26840_ (.Y(_07672_),
    .A(\cpu.gpio.r_uart_rx_src[1] ),
    .B(_07669_));
 sg13g2_a21oi_1 _26841_ (.A1(_07671_),
    .A2(_07672_),
    .Y(_02009_),
    .B1(_07647_));
 sg13g2_nand3_1 _26842_ (.B(_04927_),
    .C(net111),
    .A(_10075_),
    .Y(_07673_));
 sg13g2_nand2_1 _26843_ (.Y(_07674_),
    .A(\cpu.gpio.r_uart_rx_src[2] ),
    .B(_07669_));
 sg13g2_a21oi_1 _26844_ (.A1(_07673_),
    .A2(_07674_),
    .Y(_02010_),
    .B1(_07647_));
 sg13g2_and2_1 _26845_ (.A(\cpu.i_wstrobe_d ),
    .B(_00314_),
    .X(_02267_));
 sg13g2_a21oi_1 _26846_ (.A1(_06360_),
    .A2(_06372_),
    .Y(_02268_),
    .B1(_06383_));
 sg13g2_xor2_1 _26847_ (.B(_06367_),
    .A(_06356_),
    .X(_07675_));
 sg13g2_nor2_1 _26848_ (.A(_06383_),
    .B(_07675_),
    .Y(_02269_));
 sg13g2_nor4_1 _26849_ (.A(net695),
    .B(_10115_),
    .C(_10061_),
    .D(_04906_),
    .Y(_07676_));
 sg13g2_mux2_1 _26850_ (.A0(_05345_),
    .A1(net538),
    .S(_07676_),
    .X(_07677_));
 sg13g2_xnor2_1 _26851_ (.Y(_07678_),
    .A(\cpu.intr.r_clock_cmp[12] ),
    .B(_10200_));
 sg13g2_xnor2_1 _26852_ (.Y(_07679_),
    .A(\cpu.intr.r_clock_cmp[14] ),
    .B(_10210_));
 sg13g2_xnor2_1 _26853_ (.Y(_07680_),
    .A(\cpu.intr.r_clock_cmp[11] ),
    .B(_10193_));
 sg13g2_xnor2_1 _26854_ (.Y(_07681_),
    .A(\cpu.intr.r_clock_cmp[29] ),
    .B(_05275_));
 sg13g2_nand4_1 _26855_ (.B(_07679_),
    .C(_07680_),
    .A(_07678_),
    .Y(_07682_),
    .D(_07681_));
 sg13g2_xnor2_1 _26856_ (.Y(_07683_),
    .A(\cpu.intr.r_clock_cmp[4] ),
    .B(_10153_));
 sg13g2_xnor2_1 _26857_ (.Y(_07684_),
    .A(\cpu.intr.r_clock_cmp[26] ),
    .B(_05177_));
 sg13g2_xnor2_1 _26858_ (.Y(_07685_),
    .A(\cpu.intr.r_clock_cmp[6] ),
    .B(_10165_));
 sg13g2_xnor2_1 _26859_ (.Y(_07686_),
    .A(\cpu.intr.r_clock_cmp[19] ),
    .B(_05531_));
 sg13g2_nand4_1 _26860_ (.B(_07684_),
    .C(_07685_),
    .A(_07683_),
    .Y(_07687_),
    .D(_07686_));
 sg13g2_xnor2_1 _26861_ (.Y(_07688_),
    .A(\cpu.intr.r_clock_cmp[30] ),
    .B(_05286_));
 sg13g2_xnor2_1 _26862_ (.Y(_07689_),
    .A(\cpu.intr.r_clock_cmp[10] ),
    .B(_10188_));
 sg13g2_xnor2_1 _26863_ (.Y(_07690_),
    .A(\cpu.intr.r_clock_cmp[22] ),
    .B(_05737_));
 sg13g2_xnor2_1 _26864_ (.Y(_07691_),
    .A(\cpu.intr.r_clock_cmp[1] ),
    .B(_10129_));
 sg13g2_nand4_1 _26865_ (.B(_07689_),
    .C(_07690_),
    .A(_07688_),
    .Y(_07692_),
    .D(_07691_));
 sg13g2_xnor2_1 _26866_ (.Y(_07693_),
    .A(\cpu.intr.r_clock_cmp[24] ),
    .B(_05761_));
 sg13g2_xnor2_1 _26867_ (.Y(_07694_),
    .A(\cpu.intr.r_clock_cmp[13] ),
    .B(_10206_));
 sg13g2_xnor2_1 _26868_ (.Y(_07695_),
    .A(\cpu.intr.r_clock_cmp[9] ),
    .B(_10183_));
 sg13g2_xnor2_1 _26869_ (.Y(_07696_),
    .A(\cpu.intr.r_clock_cmp[2] ),
    .B(_10142_));
 sg13g2_nand4_1 _26870_ (.B(_07694_),
    .C(_07695_),
    .A(_07693_),
    .Y(_07697_),
    .D(_07696_));
 sg13g2_nor4_1 _26871_ (.A(_07682_),
    .B(_07687_),
    .C(_07692_),
    .D(_07697_),
    .Y(_07698_));
 sg13g2_xnor2_1 _26872_ (.Y(_07699_),
    .A(\cpu.intr.r_clock_cmp[23] ),
    .B(_05111_));
 sg13g2_xnor2_1 _26873_ (.Y(_07700_),
    .A(\cpu.intr.r_clock_cmp[7] ),
    .B(_10171_));
 sg13g2_xnor2_1 _26874_ (.Y(_07701_),
    .A(\cpu.intr.r_clock_cmp[27] ),
    .B(_05218_));
 sg13g2_xnor2_1 _26875_ (.Y(_07702_),
    .A(\cpu.intr.r_clock_cmp[3] ),
    .B(_10147_));
 sg13g2_nand4_1 _26876_ (.B(_07700_),
    .C(_07701_),
    .A(_07699_),
    .Y(_07703_),
    .D(_07702_));
 sg13g2_xnor2_1 _26877_ (.Y(_07704_),
    .A(\cpu.intr.r_clock_cmp[31] ),
    .B(_05318_));
 sg13g2_xnor2_1 _26878_ (.Y(_07705_),
    .A(\cpu.intr.r_clock_cmp[17] ),
    .B(_05352_));
 sg13g2_xnor2_1 _26879_ (.Y(_07706_),
    .A(\cpu.intr.r_clock_cmp[25] ),
    .B(_05775_));
 sg13g2_xnor2_1 _26880_ (.Y(_07707_),
    .A(\cpu.intr.r_clock_cmp[28] ),
    .B(_05233_));
 sg13g2_nand4_1 _26881_ (.B(_07705_),
    .C(_07706_),
    .A(_07704_),
    .Y(_07708_),
    .D(_07707_));
 sg13g2_xnor2_1 _26882_ (.Y(_07709_),
    .A(\cpu.intr.r_clock_cmp[18] ),
    .B(_05461_));
 sg13g2_xnor2_1 _26883_ (.Y(_07710_),
    .A(\cpu.intr.r_clock_cmp[0] ),
    .B(_10128_));
 sg13g2_xnor2_1 _26884_ (.Y(_07711_),
    .A(\cpu.intr.r_clock_cmp[16] ),
    .B(_04972_));
 sg13g2_xnor2_1 _26885_ (.Y(_07712_),
    .A(\cpu.intr.r_clock_cmp[8] ),
    .B(_10175_));
 sg13g2_nand4_1 _26886_ (.B(_07710_),
    .C(_07711_),
    .A(_07709_),
    .Y(_07713_),
    .D(_07712_));
 sg13g2_xnor2_1 _26887_ (.Y(_07714_),
    .A(\cpu.intr.r_clock_cmp[21] ),
    .B(_05621_));
 sg13g2_xnor2_1 _26888_ (.Y(_07715_),
    .A(\cpu.intr.r_clock_cmp[5] ),
    .B(_10159_));
 sg13g2_xnor2_1 _26889_ (.Y(_07716_),
    .A(\cpu.intr.r_clock_cmp[20] ),
    .B(_05558_));
 sg13g2_xnor2_1 _26890_ (.Y(_07717_),
    .A(\cpu.intr.r_clock_cmp[15] ),
    .B(_10217_));
 sg13g2_nand4_1 _26891_ (.B(_07715_),
    .C(_07716_),
    .A(_07714_),
    .Y(_07718_),
    .D(_07717_));
 sg13g2_nor4_1 _26892_ (.A(_07703_),
    .B(_07708_),
    .C(_07713_),
    .D(_07718_),
    .Y(_07719_));
 sg13g2_nand2_1 _26893_ (.Y(_07720_),
    .A(_07698_),
    .B(_07719_));
 sg13g2_a21oi_1 _26894_ (.A1(_07677_),
    .A2(_07720_),
    .Y(_02430_),
    .B1(net561));
 sg13g2_and2_1 _26895_ (.A(net171),
    .B(net397),
    .X(_07721_));
 sg13g2_buf_1 _26896_ (.A(_07721_),
    .X(_07722_));
 sg13g2_nand2_1 _26897_ (.Y(_07723_),
    .A(_06748_),
    .B(_07722_));
 sg13g2_nand2_1 _26898_ (.Y(_07724_),
    .A(net171),
    .B(_04994_));
 sg13g2_buf_1 _26899_ (.A(_07724_),
    .X(_07725_));
 sg13g2_nand2_1 _26900_ (.Y(_07726_),
    .A(\cpu.intr.r_enable[0] ),
    .B(_07725_));
 sg13g2_a21oi_1 _26901_ (.A1(_07723_),
    .A2(_07726_),
    .Y(_02479_),
    .B1(net561));
 sg13g2_nand2_1 _26902_ (.Y(_07727_),
    .A(net939),
    .B(_07722_));
 sg13g2_nand2_1 _26903_ (.Y(_07728_),
    .A(_09251_),
    .B(_07725_));
 sg13g2_a21oi_1 _26904_ (.A1(_07727_),
    .A2(_07728_),
    .Y(_02480_),
    .B1(net561));
 sg13g2_nand2_1 _26905_ (.Y(_07729_),
    .A(net1026),
    .B(_07722_));
 sg13g2_nand2_1 _26906_ (.Y(_07730_),
    .A(\cpu.intr.r_enable[2] ),
    .B(_07725_));
 sg13g2_a21oi_1 _26907_ (.A1(_07729_),
    .A2(_07730_),
    .Y(_02481_),
    .B1(net561));
 sg13g2_nand2_1 _26908_ (.Y(_07731_),
    .A(net1025),
    .B(_07722_));
 sg13g2_nand2_1 _26909_ (.Y(_07732_),
    .A(_09246_),
    .B(_07725_));
 sg13g2_buf_1 _26910_ (.A(_09351_),
    .X(_07733_));
 sg13g2_a21oi_1 _26911_ (.A1(_07731_),
    .A2(_07732_),
    .Y(_02482_),
    .B1(net560));
 sg13g2_nand2_1 _26912_ (.Y(_07734_),
    .A(net1024),
    .B(_07722_));
 sg13g2_nand2_1 _26913_ (.Y(_07735_),
    .A(_09214_),
    .B(_07725_));
 sg13g2_a21oi_1 _26914_ (.A1(_07734_),
    .A2(_07735_),
    .Y(_02483_),
    .B1(_07733_));
 sg13g2_nand2_1 _26915_ (.Y(_07736_),
    .A(net1023),
    .B(_07722_));
 sg13g2_nand2_1 _26916_ (.Y(_07737_),
    .A(_09253_),
    .B(_07725_));
 sg13g2_a21oi_1 _26917_ (.A1(_07736_),
    .A2(_07737_),
    .Y(_02484_),
    .B1(net560));
 sg13g2_nand3_1 _26918_ (.B(_10003_),
    .C(net389),
    .A(net1020),
    .Y(_07738_));
 sg13g2_nand3_1 _26919_ (.B(_10003_),
    .C(net388),
    .A(net1020),
    .Y(_07739_));
 sg13g2_nand2_1 _26920_ (.Y(_07740_),
    .A(_09991_),
    .B(_07739_));
 sg13g2_a21oi_1 _26921_ (.A1(_09245_),
    .A2(_07738_),
    .Y(_07741_),
    .B1(_07740_));
 sg13g2_nor2_1 _26922_ (.A(net562),
    .B(_07741_),
    .Y(_02485_));
 sg13g2_nor3_1 _26923_ (.A(net1114),
    .B(_09851_),
    .C(_06787_),
    .Y(_07742_));
 sg13g2_nor2b_1 _26924_ (.A(net1117),
    .B_N(_07742_),
    .Y(_07743_));
 sg13g2_nand4_1 _26925_ (.B(_09873_),
    .C(_06788_),
    .A(_09831_),
    .Y(_07744_),
    .D(_07743_));
 sg13g2_buf_1 _26926_ (.A(_07744_),
    .X(_07745_));
 sg13g2_o21ai_1 _26927_ (.B1(net764),
    .Y(_07746_),
    .A1(_06764_),
    .A2(_07745_));
 sg13g2_nor2b_1 _26928_ (.A(_09866_),
    .B_N(_09899_),
    .Y(_07747_));
 sg13g2_o21ai_1 _26929_ (.B1(net19),
    .Y(_07748_),
    .A1(_07745_),
    .A2(_07747_));
 sg13g2_nand2b_1 _26930_ (.Y(_02515_),
    .B(_07748_),
    .A_N(_07746_));
 sg13g2_nand2_1 _26931_ (.Y(_07749_),
    .A(_09833_),
    .B(\cpu.qspi.r_state[0] ));
 sg13g2_o21ai_1 _26932_ (.B1(_06764_),
    .Y(_07750_),
    .A1(_09899_),
    .A2(_07749_));
 sg13g2_nand2b_1 _26933_ (.Y(_07751_),
    .B(_07750_),
    .A_N(_07745_));
 sg13g2_nand2_1 _26934_ (.Y(_07752_),
    .A(_09899_),
    .B(_06764_));
 sg13g2_nor2_1 _26935_ (.A(net88),
    .B(_07752_),
    .Y(_07753_));
 sg13g2_o21ai_1 _26936_ (.B1(net20),
    .Y(_07754_),
    .A1(_07745_),
    .A2(_07753_));
 sg13g2_nand3_1 _26937_ (.B(_07751_),
    .C(_07754_),
    .A(net645),
    .Y(_02516_));
 sg13g2_nor2b_1 _26938_ (.A(net245),
    .B_N(_09899_),
    .Y(_07755_));
 sg13g2_buf_1 _26939_ (.A(\cpu.gpio.genblk1[3].srcs_o[11] ),
    .X(_07756_));
 sg13g2_o21ai_1 _26940_ (.B1(_07756_),
    .Y(_07757_),
    .A1(_07745_),
    .A2(_07755_));
 sg13g2_nand2b_1 _26941_ (.Y(_02517_),
    .B(_07757_),
    .A_N(_07746_));
 sg13g2_nor2_1 _26942_ (.A(\cpu.qspi.r_state[11] ),
    .B(\cpu.qspi.r_state[0] ),
    .Y(_07758_));
 sg13g2_nor4_1 _26943_ (.A(_09390_),
    .B(_09843_),
    .C(net1031),
    .D(_09844_),
    .Y(_07759_));
 sg13g2_nand3_1 _26944_ (.B(_07758_),
    .C(_07759_),
    .A(_06677_),
    .Y(_07760_));
 sg13g2_inv_1 _26945_ (.Y(_07761_),
    .A(_07760_));
 sg13g2_a21oi_1 _26946_ (.A1(_07743_),
    .A2(_07761_),
    .Y(_07762_),
    .B1(_09833_));
 sg13g2_nor2_1 _26947_ (.A(net562),
    .B(_07762_),
    .Y(_02518_));
 sg13g2_nand2_1 _26948_ (.Y(_07763_),
    .A(net1021),
    .B(_06722_));
 sg13g2_nand2_1 _26949_ (.Y(_07764_),
    .A(\cpu.qspi.r_mask[0] ),
    .B(_06725_));
 sg13g2_a21oi_1 _26950_ (.A1(_07763_),
    .A2(_07764_),
    .Y(_02519_),
    .B1(_07733_));
 sg13g2_a21oi_1 _26951_ (.A1(_04950_),
    .A2(net583),
    .Y(_07765_),
    .B1(net959));
 sg13g2_nand2_1 _26952_ (.Y(_07766_),
    .A(_06720_),
    .B(_07765_));
 sg13g2_o21ai_1 _26953_ (.B1(_09878_),
    .Y(_07767_),
    .A1(_06974_),
    .A2(_07766_));
 sg13g2_a21o_1 _26954_ (.A2(_06740_),
    .A1(\cpu.qspi.r_mask[1] ),
    .B1(_07767_),
    .X(_02520_));
 sg13g2_nor2_1 _26955_ (.A(_06974_),
    .B(_06753_),
    .Y(_07768_));
 sg13g2_a21oi_1 _26956_ (.A1(\cpu.qspi.r_mask[2] ),
    .A2(_06753_),
    .Y(_07769_),
    .B1(_07768_));
 sg13g2_nor2_1 _26957_ (.A(net562),
    .B(_07769_),
    .Y(_02521_));
 sg13g2_nand2_1 _26958_ (.Y(_07770_),
    .A(\cpu.qspi.r_quad[0] ),
    .B(_06725_));
 sg13g2_nand2_1 _26959_ (.Y(_07771_),
    .A(net1022),
    .B(_06722_));
 sg13g2_nand3_1 _26960_ (.B(_07770_),
    .C(_07771_),
    .A(net645),
    .Y(_02522_));
 sg13g2_nor2_1 _26961_ (.A(_06970_),
    .B(_07766_),
    .Y(_07772_));
 sg13g2_a21oi_1 _26962_ (.A1(\cpu.qspi.r_quad[1] ),
    .A2(_06740_),
    .Y(_07773_),
    .B1(_07772_));
 sg13g2_nor2_1 _26963_ (.A(net562),
    .B(_07773_),
    .Y(_02523_));
 sg13g2_nand2_1 _26964_ (.Y(_07774_),
    .A(_06970_),
    .B(_06750_));
 sg13g2_o21ai_1 _26965_ (.B1(_07774_),
    .Y(_07775_),
    .A1(\cpu.qspi.r_quad[2] ),
    .A2(_06750_));
 sg13g2_nand2_1 _26966_ (.Y(_02524_),
    .A(net675),
    .B(_07775_));
 sg13g2_nand2b_1 _26967_ (.Y(_07776_),
    .B(_06720_),
    .A_N(_04920_));
 sg13g2_buf_1 _26968_ (.A(_07776_),
    .X(_07777_));
 sg13g2_nor2_1 _26969_ (.A(net1029),
    .B(_07777_),
    .Y(_07778_));
 sg13g2_nor2b_1 _26970_ (.A(\cpu.qspi.r_rom_mode[0] ),
    .B_N(_07777_),
    .Y(_07779_));
 sg13g2_o21ai_1 _26971_ (.B1(net675),
    .Y(_02537_),
    .A1(_07778_),
    .A2(_07779_));
 sg13g2_nor2_1 _26972_ (.A(net1027),
    .B(_07777_),
    .Y(_07780_));
 sg13g2_nor2b_1 _26973_ (.A(_09861_),
    .B_N(_07777_),
    .Y(_07781_));
 sg13g2_o21ai_1 _26974_ (.B1(net675),
    .Y(_02538_),
    .A1(_07780_),
    .A2(_07781_));
 sg13g2_nor2_1 _26975_ (.A(_11882_),
    .B(net1117),
    .Y(_07782_));
 sg13g2_nand3_1 _26976_ (.B(_07758_),
    .C(_07782_),
    .A(_06676_),
    .Y(_07783_));
 sg13g2_nand2_1 _26977_ (.Y(_07784_),
    .A(_07758_),
    .B(_07783_));
 sg13g2_a21o_1 _26978_ (.A2(_06762_),
    .A1(_06761_),
    .B1(_11883_),
    .X(_07785_));
 sg13g2_nor3_1 _26979_ (.A(_09843_),
    .B(_09901_),
    .C(_09854_),
    .Y(_07786_));
 sg13g2_nand4_1 _26980_ (.B(_07742_),
    .C(_07785_),
    .A(_09831_),
    .Y(_07787_),
    .D(_07786_));
 sg13g2_buf_1 _26981_ (.A(_07787_),
    .X(_07788_));
 sg13g2_mux2_1 _26982_ (.A0(_07784_),
    .A1(net3),
    .S(_07788_),
    .X(_07789_));
 sg13g2_and2_1 _26983_ (.A(net644),
    .B(_07789_),
    .X(_02539_));
 sg13g2_nor2b_1 _26984_ (.A(net6),
    .B_N(_07788_),
    .Y(_07790_));
 sg13g2_o21ai_1 _26985_ (.B1(_11880_),
    .Y(_07791_),
    .A1(_09869_),
    .A2(_07783_));
 sg13g2_nor2_1 _26986_ (.A(_07788_),
    .B(_07791_),
    .Y(_07792_));
 sg13g2_nor3_1 _26987_ (.A(net618),
    .B(_07790_),
    .C(_07792_),
    .Y(_02540_));
 sg13g2_nor2_1 _26988_ (.A(_09285_),
    .B(_06984_),
    .Y(_07793_));
 sg13g2_a221oi_1 _26989_ (.B2(_09332_),
    .C1(_07793_),
    .B1(net419),
    .A1(_09195_),
    .Y(_07794_),
    .A2(net117));
 sg13g2_buf_2 _26990_ (.A(_07794_),
    .X(_07795_));
 sg13g2_nand3_1 _26991_ (.B(net1038),
    .C(_07795_),
    .A(_09299_),
    .Y(_07796_));
 sg13g2_o21ai_1 _26992_ (.B1(_07796_),
    .Y(_07797_),
    .A1(_09299_),
    .A2(_07795_));
 sg13g2_nand2_1 _26993_ (.Y(_02546_),
    .A(net675),
    .B(_07797_));
 sg13g2_nand2_1 _26994_ (.Y(_07798_),
    .A(_09299_),
    .B(_11923_));
 sg13g2_a21oi_1 _26995_ (.A1(_07795_),
    .A2(_07798_),
    .Y(_07799_),
    .B1(_09300_));
 sg13g2_inv_1 _26996_ (.Y(_07800_),
    .A(_09299_));
 sg13g2_and4_1 _26997_ (.A(_07800_),
    .B(_09300_),
    .C(_11923_),
    .D(_07795_),
    .X(_07801_));
 sg13g2_o21ai_1 _26998_ (.B1(net675),
    .Y(_02547_),
    .A1(_07799_),
    .A2(_07801_));
 sg13g2_nor2_1 _26999_ (.A(_09299_),
    .B(_09300_),
    .Y(_07802_));
 sg13g2_or2_1 _27000_ (.X(_07803_),
    .B(_07802_),
    .A(_00224_));
 sg13g2_a21oi_1 _27001_ (.A1(_07795_),
    .A2(_07803_),
    .Y(_07804_),
    .B1(\cpu.spi.r_bits[2] ));
 sg13g2_and4_1 _27002_ (.A(\cpu.spi.r_bits[2] ),
    .B(_11923_),
    .C(_07802_),
    .D(_07795_),
    .X(_07805_));
 sg13g2_o21ai_1 _27003_ (.B1(_06729_),
    .Y(_02548_),
    .A1(_07804_),
    .A2(_07805_));
 sg13g2_nor2_1 _27004_ (.A(net858),
    .B(_04943_),
    .Y(_07806_));
 sg13g2_nand4_1 _27005_ (.B(_09344_),
    .C(_10120_),
    .A(net733),
    .Y(_07807_),
    .D(_07806_));
 sg13g2_buf_1 _27006_ (.A(_07807_),
    .X(_07808_));
 sg13g2_mux2_1 _27007_ (.A0(net1029),
    .A1(\cpu.spi.r_clk_count[0][0] ),
    .S(net110),
    .X(_07809_));
 sg13g2_and2_1 _27008_ (.A(_07656_),
    .B(_07809_),
    .X(_02549_));
 sg13g2_nand2_1 _27009_ (.Y(_07810_),
    .A(\cpu.spi.r_clk_count[0][1] ),
    .B(net110));
 sg13g2_o21ai_1 _27010_ (.B1(_07810_),
    .Y(_07811_),
    .A1(net887),
    .A2(net110));
 sg13g2_and2_1 _27011_ (.A(_07656_),
    .B(_07811_),
    .X(_02550_));
 sg13g2_mux2_1 _27012_ (.A0(net1020),
    .A1(\cpu.spi.r_clk_count[0][2] ),
    .S(net110),
    .X(_07812_));
 sg13g2_and2_1 _27013_ (.A(net644),
    .B(_07812_),
    .X(_02551_));
 sg13g2_mux2_1 _27014_ (.A0(net1113),
    .A1(\cpu.spi.r_clk_count[0][3] ),
    .S(net110),
    .X(_07813_));
 sg13g2_and2_1 _27015_ (.A(net644),
    .B(_07813_),
    .X(_02552_));
 sg13g2_buf_1 _27016_ (.A(net764),
    .X(_07814_));
 sg13g2_mux2_1 _27017_ (.A0(_10085_),
    .A1(\cpu.spi.r_clk_count[0][4] ),
    .S(net110),
    .X(_07815_));
 sg13g2_and2_1 _27018_ (.A(net643),
    .B(_07815_),
    .X(_02553_));
 sg13g2_mux2_1 _27019_ (.A0(net1023),
    .A1(\cpu.spi.r_clk_count[0][5] ),
    .S(net110),
    .X(_07816_));
 sg13g2_and2_1 _27020_ (.A(net643),
    .B(_07816_),
    .X(_02554_));
 sg13g2_mux2_1 _27021_ (.A0(_10098_),
    .A1(\cpu.spi.r_clk_count[0][6] ),
    .S(_07808_),
    .X(_07817_));
 sg13g2_and2_1 _27022_ (.A(net643),
    .B(_07817_),
    .X(_02555_));
 sg13g2_mux2_1 _27023_ (.A0(_10103_),
    .A1(\cpu.spi.r_clk_count[0][7] ),
    .S(net110),
    .X(_07818_));
 sg13g2_and2_1 _27024_ (.A(_07814_),
    .B(_07818_),
    .X(_02556_));
 sg13g2_nand4_1 _27025_ (.B(_09344_),
    .C(_10120_),
    .A(net595),
    .Y(_07819_),
    .D(_07806_));
 sg13g2_buf_2 _27026_ (.A(_07819_),
    .X(_07820_));
 sg13g2_nand2_1 _27027_ (.Y(_07821_),
    .A(\cpu.spi.r_clk_count[1][0] ),
    .B(_07820_));
 sg13g2_and4_1 _27028_ (.A(net595),
    .B(_09344_),
    .C(_10120_),
    .D(_07806_),
    .X(_07822_));
 sg13g2_buf_2 _27029_ (.A(_07822_),
    .X(_07823_));
 sg13g2_nand2_1 _27030_ (.Y(_07824_),
    .A(net799),
    .B(_07823_));
 sg13g2_a21oi_1 _27031_ (.A1(_07821_),
    .A2(_07824_),
    .Y(_02557_),
    .B1(net560));
 sg13g2_nand2_1 _27032_ (.Y(_07825_),
    .A(\cpu.spi.r_clk_count[1][1] ),
    .B(_07820_));
 sg13g2_nand2_1 _27033_ (.Y(_07826_),
    .A(_10070_),
    .B(_07823_));
 sg13g2_a21oi_1 _27034_ (.A1(_07825_),
    .A2(_07826_),
    .Y(_02558_),
    .B1(net560));
 sg13g2_nand2_1 _27035_ (.Y(_07827_),
    .A(\cpu.spi.r_clk_count[1][2] ),
    .B(_07820_));
 sg13g2_nand2_1 _27036_ (.Y(_07828_),
    .A(net1026),
    .B(_07823_));
 sg13g2_a21oi_1 _27037_ (.A1(_07827_),
    .A2(_07828_),
    .Y(_02559_),
    .B1(net560));
 sg13g2_nand2_1 _27038_ (.Y(_07829_),
    .A(\cpu.spi.r_clk_count[1][3] ),
    .B(_07820_));
 sg13g2_nand2_1 _27039_ (.Y(_07830_),
    .A(net1025),
    .B(_07823_));
 sg13g2_a21oi_1 _27040_ (.A1(_07829_),
    .A2(_07830_),
    .Y(_02560_),
    .B1(net560));
 sg13g2_nand2_1 _27041_ (.Y(_07831_),
    .A(\cpu.spi.r_clk_count[1][4] ),
    .B(_07820_));
 sg13g2_nand2_1 _27042_ (.Y(_07832_),
    .A(net1024),
    .B(_07823_));
 sg13g2_a21oi_1 _27043_ (.A1(_07831_),
    .A2(_07832_),
    .Y(_02561_),
    .B1(net560));
 sg13g2_nand2_1 _27044_ (.Y(_07833_),
    .A(\cpu.spi.r_clk_count[1][5] ),
    .B(_07820_));
 sg13g2_nand2_1 _27045_ (.Y(_07834_),
    .A(net1023),
    .B(_07823_));
 sg13g2_a21oi_1 _27046_ (.A1(_07833_),
    .A2(_07834_),
    .Y(_02562_),
    .B1(net560));
 sg13g2_nand2_1 _27047_ (.Y(_07835_),
    .A(\cpu.spi.r_clk_count[1][6] ),
    .B(_07820_));
 sg13g2_nand2_1 _27048_ (.Y(_07836_),
    .A(_10098_),
    .B(_07823_));
 sg13g2_buf_1 _27049_ (.A(_09351_),
    .X(_07837_));
 sg13g2_a21oi_1 _27050_ (.A1(_07835_),
    .A2(_07836_),
    .Y(_02563_),
    .B1(net559));
 sg13g2_nand2_1 _27051_ (.Y(_07838_),
    .A(\cpu.spi.r_clk_count[1][7] ),
    .B(_07820_));
 sg13g2_nand2_1 _27052_ (.Y(_07839_),
    .A(_10104_),
    .B(_07823_));
 sg13g2_a21oi_1 _27053_ (.A1(_07838_),
    .A2(_07839_),
    .Y(_02564_),
    .B1(net559));
 sg13g2_nor3_1 _27054_ (.A(net862),
    .B(net734),
    .C(_04943_),
    .Y(_07840_));
 sg13g2_nand3_1 _27055_ (.B(_10120_),
    .C(_07840_),
    .A(_09344_),
    .Y(_07841_));
 sg13g2_buf_1 _27056_ (.A(_07841_),
    .X(_07842_));
 sg13g2_mux2_1 _27057_ (.A0(_10048_),
    .A1(_04965_),
    .S(net109),
    .X(_07843_));
 sg13g2_and2_1 _27058_ (.A(_07814_),
    .B(_07843_),
    .X(_02565_));
 sg13g2_nand2_1 _27059_ (.Y(_07844_),
    .A(_05337_),
    .B(net109));
 sg13g2_o21ai_1 _27060_ (.B1(_07844_),
    .Y(_07845_),
    .A1(net887),
    .A2(net109));
 sg13g2_and2_1 _27061_ (.A(net643),
    .B(_07845_),
    .X(_02566_));
 sg13g2_mux2_1 _27062_ (.A0(net1020),
    .A1(_05439_),
    .S(net109),
    .X(_07846_));
 sg13g2_and2_1 _27063_ (.A(net643),
    .B(_07846_),
    .X(_02567_));
 sg13g2_mux2_1 _27064_ (.A0(net1113),
    .A1(_05508_),
    .S(net109),
    .X(_07847_));
 sg13g2_and2_1 _27065_ (.A(net643),
    .B(_07847_),
    .X(_02568_));
 sg13g2_mux2_1 _27066_ (.A0(_10085_),
    .A1(_05586_),
    .S(net109),
    .X(_07848_));
 sg13g2_and2_1 _27067_ (.A(net643),
    .B(_07848_),
    .X(_02569_));
 sg13g2_mux2_1 _27068_ (.A0(_10091_),
    .A1(_05652_),
    .S(net109),
    .X(_07849_));
 sg13g2_and2_1 _27069_ (.A(net643),
    .B(_07849_),
    .X(_02570_));
 sg13g2_mux2_1 _27070_ (.A0(_10097_),
    .A1(_05741_),
    .S(net109),
    .X(_07850_));
 sg13g2_and2_1 _27071_ (.A(net659),
    .B(_07850_),
    .X(_02571_));
 sg13g2_mux2_1 _27072_ (.A0(_10103_),
    .A1(_05079_),
    .S(_07842_),
    .X(_07851_));
 sg13g2_and2_1 _27073_ (.A(net659),
    .B(_07851_),
    .X(_02572_));
 sg13g2_o21ai_1 _27074_ (.B1(_09265_),
    .Y(_07852_),
    .A1(net473),
    .A2(_09282_));
 sg13g2_nor4_1 _27075_ (.A(_09283_),
    .B(\cpu.spi.r_state[5] ),
    .C(net1121),
    .D(_11919_),
    .Y(_07853_));
 sg13g2_buf_1 _27076_ (.A(_07853_),
    .X(_07854_));
 sg13g2_nor2_1 _27077_ (.A(_06948_),
    .B(net473),
    .Y(_07855_));
 sg13g2_a22oi_1 _27078_ (.Y(_07856_),
    .B1(_07855_),
    .B2(_09354_),
    .A2(_07854_),
    .A1(_06944_));
 sg13g2_nand3_1 _27079_ (.B(_07852_),
    .C(_07856_),
    .A(_06943_),
    .Y(_07857_));
 sg13g2_buf_1 _27080_ (.A(_07857_),
    .X(_07858_));
 sg13g2_buf_1 _27081_ (.A(_07858_),
    .X(_07859_));
 sg13g2_nand2b_1 _27082_ (.Y(_07860_),
    .B(net656),
    .A_N(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_o21ai_1 _27083_ (.B1(_07860_),
    .Y(_07861_),
    .A1(net656),
    .A2(_04965_));
 sg13g2_mux2_1 _27084_ (.A0(\cpu.spi.r_clk_count[0][0] ),
    .A1(\cpu.spi.r_clk_count[1][0] ),
    .S(net655),
    .X(_07862_));
 sg13g2_nor2_1 _27085_ (.A(net657),
    .B(_07862_),
    .Y(_07863_));
 sg13g2_a21oi_1 _27086_ (.A1(net651),
    .A2(_07861_),
    .Y(_07864_),
    .B1(_07863_));
 sg13g2_nand2_1 _27087_ (.Y(_07865_),
    .A(_06948_),
    .B(_07853_));
 sg13g2_inv_1 _27088_ (.Y(_07866_),
    .A(_07865_));
 sg13g2_buf_1 _27089_ (.A(_07866_),
    .X(_07867_));
 sg13g2_nor2_1 _27090_ (.A(_11953_),
    .B(_04965_),
    .Y(_07868_));
 sg13g2_a21oi_1 _27091_ (.A1(_11953_),
    .A2(_00312_),
    .Y(_07869_),
    .B1(_07868_));
 sg13g2_nand2_1 _27092_ (.Y(_07870_),
    .A(_11950_),
    .B(_00311_));
 sg13g2_o21ai_1 _27093_ (.B1(_07870_),
    .Y(_07871_),
    .A1(net1001),
    .A2(_04955_));
 sg13g2_nor2_1 _27094_ (.A(_11947_),
    .B(_07871_),
    .Y(_07872_));
 sg13g2_a21oi_1 _27095_ (.A1(net1002),
    .A2(_07869_),
    .Y(_07873_),
    .B1(_07872_));
 sg13g2_nand2_1 _27096_ (.Y(_07874_),
    .A(net418),
    .B(_07873_));
 sg13g2_nor2_1 _27097_ (.A(_09185_),
    .B(net642),
    .Y(_07875_));
 sg13g2_mux2_1 _27098_ (.A0(_09185_),
    .A1(_07873_),
    .S(_09263_),
    .X(_07876_));
 sg13g2_nor2_1 _27099_ (.A(_09196_),
    .B(_07876_),
    .Y(_07877_));
 sg13g2_a21oi_1 _27100_ (.A1(_07874_),
    .A2(_07875_),
    .Y(_07878_),
    .B1(_07877_));
 sg13g2_nor2_1 _27101_ (.A(_07867_),
    .B(_07878_),
    .Y(_07879_));
 sg13g2_a21oi_1 _27102_ (.A1(_07864_),
    .A2(net484),
    .Y(_07880_),
    .B1(_07879_));
 sg13g2_nor2_1 _27103_ (.A(net59),
    .B(_07880_),
    .Y(_07881_));
 sg13g2_a21oi_1 _27104_ (.A1(_09185_),
    .A2(net59),
    .Y(_07882_),
    .B1(_07881_));
 sg13g2_nor2_1 _27105_ (.A(net562),
    .B(_07882_),
    .Y(_02573_));
 sg13g2_mux2_1 _27106_ (.A0(\cpu.spi.r_clk_count[0][1] ),
    .A1(\cpu.spi.r_clk_count[1][1] ),
    .S(net734),
    .X(_07883_));
 sg13g2_nor2_1 _27107_ (.A(_11926_),
    .B(_07883_),
    .Y(_07884_));
 sg13g2_mux2_1 _27108_ (.A0(_05337_),
    .A1(\cpu.spi.r_clk_count[0][1] ),
    .S(net734),
    .X(_07885_));
 sg13g2_nor2_1 _27109_ (.A(net862),
    .B(_07885_),
    .Y(_07886_));
 sg13g2_o21ai_1 _27110_ (.B1(_07866_),
    .Y(_07887_),
    .A1(_07884_),
    .A2(_07886_));
 sg13g2_and3_1 _27111_ (.X(_07888_),
    .A(_09185_),
    .B(_09265_),
    .C(_07887_));
 sg13g2_o21ai_1 _27112_ (.B1(_09186_),
    .Y(_07889_),
    .A1(_07859_),
    .A2(_07888_));
 sg13g2_nor2_1 _27113_ (.A(net732),
    .B(_05337_),
    .Y(_07890_));
 sg13g2_a21oi_1 _27114_ (.A1(net732),
    .A2(_00095_),
    .Y(_07891_),
    .B1(_07890_));
 sg13g2_nand2_1 _27115_ (.Y(_07892_),
    .A(net856),
    .B(_00094_));
 sg13g2_o21ai_1 _27116_ (.B1(_07892_),
    .Y(_07893_),
    .A1(net732),
    .A2(_05335_));
 sg13g2_nor2_1 _27117_ (.A(net857),
    .B(_07893_),
    .Y(_07894_));
 sg13g2_a21oi_1 _27118_ (.A1(net857),
    .A2(_07891_),
    .Y(_07895_),
    .B1(_07894_));
 sg13g2_nor2_1 _27119_ (.A(net143),
    .B(_09187_),
    .Y(_07896_));
 sg13g2_a21oi_1 _27120_ (.A1(net143),
    .A2(_07895_),
    .Y(_07897_),
    .B1(_07896_));
 sg13g2_nand2_1 _27121_ (.Y(_07898_),
    .A(_09185_),
    .B(_09186_));
 sg13g2_or2_1 _27122_ (.X(_07899_),
    .B(_09186_),
    .A(_09185_));
 sg13g2_a221oi_1 _27123_ (.B2(_07899_),
    .C1(_07854_),
    .B1(_07898_),
    .A1(net418),
    .Y(_07900_),
    .A2(_07895_));
 sg13g2_a221oi_1 _27124_ (.B2(net1037),
    .C1(_07900_),
    .B1(_07897_),
    .A1(_06948_),
    .Y(_07901_),
    .A2(net642));
 sg13g2_nor2_1 _27125_ (.A(_07858_),
    .B(_07901_),
    .Y(_07902_));
 sg13g2_nand2_1 _27126_ (.Y(_07903_),
    .A(_07887_),
    .B(_07902_));
 sg13g2_a21oi_1 _27127_ (.A1(_07889_),
    .A2(_07903_),
    .Y(_02574_),
    .B1(net559));
 sg13g2_nand2b_1 _27128_ (.Y(_07904_),
    .B(net655),
    .A_N(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_o21ai_1 _27129_ (.B1(_07904_),
    .Y(_07905_),
    .A1(net656),
    .A2(_05439_));
 sg13g2_mux2_1 _27130_ (.A0(\cpu.spi.r_clk_count[0][2] ),
    .A1(\cpu.spi.r_clk_count[1][2] ),
    .S(net655),
    .X(_07906_));
 sg13g2_nor2_1 _27131_ (.A(net657),
    .B(_07906_),
    .Y(_07907_));
 sg13g2_a21oi_1 _27132_ (.A1(net651),
    .A2(_07905_),
    .Y(_07908_),
    .B1(_07907_));
 sg13g2_nor2_1 _27133_ (.A(net856),
    .B(_05439_),
    .Y(_07909_));
 sg13g2_a21oi_1 _27134_ (.A1(net856),
    .A2(_00105_),
    .Y(_07910_),
    .B1(_07909_));
 sg13g2_nand2_1 _27135_ (.Y(_07911_),
    .A(net1001),
    .B(_00104_));
 sg13g2_o21ai_1 _27136_ (.B1(_07911_),
    .Y(_07912_),
    .A1(net855),
    .A2(_05434_));
 sg13g2_nor2_1 _27137_ (.A(net1002),
    .B(_07912_),
    .Y(_07913_));
 sg13g2_a21oi_1 _27138_ (.A1(net857),
    .A2(_07910_),
    .Y(_07914_),
    .B1(_07913_));
 sg13g2_nand2_1 _27139_ (.Y(_07915_),
    .A(net418),
    .B(_07914_));
 sg13g2_xnor2_1 _27140_ (.Y(_07916_),
    .A(\cpu.spi.r_count[2] ),
    .B(_09187_));
 sg13g2_nor2_1 _27141_ (.A(net642),
    .B(_07916_),
    .Y(_07917_));
 sg13g2_or2_1 _27142_ (.X(_07918_),
    .B(_07916_),
    .A(net143));
 sg13g2_o21ai_1 _27143_ (.B1(_07918_),
    .Y(_07919_),
    .A1(net117),
    .A2(_07914_));
 sg13g2_a22oi_1 _27144_ (.Y(_07920_),
    .B1(_07919_),
    .B2(net1037),
    .A2(_07917_),
    .A1(_07915_));
 sg13g2_nor2_1 _27145_ (.A(net484),
    .B(_07920_),
    .Y(_07921_));
 sg13g2_a21oi_1 _27146_ (.A1(net484),
    .A2(_07908_),
    .Y(_07922_),
    .B1(_07921_));
 sg13g2_nor2_1 _27147_ (.A(net59),
    .B(_07922_),
    .Y(_07923_));
 sg13g2_a21oi_1 _27148_ (.A1(\cpu.spi.r_count[2] ),
    .A2(net59),
    .Y(_07924_),
    .B1(_07923_));
 sg13g2_nor2_1 _27149_ (.A(net562),
    .B(_07924_),
    .Y(_02575_));
 sg13g2_buf_1 _27150_ (.A(_06734_),
    .X(_07925_));
 sg13g2_nand2b_1 _27151_ (.Y(_07926_),
    .B(net655),
    .A_N(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_o21ai_1 _27152_ (.B1(_07926_),
    .Y(_07927_),
    .A1(net656),
    .A2(_05508_));
 sg13g2_mux2_1 _27153_ (.A0(\cpu.spi.r_clk_count[0][3] ),
    .A1(\cpu.spi.r_clk_count[1][3] ),
    .S(net655),
    .X(_07928_));
 sg13g2_nor2_1 _27154_ (.A(net735),
    .B(_07928_),
    .Y(_07929_));
 sg13g2_a21oi_1 _27155_ (.A1(net651),
    .A2(_07927_),
    .Y(_07930_),
    .B1(_07929_));
 sg13g2_xor2_1 _27156_ (.B(_09188_),
    .A(_09184_),
    .X(_07931_));
 sg13g2_nor2_1 _27157_ (.A(net642),
    .B(_07931_),
    .Y(_07932_));
 sg13g2_nor2_1 _27158_ (.A(net856),
    .B(_05508_),
    .Y(_07933_));
 sg13g2_a21oi_1 _27159_ (.A1(net856),
    .A2(_00115_),
    .Y(_07934_),
    .B1(_07933_));
 sg13g2_nand2_1 _27160_ (.Y(_07935_),
    .A(net1001),
    .B(_00114_));
 sg13g2_o21ai_1 _27161_ (.B1(_07935_),
    .Y(_07936_),
    .A1(net855),
    .A2(_05507_));
 sg13g2_nor2_1 _27162_ (.A(net1002),
    .B(_07936_),
    .Y(_07937_));
 sg13g2_a21oi_1 _27163_ (.A1(net857),
    .A2(_07934_),
    .Y(_07938_),
    .B1(_07937_));
 sg13g2_nand2_1 _27164_ (.Y(_07939_),
    .A(net473),
    .B(_07938_));
 sg13g2_or2_1 _27165_ (.X(_07940_),
    .B(_07931_),
    .A(net143));
 sg13g2_o21ai_1 _27166_ (.B1(_07940_),
    .Y(_07941_),
    .A1(net117),
    .A2(_07938_));
 sg13g2_a22oi_1 _27167_ (.Y(_07942_),
    .B1(_07941_),
    .B2(net1037),
    .A2(_07939_),
    .A1(_07932_));
 sg13g2_nor2_1 _27168_ (.A(net484),
    .B(_07942_),
    .Y(_07943_));
 sg13g2_a21oi_1 _27169_ (.A1(net484),
    .A2(_07930_),
    .Y(_07944_),
    .B1(_07943_));
 sg13g2_nor2_1 _27170_ (.A(_07858_),
    .B(_07944_),
    .Y(_07945_));
 sg13g2_a21oi_1 _27171_ (.A1(_09184_),
    .A2(net59),
    .Y(_07946_),
    .B1(_07945_));
 sg13g2_nor2_1 _27172_ (.A(net558),
    .B(_07946_),
    .Y(_02576_));
 sg13g2_nand2b_1 _27173_ (.Y(_07947_),
    .B(net655),
    .A_N(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_o21ai_1 _27174_ (.B1(_07947_),
    .Y(_07948_),
    .A1(net656),
    .A2(_05586_));
 sg13g2_mux2_1 _27175_ (.A0(\cpu.spi.r_clk_count[0][4] ),
    .A1(\cpu.spi.r_clk_count[1][4] ),
    .S(net655),
    .X(_07949_));
 sg13g2_nor2_1 _27176_ (.A(net735),
    .B(_07949_),
    .Y(_07950_));
 sg13g2_a21oi_1 _27177_ (.A1(net657),
    .A2(_07948_),
    .Y(_07951_),
    .B1(_07950_));
 sg13g2_nor2_1 _27178_ (.A(_09184_),
    .B(_09188_),
    .Y(_07952_));
 sg13g2_xnor2_1 _27179_ (.Y(_07953_),
    .A(\cpu.spi.r_count[4] ),
    .B(_07952_));
 sg13g2_nor2_1 _27180_ (.A(net642),
    .B(_07953_),
    .Y(_07954_));
 sg13g2_nor2_1 _27181_ (.A(net855),
    .B(_05586_),
    .Y(_07955_));
 sg13g2_a21oi_1 _27182_ (.A1(net856),
    .A2(_00126_),
    .Y(_07956_),
    .B1(_07955_));
 sg13g2_nand2_1 _27183_ (.Y(_07957_),
    .A(net1001),
    .B(_00125_));
 sg13g2_o21ai_1 _27184_ (.B1(_07957_),
    .Y(_07958_),
    .A1(net855),
    .A2(_05585_));
 sg13g2_nor2_1 _27185_ (.A(net1002),
    .B(_07958_),
    .Y(_07959_));
 sg13g2_a21oi_1 _27186_ (.A1(net857),
    .A2(_07956_),
    .Y(_07960_),
    .B1(_07959_));
 sg13g2_nand2_1 _27187_ (.Y(_07961_),
    .A(net473),
    .B(_07960_));
 sg13g2_or2_1 _27188_ (.X(_07962_),
    .B(_07953_),
    .A(net143));
 sg13g2_o21ai_1 _27189_ (.B1(_07962_),
    .Y(_07963_),
    .A1(net117),
    .A2(_07960_));
 sg13g2_a22oi_1 _27190_ (.Y(_07964_),
    .B1(_07963_),
    .B2(net1037),
    .A2(_07961_),
    .A1(_07954_));
 sg13g2_nor2_1 _27191_ (.A(_07866_),
    .B(_07964_),
    .Y(_07965_));
 sg13g2_a21oi_1 _27192_ (.A1(net484),
    .A2(_07951_),
    .Y(_07966_),
    .B1(_07965_));
 sg13g2_nor2_1 _27193_ (.A(_07858_),
    .B(_07966_),
    .Y(_07967_));
 sg13g2_a21oi_1 _27194_ (.A1(\cpu.spi.r_count[4] ),
    .A2(net59),
    .Y(_07968_),
    .B1(_07967_));
 sg13g2_nor2_1 _27195_ (.A(net558),
    .B(_07968_),
    .Y(_02577_));
 sg13g2_nand2b_1 _27196_ (.Y(_07969_),
    .B(net655),
    .A_N(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_o21ai_1 _27197_ (.B1(_07969_),
    .Y(_07970_),
    .A1(net656),
    .A2(_05652_));
 sg13g2_mux2_1 _27198_ (.A0(\cpu.spi.r_clk_count[0][5] ),
    .A1(\cpu.spi.r_clk_count[1][5] ),
    .S(net734),
    .X(_07971_));
 sg13g2_nor2_1 _27199_ (.A(net735),
    .B(_07971_),
    .Y(_07972_));
 sg13g2_a21oi_1 _27200_ (.A1(net657),
    .A2(_07970_),
    .Y(_07973_),
    .B1(_07972_));
 sg13g2_nor2_1 _27201_ (.A(net855),
    .B(_05652_),
    .Y(_07974_));
 sg13g2_a21oi_1 _27202_ (.A1(net856),
    .A2(_00133_),
    .Y(_07975_),
    .B1(_07974_));
 sg13g2_nand2_1 _27203_ (.Y(_07976_),
    .A(net1001),
    .B(_00132_));
 sg13g2_o21ai_1 _27204_ (.B1(_07976_),
    .Y(_07977_),
    .A1(net855),
    .A2(_05651_));
 sg13g2_nor2_1 _27205_ (.A(net1002),
    .B(_07977_),
    .Y(_07978_));
 sg13g2_a21oi_1 _27206_ (.A1(net1002),
    .A2(_07975_),
    .Y(_07979_),
    .B1(_07978_));
 sg13g2_nand2_1 _27207_ (.Y(_07980_),
    .A(net473),
    .B(_07979_));
 sg13g2_xnor2_1 _27208_ (.Y(_07981_),
    .A(\cpu.spi.r_count[5] ),
    .B(_09189_));
 sg13g2_nor2_1 _27209_ (.A(net642),
    .B(_07981_),
    .Y(_07982_));
 sg13g2_or2_1 _27210_ (.X(_07983_),
    .B(_07981_),
    .A(_09263_));
 sg13g2_o21ai_1 _27211_ (.B1(_07983_),
    .Y(_07984_),
    .A1(net117),
    .A2(_07979_));
 sg13g2_a22oi_1 _27212_ (.Y(_07985_),
    .B1(_07984_),
    .B2(net1037),
    .A2(_07982_),
    .A1(_07980_));
 sg13g2_nor2_1 _27213_ (.A(_07866_),
    .B(_07985_),
    .Y(_07986_));
 sg13g2_a21oi_1 _27214_ (.A1(net484),
    .A2(_07973_),
    .Y(_07987_),
    .B1(_07986_));
 sg13g2_nor2_1 _27215_ (.A(_07858_),
    .B(_07987_),
    .Y(_07988_));
 sg13g2_a21oi_1 _27216_ (.A1(\cpu.spi.r_count[5] ),
    .A2(net59),
    .Y(_07989_),
    .B1(_07988_));
 sg13g2_nor2_1 _27217_ (.A(net558),
    .B(_07989_),
    .Y(_02578_));
 sg13g2_nand2b_1 _27218_ (.Y(_07990_),
    .B(_11943_),
    .A_N(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_o21ai_1 _27219_ (.B1(_07990_),
    .Y(_07991_),
    .A1(_11937_),
    .A2(_05741_));
 sg13g2_mux2_1 _27220_ (.A0(\cpu.spi.r_clk_count[0][6] ),
    .A1(\cpu.spi.r_clk_count[1][6] ),
    .S(net734),
    .X(_07992_));
 sg13g2_nor2_1 _27221_ (.A(net735),
    .B(_07992_),
    .Y(_07993_));
 sg13g2_a21oi_1 _27222_ (.A1(_11936_),
    .A2(_07991_),
    .Y(_07994_),
    .B1(_07993_));
 sg13g2_nor2_1 _27223_ (.A(_11955_),
    .B(_05741_),
    .Y(_07995_));
 sg13g2_a21oi_1 _27224_ (.A1(_11954_),
    .A2(_00145_),
    .Y(_07996_),
    .B1(_07995_));
 sg13g2_nand2_1 _27225_ (.Y(_07997_),
    .A(net1001),
    .B(_00144_));
 sg13g2_o21ai_1 _27226_ (.B1(_07997_),
    .Y(_07998_),
    .A1(_11955_),
    .A2(_05740_));
 sg13g2_nor2_1 _27227_ (.A(_11948_),
    .B(_07998_),
    .Y(_07999_));
 sg13g2_a21oi_1 _27228_ (.A1(_11948_),
    .A2(_07996_),
    .Y(_08000_),
    .B1(_07999_));
 sg13g2_nand2_1 _27229_ (.Y(_08001_),
    .A(net473),
    .B(_08000_));
 sg13g2_xnor2_1 _27230_ (.Y(_08002_),
    .A(\cpu.spi.r_count[6] ),
    .B(_09190_));
 sg13g2_nor2_1 _27231_ (.A(net642),
    .B(_08002_),
    .Y(_08003_));
 sg13g2_or2_1 _27232_ (.X(_08004_),
    .B(_08002_),
    .A(_09263_));
 sg13g2_o21ai_1 _27233_ (.B1(_08004_),
    .Y(_08005_),
    .A1(net117),
    .A2(_08000_));
 sg13g2_a22oi_1 _27234_ (.Y(_08006_),
    .B1(_08005_),
    .B2(net1037),
    .A2(_08003_),
    .A1(_08001_));
 sg13g2_nor2_1 _27235_ (.A(_07866_),
    .B(_08006_),
    .Y(_08007_));
 sg13g2_a21oi_1 _27236_ (.A1(net484),
    .A2(_07994_),
    .Y(_08008_),
    .B1(_08007_));
 sg13g2_nor2_1 _27237_ (.A(_07858_),
    .B(_08008_),
    .Y(_08009_));
 sg13g2_a21oi_1 _27238_ (.A1(\cpu.spi.r_count[6] ),
    .A2(net59),
    .Y(_08010_),
    .B1(_08009_));
 sg13g2_nor2_1 _27239_ (.A(_07925_),
    .B(_08010_),
    .Y(_02579_));
 sg13g2_nor2_1 _27240_ (.A(net732),
    .B(_05079_),
    .Y(_08011_));
 sg13g2_a21oi_1 _27241_ (.A1(net732),
    .A2(_00157_),
    .Y(_08012_),
    .B1(_08011_));
 sg13g2_nand2_1 _27242_ (.Y(_08013_),
    .A(net856),
    .B(_00156_));
 sg13g2_o21ai_1 _27243_ (.B1(_08013_),
    .Y(_08014_),
    .A1(net732),
    .A2(_05078_));
 sg13g2_nor2_1 _27244_ (.A(_11949_),
    .B(_08014_),
    .Y(_08015_));
 sg13g2_a21oi_1 _27245_ (.A1(_11949_),
    .A2(_08012_),
    .Y(_08016_),
    .B1(_08015_));
 sg13g2_nand2_1 _27246_ (.Y(_08017_),
    .A(net143),
    .B(_08016_));
 sg13g2_nand2b_1 _27247_ (.Y(_08018_),
    .B(_09183_),
    .A_N(_09191_));
 sg13g2_nand3_1 _27248_ (.B(_09194_),
    .C(_08018_),
    .A(net117),
    .Y(_08019_));
 sg13g2_nand4_1 _27249_ (.B(_07865_),
    .C(_08017_),
    .A(net1037),
    .Y(_08020_),
    .D(_08019_));
 sg13g2_and2_1 _27250_ (.A(_11927_),
    .B(\cpu.spi.r_clk_count[1][7] ),
    .X(_08021_));
 sg13g2_a21oi_1 _27251_ (.A1(net733),
    .A2(\cpu.spi.r_clk_count[0][7] ),
    .Y(_08022_),
    .B1(_08021_));
 sg13g2_mux2_1 _27252_ (.A0(_05079_),
    .A1(\cpu.spi.r_clk_count[0][7] ),
    .S(_11927_),
    .X(_08023_));
 sg13g2_nand2_1 _27253_ (.Y(_08024_),
    .A(_11926_),
    .B(_08023_));
 sg13g2_o21ai_1 _27254_ (.B1(_08024_),
    .Y(_08025_),
    .A1(_11936_),
    .A2(_08022_));
 sg13g2_o21ai_1 _27255_ (.B1(_08018_),
    .Y(_08026_),
    .A1(net419),
    .A2(_08016_));
 sg13g2_inv_1 _27256_ (.Y(_08027_),
    .A(net642));
 sg13g2_a22oi_1 _27257_ (.Y(_08028_),
    .B1(_08026_),
    .B2(_08027_),
    .A2(_08025_),
    .A1(_07867_));
 sg13g2_a21oi_1 _27258_ (.A1(_08020_),
    .A2(_08028_),
    .Y(_08029_),
    .B1(_07858_));
 sg13g2_a21oi_1 _27259_ (.A1(_09183_),
    .A2(_07859_),
    .Y(_08030_),
    .B1(_08029_));
 sg13g2_nor2_1 _27260_ (.A(net558),
    .B(_08030_),
    .Y(_02580_));
 sg13g2_inv_1 _27261_ (.Y(_08031_),
    .A(_09283_));
 sg13g2_nand2_1 _27262_ (.Y(_08032_),
    .A(_08031_),
    .B(_09196_));
 sg13g2_nor3_1 _27263_ (.A(_09347_),
    .B(_09335_),
    .C(_08032_),
    .Y(_08033_));
 sg13g2_a21oi_1 _27264_ (.A1(net857),
    .A2(_11963_),
    .Y(_08034_),
    .B1(net419));
 sg13g2_nor3_1 _27265_ (.A(_00276_),
    .B(_08033_),
    .C(_08034_),
    .Y(_08035_));
 sg13g2_inv_1 _27266_ (.Y(_08036_),
    .A(_00276_));
 sg13g2_a21oi_1 _27267_ (.A1(net418),
    .A2(_08032_),
    .Y(_08037_),
    .B1(_08036_));
 sg13g2_a21oi_1 _27268_ (.A1(_09346_),
    .A2(_09282_),
    .Y(_08038_),
    .B1(_06948_));
 sg13g2_nor3_1 _27269_ (.A(_08035_),
    .B(_08037_),
    .C(_08038_),
    .Y(_08039_));
 sg13g2_a21oi_1 _27270_ (.A1(_08032_),
    .A2(_08039_),
    .Y(_08040_),
    .B1(_09296_));
 sg13g2_nand2_1 _27271_ (.Y(_08041_),
    .A(_11962_),
    .B(_08039_));
 sg13g2_buf_1 _27272_ (.A(\cpu.gpio.genblk1[3].srcs_o[6] ),
    .X(_08042_));
 sg13g2_o21ai_1 _27273_ (.B1(_08042_),
    .Y(_08043_),
    .A1(_11963_),
    .A2(_08041_));
 sg13g2_nand2_1 _27274_ (.Y(_02581_),
    .A(_08040_),
    .B(_08043_));
 sg13g2_buf_1 _27275_ (.A(\cpu.gpio.genblk1[3].srcs_o[7] ),
    .X(_08044_));
 sg13g2_o21ai_1 _27276_ (.B1(_08044_),
    .Y(_08045_),
    .A1(_11951_),
    .A2(_08041_));
 sg13g2_nand2_1 _27277_ (.Y(_02582_),
    .A(_08040_),
    .B(_08045_));
 sg13g2_buf_1 _27278_ (.A(\cpu.gpio.genblk1[3].srcs_o[8] ),
    .X(_08046_));
 sg13g2_nand2_1 _27279_ (.Y(_08047_),
    .A(_11965_),
    .B(_08039_));
 sg13g2_nand2_1 _27280_ (.Y(_08048_),
    .A(_08046_),
    .B(_08047_));
 sg13g2_nand2_1 _27281_ (.Y(_02583_),
    .A(_08040_),
    .B(_08048_));
 sg13g2_nor3_1 _27282_ (.A(_06948_),
    .B(_09263_),
    .C(_09282_),
    .Y(_08049_));
 sg13g2_o21ai_1 _27283_ (.B1(_09290_),
    .Y(_08050_),
    .A1(_09285_),
    .A2(_08049_));
 sg13g2_o21ai_1 _27284_ (.B1(_08050_),
    .Y(_08051_),
    .A1(_11988_),
    .A2(_09330_));
 sg13g2_o21ai_1 _27285_ (.B1(_09252_),
    .Y(_08052_),
    .A1(_06944_),
    .A2(_08051_));
 sg13g2_nand3_1 _27286_ (.B(_09330_),
    .C(_08050_),
    .A(_09332_),
    .Y(_08053_));
 sg13g2_a21oi_1 _27287_ (.A1(_08052_),
    .A2(_08053_),
    .Y(_02592_),
    .B1(net559));
 sg13g2_nand2_1 _27288_ (.Y(_08054_),
    .A(_09344_),
    .B(_09289_));
 sg13g2_nor4_1 _27289_ (.A(net657),
    .B(net595),
    .C(_04943_),
    .D(_08054_),
    .Y(_08055_));
 sg13g2_buf_1 _27290_ (.A(_08055_),
    .X(_08056_));
 sg13g2_nand2b_1 _27291_ (.Y(_08057_),
    .B(\cpu.spi.r_mode[0][0] ),
    .A_N(_08056_));
 sg13g2_nand2_1 _27292_ (.Y(_08058_),
    .A(net799),
    .B(_08056_));
 sg13g2_a21oi_1 _27293_ (.A1(_08057_),
    .A2(_08058_),
    .Y(_02593_),
    .B1(net559));
 sg13g2_nand2b_1 _27294_ (.Y(_08059_),
    .B(_11939_),
    .A_N(_08056_));
 sg13g2_nand2_1 _27295_ (.Y(_08060_),
    .A(net1027),
    .B(_08056_));
 sg13g2_a21oi_1 _27296_ (.A1(_08059_),
    .A2(_08060_),
    .Y(_02594_),
    .B1(net559));
 sg13g2_nor4_1 _27297_ (.A(net657),
    .B(net733),
    .C(_04943_),
    .D(_08054_),
    .Y(_08061_));
 sg13g2_buf_1 _27298_ (.A(_08061_),
    .X(_08062_));
 sg13g2_nand2b_1 _27299_ (.Y(_08063_),
    .B(\cpu.spi.r_mode[1][0] ),
    .A_N(_08062_));
 sg13g2_nand2_1 _27300_ (.Y(_08064_),
    .A(net799),
    .B(_08062_));
 sg13g2_a21oi_1 _27301_ (.A1(_08063_),
    .A2(_08064_),
    .Y(_02595_),
    .B1(net559));
 sg13g2_nand2b_1 _27302_ (.Y(_08065_),
    .B(_11942_),
    .A_N(_08062_));
 sg13g2_nand2_1 _27303_ (.Y(_08066_),
    .A(_10070_),
    .B(_08062_));
 sg13g2_a21oi_1 _27304_ (.A1(_08065_),
    .A2(_08066_),
    .Y(_02596_),
    .B1(_07837_));
 sg13g2_nand3_1 _27305_ (.B(_09289_),
    .C(_07840_),
    .A(_09344_),
    .Y(_08067_));
 sg13g2_buf_1 _27306_ (.A(_08067_),
    .X(_08068_));
 sg13g2_mux2_1 _27307_ (.A0(net1029),
    .A1(\cpu.spi.r_mode[2][0] ),
    .S(_08068_),
    .X(_08069_));
 sg13g2_and2_1 _27308_ (.A(net659),
    .B(_08069_),
    .X(_02597_));
 sg13g2_nand2_1 _27309_ (.Y(_08070_),
    .A(_11938_),
    .B(_08068_));
 sg13g2_o21ai_1 _27310_ (.B1(_08070_),
    .Y(_08071_),
    .A1(net887),
    .A2(_08068_));
 sg13g2_and2_1 _27311_ (.A(net659),
    .B(_08071_),
    .X(_02598_));
 sg13g2_a21oi_1 _27312_ (.A1(_08031_),
    .A2(_07793_),
    .Y(_08072_),
    .B1(_08051_));
 sg13g2_nor2_1 _27313_ (.A(\cpu.spi.r_ready ),
    .B(net418),
    .Y(_08073_));
 sg13g2_nor4_1 _27314_ (.A(_09283_),
    .B(_09265_),
    .C(_07793_),
    .D(_08051_),
    .Y(_08074_));
 sg13g2_o21ai_1 _27315_ (.B1(_11988_),
    .Y(_08075_),
    .A1(_08073_),
    .A2(_08074_));
 sg13g2_o21ai_1 _27316_ (.B1(_08075_),
    .Y(_08076_),
    .A1(\cpu.spi.r_ready ),
    .A2(_08072_));
 sg13g2_nand2_1 _27317_ (.Y(_02607_),
    .A(net675),
    .B(_08076_));
 sg13g2_nand2_1 _27318_ (.Y(_08077_),
    .A(_09338_),
    .B(_07795_));
 sg13g2_nand2_1 _27319_ (.Y(_08078_),
    .A(\cpu.spi.r_searching ),
    .B(_08077_));
 sg13g2_nand2_1 _27320_ (.Y(_08079_),
    .A(net780),
    .B(_09289_));
 sg13g2_nand4_1 _27321_ (.B(_09338_),
    .C(_07795_),
    .A(net897),
    .Y(_08080_),
    .D(_08079_));
 sg13g2_a21oi_1 _27322_ (.A1(_08078_),
    .A2(_08080_),
    .Y(_02608_),
    .B1(net559));
 sg13g2_nand2b_1 _27323_ (.Y(_08081_),
    .B(\cpu.spi.r_src[0] ),
    .A_N(_08056_));
 sg13g2_nand2_1 _27324_ (.Y(_08082_),
    .A(net1026),
    .B(_08056_));
 sg13g2_a21oi_1 _27325_ (.A1(_08081_),
    .A2(_08082_),
    .Y(_02611_),
    .B1(_07837_));
 sg13g2_nand2b_1 _27326_ (.Y(_08083_),
    .B(\cpu.spi.r_src[1] ),
    .A_N(_08062_));
 sg13g2_nand2_1 _27327_ (.Y(_08084_),
    .A(net1026),
    .B(_08062_));
 sg13g2_buf_1 _27328_ (.A(_09351_),
    .X(_08085_));
 sg13g2_a21oi_1 _27329_ (.A1(_08083_),
    .A2(_08084_),
    .Y(_02612_),
    .B1(_08085_));
 sg13g2_mux2_1 _27330_ (.A0(net1020),
    .A1(_11932_),
    .S(_08068_),
    .X(_08086_));
 sg13g2_and2_1 _27331_ (.A(net659),
    .B(_08086_),
    .X(_02613_));
 sg13g2_and2_1 _27332_ (.A(net388),
    .B(_07042_),
    .X(_08087_));
 sg13g2_buf_2 _27333_ (.A(_08087_),
    .X(_08088_));
 sg13g2_nand2_1 _27334_ (.Y(_08089_),
    .A(net850),
    .B(_08088_));
 sg13g2_nand2_1 _27335_ (.Y(_08090_),
    .A(net388),
    .B(_07042_));
 sg13g2_buf_2 _27336_ (.A(_08090_),
    .X(_08091_));
 sg13g2_nand2_1 _27337_ (.Y(_08092_),
    .A(\cpu.uart.r_div_value[0] ),
    .B(_08091_));
 sg13g2_nand3_1 _27338_ (.B(_08089_),
    .C(_08092_),
    .A(net645),
    .Y(_02630_));
 sg13g2_buf_1 _27339_ (.A(_07042_),
    .X(_08093_));
 sg13g2_nand3_1 _27340_ (.B(net389),
    .C(net108),
    .A(net1026),
    .Y(_08094_));
 sg13g2_nand2_1 _27341_ (.Y(_08095_),
    .A(net389),
    .B(net108));
 sg13g2_nand2_1 _27342_ (.Y(_08096_),
    .A(_09952_),
    .B(_08095_));
 sg13g2_a21oi_1 _27343_ (.A1(_08094_),
    .A2(_08096_),
    .Y(_02631_),
    .B1(net557));
 sg13g2_nand3_1 _27344_ (.B(net389),
    .C(net108),
    .A(net1025),
    .Y(_08097_));
 sg13g2_nand2_1 _27345_ (.Y(_08098_),
    .A(\cpu.uart.r_div_value[11] ),
    .B(_08095_));
 sg13g2_a21oi_1 _27346_ (.A1(_08097_),
    .A2(_08098_),
    .Y(_02632_),
    .B1(net557));
 sg13g2_nand2_1 _27347_ (.Y(_08099_),
    .A(net939),
    .B(_08088_));
 sg13g2_nand2_1 _27348_ (.Y(_08100_),
    .A(\cpu.uart.r_div_value[1] ),
    .B(_08091_));
 sg13g2_a21oi_1 _27349_ (.A1(_08099_),
    .A2(_08100_),
    .Y(_02633_),
    .B1(net557));
 sg13g2_nand2_1 _27350_ (.Y(_08101_),
    .A(net1026),
    .B(_08088_));
 sg13g2_nand2_1 _27351_ (.Y(_08102_),
    .A(\cpu.uart.r_div_value[2] ),
    .B(_08091_));
 sg13g2_a21oi_1 _27352_ (.A1(_08101_),
    .A2(_08102_),
    .Y(_02634_),
    .B1(_08085_));
 sg13g2_nand2_1 _27353_ (.Y(_08103_),
    .A(net1025),
    .B(_08088_));
 sg13g2_nand2_1 _27354_ (.Y(_08104_),
    .A(\cpu.uart.r_div_value[3] ),
    .B(_08091_));
 sg13g2_a21oi_1 _27355_ (.A1(_08103_),
    .A2(_08104_),
    .Y(_02635_),
    .B1(net557));
 sg13g2_nand2_1 _27356_ (.Y(_08105_),
    .A(net1024),
    .B(_08088_));
 sg13g2_nand2_1 _27357_ (.Y(_08106_),
    .A(\cpu.uart.r_div_value[4] ),
    .B(_08091_));
 sg13g2_a21oi_1 _27358_ (.A1(_08105_),
    .A2(_08106_),
    .Y(_02636_),
    .B1(net557));
 sg13g2_nand2_1 _27359_ (.Y(_08107_),
    .A(net1023),
    .B(_08088_));
 sg13g2_nand2_1 _27360_ (.Y(_08108_),
    .A(\cpu.uart.r_div_value[5] ),
    .B(_08091_));
 sg13g2_a21oi_1 _27361_ (.A1(_08107_),
    .A2(_08108_),
    .Y(_02637_),
    .B1(net557));
 sg13g2_nand2_1 _27362_ (.Y(_08109_),
    .A(net1022),
    .B(_08088_));
 sg13g2_nand2_1 _27363_ (.Y(_08110_),
    .A(\cpu.uart.r_div_value[6] ),
    .B(_08091_));
 sg13g2_a21oi_1 _27364_ (.A1(_08109_),
    .A2(_08110_),
    .Y(_02638_),
    .B1(net557));
 sg13g2_nand2_1 _27365_ (.Y(_08111_),
    .A(net1021),
    .B(_08088_));
 sg13g2_nand2_1 _27366_ (.Y(_08112_),
    .A(\cpu.uart.r_div_value[7] ),
    .B(_08091_));
 sg13g2_a21oi_1 _27367_ (.A1(_08111_),
    .A2(_08112_),
    .Y(_02639_),
    .B1(net557));
 sg13g2_nand3_1 _27368_ (.B(net389),
    .C(_08093_),
    .A(net799),
    .Y(_08113_));
 sg13g2_nand2_1 _27369_ (.Y(_08114_),
    .A(\cpu.uart.r_div_value[8] ),
    .B(_08095_));
 sg13g2_a21oi_1 _27370_ (.A1(_08113_),
    .A2(_08114_),
    .Y(_02640_),
    .B1(net629));
 sg13g2_nand3_1 _27371_ (.B(net389),
    .C(net108),
    .A(net1027),
    .Y(_08115_));
 sg13g2_nand2_1 _27372_ (.Y(_08116_),
    .A(\cpu.uart.r_div_value[9] ),
    .B(_08095_));
 sg13g2_a21oi_1 _27373_ (.A1(_08115_),
    .A2(_08116_),
    .Y(_02641_),
    .B1(net629));
 sg13g2_nand3_1 _27374_ (.B(net397),
    .C(net108),
    .A(net1027),
    .Y(_08117_));
 sg13g2_nor2_1 _27375_ (.A(net1028),
    .B(net648),
    .Y(_08118_));
 sg13g2_nand4_1 _27376_ (.B(_05038_),
    .C(_07040_),
    .A(net651),
    .Y(_08119_),
    .D(_08118_));
 sg13g2_or2_1 _27377_ (.X(_08120_),
    .B(_08119_),
    .A(_09275_));
 sg13g2_nand4_1 _27378_ (.B(net764),
    .C(_08117_),
    .A(_09249_),
    .Y(_08121_),
    .D(_08120_));
 sg13g2_nand2b_1 _27379_ (.Y(_02665_),
    .B(_08121_),
    .A_N(net178));
 sg13g2_nand3_1 _27380_ (.B(net440),
    .C(net108),
    .A(net1027),
    .Y(_08122_));
 sg13g2_nand2_1 _27381_ (.Y(_08123_),
    .A(net440),
    .B(net108));
 sg13g2_nand2_1 _27382_ (.Y(_08124_),
    .A(\cpu.uart.r_r_invert ),
    .B(_08123_));
 sg13g2_a21oi_1 _27383_ (.A1(_08122_),
    .A2(_08124_),
    .Y(_02666_),
    .B1(net629));
 sg13g2_a21oi_1 _27384_ (.A1(_07027_),
    .A2(_09930_),
    .Y(_08125_),
    .B1(net1080));
 sg13g2_a21oi_1 _27385_ (.A1(_07028_),
    .A2(_09930_),
    .Y(_08126_),
    .B1(_07098_));
 sg13g2_a221oi_1 _27386_ (.B2(_08125_),
    .C1(_08126_),
    .B1(_07026_),
    .A1(net932),
    .Y(_08127_),
    .A2(net937));
 sg13g2_a21oi_1 _27387_ (.A1(_07020_),
    .A2(_08127_),
    .Y(_08128_),
    .B1(_07095_));
 sg13g2_buf_2 _27388_ (.A(_08128_),
    .X(_08129_));
 sg13g2_o21ai_1 _27389_ (.B1(_08129_),
    .Y(_08130_),
    .A1(net932),
    .A2(_07098_));
 sg13g2_xnor2_1 _27390_ (.Y(_08131_),
    .A(_07028_),
    .B(_08130_));
 sg13g2_nor2_1 _27391_ (.A(net558),
    .B(_08131_),
    .Y(_02669_));
 sg13g2_o21ai_1 _27392_ (.B1(_08129_),
    .Y(_08132_),
    .A1(_07027_),
    .A2(net937));
 sg13g2_nand2_1 _27393_ (.Y(_08133_),
    .A(_07024_),
    .B(_08132_));
 sg13g2_nand2b_1 _27394_ (.Y(_08134_),
    .B(net932),
    .A_N(net937));
 sg13g2_o21ai_1 _27395_ (.B1(_08134_),
    .Y(_08135_),
    .A1(net932),
    .A2(_07097_));
 sg13g2_nand3_1 _27396_ (.B(_08129_),
    .C(_08135_),
    .A(_07096_),
    .Y(_08136_));
 sg13g2_a21oi_1 _27397_ (.A1(_08133_),
    .A2(_08136_),
    .Y(_02670_),
    .B1(net629));
 sg13g2_nand2_1 _27398_ (.Y(_08137_),
    .A(_07027_),
    .B(net1079));
 sg13g2_nor3_1 _27399_ (.A(net932),
    .B(net937),
    .C(_08137_),
    .Y(_08138_));
 sg13g2_o21ai_1 _27400_ (.B1(_08129_),
    .Y(_08139_),
    .A1(net937),
    .A2(_07106_));
 sg13g2_a22oi_1 _27401_ (.Y(_08140_),
    .B1(_08139_),
    .B2(net932),
    .A2(_08138_),
    .A1(_08129_));
 sg13g2_nor2_1 _27402_ (.A(net558),
    .B(_08140_),
    .Y(_02671_));
 sg13g2_a21oi_1 _27403_ (.A1(_07106_),
    .A2(_08129_),
    .Y(_08141_),
    .B1(net937));
 sg13g2_nor2b_1 _27404_ (.A(_07092_),
    .B_N(net1079),
    .Y(_08142_));
 sg13g2_a21oi_1 _27405_ (.A1(_08129_),
    .A2(_08142_),
    .Y(_08143_),
    .B1(_06734_));
 sg13g2_nor2b_1 _27406_ (.A(_08141_),
    .B_N(_08143_),
    .Y(_02672_));
 sg13g2_or2_1 _27407_ (.X(_08144_),
    .B(_07120_),
    .A(_07039_));
 sg13g2_a21oi_1 _27408_ (.A1(_10047_),
    .A2(net397),
    .Y(_08145_),
    .B1(net391));
 sg13g2_o21ai_1 _27409_ (.B1(_04950_),
    .Y(_08146_),
    .A1(_00221_),
    .A2(net583));
 sg13g2_nand3_1 _27410_ (.B(_07144_),
    .C(_08146_),
    .A(net895),
    .Y(_08147_));
 sg13g2_o21ai_1 _27411_ (.B1(_08147_),
    .Y(_08148_),
    .A1(_07120_),
    .A2(_08145_));
 sg13g2_nand3_1 _27412_ (.B(_08144_),
    .C(_08148_),
    .A(_08093_),
    .Y(_08149_));
 sg13g2_nor2_1 _27413_ (.A(_07059_),
    .B(_08144_),
    .Y(_08150_));
 sg13g2_a21oi_1 _27414_ (.A1(_09248_),
    .A2(_08149_),
    .Y(_08151_),
    .B1(_08150_));
 sg13g2_nor2_1 _27415_ (.A(_07925_),
    .B(_08151_),
    .Y(_02674_));
 sg13g2_nand3_1 _27416_ (.B(net440),
    .C(net108),
    .A(net799),
    .Y(_08152_));
 sg13g2_nand2_1 _27417_ (.Y(_08153_),
    .A(\cpu.uart.r_x_invert ),
    .B(_08123_));
 sg13g2_a21oi_1 _27418_ (.A1(_08152_),
    .A2(_08153_),
    .Y(_02675_),
    .B1(net629));
 sg13g2_and2_1 _27419_ (.A(net936),
    .B(_07038_),
    .X(_08154_));
 sg13g2_buf_1 _27420_ (.A(_08154_),
    .X(_08155_));
 sg13g2_nand2_1 _27421_ (.Y(_08156_),
    .A(_07043_),
    .B(_08155_));
 sg13g2_nand2_1 _27422_ (.Y(_08157_),
    .A(_07046_),
    .B(_07117_));
 sg13g2_o21ai_1 _27423_ (.B1(_08157_),
    .Y(_08158_),
    .A1(net933),
    .A2(_08156_));
 sg13g2_a221oi_1 _27424_ (.B2(_07134_),
    .C1(_07138_),
    .B1(_08158_),
    .A1(_07043_),
    .Y(_08159_),
    .A2(_07144_));
 sg13g2_buf_2 _27425_ (.A(_08159_),
    .X(_08160_));
 sg13g2_nor2b_1 _27426_ (.A(_07116_),
    .B_N(_08160_),
    .Y(_08161_));
 sg13g2_nand2b_1 _27427_ (.Y(_08162_),
    .B(_07128_),
    .A_N(_07059_));
 sg13g2_nand3_1 _27428_ (.B(_08161_),
    .C(_08162_),
    .A(net935),
    .Y(_08163_));
 sg13g2_o21ai_1 _27429_ (.B1(_08163_),
    .Y(_08164_),
    .A1(net935),
    .A2(_08160_));
 sg13g2_nor2_1 _27430_ (.A(net558),
    .B(_08164_),
    .Y(_02678_));
 sg13g2_o21ai_1 _27431_ (.B1(_08160_),
    .Y(_08165_),
    .A1(net935),
    .A2(_07116_));
 sg13g2_nor2b_1 _27432_ (.A(net936),
    .B_N(net935),
    .Y(_08166_));
 sg13g2_a22oi_1 _27433_ (.Y(_08167_),
    .B1(_08166_),
    .B2(_08161_),
    .A2(_08165_),
    .A1(net936));
 sg13g2_nor2_1 _27434_ (.A(net558),
    .B(_08167_),
    .Y(_02679_));
 sg13g2_a21oi_1 _27435_ (.A1(_08155_),
    .A2(_08160_),
    .Y(_08168_),
    .B1(net933));
 sg13g2_nand2_1 _27436_ (.Y(_08169_),
    .A(net933),
    .B(_08155_));
 sg13g2_a22oi_1 _27437_ (.Y(_08170_),
    .B1(_08169_),
    .B2(_07126_),
    .A2(_07128_),
    .A1(_07059_));
 sg13g2_a21oi_1 _27438_ (.A1(_08160_),
    .A2(_08170_),
    .Y(_08171_),
    .B1(_06734_));
 sg13g2_nor2b_1 _27439_ (.A(_08168_),
    .B_N(_08171_),
    .Y(_02680_));
 sg13g2_o21ai_1 _27440_ (.B1(_08160_),
    .Y(_08172_),
    .A1(net933),
    .A2(_08155_));
 sg13g2_nand2_1 _27441_ (.Y(_08173_),
    .A(_07059_),
    .B(_07128_));
 sg13g2_o21ai_1 _27442_ (.B1(_08173_),
    .Y(_08174_),
    .A1(net934),
    .A2(_08169_));
 sg13g2_a22oi_1 _27443_ (.Y(_08175_),
    .B1(_08174_),
    .B2(_08160_),
    .A2(_08172_),
    .A1(net934));
 sg13g2_nor2_1 _27444_ (.A(_09352_),
    .B(_08175_),
    .Y(_02681_));
 sg13g2_nand2b_1 _27445_ (.Y(\cpu.ex.genblk3.c_supmode ),
    .B(_07321_),
    .A_N(_07318_));
 sg13g2_nand2_1 _27446_ (.Y(_08176_),
    .A(_09876_),
    .B(_07761_));
 sg13g2_nor4_1 _27447_ (.A(_09910_),
    .B(_09874_),
    .C(_06787_),
    .D(_08176_),
    .Y(_08177_));
 sg13g2_a22oi_1 _27448_ (.Y(_08178_),
    .B1(net142),
    .B2(_08177_),
    .A2(_09848_),
    .A1(net1118));
 sg13g2_inv_1 _27449_ (.Y(\cpu.qspi.c_rstrobe_d ),
    .A(_08178_));
 sg13g2_nor2_1 _27450_ (.A(_09848_),
    .B(_08176_),
    .Y(_08179_));
 sg13g2_a22oi_1 _27451_ (.Y(_08180_),
    .B1(_07742_),
    .B2(_08179_),
    .A2(_09848_),
    .A1(_09843_));
 sg13g2_nor2_1 _27452_ (.A(net798),
    .B(_08180_),
    .Y(\cpu.qspi.c_wstrobe_d ));
 sg13g2_nor2_1 _27453_ (.A(_08462_),
    .B(_08180_),
    .Y(\cpu.qspi.c_wstrobe_i ));
 sg13g2_mux4_1 _27454_ (.S0(_04925_),
    .A0(_09220_),
    .A1(_09226_),
    .A2(_09215_),
    .A3(_09230_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08181_));
 sg13g2_mux4_1 _27455_ (.S0(_04925_),
    .A0(_09234_),
    .A1(_09236_),
    .A2(_09222_),
    .A3(_09217_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08182_));
 sg13g2_mux2_1 _27456_ (.A0(_08181_),
    .A1(_08182_),
    .S(\cpu.gpio.r_uart_rx_src[2] ),
    .X(\cpu.gpio.uart_rx ));
 sg13g2_mux4_1 _27457_ (.S0(_04937_),
    .A0(net1099),
    .A1(net1100),
    .A2(net1076),
    .A3(net1075),
    .S1(_05361_),
    .X(_08183_));
 sg13g2_mux4_1 _27458_ (.S0(_04937_),
    .A0(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A1(net1078),
    .A2(net1097),
    .A3(net1098),
    .S1(_05361_),
    .X(_08184_));
 sg13g2_nor2b_1 _27459_ (.A(_05448_),
    .B_N(_08184_),
    .Y(_08185_));
 sg13g2_a21oi_1 _27460_ (.A1(_05448_),
    .A2(_08183_),
    .Y(_08186_),
    .B1(_08185_));
 sg13g2_nand2b_1 _27461_ (.Y(_08187_),
    .B(net1074),
    .A_N(_04937_));
 sg13g2_nand3_1 _27462_ (.B(_05361_),
    .C(net1077),
    .A(_04937_),
    .Y(_08188_));
 sg13g2_o21ai_1 _27463_ (.B1(_08188_),
    .Y(_08189_),
    .A1(_05361_),
    .A2(_08187_));
 sg13g2_nand3_1 _27464_ (.B(_00187_),
    .C(_08189_),
    .A(_05522_),
    .Y(_08190_));
 sg13g2_o21ai_1 _27465_ (.B1(_08190_),
    .Y(net15),
    .A1(_05522_),
    .A2(_08186_));
 sg13g2_mux4_1 _27466_ (.S0(_05576_),
    .A0(net1099),
    .A1(net1100),
    .A2(net1076),
    .A3(net1075),
    .S1(_05646_),
    .X(_08191_));
 sg13g2_mux4_1 _27467_ (.S0(_05576_),
    .A0(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .A1(net1078),
    .A2(net1097),
    .A3(net1098),
    .S1(_05646_),
    .X(_08192_));
 sg13g2_nor2b_1 _27468_ (.A(_05720_),
    .B_N(_08192_),
    .Y(_08193_));
 sg13g2_a21oi_1 _27469_ (.A1(_05720_),
    .A2(_08191_),
    .Y(_08194_),
    .B1(_08193_));
 sg13g2_nand2b_1 _27470_ (.Y(_08195_),
    .B(net1074),
    .A_N(_05576_));
 sg13g2_nand3_1 _27471_ (.B(_05646_),
    .C(net1077),
    .A(_05576_),
    .Y(_08196_));
 sg13g2_o21ai_1 _27472_ (.B1(_08196_),
    .Y(_08197_),
    .A1(_05646_),
    .A2(_08195_));
 sg13g2_nand3_1 _27473_ (.B(_00186_),
    .C(_08197_),
    .A(_05094_),
    .Y(_08198_));
 sg13g2_o21ai_1 _27474_ (.B1(_08198_),
    .Y(net16),
    .A1(_05094_),
    .A2(_08194_));
 sg13g2_mux4_1 _27475_ (.S0(_04923_),
    .A0(net1099),
    .A1(net1100),
    .A2(net1076),
    .A3(net1075),
    .S1(_06340_),
    .X(_08199_));
 sg13g2_mux4_1 _27476_ (.S0(_04923_),
    .A0(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A1(net1078),
    .A2(net1097),
    .A3(net1098),
    .S1(_06340_),
    .X(_08200_));
 sg13g2_nor2b_1 _27477_ (.A(\cpu.gpio.r_src_io[6][2] ),
    .B_N(_08200_),
    .Y(_08201_));
 sg13g2_a21oi_1 _27478_ (.A1(\cpu.gpio.r_src_io[6][2] ),
    .A2(_08199_),
    .Y(_08202_),
    .B1(_08201_));
 sg13g2_nand2b_1 _27479_ (.Y(_08203_),
    .B(net1074),
    .A_N(_04923_));
 sg13g2_nand3_1 _27480_ (.B(net1077),
    .C(_06340_),
    .A(_04923_),
    .Y(_08204_));
 sg13g2_o21ai_1 _27481_ (.B1(_08204_),
    .Y(_08205_),
    .A1(_06340_),
    .A2(_08203_));
 sg13g2_nand3_1 _27482_ (.B(\cpu.gpio.r_src_io[6][3] ),
    .C(_08205_),
    .A(_00106_),
    .Y(_08206_));
 sg13g2_o21ai_1 _27483_ (.B1(_08206_),
    .Y(net17),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .A2(_08202_));
 sg13g2_mux4_1 _27484_ (.S0(_05581_),
    .A0(net1099),
    .A1(net1100),
    .A2(net1076),
    .A3(net1075),
    .S1(_06342_),
    .X(_08207_));
 sg13g2_mux4_1 _27485_ (.S0(_05581_),
    .A0(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A1(net1078),
    .A2(net1097),
    .A3(net1098),
    .S1(_06342_),
    .X(_08208_));
 sg13g2_nor2b_1 _27486_ (.A(\cpu.gpio.r_src_io[7][2] ),
    .B_N(_08208_),
    .Y(_08209_));
 sg13g2_a21oi_1 _27487_ (.A1(\cpu.gpio.r_src_io[7][2] ),
    .A2(_08207_),
    .Y(_08210_),
    .B1(_08209_));
 sg13g2_nand2b_1 _27488_ (.Y(_08211_),
    .B(net1074),
    .A_N(_05581_));
 sg13g2_nand3_1 _27489_ (.B(net1077),
    .C(_06342_),
    .A(_05581_),
    .Y(_08212_));
 sg13g2_o21ai_1 _27490_ (.B1(_08212_),
    .Y(_08213_),
    .A1(_06342_),
    .A2(_08211_));
 sg13g2_nand3_1 _27491_ (.B(\cpu.gpio.r_src_io[7][3] ),
    .C(_08213_),
    .A(_00146_),
    .Y(_08214_));
 sg13g2_o21ai_1 _27492_ (.B1(_08214_),
    .Y(net18),
    .A1(\cpu.gpio.r_src_io[7][3] ),
    .A2(_08210_));
 sg13g2_xor2_1 _27493_ (.B(clknet_leaf_75_clk),
    .A(\cpu.r_clk_invert ),
    .X(net21));
 sg13g2_mux4_1 _27494_ (.S0(_05570_),
    .A0(net1099),
    .A1(net1100),
    .A2(_08042_),
    .A3(_08044_),
    .S1(_06345_),
    .X(_08215_));
 sg13g2_mux4_1 _27495_ (.S0(_05570_),
    .A0(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .A1(_07114_),
    .A2(_11998_),
    .A3(net1098),
    .S1(_06345_),
    .X(_08216_));
 sg13g2_nor2b_1 _27496_ (.A(\cpu.gpio.r_src_o[3][2] ),
    .B_N(_08216_),
    .Y(_08217_));
 sg13g2_a21oi_1 _27497_ (.A1(\cpu.gpio.r_src_o[3][2] ),
    .A2(_08215_),
    .Y(_08218_),
    .B1(_08217_));
 sg13g2_nand2b_1 _27498_ (.Y(_08219_),
    .B(_08046_),
    .A_N(_05570_));
 sg13g2_nand3_1 _27499_ (.B(_07756_),
    .C(_06345_),
    .A(_05570_),
    .Y(_08220_));
 sg13g2_o21ai_1 _27500_ (.B1(_08220_),
    .Y(_08221_),
    .A1(_06345_),
    .A2(_08219_));
 sg13g2_nand3_1 _27501_ (.B(\cpu.gpio.r_src_o[3][3] ),
    .C(_08221_),
    .A(_00149_),
    .Y(_08222_));
 sg13g2_o21ai_1 _27502_ (.B1(_08222_),
    .Y(net22),
    .A1(\cpu.gpio.r_src_o[3][3] ),
    .A2(_08218_));
 sg13g2_mux4_1 _27503_ (.S0(_04915_),
    .A0(_11977_),
    .A1(_11970_),
    .A2(net1076),
    .A3(net1075),
    .S1(_06348_),
    .X(_08223_));
 sg13g2_mux4_1 _27504_ (.S0(_04915_),
    .A0(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .A1(net1078),
    .A2(net1097),
    .A3(_11979_),
    .S1(_06348_),
    .X(_08224_));
 sg13g2_nor2b_1 _27505_ (.A(\cpu.gpio.r_src_o[4][2] ),
    .B_N(_08224_),
    .Y(_08225_));
 sg13g2_a21oi_1 _27506_ (.A1(\cpu.gpio.r_src_o[4][2] ),
    .A2(_08223_),
    .Y(_08226_),
    .B1(_08225_));
 sg13g2_nand2b_1 _27507_ (.Y(_08227_),
    .B(net1074),
    .A_N(_04915_));
 sg13g2_nand3_1 _27508_ (.B(net1077),
    .C(_06348_),
    .A(_04915_),
    .Y(_08228_));
 sg13g2_o21ai_1 _27509_ (.B1(_08228_),
    .Y(_08229_),
    .A1(_06348_),
    .A2(_08227_));
 sg13g2_nand3_1 _27510_ (.B(\cpu.gpio.r_src_o[4][3] ),
    .C(_08229_),
    .A(_00108_),
    .Y(_08230_));
 sg13g2_o21ai_1 _27511_ (.B1(_08230_),
    .Y(net23),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .A2(_08226_));
 sg13g2_mux4_1 _27512_ (.S0(_05580_),
    .A0(net1099),
    .A1(net1100),
    .A2(net1076),
    .A3(net1075),
    .S1(_06350_),
    .X(_08231_));
 sg13g2_mux4_1 _27513_ (.S0(_05580_),
    .A0(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .A1(net1078),
    .A2(net1097),
    .A3(net1098),
    .S1(_06350_),
    .X(_08232_));
 sg13g2_nor2b_1 _27514_ (.A(\cpu.gpio.r_src_o[5][2] ),
    .B_N(_08232_),
    .Y(_08233_));
 sg13g2_a21oi_1 _27515_ (.A1(\cpu.gpio.r_src_o[5][2] ),
    .A2(_08231_),
    .Y(_08234_),
    .B1(_08233_));
 sg13g2_nand2b_1 _27516_ (.Y(_08235_),
    .B(net1074),
    .A_N(_05580_));
 sg13g2_nand3_1 _27517_ (.B(net1077),
    .C(_06350_),
    .A(_05580_),
    .Y(_08236_));
 sg13g2_o21ai_1 _27518_ (.B1(_08236_),
    .Y(_08237_),
    .A1(_06350_),
    .A2(_08235_));
 sg13g2_nand3_1 _27519_ (.B(\cpu.gpio.r_src_o[5][3] ),
    .C(_08237_),
    .A(_00148_),
    .Y(_08238_));
 sg13g2_o21ai_1 _27520_ (.B1(_08238_),
    .Y(net24),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .A2(_08234_));
 sg13g2_mux4_1 _27521_ (.S0(_04933_),
    .A0(net1099),
    .A1(net1100),
    .A2(net1076),
    .A3(net1075),
    .S1(_07663_),
    .X(_08239_));
 sg13g2_mux4_1 _27522_ (.S0(_04933_),
    .A0(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .A1(net1078),
    .A2(net1097),
    .A3(net1098),
    .S1(_07663_),
    .X(_08240_));
 sg13g2_nor2b_1 _27523_ (.A(\cpu.gpio.r_src_o[6][2] ),
    .B_N(_08240_),
    .Y(_08241_));
 sg13g2_a21oi_1 _27524_ (.A1(\cpu.gpio.r_src_o[6][2] ),
    .A2(_08239_),
    .Y(_08242_),
    .B1(_08241_));
 sg13g2_nand2b_1 _27525_ (.Y(_08243_),
    .B(net1074),
    .A_N(_04933_));
 sg13g2_nand3_1 _27526_ (.B(net1077),
    .C(_07663_),
    .A(_04933_),
    .Y(_08244_));
 sg13g2_o21ai_1 _27527_ (.B1(_08244_),
    .Y(_08245_),
    .A1(_07663_),
    .A2(_08243_));
 sg13g2_nand3_1 _27528_ (.B(\cpu.gpio.r_src_o[6][3] ),
    .C(_08245_),
    .A(_00107_),
    .Y(_08246_));
 sg13g2_o21ai_1 _27529_ (.B1(_08246_),
    .Y(net25),
    .A1(\cpu.gpio.r_src_o[6][3] ),
    .A2(_08242_));
 sg13g2_mux4_1 _27530_ (.S0(_05575_),
    .A0(net1099),
    .A1(net1100),
    .A2(net1076),
    .A3(net1075),
    .S1(_06352_),
    .X(_08247_));
 sg13g2_mux4_1 _27531_ (.S0(_05575_),
    .A0(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .A1(net1078),
    .A2(net1097),
    .A3(net1098),
    .S1(_06352_),
    .X(_08248_));
 sg13g2_nor2b_1 _27532_ (.A(\cpu.gpio.r_src_o[7][2] ),
    .B_N(_08248_),
    .Y(_08249_));
 sg13g2_a21oi_1 _27533_ (.A1(\cpu.gpio.r_src_o[7][2] ),
    .A2(_08247_),
    .Y(_08250_),
    .B1(_08249_));
 sg13g2_nand2b_1 _27534_ (.Y(_08251_),
    .B(net1074),
    .A_N(_05575_));
 sg13g2_nand3_1 _27535_ (.B(net1077),
    .C(_06352_),
    .A(_05575_),
    .Y(_08252_));
 sg13g2_o21ai_1 _27536_ (.B1(_08252_),
    .Y(_08253_),
    .A1(_06352_),
    .A2(_08251_));
 sg13g2_nand3_1 _27537_ (.B(\cpu.gpio.r_src_o[7][3] ),
    .C(_08253_),
    .A(_00147_),
    .Y(_08254_));
 sg13g2_o21ai_1 _27538_ (.B1(_08254_),
    .Y(net26),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .A2(_08250_));
 sg13g2_dfrbp_1 _27539_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1131),
    .D(_00315_),
    .Q_N(_14894_),
    .Q(\cpu.intr.r_swi ));
 sg13g2_dfrbp_1 _27540_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1132),
    .D(_00316_),
    .Q_N(_14893_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[5] ));
 sg13g2_dfrbp_1 _27541_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1133),
    .D(_00317_),
    .Q_N(_14892_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[4] ));
 sg13g2_dfrbp_1 _27542_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1134),
    .D(_00318_),
    .Q_N(_14891_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[3] ));
 sg13g2_dfrbp_1 _27543_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1135),
    .D(_00319_),
    .Q_N(_14890_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[2] ));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _27545_ (.A(net6),
    .X(net4));
 sg13g2_buf_1 _27546_ (.A(net6),
    .X(net5));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1136),
    .D(_00320_),
    .Q_N(_14889_),
    .Q(\cpu.dcache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1137),
    .D(_00321_),
    .Q_N(_00103_),
    .Q(\cpu.dcache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1138),
    .D(_00322_),
    .Q_N(_00113_),
    .Q(\cpu.dcache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1139),
    .D(_00323_),
    .Q_N(_00124_),
    .Q(\cpu.dcache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1140),
    .D(_00324_),
    .Q_N(_00131_),
    .Q(\cpu.dcache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1141),
    .D(_00325_),
    .Q_N(_00143_),
    .Q(\cpu.dcache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1142),
    .D(_00326_),
    .Q_N(_00155_),
    .Q(\cpu.dcache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1143),
    .D(_00327_),
    .Q_N(_14888_),
    .Q(\cpu.dcache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1144),
    .D(_00328_),
    .Q_N(_00091_),
    .Q(\cpu.dcache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1145),
    .D(_00329_),
    .Q_N(_00101_),
    .Q(\cpu.dcache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1146),
    .D(_00330_),
    .Q_N(_00111_),
    .Q(\cpu.dcache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1147),
    .D(_00331_),
    .Q_N(_14887_),
    .Q(\cpu.dcache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1148),
    .D(_00332_),
    .Q_N(_00122_),
    .Q(\cpu.dcache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1149),
    .D(_00333_),
    .Q_N(_00129_),
    .Q(\cpu.dcache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1150),
    .D(_00334_),
    .Q_N(_00141_),
    .Q(\cpu.dcache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1151),
    .D(_00335_),
    .Q_N(_00153_),
    .Q(\cpu.dcache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1152),
    .D(_00336_),
    .Q_N(_00309_),
    .Q(\cpu.dcache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1153),
    .D(_00337_),
    .Q_N(_00092_),
    .Q(\cpu.dcache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1154),
    .D(_00338_),
    .Q_N(_00102_),
    .Q(\cpu.dcache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1155),
    .D(_00339_),
    .Q_N(_00112_),
    .Q(\cpu.dcache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1156),
    .D(_00340_),
    .Q_N(_00123_),
    .Q(\cpu.dcache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1157),
    .D(_00341_),
    .Q_N(_00130_),
    .Q(\cpu.dcache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1158),
    .D(_00342_),
    .Q_N(_14886_),
    .Q(\cpu.dcache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1159),
    .D(_00343_),
    .Q_N(_00142_),
    .Q(\cpu.dcache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1160),
    .D(_00344_),
    .Q_N(_00154_),
    .Q(\cpu.dcache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1161),
    .D(_00345_),
    .Q_N(_14885_),
    .Q(\cpu.dcache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1162),
    .D(_00346_),
    .Q_N(_00121_),
    .Q(\cpu.dcache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1163),
    .D(_00347_),
    .Q_N(_00128_),
    .Q(\cpu.dcache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1164),
    .D(_00348_),
    .Q_N(_00140_),
    .Q(\cpu.dcache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1165),
    .D(_00349_),
    .Q_N(_00152_),
    .Q(\cpu.dcache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1166),
    .D(_00350_),
    .Q_N(_00310_),
    .Q(\cpu.dcache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1167),
    .D(_00351_),
    .Q_N(_00093_),
    .Q(\cpu.dcache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1168),
    .D(_00352_),
    .Q_N(_14884_),
    .Q(\cpu.dcache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1169),
    .D(_00353_),
    .Q_N(_14883_),
    .Q(\cpu.dcache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1170),
    .D(_00354_),
    .Q_N(_14882_),
    .Q(\cpu.dcache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1171),
    .D(_00355_),
    .Q_N(_14881_),
    .Q(\cpu.dcache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1172),
    .D(_00356_),
    .Q_N(_14880_),
    .Q(\cpu.dcache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1173),
    .D(_00357_),
    .Q_N(_14879_),
    .Q(\cpu.dcache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1174),
    .D(_00358_),
    .Q_N(_14878_),
    .Q(\cpu.dcache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1175),
    .D(_00359_),
    .Q_N(_14877_),
    .Q(\cpu.dcache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1176),
    .D(_00360_),
    .Q_N(_14876_),
    .Q(\cpu.dcache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1177),
    .D(_00361_),
    .Q_N(_14875_),
    .Q(\cpu.dcache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1178),
    .D(_00362_),
    .Q_N(_14874_),
    .Q(\cpu.dcache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1179),
    .D(_00363_),
    .Q_N(_14873_),
    .Q(\cpu.dcache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1180),
    .D(_00364_),
    .Q_N(_14872_),
    .Q(\cpu.dcache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1181),
    .D(_00365_),
    .Q_N(_14871_),
    .Q(\cpu.dcache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1182),
    .D(_00366_),
    .Q_N(_14870_),
    .Q(\cpu.dcache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1183),
    .D(_00367_),
    .Q_N(_14869_),
    .Q(\cpu.dcache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1184),
    .D(_00368_),
    .Q_N(_14868_),
    .Q(\cpu.dcache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1185),
    .D(_00369_),
    .Q_N(_14867_),
    .Q(\cpu.dcache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1186),
    .D(_00370_),
    .Q_N(_14866_),
    .Q(\cpu.dcache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1187),
    .D(_00371_),
    .Q_N(_14865_),
    .Q(\cpu.dcache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1188),
    .D(_00372_),
    .Q_N(_14864_),
    .Q(\cpu.dcache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1189),
    .D(_00373_),
    .Q_N(_14863_),
    .Q(\cpu.dcache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1190),
    .D(_00374_),
    .Q_N(_14862_),
    .Q(\cpu.dcache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1191),
    .D(_00375_),
    .Q_N(_14861_),
    .Q(\cpu.dcache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1192),
    .D(_00376_),
    .Q_N(_14860_),
    .Q(\cpu.dcache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1193),
    .D(_00377_),
    .Q_N(_14859_),
    .Q(\cpu.dcache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1194),
    .D(_00378_),
    .Q_N(_14858_),
    .Q(\cpu.dcache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1195),
    .D(_00379_),
    .Q_N(_14857_),
    .Q(\cpu.dcache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1196),
    .D(_00380_),
    .Q_N(_14856_),
    .Q(\cpu.dcache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1197),
    .D(_00381_),
    .Q_N(_14855_),
    .Q(\cpu.dcache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1198),
    .D(_00382_),
    .Q_N(_14854_),
    .Q(\cpu.dcache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1199),
    .D(_00383_),
    .Q_N(_14853_),
    .Q(\cpu.dcache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1200),
    .D(_00384_),
    .Q_N(_14852_),
    .Q(\cpu.dcache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1201),
    .D(_00385_),
    .Q_N(_14851_),
    .Q(\cpu.dcache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1202),
    .D(_00386_),
    .Q_N(_14850_),
    .Q(\cpu.dcache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1203),
    .D(_00387_),
    .Q_N(_14849_),
    .Q(\cpu.dcache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1204),
    .D(_00388_),
    .Q_N(_14848_),
    .Q(\cpu.dcache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1205),
    .D(_00389_),
    .Q_N(_14847_),
    .Q(\cpu.dcache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1206),
    .D(_00390_),
    .Q_N(_14846_),
    .Q(\cpu.dcache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1207),
    .D(_00391_),
    .Q_N(_14845_),
    .Q(\cpu.dcache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1208),
    .D(_00392_),
    .Q_N(_14844_),
    .Q(\cpu.dcache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1209),
    .D(_00393_),
    .Q_N(_14843_),
    .Q(\cpu.dcache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1210),
    .D(_00394_),
    .Q_N(_14842_),
    .Q(\cpu.dcache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1211),
    .D(_00395_),
    .Q_N(_14841_),
    .Q(\cpu.dcache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1212),
    .D(_00396_),
    .Q_N(_14840_),
    .Q(\cpu.dcache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1213),
    .D(_00397_),
    .Q_N(_14839_),
    .Q(\cpu.dcache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1214),
    .D(_00398_),
    .Q_N(_14838_),
    .Q(\cpu.dcache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1215),
    .D(_00399_),
    .Q_N(_14837_),
    .Q(\cpu.dcache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1216),
    .D(_00400_),
    .Q_N(_14836_),
    .Q(\cpu.dcache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1217),
    .D(_00401_),
    .Q_N(_14835_),
    .Q(\cpu.dcache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1218),
    .D(_00402_),
    .Q_N(_14834_),
    .Q(\cpu.dcache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1219),
    .D(_00403_),
    .Q_N(_14833_),
    .Q(\cpu.dcache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1220),
    .D(_00404_),
    .Q_N(_14832_),
    .Q(\cpu.dcache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1221),
    .D(_00405_),
    .Q_N(_14831_),
    .Q(\cpu.dcache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1222),
    .D(_00406_),
    .Q_N(_14830_),
    .Q(\cpu.dcache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1223),
    .D(_00407_),
    .Q_N(_14829_),
    .Q(\cpu.dcache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1224),
    .D(_00408_),
    .Q_N(_14828_),
    .Q(\cpu.dcache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1225),
    .D(_00409_),
    .Q_N(_14827_),
    .Q(\cpu.dcache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1226),
    .D(_00410_),
    .Q_N(_14826_),
    .Q(\cpu.dcache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1227),
    .D(_00411_),
    .Q_N(_14825_),
    .Q(\cpu.dcache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1228),
    .D(_00412_),
    .Q_N(_14824_),
    .Q(\cpu.dcache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1229),
    .D(_00413_),
    .Q_N(_14823_),
    .Q(\cpu.dcache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1230),
    .D(_00414_),
    .Q_N(_14822_),
    .Q(\cpu.dcache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1231),
    .D(_00415_),
    .Q_N(_14821_),
    .Q(\cpu.dcache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1232),
    .D(_00416_),
    .Q_N(_14820_),
    .Q(\cpu.dcache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1233),
    .D(_00417_),
    .Q_N(_14819_),
    .Q(\cpu.dcache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1234),
    .D(_00418_),
    .Q_N(_14818_),
    .Q(\cpu.dcache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1235),
    .D(_00419_),
    .Q_N(_14817_),
    .Q(\cpu.dcache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1236),
    .D(_00420_),
    .Q_N(_14816_),
    .Q(\cpu.dcache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1237),
    .D(_00421_),
    .Q_N(_14815_),
    .Q(\cpu.dcache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1238),
    .D(_00422_),
    .Q_N(_14814_),
    .Q(\cpu.dcache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1239),
    .D(_00423_),
    .Q_N(_14813_),
    .Q(\cpu.dcache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1240),
    .D(_00424_),
    .Q_N(_14812_),
    .Q(\cpu.dcache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1241),
    .D(_00425_),
    .Q_N(_14811_),
    .Q(\cpu.dcache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1242),
    .D(_00426_),
    .Q_N(_14810_),
    .Q(\cpu.dcache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1243),
    .D(_00427_),
    .Q_N(_14809_),
    .Q(\cpu.dcache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1244),
    .D(_00428_),
    .Q_N(_14808_),
    .Q(\cpu.dcache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1245),
    .D(_00429_),
    .Q_N(_14807_),
    .Q(\cpu.dcache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1246),
    .D(_00430_),
    .Q_N(_14806_),
    .Q(\cpu.dcache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1247),
    .D(_00431_),
    .Q_N(_14805_),
    .Q(\cpu.dcache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1248),
    .D(_00432_),
    .Q_N(_14804_),
    .Q(\cpu.dcache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1249),
    .D(_00433_),
    .Q_N(_14803_),
    .Q(\cpu.dcache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1250),
    .D(_00434_),
    .Q_N(_14802_),
    .Q(\cpu.dcache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1251),
    .D(_00435_),
    .Q_N(_14801_),
    .Q(\cpu.dcache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1252),
    .D(_00436_),
    .Q_N(_14800_),
    .Q(\cpu.dcache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1253),
    .D(_00437_),
    .Q_N(_14799_),
    .Q(\cpu.dcache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1254),
    .D(_00438_),
    .Q_N(_14798_),
    .Q(\cpu.dcache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1255),
    .D(_00439_),
    .Q_N(_14797_),
    .Q(\cpu.dcache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1256),
    .D(_00440_),
    .Q_N(_14796_),
    .Q(\cpu.dcache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1257),
    .D(_00441_),
    .Q_N(_14795_),
    .Q(\cpu.dcache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1258),
    .D(_00442_),
    .Q_N(_14794_),
    .Q(\cpu.dcache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1259),
    .D(_00443_),
    .Q_N(_14793_),
    .Q(\cpu.dcache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1260),
    .D(_00444_),
    .Q_N(_14792_),
    .Q(\cpu.dcache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1261),
    .D(_00445_),
    .Q_N(_14791_),
    .Q(\cpu.dcache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1262),
    .D(_00446_),
    .Q_N(_14790_),
    .Q(\cpu.dcache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1263),
    .D(_00447_),
    .Q_N(_14789_),
    .Q(\cpu.dcache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1264),
    .D(_00448_),
    .Q_N(_14788_),
    .Q(\cpu.dcache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1265),
    .D(_00449_),
    .Q_N(_14787_),
    .Q(\cpu.dcache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1266),
    .D(_00450_),
    .Q_N(_14786_),
    .Q(\cpu.dcache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1267),
    .D(_00451_),
    .Q_N(_14785_),
    .Q(\cpu.dcache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1268),
    .D(_00452_),
    .Q_N(_14784_),
    .Q(\cpu.dcache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1269),
    .D(_00453_),
    .Q_N(_14783_),
    .Q(\cpu.dcache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1270),
    .D(_00454_),
    .Q_N(_14782_),
    .Q(\cpu.dcache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1271),
    .D(_00455_),
    .Q_N(_14781_),
    .Q(\cpu.dcache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1272),
    .D(_00456_),
    .Q_N(_14780_),
    .Q(\cpu.dcache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1273),
    .D(_00457_),
    .Q_N(_14779_),
    .Q(\cpu.dcache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1274),
    .D(_00458_),
    .Q_N(_14778_),
    .Q(\cpu.dcache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1275),
    .D(_00459_),
    .Q_N(_14777_),
    .Q(\cpu.dcache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1276),
    .D(_00460_),
    .Q_N(_14776_),
    .Q(\cpu.dcache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1277),
    .D(_00461_),
    .Q_N(_14775_),
    .Q(\cpu.dcache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1278),
    .D(_00462_),
    .Q_N(_14774_),
    .Q(\cpu.dcache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1279),
    .D(_00463_),
    .Q_N(_14773_),
    .Q(\cpu.dcache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1280),
    .D(_00464_),
    .Q_N(_14772_),
    .Q(\cpu.dcache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1281),
    .D(_00465_),
    .Q_N(_14771_),
    .Q(\cpu.dcache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1282),
    .D(_00466_),
    .Q_N(_14770_),
    .Q(\cpu.dcache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1283),
    .D(_00467_),
    .Q_N(_14769_),
    .Q(\cpu.dcache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1284),
    .D(_00468_),
    .Q_N(_14768_),
    .Q(\cpu.dcache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1285),
    .D(_00469_),
    .Q_N(_14767_),
    .Q(\cpu.dcache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1286),
    .D(_00470_),
    .Q_N(_14766_),
    .Q(\cpu.dcache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1287),
    .D(_00471_),
    .Q_N(_14765_),
    .Q(\cpu.dcache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1288),
    .D(_00472_),
    .Q_N(_14764_),
    .Q(\cpu.dcache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1289),
    .D(_00473_),
    .Q_N(_14763_),
    .Q(\cpu.dcache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1290),
    .D(_00474_),
    .Q_N(_14762_),
    .Q(\cpu.dcache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1291),
    .D(_00475_),
    .Q_N(_14761_),
    .Q(\cpu.dcache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1292),
    .D(_00476_),
    .Q_N(_14760_),
    .Q(\cpu.dcache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1293),
    .D(_00477_),
    .Q_N(_14759_),
    .Q(\cpu.dcache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1294),
    .D(_00478_),
    .Q_N(_14758_),
    .Q(\cpu.dcache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1295),
    .D(_00479_),
    .Q_N(_14757_),
    .Q(\cpu.dcache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1296),
    .D(_00480_),
    .Q_N(_14756_),
    .Q(\cpu.dcache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1297),
    .D(_00481_),
    .Q_N(_14755_),
    .Q(\cpu.dcache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1298),
    .D(_00482_),
    .Q_N(_14754_),
    .Q(\cpu.dcache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1299),
    .D(_00483_),
    .Q_N(_14753_),
    .Q(\cpu.dcache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1300),
    .D(_00484_),
    .Q_N(_14752_),
    .Q(\cpu.dcache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1301),
    .D(_00485_),
    .Q_N(_14751_),
    .Q(\cpu.dcache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1302),
    .D(_00486_),
    .Q_N(_14750_),
    .Q(\cpu.dcache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1303),
    .D(_00487_),
    .Q_N(_14749_),
    .Q(\cpu.dcache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1304),
    .D(_00488_),
    .Q_N(_14748_),
    .Q(\cpu.dcache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1305),
    .D(_00489_),
    .Q_N(_14747_),
    .Q(\cpu.dcache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1306),
    .D(_00490_),
    .Q_N(_14746_),
    .Q(\cpu.dcache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1307),
    .D(_00491_),
    .Q_N(_14745_),
    .Q(\cpu.dcache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1308),
    .D(_00492_),
    .Q_N(_14744_),
    .Q(\cpu.dcache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1309),
    .D(_00493_),
    .Q_N(_14743_),
    .Q(\cpu.dcache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1310),
    .D(_00494_),
    .Q_N(_14742_),
    .Q(\cpu.dcache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1311),
    .D(_00495_),
    .Q_N(_14741_),
    .Q(\cpu.dcache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1312),
    .D(_00496_),
    .Q_N(_14740_),
    .Q(\cpu.dcache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1313),
    .D(_00497_),
    .Q_N(_14739_),
    .Q(\cpu.dcache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1314),
    .D(_00498_),
    .Q_N(_14738_),
    .Q(\cpu.dcache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1315),
    .D(_00499_),
    .Q_N(_14737_),
    .Q(\cpu.dcache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1316),
    .D(_00500_),
    .Q_N(_14736_),
    .Q(\cpu.dcache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1317),
    .D(_00501_),
    .Q_N(_14735_),
    .Q(\cpu.dcache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1318),
    .D(_00502_),
    .Q_N(_14734_),
    .Q(\cpu.dcache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1319),
    .D(_00503_),
    .Q_N(_14733_),
    .Q(\cpu.dcache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1320),
    .D(_00504_),
    .Q_N(_14732_),
    .Q(\cpu.dcache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1321),
    .D(_00505_),
    .Q_N(_14731_),
    .Q(\cpu.dcache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1322),
    .D(_00506_),
    .Q_N(_14730_),
    .Q(\cpu.dcache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1323),
    .D(_00507_),
    .Q_N(_14729_),
    .Q(\cpu.dcache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1324),
    .D(_00508_),
    .Q_N(_14728_),
    .Q(\cpu.dcache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1325),
    .D(_00509_),
    .Q_N(_14727_),
    .Q(\cpu.dcache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1326),
    .D(_00510_),
    .Q_N(_14726_),
    .Q(\cpu.dcache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1327),
    .D(_00511_),
    .Q_N(_14725_),
    .Q(\cpu.dcache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1328),
    .D(_00512_),
    .Q_N(_14724_),
    .Q(\cpu.dcache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1329),
    .D(_00513_),
    .Q_N(_14723_),
    .Q(\cpu.dcache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1330),
    .D(_00514_),
    .Q_N(_14722_),
    .Q(\cpu.dcache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1331),
    .D(_00515_),
    .Q_N(_14721_),
    .Q(\cpu.dcache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1332),
    .D(_00516_),
    .Q_N(_14720_),
    .Q(\cpu.dcache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1333),
    .D(_00517_),
    .Q_N(_14719_),
    .Q(\cpu.dcache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1334),
    .D(_00518_),
    .Q_N(_14718_),
    .Q(\cpu.dcache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1335),
    .D(_00519_),
    .Q_N(_14717_),
    .Q(\cpu.dcache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1336),
    .D(_00520_),
    .Q_N(_14716_),
    .Q(\cpu.dcache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1337),
    .D(_00521_),
    .Q_N(_14715_),
    .Q(\cpu.dcache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1338),
    .D(_00522_),
    .Q_N(_14714_),
    .Q(\cpu.dcache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1339),
    .D(_00523_),
    .Q_N(_14713_),
    .Q(\cpu.dcache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1340),
    .D(_00524_),
    .Q_N(_14712_),
    .Q(\cpu.dcache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1341),
    .D(_00525_),
    .Q_N(_14711_),
    .Q(\cpu.dcache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1342),
    .D(_00526_),
    .Q_N(_14710_),
    .Q(\cpu.dcache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1343),
    .D(_00527_),
    .Q_N(_14709_),
    .Q(\cpu.dcache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1344),
    .D(_00528_),
    .Q_N(_14708_),
    .Q(\cpu.dcache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1345),
    .D(_00529_),
    .Q_N(_14707_),
    .Q(\cpu.dcache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1346),
    .D(_00530_),
    .Q_N(_14706_),
    .Q(\cpu.dcache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1347),
    .D(_00531_),
    .Q_N(_14705_),
    .Q(\cpu.dcache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1348),
    .D(_00532_),
    .Q_N(_14704_),
    .Q(\cpu.dcache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1349),
    .D(_00533_),
    .Q_N(_14703_),
    .Q(\cpu.dcache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1350),
    .D(_00534_),
    .Q_N(_14702_),
    .Q(\cpu.dcache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1351),
    .D(_00535_),
    .Q_N(_14701_),
    .Q(\cpu.dcache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1352),
    .D(_00536_),
    .Q_N(_14700_),
    .Q(\cpu.dcache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1353),
    .D(_00537_),
    .Q_N(_14699_),
    .Q(\cpu.dcache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1354),
    .D(_00538_),
    .Q_N(_14698_),
    .Q(\cpu.dcache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1355),
    .D(_00539_),
    .Q_N(_14697_),
    .Q(\cpu.dcache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1356),
    .D(_00540_),
    .Q_N(_14696_),
    .Q(\cpu.dcache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1357),
    .D(_00541_),
    .Q_N(_14695_),
    .Q(\cpu.dcache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1358),
    .D(_00542_),
    .Q_N(_14694_),
    .Q(\cpu.dcache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1359),
    .D(_00543_),
    .Q_N(_14693_),
    .Q(\cpu.dcache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1360),
    .D(_00544_),
    .Q_N(_14692_),
    .Q(\cpu.dcache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1361),
    .D(_00545_),
    .Q_N(_14691_),
    .Q(\cpu.dcache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1362),
    .D(_00546_),
    .Q_N(_14690_),
    .Q(\cpu.dcache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1363),
    .D(_00547_),
    .Q_N(_14689_),
    .Q(\cpu.dcache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1364),
    .D(_00548_),
    .Q_N(_14688_),
    .Q(\cpu.dcache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1365),
    .D(_00549_),
    .Q_N(_14687_),
    .Q(\cpu.dcache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1366),
    .D(_00550_),
    .Q_N(_14686_),
    .Q(\cpu.dcache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1367),
    .D(_00551_),
    .Q_N(_14685_),
    .Q(\cpu.dcache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1368),
    .D(_00552_),
    .Q_N(_14684_),
    .Q(\cpu.dcache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1369),
    .D(_00553_),
    .Q_N(_14683_),
    .Q(\cpu.dcache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1370),
    .D(_00554_),
    .Q_N(_14682_),
    .Q(\cpu.dcache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1371),
    .D(_00555_),
    .Q_N(_14681_),
    .Q(\cpu.dcache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1372),
    .D(_00556_),
    .Q_N(_14680_),
    .Q(\cpu.dcache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1373),
    .D(_00557_),
    .Q_N(_14679_),
    .Q(\cpu.dcache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1374),
    .D(_00558_),
    .Q_N(_14678_),
    .Q(\cpu.dcache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1375),
    .D(_00559_),
    .Q_N(_14677_),
    .Q(\cpu.dcache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1376),
    .D(_00560_),
    .Q_N(_14676_),
    .Q(\cpu.dcache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1377),
    .D(_00561_),
    .Q_N(_14675_),
    .Q(\cpu.dcache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1378),
    .D(_00562_),
    .Q_N(_14674_),
    .Q(\cpu.dcache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1379),
    .D(_00563_),
    .Q_N(_14673_),
    .Q(\cpu.dcache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1380),
    .D(_00564_),
    .Q_N(_14672_),
    .Q(\cpu.dcache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1381),
    .D(_00565_),
    .Q_N(_14671_),
    .Q(\cpu.dcache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1382),
    .D(_00566_),
    .Q_N(_14670_),
    .Q(\cpu.dcache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1383),
    .D(_00567_),
    .Q_N(_14669_),
    .Q(\cpu.dcache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1384),
    .D(_00568_),
    .Q_N(_14668_),
    .Q(\cpu.dcache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1385),
    .D(_00569_),
    .Q_N(_14667_),
    .Q(\cpu.dcache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1386),
    .D(_00570_),
    .Q_N(_14666_),
    .Q(\cpu.dcache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1387),
    .D(_00571_),
    .Q_N(_14665_),
    .Q(\cpu.dcache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1388),
    .D(_00572_),
    .Q_N(_14664_),
    .Q(\cpu.dcache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1389),
    .D(_00573_),
    .Q_N(_14663_),
    .Q(\cpu.dcache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1390),
    .D(_00574_),
    .Q_N(_14662_),
    .Q(\cpu.dcache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1391),
    .D(_00575_),
    .Q_N(_14661_),
    .Q(\cpu.dcache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1392),
    .D(_00576_),
    .Q_N(_14660_),
    .Q(\cpu.dcache.r_dirty[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1393),
    .D(_00577_),
    .Q_N(_14659_),
    .Q(\cpu.dcache.r_dirty[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1394),
    .D(_00578_),
    .Q_N(_14658_),
    .Q(\cpu.dcache.r_dirty[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1395),
    .D(_00579_),
    .Q_N(_14657_),
    .Q(\cpu.dcache.r_dirty[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1396),
    .D(_00580_),
    .Q_N(_14656_),
    .Q(\cpu.dcache.r_dirty[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1397),
    .D(_00581_),
    .Q_N(_14655_),
    .Q(\cpu.dcache.r_dirty[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1398),
    .D(_00582_),
    .Q_N(_14654_),
    .Q(\cpu.dcache.r_dirty[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1399),
    .D(_00583_),
    .Q_N(_14653_),
    .Q(\cpu.dcache.r_dirty[7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1400),
    .D(_00584_),
    .Q_N(_00313_),
    .Q(\cpu.dcache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1401),
    .D(_00585_),
    .Q_N(_14652_),
    .Q(\cpu.dcache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1402),
    .D(_00586_),
    .Q_N(_00274_),
    .Q(\cpu.dcache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1403),
    .D(_00587_),
    .Q_N(_00228_),
    .Q(\cpu.dcache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1404),
    .D(_00588_),
    .Q_N(_00244_),
    .Q(\cpu.dcache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1405),
    .D(_00589_),
    .Q_N(_00245_),
    .Q(\cpu.dcache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1406),
    .D(_00590_),
    .Q_N(_00246_),
    .Q(\cpu.dcache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1407),
    .D(_00591_),
    .Q_N(_00247_),
    .Q(\cpu.dcache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1408),
    .D(_00592_),
    .Q_N(_00248_),
    .Q(\cpu.dcache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1409),
    .D(_00593_),
    .Q_N(_14651_),
    .Q(\cpu.dcache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1410),
    .D(_00594_),
    .Q_N(_14650_),
    .Q(\cpu.dcache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1411),
    .D(_00595_),
    .Q_N(_14649_),
    .Q(\cpu.dcache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1412),
    .D(_00596_),
    .Q_N(_00249_),
    .Q(\cpu.dcache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1413),
    .D(_00597_),
    .Q_N(_00230_),
    .Q(\cpu.dcache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1414),
    .D(_00598_),
    .Q_N(_00232_),
    .Q(\cpu.dcache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1415),
    .D(_00599_),
    .Q_N(_00234_),
    .Q(\cpu.dcache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1416),
    .D(_00600_),
    .Q_N(_00236_),
    .Q(\cpu.dcache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1417),
    .D(_00601_),
    .Q_N(_00238_),
    .Q(\cpu.dcache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1418),
    .D(_00602_),
    .Q_N(_00240_),
    .Q(\cpu.dcache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1419),
    .D(_00603_),
    .Q_N(_00241_),
    .Q(\cpu.dcache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1420),
    .D(_00604_),
    .Q_N(_00242_),
    .Q(\cpu.dcache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1421),
    .D(_00605_),
    .Q_N(_00243_),
    .Q(\cpu.dcache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1422),
    .D(_00606_),
    .Q_N(_14648_),
    .Q(\cpu.dcache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1423),
    .D(_00607_),
    .Q_N(_14647_),
    .Q(\cpu.dcache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1424),
    .D(_00608_),
    .Q_N(_14646_),
    .Q(\cpu.dcache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1425),
    .D(_00609_),
    .Q_N(_14645_),
    .Q(\cpu.dcache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1426),
    .D(_00610_),
    .Q_N(_14644_),
    .Q(\cpu.dcache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1427),
    .D(_00611_),
    .Q_N(_14643_),
    .Q(\cpu.dcache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1428),
    .D(_00612_),
    .Q_N(_14642_),
    .Q(\cpu.dcache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1429),
    .D(_00613_),
    .Q_N(_14641_),
    .Q(\cpu.dcache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1430),
    .D(_00614_),
    .Q_N(_14640_),
    .Q(\cpu.dcache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1431),
    .D(_00615_),
    .Q_N(_14639_),
    .Q(\cpu.dcache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1432),
    .D(_00616_),
    .Q_N(_14638_),
    .Q(\cpu.dcache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1433),
    .D(_00617_),
    .Q_N(_14637_),
    .Q(\cpu.dcache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1434),
    .D(_00618_),
    .Q_N(_14636_),
    .Q(\cpu.dcache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1435),
    .D(_00619_),
    .Q_N(_14635_),
    .Q(\cpu.dcache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1436),
    .D(_00620_),
    .Q_N(_14634_),
    .Q(\cpu.dcache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1437),
    .D(_00621_),
    .Q_N(_14633_),
    .Q(\cpu.dcache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1438),
    .D(_00622_),
    .Q_N(_14632_),
    .Q(\cpu.dcache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1439),
    .D(_00623_),
    .Q_N(_14631_),
    .Q(\cpu.dcache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1440),
    .D(_00624_),
    .Q_N(_14630_),
    .Q(\cpu.dcache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1441),
    .D(_00625_),
    .Q_N(_14629_),
    .Q(\cpu.dcache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1442),
    .D(_00626_),
    .Q_N(_14628_),
    .Q(\cpu.dcache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1443),
    .D(_00627_),
    .Q_N(_14627_),
    .Q(\cpu.dcache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1444),
    .D(_00628_),
    .Q_N(_14626_),
    .Q(\cpu.dcache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1445),
    .D(_00629_),
    .Q_N(_14625_),
    .Q(\cpu.dcache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1446),
    .D(_00630_),
    .Q_N(_14624_),
    .Q(\cpu.dcache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1447),
    .D(_00631_),
    .Q_N(_14623_),
    .Q(\cpu.dcache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1448),
    .D(_00632_),
    .Q_N(_14622_),
    .Q(\cpu.dcache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1449),
    .D(_00633_),
    .Q_N(_14621_),
    .Q(\cpu.dcache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1450),
    .D(_00634_),
    .Q_N(_14620_),
    .Q(\cpu.dcache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1451),
    .D(_00635_),
    .Q_N(_14619_),
    .Q(\cpu.dcache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1452),
    .D(_00636_),
    .Q_N(_14618_),
    .Q(\cpu.dcache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1453),
    .D(_00637_),
    .Q_N(_14617_),
    .Q(\cpu.dcache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1454),
    .D(_00638_),
    .Q_N(_14616_),
    .Q(\cpu.dcache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1455),
    .D(_00639_),
    .Q_N(_14615_),
    .Q(\cpu.dcache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1456),
    .D(_00640_),
    .Q_N(_14614_),
    .Q(\cpu.dcache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1457),
    .D(_00641_),
    .Q_N(_14613_),
    .Q(\cpu.dcache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1458),
    .D(_00642_),
    .Q_N(_14612_),
    .Q(\cpu.dcache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1459),
    .D(_00643_),
    .Q_N(_14611_),
    .Q(\cpu.dcache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1460),
    .D(_00644_),
    .Q_N(_14610_),
    .Q(\cpu.dcache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1461),
    .D(_00645_),
    .Q_N(_14609_),
    .Q(\cpu.dcache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1462),
    .D(_00646_),
    .Q_N(_14608_),
    .Q(\cpu.dcache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1463),
    .D(_00647_),
    .Q_N(_14607_),
    .Q(\cpu.dcache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1464),
    .D(_00648_),
    .Q_N(_14606_),
    .Q(\cpu.dcache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1465),
    .D(_00649_),
    .Q_N(_14605_),
    .Q(\cpu.dcache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1466),
    .D(_00650_),
    .Q_N(_14604_),
    .Q(\cpu.dcache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1467),
    .D(_00651_),
    .Q_N(_14603_),
    .Q(\cpu.dcache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1468),
    .D(_00652_),
    .Q_N(_14602_),
    .Q(\cpu.dcache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1469),
    .D(_00653_),
    .Q_N(_14601_),
    .Q(\cpu.dcache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1470),
    .D(_00654_),
    .Q_N(_14600_),
    .Q(\cpu.dcache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1471),
    .D(_00655_),
    .Q_N(_14599_),
    .Q(\cpu.dcache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1472),
    .D(_00656_),
    .Q_N(_14598_),
    .Q(\cpu.dcache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1473),
    .D(_00657_),
    .Q_N(_14597_),
    .Q(\cpu.dcache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1474),
    .D(_00658_),
    .Q_N(_14596_),
    .Q(\cpu.dcache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1475),
    .D(_00659_),
    .Q_N(_14595_),
    .Q(\cpu.dcache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1476),
    .D(_00660_),
    .Q_N(_14594_),
    .Q(\cpu.dcache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1477),
    .D(_00661_),
    .Q_N(_14593_),
    .Q(\cpu.dcache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1478),
    .D(_00662_),
    .Q_N(_14592_),
    .Q(\cpu.dcache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1479),
    .D(_00663_),
    .Q_N(_14591_),
    .Q(\cpu.dcache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1480),
    .D(_00664_),
    .Q_N(_14590_),
    .Q(\cpu.dcache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1481),
    .D(_00665_),
    .Q_N(_14589_),
    .Q(\cpu.dcache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1482),
    .D(_00666_),
    .Q_N(_14588_),
    .Q(\cpu.dcache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1483),
    .D(_00667_),
    .Q_N(_14587_),
    .Q(\cpu.dcache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1484),
    .D(_00668_),
    .Q_N(_14586_),
    .Q(\cpu.dcache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1485),
    .D(_00669_),
    .Q_N(_14585_),
    .Q(\cpu.dcache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1486),
    .D(_00670_),
    .Q_N(_14584_),
    .Q(\cpu.dcache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1487),
    .D(_00671_),
    .Q_N(_14583_),
    .Q(\cpu.dcache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1488),
    .D(_00672_),
    .Q_N(_14582_),
    .Q(\cpu.dcache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1489),
    .D(_00673_),
    .Q_N(_14581_),
    .Q(\cpu.dcache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1490),
    .D(_00674_),
    .Q_N(_14580_),
    .Q(\cpu.dcache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1491),
    .D(_00675_),
    .Q_N(_14579_),
    .Q(\cpu.dcache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1492),
    .D(_00676_),
    .Q_N(_14578_),
    .Q(\cpu.dcache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1493),
    .D(_00677_),
    .Q_N(_14577_),
    .Q(\cpu.dcache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1494),
    .D(_00678_),
    .Q_N(_14576_),
    .Q(\cpu.dcache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1495),
    .D(_00679_),
    .Q_N(_14575_),
    .Q(\cpu.dcache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1496),
    .D(_00680_),
    .Q_N(_14574_),
    .Q(\cpu.dcache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1497),
    .D(_00681_),
    .Q_N(_14573_),
    .Q(\cpu.dcache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1498),
    .D(_00682_),
    .Q_N(_14572_),
    .Q(\cpu.dcache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1499),
    .D(_00683_),
    .Q_N(_14571_),
    .Q(\cpu.dcache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1500),
    .D(_00684_),
    .Q_N(_14570_),
    .Q(\cpu.dcache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1501),
    .D(_00685_),
    .Q_N(_14569_),
    .Q(\cpu.dcache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1502),
    .D(_00686_),
    .Q_N(_14568_),
    .Q(\cpu.dcache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1503),
    .D(_00687_),
    .Q_N(_14567_),
    .Q(\cpu.dcache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1504),
    .D(_00688_),
    .Q_N(_14566_),
    .Q(\cpu.dcache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1505),
    .D(_00689_),
    .Q_N(_14565_),
    .Q(\cpu.dcache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1506),
    .D(_00690_),
    .Q_N(_14564_),
    .Q(\cpu.dcache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1507),
    .D(_00691_),
    .Q_N(_14563_),
    .Q(\cpu.dcache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1508),
    .D(_00692_),
    .Q_N(_14562_),
    .Q(\cpu.dcache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1509),
    .D(_00693_),
    .Q_N(_14561_),
    .Q(\cpu.dcache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1510),
    .D(_00694_),
    .Q_N(_14560_),
    .Q(\cpu.dcache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1511),
    .D(_00695_),
    .Q_N(_14559_),
    .Q(\cpu.dcache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1512),
    .D(_00696_),
    .Q_N(_14558_),
    .Q(\cpu.dcache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1513),
    .D(_00697_),
    .Q_N(_14557_),
    .Q(\cpu.dcache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1514),
    .D(_00698_),
    .Q_N(_14556_),
    .Q(\cpu.dcache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1515),
    .D(_00699_),
    .Q_N(_14555_),
    .Q(\cpu.dcache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1516),
    .D(_00700_),
    .Q_N(_14554_),
    .Q(\cpu.dcache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1517),
    .D(_00701_),
    .Q_N(_14553_),
    .Q(\cpu.dcache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1518),
    .D(_00702_),
    .Q_N(_14552_),
    .Q(\cpu.dcache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1519),
    .D(_00703_),
    .Q_N(_14551_),
    .Q(\cpu.dcache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1520),
    .D(_00704_),
    .Q_N(_14550_),
    .Q(\cpu.dcache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1521),
    .D(_00705_),
    .Q_N(_14549_),
    .Q(\cpu.dcache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1522),
    .D(_00706_),
    .Q_N(_14548_),
    .Q(\cpu.dcache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1523),
    .D(_00707_),
    .Q_N(_14547_),
    .Q(\cpu.dcache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1524),
    .D(_00708_),
    .Q_N(_14546_),
    .Q(\cpu.dcache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1525),
    .D(_00709_),
    .Q_N(_14545_),
    .Q(\cpu.dcache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1526),
    .D(_00710_),
    .Q_N(_14544_),
    .Q(\cpu.dcache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1527),
    .D(_00711_),
    .Q_N(_14543_),
    .Q(\cpu.dcache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1528),
    .D(_00712_),
    .Q_N(_14542_),
    .Q(\cpu.dcache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1529),
    .D(_00713_),
    .Q_N(_14541_),
    .Q(\cpu.dcache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1530),
    .D(_00714_),
    .Q_N(_14540_),
    .Q(\cpu.dcache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1531),
    .D(_00715_),
    .Q_N(_14539_),
    .Q(\cpu.dcache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1532),
    .D(_00716_),
    .Q_N(_14538_),
    .Q(\cpu.dcache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1533),
    .D(_00717_),
    .Q_N(_14537_),
    .Q(\cpu.dcache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1534),
    .D(_00718_),
    .Q_N(_14536_),
    .Q(\cpu.dcache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1535),
    .D(_00719_),
    .Q_N(_14535_),
    .Q(\cpu.dcache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1536),
    .D(_00720_),
    .Q_N(_14534_),
    .Q(\cpu.dcache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1537),
    .D(_00721_),
    .Q_N(_14533_),
    .Q(\cpu.dcache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1538),
    .D(_00722_),
    .Q_N(_14532_),
    .Q(\cpu.dcache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1539),
    .D(_00723_),
    .Q_N(_14531_),
    .Q(\cpu.dcache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1540),
    .D(_00724_),
    .Q_N(_14530_),
    .Q(\cpu.dcache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1541),
    .D(_00725_),
    .Q_N(_14529_),
    .Q(\cpu.dcache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1542),
    .D(_00726_),
    .Q_N(_14528_),
    .Q(\cpu.dcache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1543),
    .D(_00727_),
    .Q_N(_14527_),
    .Q(\cpu.dcache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1544),
    .D(_00728_),
    .Q_N(_14526_),
    .Q(\cpu.dcache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1545),
    .D(_00729_),
    .Q_N(_14525_),
    .Q(\cpu.dcache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1546),
    .D(_00730_),
    .Q_N(_14524_),
    .Q(\cpu.dcache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1547),
    .D(_00731_),
    .Q_N(_14523_),
    .Q(\cpu.dcache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1548),
    .D(_00732_),
    .Q_N(_14522_),
    .Q(\cpu.dcache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1549),
    .D(_00733_),
    .Q_N(_14521_),
    .Q(\cpu.dcache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1550),
    .D(_00734_),
    .Q_N(_14520_),
    .Q(\cpu.dcache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1551),
    .D(_00735_),
    .Q_N(_14519_),
    .Q(\cpu.dcache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1552),
    .D(_00736_),
    .Q_N(_14518_),
    .Q(\cpu.dcache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1553),
    .D(_00737_),
    .Q_N(_14517_),
    .Q(\cpu.dcache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1554),
    .D(_00738_),
    .Q_N(_14516_),
    .Q(\cpu.dcache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1555),
    .D(_00739_),
    .Q_N(_14515_),
    .Q(\cpu.dcache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1556),
    .D(_00740_),
    .Q_N(_14514_),
    .Q(\cpu.dcache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1557),
    .D(_00741_),
    .Q_N(_14513_),
    .Q(\cpu.dcache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1558),
    .D(_00742_),
    .Q_N(_14512_),
    .Q(\cpu.dcache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1559),
    .D(_00743_),
    .Q_N(_14511_),
    .Q(\cpu.dcache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1560),
    .D(_00744_),
    .Q_N(_14510_),
    .Q(\cpu.dcache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1561),
    .D(_00745_),
    .Q_N(_14509_),
    .Q(\cpu.dcache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1562),
    .D(_00746_),
    .Q_N(_14508_),
    .Q(\cpu.dcache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_br$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1563),
    .D(_00747_),
    .Q_N(_14507_),
    .Q(\cpu.br ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[0]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1564),
    .D(_00748_),
    .Q_N(_00296_),
    .Q(\cpu.cond[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[1]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1565),
    .D(_00749_),
    .Q_N(_14506_),
    .Q(\cpu.cond[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[2]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1566),
    .D(_00750_),
    .Q_N(_00271_),
    .Q(\cpu.cond[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_div$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1567),
    .D(_00751_),
    .Q_N(_14505_),
    .Q(\cpu.dec.div ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_all$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1568),
    .D(_00752_),
    .Q_N(_14504_),
    .Q(\cpu.dec.do_flush_all ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_write$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1569),
    .D(_00753_),
    .Q_N(_14503_),
    .Q(\cpu.dec.do_flush_write ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[0]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1570),
    .D(_00754_),
    .Q_N(_14502_),
    .Q(\cpu.dec.imm[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[10]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1571),
    .D(_00755_),
    .Q_N(_14501_),
    .Q(\cpu.dec.imm[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[11]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1572),
    .D(_00756_),
    .Q_N(_14500_),
    .Q(\cpu.dec.imm[11] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[12]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1573),
    .D(_00757_),
    .Q_N(_14499_),
    .Q(\cpu.dec.imm[12] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[13]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1574),
    .D(_00758_),
    .Q_N(_14498_),
    .Q(\cpu.dec.imm[13] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[14]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1575),
    .D(_00759_),
    .Q_N(_14497_),
    .Q(\cpu.dec.imm[14] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[15]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1576),
    .D(_00760_),
    .Q_N(_14496_),
    .Q(\cpu.dec.imm[15] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[1]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1577),
    .D(_00761_),
    .Q_N(_14495_),
    .Q(\cpu.dec.imm[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[2]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1578),
    .D(_00762_),
    .Q_N(_14494_),
    .Q(\cpu.dec.imm[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[3]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1579),
    .D(_00763_),
    .Q_N(_14493_),
    .Q(\cpu.dec.imm[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[4]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1580),
    .D(_00764_),
    .Q_N(_14492_),
    .Q(\cpu.dec.imm[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[5]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1581),
    .D(_00765_),
    .Q_N(_14491_),
    .Q(\cpu.dec.imm[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[6]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1582),
    .D(_00766_),
    .Q_N(_14490_),
    .Q(\cpu.dec.imm[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[7]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1583),
    .D(_00767_),
    .Q_N(_14489_),
    .Q(\cpu.dec.imm[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[8]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1584),
    .D(_00768_),
    .Q_N(_14488_),
    .Q(\cpu.dec.imm[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[9]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1585),
    .D(_00769_),
    .Q_N(_14487_),
    .Q(\cpu.dec.imm[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_inv_mmu$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1586),
    .D(_00770_),
    .Q_N(_14486_),
    .Q(\cpu.dec.do_inv_mmu ));
 sg13g2_dfrbp_1 \cpu.dec.r_io$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1587),
    .D(_00771_),
    .Q_N(_14485_),
    .Q(\cpu.dec.io ));
 sg13g2_dfrbp_1 \cpu.dec.r_jmp$_SDFFCE_PP0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1588),
    .D(_00772_),
    .Q_N(_00256_),
    .Q(\cpu.dec.jmp ));
 sg13g2_dfrbp_1 \cpu.dec.r_load$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1589),
    .D(_00773_),
    .Q_N(_14484_),
    .Q(\cpu.dec.load ));
 sg13g2_dfrbp_1 \cpu.dec.r_mult$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1590),
    .D(_00774_),
    .Q_N(_14483_),
    .Q(\cpu.dec.mult ));
 sg13g2_dfrbp_1 \cpu.dec.r_needs_rs2$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1591),
    .D(_00775_),
    .Q_N(_14895_),
    .Q(\cpu.dec.needs_rs2 ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[10]$_DFF_P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1592),
    .D(_00011_),
    .Q_N(_14896_),
    .Q(\cpu.dec.r_op[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[1]$_DFF_P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1593),
    .D(_00012_),
    .Q_N(_14897_),
    .Q(\cpu.dec.r_op[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[2]$_DFF_P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1594),
    .D(_00013_),
    .Q_N(_14898_),
    .Q(\cpu.dec.r_op[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[3]$_DFF_P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1595),
    .D(_00014_),
    .Q_N(_14899_),
    .Q(\cpu.dec.r_op[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[4]$_DFF_P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1596),
    .D(_00015_),
    .Q_N(_14900_),
    .Q(\cpu.dec.r_op[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[5]$_DFF_P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1597),
    .D(_00016_),
    .Q_N(_14901_),
    .Q(\cpu.dec.r_op[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[6]$_DFF_P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1598),
    .D(_00017_),
    .Q_N(_14902_),
    .Q(\cpu.dec.r_op[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[7]$_DFF_P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1599),
    .D(_00018_),
    .Q_N(_14903_),
    .Q(\cpu.dec.r_op[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[8]$_DFF_P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1600),
    .D(_00019_),
    .Q_N(_14904_),
    .Q(\cpu.dec.r_op[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[9]$_DFF_P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1601),
    .D(_00020_),
    .Q_N(_14482_),
    .Q(\cpu.dec.r_op[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[0]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1602),
    .D(_00776_),
    .Q_N(_14481_),
    .Q(\cpu.dec.r_rd[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[1]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1603),
    .D(_00777_),
    .Q_N(_14480_),
    .Q(\cpu.dec.r_rd[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1604),
    .D(_00778_),
    .Q_N(_14479_),
    .Q(\cpu.dec.r_rd[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[3]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1605),
    .D(_00779_),
    .Q_N(_14905_),
    .Q(\cpu.dec.r_rd[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_ready$_DFF_P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1606),
    .D(_00052_),
    .Q_N(_14478_),
    .Q(\cpu.dec.iready ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[0]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1607),
    .D(_00780_),
    .Q_N(_14477_),
    .Q(\cpu.dec.r_rs1[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[1]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1608),
    .D(_00781_),
    .Q_N(_14476_),
    .Q(\cpu.dec.r_rs1[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[2]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1609),
    .D(_00782_),
    .Q_N(_14475_),
    .Q(\cpu.dec.r_rs1[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[3]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1610),
    .D(_00783_),
    .Q_N(_14474_),
    .Q(\cpu.dec.r_rs1[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[0]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1611),
    .D(_00784_),
    .Q_N(_14473_),
    .Q(\cpu.dec.r_rs2[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[1]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1612),
    .D(_00785_),
    .Q_N(_14472_),
    .Q(\cpu.dec.r_rs2[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[2]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1613),
    .D(_00786_),
    .Q_N(_14471_),
    .Q(\cpu.dec.r_rs2[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[3]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1614),
    .D(_00787_),
    .Q_N(_14470_),
    .Q(\cpu.dec.r_rs2[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_inv$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1615),
    .D(_00788_),
    .Q_N(_14469_),
    .Q(\cpu.dec.r_rs2_inv ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_pc$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1616),
    .D(_00789_),
    .Q_N(_14468_),
    .Q(\cpu.dec.r_rs2_pc ));
 sg13g2_dfrbp_1 \cpu.dec.r_set_cc$_SDFFCE_PP0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1617),
    .D(_00790_),
    .Q_N(_14467_),
    .Q(\cpu.dec.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.dec.r_store$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1618),
    .D(_00791_),
    .Q_N(_00308_),
    .Q(\cpu.dec.r_store ));
 sg13g2_dfrbp_1 \cpu.dec.r_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1619),
    .D(_00792_),
    .Q_N(_14466_),
    .Q(\cpu.dec.r_swapsp ));
 sg13g2_dfrbp_1 \cpu.dec.r_sys_call$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1620),
    .D(_00793_),
    .Q_N(_00272_),
    .Q(\cpu.dec.r_sys_call ));
 sg13g2_dfrbp_1 \cpu.dec.r_trap$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1621),
    .D(_00794_),
    .Q_N(_14465_),
    .Q(\cpu.dec.r_trap ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1622),
    .D(_00795_),
    .Q_N(_14464_),
    .Q(\cpu.ex.genblk3.r_mmu_d_proxy ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1623),
    .D(_00796_),
    .Q_N(_00192_),
    .Q(\cpu.ex.genblk3.r_mmu_enable ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1624),
    .D(_00797_),
    .Q_N(_14906_),
    .Q(\cpu.ex.genblk3.r_prev_supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_supmode$_DFF_P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1625),
    .D(\cpu.ex.genblk3.c_supmode ),
    .Q_N(_00193_),
    .Q(\cpu.dec.supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1626),
    .D(_00798_),
    .Q_N(_14463_),
    .Q(\cpu.dec.user_io ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1627),
    .D(_00799_),
    .Q_N(_14462_),
    .Q(\cpu.ex.r_10[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[10]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1628),
    .D(_00800_),
    .Q_N(_14461_),
    .Q(\cpu.ex.r_10[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[11]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1629),
    .D(_00801_),
    .Q_N(_14460_),
    .Q(\cpu.ex.r_10[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[12]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1630),
    .D(_00802_),
    .Q_N(_14459_),
    .Q(\cpu.ex.r_10[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[13]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1631),
    .D(_00803_),
    .Q_N(_14458_),
    .Q(\cpu.ex.r_10[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[14]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1632),
    .D(_00804_),
    .Q_N(_14457_),
    .Q(\cpu.ex.r_10[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[15]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1633),
    .D(_00805_),
    .Q_N(_14456_),
    .Q(\cpu.ex.r_10[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[1]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1634),
    .D(_00806_),
    .Q_N(_14455_),
    .Q(\cpu.ex.r_10[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[2]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1635),
    .D(_00807_),
    .Q_N(_14454_),
    .Q(\cpu.ex.r_10[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[3]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1636),
    .D(_00808_),
    .Q_N(_14453_),
    .Q(\cpu.ex.r_10[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[4]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1637),
    .D(_00809_),
    .Q_N(_14452_),
    .Q(\cpu.ex.r_10[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[5]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1638),
    .D(_00810_),
    .Q_N(_14451_),
    .Q(\cpu.ex.r_10[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[6]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1639),
    .D(_00811_),
    .Q_N(_14450_),
    .Q(\cpu.ex.r_10[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[7]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1640),
    .D(_00812_),
    .Q_N(_14449_),
    .Q(\cpu.ex.r_10[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[8]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1641),
    .D(_00813_),
    .Q_N(_14448_),
    .Q(\cpu.ex.r_10[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[9]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1642),
    .D(_00814_),
    .Q_N(_14447_),
    .Q(\cpu.ex.r_10[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1643),
    .D(_00815_),
    .Q_N(_14446_),
    .Q(\cpu.ex.r_11[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[10]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1644),
    .D(_00816_),
    .Q_N(_14445_),
    .Q(\cpu.ex.r_11[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[11]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1645),
    .D(_00817_),
    .Q_N(_14444_),
    .Q(\cpu.ex.r_11[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[12]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1646),
    .D(_00818_),
    .Q_N(_14443_),
    .Q(\cpu.ex.r_11[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[13]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1647),
    .D(_00819_),
    .Q_N(_14442_),
    .Q(\cpu.ex.r_11[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[14]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1648),
    .D(_00820_),
    .Q_N(_14441_),
    .Q(\cpu.ex.r_11[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[15]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1649),
    .D(_00821_),
    .Q_N(_14440_),
    .Q(\cpu.ex.r_11[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[1]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1650),
    .D(_00822_),
    .Q_N(_14439_),
    .Q(\cpu.ex.r_11[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[2]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1651),
    .D(_00823_),
    .Q_N(_14438_),
    .Q(\cpu.ex.r_11[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[3]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1652),
    .D(_00824_),
    .Q_N(_14437_),
    .Q(\cpu.ex.r_11[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[4]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1653),
    .D(_00825_),
    .Q_N(_14436_),
    .Q(\cpu.ex.r_11[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[5]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1654),
    .D(_00826_),
    .Q_N(_14435_),
    .Q(\cpu.ex.r_11[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[6]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1655),
    .D(_00827_),
    .Q_N(_14434_),
    .Q(\cpu.ex.r_11[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[7]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1656),
    .D(_00828_),
    .Q_N(_14433_),
    .Q(\cpu.ex.r_11[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[8]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1657),
    .D(_00829_),
    .Q_N(_14432_),
    .Q(\cpu.ex.r_11[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[9]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1658),
    .D(_00830_),
    .Q_N(_14431_),
    .Q(\cpu.ex.r_11[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[0]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1659),
    .D(_00831_),
    .Q_N(_14430_),
    .Q(\cpu.ex.r_12[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[10]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1660),
    .D(_00832_),
    .Q_N(_14429_),
    .Q(\cpu.ex.r_12[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[11]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1661),
    .D(_00833_),
    .Q_N(_14428_),
    .Q(\cpu.ex.r_12[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[12]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1662),
    .D(_00834_),
    .Q_N(_14427_),
    .Q(\cpu.ex.r_12[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[13]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1663),
    .D(_00835_),
    .Q_N(_14426_),
    .Q(\cpu.ex.r_12[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[14]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1664),
    .D(_00836_),
    .Q_N(_14425_),
    .Q(\cpu.ex.r_12[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[15]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1665),
    .D(_00837_),
    .Q_N(_14424_),
    .Q(\cpu.ex.r_12[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[1]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1666),
    .D(_00838_),
    .Q_N(_14423_),
    .Q(\cpu.ex.r_12[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[2]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1667),
    .D(_00839_),
    .Q_N(_14422_),
    .Q(\cpu.ex.r_12[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[3]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1668),
    .D(_00840_),
    .Q_N(_14421_),
    .Q(\cpu.ex.r_12[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[4]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1669),
    .D(_00841_),
    .Q_N(_14420_),
    .Q(\cpu.ex.r_12[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[5]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1670),
    .D(_00842_),
    .Q_N(_14419_),
    .Q(\cpu.ex.r_12[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[6]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1671),
    .D(_00843_),
    .Q_N(_14418_),
    .Q(\cpu.ex.r_12[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[7]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1672),
    .D(_00844_),
    .Q_N(_14417_),
    .Q(\cpu.ex.r_12[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[8]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1673),
    .D(_00845_),
    .Q_N(_14416_),
    .Q(\cpu.ex.r_12[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[9]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1674),
    .D(_00846_),
    .Q_N(_14415_),
    .Q(\cpu.ex.r_12[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[0]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1675),
    .D(_00847_),
    .Q_N(_14414_),
    .Q(\cpu.ex.r_13[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[10]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1676),
    .D(_00848_),
    .Q_N(_14413_),
    .Q(\cpu.ex.r_13[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[11]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1677),
    .D(_00849_),
    .Q_N(_14412_),
    .Q(\cpu.ex.r_13[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[12]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1678),
    .D(_00850_),
    .Q_N(_14411_),
    .Q(\cpu.ex.r_13[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[13]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1679),
    .D(_00851_),
    .Q_N(_14410_),
    .Q(\cpu.ex.r_13[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[14]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1680),
    .D(_00852_),
    .Q_N(_14409_),
    .Q(\cpu.ex.r_13[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[15]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1681),
    .D(_00853_),
    .Q_N(_14408_),
    .Q(\cpu.ex.r_13[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[1]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1682),
    .D(_00854_),
    .Q_N(_14407_),
    .Q(\cpu.ex.r_13[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[2]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1683),
    .D(_00855_),
    .Q_N(_14406_),
    .Q(\cpu.ex.r_13[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[3]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1684),
    .D(_00856_),
    .Q_N(_14405_),
    .Q(\cpu.ex.r_13[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[4]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1685),
    .D(_00857_),
    .Q_N(_14404_),
    .Q(\cpu.ex.r_13[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[5]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1686),
    .D(_00858_),
    .Q_N(_14403_),
    .Q(\cpu.ex.r_13[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[6]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1687),
    .D(_00859_),
    .Q_N(_14402_),
    .Q(\cpu.ex.r_13[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[7]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1688),
    .D(_00860_),
    .Q_N(_14401_),
    .Q(\cpu.ex.r_13[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[8]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1689),
    .D(_00861_),
    .Q_N(_14400_),
    .Q(\cpu.ex.r_13[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[9]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1690),
    .D(_00862_),
    .Q_N(_14399_),
    .Q(\cpu.ex.r_13[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1691),
    .D(_00863_),
    .Q_N(_14398_),
    .Q(\cpu.ex.r_14[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[10]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1692),
    .D(_00864_),
    .Q_N(_14397_),
    .Q(\cpu.ex.r_14[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[11]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1693),
    .D(_00865_),
    .Q_N(_14396_),
    .Q(\cpu.ex.r_14[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[12]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1694),
    .D(_00866_),
    .Q_N(_14395_),
    .Q(\cpu.ex.r_14[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[13]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1695),
    .D(_00867_),
    .Q_N(_14394_),
    .Q(\cpu.ex.r_14[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[14]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1696),
    .D(_00868_),
    .Q_N(_14393_),
    .Q(\cpu.ex.r_14[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[15]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1697),
    .D(_00869_),
    .Q_N(_14392_),
    .Q(\cpu.ex.r_14[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[1]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1698),
    .D(_00870_),
    .Q_N(_14391_),
    .Q(\cpu.ex.r_14[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[2]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1699),
    .D(_00871_),
    .Q_N(_14390_),
    .Q(\cpu.ex.r_14[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[3]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1700),
    .D(_00872_),
    .Q_N(_14389_),
    .Q(\cpu.ex.r_14[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[4]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1701),
    .D(_00873_),
    .Q_N(_14388_),
    .Q(\cpu.ex.r_14[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[5]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1702),
    .D(_00874_),
    .Q_N(_14387_),
    .Q(\cpu.ex.r_14[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[6]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1703),
    .D(_00875_),
    .Q_N(_14386_),
    .Q(\cpu.ex.r_14[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[7]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1704),
    .D(_00876_),
    .Q_N(_14385_),
    .Q(\cpu.ex.r_14[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[8]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1705),
    .D(_00877_),
    .Q_N(_14384_),
    .Q(\cpu.ex.r_14[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[9]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1706),
    .D(_00878_),
    .Q_N(_14383_),
    .Q(\cpu.ex.r_14[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[0]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1707),
    .D(_00879_),
    .Q_N(_14382_),
    .Q(\cpu.ex.r_15[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[10]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1708),
    .D(_00880_),
    .Q_N(_00266_),
    .Q(\cpu.ex.r_15[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[11]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1709),
    .D(_00881_),
    .Q_N(_00267_),
    .Q(\cpu.ex.r_15[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[12]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1710),
    .D(_00882_),
    .Q_N(_00268_),
    .Q(\cpu.ex.r_15[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[13]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1711),
    .D(_00883_),
    .Q_N(_00269_),
    .Q(\cpu.ex.r_15[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[14]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1712),
    .D(_00884_),
    .Q_N(_00270_),
    .Q(\cpu.ex.r_15[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[15]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1713),
    .D(_00885_),
    .Q_N(_14381_),
    .Q(\cpu.ex.r_15[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[1]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1714),
    .D(_00886_),
    .Q_N(_00257_),
    .Q(\cpu.ex.r_15[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[2]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1715),
    .D(_00887_),
    .Q_N(_00258_),
    .Q(\cpu.ex.r_15[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[3]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1716),
    .D(_00888_),
    .Q_N(_00259_),
    .Q(\cpu.ex.r_15[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[4]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1717),
    .D(_00889_),
    .Q_N(_00260_),
    .Q(\cpu.ex.r_15[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[5]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1718),
    .D(_00890_),
    .Q_N(_00261_),
    .Q(\cpu.ex.r_15[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[6]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1719),
    .D(_00891_),
    .Q_N(_00262_),
    .Q(\cpu.ex.r_15[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[7]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1720),
    .D(_00892_),
    .Q_N(_00263_),
    .Q(\cpu.ex.r_15[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[8]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1721),
    .D(_00893_),
    .Q_N(_00264_),
    .Q(\cpu.ex.r_15[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[9]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1722),
    .D(_00894_),
    .Q_N(_00265_),
    .Q(\cpu.ex.r_15[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[0]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1723),
    .D(_00895_),
    .Q_N(_14380_),
    .Q(\cpu.ex.r_8[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[10]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1724),
    .D(_00896_),
    .Q_N(_14379_),
    .Q(\cpu.ex.r_8[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[11]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1725),
    .D(_00897_),
    .Q_N(_14378_),
    .Q(\cpu.ex.r_8[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[12]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1726),
    .D(_00898_),
    .Q_N(_14377_),
    .Q(\cpu.ex.r_8[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1727),
    .D(_00899_),
    .Q_N(_14376_),
    .Q(\cpu.ex.r_8[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[14]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1728),
    .D(_00900_),
    .Q_N(_14375_),
    .Q(\cpu.ex.r_8[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[15]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1729),
    .D(_00901_),
    .Q_N(_14374_),
    .Q(\cpu.ex.r_8[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[1]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1730),
    .D(_00902_),
    .Q_N(_14373_),
    .Q(\cpu.ex.r_8[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[2]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1731),
    .D(_00903_),
    .Q_N(_14372_),
    .Q(\cpu.ex.r_8[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[3]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1732),
    .D(_00904_),
    .Q_N(_14371_),
    .Q(\cpu.ex.r_8[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[4]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1733),
    .D(_00905_),
    .Q_N(_14370_),
    .Q(\cpu.ex.r_8[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[5]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1734),
    .D(_00906_),
    .Q_N(_14369_),
    .Q(\cpu.ex.r_8[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[6]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1735),
    .D(_00907_),
    .Q_N(_14368_),
    .Q(\cpu.ex.r_8[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[7]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1736),
    .D(_00908_),
    .Q_N(_14367_),
    .Q(\cpu.ex.r_8[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[8]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1737),
    .D(_00909_),
    .Q_N(_14366_),
    .Q(\cpu.ex.r_8[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[9]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1738),
    .D(_00910_),
    .Q_N(_14365_),
    .Q(\cpu.ex.r_8[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1739),
    .D(_00911_),
    .Q_N(_14364_),
    .Q(\cpu.ex.r_9[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[10]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1740),
    .D(_00912_),
    .Q_N(_14363_),
    .Q(\cpu.ex.r_9[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[11]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1741),
    .D(_00913_),
    .Q_N(_14362_),
    .Q(\cpu.ex.r_9[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[12]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1742),
    .D(_00914_),
    .Q_N(_14361_),
    .Q(\cpu.ex.r_9[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[13]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1743),
    .D(_00915_),
    .Q_N(_14360_),
    .Q(\cpu.ex.r_9[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[14]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1744),
    .D(_00916_),
    .Q_N(_14359_),
    .Q(\cpu.ex.r_9[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[15]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1745),
    .D(_00917_),
    .Q_N(_14358_),
    .Q(\cpu.ex.r_9[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[1]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1746),
    .D(_00918_),
    .Q_N(_14357_),
    .Q(\cpu.ex.r_9[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[2]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1747),
    .D(_00919_),
    .Q_N(_14356_),
    .Q(\cpu.ex.r_9[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[3]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1748),
    .D(_00920_),
    .Q_N(_14355_),
    .Q(\cpu.ex.r_9[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[4]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1749),
    .D(_00921_),
    .Q_N(_14354_),
    .Q(\cpu.ex.r_9[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[5]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1750),
    .D(_00922_),
    .Q_N(_14353_),
    .Q(\cpu.ex.r_9[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[6]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1751),
    .D(_00923_),
    .Q_N(_14352_),
    .Q(\cpu.ex.r_9[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[7]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1752),
    .D(_00924_),
    .Q_N(_14351_),
    .Q(\cpu.ex.r_9[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[8]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1753),
    .D(_00925_),
    .Q_N(_14350_),
    .Q(\cpu.ex.r_9[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[9]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1754),
    .D(_00926_),
    .Q_N(_14907_),
    .Q(\cpu.ex.r_9[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_branch_stall$_DFF_P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1755),
    .D(_00053_),
    .Q_N(_14349_),
    .Q(\cpu.ex.r_branch_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_cc$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1756),
    .D(_00927_),
    .Q_N(_14348_),
    .Q(\cpu.ex.r_cc ));
 sg13g2_dfrbp_1 \cpu.ex.r_d_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1757),
    .D(_00928_),
    .Q_N(_14908_),
    .Q(\cpu.d_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_div_running$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1758),
    .D(\cpu.ex.c_div_running ),
    .Q_N(_14347_),
    .Q(\cpu.ex.r_div_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[0]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1759),
    .D(_00929_),
    .Q_N(_14346_),
    .Q(\cpu.ex.r_epc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[10]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1760),
    .D(_00930_),
    .Q_N(_14345_),
    .Q(\cpu.ex.r_epc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[11]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1761),
    .D(_00931_),
    .Q_N(_14344_),
    .Q(\cpu.ex.r_epc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[12]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1762),
    .D(_00932_),
    .Q_N(_14343_),
    .Q(\cpu.ex.r_epc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1763),
    .D(_00933_),
    .Q_N(_14342_),
    .Q(\cpu.ex.r_epc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[14]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1764),
    .D(_00934_),
    .Q_N(_14341_),
    .Q(\cpu.ex.r_epc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[1]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1765),
    .D(_00935_),
    .Q_N(_14340_),
    .Q(\cpu.ex.r_epc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[2]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1766),
    .D(_00936_),
    .Q_N(_14339_),
    .Q(\cpu.ex.r_epc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[3]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1767),
    .D(_00937_),
    .Q_N(_14338_),
    .Q(\cpu.ex.r_epc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[4]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1768),
    .D(_00938_),
    .Q_N(_14337_),
    .Q(\cpu.ex.r_epc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[5]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1769),
    .D(_00939_),
    .Q_N(_14336_),
    .Q(\cpu.ex.r_epc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[6]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1770),
    .D(_00940_),
    .Q_N(_14335_),
    .Q(\cpu.ex.r_epc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[7]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1771),
    .D(_00941_),
    .Q_N(_14334_),
    .Q(\cpu.ex.r_epc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[8]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1772),
    .D(_00942_),
    .Q_N(_14333_),
    .Q(\cpu.ex.r_epc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[9]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1773),
    .D(_00943_),
    .Q_N(_14332_),
    .Q(\cpu.ex.r_epc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_fetch$_SDFF_PN1_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1774),
    .D(_00944_),
    .Q_N(_00189_),
    .Q(\cpu.ex.ifetch ));
 sg13g2_dfrbp_1 \cpu.ex.r_flush_write$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1775),
    .D(_00945_),
    .Q_N(_14331_),
    .Q(\cpu.dcache.flush_write ));
 sg13g2_dfrbp_1 \cpu.ex.r_i_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1776),
    .D(_00946_),
    .Q_N(_14330_),
    .Q(\cpu.ex.i_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_ie$_SDFFE_PP0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1777),
    .D(_00947_),
    .Q_N(_14329_),
    .Q(\cpu.ex.r_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_io_access$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1778),
    .D(_00948_),
    .Q_N(_00197_),
    .Q(\cpu.ex.io_access ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[0]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1779),
    .D(_00949_),
    .Q_N(_14328_),
    .Q(\cpu.ex.r_lr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[10]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1780),
    .D(_00950_),
    .Q_N(_14327_),
    .Q(\cpu.ex.r_lr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[11]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1781),
    .D(_00951_),
    .Q_N(_14326_),
    .Q(\cpu.ex.r_lr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[12]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1782),
    .D(_00952_),
    .Q_N(_14325_),
    .Q(\cpu.ex.r_lr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[13]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1783),
    .D(_00953_),
    .Q_N(_14324_),
    .Q(\cpu.ex.r_lr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[14]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1784),
    .D(_00954_),
    .Q_N(_14323_),
    .Q(\cpu.ex.r_lr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[1]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1785),
    .D(_00955_),
    .Q_N(_14322_),
    .Q(\cpu.ex.r_lr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[2]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1786),
    .D(_00956_),
    .Q_N(_14321_),
    .Q(\cpu.ex.r_lr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1787),
    .D(_00957_),
    .Q_N(_14320_),
    .Q(\cpu.ex.r_lr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[4]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1788),
    .D(_00958_),
    .Q_N(_14319_),
    .Q(\cpu.ex.r_lr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[5]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1789),
    .D(_00959_),
    .Q_N(_14318_),
    .Q(\cpu.ex.r_lr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[6]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1790),
    .D(_00960_),
    .Q_N(_14317_),
    .Q(\cpu.ex.r_lr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[7]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1791),
    .D(_00961_),
    .Q_N(_14316_),
    .Q(\cpu.ex.r_lr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[8]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1792),
    .D(_00962_),
    .Q_N(_14315_),
    .Q(\cpu.ex.r_lr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[9]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1793),
    .D(_00963_),
    .Q_N(_14909_),
    .Q(\cpu.ex.r_lr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[0]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1794),
    .D(\cpu.ex.c_mult[0] ),
    .Q_N(_14910_),
    .Q(\cpu.ex.r_mult[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[10]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1795),
    .D(\cpu.ex.c_mult[10] ),
    .Q_N(_00167_),
    .Q(\cpu.ex.r_mult[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[11]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1796),
    .D(\cpu.ex.c_mult[11] ),
    .Q_N(_00168_),
    .Q(\cpu.ex.r_mult[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[12]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1797),
    .D(\cpu.ex.c_mult[12] ),
    .Q_N(_00169_),
    .Q(\cpu.ex.r_mult[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[13]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1798),
    .D(\cpu.ex.c_mult[13] ),
    .Q_N(_00170_),
    .Q(\cpu.ex.r_mult[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[14]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1799),
    .D(\cpu.ex.c_mult[14] ),
    .Q_N(_00171_),
    .Q(\cpu.ex.r_mult[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[15]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1800),
    .D(\cpu.ex.c_mult[15] ),
    .Q_N(_14314_),
    .Q(\cpu.ex.r_mult[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[16]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1801),
    .D(_00964_),
    .Q_N(_00307_),
    .Q(\cpu.ex.r_mult[16] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[17]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1802),
    .D(_00965_),
    .Q_N(_00306_),
    .Q(\cpu.ex.r_mult[17] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[18]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1803),
    .D(_00966_),
    .Q_N(_00305_),
    .Q(\cpu.ex.r_mult[18] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[19]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1804),
    .D(_00967_),
    .Q_N(_00304_),
    .Q(\cpu.ex.r_mult[19] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[1]$_DFF_P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1805),
    .D(\cpu.ex.c_mult[1] ),
    .Q_N(_14313_),
    .Q(\cpu.ex.r_mult[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[20]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1806),
    .D(_00968_),
    .Q_N(_00303_),
    .Q(\cpu.ex.r_mult[20] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[21]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1807),
    .D(_00969_),
    .Q_N(_00302_),
    .Q(\cpu.ex.r_mult[21] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[22]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1808),
    .D(_00970_),
    .Q_N(_14312_),
    .Q(\cpu.ex.r_mult[22] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[23]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1809),
    .D(_00971_),
    .Q_N(_00301_),
    .Q(\cpu.ex.r_mult[23] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[24]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1810),
    .D(_00972_),
    .Q_N(_00300_),
    .Q(\cpu.ex.r_mult[24] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[25]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1811),
    .D(_00973_),
    .Q_N(_00299_),
    .Q(\cpu.ex.r_mult[25] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[26]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1812),
    .D(_00974_),
    .Q_N(_14311_),
    .Q(\cpu.ex.r_mult[26] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[27]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1813),
    .D(_00975_),
    .Q_N(_00298_),
    .Q(\cpu.ex.r_mult[27] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[28]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1814),
    .D(_00976_),
    .Q_N(_14310_),
    .Q(\cpu.ex.r_mult[28] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[29]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1815),
    .D(_00977_),
    .Q_N(_14911_),
    .Q(\cpu.ex.r_mult[29] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[2]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1816),
    .D(\cpu.ex.c_mult[2] ),
    .Q_N(_00120_),
    .Q(\cpu.ex.r_mult[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[30]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1817),
    .D(_00978_),
    .Q_N(_00297_),
    .Q(\cpu.ex.r_mult[30] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[31]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1818),
    .D(_00979_),
    .Q_N(_14912_),
    .Q(\cpu.ex.r_mult[31] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[3]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1819),
    .D(\cpu.ex.c_mult[3] ),
    .Q_N(_00127_),
    .Q(\cpu.ex.r_mult[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[4]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1820),
    .D(\cpu.ex.c_mult[4] ),
    .Q_N(_00139_),
    .Q(\cpu.ex.r_mult[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[5]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1821),
    .D(\cpu.ex.c_mult[5] ),
    .Q_N(_00151_),
    .Q(\cpu.ex.r_mult[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[6]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1822),
    .D(\cpu.ex.c_mult[6] ),
    .Q_N(_00163_),
    .Q(\cpu.ex.r_mult[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[7]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1823),
    .D(\cpu.ex.c_mult[7] ),
    .Q_N(_00164_),
    .Q(\cpu.ex.r_mult[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[8]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1824),
    .D(\cpu.ex.c_mult[8] ),
    .Q_N(_00165_),
    .Q(\cpu.ex.r_mult[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[9]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1825),
    .D(\cpu.ex.c_mult[9] ),
    .Q_N(_00166_),
    .Q(\cpu.ex.r_mult[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[0]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1826),
    .D(\cpu.ex.c_mult_off[0] ),
    .Q_N(_14913_),
    .Q(\cpu.ex.r_mult_off[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[1]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1827),
    .D(\cpu.ex.c_mult_off[1] ),
    .Q_N(_14914_),
    .Q(\cpu.ex.r_mult_off[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[2]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1828),
    .D(\cpu.ex.c_mult_off[2] ),
    .Q_N(_14915_),
    .Q(\cpu.ex.r_mult_off[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[3]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1829),
    .D(\cpu.ex.c_mult_off[3] ),
    .Q_N(_14916_),
    .Q(\cpu.ex.r_mult_off[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_running$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1830),
    .D(\cpu.ex.c_mult_running ),
    .Q_N(_00199_),
    .Q(\cpu.ex.r_mult_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[0]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1831),
    .D(_00980_),
    .Q_N(_00200_),
    .Q(\cpu.ex.pc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[10]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1832),
    .D(_00981_),
    .Q_N(_00288_),
    .Q(\cpu.ex.pc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[11]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1833),
    .D(_00982_),
    .Q_N(_00287_),
    .Q(\cpu.ex.pc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[12]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1834),
    .D(_00983_),
    .Q_N(_00196_),
    .Q(\cpu.ex.pc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[13]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1835),
    .D(_00984_),
    .Q_N(_00195_),
    .Q(\cpu.ex.pc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[14]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1836),
    .D(_00985_),
    .Q_N(_00194_),
    .Q(\cpu.ex.pc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[1]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1837),
    .D(_00986_),
    .Q_N(_00295_),
    .Q(\cpu.ex.pc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[2]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1838),
    .D(_00987_),
    .Q_N(_00191_),
    .Q(\cpu.ex.pc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[3]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1839),
    .D(_00988_),
    .Q_N(_00190_),
    .Q(\cpu.ex.pc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[4]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1840),
    .D(_00989_),
    .Q_N(_00294_),
    .Q(\cpu.ex.pc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[5]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1841),
    .D(_00990_),
    .Q_N(_00293_),
    .Q(\cpu.ex.pc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[6]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1842),
    .D(_00991_),
    .Q_N(_00292_),
    .Q(\cpu.ex.pc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[7]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1843),
    .D(_00992_),
    .Q_N(_00291_),
    .Q(\cpu.ex.pc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[8]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1844),
    .D(_00993_),
    .Q_N(_00290_),
    .Q(\cpu.ex.pc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[9]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1845),
    .D(_00994_),
    .Q_N(_00289_),
    .Q(\cpu.ex.pc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_prev_ie$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1846),
    .D(_00995_),
    .Q_N(_14309_),
    .Q(\cpu.ex.r_prev_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_read_stall$_SDFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1847),
    .D(_00996_),
    .Q_N(_00198_),
    .Q(\cpu.ex.r_read_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_set_cc$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1848),
    .D(_00997_),
    .Q_N(_14308_),
    .Q(\cpu.ex.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[0]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1849),
    .D(_00998_),
    .Q_N(_14307_),
    .Q(\cpu.ex.r_sp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[10]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1850),
    .D(_00999_),
    .Q_N(_14306_),
    .Q(\cpu.ex.r_sp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[11]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1851),
    .D(_01000_),
    .Q_N(_14305_),
    .Q(\cpu.ex.r_sp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[12]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1852),
    .D(_01001_),
    .Q_N(_14304_),
    .Q(\cpu.ex.r_sp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[13]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1853),
    .D(_01002_),
    .Q_N(_14303_),
    .Q(\cpu.ex.r_sp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[14]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1854),
    .D(_01003_),
    .Q_N(_14302_),
    .Q(\cpu.ex.r_sp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[1]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1855),
    .D(_01004_),
    .Q_N(_14301_),
    .Q(\cpu.ex.r_sp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[2]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1856),
    .D(_01005_),
    .Q_N(_14300_),
    .Q(\cpu.ex.r_sp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[3]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1857),
    .D(_01006_),
    .Q_N(_14299_),
    .Q(\cpu.ex.r_sp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[4]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1858),
    .D(_01007_),
    .Q_N(_14298_),
    .Q(\cpu.ex.r_sp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[5]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1859),
    .D(_01008_),
    .Q_N(_14297_),
    .Q(\cpu.ex.r_sp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[6]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1860),
    .D(_01009_),
    .Q_N(_14296_),
    .Q(\cpu.ex.r_sp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[7]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1861),
    .D(_01010_),
    .Q_N(_14295_),
    .Q(\cpu.ex.r_sp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[8]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1862),
    .D(_01011_),
    .Q_N(_14294_),
    .Q(\cpu.ex.r_sp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[9]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1863),
    .D(_01012_),
    .Q_N(_14293_),
    .Q(\cpu.ex.r_sp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1864),
    .D(_01013_),
    .Q_N(_14292_),
    .Q(\cpu.ex.r_stmp[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1865),
    .D(_01014_),
    .Q_N(_14291_),
    .Q(\cpu.ex.r_stmp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1866),
    .D(_01015_),
    .Q_N(_14290_),
    .Q(\cpu.ex.r_stmp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1867),
    .D(_01016_),
    .Q_N(_14289_),
    .Q(\cpu.ex.r_stmp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1868),
    .D(_01017_),
    .Q_N(_14288_),
    .Q(\cpu.ex.r_stmp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1869),
    .D(_01018_),
    .Q_N(_14287_),
    .Q(\cpu.ex.r_stmp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1870),
    .D(_01019_),
    .Q_N(_14286_),
    .Q(\cpu.ex.r_stmp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1871),
    .D(_01020_),
    .Q_N(_14285_),
    .Q(\cpu.ex.r_stmp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1872),
    .D(_01021_),
    .Q_N(_14284_),
    .Q(\cpu.ex.r_stmp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1873),
    .D(_01022_),
    .Q_N(_14283_),
    .Q(\cpu.ex.r_stmp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1874),
    .D(_01023_),
    .Q_N(_14282_),
    .Q(\cpu.ex.r_stmp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1875),
    .D(_01024_),
    .Q_N(_14281_),
    .Q(\cpu.ex.r_stmp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1876),
    .D(_01025_),
    .Q_N(_14280_),
    .Q(\cpu.ex.r_stmp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1877),
    .D(_01026_),
    .Q_N(_14279_),
    .Q(\cpu.ex.r_stmp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1878),
    .D(_01027_),
    .Q_N(_14278_),
    .Q(\cpu.ex.r_stmp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1879),
    .D(_01028_),
    .Q_N(_14277_),
    .Q(\cpu.ex.r_stmp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[0]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1880),
    .D(_01029_),
    .Q_N(_00255_),
    .Q(\cpu.ex.mmu_reg_data[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1881),
    .D(_01030_),
    .Q_N(_00237_),
    .Q(\cpu.addr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[11]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1882),
    .D(_01031_),
    .Q_N(_00239_),
    .Q(\cpu.addr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[12]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1883),
    .D(_01032_),
    .Q_N(_14276_),
    .Q(\cpu.addr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[13]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1884),
    .D(_01033_),
    .Q_N(_14275_),
    .Q(\cpu.addr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[14]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1885),
    .D(_01034_),
    .Q_N(_14274_),
    .Q(\cpu.addr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[15]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1886),
    .D(_01035_),
    .Q_N(_14273_),
    .Q(\cpu.addr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1887),
    .D(_01036_),
    .Q_N(_00273_),
    .Q(\cpu.addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[2]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1888),
    .D(_01037_),
    .Q_N(_14272_),
    .Q(\cpu.addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[3]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1889),
    .D(_01038_),
    .Q_N(_00226_),
    .Q(\cpu.addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[4]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1890),
    .D(_01039_),
    .Q_N(_00225_),
    .Q(\cpu.addr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[5]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1891),
    .D(_01040_),
    .Q_N(_00227_),
    .Q(\cpu.addr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[6]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1892),
    .D(_01041_),
    .Q_N(_00229_),
    .Q(\cpu.addr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[7]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1893),
    .D(_01042_),
    .Q_N(_00231_),
    .Q(\cpu.addr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[8]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1894),
    .D(_01043_),
    .Q_N(_00233_),
    .Q(\cpu.addr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[9]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1895),
    .D(_01044_),
    .Q_N(_00235_),
    .Q(\cpu.addr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1896),
    .D(_01045_),
    .Q_N(_14271_),
    .Q(\cpu.ex.r_wb_addr[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1897),
    .D(_01046_),
    .Q_N(_14270_),
    .Q(\cpu.ex.r_wb_addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1898),
    .D(_01047_),
    .Q_N(_14269_),
    .Q(\cpu.ex.r_wb_addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1899),
    .D(_01048_),
    .Q_N(_14268_),
    .Q(\cpu.ex.r_wb_addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1900),
    .D(_01049_),
    .Q_N(_14917_),
    .Q(\cpu.ex.r_wb_swapsp ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_valid$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1901),
    .D(_00054_),
    .Q_N(_00254_),
    .Q(\cpu.ex.r_wb_valid ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[0]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1902),
    .D(_01050_),
    .Q_N(_00221_),
    .Q(\cpu.dcache.wdata[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[10]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1903),
    .D(_01051_),
    .Q_N(_14267_),
    .Q(\cpu.dcache.wdata[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1904),
    .D(_01052_),
    .Q_N(_14266_),
    .Q(\cpu.dcache.wdata[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[12]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1905),
    .D(_01053_),
    .Q_N(_14265_),
    .Q(\cpu.dcache.wdata[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[13]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1906),
    .D(_01054_),
    .Q_N(_14264_),
    .Q(\cpu.dcache.wdata[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[14]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1907),
    .D(_01055_),
    .Q_N(_14263_),
    .Q(\cpu.dcache.wdata[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[15]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1908),
    .D(_01056_),
    .Q_N(_14262_),
    .Q(\cpu.dcache.wdata[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[1]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1909),
    .D(_01057_),
    .Q_N(_00181_),
    .Q(\cpu.dcache.wdata[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1910),
    .D(_01058_),
    .Q_N(_00182_),
    .Q(\cpu.dcache.wdata[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[3]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1911),
    .D(_01059_),
    .Q_N(_00285_),
    .Q(\cpu.dcache.wdata[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[4]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1912),
    .D(_01060_),
    .Q_N(_00183_),
    .Q(\cpu.dcache.wdata[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[5]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1913),
    .D(_01061_),
    .Q_N(_00184_),
    .Q(\cpu.dcache.wdata[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1914),
    .D(_01062_),
    .Q_N(_00185_),
    .Q(\cpu.dcache.wdata[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[7]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1915),
    .D(_01063_),
    .Q_N(_00279_),
    .Q(\cpu.dcache.wdata[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[8]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1916),
    .D(_01064_),
    .Q_N(_14261_),
    .Q(\cpu.dcache.wdata[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[9]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1917),
    .D(_01065_),
    .Q_N(_14260_),
    .Q(\cpu.dcache.wdata[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1918),
    .D(_01066_),
    .Q_N(_14259_),
    .Q(\cpu.ex.r_wmask[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1919),
    .D(_01067_),
    .Q_N(_14258_),
    .Q(\cpu.ex.r_wmask[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1920),
    .D(_01068_),
    .Q_N(_00286_),
    .Q(\cpu.ex.mmu_read[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1921),
    .D(_01069_),
    .Q_N(_14257_),
    .Q(\cpu.ex.mmu_read[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1922),
    .D(_01070_),
    .Q_N(_00188_),
    .Q(\cpu.ex.mmu_read[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1923),
    .D(_01071_),
    .Q_N(_14256_),
    .Q(\cpu.ex.mmu_read[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1924),
    .D(_01072_),
    .Q_N(_00253_),
    .Q(\cpu.ex.mmu_read[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1925),
    .D(_01073_),
    .Q_N(_14255_),
    .Q(\cpu.ex.mmu_read[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1926),
    .D(_01074_),
    .Q_N(_14254_),
    .Q(\cpu.ex.mmu_read[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1927),
    .D(_01075_),
    .Q_N(_14253_),
    .Q(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1928),
    .D(_01076_),
    .Q_N(_14252_),
    .Q(\cpu.genblk1.mmu.r_valid_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1929),
    .D(_01077_),
    .Q_N(_14251_),
    .Q(\cpu.genblk1.mmu.r_valid_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1930),
    .D(_01078_),
    .Q_N(_14250_),
    .Q(\cpu.genblk1.mmu.r_valid_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1931),
    .D(_01079_),
    .Q_N(_14249_),
    .Q(\cpu.genblk1.mmu.r_valid_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1932),
    .D(_01080_),
    .Q_N(_14248_),
    .Q(\cpu.genblk1.mmu.r_valid_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1933),
    .D(_01081_),
    .Q_N(_14247_),
    .Q(\cpu.genblk1.mmu.r_valid_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1934),
    .D(_01082_),
    .Q_N(_14246_),
    .Q(\cpu.genblk1.mmu.r_valid_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1935),
    .D(_01083_),
    .Q_N(_14245_),
    .Q(\cpu.genblk1.mmu.r_valid_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1936),
    .D(_01084_),
    .Q_N(_14244_),
    .Q(\cpu.genblk1.mmu.r_valid_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1937),
    .D(_01085_),
    .Q_N(_14243_),
    .Q(\cpu.genblk1.mmu.r_valid_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1938),
    .D(_01086_),
    .Q_N(_14242_),
    .Q(\cpu.genblk1.mmu.r_valid_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1939),
    .D(_01087_),
    .Q_N(_14241_),
    .Q(\cpu.genblk1.mmu.r_valid_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1940),
    .D(_01088_),
    .Q_N(_14240_),
    .Q(\cpu.genblk1.mmu.r_valid_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1941),
    .D(_01089_),
    .Q_N(_14239_),
    .Q(\cpu.genblk1.mmu.r_valid_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1942),
    .D(_01090_),
    .Q_N(_14238_),
    .Q(\cpu.genblk1.mmu.r_valid_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1943),
    .D(_01091_),
    .Q_N(_14237_),
    .Q(\cpu.genblk1.mmu.r_valid_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1944),
    .D(_01092_),
    .Q_N(_14236_),
    .Q(\cpu.genblk1.mmu.r_valid_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1945),
    .D(_01093_),
    .Q_N(_14235_),
    .Q(\cpu.genblk1.mmu.r_valid_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1946),
    .D(_01094_),
    .Q_N(_14234_),
    .Q(\cpu.genblk1.mmu.r_valid_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1947),
    .D(_01095_),
    .Q_N(_14233_),
    .Q(\cpu.genblk1.mmu.r_valid_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1948),
    .D(_01096_),
    .Q_N(_14232_),
    .Q(\cpu.genblk1.mmu.r_valid_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1949),
    .D(_01097_),
    .Q_N(_14231_),
    .Q(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1950),
    .D(_01098_),
    .Q_N(_14230_),
    .Q(\cpu.genblk1.mmu.r_valid_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1951),
    .D(_01099_),
    .Q_N(_14229_),
    .Q(\cpu.genblk1.mmu.r_valid_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1952),
    .D(_01100_),
    .Q_N(_14228_),
    .Q(\cpu.genblk1.mmu.r_valid_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1953),
    .D(_01101_),
    .Q_N(_14227_),
    .Q(\cpu.genblk1.mmu.r_valid_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1954),
    .D(_01102_),
    .Q_N(_14226_),
    .Q(\cpu.genblk1.mmu.r_valid_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1955),
    .D(_01103_),
    .Q_N(_14225_),
    .Q(\cpu.genblk1.mmu.r_valid_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1956),
    .D(_01104_),
    .Q_N(_14224_),
    .Q(\cpu.genblk1.mmu.r_valid_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1957),
    .D(_01105_),
    .Q_N(_14223_),
    .Q(\cpu.genblk1.mmu.r_valid_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1958),
    .D(_01106_),
    .Q_N(_14222_),
    .Q(\cpu.genblk1.mmu.r_valid_d[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1959),
    .D(_01107_),
    .Q_N(_14221_),
    .Q(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1960),
    .D(_01108_),
    .Q_N(_14220_),
    .Q(\cpu.genblk1.mmu.r_valid_i[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1961),
    .D(_01109_),
    .Q_N(_14219_),
    .Q(\cpu.genblk1.mmu.r_valid_i[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1962),
    .D(_01110_),
    .Q_N(_14218_),
    .Q(\cpu.genblk1.mmu.r_valid_i[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1963),
    .D(_01111_),
    .Q_N(_14217_),
    .Q(\cpu.genblk1.mmu.r_valid_i[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1964),
    .D(_01112_),
    .Q_N(_14216_),
    .Q(\cpu.genblk1.mmu.r_valid_i[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1965),
    .D(_01113_),
    .Q_N(_14215_),
    .Q(\cpu.genblk1.mmu.r_valid_i[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1966),
    .D(_01114_),
    .Q_N(_14214_),
    .Q(\cpu.genblk1.mmu.r_valid_i[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1967),
    .D(_01115_),
    .Q_N(_14213_),
    .Q(\cpu.genblk1.mmu.r_valid_i[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1968),
    .D(_01116_),
    .Q_N(_14212_),
    .Q(\cpu.genblk1.mmu.r_valid_i[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1969),
    .D(_01117_),
    .Q_N(_14211_),
    .Q(\cpu.genblk1.mmu.r_valid_i[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1970),
    .D(_01118_),
    .Q_N(_14210_),
    .Q(\cpu.genblk1.mmu.r_valid_i[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1971),
    .D(_01119_),
    .Q_N(_14209_),
    .Q(\cpu.genblk1.mmu.r_valid_i[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1972),
    .D(_01120_),
    .Q_N(_14208_),
    .Q(\cpu.genblk1.mmu.r_valid_i[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1973),
    .D(_01121_),
    .Q_N(_14207_),
    .Q(\cpu.genblk1.mmu.r_valid_i[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1974),
    .D(_01122_),
    .Q_N(_14206_),
    .Q(\cpu.genblk1.mmu.r_valid_i[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1975),
    .D(_01123_),
    .Q_N(_14205_),
    .Q(\cpu.genblk1.mmu.r_valid_i[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1976),
    .D(_01124_),
    .Q_N(_14204_),
    .Q(\cpu.genblk1.mmu.r_valid_i[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1977),
    .D(_01125_),
    .Q_N(_14203_),
    .Q(\cpu.genblk1.mmu.r_valid_i[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1978),
    .D(_01126_),
    .Q_N(_14202_),
    .Q(\cpu.genblk1.mmu.r_valid_i[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1979),
    .D(_01127_),
    .Q_N(_14201_),
    .Q(\cpu.genblk1.mmu.r_valid_i[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1980),
    .D(_01128_),
    .Q_N(_14200_),
    .Q(\cpu.genblk1.mmu.r_valid_i[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1981),
    .D(_01129_),
    .Q_N(_14199_),
    .Q(\cpu.genblk1.mmu.r_valid_i[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1982),
    .D(_01130_),
    .Q_N(_14198_),
    .Q(\cpu.genblk1.mmu.r_valid_i[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1983),
    .D(_01131_),
    .Q_N(_14197_),
    .Q(\cpu.genblk1.mmu.r_valid_i[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1984),
    .D(_01132_),
    .Q_N(_14196_),
    .Q(\cpu.genblk1.mmu.r_valid_i[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1985),
    .D(_01133_),
    .Q_N(_14195_),
    .Q(\cpu.genblk1.mmu.r_valid_i[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1986),
    .D(_01134_),
    .Q_N(_14194_),
    .Q(\cpu.genblk1.mmu.r_valid_i[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1987),
    .D(_01135_),
    .Q_N(_14193_),
    .Q(\cpu.genblk1.mmu.r_valid_i[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1988),
    .D(_01136_),
    .Q_N(_14192_),
    .Q(\cpu.genblk1.mmu.r_valid_i[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1989),
    .D(_01137_),
    .Q_N(_14191_),
    .Q(\cpu.genblk1.mmu.r_valid_i[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1990),
    .D(_01138_),
    .Q_N(_14190_),
    .Q(\cpu.genblk1.mmu.r_valid_i[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1991),
    .D(_01139_),
    .Q_N(_14189_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1992),
    .D(_01140_),
    .Q_N(_14188_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1993),
    .D(_01141_),
    .Q_N(_14187_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1994),
    .D(_01142_),
    .Q_N(_14186_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1995),
    .D(_01143_),
    .Q_N(_14185_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1996),
    .D(_01144_),
    .Q_N(_14184_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1997),
    .D(_01145_),
    .Q_N(_14183_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1998),
    .D(_01146_),
    .Q_N(_14182_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1999),
    .D(_01147_),
    .Q_N(_14181_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2000),
    .D(_01148_),
    .Q_N(_14180_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2001),
    .D(_01149_),
    .Q_N(_14179_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2002),
    .D(_01150_),
    .Q_N(_14178_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2003),
    .D(_01151_),
    .Q_N(_14177_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2004),
    .D(_01152_),
    .Q_N(_14176_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2005),
    .D(_01153_),
    .Q_N(_14175_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2006),
    .D(_01154_),
    .Q_N(_14174_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2007),
    .D(_01155_),
    .Q_N(_14173_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2008),
    .D(_01156_),
    .Q_N(_14172_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2009),
    .D(_01157_),
    .Q_N(_14171_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2010),
    .D(_01158_),
    .Q_N(_14170_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2011),
    .D(_01159_),
    .Q_N(_14169_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2012),
    .D(_01160_),
    .Q_N(_14168_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2013),
    .D(_01161_),
    .Q_N(_14167_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2014),
    .D(_01162_),
    .Q_N(_14166_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2015),
    .D(_01163_),
    .Q_N(_14165_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2016),
    .D(_01164_),
    .Q_N(_14164_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2017),
    .D(_01165_),
    .Q_N(_14163_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2018),
    .D(_01166_),
    .Q_N(_14162_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2019),
    .D(_01167_),
    .Q_N(_14161_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2020),
    .D(_01168_),
    .Q_N(_14160_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2021),
    .D(_01169_),
    .Q_N(_14159_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2022),
    .D(_01170_),
    .Q_N(_14158_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2023),
    .D(_01171_),
    .Q_N(_14157_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2024),
    .D(_01172_),
    .Q_N(_14156_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2025),
    .D(_01173_),
    .Q_N(_14155_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2026),
    .D(_01174_),
    .Q_N(_14154_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2027),
    .D(_01175_),
    .Q_N(_14153_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2028),
    .D(_01176_),
    .Q_N(_14152_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2029),
    .D(_01177_),
    .Q_N(_14151_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2030),
    .D(_01178_),
    .Q_N(_14150_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2031),
    .D(_01179_),
    .Q_N(_14149_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2032),
    .D(_01180_),
    .Q_N(_14148_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2033),
    .D(_01181_),
    .Q_N(_14147_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2034),
    .D(_01182_),
    .Q_N(_14146_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2035),
    .D(_01183_),
    .Q_N(_14145_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2036),
    .D(_01184_),
    .Q_N(_14144_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2037),
    .D(_01185_),
    .Q_N(_14143_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2038),
    .D(_01186_),
    .Q_N(_14142_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2039),
    .D(_01187_),
    .Q_N(_14141_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2040),
    .D(_01188_),
    .Q_N(_14140_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2041),
    .D(_01189_),
    .Q_N(_14139_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2042),
    .D(_01190_),
    .Q_N(_14138_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2043),
    .D(_01191_),
    .Q_N(_14137_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2044),
    .D(_01192_),
    .Q_N(_14136_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2045),
    .D(_01193_),
    .Q_N(_14135_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2046),
    .D(_01194_),
    .Q_N(_14134_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2047),
    .D(_01195_),
    .Q_N(_14133_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2048),
    .D(_01196_),
    .Q_N(_14132_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2049),
    .D(_01197_),
    .Q_N(_14131_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2050),
    .D(_01198_),
    .Q_N(_14130_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2051),
    .D(_01199_),
    .Q_N(_14129_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2052),
    .D(_01200_),
    .Q_N(_14128_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2053),
    .D(_01201_),
    .Q_N(_14127_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2054),
    .D(_01202_),
    .Q_N(_14126_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2055),
    .D(_01203_),
    .Q_N(_14125_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2056),
    .D(_01204_),
    .Q_N(_14124_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2057),
    .D(_01205_),
    .Q_N(_14123_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2058),
    .D(_01206_),
    .Q_N(_14122_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2059),
    .D(_01207_),
    .Q_N(_14121_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2060),
    .D(_01208_),
    .Q_N(_14120_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2061),
    .D(_01209_),
    .Q_N(_14119_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2062),
    .D(_01210_),
    .Q_N(_14118_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2063),
    .D(_01211_),
    .Q_N(_14117_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2064),
    .D(_01212_),
    .Q_N(_14116_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2065),
    .D(_01213_),
    .Q_N(_14115_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2066),
    .D(_01214_),
    .Q_N(_14114_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2067),
    .D(_01215_),
    .Q_N(_14113_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2068),
    .D(_01216_),
    .Q_N(_14112_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2069),
    .D(_01217_),
    .Q_N(_14111_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2070),
    .D(_01218_),
    .Q_N(_14110_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2071),
    .D(_01219_),
    .Q_N(_14109_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2072),
    .D(_01220_),
    .Q_N(_14108_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2073),
    .D(_01221_),
    .Q_N(_14107_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2074),
    .D(_01222_),
    .Q_N(_14106_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2075),
    .D(_01223_),
    .Q_N(_14105_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2076),
    .D(_01224_),
    .Q_N(_14104_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2077),
    .D(_01225_),
    .Q_N(_14103_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2078),
    .D(_01226_),
    .Q_N(_14102_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2079),
    .D(_01227_),
    .Q_N(_14101_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2080),
    .D(_01228_),
    .Q_N(_14100_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2081),
    .D(_01229_),
    .Q_N(_14099_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2082),
    .D(_01230_),
    .Q_N(_14098_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2083),
    .D(_01231_),
    .Q_N(_14097_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2084),
    .D(_01232_),
    .Q_N(_14096_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2085),
    .D(_01233_),
    .Q_N(_14095_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2086),
    .D(_01234_),
    .Q_N(_14094_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2087),
    .D(_01235_),
    .Q_N(_14093_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2088),
    .D(_01236_),
    .Q_N(_14092_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2089),
    .D(_01237_),
    .Q_N(_14091_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2090),
    .D(_01238_),
    .Q_N(_14090_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2091),
    .D(_01239_),
    .Q_N(_14089_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2092),
    .D(_01240_),
    .Q_N(_14088_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2093),
    .D(_01241_),
    .Q_N(_14087_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2094),
    .D(_01242_),
    .Q_N(_14086_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2095),
    .D(_01243_),
    .Q_N(_14085_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2096),
    .D(_01244_),
    .Q_N(_14084_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2097),
    .D(_01245_),
    .Q_N(_14083_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2098),
    .D(_01246_),
    .Q_N(_14082_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2099),
    .D(_01247_),
    .Q_N(_14081_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2100),
    .D(_01248_),
    .Q_N(_14080_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2101),
    .D(_01249_),
    .Q_N(_14079_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2102),
    .D(_01250_),
    .Q_N(_14078_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2103),
    .D(_01251_),
    .Q_N(_14077_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2104),
    .D(_01252_),
    .Q_N(_14076_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2105),
    .D(_01253_),
    .Q_N(_14075_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2106),
    .D(_01254_),
    .Q_N(_14074_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2107),
    .D(_01255_),
    .Q_N(_14073_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2108),
    .D(_01256_),
    .Q_N(_14072_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2109),
    .D(_01257_),
    .Q_N(_14071_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2110),
    .D(_01258_),
    .Q_N(_14070_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2111),
    .D(_01259_),
    .Q_N(_14069_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2112),
    .D(_01260_),
    .Q_N(_14068_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2113),
    .D(_01261_),
    .Q_N(_14067_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2114),
    .D(_01262_),
    .Q_N(_14066_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2115),
    .D(_01263_),
    .Q_N(_14065_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2116),
    .D(_01264_),
    .Q_N(_14064_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2117),
    .D(_01265_),
    .Q_N(_14063_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2118),
    .D(_01266_),
    .Q_N(_14062_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2119),
    .D(_01267_),
    .Q_N(_14061_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2120),
    .D(_01268_),
    .Q_N(_14060_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2121),
    .D(_01269_),
    .Q_N(_14059_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2122),
    .D(_01270_),
    .Q_N(_14058_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2123),
    .D(_01271_),
    .Q_N(_14057_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2124),
    .D(_01272_),
    .Q_N(_14056_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2125),
    .D(_01273_),
    .Q_N(_14055_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2126),
    .D(_01274_),
    .Q_N(_14054_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2127),
    .D(_01275_),
    .Q_N(_14053_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2128),
    .D(_01276_),
    .Q_N(_14052_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2129),
    .D(_01277_),
    .Q_N(_14051_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2130),
    .D(_01278_),
    .Q_N(_14050_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2131),
    .D(_01279_),
    .Q_N(_14049_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2132),
    .D(_01280_),
    .Q_N(_14048_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2133),
    .D(_01281_),
    .Q_N(_14047_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2134),
    .D(_01282_),
    .Q_N(_14046_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2135),
    .D(_01283_),
    .Q_N(_14045_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2136),
    .D(_01284_),
    .Q_N(_14044_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2137),
    .D(_01285_),
    .Q_N(_14043_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2138),
    .D(_01286_),
    .Q_N(_14042_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2139),
    .D(_01287_),
    .Q_N(_14041_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2140),
    .D(_01288_),
    .Q_N(_14040_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2141),
    .D(_01289_),
    .Q_N(_14039_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2142),
    .D(_01290_),
    .Q_N(_14038_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2143),
    .D(_01291_),
    .Q_N(_14037_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2144),
    .D(_01292_),
    .Q_N(_14036_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2145),
    .D(_01293_),
    .Q_N(_14035_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2146),
    .D(_01294_),
    .Q_N(_14034_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2147),
    .D(_01295_),
    .Q_N(_14033_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2148),
    .D(_01296_),
    .Q_N(_14032_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2149),
    .D(_01297_),
    .Q_N(_14031_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2150),
    .D(_01298_),
    .Q_N(_14030_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2151),
    .D(_01299_),
    .Q_N(_14029_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2152),
    .D(_01300_),
    .Q_N(_14028_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2153),
    .D(_01301_),
    .Q_N(_14027_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2154),
    .D(_01302_),
    .Q_N(_14026_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2155),
    .D(_01303_),
    .Q_N(_14025_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2156),
    .D(_01304_),
    .Q_N(_14024_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2157),
    .D(_01305_),
    .Q_N(_14023_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2158),
    .D(_01306_),
    .Q_N(_14022_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2159),
    .D(_01307_),
    .Q_N(_14021_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2160),
    .D(_01308_),
    .Q_N(_14020_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2161),
    .D(_01309_),
    .Q_N(_14019_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2162),
    .D(_01310_),
    .Q_N(_14018_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2163),
    .D(_01311_),
    .Q_N(_14017_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2164),
    .D(_01312_),
    .Q_N(_14016_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2165),
    .D(_01313_),
    .Q_N(_14015_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2166),
    .D(_01314_),
    .Q_N(_14014_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2167),
    .D(_01315_),
    .Q_N(_14013_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2168),
    .D(_01316_),
    .Q_N(_14012_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2169),
    .D(_01317_),
    .Q_N(_14011_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2170),
    .D(_01318_),
    .Q_N(_14010_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2171),
    .D(_01319_),
    .Q_N(_14009_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2172),
    .D(_01320_),
    .Q_N(_14008_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2173),
    .D(_01321_),
    .Q_N(_14007_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2174),
    .D(_01322_),
    .Q_N(_14006_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2175),
    .D(_01323_),
    .Q_N(_14005_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2176),
    .D(_01324_),
    .Q_N(_14004_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2177),
    .D(_01325_),
    .Q_N(_14003_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2178),
    .D(_01326_),
    .Q_N(_14002_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2179),
    .D(_01327_),
    .Q_N(_14001_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2180),
    .D(_01328_),
    .Q_N(_14000_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2181),
    .D(_01329_),
    .Q_N(_13999_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2182),
    .D(_01330_),
    .Q_N(_13998_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2183),
    .D(_01331_),
    .Q_N(_13997_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2184),
    .D(_01332_),
    .Q_N(_13996_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2185),
    .D(_01333_),
    .Q_N(_13995_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2186),
    .D(_01334_),
    .Q_N(_13994_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2187),
    .D(_01335_),
    .Q_N(_13993_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2188),
    .D(_01336_),
    .Q_N(_13992_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2189),
    .D(_01337_),
    .Q_N(_13991_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2190),
    .D(_01338_),
    .Q_N(_13990_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2191),
    .D(_01339_),
    .Q_N(_13989_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2192),
    .D(_01340_),
    .Q_N(_13988_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2193),
    .D(_01341_),
    .Q_N(_13987_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2194),
    .D(_01342_),
    .Q_N(_13986_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2195),
    .D(_01343_),
    .Q_N(_13985_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2196),
    .D(_01344_),
    .Q_N(_13984_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2197),
    .D(_01345_),
    .Q_N(_13983_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2198),
    .D(_01346_),
    .Q_N(_13982_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2199),
    .D(_01347_),
    .Q_N(_13981_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2200),
    .D(_01348_),
    .Q_N(_13980_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2201),
    .D(_01349_),
    .Q_N(_13979_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2202),
    .D(_01350_),
    .Q_N(_13978_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2203),
    .D(_01351_),
    .Q_N(_13977_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2204),
    .D(_01352_),
    .Q_N(_13976_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2205),
    .D(_01353_),
    .Q_N(_13975_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2206),
    .D(_01354_),
    .Q_N(_13974_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2207),
    .D(_01355_),
    .Q_N(_13973_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2208),
    .D(_01356_),
    .Q_N(_13972_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2209),
    .D(_01357_),
    .Q_N(_13971_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2210),
    .D(_01358_),
    .Q_N(_13970_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2211),
    .D(_01359_),
    .Q_N(_13969_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2212),
    .D(_01360_),
    .Q_N(_13968_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2213),
    .D(_01361_),
    .Q_N(_13967_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2214),
    .D(_01362_),
    .Q_N(_13966_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2215),
    .D(_01363_),
    .Q_N(_13965_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2216),
    .D(_01364_),
    .Q_N(_13964_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2217),
    .D(_01365_),
    .Q_N(_13963_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2218),
    .D(_01366_),
    .Q_N(_13962_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2219),
    .D(_01367_),
    .Q_N(_13961_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2220),
    .D(_01368_),
    .Q_N(_13960_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2221),
    .D(_01369_),
    .Q_N(_13959_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2222),
    .D(_01370_),
    .Q_N(_13958_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2223),
    .D(_01371_),
    .Q_N(_13957_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2224),
    .D(_01372_),
    .Q_N(_13956_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2225),
    .D(_01373_),
    .Q_N(_13955_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2226),
    .D(_01374_),
    .Q_N(_13954_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2227),
    .D(_01375_),
    .Q_N(_13953_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2228),
    .D(_01376_),
    .Q_N(_13952_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2229),
    .D(_01377_),
    .Q_N(_13951_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2230),
    .D(_01378_),
    .Q_N(_13950_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2231),
    .D(_01379_),
    .Q_N(_13949_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2232),
    .D(_01380_),
    .Q_N(_13948_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2233),
    .D(_01381_),
    .Q_N(_13947_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2234),
    .D(_01382_),
    .Q_N(_13946_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2235),
    .D(_01383_),
    .Q_N(_13945_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2236),
    .D(_01384_),
    .Q_N(_13944_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2237),
    .D(_01385_),
    .Q_N(_13943_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2238),
    .D(_01386_),
    .Q_N(_13942_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2239),
    .D(_01387_),
    .Q_N(_13941_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2240),
    .D(_01388_),
    .Q_N(_13940_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2241),
    .D(_01389_),
    .Q_N(_13939_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2242),
    .D(_01390_),
    .Q_N(_13938_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2243),
    .D(_01391_),
    .Q_N(_13937_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2244),
    .D(_01392_),
    .Q_N(_13936_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2245),
    .D(_01393_),
    .Q_N(_13935_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2246),
    .D(_01394_),
    .Q_N(_13934_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2247),
    .D(_01395_),
    .Q_N(_13933_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2248),
    .D(_01396_),
    .Q_N(_13932_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2249),
    .D(_01397_),
    .Q_N(_13931_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2250),
    .D(_01398_),
    .Q_N(_13930_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2251),
    .D(_01399_),
    .Q_N(_13929_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2252),
    .D(_01400_),
    .Q_N(_13928_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2253),
    .D(_01401_),
    .Q_N(_13927_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2254),
    .D(_01402_),
    .Q_N(_13926_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2255),
    .D(_01403_),
    .Q_N(_13925_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2256),
    .D(_01404_),
    .Q_N(_13924_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2257),
    .D(_01405_),
    .Q_N(_13923_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2258),
    .D(_01406_),
    .Q_N(_13922_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2259),
    .D(_01407_),
    .Q_N(_13921_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2260),
    .D(_01408_),
    .Q_N(_13920_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2261),
    .D(_01409_),
    .Q_N(_13919_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2262),
    .D(_01410_),
    .Q_N(_13918_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2263),
    .D(_01411_),
    .Q_N(_13917_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2264),
    .D(_01412_),
    .Q_N(_13916_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2265),
    .D(_01413_),
    .Q_N(_13915_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2266),
    .D(_01414_),
    .Q_N(_13914_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2267),
    .D(_01415_),
    .Q_N(_13913_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2268),
    .D(_01416_),
    .Q_N(_13912_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2269),
    .D(_01417_),
    .Q_N(_13911_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2270),
    .D(_01418_),
    .Q_N(_13910_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2271),
    .D(_01419_),
    .Q_N(_13909_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2272),
    .D(_01420_),
    .Q_N(_13908_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2273),
    .D(_01421_),
    .Q_N(_13907_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2274),
    .D(_01422_),
    .Q_N(_13906_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2275),
    .D(_01423_),
    .Q_N(_13905_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2276),
    .D(_01424_),
    .Q_N(_13904_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2277),
    .D(_01425_),
    .Q_N(_13903_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2278),
    .D(_01426_),
    .Q_N(_13902_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2279),
    .D(_01427_),
    .Q_N(_13901_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2280),
    .D(_01428_),
    .Q_N(_13900_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2281),
    .D(_01429_),
    .Q_N(_13899_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2282),
    .D(_01430_),
    .Q_N(_13898_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2283),
    .D(_01431_),
    .Q_N(_13897_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2284),
    .D(_01432_),
    .Q_N(_13896_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2285),
    .D(_01433_),
    .Q_N(_13895_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2286),
    .D(_01434_),
    .Q_N(_13894_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2287),
    .D(_01435_),
    .Q_N(_13893_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2288),
    .D(_01436_),
    .Q_N(_13892_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2289),
    .D(_01437_),
    .Q_N(_13891_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2290),
    .D(_01438_),
    .Q_N(_13890_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2291),
    .D(_01439_),
    .Q_N(_13889_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2292),
    .D(_01440_),
    .Q_N(_13888_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2293),
    .D(_01441_),
    .Q_N(_13887_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2294),
    .D(_01442_),
    .Q_N(_13886_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2295),
    .D(_01443_),
    .Q_N(_13885_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2296),
    .D(_01444_),
    .Q_N(_13884_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2297),
    .D(_01445_),
    .Q_N(_13883_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2298),
    .D(_01446_),
    .Q_N(_13882_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2299),
    .D(_01447_),
    .Q_N(_13881_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2300),
    .D(_01448_),
    .Q_N(_13880_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2301),
    .D(_01449_),
    .Q_N(_13879_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2302),
    .D(_01450_),
    .Q_N(_13878_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2303),
    .D(_01451_),
    .Q_N(_13877_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2304),
    .D(_01452_),
    .Q_N(_13876_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2305),
    .D(_01453_),
    .Q_N(_13875_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2306),
    .D(_01454_),
    .Q_N(_13874_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2307),
    .D(_01455_),
    .Q_N(_13873_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2308),
    .D(_01456_),
    .Q_N(_13872_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2309),
    .D(_01457_),
    .Q_N(_13871_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2310),
    .D(_01458_),
    .Q_N(_13870_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2311),
    .D(_01459_),
    .Q_N(_13869_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2312),
    .D(_01460_),
    .Q_N(_13868_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2313),
    .D(_01461_),
    .Q_N(_13867_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2314),
    .D(_01462_),
    .Q_N(_13866_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2315),
    .D(_01463_),
    .Q_N(_13865_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2316),
    .D(_01464_),
    .Q_N(_13864_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2317),
    .D(_01465_),
    .Q_N(_13863_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2318),
    .D(_01466_),
    .Q_N(_13862_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2319),
    .D(_01467_),
    .Q_N(_13861_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2320),
    .D(_01468_),
    .Q_N(_13860_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2321),
    .D(_01469_),
    .Q_N(_13859_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2322),
    .D(_01470_),
    .Q_N(_13858_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2323),
    .D(_01471_),
    .Q_N(_13857_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2324),
    .D(_01472_),
    .Q_N(_13856_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2325),
    .D(_01473_),
    .Q_N(_13855_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2326),
    .D(_01474_),
    .Q_N(_13854_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2327),
    .D(_01475_),
    .Q_N(_13853_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2328),
    .D(_01476_),
    .Q_N(_13852_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2329),
    .D(_01477_),
    .Q_N(_13851_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2330),
    .D(_01478_),
    .Q_N(_13850_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2331),
    .D(_01479_),
    .Q_N(_13849_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2332),
    .D(_01480_),
    .Q_N(_13848_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2333),
    .D(_01481_),
    .Q_N(_13847_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2334),
    .D(_01482_),
    .Q_N(_13846_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2335),
    .D(_01483_),
    .Q_N(_13845_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2336),
    .D(_01484_),
    .Q_N(_13844_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2337),
    .D(_01485_),
    .Q_N(_13843_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2338),
    .D(_01486_),
    .Q_N(_13842_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2339),
    .D(_01487_),
    .Q_N(_13841_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2340),
    .D(_01488_),
    .Q_N(_13840_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2341),
    .D(_01489_),
    .Q_N(_13839_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2342),
    .D(_01490_),
    .Q_N(_13838_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2343),
    .D(_01491_),
    .Q_N(_13837_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2344),
    .D(_01492_),
    .Q_N(_13836_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2345),
    .D(_01493_),
    .Q_N(_13835_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2346),
    .D(_01494_),
    .Q_N(_13834_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2347),
    .D(_01495_),
    .Q_N(_13833_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2348),
    .D(_01496_),
    .Q_N(_13832_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2349),
    .D(_01497_),
    .Q_N(_13831_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2350),
    .D(_01498_),
    .Q_N(_13830_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2351),
    .D(_01499_),
    .Q_N(_13829_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2352),
    .D(_01500_),
    .Q_N(_13828_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2353),
    .D(_01501_),
    .Q_N(_13827_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2354),
    .D(_01502_),
    .Q_N(_13826_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2355),
    .D(_01503_),
    .Q_N(_13825_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2356),
    .D(_01504_),
    .Q_N(_13824_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2357),
    .D(_01505_),
    .Q_N(_13823_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2358),
    .D(_01506_),
    .Q_N(_13822_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2359),
    .D(_01507_),
    .Q_N(_13821_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2360),
    .D(_01508_),
    .Q_N(_13820_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2361),
    .D(_01509_),
    .Q_N(_13819_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2362),
    .D(_01510_),
    .Q_N(_13818_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2363),
    .D(_01511_),
    .Q_N(_13817_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2364),
    .D(_01512_),
    .Q_N(_13816_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2365),
    .D(_01513_),
    .Q_N(_13815_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2366),
    .D(_01514_),
    .Q_N(_13814_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2367),
    .D(_01515_),
    .Q_N(_13813_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2368),
    .D(_01516_),
    .Q_N(_13812_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2369),
    .D(_01517_),
    .Q_N(_13811_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2370),
    .D(_01518_),
    .Q_N(_13810_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2371),
    .D(_01519_),
    .Q_N(_13809_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2372),
    .D(_01520_),
    .Q_N(_13808_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2373),
    .D(_01521_),
    .Q_N(_13807_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2374),
    .D(_01522_),
    .Q_N(_13806_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2375),
    .D(_01523_),
    .Q_N(_13805_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2376),
    .D(_01524_),
    .Q_N(_13804_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2377),
    .D(_01525_),
    .Q_N(_13803_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2378),
    .D(_01526_),
    .Q_N(_13802_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2379),
    .D(_01527_),
    .Q_N(_13801_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2380),
    .D(_01528_),
    .Q_N(_13800_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2381),
    .D(_01529_),
    .Q_N(_13799_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2382),
    .D(_01530_),
    .Q_N(_13798_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2383),
    .D(_01531_),
    .Q_N(_13797_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2384),
    .D(_01532_),
    .Q_N(_13796_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2385),
    .D(_01533_),
    .Q_N(_13795_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2386),
    .D(_01534_),
    .Q_N(_13794_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2387),
    .D(_01535_),
    .Q_N(_13793_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2388),
    .D(_01536_),
    .Q_N(_13792_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2389),
    .D(_01537_),
    .Q_N(_13791_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2390),
    .D(_01538_),
    .Q_N(_13790_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2391),
    .D(_01539_),
    .Q_N(_13789_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2392),
    .D(_01540_),
    .Q_N(_13788_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2393),
    .D(_01541_),
    .Q_N(_13787_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2394),
    .D(_01542_),
    .Q_N(_13786_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2395),
    .D(_01543_),
    .Q_N(_13785_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2396),
    .D(_01544_),
    .Q_N(_13784_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2397),
    .D(_01545_),
    .Q_N(_13783_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2398),
    .D(_01546_),
    .Q_N(_13782_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2399),
    .D(_01547_),
    .Q_N(_13781_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2400),
    .D(_01548_),
    .Q_N(_13780_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2401),
    .D(_01549_),
    .Q_N(_13779_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2402),
    .D(_01550_),
    .Q_N(_13778_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2403),
    .D(_01551_),
    .Q_N(_13777_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2404),
    .D(_01552_),
    .Q_N(_13776_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2405),
    .D(_01553_),
    .Q_N(_13775_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2406),
    .D(_01554_),
    .Q_N(_13774_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2407),
    .D(_01555_),
    .Q_N(_13773_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2408),
    .D(_01556_),
    .Q_N(_13772_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2409),
    .D(_01557_),
    .Q_N(_13771_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2410),
    .D(_01558_),
    .Q_N(_13770_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2411),
    .D(_01559_),
    .Q_N(_13769_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2412),
    .D(_01560_),
    .Q_N(_13768_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2413),
    .D(_01561_),
    .Q_N(_13767_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2414),
    .D(_01562_),
    .Q_N(_13766_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2415),
    .D(_01563_),
    .Q_N(_13765_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2416),
    .D(_01564_),
    .Q_N(_13764_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2417),
    .D(_01565_),
    .Q_N(_13763_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2418),
    .D(_01566_),
    .Q_N(_13762_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2419),
    .D(_01567_),
    .Q_N(_13761_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2420),
    .D(_01568_),
    .Q_N(_13760_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2421),
    .D(_01569_),
    .Q_N(_13759_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2422),
    .D(_01570_),
    .Q_N(_13758_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2423),
    .D(_01571_),
    .Q_N(_13757_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2424),
    .D(_01572_),
    .Q_N(_13756_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2425),
    .D(_01573_),
    .Q_N(_13755_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2426),
    .D(_01574_),
    .Q_N(_13754_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2427),
    .D(_01575_),
    .Q_N(_13753_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2428),
    .D(_01576_),
    .Q_N(_13752_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2429),
    .D(_01577_),
    .Q_N(_13751_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2430),
    .D(_01578_),
    .Q_N(_13750_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2431),
    .D(_01579_),
    .Q_N(_13749_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2432),
    .D(_01580_),
    .Q_N(_13748_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2433),
    .D(_01581_),
    .Q_N(_13747_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2434),
    .D(_01582_),
    .Q_N(_13746_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2435),
    .D(_01583_),
    .Q_N(_13745_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2436),
    .D(_01584_),
    .Q_N(_13744_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2437),
    .D(_01585_),
    .Q_N(_13743_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2438),
    .D(_01586_),
    .Q_N(_13742_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2439),
    .D(_01587_),
    .Q_N(_13741_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2440),
    .D(_01588_),
    .Q_N(_13740_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2441),
    .D(_01589_),
    .Q_N(_13739_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2442),
    .D(_01590_),
    .Q_N(_13738_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2443),
    .D(_01591_),
    .Q_N(_13737_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2444),
    .D(_01592_),
    .Q_N(_13736_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2445),
    .D(_01593_),
    .Q_N(_13735_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2446),
    .D(_01594_),
    .Q_N(_13734_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2447),
    .D(_01595_),
    .Q_N(_13733_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2448),
    .D(_01596_),
    .Q_N(_13732_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2449),
    .D(_01597_),
    .Q_N(_13731_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2450),
    .D(_01598_),
    .Q_N(_13730_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2451),
    .D(_01599_),
    .Q_N(_13729_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2452),
    .D(_01600_),
    .Q_N(_13728_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2453),
    .D(_01601_),
    .Q_N(_13727_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2454),
    .D(_01602_),
    .Q_N(_13726_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2455),
    .D(_01603_),
    .Q_N(_13725_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2456),
    .D(_01604_),
    .Q_N(_13724_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2457),
    .D(_01605_),
    .Q_N(_13723_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2458),
    .D(_01606_),
    .Q_N(_13722_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2459),
    .D(_01607_),
    .Q_N(_13721_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2460),
    .D(_01608_),
    .Q_N(_13720_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2461),
    .D(_01609_),
    .Q_N(_13719_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2462),
    .D(_01610_),
    .Q_N(_13718_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2463),
    .D(_01611_),
    .Q_N(_13717_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2464),
    .D(_01612_),
    .Q_N(_13716_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2465),
    .D(_01613_),
    .Q_N(_13715_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2466),
    .D(_01614_),
    .Q_N(_13714_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2467),
    .D(_01615_),
    .Q_N(_13713_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2468),
    .D(_01616_),
    .Q_N(_13712_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2469),
    .D(_01617_),
    .Q_N(_13711_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2470),
    .D(_01618_),
    .Q_N(_13710_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2471),
    .D(_01619_),
    .Q_N(_13709_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2472),
    .D(_01620_),
    .Q_N(_13708_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2473),
    .D(_01621_),
    .Q_N(_13707_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2474),
    .D(_01622_),
    .Q_N(_13706_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2475),
    .D(_01623_),
    .Q_N(_13705_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2476),
    .D(_01624_),
    .Q_N(_13704_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2477),
    .D(_01625_),
    .Q_N(_13703_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2478),
    .D(_01626_),
    .Q_N(_13702_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2479),
    .D(_01627_),
    .Q_N(_13701_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2480),
    .D(_01628_),
    .Q_N(_13700_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2481),
    .D(_01629_),
    .Q_N(_13699_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2482),
    .D(_01630_),
    .Q_N(_13698_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2483),
    .D(_01631_),
    .Q_N(_13697_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2484),
    .D(_01632_),
    .Q_N(_13696_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2485),
    .D(_01633_),
    .Q_N(_13695_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2486),
    .D(_01634_),
    .Q_N(_13694_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2487),
    .D(_01635_),
    .Q_N(_13693_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2488),
    .D(_01636_),
    .Q_N(_13692_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2489),
    .D(_01637_),
    .Q_N(_13691_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2490),
    .D(_01638_),
    .Q_N(_13690_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2491),
    .D(_01639_),
    .Q_N(_13689_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2492),
    .D(_01640_),
    .Q_N(_13688_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2493),
    .D(_01641_),
    .Q_N(_13687_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2494),
    .D(_01642_),
    .Q_N(_13686_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2495),
    .D(_01643_),
    .Q_N(_13685_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2496),
    .D(_01644_),
    .Q_N(_13684_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2497),
    .D(_01645_),
    .Q_N(_13683_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2498),
    .D(_01646_),
    .Q_N(_13682_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2499),
    .D(_01647_),
    .Q_N(_13681_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2500),
    .D(_01648_),
    .Q_N(_13680_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2501),
    .D(_01649_),
    .Q_N(_13679_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2502),
    .D(_01650_),
    .Q_N(_13678_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2503),
    .D(_01651_),
    .Q_N(_13677_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2504),
    .D(_01652_),
    .Q_N(_13676_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2505),
    .D(_01653_),
    .Q_N(_13675_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2506),
    .D(_01654_),
    .Q_N(_13674_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2507),
    .D(_01655_),
    .Q_N(_13673_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2508),
    .D(_01656_),
    .Q_N(_13672_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2509),
    .D(_01657_),
    .Q_N(_13671_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2510),
    .D(_01658_),
    .Q_N(_13670_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2511),
    .D(_01659_),
    .Q_N(_13669_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2512),
    .D(_01660_),
    .Q_N(_13668_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2513),
    .D(_01661_),
    .Q_N(_13667_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2514),
    .D(_01662_),
    .Q_N(_13666_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2515),
    .D(_01663_),
    .Q_N(_13665_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2516),
    .D(_01664_),
    .Q_N(_13664_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2517),
    .D(_01665_),
    .Q_N(_13663_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2518),
    .D(_01666_),
    .Q_N(_13662_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2519),
    .D(_01667_),
    .Q_N(_13661_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2520),
    .D(_01668_),
    .Q_N(_13660_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2521),
    .D(_01669_),
    .Q_N(_13659_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2522),
    .D(_01670_),
    .Q_N(_13658_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2523),
    .D(_01671_),
    .Q_N(_13657_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2524),
    .D(_01672_),
    .Q_N(_13656_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2525),
    .D(_01673_),
    .Q_N(_13655_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2526),
    .D(_01674_),
    .Q_N(_13654_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net2527),
    .D(_01675_),
    .Q_N(_13653_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2528),
    .D(_01676_),
    .Q_N(_13652_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2529),
    .D(_01677_),
    .Q_N(_13651_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2530),
    .D(_01678_),
    .Q_N(_13650_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2531),
    .D(_01679_),
    .Q_N(_13649_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2532),
    .D(_01680_),
    .Q_N(_13648_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2533),
    .D(_01681_),
    .Q_N(_13647_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2534),
    .D(_01682_),
    .Q_N(_13646_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2535),
    .D(_01683_),
    .Q_N(_13645_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2536),
    .D(_01684_),
    .Q_N(_13644_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2537),
    .D(_01685_),
    .Q_N(_13643_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2538),
    .D(_01686_),
    .Q_N(_13642_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2539),
    .D(_01687_),
    .Q_N(_13641_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2540),
    .D(_01688_),
    .Q_N(_13640_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2541),
    .D(_01689_),
    .Q_N(_13639_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2542),
    .D(_01690_),
    .Q_N(_13638_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2543),
    .D(_01691_),
    .Q_N(_13637_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2544),
    .D(_01692_),
    .Q_N(_13636_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2545),
    .D(_01693_),
    .Q_N(_13635_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2546),
    .D(_01694_),
    .Q_N(_13634_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2547),
    .D(_01695_),
    .Q_N(_13633_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2548),
    .D(_01696_),
    .Q_N(_13632_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2549),
    .D(_01697_),
    .Q_N(_13631_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2550),
    .D(_01698_),
    .Q_N(_13630_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net2551),
    .D(_01699_),
    .Q_N(_13629_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2552),
    .D(_01700_),
    .Q_N(_13628_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2553),
    .D(_01701_),
    .Q_N(_13627_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2554),
    .D(_01702_),
    .Q_N(_13626_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2555),
    .D(_01703_),
    .Q_N(_13625_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2556),
    .D(_01704_),
    .Q_N(_13624_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2557),
    .D(_01705_),
    .Q_N(_13623_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2558),
    .D(_01706_),
    .Q_N(_13622_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2559),
    .D(_01707_),
    .Q_N(_13621_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2560),
    .D(_01708_),
    .Q_N(_13620_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net2561),
    .D(_01709_),
    .Q_N(_13619_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2562),
    .D(_01710_),
    .Q_N(_13618_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2563),
    .D(_01711_),
    .Q_N(_13617_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2564),
    .D(_01712_),
    .Q_N(_13616_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2565),
    .D(_01713_),
    .Q_N(_13615_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2566),
    .D(_01714_),
    .Q_N(_13614_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2567),
    .D(_01715_),
    .Q_N(_13613_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2568),
    .D(_01716_),
    .Q_N(_13612_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2569),
    .D(_01717_),
    .Q_N(_13611_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2570),
    .D(_01718_),
    .Q_N(_13610_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2571),
    .D(_01719_),
    .Q_N(_13609_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2572),
    .D(_01720_),
    .Q_N(_13608_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2573),
    .D(_01721_),
    .Q_N(_13607_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2574),
    .D(_01722_),
    .Q_N(_13606_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2575),
    .D(_01723_),
    .Q_N(_13605_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2576),
    .D(_01724_),
    .Q_N(_13604_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2577),
    .D(_01725_),
    .Q_N(_13603_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2578),
    .D(_01726_),
    .Q_N(_13602_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2579),
    .D(_01727_),
    .Q_N(_13601_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2580),
    .D(_01728_),
    .Q_N(_13600_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2581),
    .D(_01729_),
    .Q_N(_13599_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2582),
    .D(_01730_),
    .Q_N(_13598_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2583),
    .D(_01731_),
    .Q_N(_13597_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2584),
    .D(_01732_),
    .Q_N(_13596_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2585),
    .D(_01733_),
    .Q_N(_13595_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2586),
    .D(_01734_),
    .Q_N(_13594_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2587),
    .D(_01735_),
    .Q_N(_13593_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2588),
    .D(_01736_),
    .Q_N(_13592_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2589),
    .D(_01737_),
    .Q_N(_13591_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2590),
    .D(_01738_),
    .Q_N(_13590_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2591),
    .D(_01739_),
    .Q_N(_13589_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2592),
    .D(_01740_),
    .Q_N(_13588_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2593),
    .D(_01741_),
    .Q_N(_13587_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2594),
    .D(_01742_),
    .Q_N(_13586_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2595),
    .D(_01743_),
    .Q_N(_13585_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2596),
    .D(_01744_),
    .Q_N(_13584_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2597),
    .D(_01745_),
    .Q_N(_13583_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2598),
    .D(_01746_),
    .Q_N(_13582_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2599),
    .D(_01747_),
    .Q_N(_13581_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2600),
    .D(_01748_),
    .Q_N(_13580_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2601),
    .D(_01749_),
    .Q_N(_13579_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2602),
    .D(_01750_),
    .Q_N(_13578_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2603),
    .D(_01751_),
    .Q_N(_13577_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2604),
    .D(_01752_),
    .Q_N(_13576_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2605),
    .D(_01753_),
    .Q_N(_13575_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2606),
    .D(_01754_),
    .Q_N(_13574_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2607),
    .D(_01755_),
    .Q_N(_13573_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2608),
    .D(_01756_),
    .Q_N(_13572_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2609),
    .D(_01757_),
    .Q_N(_13571_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2610),
    .D(_01758_),
    .Q_N(_13570_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2611),
    .D(_01759_),
    .Q_N(_13569_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2612),
    .D(_01760_),
    .Q_N(_13568_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2613),
    .D(_01761_),
    .Q_N(_13567_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2614),
    .D(_01762_),
    .Q_N(_13566_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2615),
    .D(_01763_),
    .Q_N(_13565_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2616),
    .D(_01764_),
    .Q_N(_13564_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2617),
    .D(_01765_),
    .Q_N(_13563_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2618),
    .D(_01766_),
    .Q_N(_13562_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2619),
    .D(_01767_),
    .Q_N(_13561_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2620),
    .D(_01768_),
    .Q_N(_13560_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2621),
    .D(_01769_),
    .Q_N(_13559_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2622),
    .D(_01770_),
    .Q_N(_13558_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2623),
    .D(_01771_),
    .Q_N(_13557_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2624),
    .D(_01772_),
    .Q_N(_13556_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2625),
    .D(_01773_),
    .Q_N(_13555_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2626),
    .D(_01774_),
    .Q_N(_13554_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2627),
    .D(_01775_),
    .Q_N(_13553_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2628),
    .D(_01776_),
    .Q_N(_13552_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2629),
    .D(_01777_),
    .Q_N(_13551_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2630),
    .D(_01778_),
    .Q_N(_13550_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2631),
    .D(_01779_),
    .Q_N(_13549_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2632),
    .D(_01780_),
    .Q_N(_13548_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2633),
    .D(_01781_),
    .Q_N(_13547_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2634),
    .D(_01782_),
    .Q_N(_13546_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2635),
    .D(_01783_),
    .Q_N(_13545_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2636),
    .D(_01784_),
    .Q_N(_13544_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2637),
    .D(_01785_),
    .Q_N(_13543_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2638),
    .D(_01786_),
    .Q_N(_13542_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2639),
    .D(_01787_),
    .Q_N(_13541_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2640),
    .D(_01788_),
    .Q_N(_13540_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2641),
    .D(_01789_),
    .Q_N(_13539_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2642),
    .D(_01790_),
    .Q_N(_13538_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2643),
    .D(_01791_),
    .Q_N(_13537_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2644),
    .D(_01792_),
    .Q_N(_13536_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2645),
    .D(_01793_),
    .Q_N(_13535_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2646),
    .D(_01794_),
    .Q_N(_13534_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2647),
    .D(_01795_),
    .Q_N(_13533_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2648),
    .D(_01796_),
    .Q_N(_13532_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2649),
    .D(_01797_),
    .Q_N(_13531_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2650),
    .D(_01798_),
    .Q_N(_13530_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2651),
    .D(_01799_),
    .Q_N(_13529_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2652),
    .D(_01800_),
    .Q_N(_13528_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2653),
    .D(_01801_),
    .Q_N(_13527_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2654),
    .D(_01802_),
    .Q_N(_13526_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2655),
    .D(_01803_),
    .Q_N(_13525_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2656),
    .D(_01804_),
    .Q_N(_13524_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2657),
    .D(_01805_),
    .Q_N(_13523_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2658),
    .D(_01806_),
    .Q_N(_13522_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2659),
    .D(_01807_),
    .Q_N(_13521_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2660),
    .D(_01808_),
    .Q_N(_13520_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2661),
    .D(_01809_),
    .Q_N(_13519_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2662),
    .D(_01810_),
    .Q_N(_13518_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2663),
    .D(_01811_),
    .Q_N(_13517_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2664),
    .D(_01812_),
    .Q_N(_13516_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2665),
    .D(_01813_),
    .Q_N(_13515_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2666),
    .D(_01814_),
    .Q_N(_13514_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2667),
    .D(_01815_),
    .Q_N(_13513_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2668),
    .D(_01816_),
    .Q_N(_13512_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2669),
    .D(_01817_),
    .Q_N(_13511_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2670),
    .D(_01818_),
    .Q_N(_13510_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2671),
    .D(_01819_),
    .Q_N(_13509_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2672),
    .D(_01820_),
    .Q_N(_13508_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2673),
    .D(_01821_),
    .Q_N(_13507_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2674),
    .D(_01822_),
    .Q_N(_13506_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2675),
    .D(_01823_),
    .Q_N(_13505_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2676),
    .D(_01824_),
    .Q_N(_13504_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2677),
    .D(_01825_),
    .Q_N(_13503_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2678),
    .D(_01826_),
    .Q_N(_13502_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2679),
    .D(_01827_),
    .Q_N(_13501_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2680),
    .D(_01828_),
    .Q_N(_13500_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2681),
    .D(_01829_),
    .Q_N(_13499_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2682),
    .D(_01830_),
    .Q_N(_13498_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2683),
    .D(_01831_),
    .Q_N(_13497_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2684),
    .D(_01832_),
    .Q_N(_13496_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2685),
    .D(_01833_),
    .Q_N(_13495_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2686),
    .D(_01834_),
    .Q_N(_13494_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2687),
    .D(_01835_),
    .Q_N(_13493_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2688),
    .D(_01836_),
    .Q_N(_13492_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2689),
    .D(_01837_),
    .Q_N(_13491_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2690),
    .D(_01838_),
    .Q_N(_13490_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2691),
    .D(_01839_),
    .Q_N(_13489_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2692),
    .D(_01840_),
    .Q_N(_13488_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2693),
    .D(_01841_),
    .Q_N(_13487_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2694),
    .D(_01842_),
    .Q_N(_13486_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2695),
    .D(_01843_),
    .Q_N(_13485_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2696),
    .D(_01844_),
    .Q_N(_13484_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2697),
    .D(_01845_),
    .Q_N(_13483_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2698),
    .D(_01846_),
    .Q_N(_13482_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2699),
    .D(_01847_),
    .Q_N(_13481_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2700),
    .D(_01848_),
    .Q_N(_13480_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2701),
    .D(_01849_),
    .Q_N(_13479_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2702),
    .D(_01850_),
    .Q_N(_13478_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2703),
    .D(_01851_),
    .Q_N(_13477_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2704),
    .D(_01852_),
    .Q_N(_13476_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2705),
    .D(_01853_),
    .Q_N(_13475_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2706),
    .D(_01854_),
    .Q_N(_13474_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2707),
    .D(_01855_),
    .Q_N(_13473_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2708),
    .D(_01856_),
    .Q_N(_13472_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2709),
    .D(_01857_),
    .Q_N(_13471_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2710),
    .D(_01858_),
    .Q_N(_13470_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2711),
    .D(_01859_),
    .Q_N(_13469_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2712),
    .D(_01860_),
    .Q_N(_13468_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2713),
    .D(_01861_),
    .Q_N(_13467_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2714),
    .D(_01862_),
    .Q_N(_13466_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2715),
    .D(_01863_),
    .Q_N(_13465_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2716),
    .D(_01864_),
    .Q_N(_13464_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2717),
    .D(_01865_),
    .Q_N(_13463_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2718),
    .D(_01866_),
    .Q_N(_13462_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2719),
    .D(_01867_),
    .Q_N(_13461_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2720),
    .D(_01868_),
    .Q_N(_13460_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2721),
    .D(_01869_),
    .Q_N(_13459_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2722),
    .D(_01870_),
    .Q_N(_13458_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2723),
    .D(_01871_),
    .Q_N(_13457_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2724),
    .D(_01872_),
    .Q_N(_13456_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2725),
    .D(_01873_),
    .Q_N(_13455_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2726),
    .D(_01874_),
    .Q_N(_13454_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2727),
    .D(_01875_),
    .Q_N(_13453_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2728),
    .D(_01876_),
    .Q_N(_13452_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2729),
    .D(_01877_),
    .Q_N(_13451_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2730),
    .D(_01878_),
    .Q_N(_13450_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2731),
    .D(_01879_),
    .Q_N(_13449_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2732),
    .D(_01880_),
    .Q_N(_13448_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2733),
    .D(_01881_),
    .Q_N(_13447_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2734),
    .D(_01882_),
    .Q_N(_13446_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2735),
    .D(_01883_),
    .Q_N(_13445_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2736),
    .D(_01884_),
    .Q_N(_13444_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2737),
    .D(_01885_),
    .Q_N(_13443_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2738),
    .D(_01886_),
    .Q_N(_13442_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2739),
    .D(_01887_),
    .Q_N(_13441_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2740),
    .D(_01888_),
    .Q_N(_13440_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2741),
    .D(_01889_),
    .Q_N(_13439_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2742),
    .D(_01890_),
    .Q_N(_13438_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2743),
    .D(_01891_),
    .Q_N(_13437_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2744),
    .D(_01892_),
    .Q_N(_13436_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2745),
    .D(_01893_),
    .Q_N(_13435_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2746),
    .D(_01894_),
    .Q_N(_13434_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2747),
    .D(_01895_),
    .Q_N(_13433_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2748),
    .D(_01896_),
    .Q_N(_13432_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2749),
    .D(_01897_),
    .Q_N(_13431_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2750),
    .D(_01898_),
    .Q_N(_13430_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2751),
    .D(_01899_),
    .Q_N(_13429_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2752),
    .D(_01900_),
    .Q_N(_13428_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2753),
    .D(_01901_),
    .Q_N(_13427_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2754),
    .D(_01902_),
    .Q_N(_13426_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2755),
    .D(_01903_),
    .Q_N(_13425_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2756),
    .D(_01904_),
    .Q_N(_13424_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2757),
    .D(_01905_),
    .Q_N(_13423_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2758),
    .D(_01906_),
    .Q_N(_13422_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2759),
    .D(_01907_),
    .Q_N(_13421_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2760),
    .D(_01908_),
    .Q_N(_13420_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2761),
    .D(_01909_),
    .Q_N(_13419_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2762),
    .D(_01910_),
    .Q_N(_13418_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2763),
    .D(_01911_),
    .Q_N(_13417_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2764),
    .D(_01912_),
    .Q_N(_13416_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2765),
    .D(_01913_),
    .Q_N(_13415_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2766),
    .D(_01914_),
    .Q_N(_13414_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2767),
    .D(_01915_),
    .Q_N(_13413_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2768),
    .D(_01916_),
    .Q_N(_13412_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2769),
    .D(_01917_),
    .Q_N(_13411_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2770),
    .D(_01918_),
    .Q_N(_13410_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2771),
    .D(_01919_),
    .Q_N(_13409_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2772),
    .D(_01920_),
    .Q_N(_13408_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2773),
    .D(_01921_),
    .Q_N(_13407_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2774),
    .D(_01922_),
    .Q_N(_13406_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2775),
    .D(_01923_),
    .Q_N(_13405_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2776),
    .D(_01924_),
    .Q_N(_13404_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2777),
    .D(_01925_),
    .Q_N(_13403_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2778),
    .D(_01926_),
    .Q_N(_13402_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2779),
    .D(_01927_),
    .Q_N(_13401_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2780),
    .D(_01928_),
    .Q_N(_13400_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2781),
    .D(_01929_),
    .Q_N(_13399_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2782),
    .D(_01930_),
    .Q_N(_13398_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2783),
    .D(_01931_),
    .Q_N(_13397_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2784),
    .D(_01932_),
    .Q_N(_13396_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2785),
    .D(_01933_),
    .Q_N(_13395_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2786),
    .D(_01934_),
    .Q_N(_13394_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2787),
    .D(_01935_),
    .Q_N(_13393_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2788),
    .D(_01936_),
    .Q_N(_13392_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2789),
    .D(_01937_),
    .Q_N(_13391_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2790),
    .D(_01938_),
    .Q_N(_13390_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[9] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2791),
    .D(_01939_),
    .Q_N(_13389_),
    .Q(\cpu.gpio.r_enable_in[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2792),
    .D(_01940_),
    .Q_N(_13388_),
    .Q(\cpu.gpio.r_enable_in[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2793),
    .D(_01941_),
    .Q_N(_13387_),
    .Q(\cpu.gpio.r_enable_in[2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2794),
    .D(_01942_),
    .Q_N(_13386_),
    .Q(\cpu.gpio.r_enable_in[3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2795),
    .D(_01943_),
    .Q_N(_13385_),
    .Q(\cpu.gpio.r_enable_in[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2796),
    .D(_01944_),
    .Q_N(_13384_),
    .Q(\cpu.gpio.r_enable_in[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2797),
    .D(_01945_),
    .Q_N(_13383_),
    .Q(\cpu.gpio.r_enable_in[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2798),
    .D(_01946_),
    .Q_N(_13382_),
    .Q(\cpu.gpio.r_enable_in[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2799),
    .D(_01947_),
    .Q_N(_13381_),
    .Q(\cpu.gpio.r_enable_io[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2800),
    .D(_01948_),
    .Q_N(_13380_),
    .Q(\cpu.gpio.r_enable_io[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2801),
    .D(_01949_),
    .Q_N(_13379_),
    .Q(\cpu.gpio.r_enable_io[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2802),
    .D(_01950_),
    .Q_N(_13378_),
    .Q(\cpu.gpio.r_enable_io[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2803),
    .D(_01951_),
    .Q_N(_13377_),
    .Q(net7));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2804),
    .D(_01952_),
    .Q_N(_13376_),
    .Q(net8));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2805),
    .D(_01953_),
    .Q_N(_13375_),
    .Q(net9));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2806),
    .D(_01954_),
    .Q_N(_13374_),
    .Q(net10));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[0]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2807),
    .D(_01955_),
    .Q_N(_13373_),
    .Q(\cpu.gpio.genblk2[4].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[1]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2808),
    .D(_01956_),
    .Q_N(_13372_),
    .Q(\cpu.gpio.genblk2[5].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2809),
    .D(_01957_),
    .Q_N(_13371_),
    .Q(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2810),
    .D(_01958_),
    .Q_N(_13370_),
    .Q(\cpu.gpio.genblk2[7].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[0]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2811),
    .D(_01959_),
    .Q_N(_13369_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[1]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2812),
    .D(_01960_),
    .Q_N(_13368_),
    .Q(\cpu.gpio.genblk1[4].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[2]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2813),
    .D(_01961_),
    .Q_N(_13367_),
    .Q(\cpu.gpio.genblk1[5].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[3]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2814),
    .D(_01962_),
    .Q_N(_13366_),
    .Q(\cpu.gpio.genblk1[6].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[4]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2815),
    .D(_01963_),
    .Q_N(_13365_),
    .Q(\cpu.gpio.genblk1[7].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2816),
    .D(_01964_),
    .Q_N(_13364_),
    .Q(\cpu.gpio.r_spi_miso_src[0][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2817),
    .D(_01965_),
    .Q_N(_00100_),
    .Q(\cpu.gpio.r_spi_miso_src[0][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2818),
    .D(_01966_),
    .Q_N(_00110_),
    .Q(\cpu.gpio.r_spi_miso_src[0][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2819),
    .D(_01967_),
    .Q_N(_00119_),
    .Q(\cpu.gpio.r_spi_miso_src[0][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2820),
    .D(_01968_),
    .Q_N(_13363_),
    .Q(\cpu.gpio.r_spi_miso_src[1][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2821),
    .D(_01969_),
    .Q_N(_00138_),
    .Q(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2822),
    .D(_01970_),
    .Q_N(_00150_),
    .Q(\cpu.gpio.r_spi_miso_src[1][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2823),
    .D(_01971_),
    .Q_N(_00162_),
    .Q(\cpu.gpio.r_spi_miso_src[1][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2824),
    .D(_01972_),
    .Q_N(_13362_),
    .Q(\cpu.gpio.r_src_io[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2825),
    .D(_01973_),
    .Q_N(_13361_),
    .Q(\cpu.gpio.r_src_io[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2826),
    .D(_01974_),
    .Q_N(_00187_),
    .Q(\cpu.gpio.r_src_io[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2827),
    .D(_01975_),
    .Q_N(_13360_),
    .Q(\cpu.gpio.r_src_io[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2828),
    .D(_01976_),
    .Q_N(_13359_),
    .Q(\cpu.gpio.r_src_io[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2829),
    .D(_01977_),
    .Q_N(_13358_),
    .Q(\cpu.gpio.r_src_io[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2830),
    .D(_01978_),
    .Q_N(_00186_),
    .Q(\cpu.gpio.r_src_io[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2831),
    .D(_01979_),
    .Q_N(_13357_),
    .Q(\cpu.gpio.r_src_io[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2832),
    .D(_01980_),
    .Q_N(_13356_),
    .Q(\cpu.gpio.r_src_io[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2833),
    .D(_01981_),
    .Q_N(_00096_),
    .Q(\cpu.gpio.r_src_io[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2834),
    .D(_01982_),
    .Q_N(_00106_),
    .Q(\cpu.gpio.r_src_io[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2835),
    .D(_01983_),
    .Q_N(_00116_),
    .Q(\cpu.gpio.r_src_io[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2836),
    .D(_01984_),
    .Q_N(_13355_),
    .Q(\cpu.gpio.r_src_io[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2837),
    .D(_01985_),
    .Q_N(_00134_),
    .Q(\cpu.gpio.r_src_io[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2838),
    .D(_01986_),
    .Q_N(_00146_),
    .Q(\cpu.gpio.r_src_io[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2839),
    .D(_01987_),
    .Q_N(_00158_),
    .Q(\cpu.gpio.r_src_io[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2840),
    .D(_01988_),
    .Q_N(_13354_),
    .Q(\cpu.gpio.r_src_o[3][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2841),
    .D(_01989_),
    .Q_N(_00137_),
    .Q(\cpu.gpio.r_src_o[3][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2842),
    .D(_01990_),
    .Q_N(_00149_),
    .Q(\cpu.gpio.r_src_o[3][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2843),
    .D(_01991_),
    .Q_N(_00161_),
    .Q(\cpu.gpio.r_src_o[3][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2844),
    .D(_01992_),
    .Q_N(_13353_),
    .Q(\cpu.gpio.r_src_o[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2845),
    .D(_01993_),
    .Q_N(_00098_),
    .Q(\cpu.gpio.r_src_o[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2846),
    .D(_01994_),
    .Q_N(_00108_),
    .Q(\cpu.gpio.r_src_o[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2847),
    .D(_01995_),
    .Q_N(_00118_),
    .Q(\cpu.gpio.r_src_o[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2848),
    .D(_01996_),
    .Q_N(_13352_),
    .Q(\cpu.gpio.r_src_o[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2849),
    .D(_01997_),
    .Q_N(_00136_),
    .Q(\cpu.gpio.r_src_o[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2850),
    .D(_01998_),
    .Q_N(_00148_),
    .Q(\cpu.gpio.r_src_o[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2851),
    .D(_01999_),
    .Q_N(_00160_),
    .Q(\cpu.gpio.r_src_o[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2852),
    .D(_02000_),
    .Q_N(_13351_),
    .Q(\cpu.gpio.r_src_o[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2853),
    .D(_02001_),
    .Q_N(_00097_),
    .Q(\cpu.gpio.r_src_o[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2854),
    .D(_02002_),
    .Q_N(_00107_),
    .Q(\cpu.gpio.r_src_o[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2855),
    .D(_02003_),
    .Q_N(_00117_),
    .Q(\cpu.gpio.r_src_o[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2856),
    .D(_02004_),
    .Q_N(_13350_),
    .Q(\cpu.gpio.r_src_o[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2857),
    .D(_02005_),
    .Q_N(_00135_),
    .Q(\cpu.gpio.r_src_o[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2858),
    .D(_02006_),
    .Q_N(_00147_),
    .Q(\cpu.gpio.r_src_o[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2859),
    .D(_02007_),
    .Q_N(_00159_),
    .Q(\cpu.gpio.r_src_o[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2860),
    .D(_02008_),
    .Q_N(_13349_),
    .Q(\cpu.gpio.r_uart_rx_src[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2861),
    .D(_02009_),
    .Q_N(_00099_),
    .Q(\cpu.gpio.r_uart_rx_src[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2862),
    .D(_02010_),
    .Q_N(_00109_),
    .Q(\cpu.gpio.r_uart_rx_src[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2863),
    .D(_02011_),
    .Q_N(_13348_),
    .Q(\cpu.icache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2864),
    .D(_02012_),
    .Q_N(_00203_),
    .Q(\cpu.icache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2865),
    .D(_02013_),
    .Q_N(_00205_),
    .Q(\cpu.icache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2866),
    .D(_02014_),
    .Q_N(_00211_),
    .Q(\cpu.icache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2867),
    .D(_02015_),
    .Q_N(_13347_),
    .Q(\cpu.icache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2868),
    .D(_02016_),
    .Q_N(_13346_),
    .Q(\cpu.icache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2869),
    .D(_02017_),
    .Q_N(_00201_),
    .Q(\cpu.icache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2870),
    .D(_02018_),
    .Q_N(_13345_),
    .Q(\cpu.icache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2871),
    .D(_02019_),
    .Q_N(_13344_),
    .Q(\cpu.icache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2872),
    .D(_02020_),
    .Q_N(_00214_),
    .Q(\cpu.icache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2873),
    .D(_02021_),
    .Q_N(_00216_),
    .Q(\cpu.icache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2874),
    .D(_02022_),
    .Q_N(_13343_),
    .Q(\cpu.icache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2875),
    .D(_02023_),
    .Q_N(_00218_),
    .Q(\cpu.icache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2876),
    .D(_02024_),
    .Q_N(_00208_),
    .Q(\cpu.icache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2877),
    .D(_02025_),
    .Q_N(_00210_),
    .Q(\cpu.icache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2878),
    .D(_02026_),
    .Q_N(_00173_),
    .Q(\cpu.icache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2879),
    .D(_02027_),
    .Q_N(_00175_),
    .Q(\cpu.icache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2880),
    .D(_02028_),
    .Q_N(_00177_),
    .Q(\cpu.icache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2881),
    .D(_02029_),
    .Q_N(_00204_),
    .Q(\cpu.icache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2882),
    .D(_02030_),
    .Q_N(_00206_),
    .Q(\cpu.icache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2883),
    .D(_02031_),
    .Q_N(_00212_),
    .Q(\cpu.icache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2884),
    .D(_02032_),
    .Q_N(_13342_),
    .Q(\cpu.icache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2885),
    .D(_02033_),
    .Q_N(_00213_),
    .Q(\cpu.icache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2886),
    .D(_02034_),
    .Q_N(_13341_),
    .Q(\cpu.icache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2887),
    .D(_02035_),
    .Q_N(_00202_),
    .Q(\cpu.icache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2888),
    .D(_02036_),
    .Q_N(_00215_),
    .Q(\cpu.icache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2889),
    .D(_02037_),
    .Q_N(_00217_),
    .Q(\cpu.icache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2890),
    .D(_02038_),
    .Q_N(_00207_),
    .Q(\cpu.icache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2891),
    .D(_02039_),
    .Q_N(_00209_),
    .Q(\cpu.icache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2892),
    .D(_02040_),
    .Q_N(_00172_),
    .Q(\cpu.icache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2893),
    .D(_02041_),
    .Q_N(_00174_),
    .Q(\cpu.icache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2894),
    .D(_02042_),
    .Q_N(_00176_),
    .Q(\cpu.icache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2895),
    .D(_02043_),
    .Q_N(_13340_),
    .Q(\cpu.icache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2896),
    .D(_02044_),
    .Q_N(_13339_),
    .Q(\cpu.icache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2897),
    .D(_02045_),
    .Q_N(_13338_),
    .Q(\cpu.icache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2898),
    .D(_02046_),
    .Q_N(_13337_),
    .Q(\cpu.icache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2899),
    .D(_02047_),
    .Q_N(_13336_),
    .Q(\cpu.icache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2900),
    .D(_02048_),
    .Q_N(_13335_),
    .Q(\cpu.icache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2901),
    .D(_02049_),
    .Q_N(_13334_),
    .Q(\cpu.icache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2902),
    .D(_02050_),
    .Q_N(_13333_),
    .Q(\cpu.icache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2903),
    .D(_02051_),
    .Q_N(_13332_),
    .Q(\cpu.icache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2904),
    .D(_02052_),
    .Q_N(_13331_),
    .Q(\cpu.icache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2905),
    .D(_02053_),
    .Q_N(_13330_),
    .Q(\cpu.icache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2906),
    .D(_02054_),
    .Q_N(_13329_),
    .Q(\cpu.icache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2907),
    .D(_02055_),
    .Q_N(_13328_),
    .Q(\cpu.icache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2908),
    .D(_02056_),
    .Q_N(_13327_),
    .Q(\cpu.icache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2909),
    .D(_02057_),
    .Q_N(_13326_),
    .Q(\cpu.icache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2910),
    .D(_02058_),
    .Q_N(_13325_),
    .Q(\cpu.icache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2911),
    .D(_02059_),
    .Q_N(_13324_),
    .Q(\cpu.icache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2912),
    .D(_02060_),
    .Q_N(_13323_),
    .Q(\cpu.icache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2913),
    .D(_02061_),
    .Q_N(_13322_),
    .Q(\cpu.icache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2914),
    .D(_02062_),
    .Q_N(_13321_),
    .Q(\cpu.icache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2915),
    .D(_02063_),
    .Q_N(_13320_),
    .Q(\cpu.icache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2916),
    .D(_02064_),
    .Q_N(_13319_),
    .Q(\cpu.icache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2917),
    .D(_02065_),
    .Q_N(_13318_),
    .Q(\cpu.icache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2918),
    .D(_02066_),
    .Q_N(_13317_),
    .Q(\cpu.icache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2919),
    .D(_02067_),
    .Q_N(_13316_),
    .Q(\cpu.icache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2920),
    .D(_02068_),
    .Q_N(_13315_),
    .Q(\cpu.icache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2921),
    .D(_02069_),
    .Q_N(_13314_),
    .Q(\cpu.icache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2922),
    .D(_02070_),
    .Q_N(_13313_),
    .Q(\cpu.icache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2923),
    .D(_02071_),
    .Q_N(_13312_),
    .Q(\cpu.icache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2924),
    .D(_02072_),
    .Q_N(_13311_),
    .Q(\cpu.icache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2925),
    .D(_02073_),
    .Q_N(_13310_),
    .Q(\cpu.icache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2926),
    .D(_02074_),
    .Q_N(_13309_),
    .Q(\cpu.icache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2927),
    .D(_02075_),
    .Q_N(_13308_),
    .Q(\cpu.icache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2928),
    .D(_02076_),
    .Q_N(_13307_),
    .Q(\cpu.icache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2929),
    .D(_02077_),
    .Q_N(_13306_),
    .Q(\cpu.icache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2930),
    .D(_02078_),
    .Q_N(_13305_),
    .Q(\cpu.icache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2931),
    .D(_02079_),
    .Q_N(_13304_),
    .Q(\cpu.icache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2932),
    .D(_02080_),
    .Q_N(_13303_),
    .Q(\cpu.icache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2933),
    .D(_02081_),
    .Q_N(_13302_),
    .Q(\cpu.icache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2934),
    .D(_02082_),
    .Q_N(_13301_),
    .Q(\cpu.icache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2935),
    .D(_02083_),
    .Q_N(_13300_),
    .Q(\cpu.icache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2936),
    .D(_02084_),
    .Q_N(_13299_),
    .Q(\cpu.icache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2937),
    .D(_02085_),
    .Q_N(_13298_),
    .Q(\cpu.icache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2938),
    .D(_02086_),
    .Q_N(_13297_),
    .Q(\cpu.icache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2939),
    .D(_02087_),
    .Q_N(_13296_),
    .Q(\cpu.icache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2940),
    .D(_02088_),
    .Q_N(_13295_),
    .Q(\cpu.icache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2941),
    .D(_02089_),
    .Q_N(_13294_),
    .Q(\cpu.icache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2942),
    .D(_02090_),
    .Q_N(_13293_),
    .Q(\cpu.icache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2943),
    .D(_02091_),
    .Q_N(_13292_),
    .Q(\cpu.icache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2944),
    .D(_02092_),
    .Q_N(_13291_),
    .Q(\cpu.icache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2945),
    .D(_02093_),
    .Q_N(_13290_),
    .Q(\cpu.icache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2946),
    .D(_02094_),
    .Q_N(_13289_),
    .Q(\cpu.icache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2947),
    .D(_02095_),
    .Q_N(_13288_),
    .Q(\cpu.icache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2948),
    .D(_02096_),
    .Q_N(_13287_),
    .Q(\cpu.icache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2949),
    .D(_02097_),
    .Q_N(_13286_),
    .Q(\cpu.icache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2950),
    .D(_02098_),
    .Q_N(_13285_),
    .Q(\cpu.icache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2951),
    .D(_02099_),
    .Q_N(_13284_),
    .Q(\cpu.icache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2952),
    .D(_02100_),
    .Q_N(_13283_),
    .Q(\cpu.icache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2953),
    .D(_02101_),
    .Q_N(_13282_),
    .Q(\cpu.icache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2954),
    .D(_02102_),
    .Q_N(_13281_),
    .Q(\cpu.icache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2955),
    .D(_02103_),
    .Q_N(_13280_),
    .Q(\cpu.icache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2956),
    .D(_02104_),
    .Q_N(_13279_),
    .Q(\cpu.icache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2957),
    .D(_02105_),
    .Q_N(_13278_),
    .Q(\cpu.icache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2958),
    .D(_02106_),
    .Q_N(_13277_),
    .Q(\cpu.icache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2959),
    .D(_02107_),
    .Q_N(_13276_),
    .Q(\cpu.icache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2960),
    .D(_02108_),
    .Q_N(_13275_),
    .Q(\cpu.icache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2961),
    .D(_02109_),
    .Q_N(_13274_),
    .Q(\cpu.icache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2962),
    .D(_02110_),
    .Q_N(_13273_),
    .Q(\cpu.icache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2963),
    .D(_02111_),
    .Q_N(_13272_),
    .Q(\cpu.icache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2964),
    .D(_02112_),
    .Q_N(_13271_),
    .Q(\cpu.icache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2965),
    .D(_02113_),
    .Q_N(_13270_),
    .Q(\cpu.icache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2966),
    .D(_02114_),
    .Q_N(_13269_),
    .Q(\cpu.icache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2967),
    .D(_02115_),
    .Q_N(_13268_),
    .Q(\cpu.icache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2968),
    .D(_02116_),
    .Q_N(_13267_),
    .Q(\cpu.icache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2969),
    .D(_02117_),
    .Q_N(_13266_),
    .Q(\cpu.icache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2970),
    .D(_02118_),
    .Q_N(_13265_),
    .Q(\cpu.icache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2971),
    .D(_02119_),
    .Q_N(_13264_),
    .Q(\cpu.icache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2972),
    .D(_02120_),
    .Q_N(_13263_),
    .Q(\cpu.icache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2973),
    .D(_02121_),
    .Q_N(_13262_),
    .Q(\cpu.icache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2974),
    .D(_02122_),
    .Q_N(_13261_),
    .Q(\cpu.icache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2975),
    .D(_02123_),
    .Q_N(_13260_),
    .Q(\cpu.icache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2976),
    .D(_02124_),
    .Q_N(_13259_),
    .Q(\cpu.icache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2977),
    .D(_02125_),
    .Q_N(_13258_),
    .Q(\cpu.icache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2978),
    .D(_02126_),
    .Q_N(_13257_),
    .Q(\cpu.icache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2979),
    .D(_02127_),
    .Q_N(_13256_),
    .Q(\cpu.icache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2980),
    .D(_02128_),
    .Q_N(_13255_),
    .Q(\cpu.icache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2981),
    .D(_02129_),
    .Q_N(_13254_),
    .Q(\cpu.icache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2982),
    .D(_02130_),
    .Q_N(_13253_),
    .Q(\cpu.icache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2983),
    .D(_02131_),
    .Q_N(_13252_),
    .Q(\cpu.icache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2984),
    .D(_02132_),
    .Q_N(_13251_),
    .Q(\cpu.icache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2985),
    .D(_02133_),
    .Q_N(_13250_),
    .Q(\cpu.icache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2986),
    .D(_02134_),
    .Q_N(_13249_),
    .Q(\cpu.icache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2987),
    .D(_02135_),
    .Q_N(_13248_),
    .Q(\cpu.icache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2988),
    .D(_02136_),
    .Q_N(_13247_),
    .Q(\cpu.icache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2989),
    .D(_02137_),
    .Q_N(_13246_),
    .Q(\cpu.icache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2990),
    .D(_02138_),
    .Q_N(_13245_),
    .Q(\cpu.icache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2991),
    .D(_02139_),
    .Q_N(_13244_),
    .Q(\cpu.icache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2992),
    .D(_02140_),
    .Q_N(_13243_),
    .Q(\cpu.icache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2993),
    .D(_02141_),
    .Q_N(_13242_),
    .Q(\cpu.icache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2994),
    .D(_02142_),
    .Q_N(_13241_),
    .Q(\cpu.icache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2995),
    .D(_02143_),
    .Q_N(_13240_),
    .Q(\cpu.icache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2996),
    .D(_02144_),
    .Q_N(_13239_),
    .Q(\cpu.icache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2997),
    .D(_02145_),
    .Q_N(_13238_),
    .Q(\cpu.icache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2998),
    .D(_02146_),
    .Q_N(_13237_),
    .Q(\cpu.icache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2999),
    .D(_02147_),
    .Q_N(_13236_),
    .Q(\cpu.icache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net3000),
    .D(_02148_),
    .Q_N(_13235_),
    .Q(\cpu.icache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net3001),
    .D(_02149_),
    .Q_N(_13234_),
    .Q(\cpu.icache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net3002),
    .D(_02150_),
    .Q_N(_13233_),
    .Q(\cpu.icache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3003),
    .D(_02151_),
    .Q_N(_13232_),
    .Q(\cpu.icache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net3004),
    .D(_02152_),
    .Q_N(_13231_),
    .Q(\cpu.icache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3005),
    .D(_02153_),
    .Q_N(_13230_),
    .Q(\cpu.icache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net3006),
    .D(_02154_),
    .Q_N(_13229_),
    .Q(\cpu.icache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3007),
    .D(_02155_),
    .Q_N(_13228_),
    .Q(\cpu.icache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3008),
    .D(_02156_),
    .Q_N(_13227_),
    .Q(\cpu.icache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3009),
    .D(_02157_),
    .Q_N(_13226_),
    .Q(\cpu.icache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3010),
    .D(_02158_),
    .Q_N(_13225_),
    .Q(\cpu.icache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3011),
    .D(_02159_),
    .Q_N(_13224_),
    .Q(\cpu.icache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3012),
    .D(_02160_),
    .Q_N(_13223_),
    .Q(\cpu.icache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3013),
    .D(_02161_),
    .Q_N(_13222_),
    .Q(\cpu.icache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3014),
    .D(_02162_),
    .Q_N(_13221_),
    .Q(\cpu.icache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3015),
    .D(_02163_),
    .Q_N(_13220_),
    .Q(\cpu.icache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3016),
    .D(_02164_),
    .Q_N(_13219_),
    .Q(\cpu.icache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net3017),
    .D(_02165_),
    .Q_N(_13218_),
    .Q(\cpu.icache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net3018),
    .D(_02166_),
    .Q_N(_13217_),
    .Q(\cpu.icache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net3019),
    .D(_02167_),
    .Q_N(_13216_),
    .Q(\cpu.icache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net3020),
    .D(_02168_),
    .Q_N(_13215_),
    .Q(\cpu.icache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3021),
    .D(_02169_),
    .Q_N(_13214_),
    .Q(\cpu.icache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3022),
    .D(_02170_),
    .Q_N(_13213_),
    .Q(\cpu.icache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net3023),
    .D(_02171_),
    .Q_N(_13212_),
    .Q(\cpu.icache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3024),
    .D(_02172_),
    .Q_N(_13211_),
    .Q(\cpu.icache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3025),
    .D(_02173_),
    .Q_N(_13210_),
    .Q(\cpu.icache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net3026),
    .D(_02174_),
    .Q_N(_13209_),
    .Q(\cpu.icache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net3027),
    .D(_02175_),
    .Q_N(_13208_),
    .Q(\cpu.icache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net3028),
    .D(_02176_),
    .Q_N(_13207_),
    .Q(\cpu.icache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net3029),
    .D(_02177_),
    .Q_N(_13206_),
    .Q(\cpu.icache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net3030),
    .D(_02178_),
    .Q_N(_13205_),
    .Q(\cpu.icache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net3031),
    .D(_02179_),
    .Q_N(_13204_),
    .Q(\cpu.icache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net3032),
    .D(_02180_),
    .Q_N(_13203_),
    .Q(\cpu.icache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net3033),
    .D(_02181_),
    .Q_N(_13202_),
    .Q(\cpu.icache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net3034),
    .D(_02182_),
    .Q_N(_13201_),
    .Q(\cpu.icache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net3035),
    .D(_02183_),
    .Q_N(_13200_),
    .Q(\cpu.icache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net3036),
    .D(_02184_),
    .Q_N(_13199_),
    .Q(\cpu.icache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net3037),
    .D(_02185_),
    .Q_N(_13198_),
    .Q(\cpu.icache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net3038),
    .D(_02186_),
    .Q_N(_13197_),
    .Q(\cpu.icache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3039),
    .D(_02187_),
    .Q_N(_13196_),
    .Q(\cpu.icache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3040),
    .D(_02188_),
    .Q_N(_13195_),
    .Q(\cpu.icache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3041),
    .D(_02189_),
    .Q_N(_13194_),
    .Q(\cpu.icache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3042),
    .D(_02190_),
    .Q_N(_13193_),
    .Q(\cpu.icache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3043),
    .D(_02191_),
    .Q_N(_13192_),
    .Q(\cpu.icache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net3044),
    .D(_02192_),
    .Q_N(_13191_),
    .Q(\cpu.icache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3045),
    .D(_02193_),
    .Q_N(_13190_),
    .Q(\cpu.icache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3046),
    .D(_02194_),
    .Q_N(_13189_),
    .Q(\cpu.icache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3047),
    .D(_02195_),
    .Q_N(_13188_),
    .Q(\cpu.icache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3048),
    .D(_02196_),
    .Q_N(_13187_),
    .Q(\cpu.icache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net3049),
    .D(_02197_),
    .Q_N(_13186_),
    .Q(\cpu.icache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3050),
    .D(_02198_),
    .Q_N(_13185_),
    .Q(\cpu.icache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3051),
    .D(_02199_),
    .Q_N(_13184_),
    .Q(\cpu.icache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net3052),
    .D(_02200_),
    .Q_N(_13183_),
    .Q(\cpu.icache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3053),
    .D(_02201_),
    .Q_N(_13182_),
    .Q(\cpu.icache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3054),
    .D(_02202_),
    .Q_N(_13181_),
    .Q(\cpu.icache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net3055),
    .D(_02203_),
    .Q_N(_13180_),
    .Q(\cpu.icache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3056),
    .D(_02204_),
    .Q_N(_13179_),
    .Q(\cpu.icache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3057),
    .D(_02205_),
    .Q_N(_13178_),
    .Q(\cpu.icache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3058),
    .D(_02206_),
    .Q_N(_13177_),
    .Q(\cpu.icache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net3059),
    .D(_02207_),
    .Q_N(_13176_),
    .Q(\cpu.icache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net3060),
    .D(_02208_),
    .Q_N(_13175_),
    .Q(\cpu.icache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net3061),
    .D(_02209_),
    .Q_N(_13174_),
    .Q(\cpu.icache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net3062),
    .D(_02210_),
    .Q_N(_13173_),
    .Q(\cpu.icache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net3063),
    .D(_02211_),
    .Q_N(_13172_),
    .Q(\cpu.icache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net3064),
    .D(_02212_),
    .Q_N(_13171_),
    .Q(\cpu.icache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net3065),
    .D(_02213_),
    .Q_N(_13170_),
    .Q(\cpu.icache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3066),
    .D(_02214_),
    .Q_N(_13169_),
    .Q(\cpu.icache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net3067),
    .D(_02215_),
    .Q_N(_13168_),
    .Q(\cpu.icache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net3068),
    .D(_02216_),
    .Q_N(_13167_),
    .Q(\cpu.icache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net3069),
    .D(_02217_),
    .Q_N(_13166_),
    .Q(\cpu.icache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net3070),
    .D(_02218_),
    .Q_N(_13165_),
    .Q(\cpu.icache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3071),
    .D(_02219_),
    .Q_N(_13164_),
    .Q(\cpu.icache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3072),
    .D(_02220_),
    .Q_N(_13163_),
    .Q(\cpu.icache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3073),
    .D(_02221_),
    .Q_N(_13162_),
    .Q(\cpu.icache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3074),
    .D(_02222_),
    .Q_N(_13161_),
    .Q(\cpu.icache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3075),
    .D(_02223_),
    .Q_N(_13160_),
    .Q(\cpu.icache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3076),
    .D(_02224_),
    .Q_N(_13159_),
    .Q(\cpu.icache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3077),
    .D(_02225_),
    .Q_N(_13158_),
    .Q(\cpu.icache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3078),
    .D(_02226_),
    .Q_N(_13157_),
    .Q(\cpu.icache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3079),
    .D(_02227_),
    .Q_N(_13156_),
    .Q(\cpu.icache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3080),
    .D(_02228_),
    .Q_N(_13155_),
    .Q(\cpu.icache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3081),
    .D(_02229_),
    .Q_N(_13154_),
    .Q(\cpu.icache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3082),
    .D(_02230_),
    .Q_N(_13153_),
    .Q(\cpu.icache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3083),
    .D(_02231_),
    .Q_N(_13152_),
    .Q(\cpu.icache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3084),
    .D(_02232_),
    .Q_N(_13151_),
    .Q(\cpu.icache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3085),
    .D(_02233_),
    .Q_N(_13150_),
    .Q(\cpu.icache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3086),
    .D(_02234_),
    .Q_N(_13149_),
    .Q(\cpu.icache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net3087),
    .D(_02235_),
    .Q_N(_13148_),
    .Q(\cpu.icache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3088),
    .D(_02236_),
    .Q_N(_13147_),
    .Q(\cpu.icache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3089),
    .D(_02237_),
    .Q_N(_13146_),
    .Q(\cpu.icache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3090),
    .D(_02238_),
    .Q_N(_13145_),
    .Q(\cpu.icache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net3091),
    .D(_02239_),
    .Q_N(_13144_),
    .Q(\cpu.icache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net3092),
    .D(_02240_),
    .Q_N(_13143_),
    .Q(\cpu.icache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net3093),
    .D(_02241_),
    .Q_N(_13142_),
    .Q(\cpu.icache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3094),
    .D(_02242_),
    .Q_N(_13141_),
    .Q(\cpu.icache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net3095),
    .D(_02243_),
    .Q_N(_13140_),
    .Q(\cpu.icache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3096),
    .D(_02244_),
    .Q_N(_13139_),
    .Q(\cpu.icache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3097),
    .D(_02245_),
    .Q_N(_13138_),
    .Q(\cpu.icache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net3098),
    .D(_02246_),
    .Q_N(_13137_),
    .Q(\cpu.icache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3099),
    .D(_02247_),
    .Q_N(_13136_),
    .Q(\cpu.icache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net3100),
    .D(_02248_),
    .Q_N(_13135_),
    .Q(\cpu.icache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3101),
    .D(_02249_),
    .Q_N(_13134_),
    .Q(\cpu.icache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net3102),
    .D(_02250_),
    .Q_N(_13133_),
    .Q(\cpu.icache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3103),
    .D(_02251_),
    .Q_N(_13132_),
    .Q(\cpu.icache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3104),
    .D(_02252_),
    .Q_N(_13131_),
    .Q(\cpu.icache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3105),
    .D(_02253_),
    .Q_N(_13130_),
    .Q(\cpu.icache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3106),
    .D(_02254_),
    .Q_N(_13129_),
    .Q(\cpu.icache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3107),
    .D(_02255_),
    .Q_N(_13128_),
    .Q(\cpu.icache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3108),
    .D(_02256_),
    .Q_N(_13127_),
    .Q(\cpu.icache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net3109),
    .D(_02257_),
    .Q_N(_13126_),
    .Q(\cpu.icache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3110),
    .D(_02258_),
    .Q_N(_13125_),
    .Q(\cpu.icache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3111),
    .D(_02259_),
    .Q_N(_13124_),
    .Q(\cpu.icache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3112),
    .D(_02260_),
    .Q_N(_13123_),
    .Q(\cpu.icache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3113),
    .D(_02261_),
    .Q_N(_13122_),
    .Q(\cpu.icache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3114),
    .D(_02262_),
    .Q_N(_13121_),
    .Q(\cpu.icache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3115),
    .D(_02263_),
    .Q_N(_13120_),
    .Q(\cpu.icache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3116),
    .D(_02264_),
    .Q_N(_13119_),
    .Q(\cpu.icache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3117),
    .D(_02265_),
    .Q_N(_13118_),
    .Q(\cpu.icache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3118),
    .D(_02266_),
    .Q_N(_13117_),
    .Q(\cpu.icache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3119),
    .D(_02267_),
    .Q_N(_00314_),
    .Q(\cpu.icache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3120),
    .D(_02268_),
    .Q_N(_13116_),
    .Q(\cpu.icache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3121),
    .D(_02269_),
    .Q_N(_00252_),
    .Q(\cpu.icache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3122),
    .D(_02270_),
    .Q_N(_13115_),
    .Q(\cpu.icache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3123),
    .D(_02271_),
    .Q_N(_13114_),
    .Q(\cpu.icache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3124),
    .D(_02272_),
    .Q_N(_13113_),
    .Q(\cpu.icache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3125),
    .D(_02273_),
    .Q_N(_13112_),
    .Q(\cpu.icache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3126),
    .D(_02274_),
    .Q_N(_13111_),
    .Q(\cpu.icache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3127),
    .D(_02275_),
    .Q_N(_13110_),
    .Q(\cpu.icache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3128),
    .D(_02276_),
    .Q_N(_13109_),
    .Q(\cpu.icache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3129),
    .D(_02277_),
    .Q_N(_13108_),
    .Q(\cpu.icache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3130),
    .D(_02278_),
    .Q_N(_13107_),
    .Q(\cpu.icache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3131),
    .D(_02279_),
    .Q_N(_13106_),
    .Q(\cpu.icache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3132),
    .D(_02280_),
    .Q_N(_13105_),
    .Q(\cpu.icache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3133),
    .D(_02281_),
    .Q_N(_13104_),
    .Q(\cpu.icache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3134),
    .D(_02282_),
    .Q_N(_13103_),
    .Q(\cpu.icache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3135),
    .D(_02283_),
    .Q_N(_13102_),
    .Q(\cpu.icache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3136),
    .D(_02284_),
    .Q_N(_13101_),
    .Q(\cpu.icache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3137),
    .D(_02285_),
    .Q_N(_13100_),
    .Q(\cpu.icache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3138),
    .D(_02286_),
    .Q_N(_13099_),
    .Q(\cpu.icache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3139),
    .D(_02287_),
    .Q_N(_13098_),
    .Q(\cpu.icache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3140),
    .D(_02288_),
    .Q_N(_13097_),
    .Q(\cpu.icache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3141),
    .D(_02289_),
    .Q_N(_13096_),
    .Q(\cpu.icache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3142),
    .D(_02290_),
    .Q_N(_13095_),
    .Q(\cpu.icache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3143),
    .D(_02291_),
    .Q_N(_13094_),
    .Q(\cpu.icache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3144),
    .D(_02292_),
    .Q_N(_13093_),
    .Q(\cpu.icache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3145),
    .D(_02293_),
    .Q_N(_13092_),
    .Q(\cpu.icache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3146),
    .D(_02294_),
    .Q_N(_13091_),
    .Q(\cpu.icache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3147),
    .D(_02295_),
    .Q_N(_13090_),
    .Q(\cpu.icache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3148),
    .D(_02296_),
    .Q_N(_13089_),
    .Q(\cpu.icache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3149),
    .D(_02297_),
    .Q_N(_13088_),
    .Q(\cpu.icache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3150),
    .D(_02298_),
    .Q_N(_13087_),
    .Q(\cpu.icache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3151),
    .D(_02299_),
    .Q_N(_13086_),
    .Q(\cpu.icache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3152),
    .D(_02300_),
    .Q_N(_13085_),
    .Q(\cpu.icache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3153),
    .D(_02301_),
    .Q_N(_13084_),
    .Q(\cpu.icache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3154),
    .D(_02302_),
    .Q_N(_13083_),
    .Q(\cpu.icache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3155),
    .D(_02303_),
    .Q_N(_13082_),
    .Q(\cpu.icache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3156),
    .D(_02304_),
    .Q_N(_13081_),
    .Q(\cpu.icache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3157),
    .D(_02305_),
    .Q_N(_13080_),
    .Q(\cpu.icache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3158),
    .D(_02306_),
    .Q_N(_13079_),
    .Q(\cpu.icache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3159),
    .D(_02307_),
    .Q_N(_13078_),
    .Q(\cpu.icache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3160),
    .D(_02308_),
    .Q_N(_13077_),
    .Q(\cpu.icache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3161),
    .D(_02309_),
    .Q_N(_13076_),
    .Q(\cpu.icache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3162),
    .D(_02310_),
    .Q_N(_13075_),
    .Q(\cpu.icache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3163),
    .D(_02311_),
    .Q_N(_13074_),
    .Q(\cpu.icache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3164),
    .D(_02312_),
    .Q_N(_13073_),
    .Q(\cpu.icache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3165),
    .D(_02313_),
    .Q_N(_13072_),
    .Q(\cpu.icache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3166),
    .D(_02314_),
    .Q_N(_13071_),
    .Q(\cpu.icache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3167),
    .D(_02315_),
    .Q_N(_13070_),
    .Q(\cpu.icache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3168),
    .D(_02316_),
    .Q_N(_13069_),
    .Q(\cpu.icache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3169),
    .D(_02317_),
    .Q_N(_13068_),
    .Q(\cpu.icache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3170),
    .D(_02318_),
    .Q_N(_13067_),
    .Q(\cpu.icache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3171),
    .D(_02319_),
    .Q_N(_13066_),
    .Q(\cpu.icache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3172),
    .D(_02320_),
    .Q_N(_13065_),
    .Q(\cpu.icache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3173),
    .D(_02321_),
    .Q_N(_13064_),
    .Q(\cpu.icache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3174),
    .D(_02322_),
    .Q_N(_13063_),
    .Q(\cpu.icache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3175),
    .D(_02323_),
    .Q_N(_13062_),
    .Q(\cpu.icache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3176),
    .D(_02324_),
    .Q_N(_13061_),
    .Q(\cpu.icache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3177),
    .D(_02325_),
    .Q_N(_13060_),
    .Q(\cpu.icache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3178),
    .D(_02326_),
    .Q_N(_13059_),
    .Q(\cpu.icache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3179),
    .D(_02327_),
    .Q_N(_13058_),
    .Q(\cpu.icache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3180),
    .D(_02328_),
    .Q_N(_13057_),
    .Q(\cpu.icache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3181),
    .D(_02329_),
    .Q_N(_13056_),
    .Q(\cpu.icache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3182),
    .D(_02330_),
    .Q_N(_13055_),
    .Q(\cpu.icache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3183),
    .D(_02331_),
    .Q_N(_13054_),
    .Q(\cpu.icache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3184),
    .D(_02332_),
    .Q_N(_13053_),
    .Q(\cpu.icache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3185),
    .D(_02333_),
    .Q_N(_13052_),
    .Q(\cpu.icache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3186),
    .D(_02334_),
    .Q_N(_13051_),
    .Q(\cpu.icache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3187),
    .D(_02335_),
    .Q_N(_13050_),
    .Q(\cpu.icache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3188),
    .D(_02336_),
    .Q_N(_13049_),
    .Q(\cpu.icache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3189),
    .D(_02337_),
    .Q_N(_13048_),
    .Q(\cpu.icache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3190),
    .D(_02338_),
    .Q_N(_13047_),
    .Q(\cpu.icache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3191),
    .D(_02339_),
    .Q_N(_13046_),
    .Q(\cpu.icache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3192),
    .D(_02340_),
    .Q_N(_13045_),
    .Q(\cpu.icache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3193),
    .D(_02341_),
    .Q_N(_13044_),
    .Q(\cpu.icache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3194),
    .D(_02342_),
    .Q_N(_13043_),
    .Q(\cpu.icache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3195),
    .D(_02343_),
    .Q_N(_13042_),
    .Q(\cpu.icache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3196),
    .D(_02344_),
    .Q_N(_13041_),
    .Q(\cpu.icache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3197),
    .D(_02345_),
    .Q_N(_13040_),
    .Q(\cpu.icache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3198),
    .D(_02346_),
    .Q_N(_13039_),
    .Q(\cpu.icache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3199),
    .D(_02347_),
    .Q_N(_13038_),
    .Q(\cpu.icache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3200),
    .D(_02348_),
    .Q_N(_13037_),
    .Q(\cpu.icache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3201),
    .D(_02349_),
    .Q_N(_13036_),
    .Q(\cpu.icache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3202),
    .D(_02350_),
    .Q_N(_13035_),
    .Q(\cpu.icache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3203),
    .D(_02351_),
    .Q_N(_13034_),
    .Q(\cpu.icache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3204),
    .D(_02352_),
    .Q_N(_13033_),
    .Q(\cpu.icache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3205),
    .D(_02353_),
    .Q_N(_13032_),
    .Q(\cpu.icache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3206),
    .D(_02354_),
    .Q_N(_13031_),
    .Q(\cpu.icache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3207),
    .D(_02355_),
    .Q_N(_13030_),
    .Q(\cpu.icache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3208),
    .D(_02356_),
    .Q_N(_13029_),
    .Q(\cpu.icache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3209),
    .D(_02357_),
    .Q_N(_13028_),
    .Q(\cpu.icache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3210),
    .D(_02358_),
    .Q_N(_13027_),
    .Q(\cpu.icache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3211),
    .D(_02359_),
    .Q_N(_13026_),
    .Q(\cpu.icache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3212),
    .D(_02360_),
    .Q_N(_13025_),
    .Q(\cpu.icache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3213),
    .D(_02361_),
    .Q_N(_13024_),
    .Q(\cpu.icache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3214),
    .D(_02362_),
    .Q_N(_13023_),
    .Q(\cpu.icache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3215),
    .D(_02363_),
    .Q_N(_13022_),
    .Q(\cpu.icache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3216),
    .D(_02364_),
    .Q_N(_13021_),
    .Q(\cpu.icache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3217),
    .D(_02365_),
    .Q_N(_13020_),
    .Q(\cpu.icache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3218),
    .D(_02366_),
    .Q_N(_13019_),
    .Q(\cpu.icache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3219),
    .D(_02367_),
    .Q_N(_13018_),
    .Q(\cpu.icache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3220),
    .D(_02368_),
    .Q_N(_13017_),
    .Q(\cpu.icache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3221),
    .D(_02369_),
    .Q_N(_13016_),
    .Q(\cpu.icache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3222),
    .D(_02370_),
    .Q_N(_13015_),
    .Q(\cpu.icache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3223),
    .D(_02371_),
    .Q_N(_13014_),
    .Q(\cpu.icache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3224),
    .D(_02372_),
    .Q_N(_13013_),
    .Q(\cpu.icache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3225),
    .D(_02373_),
    .Q_N(_13012_),
    .Q(\cpu.icache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3226),
    .D(_02374_),
    .Q_N(_13011_),
    .Q(\cpu.icache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3227),
    .D(_02375_),
    .Q_N(_13010_),
    .Q(\cpu.icache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3228),
    .D(_02376_),
    .Q_N(_13009_),
    .Q(\cpu.icache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3229),
    .D(_02377_),
    .Q_N(_13008_),
    .Q(\cpu.icache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3230),
    .D(_02378_),
    .Q_N(_13007_),
    .Q(\cpu.icache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3231),
    .D(_02379_),
    .Q_N(_13006_),
    .Q(\cpu.icache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3232),
    .D(_02380_),
    .Q_N(_13005_),
    .Q(\cpu.icache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3233),
    .D(_02381_),
    .Q_N(_13004_),
    .Q(\cpu.icache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3234),
    .D(_02382_),
    .Q_N(_13003_),
    .Q(\cpu.icache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3235),
    .D(_02383_),
    .Q_N(_13002_),
    .Q(\cpu.icache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3236),
    .D(_02384_),
    .Q_N(_13001_),
    .Q(\cpu.icache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3237),
    .D(_02385_),
    .Q_N(_13000_),
    .Q(\cpu.icache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3238),
    .D(_02386_),
    .Q_N(_12999_),
    .Q(\cpu.icache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3239),
    .D(_02387_),
    .Q_N(_12998_),
    .Q(\cpu.icache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3240),
    .D(_02388_),
    .Q_N(_12997_),
    .Q(\cpu.icache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3241),
    .D(_02389_),
    .Q_N(_12996_),
    .Q(\cpu.icache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3242),
    .D(_02390_),
    .Q_N(_12995_),
    .Q(\cpu.icache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3243),
    .D(_02391_),
    .Q_N(_12994_),
    .Q(\cpu.icache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3244),
    .D(_02392_),
    .Q_N(_12993_),
    .Q(\cpu.icache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3245),
    .D(_02393_),
    .Q_N(_12992_),
    .Q(\cpu.icache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3246),
    .D(_02394_),
    .Q_N(_12991_),
    .Q(\cpu.icache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3247),
    .D(_02395_),
    .Q_N(_12990_),
    .Q(\cpu.icache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3248),
    .D(_02396_),
    .Q_N(_12989_),
    .Q(\cpu.icache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3249),
    .D(_02397_),
    .Q_N(_12988_),
    .Q(\cpu.icache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3250),
    .D(_02398_),
    .Q_N(_12987_),
    .Q(\cpu.icache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3251),
    .D(_02399_),
    .Q_N(_12986_),
    .Q(\cpu.icache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3252),
    .D(_02400_),
    .Q_N(_12985_),
    .Q(\cpu.icache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3253),
    .D(_02401_),
    .Q_N(_12984_),
    .Q(\cpu.icache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3254),
    .D(_02402_),
    .Q_N(_12983_),
    .Q(\cpu.icache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3255),
    .D(_02403_),
    .Q_N(_12982_),
    .Q(\cpu.icache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3256),
    .D(_02404_),
    .Q_N(_12981_),
    .Q(\cpu.icache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3257),
    .D(_02405_),
    .Q_N(_12980_),
    .Q(\cpu.icache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3258),
    .D(_02406_),
    .Q_N(_12979_),
    .Q(\cpu.icache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3259),
    .D(_02407_),
    .Q_N(_12978_),
    .Q(\cpu.icache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3260),
    .D(_02408_),
    .Q_N(_12977_),
    .Q(\cpu.icache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3261),
    .D(_02409_),
    .Q_N(_12976_),
    .Q(\cpu.icache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3262),
    .D(_02410_),
    .Q_N(_12975_),
    .Q(\cpu.icache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3263),
    .D(_02411_),
    .Q_N(_12974_),
    .Q(\cpu.icache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3264),
    .D(_02412_),
    .Q_N(_12973_),
    .Q(\cpu.icache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3265),
    .D(_02413_),
    .Q_N(_12972_),
    .Q(\cpu.icache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3266),
    .D(_02414_),
    .Q_N(_12971_),
    .Q(\cpu.icache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3267),
    .D(_02415_),
    .Q_N(_12970_),
    .Q(\cpu.icache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3268),
    .D(_02416_),
    .Q_N(_12969_),
    .Q(\cpu.icache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3269),
    .D(_02417_),
    .Q_N(_12968_),
    .Q(\cpu.icache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3270),
    .D(_02418_),
    .Q_N(_12967_),
    .Q(\cpu.icache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3271),
    .D(_02419_),
    .Q_N(_12966_),
    .Q(\cpu.icache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3272),
    .D(_02420_),
    .Q_N(_12965_),
    .Q(\cpu.icache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3273),
    .D(_02421_),
    .Q_N(_12964_),
    .Q(\cpu.icache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3274),
    .D(_02422_),
    .Q_N(_12963_),
    .Q(\cpu.icache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net3275),
    .D(_02423_),
    .Q_N(_12962_),
    .Q(\cpu.icache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3276),
    .D(_02424_),
    .Q_N(_12961_),
    .Q(\cpu.icache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3277),
    .D(_02425_),
    .Q_N(_12960_),
    .Q(\cpu.icache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3278),
    .D(_02426_),
    .Q_N(_12959_),
    .Q(\cpu.icache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net3279),
    .D(_02427_),
    .Q_N(_12958_),
    .Q(\cpu.icache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3280),
    .D(_02428_),
    .Q_N(_12957_),
    .Q(\cpu.icache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3281),
    .D(_02429_),
    .Q_N(_12956_),
    .Q(\cpu.icache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3282),
    .D(_02430_),
    .Q_N(_12955_),
    .Q(\cpu.intr.r_clock ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[0]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3283),
    .D(_02431_),
    .Q_N(_12954_),
    .Q(\cpu.intr.r_clock_cmp[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3284),
    .D(_02432_),
    .Q_N(_12953_),
    .Q(\cpu.intr.r_clock_cmp[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3285),
    .D(_02433_),
    .Q_N(_12952_),
    .Q(\cpu.intr.r_clock_cmp[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3286),
    .D(_02434_),
    .Q_N(_12951_),
    .Q(\cpu.intr.r_clock_cmp[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3287),
    .D(_02435_),
    .Q_N(_12950_),
    .Q(\cpu.intr.r_clock_cmp[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3288),
    .D(_02436_),
    .Q_N(_12949_),
    .Q(\cpu.intr.r_clock_cmp[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3289),
    .D(_02437_),
    .Q_N(_12948_),
    .Q(\cpu.intr.r_clock_cmp[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[16]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3290),
    .D(_02438_),
    .Q_N(_12947_),
    .Q(\cpu.intr.r_clock_cmp[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[17]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3291),
    .D(_02439_),
    .Q_N(_12946_),
    .Q(\cpu.intr.r_clock_cmp[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[18]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3292),
    .D(_02440_),
    .Q_N(_12945_),
    .Q(\cpu.intr.r_clock_cmp[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[19]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3293),
    .D(_02441_),
    .Q_N(_12944_),
    .Q(\cpu.intr.r_clock_cmp[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3294),
    .D(_02442_),
    .Q_N(_12943_),
    .Q(\cpu.intr.r_clock_cmp[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[20]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3295),
    .D(_02443_),
    .Q_N(_12942_),
    .Q(\cpu.intr.r_clock_cmp[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[21]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3296),
    .D(_02444_),
    .Q_N(_12941_),
    .Q(\cpu.intr.r_clock_cmp[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[22]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3297),
    .D(_02445_),
    .Q_N(_12940_),
    .Q(\cpu.intr.r_clock_cmp[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[23]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3298),
    .D(_02446_),
    .Q_N(_12939_),
    .Q(\cpu.intr.r_clock_cmp[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[24]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3299),
    .D(_02447_),
    .Q_N(_12938_),
    .Q(\cpu.intr.r_clock_cmp[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[25]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3300),
    .D(_02448_),
    .Q_N(_12937_),
    .Q(\cpu.intr.r_clock_cmp[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[26]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3301),
    .D(_02449_),
    .Q_N(_12936_),
    .Q(\cpu.intr.r_clock_cmp[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[27]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3302),
    .D(_02450_),
    .Q_N(_12935_),
    .Q(\cpu.intr.r_clock_cmp[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[28]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3303),
    .D(_02451_),
    .Q_N(_12934_),
    .Q(\cpu.intr.r_clock_cmp[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[29]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3304),
    .D(_02452_),
    .Q_N(_12933_),
    .Q(\cpu.intr.r_clock_cmp[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3305),
    .D(_02453_),
    .Q_N(_12932_),
    .Q(\cpu.intr.r_clock_cmp[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[30]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3306),
    .D(_02454_),
    .Q_N(_12931_),
    .Q(\cpu.intr.r_clock_cmp[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[31]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3307),
    .D(_02455_),
    .Q_N(_12930_),
    .Q(\cpu.intr.r_clock_cmp[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3308),
    .D(_02456_),
    .Q_N(_12929_),
    .Q(\cpu.intr.r_clock_cmp[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3309),
    .D(_02457_),
    .Q_N(_12928_),
    .Q(\cpu.intr.r_clock_cmp[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3310),
    .D(_02458_),
    .Q_N(_12927_),
    .Q(\cpu.intr.r_clock_cmp[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3311),
    .D(_02459_),
    .Q_N(_12926_),
    .Q(\cpu.intr.r_clock_cmp[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3312),
    .D(_02460_),
    .Q_N(_12925_),
    .Q(\cpu.intr.r_clock_cmp[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3313),
    .D(_02461_),
    .Q_N(_12924_),
    .Q(\cpu.intr.r_clock_cmp[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3314),
    .D(_02462_),
    .Q_N(_14918_),
    .Q(\cpu.intr.r_clock_cmp[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[0]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3315),
    .D(_00036_),
    .Q_N(_00284_),
    .Q(\cpu.intr.r_clock_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[10]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3316),
    .D(_00037_),
    .Q_N(_14919_),
    .Q(\cpu.intr.r_clock_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[11]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3317),
    .D(_00038_),
    .Q_N(_14920_),
    .Q(\cpu.intr.r_clock_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[12]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3318),
    .D(_00039_),
    .Q_N(_14921_),
    .Q(\cpu.intr.r_clock_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[13]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3319),
    .D(_00040_),
    .Q_N(_14922_),
    .Q(\cpu.intr.r_clock_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[14]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3320),
    .D(_00041_),
    .Q_N(_14923_),
    .Q(\cpu.intr.r_clock_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[15]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3321),
    .D(_00042_),
    .Q_N(_12923_),
    .Q(\cpu.intr.r_clock_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[16]$_DFFE_PN_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3322),
    .D(_02463_),
    .Q_N(_12922_),
    .Q(\cpu.intr.r_clock_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[17]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3323),
    .D(_02464_),
    .Q_N(_12921_),
    .Q(\cpu.intr.r_clock_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[18]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3324),
    .D(_02465_),
    .Q_N(_12920_),
    .Q(\cpu.intr.r_clock_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[19]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3325),
    .D(_02466_),
    .Q_N(_14924_),
    .Q(\cpu.intr.r_clock_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[1]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3326),
    .D(_00043_),
    .Q_N(_12919_),
    .Q(\cpu.intr.r_clock_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[20]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3327),
    .D(_02467_),
    .Q_N(_12918_),
    .Q(\cpu.intr.r_clock_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[21]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3328),
    .D(_02468_),
    .Q_N(_12917_),
    .Q(\cpu.intr.r_clock_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[22]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3329),
    .D(_02469_),
    .Q_N(_12916_),
    .Q(\cpu.intr.r_clock_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[23]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3330),
    .D(_02470_),
    .Q_N(_12915_),
    .Q(\cpu.intr.r_clock_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[24]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3331),
    .D(_02471_),
    .Q_N(_12914_),
    .Q(\cpu.intr.r_clock_count[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[25]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3332),
    .D(_02472_),
    .Q_N(_12913_),
    .Q(\cpu.intr.r_clock_count[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[26]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3333),
    .D(_02473_),
    .Q_N(_12912_),
    .Q(\cpu.intr.r_clock_count[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[27]$_DFFE_PN_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3334),
    .D(_02474_),
    .Q_N(_12911_),
    .Q(\cpu.intr.r_clock_count[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[28]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3335),
    .D(_02475_),
    .Q_N(_12910_),
    .Q(\cpu.intr.r_clock_count[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[29]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3336),
    .D(_02476_),
    .Q_N(_14925_),
    .Q(\cpu.intr.r_clock_count[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[2]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3337),
    .D(_00044_),
    .Q_N(_12909_),
    .Q(\cpu.intr.r_clock_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[30]$_DFFE_PN_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3338),
    .D(_02477_),
    .Q_N(_12908_),
    .Q(\cpu.intr.r_clock_count[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[31]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3339),
    .D(_02478_),
    .Q_N(_14926_),
    .Q(\cpu.intr.r_clock_count[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[3]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3340),
    .D(_00045_),
    .Q_N(_14927_),
    .Q(\cpu.intr.r_clock_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[4]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3341),
    .D(_00046_),
    .Q_N(_14928_),
    .Q(\cpu.intr.r_clock_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[5]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3342),
    .D(_00047_),
    .Q_N(_14929_),
    .Q(\cpu.intr.r_clock_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[6]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3343),
    .D(_00048_),
    .Q_N(_14930_),
    .Q(\cpu.intr.r_clock_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[7]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3344),
    .D(_00049_),
    .Q_N(_14931_),
    .Q(\cpu.intr.r_clock_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[8]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3345),
    .D(_00050_),
    .Q_N(_14932_),
    .Q(\cpu.intr.r_clock_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[9]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3346),
    .D(_00051_),
    .Q_N(_12907_),
    .Q(\cpu.intr.r_clock_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3347),
    .D(_02479_),
    .Q_N(_12906_),
    .Q(\cpu.intr.r_enable[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3348),
    .D(_02480_),
    .Q_N(_12905_),
    .Q(\cpu.intr.r_enable[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3349),
    .D(_02481_),
    .Q_N(_12904_),
    .Q(\cpu.intr.r_enable[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3350),
    .D(_02482_),
    .Q_N(_12903_),
    .Q(\cpu.intr.r_enable[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3351),
    .D(_02483_),
    .Q_N(_12902_),
    .Q(\cpu.intr.r_enable[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3352),
    .D(_02484_),
    .Q_N(_12901_),
    .Q(\cpu.intr.r_enable[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3353),
    .D(_02485_),
    .Q_N(_14933_),
    .Q(\cpu.intr.r_timer ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[0]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3354),
    .D(_00055_),
    .Q_N(_00283_),
    .Q(\cpu.intr.r_timer_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[10]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3355),
    .D(_00056_),
    .Q_N(_14934_),
    .Q(\cpu.intr.r_timer_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[11]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3356),
    .D(_00057_),
    .Q_N(_14935_),
    .Q(\cpu.intr.r_timer_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[12]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3357),
    .D(_00058_),
    .Q_N(_14936_),
    .Q(\cpu.intr.r_timer_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[13]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3358),
    .D(_00059_),
    .Q_N(_14937_),
    .Q(\cpu.intr.r_timer_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[14]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3359),
    .D(_00060_),
    .Q_N(_14938_),
    .Q(\cpu.intr.r_timer_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[15]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3360),
    .D(_00061_),
    .Q_N(_14939_),
    .Q(\cpu.intr.r_timer_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[16]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3361),
    .D(_00062_),
    .Q_N(_14940_),
    .Q(\cpu.intr.r_timer_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[17]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3362),
    .D(_00063_),
    .Q_N(_14941_),
    .Q(\cpu.intr.r_timer_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[18]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3363),
    .D(_00064_),
    .Q_N(_14942_),
    .Q(\cpu.intr.r_timer_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[19]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3364),
    .D(_00065_),
    .Q_N(_14943_),
    .Q(\cpu.intr.r_timer_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[1]$_DFF_P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3365),
    .D(_00066_),
    .Q_N(_14944_),
    .Q(\cpu.intr.r_timer_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[20]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3366),
    .D(_00067_),
    .Q_N(_14945_),
    .Q(\cpu.intr.r_timer_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[21]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3367),
    .D(_00068_),
    .Q_N(_14946_),
    .Q(\cpu.intr.r_timer_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[22]$_DFF_P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3368),
    .D(_00069_),
    .Q_N(_14947_),
    .Q(\cpu.intr.r_timer_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[23]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3369),
    .D(_00070_),
    .Q_N(_14948_),
    .Q(\cpu.intr.r_timer_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[2]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3370),
    .D(_00071_),
    .Q_N(_14949_),
    .Q(\cpu.intr.r_timer_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[3]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3371),
    .D(_00072_),
    .Q_N(_14950_),
    .Q(\cpu.intr.r_timer_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[4]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3372),
    .D(_00073_),
    .Q_N(_14951_),
    .Q(\cpu.intr.r_timer_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[5]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3373),
    .D(_00074_),
    .Q_N(_14952_),
    .Q(\cpu.intr.r_timer_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[6]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3374),
    .D(_00075_),
    .Q_N(_14953_),
    .Q(\cpu.intr.r_timer_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[7]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3375),
    .D(_00076_),
    .Q_N(_14954_),
    .Q(\cpu.intr.r_timer_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[8]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3376),
    .D(_00077_),
    .Q_N(_14955_),
    .Q(\cpu.intr.r_timer_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[9]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3377),
    .D(_00078_),
    .Q_N(_12900_),
    .Q(\cpu.intr.r_timer_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[0]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3378),
    .D(_02486_),
    .Q_N(_12899_),
    .Q(\cpu.intr.r_timer_reload[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[10]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3379),
    .D(_02487_),
    .Q_N(_12898_),
    .Q(\cpu.intr.r_timer_reload[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[11]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3380),
    .D(_02488_),
    .Q_N(_12897_),
    .Q(\cpu.intr.r_timer_reload[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[12]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3381),
    .D(_02489_),
    .Q_N(_12896_),
    .Q(\cpu.intr.r_timer_reload[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[13]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3382),
    .D(_02490_),
    .Q_N(_12895_),
    .Q(\cpu.intr.r_timer_reload[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[14]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3383),
    .D(_02491_),
    .Q_N(_12894_),
    .Q(\cpu.intr.r_timer_reload[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[15]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3384),
    .D(_02492_),
    .Q_N(_12893_),
    .Q(\cpu.intr.r_timer_reload[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[16]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3385),
    .D(_02493_),
    .Q_N(_12892_),
    .Q(\cpu.intr.r_timer_reload[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[17]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3386),
    .D(_02494_),
    .Q_N(_12891_),
    .Q(\cpu.intr.r_timer_reload[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[18]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3387),
    .D(_02495_),
    .Q_N(_12890_),
    .Q(\cpu.intr.r_timer_reload[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[19]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3388),
    .D(_02496_),
    .Q_N(_12889_),
    .Q(\cpu.intr.r_timer_reload[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[1]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3389),
    .D(_02497_),
    .Q_N(_12888_),
    .Q(\cpu.intr.r_timer_reload[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[20]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3390),
    .D(_02498_),
    .Q_N(_12887_),
    .Q(\cpu.intr.r_timer_reload[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[21]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3391),
    .D(_02499_),
    .Q_N(_12886_),
    .Q(\cpu.intr.r_timer_reload[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[22]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3392),
    .D(_02500_),
    .Q_N(_12885_),
    .Q(\cpu.intr.r_timer_reload[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[23]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3393),
    .D(_02501_),
    .Q_N(_12884_),
    .Q(\cpu.intr.r_timer_reload[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3394),
    .D(_02502_),
    .Q_N(_12883_),
    .Q(\cpu.intr.r_timer_reload[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3395),
    .D(_02503_),
    .Q_N(_12882_),
    .Q(\cpu.intr.r_timer_reload[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[4]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3396),
    .D(_02504_),
    .Q_N(_12881_),
    .Q(\cpu.intr.r_timer_reload[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[5]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3397),
    .D(_02505_),
    .Q_N(_12880_),
    .Q(\cpu.intr.r_timer_reload[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[6]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3398),
    .D(_02506_),
    .Q_N(_12879_),
    .Q(\cpu.intr.r_timer_reload[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[7]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3399),
    .D(_02507_),
    .Q_N(_12878_),
    .Q(\cpu.intr.r_timer_reload[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[8]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3400),
    .D(_02508_),
    .Q_N(_12877_),
    .Q(\cpu.intr.r_timer_reload[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[9]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3401),
    .D(_02509_),
    .Q_N(_12876_),
    .Q(\cpu.intr.r_timer_reload[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3402),
    .D(_02510_),
    .Q_N(_00178_),
    .Q(\cpu.qspi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net3403),
    .D(_02511_),
    .Q_N(_12875_),
    .Q(\cpu.qspi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net3404),
    .D(_02512_),
    .Q_N(_00179_),
    .Q(\cpu.qspi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net3405),
    .D(_02513_),
    .Q_N(_12874_),
    .Q(\cpu.qspi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net3406),
    .D(_02514_),
    .Q_N(_00250_),
    .Q(\cpu.qspi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3407),
    .D(_02515_),
    .Q_N(_12873_),
    .Q(net19));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3408),
    .D(_02516_),
    .Q_N(_12872_),
    .Q(net20));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3409),
    .D(_02517_),
    .Q_N(_12871_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_ind$_SDFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3410),
    .D(_02518_),
    .Q_N(_12870_),
    .Q(\cpu.qspi.r_ind ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3411),
    .D(_02519_),
    .Q_N(_12869_),
    .Q(\cpu.qspi.r_mask[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3412),
    .D(_02520_),
    .Q_N(_12868_),
    .Q(\cpu.qspi.r_mask[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3413),
    .D(_02521_),
    .Q_N(_12867_),
    .Q(\cpu.qspi.r_mask[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3414),
    .D(_02522_),
    .Q_N(_12866_),
    .Q(\cpu.qspi.r_quad[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3415),
    .D(_02523_),
    .Q_N(_12865_),
    .Q(\cpu.qspi.r_quad[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3416),
    .D(_02524_),
    .Q_N(_12864_),
    .Q(\cpu.qspi.r_quad[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net3417),
    .D(_02525_),
    .Q_N(_12863_),
    .Q(\cpu.qspi.r_read_delay[0][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3418),
    .D(_02526_),
    .Q_N(_12862_),
    .Q(\cpu.qspi.r_read_delay[0][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3419),
    .D(_02527_),
    .Q_N(_12861_),
    .Q(\cpu.qspi.r_read_delay[0][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3420),
    .D(_02528_),
    .Q_N(_12860_),
    .Q(\cpu.qspi.r_read_delay[0][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net3421),
    .D(_02529_),
    .Q_N(_12859_),
    .Q(\cpu.qspi.r_read_delay[1][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net3422),
    .D(_02530_),
    .Q_N(_12858_),
    .Q(\cpu.qspi.r_read_delay[1][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3423),
    .D(_02531_),
    .Q_N(_12857_),
    .Q(\cpu.qspi.r_read_delay[1][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3424),
    .D(_02532_),
    .Q_N(_12856_),
    .Q(\cpu.qspi.r_read_delay[1][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3425),
    .D(_02533_),
    .Q_N(_12855_),
    .Q(\cpu.qspi.r_read_delay[2][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net3426),
    .D(_02534_),
    .Q_N(_12854_),
    .Q(\cpu.qspi.r_read_delay[2][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net3427),
    .D(_02535_),
    .Q_N(_12853_),
    .Q(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3428),
    .D(_02536_),
    .Q_N(_12852_),
    .Q(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3429),
    .D(_02537_),
    .Q_N(_12851_),
    .Q(\cpu.qspi.r_rom_mode[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3430),
    .D(_02538_),
    .Q_N(_14956_),
    .Q(\cpu.qspi.r_rom_mode[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rstrobe_d$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net3431),
    .D(\cpu.qspi.c_rstrobe_d ),
    .Q_N(_14957_),
    .Q(\cpu.d_rstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3432),
    .D(_00021_),
    .Q_N(_00275_),
    .Q(\cpu.qspi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[10]$_DFF_P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net3433),
    .D(_00008_),
    .Q_N(_14958_),
    .Q(\cpu.qspi.r_state[10] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[11]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3434),
    .D(_00022_),
    .Q_N(_14959_),
    .Q(\cpu.qspi.r_state[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[12]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3435),
    .D(_00023_),
    .Q_N(_14960_),
    .Q(\cpu.qspi.r_state[12] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[13]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net3436),
    .D(_00009_),
    .Q_N(_14961_),
    .Q(\cpu.qspi.r_state[13] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[14]$_DFF_P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net3437),
    .D(_00024_),
    .Q_N(_14962_),
    .Q(\cpu.qspi.r_state[14] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[15]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net3438),
    .D(_00010_),
    .Q_N(_14963_),
    .Q(\cpu.qspi.r_state[15] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[16]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3439),
    .D(_00025_),
    .Q_N(_14964_),
    .Q(\cpu.qspi.r_state[16] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[17]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3440),
    .D(_00026_),
    .Q_N(_14965_),
    .Q(\cpu.qspi.r_state[17] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3441),
    .D(_00001_),
    .Q_N(_14966_),
    .Q(\cpu.qspi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3442),
    .D(_00027_),
    .Q_N(_14967_),
    .Q(\cpu.qspi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net3443),
    .D(_00002_),
    .Q_N(_14968_),
    .Q(\cpu.qspi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3444),
    .D(_00028_),
    .Q_N(_14969_),
    .Q(\cpu.qspi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3445),
    .D(_00003_),
    .Q_N(_14970_),
    .Q(\cpu.qspi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net3446),
    .D(_00004_),
    .Q_N(_14971_),
    .Q(\cpu.qspi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[7]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3447),
    .D(_00005_),
    .Q_N(_14972_),
    .Q(\cpu.qspi.r_state[7] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[8]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net3448),
    .D(_00006_),
    .Q_N(_00180_),
    .Q(\cpu.qspi.r_state[8] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[9]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3449),
    .D(_00007_),
    .Q_N(_12850_),
    .Q(\cpu.qspi.r_state[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3450),
    .D(_02539_),
    .Q_N(_12849_),
    .Q(net3));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3451),
    .D(_02540_),
    .Q_N(_12848_),
    .Q(net6));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3452),
    .D(_02541_),
    .Q_N(_12847_),
    .Q(net11));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3453),
    .D(_02542_),
    .Q_N(_12846_),
    .Q(net12));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3454),
    .D(_02543_),
    .Q_N(_12845_),
    .Q(net13));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3455),
    .D(_02544_),
    .Q_N(_14973_),
    .Q(net14));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_d$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net3456),
    .D(\cpu.qspi.c_wstrobe_d ),
    .Q_N(_14974_),
    .Q(\cpu.d_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_i$_DFF_P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3457),
    .D(\cpu.qspi.c_wstrobe_i ),
    .Q_N(_00251_),
    .Q(\cpu.i_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.r_clk_invert$_DFFE_PN_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3458),
    .D(_02545_),
    .Q_N(_12844_),
    .Q(\cpu.r_clk_invert ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3459),
    .D(_02546_),
    .Q_N(_12843_),
    .Q(\cpu.spi.r_bits[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3460),
    .D(_02547_),
    .Q_N(_12842_),
    .Q(\cpu.spi.r_bits[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3461),
    .D(_02548_),
    .Q_N(_12841_),
    .Q(\cpu.spi.r_bits[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3462),
    .D(_02549_),
    .Q_N(_00312_),
    .Q(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3463),
    .D(_02550_),
    .Q_N(_00095_),
    .Q(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3464),
    .D(_02551_),
    .Q_N(_00105_),
    .Q(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3465),
    .D(_02552_),
    .Q_N(_00115_),
    .Q(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3466),
    .D(_02553_),
    .Q_N(_00126_),
    .Q(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3467),
    .D(_02554_),
    .Q_N(_00133_),
    .Q(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3468),
    .D(_02555_),
    .Q_N(_00145_),
    .Q(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3469),
    .D(_02556_),
    .Q_N(_00157_),
    .Q(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3470),
    .D(_02557_),
    .Q_N(_00311_),
    .Q(\cpu.spi.r_clk_count[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3471),
    .D(_02558_),
    .Q_N(_00094_),
    .Q(\cpu.spi.r_clk_count[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3472),
    .D(_02559_),
    .Q_N(_00104_),
    .Q(\cpu.spi.r_clk_count[1][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3473),
    .D(_02560_),
    .Q_N(_00114_),
    .Q(\cpu.spi.r_clk_count[1][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3474),
    .D(_02561_),
    .Q_N(_00125_),
    .Q(\cpu.spi.r_clk_count[1][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3475),
    .D(_02562_),
    .Q_N(_00132_),
    .Q(\cpu.spi.r_clk_count[1][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3476),
    .D(_02563_),
    .Q_N(_00144_),
    .Q(\cpu.spi.r_clk_count[1][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3477),
    .D(_02564_),
    .Q_N(_00156_),
    .Q(\cpu.spi.r_clk_count[1][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3478),
    .D(_02565_),
    .Q_N(_12840_),
    .Q(\cpu.spi.r_clk_count[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3479),
    .D(_02566_),
    .Q_N(_12839_),
    .Q(\cpu.spi.r_clk_count[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3480),
    .D(_02567_),
    .Q_N(_12838_),
    .Q(\cpu.spi.r_clk_count[2][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3481),
    .D(_02568_),
    .Q_N(_12837_),
    .Q(\cpu.spi.r_clk_count[2][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3482),
    .D(_02569_),
    .Q_N(_12836_),
    .Q(\cpu.spi.r_clk_count[2][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3483),
    .D(_02570_),
    .Q_N(_12835_),
    .Q(\cpu.spi.r_clk_count[2][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3484),
    .D(_02571_),
    .Q_N(_12834_),
    .Q(\cpu.spi.r_clk_count[2][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3485),
    .D(_02572_),
    .Q_N(_12833_),
    .Q(\cpu.spi.r_clk_count[2][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3486),
    .D(_02573_),
    .Q_N(_12832_),
    .Q(\cpu.spi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3487),
    .D(_02574_),
    .Q_N(_12831_),
    .Q(\cpu.spi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3488),
    .D(_02575_),
    .Q_N(_12830_),
    .Q(\cpu.spi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3489),
    .D(_02576_),
    .Q_N(_12829_),
    .Q(\cpu.spi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3490),
    .D(_02577_),
    .Q_N(_12828_),
    .Q(\cpu.spi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3491),
    .D(_02578_),
    .Q_N(_12827_),
    .Q(\cpu.spi.r_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3492),
    .D(_02579_),
    .Q_N(_12826_),
    .Q(\cpu.spi.r_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3493),
    .D(_02580_),
    .Q_N(_12825_),
    .Q(\cpu.spi.r_count[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3494),
    .D(_02581_),
    .Q_N(_12824_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3495),
    .D(_02582_),
    .Q_N(_12823_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3496),
    .D(_02583_),
    .Q_N(_12822_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[8] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3497),
    .D(_02584_),
    .Q_N(_12821_),
    .Q(\cpu.spi.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3498),
    .D(_02585_),
    .Q_N(_12820_),
    .Q(\cpu.spi.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3499),
    .D(_02586_),
    .Q_N(_12819_),
    .Q(\cpu.spi.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3500),
    .D(_02587_),
    .Q_N(_12818_),
    .Q(\cpu.spi.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3501),
    .D(_02588_),
    .Q_N(_12817_),
    .Q(\cpu.spi.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3502),
    .D(_02589_),
    .Q_N(_12816_),
    .Q(\cpu.spi.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3503),
    .D(_02590_),
    .Q_N(_12815_),
    .Q(\cpu.spi.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3504),
    .D(_02591_),
    .Q_N(_00220_),
    .Q(\cpu.spi.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_interrupt$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3505),
    .D(_02592_),
    .Q_N(_12814_),
    .Q(\cpu.intr.spi_intr ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3506),
    .D(_02593_),
    .Q_N(_00222_),
    .Q(\cpu.spi.r_mode[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3507),
    .D(_02594_),
    .Q_N(_12813_),
    .Q(\cpu.spi.r_mode[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3508),
    .D(_02595_),
    .Q_N(_12812_),
    .Q(\cpu.spi.r_mode[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3509),
    .D(_02596_),
    .Q_N(_12811_),
    .Q(\cpu.spi.r_mode[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3510),
    .D(_02597_),
    .Q_N(_12810_),
    .Q(\cpu.spi.r_mode[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3511),
    .D(_02598_),
    .Q_N(_12809_),
    .Q(\cpu.spi.r_mode[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3512),
    .D(_02599_),
    .Q_N(_12808_),
    .Q(\cpu.spi.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3513),
    .D(_02600_),
    .Q_N(_12807_),
    .Q(\cpu.spi.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3514),
    .D(_02601_),
    .Q_N(_12806_),
    .Q(\cpu.spi.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3515),
    .D(_02602_),
    .Q_N(_12805_),
    .Q(\cpu.spi.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3516),
    .D(_02603_),
    .Q_N(_12804_),
    .Q(\cpu.spi.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3517),
    .D(_02604_),
    .Q_N(_12803_),
    .Q(\cpu.spi.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3518),
    .D(_02605_),
    .Q_N(_12802_),
    .Q(\cpu.spi.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3519),
    .D(_02606_),
    .Q_N(_12801_),
    .Q(\cpu.spi.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_ready$_SDFFE_PN1P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3520),
    .D(_02607_),
    .Q_N(_12800_),
    .Q(\cpu.spi.r_ready ));
 sg13g2_dfrbp_1 \cpu.spi.r_searching$_SDFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3521),
    .D(_02608_),
    .Q_N(_00219_),
    .Q(\cpu.spi.r_searching ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[0]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3522),
    .D(_02609_),
    .Q_N(_12799_),
    .Q(\cpu.spi.r_sel[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[1]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3523),
    .D(_02610_),
    .Q_N(_12798_),
    .Q(\cpu.spi.r_sel[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3524),
    .D(_02611_),
    .Q_N(_00280_),
    .Q(\cpu.spi.r_src[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3525),
    .D(_02612_),
    .Q_N(_00281_),
    .Q(\cpu.spi.r_src[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3526),
    .D(_02613_),
    .Q_N(_14975_),
    .Q(\cpu.spi.r_src[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3527),
    .D(_00029_),
    .Q_N(_14976_),
    .Q(\cpu.spi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3528),
    .D(_00030_),
    .Q_N(_00223_),
    .Q(\cpu.spi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3529),
    .D(_00031_),
    .Q_N(_14977_),
    .Q(\cpu.spi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3530),
    .D(_00032_),
    .Q_N(_14978_),
    .Q(\cpu.spi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3531),
    .D(_00033_),
    .Q_N(_00276_),
    .Q(\cpu.spi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3532),
    .D(_00034_),
    .Q_N(_14979_),
    .Q(\cpu.spi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3533),
    .D(_00035_),
    .Q_N(_00224_),
    .Q(\cpu.spi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3534),
    .D(_02614_),
    .Q_N(_12797_),
    .Q(\cpu.spi.r_timeout[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3535),
    .D(_02615_),
    .Q_N(_12796_),
    .Q(\cpu.spi.r_timeout[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3536),
    .D(_02616_),
    .Q_N(_12795_),
    .Q(\cpu.spi.r_timeout[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[3]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3537),
    .D(_02617_),
    .Q_N(_12794_),
    .Q(\cpu.spi.r_timeout[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[4]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3538),
    .D(_02618_),
    .Q_N(_12793_),
    .Q(\cpu.spi.r_timeout[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[5]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3539),
    .D(_02619_),
    .Q_N(_12792_),
    .Q(\cpu.spi.r_timeout[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[6]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3540),
    .D(_02620_),
    .Q_N(_12791_),
    .Q(\cpu.spi.r_timeout[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[7]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3541),
    .D(_02621_),
    .Q_N(_12790_),
    .Q(\cpu.spi.r_timeout[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3542),
    .D(_02622_),
    .Q_N(_00282_),
    .Q(\cpu.spi.r_timeout_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3543),
    .D(_02623_),
    .Q_N(_12789_),
    .Q(\cpu.spi.r_timeout_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3544),
    .D(_02624_),
    .Q_N(_12788_),
    .Q(\cpu.spi.r_timeout_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3545),
    .D(_02625_),
    .Q_N(_12787_),
    .Q(\cpu.spi.r_timeout_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3546),
    .D(_02626_),
    .Q_N(_12786_),
    .Q(\cpu.spi.r_timeout_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3547),
    .D(_02627_),
    .Q_N(_12785_),
    .Q(\cpu.spi.r_timeout_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3548),
    .D(_02628_),
    .Q_N(_12784_),
    .Q(\cpu.spi.r_timeout_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3549),
    .D(_02629_),
    .Q_N(_14980_),
    .Q(\cpu.spi.r_timeout_count[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[0]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3550),
    .D(_00079_),
    .Q_N(_00277_),
    .Q(\cpu.uart.r_div[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[10]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3551),
    .D(_00080_),
    .Q_N(_14981_),
    .Q(\cpu.uart.r_div[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[11]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3552),
    .D(_00081_),
    .Q_N(_14982_),
    .Q(\cpu.uart.r_div[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[1]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3553),
    .D(_00082_),
    .Q_N(_14983_),
    .Q(\cpu.uart.r_div[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[2]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3554),
    .D(_00083_),
    .Q_N(_14984_),
    .Q(\cpu.uart.r_div[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[3]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3555),
    .D(_00084_),
    .Q_N(_14985_),
    .Q(\cpu.uart.r_div[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[4]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3556),
    .D(_00085_),
    .Q_N(_14986_),
    .Q(\cpu.uart.r_div[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[5]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3557),
    .D(_00086_),
    .Q_N(_14987_),
    .Q(\cpu.uart.r_div[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[6]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3558),
    .D(_00087_),
    .Q_N(_14988_),
    .Q(\cpu.uart.r_div[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[7]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3559),
    .D(_00088_),
    .Q_N(_14989_),
    .Q(\cpu.uart.r_div[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[8]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3560),
    .D(_00089_),
    .Q_N(_14990_),
    .Q(\cpu.uart.r_div[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[9]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3561),
    .D(_00090_),
    .Q_N(_12783_),
    .Q(\cpu.uart.r_div[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3562),
    .D(_02630_),
    .Q_N(_12782_),
    .Q(\cpu.uart.r_div_value[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3563),
    .D(_02631_),
    .Q_N(_12781_),
    .Q(\cpu.uart.r_div_value[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3564),
    .D(_02632_),
    .Q_N(_12780_),
    .Q(\cpu.uart.r_div_value[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3565),
    .D(_02633_),
    .Q_N(_12779_),
    .Q(\cpu.uart.r_div_value[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3566),
    .D(_02634_),
    .Q_N(_12778_),
    .Q(\cpu.uart.r_div_value[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3567),
    .D(_02635_),
    .Q_N(_12777_),
    .Q(\cpu.uart.r_div_value[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3568),
    .D(_02636_),
    .Q_N(_12776_),
    .Q(\cpu.uart.r_div_value[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3569),
    .D(_02637_),
    .Q_N(_12775_),
    .Q(\cpu.uart.r_div_value[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3570),
    .D(_02638_),
    .Q_N(_12774_),
    .Q(\cpu.uart.r_div_value[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3571),
    .D(_02639_),
    .Q_N(_12773_),
    .Q(\cpu.uart.r_div_value[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3572),
    .D(_02640_),
    .Q_N(_12772_),
    .Q(\cpu.uart.r_div_value[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3573),
    .D(_02641_),
    .Q_N(_12771_),
    .Q(\cpu.uart.r_div_value[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[0]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3574),
    .D(_02642_),
    .Q_N(_12770_),
    .Q(\cpu.uart.r_ib[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[1]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3575),
    .D(_02643_),
    .Q_N(_12769_),
    .Q(\cpu.uart.r_ib[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3576),
    .D(_02644_),
    .Q_N(_12768_),
    .Q(\cpu.uart.r_ib[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[3]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3577),
    .D(_02645_),
    .Q_N(_12767_),
    .Q(\cpu.uart.r_ib[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[4]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3578),
    .D(_02646_),
    .Q_N(_12766_),
    .Q(\cpu.uart.r_ib[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3579),
    .D(_02647_),
    .Q_N(_12765_),
    .Q(\cpu.uart.r_ib[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[6]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3580),
    .D(_02648_),
    .Q_N(_12764_),
    .Q(\cpu.uart.r_ib[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3581),
    .D(_02649_),
    .Q_N(_12763_),
    .Q(\cpu.uart.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3582),
    .D(_02650_),
    .Q_N(_12762_),
    .Q(\cpu.uart.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3583),
    .D(_02651_),
    .Q_N(_12761_),
    .Q(\cpu.uart.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3584),
    .D(_02652_),
    .Q_N(_12760_),
    .Q(\cpu.uart.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3585),
    .D(_02653_),
    .Q_N(_12759_),
    .Q(\cpu.uart.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3586),
    .D(_02654_),
    .Q_N(_12758_),
    .Q(\cpu.uart.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3587),
    .D(_02655_),
    .Q_N(_12757_),
    .Q(\cpu.uart.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3588),
    .D(_02656_),
    .Q_N(_12756_),
    .Q(\cpu.uart.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3589),
    .D(_02657_),
    .Q_N(_12755_),
    .Q(\cpu.uart.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3590),
    .D(_02658_),
    .Q_N(_12754_),
    .Q(\cpu.uart.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3591),
    .D(_02659_),
    .Q_N(_12753_),
    .Q(\cpu.uart.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3592),
    .D(_02660_),
    .Q_N(_12752_),
    .Q(\cpu.uart.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3593),
    .D(_02661_),
    .Q_N(_12751_),
    .Q(\cpu.uart.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3594),
    .D(_02662_),
    .Q_N(_12750_),
    .Q(\cpu.uart.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3595),
    .D(_02663_),
    .Q_N(_12749_),
    .Q(\cpu.uart.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3596),
    .D(_02664_),
    .Q_N(_14991_),
    .Q(\cpu.uart.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_r$_DFF_P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3597),
    .D(\cpu.gpio.uart_rx ),
    .Q_N(_12748_),
    .Q(\cpu.uart.r_r ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3598),
    .D(_02665_),
    .Q_N(_12747_),
    .Q(\cpu.uart.r_r_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3599),
    .D(_02666_),
    .Q_N(_12746_),
    .Q(\cpu.uart.r_r_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3600),
    .D(_02667_),
    .Q_N(_12745_),
    .Q(\cpu.uart.r_rcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3601),
    .D(_02668_),
    .Q_N(_12744_),
    .Q(\cpu.uart.r_rcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3602),
    .D(_02669_),
    .Q_N(_12743_),
    .Q(\cpu.uart.r_rstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3603),
    .D(_02670_),
    .Q_N(_12742_),
    .Q(\cpu.uart.r_rstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3604),
    .D(_02671_),
    .Q_N(_12741_),
    .Q(\cpu.uart.r_rstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3605),
    .D(_02672_),
    .Q_N(_12740_),
    .Q(\cpu.uart.r_rstate[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3606),
    .D(_02673_),
    .Q_N(_12739_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3607),
    .D(_02674_),
    .Q_N(_12738_),
    .Q(\cpu.uart.r_x_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3608),
    .D(_02675_),
    .Q_N(_00278_),
    .Q(\cpu.uart.r_x_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3609),
    .D(_02676_),
    .Q_N(_12737_),
    .Q(\cpu.uart.r_xcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3610),
    .D(_02677_),
    .Q_N(_12736_),
    .Q(\cpu.uart.r_xcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3611),
    .D(_02678_),
    .Q_N(_12735_),
    .Q(\cpu.uart.r_xstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3612),
    .D(_02679_),
    .Q_N(_12734_),
    .Q(\cpu.uart.r_xstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3613),
    .D(_02680_),
    .Q_N(_12733_),
    .Q(\cpu.uart.r_xstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3614),
    .D(_02681_),
    .Q_N(_14992_),
    .Q(\cpu.uart.r_xstate[3] ));
 sg13g2_dfrbp_1 \r_reset$_DFF_P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net3615),
    .D(_00000_),
    .Q_N(_12732_),
    .Q(r_reset));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_oe[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_oe[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_oe[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_oe[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[7]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[0]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[1]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[2]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[3]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[4]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[5]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[6]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout27 (.A(_03872_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_11481_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_06680_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_07063_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_03897_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_02909_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_02866_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_02803_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_02771_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_02751_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_02743_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_02687_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_12703_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_12681_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_12671_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_12593_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_12572_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_12564_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_12519_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_12475_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_12410_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_12378_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_12358_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_12350_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_12293_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_12254_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_12228_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_12218_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_12102_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_12043_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_12020_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_11727_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_07859_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_06990_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_04268_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_02885_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_02858_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_12627_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_12494_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_12467_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_12155_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_10020_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_10009_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_10008_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_07157_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_06947_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_06347_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_06339_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_06336_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_06331_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_05310_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_04885_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_09017_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_07156_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_04345_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_04141_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_03635_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_11508_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_11500_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_10141_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_10118_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_09863_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_09016_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_07177_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_07158_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_06774_),
    .X(net92));
 sg13g2_buf_4 fanout93 (.X(net93),
    .A(_06669_));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(_06665_));
 sg13g2_buf_4 fanout95 (.X(net95),
    .A(_06662_));
 sg13g2_buf_2 fanout96 (.A(_04255_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_03345_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_03233_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_11507_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_10140_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_10137_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_10127_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_10113_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_10064_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_09918_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_09892_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_09104_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_08093_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_07842_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_07808_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_07641_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_07537_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_06770_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_03644_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_11548_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_10136_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_09346_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_09103_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_09000_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_07374_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_05416_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_04364_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_04326_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_04324_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_04322_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_04319_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_04316_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_04301_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_04214_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_04196_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_04189_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_04187_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_04180_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_04163_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_04155_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_03774_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_03752_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_03643_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_03204_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_03181_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_11833_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_09850_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_09354_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_09175_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_07586_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_07543_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_07542_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_07385_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_07384_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_05694_),
    .X(net150));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(_05334_));
 sg13g2_buf_2 fanout152 (.A(_05309_),
    .X(net152));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(_05232_));
 sg13g2_buf_2 fanout154 (.A(_04321_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_04307_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_04208_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_04200_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_04195_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_04175_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_04162_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_04152_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_04149_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_03803_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_03757_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_03753_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_03751_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_03682_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_11614_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_11442_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_10330_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_10003_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_08381_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_07564_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_07561_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_07426_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_07413_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_07367_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_07035_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_04192_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_04174_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_04161_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_04159_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_03139_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_03063_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_03052_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_03047_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_03022_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_11731_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_11719_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_11667_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_11537_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_11470_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_11393_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_11379_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_09893_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_05229_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_04860_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_04231_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_04158_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_03640_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_03334_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_03145_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_03141_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_03138_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_03061_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_03054_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_03053_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_03051_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_03046_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_03044_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_11767_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_11411_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_11400_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_11376_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_11372_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_11295_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_11227_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_09933_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_09914_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_09904_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_09127_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_09093_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_08379_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_06564_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_04230_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_04138_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_03360_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_03199_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_03149_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_03137_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_03122_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_03068_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_03048_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_03045_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_03043_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_03029_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_11594_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_11551_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_11301_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_11122_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_10665_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_09932_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_09913_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_09882_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_09865_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_09162_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_06563_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_06562_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_06451_),
    .X(net249));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(_06313_));
 sg13g2_buf_2 fanout251 (.A(_06278_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_06243_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_06236_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_06202_),
    .X(net254));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(_06173_));
 sg13g2_buf_4 fanout256 (.X(net256),
    .A(_06166_));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(_06158_));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(_06132_));
 sg13g2_buf_2 fanout259 (.A(_06095_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_06086_),
    .X(net260));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(_06063_));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(_06054_));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(_06032_));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(_06022_));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(_06018_));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(_06013_));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(_06009_));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(_05990_));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(_05976_));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(_05973_));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(_05969_));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(_05962_));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(_05944_));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(_05926_));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(_05921_));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(_05916_));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(_05890_));
 sg13g2_buf_2 fanout278 (.A(_04270_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_03915_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_03654_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_03638_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_03039_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_03038_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_03023_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_11563_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_11510_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_11332_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_09097_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_09091_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_09071_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_09044_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_09040_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_09036_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_08616_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_08460_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_06547_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_06545_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_06544_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_06299_),
    .X(net299));
 sg13g2_buf_4 fanout300 (.X(net300),
    .A(_06292_));
 sg13g2_buf_2 fanout301 (.A(_06285_),
    .X(net301));
 sg13g2_buf_4 fanout302 (.X(net302),
    .A(_06271_));
 sg13g2_buf_2 fanout303 (.A(_06264_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_06224_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_06216_),
    .X(net305));
 sg13g2_buf_4 fanout306 (.X(net306),
    .A(_06187_));
 sg13g2_buf_4 fanout307 (.X(net307),
    .A(_06151_));
 sg13g2_buf_4 fanout308 (.X(net308),
    .A(_06140_));
 sg13g2_buf_2 fanout309 (.A(_06110_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_06102_),
    .X(net310));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(_06078_));
 sg13g2_buf_4 fanout312 (.X(net312),
    .A(_06071_));
 sg13g2_buf_4 fanout313 (.X(net313),
    .A(_06051_));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(_06048_));
 sg13g2_buf_4 fanout315 (.X(net315),
    .A(_06043_));
 sg13g2_buf_4 fanout316 (.X(net316),
    .A(_06037_));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(_06028_));
 sg13g2_buf_4 fanout318 (.X(net318),
    .A(_06025_));
 sg13g2_buf_4 fanout319 (.X(net319),
    .A(_06000_));
 sg13g2_buf_4 fanout320 (.X(net320),
    .A(_05996_));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(_05985_));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(_05980_));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(_05958_));
 sg13g2_buf_4 fanout324 (.X(net324),
    .A(_05948_));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(_05939_));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(_05932_));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(_05909_));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(_05899_));
 sg13g2_buf_2 fanout329 (.A(_05181_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_04257_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_04246_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_03903_),
    .X(net332));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(_03003_));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(_03002_));
 sg13g2_buf_2 fanout335 (.A(_09997_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_08459_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_07475_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_06645_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_06643_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_06642_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_06625_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_06623_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_06622_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_06605_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_06603_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_06602_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_06585_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_06583_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_06582_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_06527_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_06525_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_06524_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_06504_),
    .X(net353));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(_06306_));
 sg13g2_buf_2 fanout355 (.A(_06257_),
    .X(net355));
 sg13g2_buf_4 fanout356 (.X(net356),
    .A(_06250_));
 sg13g2_buf_2 fanout357 (.A(_06195_),
    .X(net357));
 sg13g2_buf_4 fanout358 (.X(net358),
    .A(_06180_));
 sg13g2_buf_2 fanout359 (.A(_06118_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_05180_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_04978_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_04910_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_03921_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_03910_),
    .X(net364));
 sg13g2_buf_4 fanout365 (.X(net365),
    .A(_03017_));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(_03015_));
 sg13g2_buf_2 fanout367 (.A(_12412_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_12181_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_12178_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_12171_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_12165_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_12161_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_10124_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_09996_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_09799_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_09776_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_09754_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_09640_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_09553_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_09513_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_09489_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_09464_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_08681_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_08648_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_06503_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_06502_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_06388_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_05436_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_05435_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_05382_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_05346_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_05336_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_05213_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_05209_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_05028_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_04997_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_04994_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_04989_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_04977_),
    .X(net399));
 sg13g2_buf_4 fanout400 (.X(net400),
    .A(_03014_));
 sg13g2_buf_4 fanout401 (.X(net401),
    .A(_03013_));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(_03005_));
 sg13g2_buf_4 fanout403 (.X(net403),
    .A(_03004_));
 sg13g2_buf_4 fanout404 (.X(net404),
    .A(_02973_));
 sg13g2_buf_2 fanout405 (.A(_02972_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_02911_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_12347_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_12164_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_12151_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_12059_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_11660_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_10123_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_09995_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_09728_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_09713_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_09686_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_09665_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_09336_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_09194_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_08966_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_08944_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_08920_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_08855_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_08735_),
    .X(net424));
 sg13g2_buf_4 fanout425 (.X(net425),
    .A(_08655_));
 sg13g2_buf_2 fanout426 (.A(_07450_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_06232_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_06231_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_06226_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_06148_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_06147_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_06142_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_06068_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_05892_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_05178_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_05045_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_05031_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_05027_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_05017_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_05008_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_04988_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_04976_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_04936_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_04928_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_04927_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_04922_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_04908_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_04825_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_04822_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_04810_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_03860_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_03859_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_03858_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_03630_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_03629_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_03606_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_03589_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_03585_),
    .X(net458));
 sg13g2_buf_1 fanout459 (.A(_03583_),
    .X(net459));
 sg13g2_buf_4 fanout460 (.X(net460),
    .A(_03012_));
 sg13g2_buf_4 fanout461 (.X(net461),
    .A(_03011_));
 sg13g2_buf_4 fanout462 (.X(net462),
    .A(_03008_));
 sg13g2_buf_2 fanout463 (.A(_03006_),
    .X(net463));
 sg13g2_buf_4 fanout464 (.X(net464),
    .A(_02995_));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(_02993_));
 sg13g2_buf_2 fanout466 (.A(_02856_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_02805_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_12521_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_12147_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_11519_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_10557_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_09994_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(_09335_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(_08988_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_08900_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_08879_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_08758_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_08736_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_08713_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_08685_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_08654_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_08649_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_08345_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_07867_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_07422_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_06320_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_06319_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_06318_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_06058_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_06004_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_06001_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_05992_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_05991_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_05952_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_05949_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_05941_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_05940_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_05878_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_05534_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_05160_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_05100_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_05044_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_05030_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_05026_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_05016_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_04987_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_04975_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_04859_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_04827_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_04815_),
    .X(net510));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(_04808_));
 sg13g2_buf_4 fanout512 (.X(net512),
    .A(_03628_));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(_03624_));
 sg13g2_buf_4 fanout514 (.X(net514),
    .A(_03616_));
 sg13g2_buf_4 fanout515 (.X(net515),
    .A(_03613_));
 sg13g2_buf_4 fanout516 (.X(net516),
    .A(_03599_));
 sg13g2_buf_2 fanout517 (.A(_03594_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_03592_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_03591_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_03586_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_03584_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_03582_),
    .X(net522));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(_03581_));
 sg13g2_buf_2 fanout524 (.A(_02992_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_02740_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_02689_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_12624_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_12465_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_12295_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_11585_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_10748_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_10659_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_10336_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_10253_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_10237_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_10180_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_10134_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_10107_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_10056_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_09757_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(_09533_),
    .X(net541));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(_09078_));
 sg13g2_buf_2 fanout543 (.A(_08947_),
    .X(net543));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(_08922_));
 sg13g2_buf_4 fanout545 (.X(net545),
    .A(_08683_));
 sg13g2_buf_2 fanout546 (.A(_08682_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_08653_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_08650_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_08392_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_08364_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_08357_),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_08348_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(_08344_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_08333_),
    .X(net554));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(_08329_));
 sg13g2_buf_2 fanout556 (.A(_08323_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_08085_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_07925_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_07837_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_07733_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_07647_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_07611_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_07601_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_07572_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_07518_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_07501_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_07459_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_07421_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_07365_),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(_07355_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_07348_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_07281_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_07064_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_06735_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_06227_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_06221_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_06143_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_06137_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_05977_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_05922_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_05195_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_05003_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_04898_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_04858_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_03888_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_03866_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_03861_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_03856_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_03855_),
    .X(net589));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(_03851_));
 sg13g2_buf_2 fanout591 (.A(_03627_),
    .X(net591));
 sg13g2_buf_4 fanout592 (.X(net592),
    .A(_03621_));
 sg13g2_buf_2 fanout593 (.A(_03617_),
    .X(net593));
 sg13g2_buf_4 fanout594 (.X(net594),
    .A(_03605_));
 sg13g2_buf_2 fanout595 (.A(_03593_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_03590_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_03580_),
    .X(net597));
 sg13g2_buf_4 fanout598 (.X(net598),
    .A(_02991_));
 sg13g2_buf_2 fanout599 (.A(_12668_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_12561_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_12212_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_12056_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_12024_),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_11993_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_11895_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_11553_),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_11494_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_10648_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_10561_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_10296_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_10286_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_10258_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_10252_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_10238_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_10106_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_10054_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_09993_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_09954_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_09641_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_09461_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_09433_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_09424_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_09419_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_09413_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_09409_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_09403_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_09397_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_09379_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_09353_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_09352_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_09297_),
    .X(net631));
 sg13g2_buf_4 fanout632 (.X(net632),
    .A(_09266_));
 sg13g2_buf_2 fanout633 (.A(_08651_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_08393_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_08382_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_08347_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_08332_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_08328_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_08327_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_08322_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_08321_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_07854_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_07814_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_07656_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_06729_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_06205_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_06121_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_04913_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_03887_),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_03865_),
    .X(net650));
 sg13g2_buf_4 fanout651 (.X(net651),
    .A(_02990_));
 sg13g2_buf_2 fanout652 (.A(_02971_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_12667_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_12009_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_11943_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_11937_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_11936_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_11913_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_11885_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_11493_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_11416_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_10686_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_10634_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_10631_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_10586_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_10353_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_10295_),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(_10288_),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(_10285_),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(_10266_),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_10262_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_10257_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_10053_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_09992_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_09879_),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(_09744_),
    .X(net676));
 sg13g2_buf_4 fanout677 (.X(net677),
    .A(_09739_));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(_09538_));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(_09501_));
 sg13g2_buf_8 fanout680 (.A(_09500_),
    .X(net680));
 sg13g2_buf_4 fanout681 (.X(net681),
    .A(_09497_));
 sg13g2_buf_8 fanout682 (.A(_09496_),
    .X(net682));
 sg13g2_buf_4 fanout683 (.X(net683),
    .A(_09494_));
 sg13g2_buf_8 fanout684 (.A(_09493_),
    .X(net684));
 sg13g2_buf_4 fanout685 (.X(net685),
    .A(_09460_));
 sg13g2_buf_2 fanout686 (.A(_09449_),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_09436_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_09430_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_09418_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(_09412_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_09408_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(_09402_),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_09386_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_09378_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(_09286_),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_09201_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_08780_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(_08399_),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(_08370_),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(_08355_),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_08342_),
    .X(net701));
 sg13g2_buf_4 fanout702 (.X(net702),
    .A(_08338_));
 sg13g2_buf_2 fanout703 (.A(_08320_),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(_08315_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_08314_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_06768_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(_06210_),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(_06208_),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(_06207_),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(_06126_),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(_06124_),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(_06123_),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(_06019_),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(_05970_),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(_05910_),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(_05900_),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(_05065_),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(_04812_),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(_03618_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(_03588_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_03385_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_03018_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_03016_),
    .X(net723));
 sg13g2_buf_1 fanout724 (.A(_02998_),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_02997_),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_02994_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(_02983_),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(_02980_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(_02978_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_02970_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_12111_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_11963_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_11931_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(_11927_),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_11926_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_10883_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_10817_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_10714_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_10695_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_10683_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_10669_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_10630_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_10620_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_10613_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_10603_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_10601_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_10597_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_10585_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_10428_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_10414_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_10360_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_10352_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_10345_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_10341_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_10291_),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_10287_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(_10284_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_10279_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_10277_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_10261_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_10256_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_10116_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_10052_),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_09878_),
    .X(net764));
 sg13g2_buf_4 fanout765 (.X(net765),
    .A(_09653_));
 sg13g2_buf_8 fanout766 (.A(_09539_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_09524_),
    .X(net767));
 sg13g2_buf_8 fanout768 (.A(_09499_),
    .X(net768));
 sg13g2_buf_8 fanout769 (.A(_09478_),
    .X(net769));
 sg13g2_buf_4 fanout770 (.X(net770),
    .A(_09476_));
 sg13g2_buf_4 fanout771 (.X(net771),
    .A(_09473_));
 sg13g2_buf_8 fanout772 (.A(_09472_),
    .X(net772));
 sg13g2_buf_8 fanout773 (.A(_09456_),
    .X(net773));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(_09450_));
 sg13g2_buf_4 fanout775 (.X(net775),
    .A(_09447_));
 sg13g2_buf_8 fanout776 (.A(_09446_),
    .X(net776));
 sg13g2_buf_4 fanout777 (.X(net777),
    .A(_09442_));
 sg13g2_buf_2 fanout778 (.A(_09440_),
    .X(net778));
 sg13g2_buf_4 fanout779 (.X(net779),
    .A(_09438_));
 sg13g2_buf_2 fanout780 (.A(_09342_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_09294_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_09287_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_09270_),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(_09200_),
    .X(net784));
 sg13g2_buf_8 fanout785 (.A(_08721_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_08657_),
    .X(net786));
 sg13g2_buf_8 fanout787 (.A(_08639_),
    .X(net787));
 sg13g2_buf_8 fanout788 (.A(_08628_),
    .X(net788));
 sg13g2_buf_8 fanout789 (.A(_08623_),
    .X(net789));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(_08618_));
 sg13g2_buf_4 fanout791 (.X(net791),
    .A(_08397_));
 sg13g2_buf_4 fanout792 (.X(net792),
    .A(_08341_));
 sg13g2_buf_2 fanout793 (.A(_08337_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(_08313_),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_08300_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(_08290_),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_08276_));
 sg13g2_buf_2 fanout798 (.A(_06779_),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(_06748_),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(_06467_),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(_06466_),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(_06465_),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(_06463_),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(_06448_),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(_06447_),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(_06445_),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(_06443_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_06434_),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(_06410_),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(_06404_),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(_06401_),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(_06398_),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(_06395_),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(_06376_),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(_06371_),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(_06364_),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(_06353_),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(_06213_),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(_06212_),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(_06211_),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_06129_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(_06128_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(_06127_),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(_06014_),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(_06002_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_05981_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_05963_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_05950_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_05927_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_05891_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_04809_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_03844_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_03573_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_03035_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(_03021_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_03020_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_03019_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_03001_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_03000_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_02999_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_02996_),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_02989_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_02987_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_02985_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(_02982_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_02979_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_02977_),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_02952_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_02709_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_12677_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_12516_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_12176_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_12037_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_11974_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_11955_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_11954_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_11949_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_11925_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_11909_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_11905_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_11525_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_10889_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_10688_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_10637_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_10635_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_10622_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_10614_),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(_10612_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_10602_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(_10600_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_10584_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_10565_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_10409_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(_10390_),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(_10348_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_10326_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_10283_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_10278_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_10276_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_10268_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_10255_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_10164_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_10158_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_10152_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_10146_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_10133_),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(_10115_),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(_10105_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(_10051_),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_10049_),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_09877_),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(_09856_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(_09811_),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_09555_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_09515_),
    .X(net895));
 sg13g2_buf_8 fanout896 (.A(_09452_),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_09358_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_09340_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(_09293_),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(_09273_),
    .X(net900));
 sg13g2_buf_4 fanout901 (.X(net901),
    .A(_09269_));
 sg13g2_buf_2 fanout902 (.A(_09199_),
    .X(net902));
 sg13g2_buf_8 fanout903 (.A(_08865_),
    .X(net903));
 sg13g2_buf_4 fanout904 (.X(net904),
    .A(_08844_));
 sg13g2_buf_8 fanout905 (.A(_08843_),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(_08788_),
    .X(net906));
 sg13g2_buf_4 fanout907 (.X(net907),
    .A(_08722_));
 sg13g2_buf_8 fanout908 (.A(_08703_),
    .X(net908));
 sg13g2_buf_8 fanout909 (.A(_08700_),
    .X(net909));
 sg13g2_buf_4 fanout910 (.X(net910),
    .A(_08697_));
 sg13g2_buf_8 fanout911 (.A(_08696_),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_08666_),
    .X(net912));
 sg13g2_buf_4 fanout913 (.X(net913),
    .A(_08643_));
 sg13g2_buf_4 fanout914 (.X(net914),
    .A(_08640_));
 sg13g2_buf_4 fanout915 (.X(net915),
    .A(_08634_));
 sg13g2_buf_4 fanout916 (.X(net916),
    .A(_08633_));
 sg13g2_buf_4 fanout917 (.X(net917),
    .A(_08630_));
 sg13g2_buf_4 fanout918 (.X(net918),
    .A(_08625_));
 sg13g2_buf_4 fanout919 (.X(net919),
    .A(_08622_));
 sg13g2_buf_2 fanout920 (.A(_08621_),
    .X(net920));
 sg13g2_buf_4 fanout921 (.X(net921),
    .A(_08617_));
 sg13g2_buf_4 fanout922 (.X(net922),
    .A(_08599_));
 sg13g2_buf_2 fanout923 (.A(_08390_),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(_08366_),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(_08340_),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(_08335_),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(_08317_),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(_08312_),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(_08283_),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(_08279_),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(_08275_),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(_07092_),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(_07052_),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(_07045_),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(_07039_),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_07037_),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(_07023_),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(_06778_),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_06666_),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(_06436_),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(_06435_),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(_06431_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_06412_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(_06411_),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_06407_),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(_06015_),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(_06010_),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_06003_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_05964_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(_05959_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(_05951_),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(_05902_),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_05901_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_05881_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(_05880_),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_05867_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_05858_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_05842_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_05406_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_04911_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_04801_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_04704_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_04675_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_04644_),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(_03572_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(_03034_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_02988_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_02986_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_02984_),
    .X(net969));
 sg13g2_buf_4 fanout970 (.X(net970),
    .A(_02835_));
 sg13g2_buf_4 fanout971 (.X(net971),
    .A(_02831_));
 sg13g2_buf_4 fanout972 (.X(net972),
    .A(_02823_));
 sg13g2_buf_2 fanout973 (.A(_12725_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_12716_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(_12688_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_12682_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_12672_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_12456_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_12452_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_12448_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_12341_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_12333_),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(_12281_),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(_12267_),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(_12263_),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(_12255_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_12193_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(_12144_),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(_12140_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_12136_),
    .X(net990));
 sg13g2_buf_4 fanout991 (.X(net991),
    .A(_12133_));
 sg13g2_buf_2 fanout992 (.A(_12130_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_12119_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_12103_),
    .X(net994));
 sg13g2_buf_4 fanout995 (.X(net995),
    .A(_12063_));
 sg13g2_buf_4 fanout996 (.X(net996),
    .A(_12046_));
 sg13g2_buf_2 fanout997 (.A(_12039_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_12028_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_12027_),
    .X(net999));
 sg13g2_buf_4 fanout1000 (.X(net1000),
    .A(_12023_));
 sg13g2_buf_2 fanout1001 (.A(_11953_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_11948_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_11264_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_10662_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_10621_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_10607_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(_10595_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_10588_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(_10587_),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(_10583_),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(_10424_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(_10325_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_10319_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_10273_),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_10263_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(_10259_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_10254_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_10232_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_10230_),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_10132_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(_10104_),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(_10098_),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(_10092_),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_10086_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_10080_),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(_10075_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(_10070_),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_10057_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_10048_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_09999_),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_09901_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(_09890_),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(_09887_),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_09568_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_09526_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_09365_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(_09357_),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(_09332_),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(_09272_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_09268_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_09209_),
    .X(net1041));
 sg13g2_buf_4 fanout1042 (.X(net1042),
    .A(_09205_));
 sg13g2_buf_4 fanout1043 (.X(net1043),
    .A(_09203_));
 sg13g2_buf_2 fanout1044 (.A(_09198_),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(_09181_),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(_09167_),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_09101_),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(_09002_),
    .X(net1048));
 sg13g2_buf_4 fanout1049 (.X(net1049),
    .A(_08866_));
 sg13g2_buf_2 fanout1050 (.A(_08820_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(_08769_),
    .X(net1051));
 sg13g2_buf_4 fanout1052 (.X(net1052),
    .A(_08707_));
 sg13g2_buf_2 fanout1053 (.A(_08695_),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(_08629_),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_08624_),
    .X(net1055));
 sg13g2_buf_4 fanout1056 (.X(net1056),
    .A(_08620_));
 sg13g2_buf_2 fanout1057 (.A(_08619_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(_08610_),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_08588_),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_08579_),
    .X(net1060));
 sg13g2_buf_4 fanout1061 (.X(net1061),
    .A(_08560_));
 sg13g2_buf_4 fanout1062 (.X(net1062),
    .A(_08540_));
 sg13g2_buf_2 fanout1063 (.A(_08495_),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(_08492_),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(_08491_),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(_08485_),
    .X(net1066));
 sg13g2_buf_4 fanout1067 (.X(net1067),
    .A(_08481_));
 sg13g2_buf_4 fanout1068 (.X(net1068),
    .A(_08316_));
 sg13g2_buf_2 fanout1069 (.A(_08267_),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(_08263_),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(_08261_),
    .X(net1071));
 sg13g2_buf_2 fanout1072 (.A(_08258_),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(_08256_),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(_08046_),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(_08044_),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(_08042_),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_07756_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(_07114_),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(_07024_),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(_07022_),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(_05835_),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(_12584_),
    .X(net1082));
 sg13g2_buf_2 fanout1083 (.A(_12271_),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(_12246_),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(_12243_),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(_12237_),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_12132_),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(_12096_),
    .X(net1088));
 sg13g2_buf_2 fanout1089 (.A(_12090_),
    .X(net1089));
 sg13g2_buf_2 fanout1090 (.A(_12084_),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(_12073_),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(_12062_),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(_12045_),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(_12025_),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(_12022_),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(_12005_),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(_11998_),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(_11979_),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(_11977_),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(_11970_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(_11232_),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(_11159_),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(_10815_),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(_10703_),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(_10508_),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(_10418_),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(_10386_),
    .X(net1107));
 sg13g2_buf_2 fanout1108 (.A(_10371_),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(_10318_),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(_10227_),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(_10225_),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(_10222_),
    .X(net1112));
 sg13g2_buf_2 fanout1113 (.A(_10079_),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(_09910_),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(_09886_),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(_09880_),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(_09874_),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(_09846_),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(_09398_),
    .X(net1119));
 sg13g2_buf_2 fanout1120 (.A(_09383_),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(_09347_),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(_09339_),
    .X(net1122));
 sg13g2_buf_2 fanout1123 (.A(_09210_),
    .X(net1123));
 sg13g2_buf_2 fanout1124 (.A(_09100_),
    .X(net1124));
 sg13g2_buf_2 fanout1125 (.A(_08583_),
    .X(net1125));
 sg13g2_buf_2 fanout1126 (.A(_08582_),
    .X(net1126));
 sg13g2_buf_2 fanout1127 (.A(_08549_),
    .X(net1127));
 sg13g2_buf_2 fanout1128 (.A(_08473_),
    .X(net1128));
 sg13g2_buf_2 fanout1129 (.A(_08463_),
    .X(net1129));
 sg13g2_buf_2 fanout1130 (.A(_08260_),
    .X(net1130));
 sg13g2_tiehi _27539__1131 (.L_HI(net1131));
 sg13g2_tiehi _27540__1132 (.L_HI(net1132));
 sg13g2_tiehi _27541__1133 (.L_HI(net1133));
 sg13g2_tiehi _27542__1134 (.L_HI(net1134));
 sg13g2_tiehi _27543__1135 (.L_HI(net1135));
 sg13g2_tiehi \cpu.dcache.r_data[0][0]$_DFFE_PP__1136  (.L_HI(net1136));
 sg13g2_tiehi \cpu.dcache.r_data[0][10]$_DFFE_PP__1137  (.L_HI(net1137));
 sg13g2_tiehi \cpu.dcache.r_data[0][11]$_DFFE_PP__1138  (.L_HI(net1138));
 sg13g2_tiehi \cpu.dcache.r_data[0][12]$_DFFE_PP__1139  (.L_HI(net1139));
 sg13g2_tiehi \cpu.dcache.r_data[0][13]$_DFFE_PP__1140  (.L_HI(net1140));
 sg13g2_tiehi \cpu.dcache.r_data[0][14]$_DFFE_PP__1141  (.L_HI(net1141));
 sg13g2_tiehi \cpu.dcache.r_data[0][15]$_DFFE_PP__1142  (.L_HI(net1142));
 sg13g2_tiehi \cpu.dcache.r_data[0][16]$_DFFE_PP__1143  (.L_HI(net1143));
 sg13g2_tiehi \cpu.dcache.r_data[0][17]$_DFFE_PP__1144  (.L_HI(net1144));
 sg13g2_tiehi \cpu.dcache.r_data[0][18]$_DFFE_PP__1145  (.L_HI(net1145));
 sg13g2_tiehi \cpu.dcache.r_data[0][19]$_DFFE_PP__1146  (.L_HI(net1146));
 sg13g2_tiehi \cpu.dcache.r_data[0][1]$_DFFE_PP__1147  (.L_HI(net1147));
 sg13g2_tiehi \cpu.dcache.r_data[0][20]$_DFFE_PP__1148  (.L_HI(net1148));
 sg13g2_tiehi \cpu.dcache.r_data[0][21]$_DFFE_PP__1149  (.L_HI(net1149));
 sg13g2_tiehi \cpu.dcache.r_data[0][22]$_DFFE_PP__1150  (.L_HI(net1150));
 sg13g2_tiehi \cpu.dcache.r_data[0][23]$_DFFE_PP__1151  (.L_HI(net1151));
 sg13g2_tiehi \cpu.dcache.r_data[0][24]$_DFFE_PP__1152  (.L_HI(net1152));
 sg13g2_tiehi \cpu.dcache.r_data[0][25]$_DFFE_PP__1153  (.L_HI(net1153));
 sg13g2_tiehi \cpu.dcache.r_data[0][26]$_DFFE_PP__1154  (.L_HI(net1154));
 sg13g2_tiehi \cpu.dcache.r_data[0][27]$_DFFE_PP__1155  (.L_HI(net1155));
 sg13g2_tiehi \cpu.dcache.r_data[0][28]$_DFFE_PP__1156  (.L_HI(net1156));
 sg13g2_tiehi \cpu.dcache.r_data[0][29]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \cpu.dcache.r_data[0][2]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \cpu.dcache.r_data[0][30]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \cpu.dcache.r_data[0][31]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \cpu.dcache.r_data[0][3]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \cpu.dcache.r_data[0][4]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \cpu.dcache.r_data[0][5]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \cpu.dcache.r_data[0][6]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \cpu.dcache.r_data[0][7]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \cpu.dcache.r_data[0][8]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \cpu.dcache.r_data[0][9]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \cpu.dcache.r_data[1][0]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \cpu.dcache.r_data[1][10]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \cpu.dcache.r_data[1][11]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \cpu.dcache.r_data[1][12]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \cpu.dcache.r_data[1][13]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \cpu.dcache.r_data[1][14]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \cpu.dcache.r_data[1][15]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \cpu.dcache.r_data[1][16]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \cpu.dcache.r_data[1][17]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \cpu.dcache.r_data[1][18]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \cpu.dcache.r_data[1][19]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \cpu.dcache.r_data[1][1]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \cpu.dcache.r_data[1][20]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \cpu.dcache.r_data[1][21]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \cpu.dcache.r_data[1][22]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \cpu.dcache.r_data[1][23]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \cpu.dcache.r_data[1][24]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \cpu.dcache.r_data[1][25]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \cpu.dcache.r_data[1][26]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \cpu.dcache.r_data[1][27]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \cpu.dcache.r_data[1][28]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \cpu.dcache.r_data[1][29]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \cpu.dcache.r_data[1][2]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \cpu.dcache.r_data[1][30]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \cpu.dcache.r_data[1][31]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \cpu.dcache.r_data[1][3]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \cpu.dcache.r_data[1][4]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \cpu.dcache.r_data[1][5]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \cpu.dcache.r_data[1][6]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \cpu.dcache.r_data[1][7]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \cpu.dcache.r_data[1][8]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \cpu.dcache.r_data[1][9]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \cpu.dcache.r_data[2][0]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \cpu.dcache.r_data[2][10]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \cpu.dcache.r_data[2][11]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \cpu.dcache.r_data[2][12]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \cpu.dcache.r_data[2][13]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \cpu.dcache.r_data[2][14]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \cpu.dcache.r_data[2][15]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \cpu.dcache.r_data[2][16]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \cpu.dcache.r_data[2][17]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \cpu.dcache.r_data[2][18]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \cpu.dcache.r_data[2][19]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \cpu.dcache.r_data[2][1]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \cpu.dcache.r_data[2][20]$_DFFE_PP__1212  (.L_HI(net1212));
 sg13g2_tiehi \cpu.dcache.r_data[2][21]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \cpu.dcache.r_data[2][22]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \cpu.dcache.r_data[2][23]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \cpu.dcache.r_data[2][24]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \cpu.dcache.r_data[2][25]$_DFFE_PP__1217  (.L_HI(net1217));
 sg13g2_tiehi \cpu.dcache.r_data[2][26]$_DFFE_PP__1218  (.L_HI(net1218));
 sg13g2_tiehi \cpu.dcache.r_data[2][27]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \cpu.dcache.r_data[2][28]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \cpu.dcache.r_data[2][29]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \cpu.dcache.r_data[2][2]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \cpu.dcache.r_data[2][30]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \cpu.dcache.r_data[2][31]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \cpu.dcache.r_data[2][3]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \cpu.dcache.r_data[2][4]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \cpu.dcache.r_data[2][5]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \cpu.dcache.r_data[2][6]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \cpu.dcache.r_data[2][7]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \cpu.dcache.r_data[2][8]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \cpu.dcache.r_data[2][9]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \cpu.dcache.r_data[3][0]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \cpu.dcache.r_data[3][10]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \cpu.dcache.r_data[3][11]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \cpu.dcache.r_data[3][12]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \cpu.dcache.r_data[3][13]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \cpu.dcache.r_data[3][14]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \cpu.dcache.r_data[3][15]$_DFFE_PP__1238  (.L_HI(net1238));
 sg13g2_tiehi \cpu.dcache.r_data[3][16]$_DFFE_PP__1239  (.L_HI(net1239));
 sg13g2_tiehi \cpu.dcache.r_data[3][17]$_DFFE_PP__1240  (.L_HI(net1240));
 sg13g2_tiehi \cpu.dcache.r_data[3][18]$_DFFE_PP__1241  (.L_HI(net1241));
 sg13g2_tiehi \cpu.dcache.r_data[3][19]$_DFFE_PP__1242  (.L_HI(net1242));
 sg13g2_tiehi \cpu.dcache.r_data[3][1]$_DFFE_PP__1243  (.L_HI(net1243));
 sg13g2_tiehi \cpu.dcache.r_data[3][20]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \cpu.dcache.r_data[3][21]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \cpu.dcache.r_data[3][22]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \cpu.dcache.r_data[3][23]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \cpu.dcache.r_data[3][24]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \cpu.dcache.r_data[3][25]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \cpu.dcache.r_data[3][26]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \cpu.dcache.r_data[3][27]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \cpu.dcache.r_data[3][28]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \cpu.dcache.r_data[3][29]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \cpu.dcache.r_data[3][2]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \cpu.dcache.r_data[3][30]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \cpu.dcache.r_data[3][31]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \cpu.dcache.r_data[3][3]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \cpu.dcache.r_data[3][4]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \cpu.dcache.r_data[3][5]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \cpu.dcache.r_data[3][6]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \cpu.dcache.r_data[3][7]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \cpu.dcache.r_data[3][8]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \cpu.dcache.r_data[3][9]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \cpu.dcache.r_data[4][0]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \cpu.dcache.r_data[4][10]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \cpu.dcache.r_data[4][11]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \cpu.dcache.r_data[4][12]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \cpu.dcache.r_data[4][13]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \cpu.dcache.r_data[4][14]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \cpu.dcache.r_data[4][15]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \cpu.dcache.r_data[4][16]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \cpu.dcache.r_data[4][17]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \cpu.dcache.r_data[4][18]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \cpu.dcache.r_data[4][19]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \cpu.dcache.r_data[4][1]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \cpu.dcache.r_data[4][20]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \cpu.dcache.r_data[4][21]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \cpu.dcache.r_data[4][22]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \cpu.dcache.r_data[4][23]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \cpu.dcache.r_data[4][24]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \cpu.dcache.r_data[4][25]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \cpu.dcache.r_data[4][26]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \cpu.dcache.r_data[4][27]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \cpu.dcache.r_data[4][28]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \cpu.dcache.r_data[4][29]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \cpu.dcache.r_data[4][2]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \cpu.dcache.r_data[4][30]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \cpu.dcache.r_data[4][31]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \cpu.dcache.r_data[4][3]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \cpu.dcache.r_data[4][4]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \cpu.dcache.r_data[4][5]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \cpu.dcache.r_data[4][6]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \cpu.dcache.r_data[4][7]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \cpu.dcache.r_data[4][8]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \cpu.dcache.r_data[4][9]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \cpu.dcache.r_data[5][0]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \cpu.dcache.r_data[5][10]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \cpu.dcache.r_data[5][11]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \cpu.dcache.r_data[5][12]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \cpu.dcache.r_data[5][13]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \cpu.dcache.r_data[5][14]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \cpu.dcache.r_data[5][15]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \cpu.dcache.r_data[5][16]$_DFFE_PP__1303  (.L_HI(net1303));
 sg13g2_tiehi \cpu.dcache.r_data[5][17]$_DFFE_PP__1304  (.L_HI(net1304));
 sg13g2_tiehi \cpu.dcache.r_data[5][18]$_DFFE_PP__1305  (.L_HI(net1305));
 sg13g2_tiehi \cpu.dcache.r_data[5][19]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \cpu.dcache.r_data[5][1]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \cpu.dcache.r_data[5][20]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \cpu.dcache.r_data[5][21]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \cpu.dcache.r_data[5][22]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \cpu.dcache.r_data[5][23]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \cpu.dcache.r_data[5][24]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \cpu.dcache.r_data[5][25]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \cpu.dcache.r_data[5][26]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \cpu.dcache.r_data[5][27]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \cpu.dcache.r_data[5][28]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \cpu.dcache.r_data[5][29]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \cpu.dcache.r_data[5][2]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \cpu.dcache.r_data[5][30]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \cpu.dcache.r_data[5][31]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \cpu.dcache.r_data[5][3]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \cpu.dcache.r_data[5][4]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \cpu.dcache.r_data[5][5]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \cpu.dcache.r_data[5][6]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \cpu.dcache.r_data[5][7]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \cpu.dcache.r_data[5][8]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \cpu.dcache.r_data[5][9]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \cpu.dcache.r_data[6][0]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \cpu.dcache.r_data[6][10]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \cpu.dcache.r_data[6][11]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \cpu.dcache.r_data[6][12]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \cpu.dcache.r_data[6][13]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \cpu.dcache.r_data[6][14]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \cpu.dcache.r_data[6][15]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \cpu.dcache.r_data[6][16]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \cpu.dcache.r_data[6][17]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \cpu.dcache.r_data[6][18]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \cpu.dcache.r_data[6][19]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \cpu.dcache.r_data[6][1]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \cpu.dcache.r_data[6][20]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \cpu.dcache.r_data[6][21]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \cpu.dcache.r_data[6][22]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \cpu.dcache.r_data[6][23]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \cpu.dcache.r_data[6][24]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \cpu.dcache.r_data[6][25]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \cpu.dcache.r_data[6][26]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \cpu.dcache.r_data[6][27]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \cpu.dcache.r_data[6][28]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \cpu.dcache.r_data[6][29]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \cpu.dcache.r_data[6][2]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \cpu.dcache.r_data[6][30]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \cpu.dcache.r_data[6][31]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \cpu.dcache.r_data[6][3]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \cpu.dcache.r_data[6][4]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \cpu.dcache.r_data[6][5]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \cpu.dcache.r_data[6][6]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \cpu.dcache.r_data[6][7]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \cpu.dcache.r_data[6][8]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \cpu.dcache.r_data[6][9]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \cpu.dcache.r_data[7][0]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \cpu.dcache.r_data[7][10]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \cpu.dcache.r_data[7][11]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \cpu.dcache.r_data[7][12]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \cpu.dcache.r_data[7][13]$_DFFE_PP__1364  (.L_HI(net1364));
 sg13g2_tiehi \cpu.dcache.r_data[7][14]$_DFFE_PP__1365  (.L_HI(net1365));
 sg13g2_tiehi \cpu.dcache.r_data[7][15]$_DFFE_PP__1366  (.L_HI(net1366));
 sg13g2_tiehi \cpu.dcache.r_data[7][16]$_DFFE_PP__1367  (.L_HI(net1367));
 sg13g2_tiehi \cpu.dcache.r_data[7][17]$_DFFE_PP__1368  (.L_HI(net1368));
 sg13g2_tiehi \cpu.dcache.r_data[7][18]$_DFFE_PP__1369  (.L_HI(net1369));
 sg13g2_tiehi \cpu.dcache.r_data[7][19]$_DFFE_PP__1370  (.L_HI(net1370));
 sg13g2_tiehi \cpu.dcache.r_data[7][1]$_DFFE_PP__1371  (.L_HI(net1371));
 sg13g2_tiehi \cpu.dcache.r_data[7][20]$_DFFE_PP__1372  (.L_HI(net1372));
 sg13g2_tiehi \cpu.dcache.r_data[7][21]$_DFFE_PP__1373  (.L_HI(net1373));
 sg13g2_tiehi \cpu.dcache.r_data[7][22]$_DFFE_PP__1374  (.L_HI(net1374));
 sg13g2_tiehi \cpu.dcache.r_data[7][23]$_DFFE_PP__1375  (.L_HI(net1375));
 sg13g2_tiehi \cpu.dcache.r_data[7][24]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \cpu.dcache.r_data[7][25]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \cpu.dcache.r_data[7][26]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \cpu.dcache.r_data[7][27]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \cpu.dcache.r_data[7][28]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \cpu.dcache.r_data[7][29]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \cpu.dcache.r_data[7][2]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \cpu.dcache.r_data[7][30]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \cpu.dcache.r_data[7][31]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \cpu.dcache.r_data[7][3]$_DFFE_PP__1385  (.L_HI(net1385));
 sg13g2_tiehi \cpu.dcache.r_data[7][4]$_DFFE_PP__1386  (.L_HI(net1386));
 sg13g2_tiehi \cpu.dcache.r_data[7][5]$_DFFE_PP__1387  (.L_HI(net1387));
 sg13g2_tiehi \cpu.dcache.r_data[7][6]$_DFFE_PP__1388  (.L_HI(net1388));
 sg13g2_tiehi \cpu.dcache.r_data[7][7]$_DFFE_PP__1389  (.L_HI(net1389));
 sg13g2_tiehi \cpu.dcache.r_data[7][8]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \cpu.dcache.r_data[7][9]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P__1392  (.L_HI(net1392));
 sg13g2_tiehi \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P__1393  (.L_HI(net1393));
 sg13g2_tiehi \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P__1394  (.L_HI(net1394));
 sg13g2_tiehi \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P__1395  (.L_HI(net1395));
 sg13g2_tiehi \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P__1396  (.L_HI(net1396));
 sg13g2_tiehi \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P__1397  (.L_HI(net1397));
 sg13g2_tiehi \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P__1398  (.L_HI(net1398));
 sg13g2_tiehi \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P__1399  (.L_HI(net1399));
 sg13g2_tiehi \cpu.dcache.r_offset[0]$_SDFF_PN0__1400  (.L_HI(net1400));
 sg13g2_tiehi \cpu.dcache.r_offset[1]$_SDFF_PN0__1401  (.L_HI(net1401));
 sg13g2_tiehi \cpu.dcache.r_offset[2]$_SDFF_PN0__1402  (.L_HI(net1402));
 sg13g2_tiehi \cpu.dcache.r_tag[0][0]$_DFFE_PP__1403  (.L_HI(net1403));
 sg13g2_tiehi \cpu.dcache.r_tag[0][10]$_DFFE_PP__1404  (.L_HI(net1404));
 sg13g2_tiehi \cpu.dcache.r_tag[0][11]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \cpu.dcache.r_tag[0][12]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \cpu.dcache.r_tag[0][13]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \cpu.dcache.r_tag[0][14]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \cpu.dcache.r_tag[0][15]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \cpu.dcache.r_tag[0][16]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \cpu.dcache.r_tag[0][17]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \cpu.dcache.r_tag[0][18]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \cpu.dcache.r_tag[0][1]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \cpu.dcache.r_tag[0][2]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \cpu.dcache.r_tag[0][3]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \cpu.dcache.r_tag[0][4]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \cpu.dcache.r_tag[0][5]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \cpu.dcache.r_tag[0][6]$_DFFE_PP__1418  (.L_HI(net1418));
 sg13g2_tiehi \cpu.dcache.r_tag[0][7]$_DFFE_PP__1419  (.L_HI(net1419));
 sg13g2_tiehi \cpu.dcache.r_tag[0][8]$_DFFE_PP__1420  (.L_HI(net1420));
 sg13g2_tiehi \cpu.dcache.r_tag[0][9]$_DFFE_PP__1421  (.L_HI(net1421));
 sg13g2_tiehi \cpu.dcache.r_tag[1][0]$_DFFE_PP__1422  (.L_HI(net1422));
 sg13g2_tiehi \cpu.dcache.r_tag[1][10]$_DFFE_PP__1423  (.L_HI(net1423));
 sg13g2_tiehi \cpu.dcache.r_tag[1][11]$_DFFE_PP__1424  (.L_HI(net1424));
 sg13g2_tiehi \cpu.dcache.r_tag[1][12]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \cpu.dcache.r_tag[1][13]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \cpu.dcache.r_tag[1][14]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \cpu.dcache.r_tag[1][15]$_DFFE_PP__1428  (.L_HI(net1428));
 sg13g2_tiehi \cpu.dcache.r_tag[1][16]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \cpu.dcache.r_tag[1][17]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \cpu.dcache.r_tag[1][18]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \cpu.dcache.r_tag[1][1]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \cpu.dcache.r_tag[1][2]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \cpu.dcache.r_tag[1][3]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \cpu.dcache.r_tag[1][4]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \cpu.dcache.r_tag[1][5]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \cpu.dcache.r_tag[1][6]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \cpu.dcache.r_tag[1][7]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \cpu.dcache.r_tag[1][8]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \cpu.dcache.r_tag[1][9]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \cpu.dcache.r_tag[2][0]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \cpu.dcache.r_tag[2][10]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \cpu.dcache.r_tag[2][11]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \cpu.dcache.r_tag[2][12]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \cpu.dcache.r_tag[2][13]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \cpu.dcache.r_tag[2][14]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \cpu.dcache.r_tag[2][15]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \cpu.dcache.r_tag[2][16]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \cpu.dcache.r_tag[2][17]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \cpu.dcache.r_tag[2][18]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \cpu.dcache.r_tag[2][1]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \cpu.dcache.r_tag[2][2]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \cpu.dcache.r_tag[2][3]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \cpu.dcache.r_tag[2][4]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \cpu.dcache.r_tag[2][5]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \cpu.dcache.r_tag[2][6]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \cpu.dcache.r_tag[2][7]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \cpu.dcache.r_tag[2][8]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \cpu.dcache.r_tag[2][9]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \cpu.dcache.r_tag[3][0]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \cpu.dcache.r_tag[3][10]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \cpu.dcache.r_tag[3][11]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \cpu.dcache.r_tag[3][12]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \cpu.dcache.r_tag[3][13]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \cpu.dcache.r_tag[3][14]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \cpu.dcache.r_tag[3][15]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \cpu.dcache.r_tag[3][16]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \cpu.dcache.r_tag[3][17]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \cpu.dcache.r_tag[3][18]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \cpu.dcache.r_tag[3][1]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \cpu.dcache.r_tag[3][2]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \cpu.dcache.r_tag[3][3]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \cpu.dcache.r_tag[3][4]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \cpu.dcache.r_tag[3][5]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \cpu.dcache.r_tag[3][6]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \cpu.dcache.r_tag[3][7]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \cpu.dcache.r_tag[3][8]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \cpu.dcache.r_tag[3][9]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \cpu.dcache.r_tag[4][0]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \cpu.dcache.r_tag[4][10]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \cpu.dcache.r_tag[4][11]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \cpu.dcache.r_tag[4][12]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \cpu.dcache.r_tag[4][13]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \cpu.dcache.r_tag[4][14]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \cpu.dcache.r_tag[4][15]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \cpu.dcache.r_tag[4][16]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \cpu.dcache.r_tag[4][17]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \cpu.dcache.r_tag[4][18]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \cpu.dcache.r_tag[4][1]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \cpu.dcache.r_tag[4][2]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \cpu.dcache.r_tag[4][3]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \cpu.dcache.r_tag[4][4]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \cpu.dcache.r_tag[4][5]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \cpu.dcache.r_tag[4][6]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \cpu.dcache.r_tag[4][7]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \cpu.dcache.r_tag[4][8]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \cpu.dcache.r_tag[4][9]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \cpu.dcache.r_tag[5][0]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \cpu.dcache.r_tag[5][10]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \cpu.dcache.r_tag[5][11]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \cpu.dcache.r_tag[5][12]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \cpu.dcache.r_tag[5][13]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \cpu.dcache.r_tag[5][14]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \cpu.dcache.r_tag[5][15]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \cpu.dcache.r_tag[5][16]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \cpu.dcache.r_tag[5][17]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \cpu.dcache.r_tag[5][18]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \cpu.dcache.r_tag[5][1]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \cpu.dcache.r_tag[5][2]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \cpu.dcache.r_tag[5][3]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \cpu.dcache.r_tag[5][4]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \cpu.dcache.r_tag[5][5]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \cpu.dcache.r_tag[5][6]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \cpu.dcache.r_tag[5][7]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \cpu.dcache.r_tag[5][8]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \cpu.dcache.r_tag[5][9]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \cpu.dcache.r_tag[6][0]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \cpu.dcache.r_tag[6][10]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \cpu.dcache.r_tag[6][11]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \cpu.dcache.r_tag[6][12]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \cpu.dcache.r_tag[6][13]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \cpu.dcache.r_tag[6][14]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \cpu.dcache.r_tag[6][15]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \cpu.dcache.r_tag[6][16]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \cpu.dcache.r_tag[6][17]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \cpu.dcache.r_tag[6][18]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \cpu.dcache.r_tag[6][1]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \cpu.dcache.r_tag[6][2]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \cpu.dcache.r_tag[6][3]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \cpu.dcache.r_tag[6][4]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \cpu.dcache.r_tag[6][5]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \cpu.dcache.r_tag[6][6]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \cpu.dcache.r_tag[6][7]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \cpu.dcache.r_tag[6][8]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \cpu.dcache.r_tag[6][9]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \cpu.dcache.r_tag[7][0]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \cpu.dcache.r_tag[7][10]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \cpu.dcache.r_tag[7][11]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \cpu.dcache.r_tag[7][12]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \cpu.dcache.r_tag[7][13]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \cpu.dcache.r_tag[7][14]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \cpu.dcache.r_tag[7][15]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \cpu.dcache.r_tag[7][16]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \cpu.dcache.r_tag[7][17]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \cpu.dcache.r_tag[7][18]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \cpu.dcache.r_tag[7][1]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \cpu.dcache.r_tag[7][2]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \cpu.dcache.r_tag[7][3]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \cpu.dcache.r_tag[7][4]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \cpu.dcache.r_tag[7][5]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \cpu.dcache.r_tag[7][6]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \cpu.dcache.r_tag[7][7]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \cpu.dcache.r_tag[7][8]$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \cpu.dcache.r_tag[7][9]$_DFFE_PP__1554  (.L_HI(net1554));
 sg13g2_tiehi \cpu.dcache.r_valid[0]$_SDFFE_PP0P__1555  (.L_HI(net1555));
 sg13g2_tiehi \cpu.dcache.r_valid[1]$_SDFFE_PP0P__1556  (.L_HI(net1556));
 sg13g2_tiehi \cpu.dcache.r_valid[2]$_SDFFE_PP0P__1557  (.L_HI(net1557));
 sg13g2_tiehi \cpu.dcache.r_valid[3]$_SDFFE_PP0P__1558  (.L_HI(net1558));
 sg13g2_tiehi \cpu.dcache.r_valid[4]$_SDFFE_PP0P__1559  (.L_HI(net1559));
 sg13g2_tiehi \cpu.dcache.r_valid[5]$_SDFFE_PP0P__1560  (.L_HI(net1560));
 sg13g2_tiehi \cpu.dcache.r_valid[6]$_SDFFE_PP0P__1561  (.L_HI(net1561));
 sg13g2_tiehi \cpu.dcache.r_valid[7]$_SDFFE_PP0P__1562  (.L_HI(net1562));
 sg13g2_tiehi \cpu.dec.r_br$_DFFE_PP__1563  (.L_HI(net1563));
 sg13g2_tiehi \cpu.dec.r_cond[0]$_DFFE_PP__1564  (.L_HI(net1564));
 sg13g2_tiehi \cpu.dec.r_cond[1]$_DFFE_PP__1565  (.L_HI(net1565));
 sg13g2_tiehi \cpu.dec.r_cond[2]$_DFFE_PP__1566  (.L_HI(net1566));
 sg13g2_tiehi \cpu.dec.r_div$_DFFE_PP__1567  (.L_HI(net1567));
 sg13g2_tiehi \cpu.dec.r_flush_all$_DFFE_PP__1568  (.L_HI(net1568));
 sg13g2_tiehi \cpu.dec.r_flush_write$_DFFE_PP__1569  (.L_HI(net1569));
 sg13g2_tiehi \cpu.dec.r_imm[0]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \cpu.dec.r_imm[10]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \cpu.dec.r_imm[11]$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \cpu.dec.r_imm[12]$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \cpu.dec.r_imm[13]$_DFFE_PP__1574  (.L_HI(net1574));
 sg13g2_tiehi \cpu.dec.r_imm[14]$_DFFE_PP__1575  (.L_HI(net1575));
 sg13g2_tiehi \cpu.dec.r_imm[15]$_DFFE_PP__1576  (.L_HI(net1576));
 sg13g2_tiehi \cpu.dec.r_imm[1]$_DFFE_PP__1577  (.L_HI(net1577));
 sg13g2_tiehi \cpu.dec.r_imm[2]$_DFFE_PP__1578  (.L_HI(net1578));
 sg13g2_tiehi \cpu.dec.r_imm[3]$_DFFE_PP__1579  (.L_HI(net1579));
 sg13g2_tiehi \cpu.dec.r_imm[4]$_DFFE_PP__1580  (.L_HI(net1580));
 sg13g2_tiehi \cpu.dec.r_imm[5]$_DFFE_PP__1581  (.L_HI(net1581));
 sg13g2_tiehi \cpu.dec.r_imm[6]$_DFFE_PP__1582  (.L_HI(net1582));
 sg13g2_tiehi \cpu.dec.r_imm[7]$_DFFE_PP__1583  (.L_HI(net1583));
 sg13g2_tiehi \cpu.dec.r_imm[8]$_DFFE_PP__1584  (.L_HI(net1584));
 sg13g2_tiehi \cpu.dec.r_imm[9]$_DFFE_PP__1585  (.L_HI(net1585));
 sg13g2_tiehi \cpu.dec.r_inv_mmu$_DFFE_PP__1586  (.L_HI(net1586));
 sg13g2_tiehi \cpu.dec.r_io$_DFFE_PP__1587  (.L_HI(net1587));
 sg13g2_tiehi \cpu.dec.r_jmp$_SDFFCE_PP0P__1588  (.L_HI(net1588));
 sg13g2_tiehi \cpu.dec.r_load$_DFFE_PP__1589  (.L_HI(net1589));
 sg13g2_tiehi \cpu.dec.r_mult$_DFFE_PP__1590  (.L_HI(net1590));
 sg13g2_tiehi \cpu.dec.r_needs_rs2$_DFFE_PP__1591  (.L_HI(net1591));
 sg13g2_tiehi \cpu.dec.r_op[10]$_DFF_P__1592  (.L_HI(net1592));
 sg13g2_tiehi \cpu.dec.r_op[1]$_DFF_P__1593  (.L_HI(net1593));
 sg13g2_tiehi \cpu.dec.r_op[2]$_DFF_P__1594  (.L_HI(net1594));
 sg13g2_tiehi \cpu.dec.r_op[3]$_DFF_P__1595  (.L_HI(net1595));
 sg13g2_tiehi \cpu.dec.r_op[4]$_DFF_P__1596  (.L_HI(net1596));
 sg13g2_tiehi \cpu.dec.r_op[5]$_DFF_P__1597  (.L_HI(net1597));
 sg13g2_tiehi \cpu.dec.r_op[6]$_DFF_P__1598  (.L_HI(net1598));
 sg13g2_tiehi \cpu.dec.r_op[7]$_DFF_P__1599  (.L_HI(net1599));
 sg13g2_tiehi \cpu.dec.r_op[8]$_DFF_P__1600  (.L_HI(net1600));
 sg13g2_tiehi \cpu.dec.r_op[9]$_DFF_P__1601  (.L_HI(net1601));
 sg13g2_tiehi \cpu.dec.r_rd[0]$_DFFE_PP__1602  (.L_HI(net1602));
 sg13g2_tiehi \cpu.dec.r_rd[1]$_DFFE_PP__1603  (.L_HI(net1603));
 sg13g2_tiehi \cpu.dec.r_rd[2]$_DFFE_PP__1604  (.L_HI(net1604));
 sg13g2_tiehi \cpu.dec.r_rd[3]$_DFFE_PP__1605  (.L_HI(net1605));
 sg13g2_tiehi \cpu.dec.r_ready$_DFF_P__1606  (.L_HI(net1606));
 sg13g2_tiehi \cpu.dec.r_rs1[0]$_DFFE_PP__1607  (.L_HI(net1607));
 sg13g2_tiehi \cpu.dec.r_rs1[1]$_DFFE_PP__1608  (.L_HI(net1608));
 sg13g2_tiehi \cpu.dec.r_rs1[2]$_DFFE_PP__1609  (.L_HI(net1609));
 sg13g2_tiehi \cpu.dec.r_rs1[3]$_DFFE_PP__1610  (.L_HI(net1610));
 sg13g2_tiehi \cpu.dec.r_rs2[0]$_DFFE_PP__1611  (.L_HI(net1611));
 sg13g2_tiehi \cpu.dec.r_rs2[1]$_DFFE_PP__1612  (.L_HI(net1612));
 sg13g2_tiehi \cpu.dec.r_rs2[2]$_DFFE_PP__1613  (.L_HI(net1613));
 sg13g2_tiehi \cpu.dec.r_rs2[3]$_DFFE_PP__1614  (.L_HI(net1614));
 sg13g2_tiehi \cpu.dec.r_rs2_inv$_DFFE_PP__1615  (.L_HI(net1615));
 sg13g2_tiehi \cpu.dec.r_rs2_pc$_DFFE_PP__1616  (.L_HI(net1616));
 sg13g2_tiehi \cpu.dec.r_set_cc$_SDFFCE_PP0P__1617  (.L_HI(net1617));
 sg13g2_tiehi \cpu.dec.r_store$_DFFE_PP__1618  (.L_HI(net1618));
 sg13g2_tiehi \cpu.dec.r_swapsp$_DFFE_PP__1619  (.L_HI(net1619));
 sg13g2_tiehi \cpu.dec.r_sys_call$_DFFE_PP__1620  (.L_HI(net1620));
 sg13g2_tiehi \cpu.dec.r_trap$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P__1622  (.L_HI(net1622));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P__1623  (.L_HI(net1623));
 sg13g2_tiehi \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P__1624  (.L_HI(net1624));
 sg13g2_tiehi \cpu.ex.genblk3.r_supmode$_DFF_P__1625  (.L_HI(net1625));
 sg13g2_tiehi \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P__1626  (.L_HI(net1626));
 sg13g2_tiehi \cpu.ex.r_10[0]$_DFFE_PP__1627  (.L_HI(net1627));
 sg13g2_tiehi \cpu.ex.r_10[10]$_DFFE_PP__1628  (.L_HI(net1628));
 sg13g2_tiehi \cpu.ex.r_10[11]$_DFFE_PP__1629  (.L_HI(net1629));
 sg13g2_tiehi \cpu.ex.r_10[12]$_DFFE_PP__1630  (.L_HI(net1630));
 sg13g2_tiehi \cpu.ex.r_10[13]$_DFFE_PP__1631  (.L_HI(net1631));
 sg13g2_tiehi \cpu.ex.r_10[14]$_DFFE_PP__1632  (.L_HI(net1632));
 sg13g2_tiehi \cpu.ex.r_10[15]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \cpu.ex.r_10[1]$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \cpu.ex.r_10[2]$_DFFE_PP__1635  (.L_HI(net1635));
 sg13g2_tiehi \cpu.ex.r_10[3]$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \cpu.ex.r_10[4]$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \cpu.ex.r_10[5]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \cpu.ex.r_10[6]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \cpu.ex.r_10[7]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \cpu.ex.r_10[8]$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \cpu.ex.r_10[9]$_DFFE_PP__1642  (.L_HI(net1642));
 sg13g2_tiehi \cpu.ex.r_11[0]$_DFFE_PP__1643  (.L_HI(net1643));
 sg13g2_tiehi \cpu.ex.r_11[10]$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \cpu.ex.r_11[11]$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \cpu.ex.r_11[12]$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \cpu.ex.r_11[13]$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \cpu.ex.r_11[14]$_DFFE_PP__1648  (.L_HI(net1648));
 sg13g2_tiehi \cpu.ex.r_11[15]$_DFFE_PP__1649  (.L_HI(net1649));
 sg13g2_tiehi \cpu.ex.r_11[1]$_DFFE_PP__1650  (.L_HI(net1650));
 sg13g2_tiehi \cpu.ex.r_11[2]$_DFFE_PP__1651  (.L_HI(net1651));
 sg13g2_tiehi \cpu.ex.r_11[3]$_DFFE_PP__1652  (.L_HI(net1652));
 sg13g2_tiehi \cpu.ex.r_11[4]$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \cpu.ex.r_11[5]$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \cpu.ex.r_11[6]$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \cpu.ex.r_11[7]$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \cpu.ex.r_11[8]$_DFFE_PP__1657  (.L_HI(net1657));
 sg13g2_tiehi \cpu.ex.r_11[9]$_DFFE_PP__1658  (.L_HI(net1658));
 sg13g2_tiehi \cpu.ex.r_12[0]$_DFFE_PP__1659  (.L_HI(net1659));
 sg13g2_tiehi \cpu.ex.r_12[10]$_DFFE_PP__1660  (.L_HI(net1660));
 sg13g2_tiehi \cpu.ex.r_12[11]$_DFFE_PP__1661  (.L_HI(net1661));
 sg13g2_tiehi \cpu.ex.r_12[12]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \cpu.ex.r_12[13]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \cpu.ex.r_12[14]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \cpu.ex.r_12[15]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \cpu.ex.r_12[1]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \cpu.ex.r_12[2]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \cpu.ex.r_12[3]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \cpu.ex.r_12[4]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \cpu.ex.r_12[5]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \cpu.ex.r_12[6]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \cpu.ex.r_12[7]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \cpu.ex.r_12[8]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \cpu.ex.r_12[9]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \cpu.ex.r_13[0]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \cpu.ex.r_13[10]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \cpu.ex.r_13[11]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \cpu.ex.r_13[12]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \cpu.ex.r_13[13]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \cpu.ex.r_13[14]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \cpu.ex.r_13[15]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \cpu.ex.r_13[1]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \cpu.ex.r_13[2]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \cpu.ex.r_13[3]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \cpu.ex.r_13[4]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \cpu.ex.r_13[5]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \cpu.ex.r_13[6]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \cpu.ex.r_13[7]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \cpu.ex.r_13[8]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \cpu.ex.r_13[9]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \cpu.ex.r_14[0]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \cpu.ex.r_14[10]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \cpu.ex.r_14[11]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \cpu.ex.r_14[12]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \cpu.ex.r_14[13]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \cpu.ex.r_14[14]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \cpu.ex.r_14[15]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \cpu.ex.r_14[1]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \cpu.ex.r_14[2]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \cpu.ex.r_14[3]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \cpu.ex.r_14[4]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \cpu.ex.r_14[5]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \cpu.ex.r_14[6]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \cpu.ex.r_14[7]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \cpu.ex.r_14[8]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \cpu.ex.r_14[9]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \cpu.ex.r_15[0]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \cpu.ex.r_15[10]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \cpu.ex.r_15[11]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \cpu.ex.r_15[12]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \cpu.ex.r_15[13]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \cpu.ex.r_15[14]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \cpu.ex.r_15[15]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \cpu.ex.r_15[1]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \cpu.ex.r_15[2]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \cpu.ex.r_15[3]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \cpu.ex.r_15[4]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \cpu.ex.r_15[5]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \cpu.ex.r_15[6]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \cpu.ex.r_15[7]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \cpu.ex.r_15[8]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \cpu.ex.r_15[9]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \cpu.ex.r_8[0]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \cpu.ex.r_8[10]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \cpu.ex.r_8[11]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \cpu.ex.r_8[12]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \cpu.ex.r_8[13]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \cpu.ex.r_8[14]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \cpu.ex.r_8[15]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \cpu.ex.r_8[1]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \cpu.ex.r_8[2]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \cpu.ex.r_8[3]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \cpu.ex.r_8[4]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \cpu.ex.r_8[5]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \cpu.ex.r_8[6]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \cpu.ex.r_8[7]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \cpu.ex.r_8[8]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \cpu.ex.r_8[9]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \cpu.ex.r_9[0]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \cpu.ex.r_9[10]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \cpu.ex.r_9[11]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \cpu.ex.r_9[12]$_DFFE_PP__1742  (.L_HI(net1742));
 sg13g2_tiehi \cpu.ex.r_9[13]$_DFFE_PP__1743  (.L_HI(net1743));
 sg13g2_tiehi \cpu.ex.r_9[14]$_DFFE_PP__1744  (.L_HI(net1744));
 sg13g2_tiehi \cpu.ex.r_9[15]$_DFFE_PP__1745  (.L_HI(net1745));
 sg13g2_tiehi \cpu.ex.r_9[1]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \cpu.ex.r_9[2]$_DFFE_PP__1747  (.L_HI(net1747));
 sg13g2_tiehi \cpu.ex.r_9[3]$_DFFE_PP__1748  (.L_HI(net1748));
 sg13g2_tiehi \cpu.ex.r_9[4]$_DFFE_PP__1749  (.L_HI(net1749));
 sg13g2_tiehi \cpu.ex.r_9[5]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \cpu.ex.r_9[6]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \cpu.ex.r_9[7]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \cpu.ex.r_9[8]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \cpu.ex.r_9[9]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \cpu.ex.r_branch_stall$_DFF_P__1755  (.L_HI(net1755));
 sg13g2_tiehi \cpu.ex.r_cc$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \cpu.ex.r_d_flush_all$_SDFF_PP0__1757  (.L_HI(net1757));
 sg13g2_tiehi \cpu.ex.r_div_running$_DFF_P__1758  (.L_HI(net1758));
 sg13g2_tiehi \cpu.ex.r_epc[0]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \cpu.ex.r_epc[10]$_DFFE_PP__1760  (.L_HI(net1760));
 sg13g2_tiehi \cpu.ex.r_epc[11]$_DFFE_PP__1761  (.L_HI(net1761));
 sg13g2_tiehi \cpu.ex.r_epc[12]$_DFFE_PP__1762  (.L_HI(net1762));
 sg13g2_tiehi \cpu.ex.r_epc[13]$_DFFE_PP__1763  (.L_HI(net1763));
 sg13g2_tiehi \cpu.ex.r_epc[14]$_DFFE_PP__1764  (.L_HI(net1764));
 sg13g2_tiehi \cpu.ex.r_epc[1]$_DFFE_PP__1765  (.L_HI(net1765));
 sg13g2_tiehi \cpu.ex.r_epc[2]$_DFFE_PP__1766  (.L_HI(net1766));
 sg13g2_tiehi \cpu.ex.r_epc[3]$_DFFE_PP__1767  (.L_HI(net1767));
 sg13g2_tiehi \cpu.ex.r_epc[4]$_DFFE_PP__1768  (.L_HI(net1768));
 sg13g2_tiehi \cpu.ex.r_epc[5]$_DFFE_PP__1769  (.L_HI(net1769));
 sg13g2_tiehi \cpu.ex.r_epc[6]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \cpu.ex.r_epc[7]$_DFFE_PP__1771  (.L_HI(net1771));
 sg13g2_tiehi \cpu.ex.r_epc[8]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \cpu.ex.r_epc[9]$_DFFE_PP__1773  (.L_HI(net1773));
 sg13g2_tiehi \cpu.ex.r_fetch$_SDFF_PN1__1774  (.L_HI(net1774));
 sg13g2_tiehi \cpu.ex.r_flush_write$_SDFFE_PN0P__1775  (.L_HI(net1775));
 sg13g2_tiehi \cpu.ex.r_i_flush_all$_SDFF_PP0__1776  (.L_HI(net1776));
 sg13g2_tiehi \cpu.ex.r_ie$_SDFFE_PP0P__1777  (.L_HI(net1777));
 sg13g2_tiehi \cpu.ex.r_io_access$_SDFFE_PN0P__1778  (.L_HI(net1778));
 sg13g2_tiehi \cpu.ex.r_lr[0]$_DFFE_PP__1779  (.L_HI(net1779));
 sg13g2_tiehi \cpu.ex.r_lr[10]$_DFFE_PP__1780  (.L_HI(net1780));
 sg13g2_tiehi \cpu.ex.r_lr[11]$_DFFE_PP__1781  (.L_HI(net1781));
 sg13g2_tiehi \cpu.ex.r_lr[12]$_DFFE_PP__1782  (.L_HI(net1782));
 sg13g2_tiehi \cpu.ex.r_lr[13]$_DFFE_PP__1783  (.L_HI(net1783));
 sg13g2_tiehi \cpu.ex.r_lr[14]$_DFFE_PP__1784  (.L_HI(net1784));
 sg13g2_tiehi \cpu.ex.r_lr[1]$_DFFE_PP__1785  (.L_HI(net1785));
 sg13g2_tiehi \cpu.ex.r_lr[2]$_DFFE_PP__1786  (.L_HI(net1786));
 sg13g2_tiehi \cpu.ex.r_lr[3]$_DFFE_PP__1787  (.L_HI(net1787));
 sg13g2_tiehi \cpu.ex.r_lr[4]$_DFFE_PP__1788  (.L_HI(net1788));
 sg13g2_tiehi \cpu.ex.r_lr[5]$_DFFE_PP__1789  (.L_HI(net1789));
 sg13g2_tiehi \cpu.ex.r_lr[6]$_DFFE_PP__1790  (.L_HI(net1790));
 sg13g2_tiehi \cpu.ex.r_lr[7]$_DFFE_PP__1791  (.L_HI(net1791));
 sg13g2_tiehi \cpu.ex.r_lr[8]$_DFFE_PP__1792  (.L_HI(net1792));
 sg13g2_tiehi \cpu.ex.r_lr[9]$_DFFE_PP__1793  (.L_HI(net1793));
 sg13g2_tiehi \cpu.ex.r_mult[0]$_DFF_P__1794  (.L_HI(net1794));
 sg13g2_tiehi \cpu.ex.r_mult[10]$_DFF_P__1795  (.L_HI(net1795));
 sg13g2_tiehi \cpu.ex.r_mult[11]$_DFF_P__1796  (.L_HI(net1796));
 sg13g2_tiehi \cpu.ex.r_mult[12]$_DFF_P__1797  (.L_HI(net1797));
 sg13g2_tiehi \cpu.ex.r_mult[13]$_DFF_P__1798  (.L_HI(net1798));
 sg13g2_tiehi \cpu.ex.r_mult[14]$_DFF_P__1799  (.L_HI(net1799));
 sg13g2_tiehi \cpu.ex.r_mult[15]$_DFF_P__1800  (.L_HI(net1800));
 sg13g2_tiehi \cpu.ex.r_mult[16]$_DFFE_PP__1801  (.L_HI(net1801));
 sg13g2_tiehi \cpu.ex.r_mult[17]$_DFFE_PP__1802  (.L_HI(net1802));
 sg13g2_tiehi \cpu.ex.r_mult[18]$_DFFE_PP__1803  (.L_HI(net1803));
 sg13g2_tiehi \cpu.ex.r_mult[19]$_DFFE_PP__1804  (.L_HI(net1804));
 sg13g2_tiehi \cpu.ex.r_mult[1]$_DFF_P__1805  (.L_HI(net1805));
 sg13g2_tiehi \cpu.ex.r_mult[20]$_DFFE_PP__1806  (.L_HI(net1806));
 sg13g2_tiehi \cpu.ex.r_mult[21]$_DFFE_PP__1807  (.L_HI(net1807));
 sg13g2_tiehi \cpu.ex.r_mult[22]$_DFFE_PP__1808  (.L_HI(net1808));
 sg13g2_tiehi \cpu.ex.r_mult[23]$_DFFE_PP__1809  (.L_HI(net1809));
 sg13g2_tiehi \cpu.ex.r_mult[24]$_DFFE_PP__1810  (.L_HI(net1810));
 sg13g2_tiehi \cpu.ex.r_mult[25]$_DFFE_PP__1811  (.L_HI(net1811));
 sg13g2_tiehi \cpu.ex.r_mult[26]$_DFFE_PP__1812  (.L_HI(net1812));
 sg13g2_tiehi \cpu.ex.r_mult[27]$_DFFE_PP__1813  (.L_HI(net1813));
 sg13g2_tiehi \cpu.ex.r_mult[28]$_DFFE_PP__1814  (.L_HI(net1814));
 sg13g2_tiehi \cpu.ex.r_mult[29]$_DFFE_PP__1815  (.L_HI(net1815));
 sg13g2_tiehi \cpu.ex.r_mult[2]$_DFF_P__1816  (.L_HI(net1816));
 sg13g2_tiehi \cpu.ex.r_mult[30]$_DFFE_PP__1817  (.L_HI(net1817));
 sg13g2_tiehi \cpu.ex.r_mult[31]$_DFFE_PP__1818  (.L_HI(net1818));
 sg13g2_tiehi \cpu.ex.r_mult[3]$_DFF_P__1819  (.L_HI(net1819));
 sg13g2_tiehi \cpu.ex.r_mult[4]$_DFF_P__1820  (.L_HI(net1820));
 sg13g2_tiehi \cpu.ex.r_mult[5]$_DFF_P__1821  (.L_HI(net1821));
 sg13g2_tiehi \cpu.ex.r_mult[6]$_DFF_P__1822  (.L_HI(net1822));
 sg13g2_tiehi \cpu.ex.r_mult[7]$_DFF_P__1823  (.L_HI(net1823));
 sg13g2_tiehi \cpu.ex.r_mult[8]$_DFF_P__1824  (.L_HI(net1824));
 sg13g2_tiehi \cpu.ex.r_mult[9]$_DFF_P__1825  (.L_HI(net1825));
 sg13g2_tiehi \cpu.ex.r_mult_off[0]$_DFF_P__1826  (.L_HI(net1826));
 sg13g2_tiehi \cpu.ex.r_mult_off[1]$_DFF_P__1827  (.L_HI(net1827));
 sg13g2_tiehi \cpu.ex.r_mult_off[2]$_DFF_P__1828  (.L_HI(net1828));
 sg13g2_tiehi \cpu.ex.r_mult_off[3]$_DFF_P__1829  (.L_HI(net1829));
 sg13g2_tiehi \cpu.ex.r_mult_running$_DFF_P__1830  (.L_HI(net1830));
 sg13g2_tiehi \cpu.ex.r_pc[0]$_DFFE_PP__1831  (.L_HI(net1831));
 sg13g2_tiehi \cpu.ex.r_pc[10]$_DFFE_PP__1832  (.L_HI(net1832));
 sg13g2_tiehi \cpu.ex.r_pc[11]$_DFFE_PP__1833  (.L_HI(net1833));
 sg13g2_tiehi \cpu.ex.r_pc[12]$_DFFE_PP__1834  (.L_HI(net1834));
 sg13g2_tiehi \cpu.ex.r_pc[13]$_DFFE_PP__1835  (.L_HI(net1835));
 sg13g2_tiehi \cpu.ex.r_pc[14]$_DFFE_PP__1836  (.L_HI(net1836));
 sg13g2_tiehi \cpu.ex.r_pc[1]$_DFFE_PP__1837  (.L_HI(net1837));
 sg13g2_tiehi \cpu.ex.r_pc[2]$_DFFE_PP__1838  (.L_HI(net1838));
 sg13g2_tiehi \cpu.ex.r_pc[3]$_DFFE_PP__1839  (.L_HI(net1839));
 sg13g2_tiehi \cpu.ex.r_pc[4]$_DFFE_PP__1840  (.L_HI(net1840));
 sg13g2_tiehi \cpu.ex.r_pc[5]$_DFFE_PP__1841  (.L_HI(net1841));
 sg13g2_tiehi \cpu.ex.r_pc[6]$_DFFE_PP__1842  (.L_HI(net1842));
 sg13g2_tiehi \cpu.ex.r_pc[7]$_DFFE_PP__1843  (.L_HI(net1843));
 sg13g2_tiehi \cpu.ex.r_pc[8]$_DFFE_PP__1844  (.L_HI(net1844));
 sg13g2_tiehi \cpu.ex.r_pc[9]$_DFFE_PP__1845  (.L_HI(net1845));
 sg13g2_tiehi \cpu.ex.r_prev_ie$_SDFFE_PN0P__1846  (.L_HI(net1846));
 sg13g2_tiehi \cpu.ex.r_read_stall$_SDFFE_PN0P__1847  (.L_HI(net1847));
 sg13g2_tiehi \cpu.ex.r_set_cc$_DFFE_PP__1848  (.L_HI(net1848));
 sg13g2_tiehi \cpu.ex.r_sp[0]$_DFFE_PP__1849  (.L_HI(net1849));
 sg13g2_tiehi \cpu.ex.r_sp[10]$_DFFE_PP__1850  (.L_HI(net1850));
 sg13g2_tiehi \cpu.ex.r_sp[11]$_DFFE_PP__1851  (.L_HI(net1851));
 sg13g2_tiehi \cpu.ex.r_sp[12]$_DFFE_PP__1852  (.L_HI(net1852));
 sg13g2_tiehi \cpu.ex.r_sp[13]$_DFFE_PP__1853  (.L_HI(net1853));
 sg13g2_tiehi \cpu.ex.r_sp[14]$_DFFE_PP__1854  (.L_HI(net1854));
 sg13g2_tiehi \cpu.ex.r_sp[1]$_DFFE_PP__1855  (.L_HI(net1855));
 sg13g2_tiehi \cpu.ex.r_sp[2]$_DFFE_PP__1856  (.L_HI(net1856));
 sg13g2_tiehi \cpu.ex.r_sp[3]$_DFFE_PP__1857  (.L_HI(net1857));
 sg13g2_tiehi \cpu.ex.r_sp[4]$_DFFE_PP__1858  (.L_HI(net1858));
 sg13g2_tiehi \cpu.ex.r_sp[5]$_DFFE_PP__1859  (.L_HI(net1859));
 sg13g2_tiehi \cpu.ex.r_sp[6]$_DFFE_PP__1860  (.L_HI(net1860));
 sg13g2_tiehi \cpu.ex.r_sp[7]$_DFFE_PP__1861  (.L_HI(net1861));
 sg13g2_tiehi \cpu.ex.r_sp[8]$_DFFE_PP__1862  (.L_HI(net1862));
 sg13g2_tiehi \cpu.ex.r_sp[9]$_DFFE_PP__1863  (.L_HI(net1863));
 sg13g2_tiehi \cpu.ex.r_stmp[0]$_SDFFCE_PN0P__1864  (.L_HI(net1864));
 sg13g2_tiehi \cpu.ex.r_stmp[10]$_DFFE_PP__1865  (.L_HI(net1865));
 sg13g2_tiehi \cpu.ex.r_stmp[11]$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \cpu.ex.r_stmp[12]$_DFFE_PP__1867  (.L_HI(net1867));
 sg13g2_tiehi \cpu.ex.r_stmp[13]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \cpu.ex.r_stmp[14]$_DFFE_PP__1869  (.L_HI(net1869));
 sg13g2_tiehi \cpu.ex.r_stmp[15]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \cpu.ex.r_stmp[1]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \cpu.ex.r_stmp[2]$_DFFE_PP__1872  (.L_HI(net1872));
 sg13g2_tiehi \cpu.ex.r_stmp[3]$_DFFE_PP__1873  (.L_HI(net1873));
 sg13g2_tiehi \cpu.ex.r_stmp[4]$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \cpu.ex.r_stmp[5]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \cpu.ex.r_stmp[6]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \cpu.ex.r_stmp[7]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \cpu.ex.r_stmp[8]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \cpu.ex.r_stmp[9]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \cpu.ex.r_wb[0]$_DFFE_PP__1880  (.L_HI(net1880));
 sg13g2_tiehi \cpu.ex.r_wb[10]$_DFFE_PP__1881  (.L_HI(net1881));
 sg13g2_tiehi \cpu.ex.r_wb[11]$_DFFE_PP__1882  (.L_HI(net1882));
 sg13g2_tiehi \cpu.ex.r_wb[12]$_DFFE_PP__1883  (.L_HI(net1883));
 sg13g2_tiehi \cpu.ex.r_wb[13]$_DFFE_PP__1884  (.L_HI(net1884));
 sg13g2_tiehi \cpu.ex.r_wb[14]$_DFFE_PP__1885  (.L_HI(net1885));
 sg13g2_tiehi \cpu.ex.r_wb[15]$_DFFE_PP__1886  (.L_HI(net1886));
 sg13g2_tiehi \cpu.ex.r_wb[1]$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \cpu.ex.r_wb[2]$_DFFE_PP__1888  (.L_HI(net1888));
 sg13g2_tiehi \cpu.ex.r_wb[3]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \cpu.ex.r_wb[4]$_DFFE_PP__1890  (.L_HI(net1890));
 sg13g2_tiehi \cpu.ex.r_wb[5]$_DFFE_PP__1891  (.L_HI(net1891));
 sg13g2_tiehi \cpu.ex.r_wb[6]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \cpu.ex.r_wb[7]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \cpu.ex.r_wb[8]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \cpu.ex.r_wb[9]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P__1896  (.L_HI(net1896));
 sg13g2_tiehi \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P__1897  (.L_HI(net1897));
 sg13g2_tiehi \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P__1898  (.L_HI(net1898));
 sg13g2_tiehi \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P__1899  (.L_HI(net1899));
 sg13g2_tiehi \cpu.ex.r_wb_swapsp$_DFFE_PP__1900  (.L_HI(net1900));
 sg13g2_tiehi \cpu.ex.r_wb_valid$_DFF_P__1901  (.L_HI(net1901));
 sg13g2_tiehi \cpu.ex.r_wdata[0]$_DFFE_PP__1902  (.L_HI(net1902));
 sg13g2_tiehi \cpu.ex.r_wdata[10]$_DFFE_PP__1903  (.L_HI(net1903));
 sg13g2_tiehi \cpu.ex.r_wdata[11]$_DFFE_PP__1904  (.L_HI(net1904));
 sg13g2_tiehi \cpu.ex.r_wdata[12]$_DFFE_PP__1905  (.L_HI(net1905));
 sg13g2_tiehi \cpu.ex.r_wdata[13]$_DFFE_PP__1906  (.L_HI(net1906));
 sg13g2_tiehi \cpu.ex.r_wdata[14]$_DFFE_PP__1907  (.L_HI(net1907));
 sg13g2_tiehi \cpu.ex.r_wdata[15]$_DFFE_PP__1908  (.L_HI(net1908));
 sg13g2_tiehi \cpu.ex.r_wdata[1]$_DFFE_PP__1909  (.L_HI(net1909));
 sg13g2_tiehi \cpu.ex.r_wdata[2]$_DFFE_PP__1910  (.L_HI(net1910));
 sg13g2_tiehi \cpu.ex.r_wdata[3]$_DFFE_PP__1911  (.L_HI(net1911));
 sg13g2_tiehi \cpu.ex.r_wdata[4]$_DFFE_PP__1912  (.L_HI(net1912));
 sg13g2_tiehi \cpu.ex.r_wdata[5]$_DFFE_PP__1913  (.L_HI(net1913));
 sg13g2_tiehi \cpu.ex.r_wdata[6]$_DFFE_PP__1914  (.L_HI(net1914));
 sg13g2_tiehi \cpu.ex.r_wdata[7]$_DFFE_PP__1915  (.L_HI(net1915));
 sg13g2_tiehi \cpu.ex.r_wdata[8]$_DFFE_PP__1916  (.L_HI(net1916));
 sg13g2_tiehi \cpu.ex.r_wdata[9]$_DFFE_PP__1917  (.L_HI(net1917));
 sg13g2_tiehi \cpu.ex.r_wmask[0]$_SDFFE_PP0P__1918  (.L_HI(net1918));
 sg13g2_tiehi \cpu.ex.r_wmask[1]$_SDFFE_PP0P__1919  (.L_HI(net1919));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP__1920  (.L_HI(net1920));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP__1921  (.L_HI(net1921));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP__1922  (.L_HI(net1922));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP__1923  (.L_HI(net1923));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P__1924  (.L_HI(net1924));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P__1925  (.L_HI(net1925));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P__1926  (.L_HI(net1926));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P__1927  (.L_HI(net1927));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P__1928  (.L_HI(net1928));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P__1929  (.L_HI(net1929));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P__1930  (.L_HI(net1930));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P__1931  (.L_HI(net1931));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P__1932  (.L_HI(net1932));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P__1933  (.L_HI(net1933));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P__1934  (.L_HI(net1934));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P__1935  (.L_HI(net1935));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P__1936  (.L_HI(net1936));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P__1937  (.L_HI(net1937));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P__1938  (.L_HI(net1938));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P__1939  (.L_HI(net1939));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P__1940  (.L_HI(net1940));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P__1941  (.L_HI(net1941));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P__1942  (.L_HI(net1942));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P__1943  (.L_HI(net1943));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P__1944  (.L_HI(net1944));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P__1945  (.L_HI(net1945));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P__1946  (.L_HI(net1946));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P__1947  (.L_HI(net1947));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P__1948  (.L_HI(net1948));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P__1949  (.L_HI(net1949));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P__1950  (.L_HI(net1950));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P__1951  (.L_HI(net1951));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P__1952  (.L_HI(net1952));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P__1953  (.L_HI(net1953));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P__1954  (.L_HI(net1954));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P__1955  (.L_HI(net1955));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P__1956  (.L_HI(net1956));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P__1957  (.L_HI(net1957));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P__1958  (.L_HI(net1958));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P__1959  (.L_HI(net1959));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P__1964  (.L_HI(net1964));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P__1965  (.L_HI(net1965));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P__1966  (.L_HI(net1966));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P__1967  (.L_HI(net1967));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P__1978  (.L_HI(net1978));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P__1979  (.L_HI(net1979));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P__1980  (.L_HI(net1980));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P__1981  (.L_HI(net1981));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P__1982  (.L_HI(net1982));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P__1983  (.L_HI(net1983));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P__1984  (.L_HI(net1984));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P__1985  (.L_HI(net1985));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P__1986  (.L_HI(net1986));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P__1987  (.L_HI(net1987));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P__1988  (.L_HI(net1988));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P__1989  (.L_HI(net1989));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P__1990  (.L_HI(net1990));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP__1991  (.L_HI(net1991));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP__1992  (.L_HI(net1992));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP__1993  (.L_HI(net1993));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP__1994  (.L_HI(net1994));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP__1995  (.L_HI(net1995));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP__1996  (.L_HI(net1996));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP__1997  (.L_HI(net1997));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP__1998  (.L_HI(net1998));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP__1999  (.L_HI(net1999));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP__2000  (.L_HI(net2000));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP__2001  (.L_HI(net2001));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP__2002  (.L_HI(net2002));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP__2003  (.L_HI(net2003));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP__2004  (.L_HI(net2004));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP__2005  (.L_HI(net2005));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP__2006  (.L_HI(net2006));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP__2007  (.L_HI(net2007));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP__2008  (.L_HI(net2008));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP__2009  (.L_HI(net2009));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP__2010  (.L_HI(net2010));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP__2011  (.L_HI(net2011));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP__2012  (.L_HI(net2012));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP__2013  (.L_HI(net2013));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP__2014  (.L_HI(net2014));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP__2015  (.L_HI(net2015));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP__2016  (.L_HI(net2016));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP__2017  (.L_HI(net2017));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP__2018  (.L_HI(net2018));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP__2019  (.L_HI(net2019));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP__2020  (.L_HI(net2020));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP__2021  (.L_HI(net2021));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP__2022  (.L_HI(net2022));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP__2023  (.L_HI(net2023));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP__2024  (.L_HI(net2024));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP__2025  (.L_HI(net2025));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP__2026  (.L_HI(net2026));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP__2027  (.L_HI(net2027));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP__2028  (.L_HI(net2028));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP__2029  (.L_HI(net2029));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP__2030  (.L_HI(net2030));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP__2031  (.L_HI(net2031));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP__2032  (.L_HI(net2032));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP__2033  (.L_HI(net2033));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP__2034  (.L_HI(net2034));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP__2035  (.L_HI(net2035));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP__2036  (.L_HI(net2036));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP__2037  (.L_HI(net2037));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP__2038  (.L_HI(net2038));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP__2039  (.L_HI(net2039));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP__2040  (.L_HI(net2040));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP__2041  (.L_HI(net2041));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP__2042  (.L_HI(net2042));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP__2043  (.L_HI(net2043));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP__2044  (.L_HI(net2044));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP__2045  (.L_HI(net2045));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP__2046  (.L_HI(net2046));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP__2047  (.L_HI(net2047));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP__2048  (.L_HI(net2048));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP__2049  (.L_HI(net2049));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP__2050  (.L_HI(net2050));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP__2051  (.L_HI(net2051));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP__2052  (.L_HI(net2052));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP__2053  (.L_HI(net2053));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP__2054  (.L_HI(net2054));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP__2055  (.L_HI(net2055));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP__2056  (.L_HI(net2056));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP__2057  (.L_HI(net2057));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP__2058  (.L_HI(net2058));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP__2059  (.L_HI(net2059));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP__2060  (.L_HI(net2060));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP__2061  (.L_HI(net2061));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP__2062  (.L_HI(net2062));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP__2063  (.L_HI(net2063));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP__2064  (.L_HI(net2064));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP__2065  (.L_HI(net2065));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP__2066  (.L_HI(net2066));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP__2067  (.L_HI(net2067));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP__2068  (.L_HI(net2068));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP__2069  (.L_HI(net2069));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP__2070  (.L_HI(net2070));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP__2071  (.L_HI(net2071));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP__2072  (.L_HI(net2072));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP__2073  (.L_HI(net2073));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP__2074  (.L_HI(net2074));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP__2075  (.L_HI(net2075));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP__2076  (.L_HI(net2076));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP__2077  (.L_HI(net2077));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP__2078  (.L_HI(net2078));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP__2079  (.L_HI(net2079));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP__2080  (.L_HI(net2080));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP__2081  (.L_HI(net2081));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP__2082  (.L_HI(net2082));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP__2083  (.L_HI(net2083));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP__2084  (.L_HI(net2084));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP__2085  (.L_HI(net2085));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP__2086  (.L_HI(net2086));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP__2087  (.L_HI(net2087));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP__2088  (.L_HI(net2088));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP__2089  (.L_HI(net2089));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP__2090  (.L_HI(net2090));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP__2091  (.L_HI(net2091));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP__2092  (.L_HI(net2092));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP__2093  (.L_HI(net2093));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP__2094  (.L_HI(net2094));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP__2095  (.L_HI(net2095));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP__2096  (.L_HI(net2096));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP__2097  (.L_HI(net2097));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP__2098  (.L_HI(net2098));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP__2099  (.L_HI(net2099));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP__2100  (.L_HI(net2100));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP__2101  (.L_HI(net2101));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP__2102  (.L_HI(net2102));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP__2103  (.L_HI(net2103));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP__2104  (.L_HI(net2104));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP__2105  (.L_HI(net2105));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP__2106  (.L_HI(net2106));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP__2107  (.L_HI(net2107));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP__2108  (.L_HI(net2108));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP__2109  (.L_HI(net2109));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP__2110  (.L_HI(net2110));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP__2111  (.L_HI(net2111));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP__2112  (.L_HI(net2112));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP__2113  (.L_HI(net2113));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP__2114  (.L_HI(net2114));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP__2115  (.L_HI(net2115));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP__2116  (.L_HI(net2116));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP__2117  (.L_HI(net2117));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP__2118  (.L_HI(net2118));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP__2119  (.L_HI(net2119));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP__2120  (.L_HI(net2120));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP__2121  (.L_HI(net2121));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP__2122  (.L_HI(net2122));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP__2123  (.L_HI(net2123));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP__2124  (.L_HI(net2124));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP__2125  (.L_HI(net2125));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP__2126  (.L_HI(net2126));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP__2127  (.L_HI(net2127));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP__2128  (.L_HI(net2128));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP__2129  (.L_HI(net2129));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP__2130  (.L_HI(net2130));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP__2131  (.L_HI(net2131));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP__2132  (.L_HI(net2132));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP__2133  (.L_HI(net2133));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP__2134  (.L_HI(net2134));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP__2135  (.L_HI(net2135));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP__2136  (.L_HI(net2136));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP__2137  (.L_HI(net2137));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP__2138  (.L_HI(net2138));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP__2139  (.L_HI(net2139));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP__2140  (.L_HI(net2140));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP__2141  (.L_HI(net2141));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP__2142  (.L_HI(net2142));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP__2143  (.L_HI(net2143));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP__2144  (.L_HI(net2144));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP__2145  (.L_HI(net2145));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP__2146  (.L_HI(net2146));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP__2147  (.L_HI(net2147));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP__2148  (.L_HI(net2148));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP__2149  (.L_HI(net2149));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP__2150  (.L_HI(net2150));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP__2151  (.L_HI(net2151));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP__2152  (.L_HI(net2152));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP__2153  (.L_HI(net2153));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP__2154  (.L_HI(net2154));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP__2155  (.L_HI(net2155));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP__2156  (.L_HI(net2156));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP__2157  (.L_HI(net2157));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP__2158  (.L_HI(net2158));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP__2159  (.L_HI(net2159));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP__2160  (.L_HI(net2160));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP__2161  (.L_HI(net2161));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP__2162  (.L_HI(net2162));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP__2163  (.L_HI(net2163));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP__2164  (.L_HI(net2164));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP__2165  (.L_HI(net2165));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP__2166  (.L_HI(net2166));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP__2167  (.L_HI(net2167));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP__2168  (.L_HI(net2168));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP__2169  (.L_HI(net2169));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP__2170  (.L_HI(net2170));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP__2171  (.L_HI(net2171));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP__2172  (.L_HI(net2172));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP__2173  (.L_HI(net2173));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP__2174  (.L_HI(net2174));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP__2175  (.L_HI(net2175));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP__2176  (.L_HI(net2176));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP__2177  (.L_HI(net2177));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP__2178  (.L_HI(net2178));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP__2179  (.L_HI(net2179));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP__2180  (.L_HI(net2180));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP__2181  (.L_HI(net2181));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP__2182  (.L_HI(net2182));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP__2183  (.L_HI(net2183));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP__2184  (.L_HI(net2184));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP__2185  (.L_HI(net2185));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP__2186  (.L_HI(net2186));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP__2187  (.L_HI(net2187));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP__2188  (.L_HI(net2188));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP__2189  (.L_HI(net2189));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP__2190  (.L_HI(net2190));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP__2191  (.L_HI(net2191));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP__2192  (.L_HI(net2192));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP__2193  (.L_HI(net2193));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP__2194  (.L_HI(net2194));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP__2195  (.L_HI(net2195));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP__2196  (.L_HI(net2196));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP__2197  (.L_HI(net2197));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP__2198  (.L_HI(net2198));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP__2199  (.L_HI(net2199));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP__2200  (.L_HI(net2200));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP__2201  (.L_HI(net2201));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP__2202  (.L_HI(net2202));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP__2203  (.L_HI(net2203));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP__2204  (.L_HI(net2204));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP__2205  (.L_HI(net2205));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP__2206  (.L_HI(net2206));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP__2207  (.L_HI(net2207));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP__2208  (.L_HI(net2208));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP__2209  (.L_HI(net2209));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP__2210  (.L_HI(net2210));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP__2211  (.L_HI(net2211));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP__2212  (.L_HI(net2212));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP__2213  (.L_HI(net2213));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP__2214  (.L_HI(net2214));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP__2215  (.L_HI(net2215));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP__2216  (.L_HI(net2216));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP__2217  (.L_HI(net2217));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP__2218  (.L_HI(net2218));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP__2219  (.L_HI(net2219));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP__2220  (.L_HI(net2220));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP__2221  (.L_HI(net2221));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP__2222  (.L_HI(net2222));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP__2223  (.L_HI(net2223));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP__2224  (.L_HI(net2224));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP__2225  (.L_HI(net2225));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP__2226  (.L_HI(net2226));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP__2227  (.L_HI(net2227));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP__2228  (.L_HI(net2228));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP__2229  (.L_HI(net2229));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP__2230  (.L_HI(net2230));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP__2231  (.L_HI(net2231));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP__2232  (.L_HI(net2232));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP__2233  (.L_HI(net2233));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP__2234  (.L_HI(net2234));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP__2235  (.L_HI(net2235));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP__2236  (.L_HI(net2236));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP__2237  (.L_HI(net2237));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP__2238  (.L_HI(net2238));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP__2239  (.L_HI(net2239));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP__2240  (.L_HI(net2240));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP__2241  (.L_HI(net2241));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP__2242  (.L_HI(net2242));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP__2243  (.L_HI(net2243));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP__2244  (.L_HI(net2244));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP__2245  (.L_HI(net2245));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP__2246  (.L_HI(net2246));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP__2247  (.L_HI(net2247));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP__2248  (.L_HI(net2248));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP__2249  (.L_HI(net2249));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP__2250  (.L_HI(net2250));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP__2251  (.L_HI(net2251));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP__2252  (.L_HI(net2252));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP__2253  (.L_HI(net2253));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP__2254  (.L_HI(net2254));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP__2255  (.L_HI(net2255));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP__2256  (.L_HI(net2256));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP__2257  (.L_HI(net2257));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP__2258  (.L_HI(net2258));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP__2259  (.L_HI(net2259));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP__2260  (.L_HI(net2260));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP__2261  (.L_HI(net2261));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP__2262  (.L_HI(net2262));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP__2263  (.L_HI(net2263));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP__2264  (.L_HI(net2264));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP__2265  (.L_HI(net2265));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP__2266  (.L_HI(net2266));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP__2267  (.L_HI(net2267));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP__2268  (.L_HI(net2268));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP__2269  (.L_HI(net2269));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP__2270  (.L_HI(net2270));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP__2271  (.L_HI(net2271));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP__2272  (.L_HI(net2272));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP__2273  (.L_HI(net2273));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP__2274  (.L_HI(net2274));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP__2275  (.L_HI(net2275));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP__2276  (.L_HI(net2276));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP__2277  (.L_HI(net2277));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP__2278  (.L_HI(net2278));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP__2279  (.L_HI(net2279));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP__2280  (.L_HI(net2280));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP__2281  (.L_HI(net2281));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP__2282  (.L_HI(net2282));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP__2283  (.L_HI(net2283));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP__2284  (.L_HI(net2284));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP__2285  (.L_HI(net2285));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP__2286  (.L_HI(net2286));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP__2287  (.L_HI(net2287));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP__2288  (.L_HI(net2288));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP__2289  (.L_HI(net2289));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP__2290  (.L_HI(net2290));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP__2291  (.L_HI(net2291));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP__2292  (.L_HI(net2292));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP__2293  (.L_HI(net2293));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP__2294  (.L_HI(net2294));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP__2295  (.L_HI(net2295));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP__2296  (.L_HI(net2296));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP__2297  (.L_HI(net2297));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP__2298  (.L_HI(net2298));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP__2299  (.L_HI(net2299));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP__2300  (.L_HI(net2300));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP__2301  (.L_HI(net2301));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP__2302  (.L_HI(net2302));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP__2303  (.L_HI(net2303));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP__2304  (.L_HI(net2304));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP__2305  (.L_HI(net2305));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP__2306  (.L_HI(net2306));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP__2307  (.L_HI(net2307));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP__2308  (.L_HI(net2308));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP__2309  (.L_HI(net2309));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP__2310  (.L_HI(net2310));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP__2311  (.L_HI(net2311));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP__2312  (.L_HI(net2312));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP__2313  (.L_HI(net2313));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP__2314  (.L_HI(net2314));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP__2315  (.L_HI(net2315));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP__2316  (.L_HI(net2316));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP__2317  (.L_HI(net2317));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP__2318  (.L_HI(net2318));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP__2319  (.L_HI(net2319));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP__2320  (.L_HI(net2320));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP__2321  (.L_HI(net2321));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP__2322  (.L_HI(net2322));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP__2323  (.L_HI(net2323));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP__2324  (.L_HI(net2324));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP__2325  (.L_HI(net2325));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP__2326  (.L_HI(net2326));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP__2327  (.L_HI(net2327));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP__2328  (.L_HI(net2328));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP__2329  (.L_HI(net2329));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP__2330  (.L_HI(net2330));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP__2331  (.L_HI(net2331));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP__2332  (.L_HI(net2332));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP__2333  (.L_HI(net2333));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP__2334  (.L_HI(net2334));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP__2335  (.L_HI(net2335));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP__2336  (.L_HI(net2336));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP__2337  (.L_HI(net2337));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP__2338  (.L_HI(net2338));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP__2339  (.L_HI(net2339));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP__2340  (.L_HI(net2340));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP__2341  (.L_HI(net2341));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP__2342  (.L_HI(net2342));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP__2343  (.L_HI(net2343));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP__2344  (.L_HI(net2344));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP__2345  (.L_HI(net2345));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP__2346  (.L_HI(net2346));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP__2347  (.L_HI(net2347));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP__2348  (.L_HI(net2348));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP__2349  (.L_HI(net2349));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP__2350  (.L_HI(net2350));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP__2351  (.L_HI(net2351));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP__2352  (.L_HI(net2352));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP__2353  (.L_HI(net2353));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP__2354  (.L_HI(net2354));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP__2355  (.L_HI(net2355));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP__2356  (.L_HI(net2356));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP__2357  (.L_HI(net2357));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP__2358  (.L_HI(net2358));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP__2359  (.L_HI(net2359));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP__2360  (.L_HI(net2360));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP__2361  (.L_HI(net2361));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP__2362  (.L_HI(net2362));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP__2363  (.L_HI(net2363));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP__2364  (.L_HI(net2364));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP__2365  (.L_HI(net2365));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP__2366  (.L_HI(net2366));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP__2367  (.L_HI(net2367));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP__2368  (.L_HI(net2368));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP__2369  (.L_HI(net2369));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP__2370  (.L_HI(net2370));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP__2371  (.L_HI(net2371));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP__2372  (.L_HI(net2372));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP__2373  (.L_HI(net2373));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP__2374  (.L_HI(net2374));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP__2375  (.L_HI(net2375));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP__2376  (.L_HI(net2376));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP__2377  (.L_HI(net2377));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP__2378  (.L_HI(net2378));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP__2379  (.L_HI(net2379));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP__2380  (.L_HI(net2380));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP__2381  (.L_HI(net2381));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP__2382  (.L_HI(net2382));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP__2383  (.L_HI(net2383));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP__2384  (.L_HI(net2384));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP__2385  (.L_HI(net2385));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP__2386  (.L_HI(net2386));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP__2387  (.L_HI(net2387));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP__2388  (.L_HI(net2388));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP__2389  (.L_HI(net2389));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP__2390  (.L_HI(net2390));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP__2391  (.L_HI(net2391));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP__2392  (.L_HI(net2392));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP__2393  (.L_HI(net2393));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP__2394  (.L_HI(net2394));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP__2395  (.L_HI(net2395));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP__2396  (.L_HI(net2396));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP__2397  (.L_HI(net2397));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP__2398  (.L_HI(net2398));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP__2399  (.L_HI(net2399));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP__2400  (.L_HI(net2400));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP__2401  (.L_HI(net2401));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP__2402  (.L_HI(net2402));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP__2403  (.L_HI(net2403));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP__2404  (.L_HI(net2404));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP__2405  (.L_HI(net2405));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP__2406  (.L_HI(net2406));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP__2407  (.L_HI(net2407));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP__2408  (.L_HI(net2408));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP__2409  (.L_HI(net2409));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP__2410  (.L_HI(net2410));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP__2411  (.L_HI(net2411));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP__2412  (.L_HI(net2412));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP__2413  (.L_HI(net2413));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP__2414  (.L_HI(net2414));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP__2415  (.L_HI(net2415));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP__2416  (.L_HI(net2416));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP__2417  (.L_HI(net2417));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP__2418  (.L_HI(net2418));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP__2419  (.L_HI(net2419));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP__2420  (.L_HI(net2420));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP__2421  (.L_HI(net2421));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP__2422  (.L_HI(net2422));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP__2423  (.L_HI(net2423));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP__2424  (.L_HI(net2424));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP__2425  (.L_HI(net2425));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP__2426  (.L_HI(net2426));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP__2427  (.L_HI(net2427));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP__2428  (.L_HI(net2428));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP__2429  (.L_HI(net2429));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP__2430  (.L_HI(net2430));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP__2431  (.L_HI(net2431));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP__2432  (.L_HI(net2432));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP__2433  (.L_HI(net2433));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP__2434  (.L_HI(net2434));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP__2435  (.L_HI(net2435));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP__2436  (.L_HI(net2436));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP__2437  (.L_HI(net2437));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP__2438  (.L_HI(net2438));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP__2439  (.L_HI(net2439));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP__2440  (.L_HI(net2440));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP__2441  (.L_HI(net2441));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP__2442  (.L_HI(net2442));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP__2443  (.L_HI(net2443));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP__2444  (.L_HI(net2444));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP__2445  (.L_HI(net2445));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP__2446  (.L_HI(net2446));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP__2447  (.L_HI(net2447));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP__2448  (.L_HI(net2448));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP__2449  (.L_HI(net2449));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP__2450  (.L_HI(net2450));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP__2451  (.L_HI(net2451));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP__2452  (.L_HI(net2452));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP__2453  (.L_HI(net2453));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP__2454  (.L_HI(net2454));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP__2455  (.L_HI(net2455));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP__2456  (.L_HI(net2456));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP__2457  (.L_HI(net2457));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP__2458  (.L_HI(net2458));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP__2459  (.L_HI(net2459));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP__2460  (.L_HI(net2460));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP__2461  (.L_HI(net2461));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP__2462  (.L_HI(net2462));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP__2463  (.L_HI(net2463));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP__2464  (.L_HI(net2464));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP__2465  (.L_HI(net2465));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP__2466  (.L_HI(net2466));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP__2467  (.L_HI(net2467));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP__2468  (.L_HI(net2468));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP__2469  (.L_HI(net2469));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP__2470  (.L_HI(net2470));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP__2471  (.L_HI(net2471));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP__2472  (.L_HI(net2472));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP__2473  (.L_HI(net2473));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP__2474  (.L_HI(net2474));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP__2475  (.L_HI(net2475));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP__2476  (.L_HI(net2476));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP__2477  (.L_HI(net2477));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP__2478  (.L_HI(net2478));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP__2479  (.L_HI(net2479));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP__2480  (.L_HI(net2480));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP__2481  (.L_HI(net2481));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP__2482  (.L_HI(net2482));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP__2483  (.L_HI(net2483));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP__2484  (.L_HI(net2484));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP__2485  (.L_HI(net2485));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP__2486  (.L_HI(net2486));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP__2487  (.L_HI(net2487));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP__2488  (.L_HI(net2488));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP__2489  (.L_HI(net2489));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP__2490  (.L_HI(net2490));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP__2491  (.L_HI(net2491));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP__2492  (.L_HI(net2492));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP__2493  (.L_HI(net2493));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP__2494  (.L_HI(net2494));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP__2495  (.L_HI(net2495));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP__2496  (.L_HI(net2496));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP__2497  (.L_HI(net2497));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP__2498  (.L_HI(net2498));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP__2499  (.L_HI(net2499));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP__2500  (.L_HI(net2500));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP__2501  (.L_HI(net2501));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP__2502  (.L_HI(net2502));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP__2503  (.L_HI(net2503));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP__2504  (.L_HI(net2504));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP__2505  (.L_HI(net2505));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP__2506  (.L_HI(net2506));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP__2507  (.L_HI(net2507));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP__2508  (.L_HI(net2508));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP__2509  (.L_HI(net2509));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP__2510  (.L_HI(net2510));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP__2511  (.L_HI(net2511));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP__2512  (.L_HI(net2512));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP__2513  (.L_HI(net2513));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP__2514  (.L_HI(net2514));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP__2515  (.L_HI(net2515));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP__2516  (.L_HI(net2516));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP__2517  (.L_HI(net2517));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP__2518  (.L_HI(net2518));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP__2519  (.L_HI(net2519));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP__2520  (.L_HI(net2520));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP__2521  (.L_HI(net2521));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP__2522  (.L_HI(net2522));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP__2523  (.L_HI(net2523));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP__2524  (.L_HI(net2524));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP__2525  (.L_HI(net2525));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP__2526  (.L_HI(net2526));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP__2527  (.L_HI(net2527));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP__2528  (.L_HI(net2528));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP__2529  (.L_HI(net2529));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP__2530  (.L_HI(net2530));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP__2531  (.L_HI(net2531));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP__2532  (.L_HI(net2532));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP__2533  (.L_HI(net2533));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP__2534  (.L_HI(net2534));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP__2535  (.L_HI(net2535));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP__2536  (.L_HI(net2536));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP__2537  (.L_HI(net2537));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP__2538  (.L_HI(net2538));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP__2539  (.L_HI(net2539));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP__2540  (.L_HI(net2540));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP__2541  (.L_HI(net2541));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP__2542  (.L_HI(net2542));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP__2543  (.L_HI(net2543));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP__2544  (.L_HI(net2544));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP__2545  (.L_HI(net2545));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP__2546  (.L_HI(net2546));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP__2547  (.L_HI(net2547));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP__2548  (.L_HI(net2548));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP__2549  (.L_HI(net2549));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP__2550  (.L_HI(net2550));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP__2551  (.L_HI(net2551));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP__2552  (.L_HI(net2552));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP__2553  (.L_HI(net2553));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP__2554  (.L_HI(net2554));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP__2555  (.L_HI(net2555));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP__2556  (.L_HI(net2556));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP__2557  (.L_HI(net2557));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP__2558  (.L_HI(net2558));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP__2559  (.L_HI(net2559));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP__2560  (.L_HI(net2560));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP__2561  (.L_HI(net2561));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP__2562  (.L_HI(net2562));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP__2563  (.L_HI(net2563));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP__2564  (.L_HI(net2564));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP__2565  (.L_HI(net2565));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP__2566  (.L_HI(net2566));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP__2567  (.L_HI(net2567));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP__2568  (.L_HI(net2568));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP__2569  (.L_HI(net2569));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP__2570  (.L_HI(net2570));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP__2571  (.L_HI(net2571));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP__2572  (.L_HI(net2572));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP__2573  (.L_HI(net2573));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP__2574  (.L_HI(net2574));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP__2575  (.L_HI(net2575));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP__2576  (.L_HI(net2576));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP__2577  (.L_HI(net2577));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP__2578  (.L_HI(net2578));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP__2579  (.L_HI(net2579));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP__2580  (.L_HI(net2580));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP__2581  (.L_HI(net2581));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP__2582  (.L_HI(net2582));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP__2583  (.L_HI(net2583));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP__2584  (.L_HI(net2584));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP__2585  (.L_HI(net2585));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP__2586  (.L_HI(net2586));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP__2587  (.L_HI(net2587));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP__2588  (.L_HI(net2588));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP__2589  (.L_HI(net2589));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP__2590  (.L_HI(net2590));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP__2591  (.L_HI(net2591));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP__2592  (.L_HI(net2592));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP__2593  (.L_HI(net2593));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP__2594  (.L_HI(net2594));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP__2595  (.L_HI(net2595));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP__2596  (.L_HI(net2596));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP__2597  (.L_HI(net2597));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP__2598  (.L_HI(net2598));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP__2599  (.L_HI(net2599));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP__2600  (.L_HI(net2600));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP__2601  (.L_HI(net2601));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP__2602  (.L_HI(net2602));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP__2603  (.L_HI(net2603));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP__2604  (.L_HI(net2604));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP__2605  (.L_HI(net2605));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP__2606  (.L_HI(net2606));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP__2607  (.L_HI(net2607));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP__2608  (.L_HI(net2608));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP__2609  (.L_HI(net2609));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP__2610  (.L_HI(net2610));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP__2611  (.L_HI(net2611));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP__2612  (.L_HI(net2612));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP__2613  (.L_HI(net2613));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP__2614  (.L_HI(net2614));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP__2615  (.L_HI(net2615));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP__2616  (.L_HI(net2616));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP__2617  (.L_HI(net2617));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP__2618  (.L_HI(net2618));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP__2619  (.L_HI(net2619));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP__2620  (.L_HI(net2620));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP__2621  (.L_HI(net2621));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP__2622  (.L_HI(net2622));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP__2623  (.L_HI(net2623));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP__2624  (.L_HI(net2624));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP__2625  (.L_HI(net2625));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP__2626  (.L_HI(net2626));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP__2627  (.L_HI(net2627));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP__2628  (.L_HI(net2628));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP__2629  (.L_HI(net2629));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP__2630  (.L_HI(net2630));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP__2631  (.L_HI(net2631));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP__2632  (.L_HI(net2632));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP__2633  (.L_HI(net2633));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP__2634  (.L_HI(net2634));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP__2635  (.L_HI(net2635));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP__2636  (.L_HI(net2636));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP__2637  (.L_HI(net2637));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP__2638  (.L_HI(net2638));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP__2639  (.L_HI(net2639));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP__2640  (.L_HI(net2640));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP__2641  (.L_HI(net2641));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP__2642  (.L_HI(net2642));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP__2643  (.L_HI(net2643));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP__2644  (.L_HI(net2644));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP__2645  (.L_HI(net2645));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP__2646  (.L_HI(net2646));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP__2647  (.L_HI(net2647));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP__2648  (.L_HI(net2648));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP__2649  (.L_HI(net2649));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP__2650  (.L_HI(net2650));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP__2651  (.L_HI(net2651));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP__2652  (.L_HI(net2652));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP__2653  (.L_HI(net2653));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP__2654  (.L_HI(net2654));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP__2655  (.L_HI(net2655));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP__2656  (.L_HI(net2656));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP__2657  (.L_HI(net2657));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP__2658  (.L_HI(net2658));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP__2659  (.L_HI(net2659));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP__2660  (.L_HI(net2660));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP__2661  (.L_HI(net2661));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP__2662  (.L_HI(net2662));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP__2663  (.L_HI(net2663));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP__2664  (.L_HI(net2664));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP__2665  (.L_HI(net2665));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP__2666  (.L_HI(net2666));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP__2667  (.L_HI(net2667));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP__2668  (.L_HI(net2668));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP__2669  (.L_HI(net2669));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP__2670  (.L_HI(net2670));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP__2671  (.L_HI(net2671));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP__2672  (.L_HI(net2672));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP__2673  (.L_HI(net2673));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP__2674  (.L_HI(net2674));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP__2675  (.L_HI(net2675));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP__2676  (.L_HI(net2676));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP__2677  (.L_HI(net2677));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP__2678  (.L_HI(net2678));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP__2679  (.L_HI(net2679));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP__2680  (.L_HI(net2680));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP__2681  (.L_HI(net2681));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP__2682  (.L_HI(net2682));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP__2683  (.L_HI(net2683));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP__2684  (.L_HI(net2684));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP__2685  (.L_HI(net2685));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP__2686  (.L_HI(net2686));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP__2687  (.L_HI(net2687));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP__2688  (.L_HI(net2688));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP__2689  (.L_HI(net2689));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP__2690  (.L_HI(net2690));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP__2691  (.L_HI(net2691));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP__2692  (.L_HI(net2692));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP__2693  (.L_HI(net2693));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP__2694  (.L_HI(net2694));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP__2695  (.L_HI(net2695));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP__2696  (.L_HI(net2696));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP__2697  (.L_HI(net2697));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP__2698  (.L_HI(net2698));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP__2699  (.L_HI(net2699));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP__2700  (.L_HI(net2700));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP__2701  (.L_HI(net2701));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP__2702  (.L_HI(net2702));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP__2703  (.L_HI(net2703));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP__2704  (.L_HI(net2704));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP__2705  (.L_HI(net2705));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP__2706  (.L_HI(net2706));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP__2707  (.L_HI(net2707));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP__2708  (.L_HI(net2708));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP__2709  (.L_HI(net2709));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP__2710  (.L_HI(net2710));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP__2711  (.L_HI(net2711));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP__2712  (.L_HI(net2712));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP__2713  (.L_HI(net2713));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP__2714  (.L_HI(net2714));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP__2715  (.L_HI(net2715));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP__2716  (.L_HI(net2716));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP__2717  (.L_HI(net2717));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP__2718  (.L_HI(net2718));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP__2719  (.L_HI(net2719));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP__2720  (.L_HI(net2720));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP__2721  (.L_HI(net2721));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP__2722  (.L_HI(net2722));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP__2723  (.L_HI(net2723));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP__2724  (.L_HI(net2724));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP__2725  (.L_HI(net2725));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP__2726  (.L_HI(net2726));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP__2727  (.L_HI(net2727));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP__2728  (.L_HI(net2728));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP__2729  (.L_HI(net2729));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP__2730  (.L_HI(net2730));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP__2731  (.L_HI(net2731));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP__2732  (.L_HI(net2732));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP__2733  (.L_HI(net2733));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP__2734  (.L_HI(net2734));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP__2735  (.L_HI(net2735));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP__2736  (.L_HI(net2736));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP__2737  (.L_HI(net2737));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP__2738  (.L_HI(net2738));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP__2739  (.L_HI(net2739));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP__2740  (.L_HI(net2740));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP__2741  (.L_HI(net2741));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP__2742  (.L_HI(net2742));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP__2743  (.L_HI(net2743));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP__2744  (.L_HI(net2744));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP__2745  (.L_HI(net2745));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP__2746  (.L_HI(net2746));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP__2747  (.L_HI(net2747));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP__2748  (.L_HI(net2748));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP__2749  (.L_HI(net2749));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP__2750  (.L_HI(net2750));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP__2751  (.L_HI(net2751));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP__2752  (.L_HI(net2752));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP__2753  (.L_HI(net2753));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP__2754  (.L_HI(net2754));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP__2755  (.L_HI(net2755));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP__2756  (.L_HI(net2756));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP__2757  (.L_HI(net2757));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP__2758  (.L_HI(net2758));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP__2759  (.L_HI(net2759));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP__2760  (.L_HI(net2760));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP__2761  (.L_HI(net2761));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP__2762  (.L_HI(net2762));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP__2763  (.L_HI(net2763));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP__2764  (.L_HI(net2764));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP__2765  (.L_HI(net2765));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP__2766  (.L_HI(net2766));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP__2767  (.L_HI(net2767));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP__2768  (.L_HI(net2768));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP__2769  (.L_HI(net2769));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP__2770  (.L_HI(net2770));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP__2771  (.L_HI(net2771));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP__2772  (.L_HI(net2772));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP__2773  (.L_HI(net2773));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP__2774  (.L_HI(net2774));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP__2775  (.L_HI(net2775));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP__2776  (.L_HI(net2776));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP__2777  (.L_HI(net2777));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP__2778  (.L_HI(net2778));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP__2779  (.L_HI(net2779));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP__2780  (.L_HI(net2780));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP__2781  (.L_HI(net2781));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP__2782  (.L_HI(net2782));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP__2783  (.L_HI(net2783));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP__2784  (.L_HI(net2784));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP__2785  (.L_HI(net2785));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP__2786  (.L_HI(net2786));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP__2787  (.L_HI(net2787));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP__2788  (.L_HI(net2788));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP__2789  (.L_HI(net2789));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP__2790  (.L_HI(net2790));
 sg13g2_tiehi \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P__2791  (.L_HI(net2791));
 sg13g2_tiehi \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P__2792  (.L_HI(net2792));
 sg13g2_tiehi \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P__2793  (.L_HI(net2793));
 sg13g2_tiehi \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P__2794  (.L_HI(net2794));
 sg13g2_tiehi \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P__2795  (.L_HI(net2795));
 sg13g2_tiehi \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P__2796  (.L_HI(net2796));
 sg13g2_tiehi \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P__2797  (.L_HI(net2797));
 sg13g2_tiehi \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P__2798  (.L_HI(net2798));
 sg13g2_tiehi \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P__2799  (.L_HI(net2799));
 sg13g2_tiehi \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P__2800  (.L_HI(net2800));
 sg13g2_tiehi \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P__2801  (.L_HI(net2801));
 sg13g2_tiehi \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P__2802  (.L_HI(net2802));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P__2803  (.L_HI(net2803));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P__2804  (.L_HI(net2804));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P__2805  (.L_HI(net2805));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P__2806  (.L_HI(net2806));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[0]$_DFFE_PP__2807  (.L_HI(net2807));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[1]$_DFFE_PP__2808  (.L_HI(net2808));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[2]$_DFFE_PP__2809  (.L_HI(net2809));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[3]$_DFFE_PP__2810  (.L_HI(net2810));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[0]$_DFFE_PP__2811  (.L_HI(net2811));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[1]$_DFFE_PP__2812  (.L_HI(net2812));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[2]$_DFFE_PP__2813  (.L_HI(net2813));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[3]$_DFFE_PP__2814  (.L_HI(net2814));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[4]$_DFFE_PP__2815  (.L_HI(net2815));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP__2816  (.L_HI(net2816));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP__2817  (.L_HI(net2817));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP__2818  (.L_HI(net2818));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP__2819  (.L_HI(net2819));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP__2820  (.L_HI(net2820));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP__2821  (.L_HI(net2821));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP__2822  (.L_HI(net2822));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP__2823  (.L_HI(net2823));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][0]$_DFFE_PP__2824  (.L_HI(net2824));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][1]$_DFFE_PP__2825  (.L_HI(net2825));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][2]$_DFFE_PP__2826  (.L_HI(net2826));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][3]$_DFFE_PP__2827  (.L_HI(net2827));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][0]$_DFFE_PP__2828  (.L_HI(net2828));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][1]$_DFFE_PP__2829  (.L_HI(net2829));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][2]$_DFFE_PP__2830  (.L_HI(net2830));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][3]$_DFFE_PP__2831  (.L_HI(net2831));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][0]$_DFFE_PP__2832  (.L_HI(net2832));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][1]$_DFFE_PP__2833  (.L_HI(net2833));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][2]$_DFFE_PP__2834  (.L_HI(net2834));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][3]$_DFFE_PP__2835  (.L_HI(net2835));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][0]$_DFFE_PP__2836  (.L_HI(net2836));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][1]$_DFFE_PP__2837  (.L_HI(net2837));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][2]$_DFFE_PP__2838  (.L_HI(net2838));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][3]$_DFFE_PP__2839  (.L_HI(net2839));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][0]$_DFFE_PP__2840  (.L_HI(net2840));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][1]$_DFFE_PP__2841  (.L_HI(net2841));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][2]$_DFFE_PP__2842  (.L_HI(net2842));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][3]$_DFFE_PP__2843  (.L_HI(net2843));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][0]$_DFFE_PP__2844  (.L_HI(net2844));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][1]$_DFFE_PP__2845  (.L_HI(net2845));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][2]$_DFFE_PP__2846  (.L_HI(net2846));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][3]$_DFFE_PP__2847  (.L_HI(net2847));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][0]$_DFFE_PP__2848  (.L_HI(net2848));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][1]$_DFFE_PP__2849  (.L_HI(net2849));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][2]$_DFFE_PP__2850  (.L_HI(net2850));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][3]$_DFFE_PP__2851  (.L_HI(net2851));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P__2852  (.L_HI(net2852));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P__2853  (.L_HI(net2853));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P__2854  (.L_HI(net2854));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P__2855  (.L_HI(net2855));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][0]$_DFFE_PP__2856  (.L_HI(net2856));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][1]$_DFFE_PP__2857  (.L_HI(net2857));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][2]$_DFFE_PP__2858  (.L_HI(net2858));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][3]$_DFFE_PP__2859  (.L_HI(net2859));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P__2860  (.L_HI(net2860));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P__2861  (.L_HI(net2861));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P__2862  (.L_HI(net2862));
 sg13g2_tiehi \cpu.icache.r_data[0][0]$_DFFE_PP__2863  (.L_HI(net2863));
 sg13g2_tiehi \cpu.icache.r_data[0][10]$_DFFE_PP__2864  (.L_HI(net2864));
 sg13g2_tiehi \cpu.icache.r_data[0][11]$_DFFE_PP__2865  (.L_HI(net2865));
 sg13g2_tiehi \cpu.icache.r_data[0][12]$_DFFE_PP__2866  (.L_HI(net2866));
 sg13g2_tiehi \cpu.icache.r_data[0][13]$_DFFE_PP__2867  (.L_HI(net2867));
 sg13g2_tiehi \cpu.icache.r_data[0][14]$_DFFE_PP__2868  (.L_HI(net2868));
 sg13g2_tiehi \cpu.icache.r_data[0][15]$_DFFE_PP__2869  (.L_HI(net2869));
 sg13g2_tiehi \cpu.icache.r_data[0][16]$_DFFE_PP__2870  (.L_HI(net2870));
 sg13g2_tiehi \cpu.icache.r_data[0][17]$_DFFE_PP__2871  (.L_HI(net2871));
 sg13g2_tiehi \cpu.icache.r_data[0][18]$_DFFE_PP__2872  (.L_HI(net2872));
 sg13g2_tiehi \cpu.icache.r_data[0][19]$_DFFE_PP__2873  (.L_HI(net2873));
 sg13g2_tiehi \cpu.icache.r_data[0][1]$_DFFE_PP__2874  (.L_HI(net2874));
 sg13g2_tiehi \cpu.icache.r_data[0][20]$_DFFE_PP__2875  (.L_HI(net2875));
 sg13g2_tiehi \cpu.icache.r_data[0][21]$_DFFE_PP__2876  (.L_HI(net2876));
 sg13g2_tiehi \cpu.icache.r_data[0][22]$_DFFE_PP__2877  (.L_HI(net2877));
 sg13g2_tiehi \cpu.icache.r_data[0][23]$_DFFE_PP__2878  (.L_HI(net2878));
 sg13g2_tiehi \cpu.icache.r_data[0][24]$_DFFE_PP__2879  (.L_HI(net2879));
 sg13g2_tiehi \cpu.icache.r_data[0][25]$_DFFE_PP__2880  (.L_HI(net2880));
 sg13g2_tiehi \cpu.icache.r_data[0][26]$_DFFE_PP__2881  (.L_HI(net2881));
 sg13g2_tiehi \cpu.icache.r_data[0][27]$_DFFE_PP__2882  (.L_HI(net2882));
 sg13g2_tiehi \cpu.icache.r_data[0][28]$_DFFE_PP__2883  (.L_HI(net2883));
 sg13g2_tiehi \cpu.icache.r_data[0][29]$_DFFE_PP__2884  (.L_HI(net2884));
 sg13g2_tiehi \cpu.icache.r_data[0][2]$_DFFE_PP__2885  (.L_HI(net2885));
 sg13g2_tiehi \cpu.icache.r_data[0][30]$_DFFE_PP__2886  (.L_HI(net2886));
 sg13g2_tiehi \cpu.icache.r_data[0][31]$_DFFE_PP__2887  (.L_HI(net2887));
 sg13g2_tiehi \cpu.icache.r_data[0][3]$_DFFE_PP__2888  (.L_HI(net2888));
 sg13g2_tiehi \cpu.icache.r_data[0][4]$_DFFE_PP__2889  (.L_HI(net2889));
 sg13g2_tiehi \cpu.icache.r_data[0][5]$_DFFE_PP__2890  (.L_HI(net2890));
 sg13g2_tiehi \cpu.icache.r_data[0][6]$_DFFE_PP__2891  (.L_HI(net2891));
 sg13g2_tiehi \cpu.icache.r_data[0][7]$_DFFE_PP__2892  (.L_HI(net2892));
 sg13g2_tiehi \cpu.icache.r_data[0][8]$_DFFE_PP__2893  (.L_HI(net2893));
 sg13g2_tiehi \cpu.icache.r_data[0][9]$_DFFE_PP__2894  (.L_HI(net2894));
 sg13g2_tiehi \cpu.icache.r_data[1][0]$_DFFE_PP__2895  (.L_HI(net2895));
 sg13g2_tiehi \cpu.icache.r_data[1][10]$_DFFE_PP__2896  (.L_HI(net2896));
 sg13g2_tiehi \cpu.icache.r_data[1][11]$_DFFE_PP__2897  (.L_HI(net2897));
 sg13g2_tiehi \cpu.icache.r_data[1][12]$_DFFE_PP__2898  (.L_HI(net2898));
 sg13g2_tiehi \cpu.icache.r_data[1][13]$_DFFE_PP__2899  (.L_HI(net2899));
 sg13g2_tiehi \cpu.icache.r_data[1][14]$_DFFE_PP__2900  (.L_HI(net2900));
 sg13g2_tiehi \cpu.icache.r_data[1][15]$_DFFE_PP__2901  (.L_HI(net2901));
 sg13g2_tiehi \cpu.icache.r_data[1][16]$_DFFE_PP__2902  (.L_HI(net2902));
 sg13g2_tiehi \cpu.icache.r_data[1][17]$_DFFE_PP__2903  (.L_HI(net2903));
 sg13g2_tiehi \cpu.icache.r_data[1][18]$_DFFE_PP__2904  (.L_HI(net2904));
 sg13g2_tiehi \cpu.icache.r_data[1][19]$_DFFE_PP__2905  (.L_HI(net2905));
 sg13g2_tiehi \cpu.icache.r_data[1][1]$_DFFE_PP__2906  (.L_HI(net2906));
 sg13g2_tiehi \cpu.icache.r_data[1][20]$_DFFE_PP__2907  (.L_HI(net2907));
 sg13g2_tiehi \cpu.icache.r_data[1][21]$_DFFE_PP__2908  (.L_HI(net2908));
 sg13g2_tiehi \cpu.icache.r_data[1][22]$_DFFE_PP__2909  (.L_HI(net2909));
 sg13g2_tiehi \cpu.icache.r_data[1][23]$_DFFE_PP__2910  (.L_HI(net2910));
 sg13g2_tiehi \cpu.icache.r_data[1][24]$_DFFE_PP__2911  (.L_HI(net2911));
 sg13g2_tiehi \cpu.icache.r_data[1][25]$_DFFE_PP__2912  (.L_HI(net2912));
 sg13g2_tiehi \cpu.icache.r_data[1][26]$_DFFE_PP__2913  (.L_HI(net2913));
 sg13g2_tiehi \cpu.icache.r_data[1][27]$_DFFE_PP__2914  (.L_HI(net2914));
 sg13g2_tiehi \cpu.icache.r_data[1][28]$_DFFE_PP__2915  (.L_HI(net2915));
 sg13g2_tiehi \cpu.icache.r_data[1][29]$_DFFE_PP__2916  (.L_HI(net2916));
 sg13g2_tiehi \cpu.icache.r_data[1][2]$_DFFE_PP__2917  (.L_HI(net2917));
 sg13g2_tiehi \cpu.icache.r_data[1][30]$_DFFE_PP__2918  (.L_HI(net2918));
 sg13g2_tiehi \cpu.icache.r_data[1][31]$_DFFE_PP__2919  (.L_HI(net2919));
 sg13g2_tiehi \cpu.icache.r_data[1][3]$_DFFE_PP__2920  (.L_HI(net2920));
 sg13g2_tiehi \cpu.icache.r_data[1][4]$_DFFE_PP__2921  (.L_HI(net2921));
 sg13g2_tiehi \cpu.icache.r_data[1][5]$_DFFE_PP__2922  (.L_HI(net2922));
 sg13g2_tiehi \cpu.icache.r_data[1][6]$_DFFE_PP__2923  (.L_HI(net2923));
 sg13g2_tiehi \cpu.icache.r_data[1][7]$_DFFE_PP__2924  (.L_HI(net2924));
 sg13g2_tiehi \cpu.icache.r_data[1][8]$_DFFE_PP__2925  (.L_HI(net2925));
 sg13g2_tiehi \cpu.icache.r_data[1][9]$_DFFE_PP__2926  (.L_HI(net2926));
 sg13g2_tiehi \cpu.icache.r_data[2][0]$_DFFE_PP__2927  (.L_HI(net2927));
 sg13g2_tiehi \cpu.icache.r_data[2][10]$_DFFE_PP__2928  (.L_HI(net2928));
 sg13g2_tiehi \cpu.icache.r_data[2][11]$_DFFE_PP__2929  (.L_HI(net2929));
 sg13g2_tiehi \cpu.icache.r_data[2][12]$_DFFE_PP__2930  (.L_HI(net2930));
 sg13g2_tiehi \cpu.icache.r_data[2][13]$_DFFE_PP__2931  (.L_HI(net2931));
 sg13g2_tiehi \cpu.icache.r_data[2][14]$_DFFE_PP__2932  (.L_HI(net2932));
 sg13g2_tiehi \cpu.icache.r_data[2][15]$_DFFE_PP__2933  (.L_HI(net2933));
 sg13g2_tiehi \cpu.icache.r_data[2][16]$_DFFE_PP__2934  (.L_HI(net2934));
 sg13g2_tiehi \cpu.icache.r_data[2][17]$_DFFE_PP__2935  (.L_HI(net2935));
 sg13g2_tiehi \cpu.icache.r_data[2][18]$_DFFE_PP__2936  (.L_HI(net2936));
 sg13g2_tiehi \cpu.icache.r_data[2][19]$_DFFE_PP__2937  (.L_HI(net2937));
 sg13g2_tiehi \cpu.icache.r_data[2][1]$_DFFE_PP__2938  (.L_HI(net2938));
 sg13g2_tiehi \cpu.icache.r_data[2][20]$_DFFE_PP__2939  (.L_HI(net2939));
 sg13g2_tiehi \cpu.icache.r_data[2][21]$_DFFE_PP__2940  (.L_HI(net2940));
 sg13g2_tiehi \cpu.icache.r_data[2][22]$_DFFE_PP__2941  (.L_HI(net2941));
 sg13g2_tiehi \cpu.icache.r_data[2][23]$_DFFE_PP__2942  (.L_HI(net2942));
 sg13g2_tiehi \cpu.icache.r_data[2][24]$_DFFE_PP__2943  (.L_HI(net2943));
 sg13g2_tiehi \cpu.icache.r_data[2][25]$_DFFE_PP__2944  (.L_HI(net2944));
 sg13g2_tiehi \cpu.icache.r_data[2][26]$_DFFE_PP__2945  (.L_HI(net2945));
 sg13g2_tiehi \cpu.icache.r_data[2][27]$_DFFE_PP__2946  (.L_HI(net2946));
 sg13g2_tiehi \cpu.icache.r_data[2][28]$_DFFE_PP__2947  (.L_HI(net2947));
 sg13g2_tiehi \cpu.icache.r_data[2][29]$_DFFE_PP__2948  (.L_HI(net2948));
 sg13g2_tiehi \cpu.icache.r_data[2][2]$_DFFE_PP__2949  (.L_HI(net2949));
 sg13g2_tiehi \cpu.icache.r_data[2][30]$_DFFE_PP__2950  (.L_HI(net2950));
 sg13g2_tiehi \cpu.icache.r_data[2][31]$_DFFE_PP__2951  (.L_HI(net2951));
 sg13g2_tiehi \cpu.icache.r_data[2][3]$_DFFE_PP__2952  (.L_HI(net2952));
 sg13g2_tiehi \cpu.icache.r_data[2][4]$_DFFE_PP__2953  (.L_HI(net2953));
 sg13g2_tiehi \cpu.icache.r_data[2][5]$_DFFE_PP__2954  (.L_HI(net2954));
 sg13g2_tiehi \cpu.icache.r_data[2][6]$_DFFE_PP__2955  (.L_HI(net2955));
 sg13g2_tiehi \cpu.icache.r_data[2][7]$_DFFE_PP__2956  (.L_HI(net2956));
 sg13g2_tiehi \cpu.icache.r_data[2][8]$_DFFE_PP__2957  (.L_HI(net2957));
 sg13g2_tiehi \cpu.icache.r_data[2][9]$_DFFE_PP__2958  (.L_HI(net2958));
 sg13g2_tiehi \cpu.icache.r_data[3][0]$_DFFE_PP__2959  (.L_HI(net2959));
 sg13g2_tiehi \cpu.icache.r_data[3][10]$_DFFE_PP__2960  (.L_HI(net2960));
 sg13g2_tiehi \cpu.icache.r_data[3][11]$_DFFE_PP__2961  (.L_HI(net2961));
 sg13g2_tiehi \cpu.icache.r_data[3][12]$_DFFE_PP__2962  (.L_HI(net2962));
 sg13g2_tiehi \cpu.icache.r_data[3][13]$_DFFE_PP__2963  (.L_HI(net2963));
 sg13g2_tiehi \cpu.icache.r_data[3][14]$_DFFE_PP__2964  (.L_HI(net2964));
 sg13g2_tiehi \cpu.icache.r_data[3][15]$_DFFE_PP__2965  (.L_HI(net2965));
 sg13g2_tiehi \cpu.icache.r_data[3][16]$_DFFE_PP__2966  (.L_HI(net2966));
 sg13g2_tiehi \cpu.icache.r_data[3][17]$_DFFE_PP__2967  (.L_HI(net2967));
 sg13g2_tiehi \cpu.icache.r_data[3][18]$_DFFE_PP__2968  (.L_HI(net2968));
 sg13g2_tiehi \cpu.icache.r_data[3][19]$_DFFE_PP__2969  (.L_HI(net2969));
 sg13g2_tiehi \cpu.icache.r_data[3][1]$_DFFE_PP__2970  (.L_HI(net2970));
 sg13g2_tiehi \cpu.icache.r_data[3][20]$_DFFE_PP__2971  (.L_HI(net2971));
 sg13g2_tiehi \cpu.icache.r_data[3][21]$_DFFE_PP__2972  (.L_HI(net2972));
 sg13g2_tiehi \cpu.icache.r_data[3][22]$_DFFE_PP__2973  (.L_HI(net2973));
 sg13g2_tiehi \cpu.icache.r_data[3][23]$_DFFE_PP__2974  (.L_HI(net2974));
 sg13g2_tiehi \cpu.icache.r_data[3][24]$_DFFE_PP__2975  (.L_HI(net2975));
 sg13g2_tiehi \cpu.icache.r_data[3][25]$_DFFE_PP__2976  (.L_HI(net2976));
 sg13g2_tiehi \cpu.icache.r_data[3][26]$_DFFE_PP__2977  (.L_HI(net2977));
 sg13g2_tiehi \cpu.icache.r_data[3][27]$_DFFE_PP__2978  (.L_HI(net2978));
 sg13g2_tiehi \cpu.icache.r_data[3][28]$_DFFE_PP__2979  (.L_HI(net2979));
 sg13g2_tiehi \cpu.icache.r_data[3][29]$_DFFE_PP__2980  (.L_HI(net2980));
 sg13g2_tiehi \cpu.icache.r_data[3][2]$_DFFE_PP__2981  (.L_HI(net2981));
 sg13g2_tiehi \cpu.icache.r_data[3][30]$_DFFE_PP__2982  (.L_HI(net2982));
 sg13g2_tiehi \cpu.icache.r_data[3][31]$_DFFE_PP__2983  (.L_HI(net2983));
 sg13g2_tiehi \cpu.icache.r_data[3][3]$_DFFE_PP__2984  (.L_HI(net2984));
 sg13g2_tiehi \cpu.icache.r_data[3][4]$_DFFE_PP__2985  (.L_HI(net2985));
 sg13g2_tiehi \cpu.icache.r_data[3][5]$_DFFE_PP__2986  (.L_HI(net2986));
 sg13g2_tiehi \cpu.icache.r_data[3][6]$_DFFE_PP__2987  (.L_HI(net2987));
 sg13g2_tiehi \cpu.icache.r_data[3][7]$_DFFE_PP__2988  (.L_HI(net2988));
 sg13g2_tiehi \cpu.icache.r_data[3][8]$_DFFE_PP__2989  (.L_HI(net2989));
 sg13g2_tiehi \cpu.icache.r_data[3][9]$_DFFE_PP__2990  (.L_HI(net2990));
 sg13g2_tiehi \cpu.icache.r_data[4][0]$_DFFE_PP__2991  (.L_HI(net2991));
 sg13g2_tiehi \cpu.icache.r_data[4][10]$_DFFE_PP__2992  (.L_HI(net2992));
 sg13g2_tiehi \cpu.icache.r_data[4][11]$_DFFE_PP__2993  (.L_HI(net2993));
 sg13g2_tiehi \cpu.icache.r_data[4][12]$_DFFE_PP__2994  (.L_HI(net2994));
 sg13g2_tiehi \cpu.icache.r_data[4][13]$_DFFE_PP__2995  (.L_HI(net2995));
 sg13g2_tiehi \cpu.icache.r_data[4][14]$_DFFE_PP__2996  (.L_HI(net2996));
 sg13g2_tiehi \cpu.icache.r_data[4][15]$_DFFE_PP__2997  (.L_HI(net2997));
 sg13g2_tiehi \cpu.icache.r_data[4][16]$_DFFE_PP__2998  (.L_HI(net2998));
 sg13g2_tiehi \cpu.icache.r_data[4][17]$_DFFE_PP__2999  (.L_HI(net2999));
 sg13g2_tiehi \cpu.icache.r_data[4][18]$_DFFE_PP__3000  (.L_HI(net3000));
 sg13g2_tiehi \cpu.icache.r_data[4][19]$_DFFE_PP__3001  (.L_HI(net3001));
 sg13g2_tiehi \cpu.icache.r_data[4][1]$_DFFE_PP__3002  (.L_HI(net3002));
 sg13g2_tiehi \cpu.icache.r_data[4][20]$_DFFE_PP__3003  (.L_HI(net3003));
 sg13g2_tiehi \cpu.icache.r_data[4][21]$_DFFE_PP__3004  (.L_HI(net3004));
 sg13g2_tiehi \cpu.icache.r_data[4][22]$_DFFE_PP__3005  (.L_HI(net3005));
 sg13g2_tiehi \cpu.icache.r_data[4][23]$_DFFE_PP__3006  (.L_HI(net3006));
 sg13g2_tiehi \cpu.icache.r_data[4][24]$_DFFE_PP__3007  (.L_HI(net3007));
 sg13g2_tiehi \cpu.icache.r_data[4][25]$_DFFE_PP__3008  (.L_HI(net3008));
 sg13g2_tiehi \cpu.icache.r_data[4][26]$_DFFE_PP__3009  (.L_HI(net3009));
 sg13g2_tiehi \cpu.icache.r_data[4][27]$_DFFE_PP__3010  (.L_HI(net3010));
 sg13g2_tiehi \cpu.icache.r_data[4][28]$_DFFE_PP__3011  (.L_HI(net3011));
 sg13g2_tiehi \cpu.icache.r_data[4][29]$_DFFE_PP__3012  (.L_HI(net3012));
 sg13g2_tiehi \cpu.icache.r_data[4][2]$_DFFE_PP__3013  (.L_HI(net3013));
 sg13g2_tiehi \cpu.icache.r_data[4][30]$_DFFE_PP__3014  (.L_HI(net3014));
 sg13g2_tiehi \cpu.icache.r_data[4][31]$_DFFE_PP__3015  (.L_HI(net3015));
 sg13g2_tiehi \cpu.icache.r_data[4][3]$_DFFE_PP__3016  (.L_HI(net3016));
 sg13g2_tiehi \cpu.icache.r_data[4][4]$_DFFE_PP__3017  (.L_HI(net3017));
 sg13g2_tiehi \cpu.icache.r_data[4][5]$_DFFE_PP__3018  (.L_HI(net3018));
 sg13g2_tiehi \cpu.icache.r_data[4][6]$_DFFE_PP__3019  (.L_HI(net3019));
 sg13g2_tiehi \cpu.icache.r_data[4][7]$_DFFE_PP__3020  (.L_HI(net3020));
 sg13g2_tiehi \cpu.icache.r_data[4][8]$_DFFE_PP__3021  (.L_HI(net3021));
 sg13g2_tiehi \cpu.icache.r_data[4][9]$_DFFE_PP__3022  (.L_HI(net3022));
 sg13g2_tiehi \cpu.icache.r_data[5][0]$_DFFE_PP__3023  (.L_HI(net3023));
 sg13g2_tiehi \cpu.icache.r_data[5][10]$_DFFE_PP__3024  (.L_HI(net3024));
 sg13g2_tiehi \cpu.icache.r_data[5][11]$_DFFE_PP__3025  (.L_HI(net3025));
 sg13g2_tiehi \cpu.icache.r_data[5][12]$_DFFE_PP__3026  (.L_HI(net3026));
 sg13g2_tiehi \cpu.icache.r_data[5][13]$_DFFE_PP__3027  (.L_HI(net3027));
 sg13g2_tiehi \cpu.icache.r_data[5][14]$_DFFE_PP__3028  (.L_HI(net3028));
 sg13g2_tiehi \cpu.icache.r_data[5][15]$_DFFE_PP__3029  (.L_HI(net3029));
 sg13g2_tiehi \cpu.icache.r_data[5][16]$_DFFE_PP__3030  (.L_HI(net3030));
 sg13g2_tiehi \cpu.icache.r_data[5][17]$_DFFE_PP__3031  (.L_HI(net3031));
 sg13g2_tiehi \cpu.icache.r_data[5][18]$_DFFE_PP__3032  (.L_HI(net3032));
 sg13g2_tiehi \cpu.icache.r_data[5][19]$_DFFE_PP__3033  (.L_HI(net3033));
 sg13g2_tiehi \cpu.icache.r_data[5][1]$_DFFE_PP__3034  (.L_HI(net3034));
 sg13g2_tiehi \cpu.icache.r_data[5][20]$_DFFE_PP__3035  (.L_HI(net3035));
 sg13g2_tiehi \cpu.icache.r_data[5][21]$_DFFE_PP__3036  (.L_HI(net3036));
 sg13g2_tiehi \cpu.icache.r_data[5][22]$_DFFE_PP__3037  (.L_HI(net3037));
 sg13g2_tiehi \cpu.icache.r_data[5][23]$_DFFE_PP__3038  (.L_HI(net3038));
 sg13g2_tiehi \cpu.icache.r_data[5][24]$_DFFE_PP__3039  (.L_HI(net3039));
 sg13g2_tiehi \cpu.icache.r_data[5][25]$_DFFE_PP__3040  (.L_HI(net3040));
 sg13g2_tiehi \cpu.icache.r_data[5][26]$_DFFE_PP__3041  (.L_HI(net3041));
 sg13g2_tiehi \cpu.icache.r_data[5][27]$_DFFE_PP__3042  (.L_HI(net3042));
 sg13g2_tiehi \cpu.icache.r_data[5][28]$_DFFE_PP__3043  (.L_HI(net3043));
 sg13g2_tiehi \cpu.icache.r_data[5][29]$_DFFE_PP__3044  (.L_HI(net3044));
 sg13g2_tiehi \cpu.icache.r_data[5][2]$_DFFE_PP__3045  (.L_HI(net3045));
 sg13g2_tiehi \cpu.icache.r_data[5][30]$_DFFE_PP__3046  (.L_HI(net3046));
 sg13g2_tiehi \cpu.icache.r_data[5][31]$_DFFE_PP__3047  (.L_HI(net3047));
 sg13g2_tiehi \cpu.icache.r_data[5][3]$_DFFE_PP__3048  (.L_HI(net3048));
 sg13g2_tiehi \cpu.icache.r_data[5][4]$_DFFE_PP__3049  (.L_HI(net3049));
 sg13g2_tiehi \cpu.icache.r_data[5][5]$_DFFE_PP__3050  (.L_HI(net3050));
 sg13g2_tiehi \cpu.icache.r_data[5][6]$_DFFE_PP__3051  (.L_HI(net3051));
 sg13g2_tiehi \cpu.icache.r_data[5][7]$_DFFE_PP__3052  (.L_HI(net3052));
 sg13g2_tiehi \cpu.icache.r_data[5][8]$_DFFE_PP__3053  (.L_HI(net3053));
 sg13g2_tiehi \cpu.icache.r_data[5][9]$_DFFE_PP__3054  (.L_HI(net3054));
 sg13g2_tiehi \cpu.icache.r_data[6][0]$_DFFE_PP__3055  (.L_HI(net3055));
 sg13g2_tiehi \cpu.icache.r_data[6][10]$_DFFE_PP__3056  (.L_HI(net3056));
 sg13g2_tiehi \cpu.icache.r_data[6][11]$_DFFE_PP__3057  (.L_HI(net3057));
 sg13g2_tiehi \cpu.icache.r_data[6][12]$_DFFE_PP__3058  (.L_HI(net3058));
 sg13g2_tiehi \cpu.icache.r_data[6][13]$_DFFE_PP__3059  (.L_HI(net3059));
 sg13g2_tiehi \cpu.icache.r_data[6][14]$_DFFE_PP__3060  (.L_HI(net3060));
 sg13g2_tiehi \cpu.icache.r_data[6][15]$_DFFE_PP__3061  (.L_HI(net3061));
 sg13g2_tiehi \cpu.icache.r_data[6][16]$_DFFE_PP__3062  (.L_HI(net3062));
 sg13g2_tiehi \cpu.icache.r_data[6][17]$_DFFE_PP__3063  (.L_HI(net3063));
 sg13g2_tiehi \cpu.icache.r_data[6][18]$_DFFE_PP__3064  (.L_HI(net3064));
 sg13g2_tiehi \cpu.icache.r_data[6][19]$_DFFE_PP__3065  (.L_HI(net3065));
 sg13g2_tiehi \cpu.icache.r_data[6][1]$_DFFE_PP__3066  (.L_HI(net3066));
 sg13g2_tiehi \cpu.icache.r_data[6][20]$_DFFE_PP__3067  (.L_HI(net3067));
 sg13g2_tiehi \cpu.icache.r_data[6][21]$_DFFE_PP__3068  (.L_HI(net3068));
 sg13g2_tiehi \cpu.icache.r_data[6][22]$_DFFE_PP__3069  (.L_HI(net3069));
 sg13g2_tiehi \cpu.icache.r_data[6][23]$_DFFE_PP__3070  (.L_HI(net3070));
 sg13g2_tiehi \cpu.icache.r_data[6][24]$_DFFE_PP__3071  (.L_HI(net3071));
 sg13g2_tiehi \cpu.icache.r_data[6][25]$_DFFE_PP__3072  (.L_HI(net3072));
 sg13g2_tiehi \cpu.icache.r_data[6][26]$_DFFE_PP__3073  (.L_HI(net3073));
 sg13g2_tiehi \cpu.icache.r_data[6][27]$_DFFE_PP__3074  (.L_HI(net3074));
 sg13g2_tiehi \cpu.icache.r_data[6][28]$_DFFE_PP__3075  (.L_HI(net3075));
 sg13g2_tiehi \cpu.icache.r_data[6][29]$_DFFE_PP__3076  (.L_HI(net3076));
 sg13g2_tiehi \cpu.icache.r_data[6][2]$_DFFE_PP__3077  (.L_HI(net3077));
 sg13g2_tiehi \cpu.icache.r_data[6][30]$_DFFE_PP__3078  (.L_HI(net3078));
 sg13g2_tiehi \cpu.icache.r_data[6][31]$_DFFE_PP__3079  (.L_HI(net3079));
 sg13g2_tiehi \cpu.icache.r_data[6][3]$_DFFE_PP__3080  (.L_HI(net3080));
 sg13g2_tiehi \cpu.icache.r_data[6][4]$_DFFE_PP__3081  (.L_HI(net3081));
 sg13g2_tiehi \cpu.icache.r_data[6][5]$_DFFE_PP__3082  (.L_HI(net3082));
 sg13g2_tiehi \cpu.icache.r_data[6][6]$_DFFE_PP__3083  (.L_HI(net3083));
 sg13g2_tiehi \cpu.icache.r_data[6][7]$_DFFE_PP__3084  (.L_HI(net3084));
 sg13g2_tiehi \cpu.icache.r_data[6][8]$_DFFE_PP__3085  (.L_HI(net3085));
 sg13g2_tiehi \cpu.icache.r_data[6][9]$_DFFE_PP__3086  (.L_HI(net3086));
 sg13g2_tiehi \cpu.icache.r_data[7][0]$_DFFE_PP__3087  (.L_HI(net3087));
 sg13g2_tiehi \cpu.icache.r_data[7][10]$_DFFE_PP__3088  (.L_HI(net3088));
 sg13g2_tiehi \cpu.icache.r_data[7][11]$_DFFE_PP__3089  (.L_HI(net3089));
 sg13g2_tiehi \cpu.icache.r_data[7][12]$_DFFE_PP__3090  (.L_HI(net3090));
 sg13g2_tiehi \cpu.icache.r_data[7][13]$_DFFE_PP__3091  (.L_HI(net3091));
 sg13g2_tiehi \cpu.icache.r_data[7][14]$_DFFE_PP__3092  (.L_HI(net3092));
 sg13g2_tiehi \cpu.icache.r_data[7][15]$_DFFE_PP__3093  (.L_HI(net3093));
 sg13g2_tiehi \cpu.icache.r_data[7][16]$_DFFE_PP__3094  (.L_HI(net3094));
 sg13g2_tiehi \cpu.icache.r_data[7][17]$_DFFE_PP__3095  (.L_HI(net3095));
 sg13g2_tiehi \cpu.icache.r_data[7][18]$_DFFE_PP__3096  (.L_HI(net3096));
 sg13g2_tiehi \cpu.icache.r_data[7][19]$_DFFE_PP__3097  (.L_HI(net3097));
 sg13g2_tiehi \cpu.icache.r_data[7][1]$_DFFE_PP__3098  (.L_HI(net3098));
 sg13g2_tiehi \cpu.icache.r_data[7][20]$_DFFE_PP__3099  (.L_HI(net3099));
 sg13g2_tiehi \cpu.icache.r_data[7][21]$_DFFE_PP__3100  (.L_HI(net3100));
 sg13g2_tiehi \cpu.icache.r_data[7][22]$_DFFE_PP__3101  (.L_HI(net3101));
 sg13g2_tiehi \cpu.icache.r_data[7][23]$_DFFE_PP__3102  (.L_HI(net3102));
 sg13g2_tiehi \cpu.icache.r_data[7][24]$_DFFE_PP__3103  (.L_HI(net3103));
 sg13g2_tiehi \cpu.icache.r_data[7][25]$_DFFE_PP__3104  (.L_HI(net3104));
 sg13g2_tiehi \cpu.icache.r_data[7][26]$_DFFE_PP__3105  (.L_HI(net3105));
 sg13g2_tiehi \cpu.icache.r_data[7][27]$_DFFE_PP__3106  (.L_HI(net3106));
 sg13g2_tiehi \cpu.icache.r_data[7][28]$_DFFE_PP__3107  (.L_HI(net3107));
 sg13g2_tiehi \cpu.icache.r_data[7][29]$_DFFE_PP__3108  (.L_HI(net3108));
 sg13g2_tiehi \cpu.icache.r_data[7][2]$_DFFE_PP__3109  (.L_HI(net3109));
 sg13g2_tiehi \cpu.icache.r_data[7][30]$_DFFE_PP__3110  (.L_HI(net3110));
 sg13g2_tiehi \cpu.icache.r_data[7][31]$_DFFE_PP__3111  (.L_HI(net3111));
 sg13g2_tiehi \cpu.icache.r_data[7][3]$_DFFE_PP__3112  (.L_HI(net3112));
 sg13g2_tiehi \cpu.icache.r_data[7][4]$_DFFE_PP__3113  (.L_HI(net3113));
 sg13g2_tiehi \cpu.icache.r_data[7][5]$_DFFE_PP__3114  (.L_HI(net3114));
 sg13g2_tiehi \cpu.icache.r_data[7][6]$_DFFE_PP__3115  (.L_HI(net3115));
 sg13g2_tiehi \cpu.icache.r_data[7][7]$_DFFE_PP__3116  (.L_HI(net3116));
 sg13g2_tiehi \cpu.icache.r_data[7][8]$_DFFE_PP__3117  (.L_HI(net3117));
 sg13g2_tiehi \cpu.icache.r_data[7][9]$_DFFE_PP__3118  (.L_HI(net3118));
 sg13g2_tiehi \cpu.icache.r_offset[0]$_SDFF_PN0__3119  (.L_HI(net3119));
 sg13g2_tiehi \cpu.icache.r_offset[1]$_SDFF_PN0__3120  (.L_HI(net3120));
 sg13g2_tiehi \cpu.icache.r_offset[2]$_SDFF_PN0__3121  (.L_HI(net3121));
 sg13g2_tiehi \cpu.icache.r_tag[0][0]$_DFFE_PP__3122  (.L_HI(net3122));
 sg13g2_tiehi \cpu.icache.r_tag[0][10]$_DFFE_PP__3123  (.L_HI(net3123));
 sg13g2_tiehi \cpu.icache.r_tag[0][11]$_DFFE_PP__3124  (.L_HI(net3124));
 sg13g2_tiehi \cpu.icache.r_tag[0][12]$_DFFE_PP__3125  (.L_HI(net3125));
 sg13g2_tiehi \cpu.icache.r_tag[0][13]$_DFFE_PP__3126  (.L_HI(net3126));
 sg13g2_tiehi \cpu.icache.r_tag[0][14]$_DFFE_PP__3127  (.L_HI(net3127));
 sg13g2_tiehi \cpu.icache.r_tag[0][15]$_DFFE_PP__3128  (.L_HI(net3128));
 sg13g2_tiehi \cpu.icache.r_tag[0][16]$_DFFE_PP__3129  (.L_HI(net3129));
 sg13g2_tiehi \cpu.icache.r_tag[0][17]$_DFFE_PP__3130  (.L_HI(net3130));
 sg13g2_tiehi \cpu.icache.r_tag[0][18]$_DFFE_PP__3131  (.L_HI(net3131));
 sg13g2_tiehi \cpu.icache.r_tag[0][1]$_DFFE_PP__3132  (.L_HI(net3132));
 sg13g2_tiehi \cpu.icache.r_tag[0][2]$_DFFE_PP__3133  (.L_HI(net3133));
 sg13g2_tiehi \cpu.icache.r_tag[0][3]$_DFFE_PP__3134  (.L_HI(net3134));
 sg13g2_tiehi \cpu.icache.r_tag[0][4]$_DFFE_PP__3135  (.L_HI(net3135));
 sg13g2_tiehi \cpu.icache.r_tag[0][5]$_DFFE_PP__3136  (.L_HI(net3136));
 sg13g2_tiehi \cpu.icache.r_tag[0][6]$_DFFE_PP__3137  (.L_HI(net3137));
 sg13g2_tiehi \cpu.icache.r_tag[0][7]$_DFFE_PP__3138  (.L_HI(net3138));
 sg13g2_tiehi \cpu.icache.r_tag[0][8]$_DFFE_PP__3139  (.L_HI(net3139));
 sg13g2_tiehi \cpu.icache.r_tag[0][9]$_DFFE_PP__3140  (.L_HI(net3140));
 sg13g2_tiehi \cpu.icache.r_tag[1][0]$_DFFE_PP__3141  (.L_HI(net3141));
 sg13g2_tiehi \cpu.icache.r_tag[1][10]$_DFFE_PP__3142  (.L_HI(net3142));
 sg13g2_tiehi \cpu.icache.r_tag[1][11]$_DFFE_PP__3143  (.L_HI(net3143));
 sg13g2_tiehi \cpu.icache.r_tag[1][12]$_DFFE_PP__3144  (.L_HI(net3144));
 sg13g2_tiehi \cpu.icache.r_tag[1][13]$_DFFE_PP__3145  (.L_HI(net3145));
 sg13g2_tiehi \cpu.icache.r_tag[1][14]$_DFFE_PP__3146  (.L_HI(net3146));
 sg13g2_tiehi \cpu.icache.r_tag[1][15]$_DFFE_PP__3147  (.L_HI(net3147));
 sg13g2_tiehi \cpu.icache.r_tag[1][16]$_DFFE_PP__3148  (.L_HI(net3148));
 sg13g2_tiehi \cpu.icache.r_tag[1][17]$_DFFE_PP__3149  (.L_HI(net3149));
 sg13g2_tiehi \cpu.icache.r_tag[1][18]$_DFFE_PP__3150  (.L_HI(net3150));
 sg13g2_tiehi \cpu.icache.r_tag[1][1]$_DFFE_PP__3151  (.L_HI(net3151));
 sg13g2_tiehi \cpu.icache.r_tag[1][2]$_DFFE_PP__3152  (.L_HI(net3152));
 sg13g2_tiehi \cpu.icache.r_tag[1][3]$_DFFE_PP__3153  (.L_HI(net3153));
 sg13g2_tiehi \cpu.icache.r_tag[1][4]$_DFFE_PP__3154  (.L_HI(net3154));
 sg13g2_tiehi \cpu.icache.r_tag[1][5]$_DFFE_PP__3155  (.L_HI(net3155));
 sg13g2_tiehi \cpu.icache.r_tag[1][6]$_DFFE_PP__3156  (.L_HI(net3156));
 sg13g2_tiehi \cpu.icache.r_tag[1][7]$_DFFE_PP__3157  (.L_HI(net3157));
 sg13g2_tiehi \cpu.icache.r_tag[1][8]$_DFFE_PP__3158  (.L_HI(net3158));
 sg13g2_tiehi \cpu.icache.r_tag[1][9]$_DFFE_PP__3159  (.L_HI(net3159));
 sg13g2_tiehi \cpu.icache.r_tag[2][0]$_DFFE_PP__3160  (.L_HI(net3160));
 sg13g2_tiehi \cpu.icache.r_tag[2][10]$_DFFE_PP__3161  (.L_HI(net3161));
 sg13g2_tiehi \cpu.icache.r_tag[2][11]$_DFFE_PP__3162  (.L_HI(net3162));
 sg13g2_tiehi \cpu.icache.r_tag[2][12]$_DFFE_PP__3163  (.L_HI(net3163));
 sg13g2_tiehi \cpu.icache.r_tag[2][13]$_DFFE_PP__3164  (.L_HI(net3164));
 sg13g2_tiehi \cpu.icache.r_tag[2][14]$_DFFE_PP__3165  (.L_HI(net3165));
 sg13g2_tiehi \cpu.icache.r_tag[2][15]$_DFFE_PP__3166  (.L_HI(net3166));
 sg13g2_tiehi \cpu.icache.r_tag[2][16]$_DFFE_PP__3167  (.L_HI(net3167));
 sg13g2_tiehi \cpu.icache.r_tag[2][17]$_DFFE_PP__3168  (.L_HI(net3168));
 sg13g2_tiehi \cpu.icache.r_tag[2][18]$_DFFE_PP__3169  (.L_HI(net3169));
 sg13g2_tiehi \cpu.icache.r_tag[2][1]$_DFFE_PP__3170  (.L_HI(net3170));
 sg13g2_tiehi \cpu.icache.r_tag[2][2]$_DFFE_PP__3171  (.L_HI(net3171));
 sg13g2_tiehi \cpu.icache.r_tag[2][3]$_DFFE_PP__3172  (.L_HI(net3172));
 sg13g2_tiehi \cpu.icache.r_tag[2][4]$_DFFE_PP__3173  (.L_HI(net3173));
 sg13g2_tiehi \cpu.icache.r_tag[2][5]$_DFFE_PP__3174  (.L_HI(net3174));
 sg13g2_tiehi \cpu.icache.r_tag[2][6]$_DFFE_PP__3175  (.L_HI(net3175));
 sg13g2_tiehi \cpu.icache.r_tag[2][7]$_DFFE_PP__3176  (.L_HI(net3176));
 sg13g2_tiehi \cpu.icache.r_tag[2][8]$_DFFE_PP__3177  (.L_HI(net3177));
 sg13g2_tiehi \cpu.icache.r_tag[2][9]$_DFFE_PP__3178  (.L_HI(net3178));
 sg13g2_tiehi \cpu.icache.r_tag[3][0]$_DFFE_PP__3179  (.L_HI(net3179));
 sg13g2_tiehi \cpu.icache.r_tag[3][10]$_DFFE_PP__3180  (.L_HI(net3180));
 sg13g2_tiehi \cpu.icache.r_tag[3][11]$_DFFE_PP__3181  (.L_HI(net3181));
 sg13g2_tiehi \cpu.icache.r_tag[3][12]$_DFFE_PP__3182  (.L_HI(net3182));
 sg13g2_tiehi \cpu.icache.r_tag[3][13]$_DFFE_PP__3183  (.L_HI(net3183));
 sg13g2_tiehi \cpu.icache.r_tag[3][14]$_DFFE_PP__3184  (.L_HI(net3184));
 sg13g2_tiehi \cpu.icache.r_tag[3][15]$_DFFE_PP__3185  (.L_HI(net3185));
 sg13g2_tiehi \cpu.icache.r_tag[3][16]$_DFFE_PP__3186  (.L_HI(net3186));
 sg13g2_tiehi \cpu.icache.r_tag[3][17]$_DFFE_PP__3187  (.L_HI(net3187));
 sg13g2_tiehi \cpu.icache.r_tag[3][18]$_DFFE_PP__3188  (.L_HI(net3188));
 sg13g2_tiehi \cpu.icache.r_tag[3][1]$_DFFE_PP__3189  (.L_HI(net3189));
 sg13g2_tiehi \cpu.icache.r_tag[3][2]$_DFFE_PP__3190  (.L_HI(net3190));
 sg13g2_tiehi \cpu.icache.r_tag[3][3]$_DFFE_PP__3191  (.L_HI(net3191));
 sg13g2_tiehi \cpu.icache.r_tag[3][4]$_DFFE_PP__3192  (.L_HI(net3192));
 sg13g2_tiehi \cpu.icache.r_tag[3][5]$_DFFE_PP__3193  (.L_HI(net3193));
 sg13g2_tiehi \cpu.icache.r_tag[3][6]$_DFFE_PP__3194  (.L_HI(net3194));
 sg13g2_tiehi \cpu.icache.r_tag[3][7]$_DFFE_PP__3195  (.L_HI(net3195));
 sg13g2_tiehi \cpu.icache.r_tag[3][8]$_DFFE_PP__3196  (.L_HI(net3196));
 sg13g2_tiehi \cpu.icache.r_tag[3][9]$_DFFE_PP__3197  (.L_HI(net3197));
 sg13g2_tiehi \cpu.icache.r_tag[4][0]$_DFFE_PP__3198  (.L_HI(net3198));
 sg13g2_tiehi \cpu.icache.r_tag[4][10]$_DFFE_PP__3199  (.L_HI(net3199));
 sg13g2_tiehi \cpu.icache.r_tag[4][11]$_DFFE_PP__3200  (.L_HI(net3200));
 sg13g2_tiehi \cpu.icache.r_tag[4][12]$_DFFE_PP__3201  (.L_HI(net3201));
 sg13g2_tiehi \cpu.icache.r_tag[4][13]$_DFFE_PP__3202  (.L_HI(net3202));
 sg13g2_tiehi \cpu.icache.r_tag[4][14]$_DFFE_PP__3203  (.L_HI(net3203));
 sg13g2_tiehi \cpu.icache.r_tag[4][15]$_DFFE_PP__3204  (.L_HI(net3204));
 sg13g2_tiehi \cpu.icache.r_tag[4][16]$_DFFE_PP__3205  (.L_HI(net3205));
 sg13g2_tiehi \cpu.icache.r_tag[4][17]$_DFFE_PP__3206  (.L_HI(net3206));
 sg13g2_tiehi \cpu.icache.r_tag[4][18]$_DFFE_PP__3207  (.L_HI(net3207));
 sg13g2_tiehi \cpu.icache.r_tag[4][1]$_DFFE_PP__3208  (.L_HI(net3208));
 sg13g2_tiehi \cpu.icache.r_tag[4][2]$_DFFE_PP__3209  (.L_HI(net3209));
 sg13g2_tiehi \cpu.icache.r_tag[4][3]$_DFFE_PP__3210  (.L_HI(net3210));
 sg13g2_tiehi \cpu.icache.r_tag[4][4]$_DFFE_PP__3211  (.L_HI(net3211));
 sg13g2_tiehi \cpu.icache.r_tag[4][5]$_DFFE_PP__3212  (.L_HI(net3212));
 sg13g2_tiehi \cpu.icache.r_tag[4][6]$_DFFE_PP__3213  (.L_HI(net3213));
 sg13g2_tiehi \cpu.icache.r_tag[4][7]$_DFFE_PP__3214  (.L_HI(net3214));
 sg13g2_tiehi \cpu.icache.r_tag[4][8]$_DFFE_PP__3215  (.L_HI(net3215));
 sg13g2_tiehi \cpu.icache.r_tag[4][9]$_DFFE_PP__3216  (.L_HI(net3216));
 sg13g2_tiehi \cpu.icache.r_tag[5][0]$_DFFE_PP__3217  (.L_HI(net3217));
 sg13g2_tiehi \cpu.icache.r_tag[5][10]$_DFFE_PP__3218  (.L_HI(net3218));
 sg13g2_tiehi \cpu.icache.r_tag[5][11]$_DFFE_PP__3219  (.L_HI(net3219));
 sg13g2_tiehi \cpu.icache.r_tag[5][12]$_DFFE_PP__3220  (.L_HI(net3220));
 sg13g2_tiehi \cpu.icache.r_tag[5][13]$_DFFE_PP__3221  (.L_HI(net3221));
 sg13g2_tiehi \cpu.icache.r_tag[5][14]$_DFFE_PP__3222  (.L_HI(net3222));
 sg13g2_tiehi \cpu.icache.r_tag[5][15]$_DFFE_PP__3223  (.L_HI(net3223));
 sg13g2_tiehi \cpu.icache.r_tag[5][16]$_DFFE_PP__3224  (.L_HI(net3224));
 sg13g2_tiehi \cpu.icache.r_tag[5][17]$_DFFE_PP__3225  (.L_HI(net3225));
 sg13g2_tiehi \cpu.icache.r_tag[5][18]$_DFFE_PP__3226  (.L_HI(net3226));
 sg13g2_tiehi \cpu.icache.r_tag[5][1]$_DFFE_PP__3227  (.L_HI(net3227));
 sg13g2_tiehi \cpu.icache.r_tag[5][2]$_DFFE_PP__3228  (.L_HI(net3228));
 sg13g2_tiehi \cpu.icache.r_tag[5][3]$_DFFE_PP__3229  (.L_HI(net3229));
 sg13g2_tiehi \cpu.icache.r_tag[5][4]$_DFFE_PP__3230  (.L_HI(net3230));
 sg13g2_tiehi \cpu.icache.r_tag[5][5]$_DFFE_PP__3231  (.L_HI(net3231));
 sg13g2_tiehi \cpu.icache.r_tag[5][6]$_DFFE_PP__3232  (.L_HI(net3232));
 sg13g2_tiehi \cpu.icache.r_tag[5][7]$_DFFE_PP__3233  (.L_HI(net3233));
 sg13g2_tiehi \cpu.icache.r_tag[5][8]$_DFFE_PP__3234  (.L_HI(net3234));
 sg13g2_tiehi \cpu.icache.r_tag[5][9]$_DFFE_PP__3235  (.L_HI(net3235));
 sg13g2_tiehi \cpu.icache.r_tag[6][0]$_DFFE_PP__3236  (.L_HI(net3236));
 sg13g2_tiehi \cpu.icache.r_tag[6][10]$_DFFE_PP__3237  (.L_HI(net3237));
 sg13g2_tiehi \cpu.icache.r_tag[6][11]$_DFFE_PP__3238  (.L_HI(net3238));
 sg13g2_tiehi \cpu.icache.r_tag[6][12]$_DFFE_PP__3239  (.L_HI(net3239));
 sg13g2_tiehi \cpu.icache.r_tag[6][13]$_DFFE_PP__3240  (.L_HI(net3240));
 sg13g2_tiehi \cpu.icache.r_tag[6][14]$_DFFE_PP__3241  (.L_HI(net3241));
 sg13g2_tiehi \cpu.icache.r_tag[6][15]$_DFFE_PP__3242  (.L_HI(net3242));
 sg13g2_tiehi \cpu.icache.r_tag[6][16]$_DFFE_PP__3243  (.L_HI(net3243));
 sg13g2_tiehi \cpu.icache.r_tag[6][17]$_DFFE_PP__3244  (.L_HI(net3244));
 sg13g2_tiehi \cpu.icache.r_tag[6][18]$_DFFE_PP__3245  (.L_HI(net3245));
 sg13g2_tiehi \cpu.icache.r_tag[6][1]$_DFFE_PP__3246  (.L_HI(net3246));
 sg13g2_tiehi \cpu.icache.r_tag[6][2]$_DFFE_PP__3247  (.L_HI(net3247));
 sg13g2_tiehi \cpu.icache.r_tag[6][3]$_DFFE_PP__3248  (.L_HI(net3248));
 sg13g2_tiehi \cpu.icache.r_tag[6][4]$_DFFE_PP__3249  (.L_HI(net3249));
 sg13g2_tiehi \cpu.icache.r_tag[6][5]$_DFFE_PP__3250  (.L_HI(net3250));
 sg13g2_tiehi \cpu.icache.r_tag[6][6]$_DFFE_PP__3251  (.L_HI(net3251));
 sg13g2_tiehi \cpu.icache.r_tag[6][7]$_DFFE_PP__3252  (.L_HI(net3252));
 sg13g2_tiehi \cpu.icache.r_tag[6][8]$_DFFE_PP__3253  (.L_HI(net3253));
 sg13g2_tiehi \cpu.icache.r_tag[6][9]$_DFFE_PP__3254  (.L_HI(net3254));
 sg13g2_tiehi \cpu.icache.r_tag[7][0]$_DFFE_PP__3255  (.L_HI(net3255));
 sg13g2_tiehi \cpu.icache.r_tag[7][10]$_DFFE_PP__3256  (.L_HI(net3256));
 sg13g2_tiehi \cpu.icache.r_tag[7][11]$_DFFE_PP__3257  (.L_HI(net3257));
 sg13g2_tiehi \cpu.icache.r_tag[7][12]$_DFFE_PP__3258  (.L_HI(net3258));
 sg13g2_tiehi \cpu.icache.r_tag[7][13]$_DFFE_PP__3259  (.L_HI(net3259));
 sg13g2_tiehi \cpu.icache.r_tag[7][14]$_DFFE_PP__3260  (.L_HI(net3260));
 sg13g2_tiehi \cpu.icache.r_tag[7][15]$_DFFE_PP__3261  (.L_HI(net3261));
 sg13g2_tiehi \cpu.icache.r_tag[7][16]$_DFFE_PP__3262  (.L_HI(net3262));
 sg13g2_tiehi \cpu.icache.r_tag[7][17]$_DFFE_PP__3263  (.L_HI(net3263));
 sg13g2_tiehi \cpu.icache.r_tag[7][18]$_DFFE_PP__3264  (.L_HI(net3264));
 sg13g2_tiehi \cpu.icache.r_tag[7][1]$_DFFE_PP__3265  (.L_HI(net3265));
 sg13g2_tiehi \cpu.icache.r_tag[7][2]$_DFFE_PP__3266  (.L_HI(net3266));
 sg13g2_tiehi \cpu.icache.r_tag[7][3]$_DFFE_PP__3267  (.L_HI(net3267));
 sg13g2_tiehi \cpu.icache.r_tag[7][4]$_DFFE_PP__3268  (.L_HI(net3268));
 sg13g2_tiehi \cpu.icache.r_tag[7][5]$_DFFE_PP__3269  (.L_HI(net3269));
 sg13g2_tiehi \cpu.icache.r_tag[7][6]$_DFFE_PP__3270  (.L_HI(net3270));
 sg13g2_tiehi \cpu.icache.r_tag[7][7]$_DFFE_PP__3271  (.L_HI(net3271));
 sg13g2_tiehi \cpu.icache.r_tag[7][8]$_DFFE_PP__3272  (.L_HI(net3272));
 sg13g2_tiehi \cpu.icache.r_tag[7][9]$_DFFE_PP__3273  (.L_HI(net3273));
 sg13g2_tiehi \cpu.icache.r_valid[0]$_SDFFE_PP0P__3274  (.L_HI(net3274));
 sg13g2_tiehi \cpu.icache.r_valid[1]$_SDFFE_PP0P__3275  (.L_HI(net3275));
 sg13g2_tiehi \cpu.icache.r_valid[2]$_SDFFE_PP0P__3276  (.L_HI(net3276));
 sg13g2_tiehi \cpu.icache.r_valid[3]$_SDFFE_PP0P__3277  (.L_HI(net3277));
 sg13g2_tiehi \cpu.icache.r_valid[4]$_SDFFE_PP0P__3278  (.L_HI(net3278));
 sg13g2_tiehi \cpu.icache.r_valid[5]$_SDFFE_PP0P__3279  (.L_HI(net3279));
 sg13g2_tiehi \cpu.icache.r_valid[6]$_SDFFE_PP0P__3280  (.L_HI(net3280));
 sg13g2_tiehi \cpu.icache.r_valid[7]$_SDFFE_PP0P__3281  (.L_HI(net3281));
 sg13g2_tiehi \cpu.intr.r_clock$_SDFFE_PN0P__3282  (.L_HI(net3282));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[0]$_DFFE_PP__3283  (.L_HI(net3283));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[10]$_DFFE_PP__3284  (.L_HI(net3284));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[11]$_DFFE_PP__3285  (.L_HI(net3285));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[12]$_DFFE_PP__3286  (.L_HI(net3286));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[13]$_DFFE_PP__3287  (.L_HI(net3287));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[14]$_DFFE_PP__3288  (.L_HI(net3288));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[15]$_DFFE_PP__3289  (.L_HI(net3289));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[16]$_DFFE_PP__3290  (.L_HI(net3290));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[17]$_DFFE_PP__3291  (.L_HI(net3291));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[18]$_DFFE_PP__3292  (.L_HI(net3292));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[19]$_DFFE_PP__3293  (.L_HI(net3293));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[1]$_DFFE_PP__3294  (.L_HI(net3294));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[20]$_DFFE_PP__3295  (.L_HI(net3295));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[21]$_DFFE_PP__3296  (.L_HI(net3296));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[22]$_DFFE_PP__3297  (.L_HI(net3297));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[23]$_DFFE_PP__3298  (.L_HI(net3298));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[24]$_DFFE_PP__3299  (.L_HI(net3299));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[25]$_DFFE_PP__3300  (.L_HI(net3300));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[26]$_DFFE_PP__3301  (.L_HI(net3301));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[27]$_DFFE_PP__3302  (.L_HI(net3302));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[28]$_DFFE_PP__3303  (.L_HI(net3303));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[29]$_DFFE_PP__3304  (.L_HI(net3304));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[2]$_DFFE_PP__3305  (.L_HI(net3305));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[30]$_DFFE_PP__3306  (.L_HI(net3306));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[31]$_DFFE_PP__3307  (.L_HI(net3307));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[3]$_DFFE_PP__3308  (.L_HI(net3308));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[4]$_DFFE_PP__3309  (.L_HI(net3309));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[5]$_DFFE_PP__3310  (.L_HI(net3310));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[6]$_DFFE_PP__3311  (.L_HI(net3311));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[7]$_DFFE_PP__3312  (.L_HI(net3312));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[8]$_DFFE_PP__3313  (.L_HI(net3313));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[9]$_DFFE_PP__3314  (.L_HI(net3314));
 sg13g2_tiehi \cpu.intr.r_clock_count[0]$_DFF_P__3315  (.L_HI(net3315));
 sg13g2_tiehi \cpu.intr.r_clock_count[10]$_DFF_P__3316  (.L_HI(net3316));
 sg13g2_tiehi \cpu.intr.r_clock_count[11]$_DFF_P__3317  (.L_HI(net3317));
 sg13g2_tiehi \cpu.intr.r_clock_count[12]$_DFF_P__3318  (.L_HI(net3318));
 sg13g2_tiehi \cpu.intr.r_clock_count[13]$_DFF_P__3319  (.L_HI(net3319));
 sg13g2_tiehi \cpu.intr.r_clock_count[14]$_DFF_P__3320  (.L_HI(net3320));
 sg13g2_tiehi \cpu.intr.r_clock_count[15]$_DFF_P__3321  (.L_HI(net3321));
 sg13g2_tiehi \cpu.intr.r_clock_count[16]$_DFFE_PN__3322  (.L_HI(net3322));
 sg13g2_tiehi \cpu.intr.r_clock_count[17]$_DFFE_PN__3323  (.L_HI(net3323));
 sg13g2_tiehi \cpu.intr.r_clock_count[18]$_DFFE_PN__3324  (.L_HI(net3324));
 sg13g2_tiehi \cpu.intr.r_clock_count[19]$_DFFE_PN__3325  (.L_HI(net3325));
 sg13g2_tiehi \cpu.intr.r_clock_count[1]$_DFF_P__3326  (.L_HI(net3326));
 sg13g2_tiehi \cpu.intr.r_clock_count[20]$_DFFE_PN__3327  (.L_HI(net3327));
 sg13g2_tiehi \cpu.intr.r_clock_count[21]$_DFFE_PN__3328  (.L_HI(net3328));
 sg13g2_tiehi \cpu.intr.r_clock_count[22]$_DFFE_PN__3329  (.L_HI(net3329));
 sg13g2_tiehi \cpu.intr.r_clock_count[23]$_DFFE_PN__3330  (.L_HI(net3330));
 sg13g2_tiehi \cpu.intr.r_clock_count[24]$_DFFE_PN__3331  (.L_HI(net3331));
 sg13g2_tiehi \cpu.intr.r_clock_count[25]$_DFFE_PN__3332  (.L_HI(net3332));
 sg13g2_tiehi \cpu.intr.r_clock_count[26]$_DFFE_PN__3333  (.L_HI(net3333));
 sg13g2_tiehi \cpu.intr.r_clock_count[27]$_DFFE_PN__3334  (.L_HI(net3334));
 sg13g2_tiehi \cpu.intr.r_clock_count[28]$_DFFE_PN__3335  (.L_HI(net3335));
 sg13g2_tiehi \cpu.intr.r_clock_count[29]$_DFFE_PN__3336  (.L_HI(net3336));
 sg13g2_tiehi \cpu.intr.r_clock_count[2]$_DFF_P__3337  (.L_HI(net3337));
 sg13g2_tiehi \cpu.intr.r_clock_count[30]$_DFFE_PN__3338  (.L_HI(net3338));
 sg13g2_tiehi \cpu.intr.r_clock_count[31]$_DFFE_PN__3339  (.L_HI(net3339));
 sg13g2_tiehi \cpu.intr.r_clock_count[3]$_DFF_P__3340  (.L_HI(net3340));
 sg13g2_tiehi \cpu.intr.r_clock_count[4]$_DFF_P__3341  (.L_HI(net3341));
 sg13g2_tiehi \cpu.intr.r_clock_count[5]$_DFF_P__3342  (.L_HI(net3342));
 sg13g2_tiehi \cpu.intr.r_clock_count[6]$_DFF_P__3343  (.L_HI(net3343));
 sg13g2_tiehi \cpu.intr.r_clock_count[7]$_DFF_P__3344  (.L_HI(net3344));
 sg13g2_tiehi \cpu.intr.r_clock_count[8]$_DFF_P__3345  (.L_HI(net3345));
 sg13g2_tiehi \cpu.intr.r_clock_count[9]$_DFF_P__3346  (.L_HI(net3346));
 sg13g2_tiehi \cpu.intr.r_enable[0]$_SDFFE_PN0P__3347  (.L_HI(net3347));
 sg13g2_tiehi \cpu.intr.r_enable[1]$_SDFFE_PN0P__3348  (.L_HI(net3348));
 sg13g2_tiehi \cpu.intr.r_enable[2]$_SDFFE_PN0P__3349  (.L_HI(net3349));
 sg13g2_tiehi \cpu.intr.r_enable[3]$_SDFFE_PN0P__3350  (.L_HI(net3350));
 sg13g2_tiehi \cpu.intr.r_enable[4]$_SDFFE_PN0P__3351  (.L_HI(net3351));
 sg13g2_tiehi \cpu.intr.r_enable[5]$_SDFFE_PN0P__3352  (.L_HI(net3352));
 sg13g2_tiehi \cpu.intr.r_timer$_SDFFE_PN0P__3353  (.L_HI(net3353));
 sg13g2_tiehi \cpu.intr.r_timer_count[0]$_DFF_P__3354  (.L_HI(net3354));
 sg13g2_tiehi \cpu.intr.r_timer_count[10]$_DFF_P__3355  (.L_HI(net3355));
 sg13g2_tiehi \cpu.intr.r_timer_count[11]$_DFF_P__3356  (.L_HI(net3356));
 sg13g2_tiehi \cpu.intr.r_timer_count[12]$_DFF_P__3357  (.L_HI(net3357));
 sg13g2_tiehi \cpu.intr.r_timer_count[13]$_DFF_P__3358  (.L_HI(net3358));
 sg13g2_tiehi \cpu.intr.r_timer_count[14]$_DFF_P__3359  (.L_HI(net3359));
 sg13g2_tiehi \cpu.intr.r_timer_count[15]$_DFF_P__3360  (.L_HI(net3360));
 sg13g2_tiehi \cpu.intr.r_timer_count[16]$_DFF_P__3361  (.L_HI(net3361));
 sg13g2_tiehi \cpu.intr.r_timer_count[17]$_DFF_P__3362  (.L_HI(net3362));
 sg13g2_tiehi \cpu.intr.r_timer_count[18]$_DFF_P__3363  (.L_HI(net3363));
 sg13g2_tiehi \cpu.intr.r_timer_count[19]$_DFF_P__3364  (.L_HI(net3364));
 sg13g2_tiehi \cpu.intr.r_timer_count[1]$_DFF_P__3365  (.L_HI(net3365));
 sg13g2_tiehi \cpu.intr.r_timer_count[20]$_DFF_P__3366  (.L_HI(net3366));
 sg13g2_tiehi \cpu.intr.r_timer_count[21]$_DFF_P__3367  (.L_HI(net3367));
 sg13g2_tiehi \cpu.intr.r_timer_count[22]$_DFF_P__3368  (.L_HI(net3368));
 sg13g2_tiehi \cpu.intr.r_timer_count[23]$_DFF_P__3369  (.L_HI(net3369));
 sg13g2_tiehi \cpu.intr.r_timer_count[2]$_DFF_P__3370  (.L_HI(net3370));
 sg13g2_tiehi \cpu.intr.r_timer_count[3]$_DFF_P__3371  (.L_HI(net3371));
 sg13g2_tiehi \cpu.intr.r_timer_count[4]$_DFF_P__3372  (.L_HI(net3372));
 sg13g2_tiehi \cpu.intr.r_timer_count[5]$_DFF_P__3373  (.L_HI(net3373));
 sg13g2_tiehi \cpu.intr.r_timer_count[6]$_DFF_P__3374  (.L_HI(net3374));
 sg13g2_tiehi \cpu.intr.r_timer_count[7]$_DFF_P__3375  (.L_HI(net3375));
 sg13g2_tiehi \cpu.intr.r_timer_count[8]$_DFF_P__3376  (.L_HI(net3376));
 sg13g2_tiehi \cpu.intr.r_timer_count[9]$_DFF_P__3377  (.L_HI(net3377));
 sg13g2_tiehi \cpu.intr.r_timer_reload[0]$_DFFE_PP__3378  (.L_HI(net3378));
 sg13g2_tiehi \cpu.intr.r_timer_reload[10]$_DFFE_PP__3379  (.L_HI(net3379));
 sg13g2_tiehi \cpu.intr.r_timer_reload[11]$_DFFE_PP__3380  (.L_HI(net3380));
 sg13g2_tiehi \cpu.intr.r_timer_reload[12]$_DFFE_PP__3381  (.L_HI(net3381));
 sg13g2_tiehi \cpu.intr.r_timer_reload[13]$_DFFE_PP__3382  (.L_HI(net3382));
 sg13g2_tiehi \cpu.intr.r_timer_reload[14]$_DFFE_PP__3383  (.L_HI(net3383));
 sg13g2_tiehi \cpu.intr.r_timer_reload[15]$_DFFE_PP__3384  (.L_HI(net3384));
 sg13g2_tiehi \cpu.intr.r_timer_reload[16]$_DFFE_PP__3385  (.L_HI(net3385));
 sg13g2_tiehi \cpu.intr.r_timer_reload[17]$_DFFE_PP__3386  (.L_HI(net3386));
 sg13g2_tiehi \cpu.intr.r_timer_reload[18]$_DFFE_PP__3387  (.L_HI(net3387));
 sg13g2_tiehi \cpu.intr.r_timer_reload[19]$_DFFE_PP__3388  (.L_HI(net3388));
 sg13g2_tiehi \cpu.intr.r_timer_reload[1]$_DFFE_PP__3389  (.L_HI(net3389));
 sg13g2_tiehi \cpu.intr.r_timer_reload[20]$_DFFE_PP__3390  (.L_HI(net3390));
 sg13g2_tiehi \cpu.intr.r_timer_reload[21]$_DFFE_PP__3391  (.L_HI(net3391));
 sg13g2_tiehi \cpu.intr.r_timer_reload[22]$_DFFE_PP__3392  (.L_HI(net3392));
 sg13g2_tiehi \cpu.intr.r_timer_reload[23]$_DFFE_PP__3393  (.L_HI(net3393));
 sg13g2_tiehi \cpu.intr.r_timer_reload[2]$_DFFE_PP__3394  (.L_HI(net3394));
 sg13g2_tiehi \cpu.intr.r_timer_reload[3]$_DFFE_PP__3395  (.L_HI(net3395));
 sg13g2_tiehi \cpu.intr.r_timer_reload[4]$_DFFE_PP__3396  (.L_HI(net3396));
 sg13g2_tiehi \cpu.intr.r_timer_reload[5]$_DFFE_PP__3397  (.L_HI(net3397));
 sg13g2_tiehi \cpu.intr.r_timer_reload[6]$_DFFE_PP__3398  (.L_HI(net3398));
 sg13g2_tiehi \cpu.intr.r_timer_reload[7]$_DFFE_PP__3399  (.L_HI(net3399));
 sg13g2_tiehi \cpu.intr.r_timer_reload[8]$_DFFE_PP__3400  (.L_HI(net3400));
 sg13g2_tiehi \cpu.intr.r_timer_reload[9]$_DFFE_PP__3401  (.L_HI(net3401));
 sg13g2_tiehi \cpu.qspi.r_count[0]$_DFFE_PP__3402  (.L_HI(net3402));
 sg13g2_tiehi \cpu.qspi.r_count[1]$_DFFE_PP__3403  (.L_HI(net3403));
 sg13g2_tiehi \cpu.qspi.r_count[2]$_DFFE_PP__3404  (.L_HI(net3404));
 sg13g2_tiehi \cpu.qspi.r_count[3]$_DFFE_PP__3405  (.L_HI(net3405));
 sg13g2_tiehi \cpu.qspi.r_count[4]$_DFFE_PP__3406  (.L_HI(net3406));
 sg13g2_tiehi \cpu.qspi.r_cs[0]$_SDFFE_PN1P__3407  (.L_HI(net3407));
 sg13g2_tiehi \cpu.qspi.r_cs[1]$_SDFFE_PN1P__3408  (.L_HI(net3408));
 sg13g2_tiehi \cpu.qspi.r_cs[2]$_SDFFE_PN1P__3409  (.L_HI(net3409));
 sg13g2_tiehi \cpu.qspi.r_ind$_SDFFE_PN0N__3410  (.L_HI(net3410));
 sg13g2_tiehi \cpu.qspi.r_mask[0]$_SDFFE_PN0P__3411  (.L_HI(net3411));
 sg13g2_tiehi \cpu.qspi.r_mask[1]$_SDFFE_PN1P__3412  (.L_HI(net3412));
 sg13g2_tiehi \cpu.qspi.r_mask[2]$_SDFFE_PN0P__3413  (.L_HI(net3413));
 sg13g2_tiehi \cpu.qspi.r_quad[0]$_SDFFE_PN1P__3414  (.L_HI(net3414));
 sg13g2_tiehi \cpu.qspi.r_quad[1]$_SDFFE_PN0P__3415  (.L_HI(net3415));
 sg13g2_tiehi \cpu.qspi.r_quad[2]$_SDFFE_PN1P__3416  (.L_HI(net3416));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P__3417  (.L_HI(net3417));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P__3418  (.L_HI(net3418));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P__3419  (.L_HI(net3419));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P__3420  (.L_HI(net3420));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P__3421  (.L_HI(net3421));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P__3422  (.L_HI(net3422));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P__3423  (.L_HI(net3423));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P__3424  (.L_HI(net3424));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P__3425  (.L_HI(net3425));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P__3426  (.L_HI(net3426));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P__3427  (.L_HI(net3427));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P__3428  (.L_HI(net3428));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P__3429  (.L_HI(net3429));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P__3430  (.L_HI(net3430));
 sg13g2_tiehi \cpu.qspi.r_rstrobe_d$_DFF_P__3431  (.L_HI(net3431));
 sg13g2_tiehi \cpu.qspi.r_state[0]$_DFF_P__3432  (.L_HI(net3432));
 sg13g2_tiehi \cpu.qspi.r_state[10]$_DFF_P__3433  (.L_HI(net3433));
 sg13g2_tiehi \cpu.qspi.r_state[11]$_DFF_P__3434  (.L_HI(net3434));
 sg13g2_tiehi \cpu.qspi.r_state[12]$_DFF_P__3435  (.L_HI(net3435));
 sg13g2_tiehi \cpu.qspi.r_state[13]$_DFF_P__3436  (.L_HI(net3436));
 sg13g2_tiehi \cpu.qspi.r_state[14]$_DFF_P__3437  (.L_HI(net3437));
 sg13g2_tiehi \cpu.qspi.r_state[15]$_DFF_P__3438  (.L_HI(net3438));
 sg13g2_tiehi \cpu.qspi.r_state[16]$_DFF_P__3439  (.L_HI(net3439));
 sg13g2_tiehi \cpu.qspi.r_state[17]$_DFF_P__3440  (.L_HI(net3440));
 sg13g2_tiehi \cpu.qspi.r_state[1]$_DFF_P__3441  (.L_HI(net3441));
 sg13g2_tiehi \cpu.qspi.r_state[2]$_DFF_P__3442  (.L_HI(net3442));
 sg13g2_tiehi \cpu.qspi.r_state[3]$_DFF_P__3443  (.L_HI(net3443));
 sg13g2_tiehi \cpu.qspi.r_state[4]$_DFF_P__3444  (.L_HI(net3444));
 sg13g2_tiehi \cpu.qspi.r_state[5]$_DFF_P__3445  (.L_HI(net3445));
 sg13g2_tiehi \cpu.qspi.r_state[6]$_DFF_P__3446  (.L_HI(net3446));
 sg13g2_tiehi \cpu.qspi.r_state[7]$_DFF_P__3447  (.L_HI(net3447));
 sg13g2_tiehi \cpu.qspi.r_state[8]$_DFF_P__3448  (.L_HI(net3448));
 sg13g2_tiehi \cpu.qspi.r_state[9]$_DFF_P__3449  (.L_HI(net3449));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P__3450  (.L_HI(net3450));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P__3451  (.L_HI(net3451));
 sg13g2_tiehi \cpu.qspi.r_uio_out[0]$_DFFE_PP__3452  (.L_HI(net3452));
 sg13g2_tiehi \cpu.qspi.r_uio_out[1]$_DFFE_PP__3453  (.L_HI(net3453));
 sg13g2_tiehi \cpu.qspi.r_uio_out[2]$_DFFE_PP__3454  (.L_HI(net3454));
 sg13g2_tiehi \cpu.qspi.r_uio_out[3]$_DFFE_PP__3455  (.L_HI(net3455));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_d$_DFF_P__3456  (.L_HI(net3456));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_i$_DFF_P__3457  (.L_HI(net3457));
 sg13g2_tiehi \cpu.r_clk_invert$_DFFE_PN__3458  (.L_HI(net3458));
 sg13g2_tiehi \cpu.spi.r_bits[0]$_SDFFE_PN1P__3459  (.L_HI(net3459));
 sg13g2_tiehi \cpu.spi.r_bits[1]$_SDFFE_PN1P__3460  (.L_HI(net3460));
 sg13g2_tiehi \cpu.spi.r_bits[2]$_SDFFE_PN1P__3461  (.L_HI(net3461));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][0]$_SDFFE_PN0P__3462  (.L_HI(net3462));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][1]$_SDFFE_PN0P__3463  (.L_HI(net3463));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][2]$_SDFFE_PN0P__3464  (.L_HI(net3464));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][3]$_SDFFE_PN0P__3465  (.L_HI(net3465));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][4]$_SDFFE_PN0P__3466  (.L_HI(net3466));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][5]$_SDFFE_PN0P__3467  (.L_HI(net3467));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][6]$_SDFFE_PN0P__3468  (.L_HI(net3468));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][7]$_SDFFE_PN0P__3469  (.L_HI(net3469));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][0]$_SDFFE_PN0P__3470  (.L_HI(net3470));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][1]$_SDFFE_PN0P__3471  (.L_HI(net3471));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][2]$_SDFFE_PN0P__3472  (.L_HI(net3472));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][3]$_SDFFE_PN0P__3473  (.L_HI(net3473));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][4]$_SDFFE_PN0P__3474  (.L_HI(net3474));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][5]$_SDFFE_PN0P__3475  (.L_HI(net3475));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][6]$_SDFFE_PN0P__3476  (.L_HI(net3476));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][7]$_SDFFE_PN0P__3477  (.L_HI(net3477));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][0]$_SDFFE_PN0P__3478  (.L_HI(net3478));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][1]$_SDFFE_PN0P__3479  (.L_HI(net3479));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][2]$_SDFFE_PN0P__3480  (.L_HI(net3480));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][3]$_SDFFE_PN0P__3481  (.L_HI(net3481));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][4]$_SDFFE_PN0P__3482  (.L_HI(net3482));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][5]$_SDFFE_PN0P__3483  (.L_HI(net3483));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][6]$_SDFFE_PN0P__3484  (.L_HI(net3484));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][7]$_SDFFE_PN0P__3485  (.L_HI(net3485));
 sg13g2_tiehi \cpu.spi.r_count[0]$_SDFFE_PN0P__3486  (.L_HI(net3486));
 sg13g2_tiehi \cpu.spi.r_count[1]$_SDFFE_PN0P__3487  (.L_HI(net3487));
 sg13g2_tiehi \cpu.spi.r_count[2]$_SDFFE_PN0P__3488  (.L_HI(net3488));
 sg13g2_tiehi \cpu.spi.r_count[3]$_SDFFE_PN0P__3489  (.L_HI(net3489));
 sg13g2_tiehi \cpu.spi.r_count[4]$_SDFFE_PN0P__3490  (.L_HI(net3490));
 sg13g2_tiehi \cpu.spi.r_count[5]$_SDFFE_PN0P__3491  (.L_HI(net3491));
 sg13g2_tiehi \cpu.spi.r_count[6]$_SDFFE_PN0P__3492  (.L_HI(net3492));
 sg13g2_tiehi \cpu.spi.r_count[7]$_SDFFE_PN0P__3493  (.L_HI(net3493));
 sg13g2_tiehi \cpu.spi.r_cs[0]$_SDFFE_PN1P__3494  (.L_HI(net3494));
 sg13g2_tiehi \cpu.spi.r_cs[1]$_SDFFE_PN1P__3495  (.L_HI(net3495));
 sg13g2_tiehi \cpu.spi.r_cs[2]$_SDFFE_PN1P__3496  (.L_HI(net3496));
 sg13g2_tiehi \cpu.spi.r_in[0]$_DFFE_PP__3497  (.L_HI(net3497));
 sg13g2_tiehi \cpu.spi.r_in[1]$_DFFE_PP__3498  (.L_HI(net3498));
 sg13g2_tiehi \cpu.spi.r_in[2]$_DFFE_PP__3499  (.L_HI(net3499));
 sg13g2_tiehi \cpu.spi.r_in[3]$_DFFE_PP__3500  (.L_HI(net3500));
 sg13g2_tiehi \cpu.spi.r_in[4]$_DFFE_PP__3501  (.L_HI(net3501));
 sg13g2_tiehi \cpu.spi.r_in[5]$_DFFE_PP__3502  (.L_HI(net3502));
 sg13g2_tiehi \cpu.spi.r_in[6]$_DFFE_PP__3503  (.L_HI(net3503));
 sg13g2_tiehi \cpu.spi.r_in[7]$_DFFE_PP__3504  (.L_HI(net3504));
 sg13g2_tiehi \cpu.spi.r_interrupt$_SDFFE_PN0P__3505  (.L_HI(net3505));
 sg13g2_tiehi \cpu.spi.r_mode[0][0]$_SDFFE_PN0P__3506  (.L_HI(net3506));
 sg13g2_tiehi \cpu.spi.r_mode[0][1]$_SDFFE_PN0P__3507  (.L_HI(net3507));
 sg13g2_tiehi \cpu.spi.r_mode[1][0]$_SDFFE_PN0P__3508  (.L_HI(net3508));
 sg13g2_tiehi \cpu.spi.r_mode[1][1]$_SDFFE_PN0P__3509  (.L_HI(net3509));
 sg13g2_tiehi \cpu.spi.r_mode[2][0]$_SDFFE_PN0P__3510  (.L_HI(net3510));
 sg13g2_tiehi \cpu.spi.r_mode[2][1]$_SDFFE_PN0P__3511  (.L_HI(net3511));
 sg13g2_tiehi \cpu.spi.r_out[0]$_DFFE_PP__3512  (.L_HI(net3512));
 sg13g2_tiehi \cpu.spi.r_out[1]$_DFFE_PP__3513  (.L_HI(net3513));
 sg13g2_tiehi \cpu.spi.r_out[2]$_DFFE_PP__3514  (.L_HI(net3514));
 sg13g2_tiehi \cpu.spi.r_out[3]$_DFFE_PP__3515  (.L_HI(net3515));
 sg13g2_tiehi \cpu.spi.r_out[4]$_DFFE_PP__3516  (.L_HI(net3516));
 sg13g2_tiehi \cpu.spi.r_out[5]$_DFFE_PP__3517  (.L_HI(net3517));
 sg13g2_tiehi \cpu.spi.r_out[6]$_DFFE_PP__3518  (.L_HI(net3518));
 sg13g2_tiehi \cpu.spi.r_out[7]$_DFFE_PP__3519  (.L_HI(net3519));
 sg13g2_tiehi \cpu.spi.r_ready$_SDFFE_PN1P__3520  (.L_HI(net3520));
 sg13g2_tiehi \cpu.spi.r_searching$_SDFFE_PN0P__3521  (.L_HI(net3521));
 sg13g2_tiehi \cpu.spi.r_sel[0]$_DFFE_PP__3522  (.L_HI(net3522));
 sg13g2_tiehi \cpu.spi.r_sel[1]$_DFFE_PP__3523  (.L_HI(net3523));
 sg13g2_tiehi \cpu.spi.r_src[0]$_SDFFE_PN0P__3524  (.L_HI(net3524));
 sg13g2_tiehi \cpu.spi.r_src[1]$_SDFFE_PN0P__3525  (.L_HI(net3525));
 sg13g2_tiehi \cpu.spi.r_src[2]$_SDFFE_PN0P__3526  (.L_HI(net3526));
 sg13g2_tiehi \cpu.spi.r_state[0]$_DFF_P__3527  (.L_HI(net3527));
 sg13g2_tiehi \cpu.spi.r_state[1]$_DFF_P__3528  (.L_HI(net3528));
 sg13g2_tiehi \cpu.spi.r_state[2]$_DFF_P__3529  (.L_HI(net3529));
 sg13g2_tiehi \cpu.spi.r_state[3]$_DFF_P__3530  (.L_HI(net3530));
 sg13g2_tiehi \cpu.spi.r_state[4]$_DFF_P__3531  (.L_HI(net3531));
 sg13g2_tiehi \cpu.spi.r_state[5]$_DFF_P__3532  (.L_HI(net3532));
 sg13g2_tiehi \cpu.spi.r_state[6]$_DFF_P__3533  (.L_HI(net3533));
 sg13g2_tiehi \cpu.spi.r_timeout[0]$_DFFE_PP__3534  (.L_HI(net3534));
 sg13g2_tiehi \cpu.spi.r_timeout[1]$_DFFE_PP__3535  (.L_HI(net3535));
 sg13g2_tiehi \cpu.spi.r_timeout[2]$_DFFE_PP__3536  (.L_HI(net3536));
 sg13g2_tiehi \cpu.spi.r_timeout[3]$_DFFE_PP__3537  (.L_HI(net3537));
 sg13g2_tiehi \cpu.spi.r_timeout[4]$_DFFE_PP__3538  (.L_HI(net3538));
 sg13g2_tiehi \cpu.spi.r_timeout[5]$_DFFE_PP__3539  (.L_HI(net3539));
 sg13g2_tiehi \cpu.spi.r_timeout[6]$_DFFE_PP__3540  (.L_HI(net3540));
 sg13g2_tiehi \cpu.spi.r_timeout[7]$_DFFE_PP__3541  (.L_HI(net3541));
 sg13g2_tiehi \cpu.spi.r_timeout_count[0]$_DFFE_PP__3542  (.L_HI(net3542));
 sg13g2_tiehi \cpu.spi.r_timeout_count[1]$_DFFE_PP__3543  (.L_HI(net3543));
 sg13g2_tiehi \cpu.spi.r_timeout_count[2]$_DFFE_PP__3544  (.L_HI(net3544));
 sg13g2_tiehi \cpu.spi.r_timeout_count[3]$_DFFE_PP__3545  (.L_HI(net3545));
 sg13g2_tiehi \cpu.spi.r_timeout_count[4]$_DFFE_PP__3546  (.L_HI(net3546));
 sg13g2_tiehi \cpu.spi.r_timeout_count[5]$_DFFE_PP__3547  (.L_HI(net3547));
 sg13g2_tiehi \cpu.spi.r_timeout_count[6]$_DFFE_PP__3548  (.L_HI(net3548));
 sg13g2_tiehi \cpu.spi.r_timeout_count[7]$_DFFE_PP__3549  (.L_HI(net3549));
 sg13g2_tiehi \cpu.uart.r_div[0]$_DFF_P__3550  (.L_HI(net3550));
 sg13g2_tiehi \cpu.uart.r_div[10]$_DFF_P__3551  (.L_HI(net3551));
 sg13g2_tiehi \cpu.uart.r_div[11]$_DFF_P__3552  (.L_HI(net3552));
 sg13g2_tiehi \cpu.uart.r_div[1]$_DFF_P__3553  (.L_HI(net3553));
 sg13g2_tiehi \cpu.uart.r_div[2]$_DFF_P__3554  (.L_HI(net3554));
 sg13g2_tiehi \cpu.uart.r_div[3]$_DFF_P__3555  (.L_HI(net3555));
 sg13g2_tiehi \cpu.uart.r_div[4]$_DFF_P__3556  (.L_HI(net3556));
 sg13g2_tiehi \cpu.uart.r_div[5]$_DFF_P__3557  (.L_HI(net3557));
 sg13g2_tiehi \cpu.uart.r_div[6]$_DFF_P__3558  (.L_HI(net3558));
 sg13g2_tiehi \cpu.uart.r_div[7]$_DFF_P__3559  (.L_HI(net3559));
 sg13g2_tiehi \cpu.uart.r_div[8]$_DFF_P__3560  (.L_HI(net3560));
 sg13g2_tiehi \cpu.uart.r_div[9]$_DFF_P__3561  (.L_HI(net3561));
 sg13g2_tiehi \cpu.uart.r_div_value[0]$_SDFFE_PN1P__3562  (.L_HI(net3562));
 sg13g2_tiehi \cpu.uart.r_div_value[10]$_SDFFE_PN0P__3563  (.L_HI(net3563));
 sg13g2_tiehi \cpu.uart.r_div_value[11]$_SDFFE_PN0P__3564  (.L_HI(net3564));
 sg13g2_tiehi \cpu.uart.r_div_value[1]$_SDFFE_PN0P__3565  (.L_HI(net3565));
 sg13g2_tiehi \cpu.uart.r_div_value[2]$_SDFFE_PN0P__3566  (.L_HI(net3566));
 sg13g2_tiehi \cpu.uart.r_div_value[3]$_SDFFE_PN0P__3567  (.L_HI(net3567));
 sg13g2_tiehi \cpu.uart.r_div_value[4]$_SDFFE_PN0P__3568  (.L_HI(net3568));
 sg13g2_tiehi \cpu.uart.r_div_value[5]$_SDFFE_PN0P__3569  (.L_HI(net3569));
 sg13g2_tiehi \cpu.uart.r_div_value[6]$_SDFFE_PN0P__3570  (.L_HI(net3570));
 sg13g2_tiehi \cpu.uart.r_div_value[7]$_SDFFE_PN0P__3571  (.L_HI(net3571));
 sg13g2_tiehi \cpu.uart.r_div_value[8]$_SDFFE_PN0P__3572  (.L_HI(net3572));
 sg13g2_tiehi \cpu.uart.r_div_value[9]$_SDFFE_PN0P__3573  (.L_HI(net3573));
 sg13g2_tiehi \cpu.uart.r_ib[0]$_DFFE_PP__3574  (.L_HI(net3574));
 sg13g2_tiehi \cpu.uart.r_ib[1]$_DFFE_PP__3575  (.L_HI(net3575));
 sg13g2_tiehi \cpu.uart.r_ib[2]$_DFFE_PP__3576  (.L_HI(net3576));
 sg13g2_tiehi \cpu.uart.r_ib[3]$_DFFE_PP__3577  (.L_HI(net3577));
 sg13g2_tiehi \cpu.uart.r_ib[4]$_DFFE_PP__3578  (.L_HI(net3578));
 sg13g2_tiehi \cpu.uart.r_ib[5]$_DFFE_PP__3579  (.L_HI(net3579));
 sg13g2_tiehi \cpu.uart.r_ib[6]$_DFFE_PP__3580  (.L_HI(net3580));
 sg13g2_tiehi \cpu.uart.r_in[0]$_DFFE_PP__3581  (.L_HI(net3581));
 sg13g2_tiehi \cpu.uart.r_in[1]$_DFFE_PP__3582  (.L_HI(net3582));
 sg13g2_tiehi \cpu.uart.r_in[2]$_DFFE_PP__3583  (.L_HI(net3583));
 sg13g2_tiehi \cpu.uart.r_in[3]$_DFFE_PP__3584  (.L_HI(net3584));
 sg13g2_tiehi \cpu.uart.r_in[4]$_DFFE_PP__3585  (.L_HI(net3585));
 sg13g2_tiehi \cpu.uart.r_in[5]$_DFFE_PP__3586  (.L_HI(net3586));
 sg13g2_tiehi \cpu.uart.r_in[6]$_DFFE_PP__3587  (.L_HI(net3587));
 sg13g2_tiehi \cpu.uart.r_in[7]$_DFFE_PP__3588  (.L_HI(net3588));
 sg13g2_tiehi \cpu.uart.r_out[0]$_DFFE_PP__3589  (.L_HI(net3589));
 sg13g2_tiehi \cpu.uart.r_out[1]$_DFFE_PP__3590  (.L_HI(net3590));
 sg13g2_tiehi \cpu.uart.r_out[2]$_DFFE_PP__3591  (.L_HI(net3591));
 sg13g2_tiehi \cpu.uart.r_out[3]$_DFFE_PP__3592  (.L_HI(net3592));
 sg13g2_tiehi \cpu.uart.r_out[4]$_DFFE_PP__3593  (.L_HI(net3593));
 sg13g2_tiehi \cpu.uart.r_out[5]$_DFFE_PP__3594  (.L_HI(net3594));
 sg13g2_tiehi \cpu.uart.r_out[6]$_DFFE_PP__3595  (.L_HI(net3595));
 sg13g2_tiehi \cpu.uart.r_out[7]$_DFFE_PP__3596  (.L_HI(net3596));
 sg13g2_tiehi \cpu.uart.r_r$_DFF_P__3597  (.L_HI(net3597));
 sg13g2_tiehi \cpu.uart.r_r_int$_SDFFE_PN0P__3598  (.L_HI(net3598));
 sg13g2_tiehi \cpu.uart.r_r_invert$_SDFFE_PN0P__3599  (.L_HI(net3599));
 sg13g2_tiehi \cpu.uart.r_rcnt[0]$_DFFE_PP__3600  (.L_HI(net3600));
 sg13g2_tiehi \cpu.uart.r_rcnt[1]$_DFFE_PP__3601  (.L_HI(net3601));
 sg13g2_tiehi \cpu.uart.r_rstate[0]$_SDFFE_PN0P__3602  (.L_HI(net3602));
 sg13g2_tiehi \cpu.uart.r_rstate[1]$_SDFFE_PN0P__3603  (.L_HI(net3603));
 sg13g2_tiehi \cpu.uart.r_rstate[2]$_SDFFE_PN0P__3604  (.L_HI(net3604));
 sg13g2_tiehi \cpu.uart.r_rstate[3]$_SDFFE_PN0P__3605  (.L_HI(net3605));
 sg13g2_tiehi \cpu.uart.r_x$_DFFE_PP__3606  (.L_HI(net3606));
 sg13g2_tiehi \cpu.uart.r_x_int$_SDFFE_PN0P__3607  (.L_HI(net3607));
 sg13g2_tiehi \cpu.uart.r_x_invert$_SDFFE_PN0P__3608  (.L_HI(net3608));
 sg13g2_tiehi \cpu.uart.r_xcnt[0]$_DFFE_PP__3609  (.L_HI(net3609));
 sg13g2_tiehi \cpu.uart.r_xcnt[1]$_DFFE_PP__3610  (.L_HI(net3610));
 sg13g2_tiehi \cpu.uart.r_xstate[0]$_SDFFE_PN0P__3611  (.L_HI(net3611));
 sg13g2_tiehi \cpu.uart.r_xstate[1]$_SDFFE_PN0P__3612  (.L_HI(net3612));
 sg13g2_tiehi \cpu.uart.r_xstate[2]$_SDFFE_PN0P__3613  (.L_HI(net3613));
 sg13g2_tiehi \cpu.uart.r_xstate[3]$_SDFFE_PN0P__3614  (.L_HI(net3614));
 sg13g2_tiehi \r_reset$_DFF_P__3615  (.L_HI(net3615));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_8 clkbuf_leaf_311_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_8 clkbuf_leaf_312_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_0__f_clk (.X(clknet_6_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_1__f_clk (.X(clknet_6_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_2__f_clk (.X(clknet_6_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_3__f_clk (.X(clknet_6_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_4__f_clk (.X(clknet_6_4__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_5__f_clk (.X(clknet_6_5__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_6__f_clk (.X(clknet_6_6__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_7__f_clk (.X(clknet_6_7__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_8__f_clk (.X(clknet_6_8__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_9__f_clk (.X(clknet_6_9__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_10__f_clk (.X(clknet_6_10__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_11__f_clk (.X(clknet_6_11__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_12__f_clk (.X(clknet_6_12__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_13__f_clk (.X(clknet_6_13__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_14__f_clk (.X(clknet_6_14__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_15__f_clk (.X(clknet_6_15__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_16__f_clk (.X(clknet_6_16__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_17__f_clk (.X(clknet_6_17__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_18__f_clk (.X(clknet_6_18__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_19__f_clk (.X(clknet_6_19__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_20__f_clk (.X(clknet_6_20__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_21__f_clk (.X(clknet_6_21__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_22__f_clk (.X(clknet_6_22__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_23__f_clk (.X(clknet_6_23__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_24__f_clk (.X(clknet_6_24__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_25__f_clk (.X(clknet_6_25__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_26__f_clk (.X(clknet_6_26__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_27__f_clk (.X(clknet_6_27__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_28__f_clk (.X(clknet_6_28__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_29__f_clk (.X(clknet_6_29__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_30__f_clk (.X(clknet_6_30__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_31__f_clk (.X(clknet_6_31__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_32__f_clk (.X(clknet_6_32__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_33__f_clk (.X(clknet_6_33__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_34__f_clk (.X(clknet_6_34__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_35__f_clk (.X(clknet_6_35__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_36__f_clk (.X(clknet_6_36__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_37__f_clk (.X(clknet_6_37__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_38__f_clk (.X(clknet_6_38__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_39__f_clk (.X(clknet_6_39__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_40__f_clk (.X(clknet_6_40__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_41__f_clk (.X(clknet_6_41__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_42__f_clk (.X(clknet_6_42__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_43__f_clk (.X(clknet_6_43__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_44__f_clk (.X(clknet_6_44__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_45__f_clk (.X(clknet_6_45__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_46__f_clk (.X(clknet_6_46__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_47__f_clk (.X(clknet_6_47__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_48__f_clk (.X(clknet_6_48__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_49__f_clk (.X(clknet_6_49__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_50__f_clk (.X(clknet_6_50__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_51__f_clk (.X(clknet_6_51__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_52__f_clk (.X(clknet_6_52__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_53__f_clk (.X(clknet_6_53__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_54__f_clk (.X(clknet_6_54__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_55__f_clk (.X(clknet_6_55__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_56__f_clk (.X(clknet_6_56__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_57__f_clk (.X(clknet_6_57__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_58__f_clk (.X(clknet_6_58__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_59__f_clk (.X(clknet_6_59__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_60__f_clk (.X(clknet_6_60__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_61__f_clk (.X(clknet_6_61__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_62__f_clk (.X(clknet_6_62__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_63__f_clk (.X(clknet_6_63__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_63__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_leaf_312_clk));
 sg13g2_buf_16 clkload8 (.A(clknet_leaf_119_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_120_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_257_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_189_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_179_clk));
 sg13g2_buf_16 clkload13 (.A(clknet_leaf_178_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00928_));
 sg13g2_antennanp ANTENNA_2 (.A(_01057_));
 sg13g2_antennanp ANTENNA_3 (.A(_02823_));
 sg13g2_antennanp ANTENNA_4 (.A(_02823_));
 sg13g2_antennanp ANTENNA_5 (.A(_02823_));
 sg13g2_antennanp ANTENNA_6 (.A(_02823_));
 sg13g2_antennanp ANTENNA_7 (.A(_02823_));
 sg13g2_antennanp ANTENNA_8 (.A(_02823_));
 sg13g2_antennanp ANTENNA_9 (.A(_02823_));
 sg13g2_antennanp ANTENNA_10 (.A(_02823_));
 sg13g2_antennanp ANTENNA_11 (.A(_02823_));
 sg13g2_antennanp ANTENNA_12 (.A(_02831_));
 sg13g2_antennanp ANTENNA_13 (.A(_02831_));
 sg13g2_antennanp ANTENNA_14 (.A(_02831_));
 sg13g2_antennanp ANTENNA_15 (.A(_02831_));
 sg13g2_antennanp ANTENNA_16 (.A(_02831_));
 sg13g2_antennanp ANTENNA_17 (.A(_02831_));
 sg13g2_antennanp ANTENNA_18 (.A(_02831_));
 sg13g2_antennanp ANTENNA_19 (.A(_02831_));
 sg13g2_antennanp ANTENNA_20 (.A(_02831_));
 sg13g2_antennanp ANTENNA_21 (.A(_02835_));
 sg13g2_antennanp ANTENNA_22 (.A(_02835_));
 sg13g2_antennanp ANTENNA_23 (.A(_02835_));
 sg13g2_antennanp ANTENNA_24 (.A(_02835_));
 sg13g2_antennanp ANTENNA_25 (.A(_02835_));
 sg13g2_antennanp ANTENNA_26 (.A(_02835_));
 sg13g2_antennanp ANTENNA_27 (.A(_02835_));
 sg13g2_antennanp ANTENNA_28 (.A(_02835_));
 sg13g2_antennanp ANTENNA_29 (.A(_02835_));
 sg13g2_antennanp ANTENNA_30 (.A(_02990_));
 sg13g2_antennanp ANTENNA_31 (.A(_02990_));
 sg13g2_antennanp ANTENNA_32 (.A(_02990_));
 sg13g2_antennanp ANTENNA_33 (.A(_02990_));
 sg13g2_antennanp ANTENNA_34 (.A(_02990_));
 sg13g2_antennanp ANTENNA_35 (.A(_02990_));
 sg13g2_antennanp ANTENNA_36 (.A(_02990_));
 sg13g2_antennanp ANTENNA_37 (.A(_02990_));
 sg13g2_antennanp ANTENNA_38 (.A(_02990_));
 sg13g2_antennanp ANTENNA_39 (.A(_03019_));
 sg13g2_antennanp ANTENNA_40 (.A(_03019_));
 sg13g2_antennanp ANTENNA_41 (.A(_03019_));
 sg13g2_antennanp ANTENNA_42 (.A(_03865_));
 sg13g2_antennanp ANTENNA_43 (.A(_03865_));
 sg13g2_antennanp ANTENNA_44 (.A(_03865_));
 sg13g2_antennanp ANTENNA_45 (.A(_03865_));
 sg13g2_antennanp ANTENNA_46 (.A(_03865_));
 sg13g2_antennanp ANTENNA_47 (.A(_03865_));
 sg13g2_antennanp ANTENNA_48 (.A(_04809_));
 sg13g2_antennanp ANTENNA_49 (.A(_04809_));
 sg13g2_antennanp ANTENNA_50 (.A(_04809_));
 sg13g2_antennanp ANTENNA_51 (.A(_04809_));
 sg13g2_antennanp ANTENNA_52 (.A(_04943_));
 sg13g2_antennanp ANTENNA_53 (.A(_04943_));
 sg13g2_antennanp ANTENNA_54 (.A(_04943_));
 sg13g2_antennanp ANTENNA_55 (.A(_04943_));
 sg13g2_antennanp ANTENNA_56 (.A(_04943_));
 sg13g2_antennanp ANTENNA_57 (.A(_04943_));
 sg13g2_antennanp ANTENNA_58 (.A(_04943_));
 sg13g2_antennanp ANTENNA_59 (.A(_05015_));
 sg13g2_antennanp ANTENNA_60 (.A(_05189_));
 sg13g2_antennanp ANTENNA_61 (.A(_05223_));
 sg13g2_antennanp ANTENNA_62 (.A(_05238_));
 sg13g2_antennanp ANTENNA_63 (.A(_05254_));
 sg13g2_antennanp ANTENNA_64 (.A(_05278_));
 sg13g2_antennanp ANTENNA_65 (.A(_05279_));
 sg13g2_antennanp ANTENNA_66 (.A(_05291_));
 sg13g2_antennanp ANTENNA_67 (.A(_05306_));
 sg13g2_antennanp ANTENNA_68 (.A(_05323_));
 sg13g2_antennanp ANTENNA_69 (.A(_05333_));
 sg13g2_antennanp ANTENNA_70 (.A(_05333_));
 sg13g2_antennanp ANTENNA_71 (.A(_05406_));
 sg13g2_antennanp ANTENNA_72 (.A(_05406_));
 sg13g2_antennanp ANTENNA_73 (.A(_05406_));
 sg13g2_antennanp ANTENNA_74 (.A(_05406_));
 sg13g2_antennanp ANTENNA_75 (.A(_05478_));
 sg13g2_antennanp ANTENNA_76 (.A(_05483_));
 sg13g2_antennanp ANTENNA_77 (.A(_05545_));
 sg13g2_antennanp ANTENNA_78 (.A(_05551_));
 sg13g2_antennanp ANTENNA_79 (.A(_05688_));
 sg13g2_antennanp ANTENNA_80 (.A(_05693_));
 sg13g2_antennanp ANTENNA_81 (.A(_05781_));
 sg13g2_antennanp ANTENNA_82 (.A(_05797_));
 sg13g2_antennanp ANTENNA_83 (.A(_05797_));
 sg13g2_antennanp ANTENNA_84 (.A(_05798_));
 sg13g2_antennanp ANTENNA_85 (.A(_05798_));
 sg13g2_antennanp ANTENNA_86 (.A(_05798_));
 sg13g2_antennanp ANTENNA_87 (.A(_05798_));
 sg13g2_antennanp ANTENNA_88 (.A(_05798_));
 sg13g2_antennanp ANTENNA_89 (.A(_05798_));
 sg13g2_antennanp ANTENNA_90 (.A(_05801_));
 sg13g2_antennanp ANTENNA_91 (.A(_05801_));
 sg13g2_antennanp ANTENNA_92 (.A(_05801_));
 sg13g2_antennanp ANTENNA_93 (.A(_05811_));
 sg13g2_antennanp ANTENNA_94 (.A(_05815_));
 sg13g2_antennanp ANTENNA_95 (.A(_05818_));
 sg13g2_antennanp ANTENNA_96 (.A(_05818_));
 sg13g2_antennanp ANTENNA_97 (.A(_06734_));
 sg13g2_antennanp ANTENNA_98 (.A(_06734_));
 sg13g2_antennanp ANTENNA_99 (.A(_06734_));
 sg13g2_antennanp ANTENNA_100 (.A(_06734_));
 sg13g2_antennanp ANTENNA_101 (.A(_06734_));
 sg13g2_antennanp ANTENNA_102 (.A(_06734_));
 sg13g2_antennanp ANTENNA_103 (.A(_06734_));
 sg13g2_antennanp ANTENNA_104 (.A(_06734_));
 sg13g2_antennanp ANTENNA_105 (.A(_06734_));
 sg13g2_antennanp ANTENNA_106 (.A(_06734_));
 sg13g2_antennanp ANTENNA_107 (.A(_06734_));
 sg13g2_antennanp ANTENNA_108 (.A(_06734_));
 sg13g2_antennanp ANTENNA_109 (.A(_06734_));
 sg13g2_antennanp ANTENNA_110 (.A(_06734_));
 sg13g2_antennanp ANTENNA_111 (.A(_06735_));
 sg13g2_antennanp ANTENNA_112 (.A(_06735_));
 sg13g2_antennanp ANTENNA_113 (.A(_06735_));
 sg13g2_antennanp ANTENNA_114 (.A(_07301_));
 sg13g2_antennanp ANTENNA_115 (.A(_07601_));
 sg13g2_antennanp ANTENNA_116 (.A(_07601_));
 sg13g2_antennanp ANTENNA_117 (.A(_07601_));
 sg13g2_antennanp ANTENNA_118 (.A(_07601_));
 sg13g2_antennanp ANTENNA_119 (.A(_07601_));
 sg13g2_antennanp ANTENNA_120 (.A(_07601_));
 sg13g2_antennanp ANTENNA_121 (.A(_07601_));
 sg13g2_antennanp ANTENNA_122 (.A(_07601_));
 sg13g2_antennanp ANTENNA_123 (.A(_07601_));
 sg13g2_antennanp ANTENNA_124 (.A(_07601_));
 sg13g2_antennanp ANTENNA_125 (.A(_07611_));
 sg13g2_antennanp ANTENNA_126 (.A(_07611_));
 sg13g2_antennanp ANTENNA_127 (.A(_07611_));
 sg13g2_antennanp ANTENNA_128 (.A(_07611_));
 sg13g2_antennanp ANTENNA_129 (.A(_07756_));
 sg13g2_antennanp ANTENNA_130 (.A(_07756_));
 sg13g2_antennanp ANTENNA_131 (.A(_07756_));
 sg13g2_antennanp ANTENNA_132 (.A(_08260_));
 sg13g2_antennanp ANTENNA_133 (.A(_08260_));
 sg13g2_antennanp ANTENNA_134 (.A(_08260_));
 sg13g2_antennanp ANTENNA_135 (.A(_08260_));
 sg13g2_antennanp ANTENNA_136 (.A(_08260_));
 sg13g2_antennanp ANTENNA_137 (.A(_08260_));
 sg13g2_antennanp ANTENNA_138 (.A(_08260_));
 sg13g2_antennanp ANTENNA_139 (.A(_08260_));
 sg13g2_antennanp ANTENNA_140 (.A(_08278_));
 sg13g2_antennanp ANTENNA_141 (.A(_08278_));
 sg13g2_antennanp ANTENNA_142 (.A(_08278_));
 sg13g2_antennanp ANTENNA_143 (.A(_08278_));
 sg13g2_antennanp ANTENNA_144 (.A(_08648_));
 sg13g2_antennanp ANTENNA_145 (.A(_08648_));
 sg13g2_antennanp ANTENNA_146 (.A(_08648_));
 sg13g2_antennanp ANTENNA_147 (.A(_08648_));
 sg13g2_antennanp ANTENNA_148 (.A(_08648_));
 sg13g2_antennanp ANTENNA_149 (.A(_08648_));
 sg13g2_antennanp ANTENNA_150 (.A(_08681_));
 sg13g2_antennanp ANTENNA_151 (.A(_08681_));
 sg13g2_antennanp ANTENNA_152 (.A(_08681_));
 sg13g2_antennanp ANTENNA_153 (.A(_08681_));
 sg13g2_antennanp ANTENNA_154 (.A(_08681_));
 sg13g2_antennanp ANTENNA_155 (.A(_08681_));
 sg13g2_antennanp ANTENNA_156 (.A(_08681_));
 sg13g2_antennanp ANTENNA_157 (.A(_08681_));
 sg13g2_antennanp ANTENNA_158 (.A(_08681_));
 sg13g2_antennanp ANTENNA_159 (.A(_08712_));
 sg13g2_antennanp ANTENNA_160 (.A(_08735_));
 sg13g2_antennanp ANTENNA_161 (.A(_08735_));
 sg13g2_antennanp ANTENNA_162 (.A(_08735_));
 sg13g2_antennanp ANTENNA_163 (.A(_08735_));
 sg13g2_antennanp ANTENNA_164 (.A(_08735_));
 sg13g2_antennanp ANTENNA_165 (.A(_08735_));
 sg13g2_antennanp ANTENNA_166 (.A(_08735_));
 sg13g2_antennanp ANTENNA_167 (.A(_08735_));
 sg13g2_antennanp ANTENNA_168 (.A(_08735_));
 sg13g2_antennanp ANTENNA_169 (.A(_08735_));
 sg13g2_antennanp ANTENNA_170 (.A(_08758_));
 sg13g2_antennanp ANTENNA_171 (.A(_08758_));
 sg13g2_antennanp ANTENNA_172 (.A(_08758_));
 sg13g2_antennanp ANTENNA_173 (.A(_08758_));
 sg13g2_antennanp ANTENNA_174 (.A(_08758_));
 sg13g2_antennanp ANTENNA_175 (.A(_08758_));
 sg13g2_antennanp ANTENNA_176 (.A(_08758_));
 sg13g2_antennanp ANTENNA_177 (.A(_08758_));
 sg13g2_antennanp ANTENNA_178 (.A(_08758_));
 sg13g2_antennanp ANTENNA_179 (.A(_08758_));
 sg13g2_antennanp ANTENNA_180 (.A(_08769_));
 sg13g2_antennanp ANTENNA_181 (.A(_08769_));
 sg13g2_antennanp ANTENNA_182 (.A(_08769_));
 sg13g2_antennanp ANTENNA_183 (.A(_08788_));
 sg13g2_antennanp ANTENNA_184 (.A(_08788_));
 sg13g2_antennanp ANTENNA_185 (.A(_08788_));
 sg13g2_antennanp ANTENNA_186 (.A(_08788_));
 sg13g2_antennanp ANTENNA_187 (.A(_08797_));
 sg13g2_antennanp ANTENNA_188 (.A(_08797_));
 sg13g2_antennanp ANTENNA_189 (.A(_08797_));
 sg13g2_antennanp ANTENNA_190 (.A(_08797_));
 sg13g2_antennanp ANTENNA_191 (.A(_08797_));
 sg13g2_antennanp ANTENNA_192 (.A(_08807_));
 sg13g2_antennanp ANTENNA_193 (.A(_08807_));
 sg13g2_antennanp ANTENNA_194 (.A(_08807_));
 sg13g2_antennanp ANTENNA_195 (.A(_08807_));
 sg13g2_antennanp ANTENNA_196 (.A(_08807_));
 sg13g2_antennanp ANTENNA_197 (.A(_08817_));
 sg13g2_antennanp ANTENNA_198 (.A(_08817_));
 sg13g2_antennanp ANTENNA_199 (.A(_08817_));
 sg13g2_antennanp ANTENNA_200 (.A(_08817_));
 sg13g2_antennanp ANTENNA_201 (.A(_08817_));
 sg13g2_antennanp ANTENNA_202 (.A(_08829_));
 sg13g2_antennanp ANTENNA_203 (.A(_08829_));
 sg13g2_antennanp ANTENNA_204 (.A(_08829_));
 sg13g2_antennanp ANTENNA_205 (.A(_08829_));
 sg13g2_antennanp ANTENNA_206 (.A(_08829_));
 sg13g2_antennanp ANTENNA_207 (.A(_08829_));
 sg13g2_antennanp ANTENNA_208 (.A(_08829_));
 sg13g2_antennanp ANTENNA_209 (.A(_08829_));
 sg13g2_antennanp ANTENNA_210 (.A(_08840_));
 sg13g2_antennanp ANTENNA_211 (.A(_08879_));
 sg13g2_antennanp ANTENNA_212 (.A(_08879_));
 sg13g2_antennanp ANTENNA_213 (.A(_08879_));
 sg13g2_antennanp ANTENNA_214 (.A(_08879_));
 sg13g2_antennanp ANTENNA_215 (.A(_08879_));
 sg13g2_antennanp ANTENNA_216 (.A(_08879_));
 sg13g2_antennanp ANTENNA_217 (.A(_08879_));
 sg13g2_antennanp ANTENNA_218 (.A(_08879_));
 sg13g2_antennanp ANTENNA_219 (.A(_08879_));
 sg13g2_antennanp ANTENNA_220 (.A(_08879_));
 sg13g2_antennanp ANTENNA_221 (.A(_08900_));
 sg13g2_antennanp ANTENNA_222 (.A(_08900_));
 sg13g2_antennanp ANTENNA_223 (.A(_08900_));
 sg13g2_antennanp ANTENNA_224 (.A(_08919_));
 sg13g2_antennanp ANTENNA_225 (.A(_08944_));
 sg13g2_antennanp ANTENNA_226 (.A(_08944_));
 sg13g2_antennanp ANTENNA_227 (.A(_08944_));
 sg13g2_antennanp ANTENNA_228 (.A(_08944_));
 sg13g2_antennanp ANTENNA_229 (.A(_08944_));
 sg13g2_antennanp ANTENNA_230 (.A(_08944_));
 sg13g2_antennanp ANTENNA_231 (.A(_08964_));
 sg13g2_antennanp ANTENNA_232 (.A(_08965_));
 sg13g2_antennanp ANTENNA_233 (.A(_08988_));
 sg13g2_antennanp ANTENNA_234 (.A(_08988_));
 sg13g2_antennanp ANTENNA_235 (.A(_08988_));
 sg13g2_antennanp ANTENNA_236 (.A(_08988_));
 sg13g2_antennanp ANTENNA_237 (.A(_08988_));
 sg13g2_antennanp ANTENNA_238 (.A(_08988_));
 sg13g2_antennanp ANTENNA_239 (.A(_08997_));
 sg13g2_antennanp ANTENNA_240 (.A(_09012_));
 sg13g2_antennanp ANTENNA_241 (.A(_09012_));
 sg13g2_antennanp ANTENNA_242 (.A(_09012_));
 sg13g2_antennanp ANTENNA_243 (.A(_09012_));
 sg13g2_antennanp ANTENNA_244 (.A(_09090_));
 sg13g2_antennanp ANTENNA_245 (.A(_09090_));
 sg13g2_antennanp ANTENNA_246 (.A(_09090_));
 sg13g2_antennanp ANTENNA_247 (.A(_09090_));
 sg13g2_antennanp ANTENNA_248 (.A(_09203_));
 sg13g2_antennanp ANTENNA_249 (.A(_09203_));
 sg13g2_antennanp ANTENNA_250 (.A(_09203_));
 sg13g2_antennanp ANTENNA_251 (.A(_09205_));
 sg13g2_antennanp ANTENNA_252 (.A(_09205_));
 sg13g2_antennanp ANTENNA_253 (.A(_09205_));
 sg13g2_antennanp ANTENNA_254 (.A(_09205_));
 sg13g2_antennanp ANTENNA_255 (.A(_09255_));
 sg13g2_antennanp ANTENNA_256 (.A(_09255_));
 sg13g2_antennanp ANTENNA_257 (.A(_09255_));
 sg13g2_antennanp ANTENNA_258 (.A(_09255_));
 sg13g2_antennanp ANTENNA_259 (.A(_09258_));
 sg13g2_antennanp ANTENNA_260 (.A(_09258_));
 sg13g2_antennanp ANTENNA_261 (.A(_09258_));
 sg13g2_antennanp ANTENNA_262 (.A(_09258_));
 sg13g2_antennanp ANTENNA_263 (.A(_09260_));
 sg13g2_antennanp ANTENNA_264 (.A(_09266_));
 sg13g2_antennanp ANTENNA_265 (.A(_09266_));
 sg13g2_antennanp ANTENNA_266 (.A(_09266_));
 sg13g2_antennanp ANTENNA_267 (.A(_09266_));
 sg13g2_antennanp ANTENNA_268 (.A(_09266_));
 sg13g2_antennanp ANTENNA_269 (.A(_09266_));
 sg13g2_antennanp ANTENNA_270 (.A(_09294_));
 sg13g2_antennanp ANTENNA_271 (.A(_09294_));
 sg13g2_antennanp ANTENNA_272 (.A(_09294_));
 sg13g2_antennanp ANTENNA_273 (.A(_09294_));
 sg13g2_antennanp ANTENNA_274 (.A(_09297_));
 sg13g2_antennanp ANTENNA_275 (.A(_09297_));
 sg13g2_antennanp ANTENNA_276 (.A(_09297_));
 sg13g2_antennanp ANTENNA_277 (.A(_09297_));
 sg13g2_antennanp ANTENNA_278 (.A(_09463_));
 sg13g2_antennanp ANTENNA_279 (.A(_09488_));
 sg13g2_antennanp ANTENNA_280 (.A(_09512_));
 sg13g2_antennanp ANTENNA_281 (.A(_09524_));
 sg13g2_antennanp ANTENNA_282 (.A(_09524_));
 sg13g2_antennanp ANTENNA_283 (.A(_09524_));
 sg13g2_antennanp ANTENNA_284 (.A(_09544_));
 sg13g2_antennanp ANTENNA_285 (.A(_09552_));
 sg13g2_antennanp ANTENNA_286 (.A(_09639_));
 sg13g2_antennanp ANTENNA_287 (.A(_09664_));
 sg13g2_antennanp ANTENNA_288 (.A(_09685_));
 sg13g2_antennanp ANTENNA_289 (.A(_09712_));
 sg13g2_antennanp ANTENNA_290 (.A(_09727_));
 sg13g2_antennanp ANTENNA_291 (.A(_09744_));
 sg13g2_antennanp ANTENNA_292 (.A(_09744_));
 sg13g2_antennanp ANTENNA_293 (.A(_09744_));
 sg13g2_antennanp ANTENNA_294 (.A(_09744_));
 sg13g2_antennanp ANTENNA_295 (.A(_09744_));
 sg13g2_antennanp ANTENNA_296 (.A(_09753_));
 sg13g2_antennanp ANTENNA_297 (.A(_09775_));
 sg13g2_antennanp ANTENNA_298 (.A(_09798_));
 sg13g2_antennanp ANTENNA_299 (.A(_09954_));
 sg13g2_antennanp ANTENNA_300 (.A(_09954_));
 sg13g2_antennanp ANTENNA_301 (.A(_09954_));
 sg13g2_antennanp ANTENNA_302 (.A(_10047_));
 sg13g2_antennanp ANTENNA_303 (.A(_10047_));
 sg13g2_antennanp ANTENNA_304 (.A(_10047_));
 sg13g2_antennanp ANTENNA_305 (.A(_10047_));
 sg13g2_antennanp ANTENNA_306 (.A(_10047_));
 sg13g2_antennanp ANTENNA_307 (.A(_10047_));
 sg13g2_antennanp ANTENNA_308 (.A(_10047_));
 sg13g2_antennanp ANTENNA_309 (.A(_10047_));
 sg13g2_antennanp ANTENNA_310 (.A(_10047_));
 sg13g2_antennanp ANTENNA_311 (.A(_10054_));
 sg13g2_antennanp ANTENNA_312 (.A(_10054_));
 sg13g2_antennanp ANTENNA_313 (.A(_10054_));
 sg13g2_antennanp ANTENNA_314 (.A(_10054_));
 sg13g2_antennanp ANTENNA_315 (.A(_10054_));
 sg13g2_antennanp ANTENNA_316 (.A(_10054_));
 sg13g2_antennanp ANTENNA_317 (.A(_10054_));
 sg13g2_antennanp ANTENNA_318 (.A(_10054_));
 sg13g2_antennanp ANTENNA_319 (.A(_10054_));
 sg13g2_antennanp ANTENNA_320 (.A(_10054_));
 sg13g2_antennanp ANTENNA_321 (.A(_10057_));
 sg13g2_antennanp ANTENNA_322 (.A(_10057_));
 sg13g2_antennanp ANTENNA_323 (.A(_10057_));
 sg13g2_antennanp ANTENNA_324 (.A(_10057_));
 sg13g2_antennanp ANTENNA_325 (.A(_10057_));
 sg13g2_antennanp ANTENNA_326 (.A(_10057_));
 sg13g2_antennanp ANTENNA_327 (.A(_10057_));
 sg13g2_antennanp ANTENNA_328 (.A(_10057_));
 sg13g2_antennanp ANTENNA_329 (.A(_10057_));
 sg13g2_antennanp ANTENNA_330 (.A(_10085_));
 sg13g2_antennanp ANTENNA_331 (.A(_10085_));
 sg13g2_antennanp ANTENNA_332 (.A(_10085_));
 sg13g2_antennanp ANTENNA_333 (.A(_10085_));
 sg13g2_antennanp ANTENNA_334 (.A(_10085_));
 sg13g2_antennanp ANTENNA_335 (.A(_10085_));
 sg13g2_antennanp ANTENNA_336 (.A(_10085_));
 sg13g2_antennanp ANTENNA_337 (.A(_10085_));
 sg13g2_antennanp ANTENNA_338 (.A(_10105_));
 sg13g2_antennanp ANTENNA_339 (.A(_10105_));
 sg13g2_antennanp ANTENNA_340 (.A(_10105_));
 sg13g2_antennanp ANTENNA_341 (.A(_10107_));
 sg13g2_antennanp ANTENNA_342 (.A(_10107_));
 sg13g2_antennanp ANTENNA_343 (.A(_10107_));
 sg13g2_antennanp ANTENNA_344 (.A(_10107_));
 sg13g2_antennanp ANTENNA_345 (.A(_10107_));
 sg13g2_antennanp ANTENNA_346 (.A(_10107_));
 sg13g2_antennanp ANTENNA_347 (.A(_10107_));
 sg13g2_antennanp ANTENNA_348 (.A(_10107_));
 sg13g2_antennanp ANTENNA_349 (.A(_10107_));
 sg13g2_antennanp ANTENNA_350 (.A(_10107_));
 sg13g2_antennanp ANTENNA_351 (.A(_10181_));
 sg13g2_antennanp ANTENNA_352 (.A(_10181_));
 sg13g2_antennanp ANTENNA_353 (.A(_10181_));
 sg13g2_antennanp ANTENNA_354 (.A(_10181_));
 sg13g2_antennanp ANTENNA_355 (.A(_10181_));
 sg13g2_antennanp ANTENNA_356 (.A(_10181_));
 sg13g2_antennanp ANTENNA_357 (.A(_10181_));
 sg13g2_antennanp ANTENNA_358 (.A(_10191_));
 sg13g2_antennanp ANTENNA_359 (.A(_10191_));
 sg13g2_antennanp ANTENNA_360 (.A(_10191_));
 sg13g2_antennanp ANTENNA_361 (.A(_10191_));
 sg13g2_antennanp ANTENNA_362 (.A(_10191_));
 sg13g2_antennanp ANTENNA_363 (.A(_10191_));
 sg13g2_antennanp ANTENNA_364 (.A(_10191_));
 sg13g2_antennanp ANTENNA_365 (.A(_10191_));
 sg13g2_antennanp ANTENNA_366 (.A(_10338_));
 sg13g2_antennanp ANTENNA_367 (.A(_10338_));
 sg13g2_antennanp ANTENNA_368 (.A(_10338_));
 sg13g2_antennanp ANTENNA_369 (.A(_10386_));
 sg13g2_antennanp ANTENNA_370 (.A(_10386_));
 sg13g2_antennanp ANTENNA_371 (.A(_10572_));
 sg13g2_antennanp ANTENNA_372 (.A(_10572_));
 sg13g2_antennanp ANTENNA_373 (.A(_10572_));
 sg13g2_antennanp ANTENNA_374 (.A(_10572_));
 sg13g2_antennanp ANTENNA_375 (.A(_10703_));
 sg13g2_antennanp ANTENNA_376 (.A(_10703_));
 sg13g2_antennanp ANTENNA_377 (.A(_10703_));
 sg13g2_antennanp ANTENNA_378 (.A(_10889_));
 sg13g2_antennanp ANTENNA_379 (.A(_10889_));
 sg13g2_antennanp ANTENNA_380 (.A(_10889_));
 sg13g2_antennanp ANTENNA_381 (.A(_11284_));
 sg13g2_antennanp ANTENNA_382 (.A(_11284_));
 sg13g2_antennanp ANTENNA_383 (.A(_11284_));
 sg13g2_antennanp ANTENNA_384 (.A(_11284_));
 sg13g2_antennanp ANTENNA_385 (.A(_11284_));
 sg13g2_antennanp ANTENNA_386 (.A(_11284_));
 sg13g2_antennanp ANTENNA_387 (.A(_11885_));
 sg13g2_antennanp ANTENNA_388 (.A(_11885_));
 sg13g2_antennanp ANTENNA_389 (.A(_11885_));
 sg13g2_antennanp ANTENNA_390 (.A(_11970_));
 sg13g2_antennanp ANTENNA_391 (.A(_11970_));
 sg13g2_antennanp ANTENNA_392 (.A(_11970_));
 sg13g2_antennanp ANTENNA_393 (.A(_12023_));
 sg13g2_antennanp ANTENNA_394 (.A(_12023_));
 sg13g2_antennanp ANTENNA_395 (.A(_12023_));
 sg13g2_antennanp ANTENNA_396 (.A(_12023_));
 sg13g2_antennanp ANTENNA_397 (.A(_12023_));
 sg13g2_antennanp ANTENNA_398 (.A(_12023_));
 sg13g2_antennanp ANTENNA_399 (.A(_12023_));
 sg13g2_antennanp ANTENNA_400 (.A(_12023_));
 sg13g2_antennanp ANTENNA_401 (.A(_12023_));
 sg13g2_antennanp ANTENNA_402 (.A(_12046_));
 sg13g2_antennanp ANTENNA_403 (.A(_12046_));
 sg13g2_antennanp ANTENNA_404 (.A(_12046_));
 sg13g2_antennanp ANTENNA_405 (.A(_12046_));
 sg13g2_antennanp ANTENNA_406 (.A(_12046_));
 sg13g2_antennanp ANTENNA_407 (.A(_12046_));
 sg13g2_antennanp ANTENNA_408 (.A(_12046_));
 sg13g2_antennanp ANTENNA_409 (.A(_12046_));
 sg13g2_antennanp ANTENNA_410 (.A(_12046_));
 sg13g2_antennanp ANTENNA_411 (.A(_12063_));
 sg13g2_antennanp ANTENNA_412 (.A(_12063_));
 sg13g2_antennanp ANTENNA_413 (.A(_12063_));
 sg13g2_antennanp ANTENNA_414 (.A(_12063_));
 sg13g2_antennanp ANTENNA_415 (.A(_12063_));
 sg13g2_antennanp ANTENNA_416 (.A(_12063_));
 sg13g2_antennanp ANTENNA_417 (.A(_12063_));
 sg13g2_antennanp ANTENNA_418 (.A(_12063_));
 sg13g2_antennanp ANTENNA_419 (.A(_12063_));
 sg13g2_antennanp ANTENNA_420 (.A(_12073_));
 sg13g2_antennanp ANTENNA_421 (.A(_12073_));
 sg13g2_antennanp ANTENNA_422 (.A(_12073_));
 sg13g2_antennanp ANTENNA_423 (.A(_12073_));
 sg13g2_antennanp ANTENNA_424 (.A(_12073_));
 sg13g2_antennanp ANTENNA_425 (.A(_12073_));
 sg13g2_antennanp ANTENNA_426 (.A(_12073_));
 sg13g2_antennanp ANTENNA_427 (.A(_12073_));
 sg13g2_antennanp ANTENNA_428 (.A(_12073_));
 sg13g2_antennanp ANTENNA_429 (.A(_12084_));
 sg13g2_antennanp ANTENNA_430 (.A(_12084_));
 sg13g2_antennanp ANTENNA_431 (.A(_12084_));
 sg13g2_antennanp ANTENNA_432 (.A(_12096_));
 sg13g2_antennanp ANTENNA_433 (.A(_12096_));
 sg13g2_antennanp ANTENNA_434 (.A(_12096_));
 sg13g2_antennanp ANTENNA_435 (.A(_12096_));
 sg13g2_antennanp ANTENNA_436 (.A(_12096_));
 sg13g2_antennanp ANTENNA_437 (.A(_12096_));
 sg13g2_antennanp ANTENNA_438 (.A(_12096_));
 sg13g2_antennanp ANTENNA_439 (.A(_12096_));
 sg13g2_antennanp ANTENNA_440 (.A(_12096_));
 sg13g2_antennanp ANTENNA_441 (.A(_12133_));
 sg13g2_antennanp ANTENNA_442 (.A(_12133_));
 sg13g2_antennanp ANTENNA_443 (.A(_12133_));
 sg13g2_antennanp ANTENNA_444 (.A(_12133_));
 sg13g2_antennanp ANTENNA_445 (.A(_12133_));
 sg13g2_antennanp ANTENNA_446 (.A(_12133_));
 sg13g2_antennanp ANTENNA_447 (.A(_12133_));
 sg13g2_antennanp ANTENNA_448 (.A(_12133_));
 sg13g2_antennanp ANTENNA_449 (.A(_12133_));
 sg13g2_antennanp ANTENNA_450 (.A(_12133_));
 sg13g2_antennanp ANTENNA_451 (.A(clk));
 sg13g2_antennanp ANTENNA_452 (.A(clk));
 sg13g2_antennanp ANTENNA_453 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_454 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_455 (.A(\cpu.ex.r_cc ));
 sg13g2_antennanp ANTENNA_456 (.A(\cpu.ex.r_cc ));
 sg13g2_antennanp ANTENNA_457 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_458 (.A(r_reset));
 sg13g2_antennanp ANTENNA_459 (.A(r_reset));
 sg13g2_antennanp ANTENNA_460 (.A(r_reset));
 sg13g2_antennanp ANTENNA_461 (.A(net1));
 sg13g2_antennanp ANTENNA_462 (.A(net1));
 sg13g2_antennanp ANTENNA_463 (.A(net1));
 sg13g2_antennanp ANTENNA_464 (.A(net2));
 sg13g2_antennanp ANTENNA_465 (.A(net2));
 sg13g2_antennanp ANTENNA_466 (.A(net3));
 sg13g2_antennanp ANTENNA_467 (.A(net3));
 sg13g2_antennanp ANTENNA_468 (.A(net3));
 sg13g2_antennanp ANTENNA_469 (.A(net11));
 sg13g2_antennanp ANTENNA_470 (.A(net11));
 sg13g2_antennanp ANTENNA_471 (.A(net11));
 sg13g2_antennanp ANTENNA_472 (.A(net12));
 sg13g2_antennanp ANTENNA_473 (.A(net12));
 sg13g2_antennanp ANTENNA_474 (.A(net13));
 sg13g2_antennanp ANTENNA_475 (.A(net13));
 sg13g2_antennanp ANTENNA_476 (.A(net14));
 sg13g2_antennanp ANTENNA_477 (.A(net14));
 sg13g2_antennanp ANTENNA_478 (.A(net14));
 sg13g2_antennanp ANTENNA_479 (.A(net19));
 sg13g2_antennanp ANTENNA_480 (.A(net19));
 sg13g2_antennanp ANTENNA_481 (.A(net19));
 sg13g2_antennanp ANTENNA_482 (.A(net20));
 sg13g2_antennanp ANTENNA_483 (.A(net20));
 sg13g2_antennanp ANTENNA_484 (.A(net153));
 sg13g2_antennanp ANTENNA_485 (.A(net153));
 sg13g2_antennanp ANTENNA_486 (.A(net153));
 sg13g2_antennanp ANTENNA_487 (.A(net153));
 sg13g2_antennanp ANTENNA_488 (.A(net153));
 sg13g2_antennanp ANTENNA_489 (.A(net153));
 sg13g2_antennanp ANTENNA_490 (.A(net153));
 sg13g2_antennanp ANTENNA_491 (.A(net153));
 sg13g2_antennanp ANTENNA_492 (.A(net153));
 sg13g2_antennanp ANTENNA_493 (.A(net153));
 sg13g2_antennanp ANTENNA_494 (.A(net153));
 sg13g2_antennanp ANTENNA_495 (.A(net520));
 sg13g2_antennanp ANTENNA_496 (.A(net520));
 sg13g2_antennanp ANTENNA_497 (.A(net520));
 sg13g2_antennanp ANTENNA_498 (.A(net520));
 sg13g2_antennanp ANTENNA_499 (.A(net520));
 sg13g2_antennanp ANTENNA_500 (.A(net520));
 sg13g2_antennanp ANTENNA_501 (.A(net520));
 sg13g2_antennanp ANTENNA_502 (.A(net520));
 sg13g2_antennanp ANTENNA_503 (.A(net520));
 sg13g2_antennanp ANTENNA_504 (.A(net520));
 sg13g2_antennanp ANTENNA_505 (.A(net520));
 sg13g2_antennanp ANTENNA_506 (.A(net520));
 sg13g2_antennanp ANTENNA_507 (.A(net520));
 sg13g2_antennanp ANTENNA_508 (.A(net520));
 sg13g2_antennanp ANTENNA_509 (.A(net520));
 sg13g2_antennanp ANTENNA_510 (.A(net520));
 sg13g2_antennanp ANTENNA_511 (.A(net536));
 sg13g2_antennanp ANTENNA_512 (.A(net536));
 sg13g2_antennanp ANTENNA_513 (.A(net536));
 sg13g2_antennanp ANTENNA_514 (.A(net536));
 sg13g2_antennanp ANTENNA_515 (.A(net536));
 sg13g2_antennanp ANTENNA_516 (.A(net536));
 sg13g2_antennanp ANTENNA_517 (.A(net536));
 sg13g2_antennanp ANTENNA_518 (.A(net536));
 sg13g2_antennanp ANTENNA_519 (.A(net536));
 sg13g2_antennanp ANTENNA_520 (.A(net593));
 sg13g2_antennanp ANTENNA_521 (.A(net593));
 sg13g2_antennanp ANTENNA_522 (.A(net593));
 sg13g2_antennanp ANTENNA_523 (.A(net593));
 sg13g2_antennanp ANTENNA_524 (.A(net593));
 sg13g2_antennanp ANTENNA_525 (.A(net593));
 sg13g2_antennanp ANTENNA_526 (.A(net593));
 sg13g2_antennanp ANTENNA_527 (.A(net593));
 sg13g2_antennanp ANTENNA_528 (.A(net593));
 sg13g2_antennanp ANTENNA_529 (.A(net596));
 sg13g2_antennanp ANTENNA_530 (.A(net596));
 sg13g2_antennanp ANTENNA_531 (.A(net596));
 sg13g2_antennanp ANTENNA_532 (.A(net596));
 sg13g2_antennanp ANTENNA_533 (.A(net596));
 sg13g2_antennanp ANTENNA_534 (.A(net596));
 sg13g2_antennanp ANTENNA_535 (.A(net596));
 sg13g2_antennanp ANTENNA_536 (.A(net596));
 sg13g2_antennanp ANTENNA_537 (.A(net618));
 sg13g2_antennanp ANTENNA_538 (.A(net618));
 sg13g2_antennanp ANTENNA_539 (.A(net618));
 sg13g2_antennanp ANTENNA_540 (.A(net618));
 sg13g2_antennanp ANTENNA_541 (.A(net618));
 sg13g2_antennanp ANTENNA_542 (.A(net618));
 sg13g2_antennanp ANTENNA_543 (.A(net618));
 sg13g2_antennanp ANTENNA_544 (.A(net618));
 sg13g2_antennanp ANTENNA_545 (.A(net618));
 sg13g2_antennanp ANTENNA_546 (.A(net618));
 sg13g2_antennanp ANTENNA_547 (.A(net618));
 sg13g2_antennanp ANTENNA_548 (.A(net618));
 sg13g2_antennanp ANTENNA_549 (.A(net618));
 sg13g2_antennanp ANTENNA_550 (.A(net618));
 sg13g2_antennanp ANTENNA_551 (.A(net618));
 sg13g2_antennanp ANTENNA_552 (.A(net623));
 sg13g2_antennanp ANTENNA_553 (.A(net623));
 sg13g2_antennanp ANTENNA_554 (.A(net623));
 sg13g2_antennanp ANTENNA_555 (.A(net623));
 sg13g2_antennanp ANTENNA_556 (.A(net623));
 sg13g2_antennanp ANTENNA_557 (.A(net623));
 sg13g2_antennanp ANTENNA_558 (.A(net623));
 sg13g2_antennanp ANTENNA_559 (.A(net623));
 sg13g2_antennanp ANTENNA_560 (.A(net625));
 sg13g2_antennanp ANTENNA_561 (.A(net625));
 sg13g2_antennanp ANTENNA_562 (.A(net625));
 sg13g2_antennanp ANTENNA_563 (.A(net625));
 sg13g2_antennanp ANTENNA_564 (.A(net625));
 sg13g2_antennanp ANTENNA_565 (.A(net625));
 sg13g2_antennanp ANTENNA_566 (.A(net625));
 sg13g2_antennanp ANTENNA_567 (.A(net625));
 sg13g2_antennanp ANTENNA_568 (.A(net631));
 sg13g2_antennanp ANTENNA_569 (.A(net631));
 sg13g2_antennanp ANTENNA_570 (.A(net631));
 sg13g2_antennanp ANTENNA_571 (.A(net631));
 sg13g2_antennanp ANTENNA_572 (.A(net631));
 sg13g2_antennanp ANTENNA_573 (.A(net631));
 sg13g2_antennanp ANTENNA_574 (.A(net631));
 sg13g2_antennanp ANTENNA_575 (.A(net631));
 sg13g2_antennanp ANTENNA_576 (.A(net631));
 sg13g2_antennanp ANTENNA_577 (.A(net632));
 sg13g2_antennanp ANTENNA_578 (.A(net632));
 sg13g2_antennanp ANTENNA_579 (.A(net632));
 sg13g2_antennanp ANTENNA_580 (.A(net632));
 sg13g2_antennanp ANTENNA_581 (.A(net632));
 sg13g2_antennanp ANTENNA_582 (.A(net632));
 sg13g2_antennanp ANTENNA_583 (.A(net632));
 sg13g2_antennanp ANTENNA_584 (.A(net632));
 sg13g2_antennanp ANTENNA_585 (.A(net632));
 sg13g2_antennanp ANTENNA_586 (.A(net632));
 sg13g2_antennanp ANTENNA_587 (.A(net632));
 sg13g2_antennanp ANTENNA_588 (.A(net632));
 sg13g2_antennanp ANTENNA_589 (.A(net632));
 sg13g2_antennanp ANTENNA_590 (.A(net651));
 sg13g2_antennanp ANTENNA_591 (.A(net651));
 sg13g2_antennanp ANTENNA_592 (.A(net651));
 sg13g2_antennanp ANTENNA_593 (.A(net651));
 sg13g2_antennanp ANTENNA_594 (.A(net651));
 sg13g2_antennanp ANTENNA_595 (.A(net651));
 sg13g2_antennanp ANTENNA_596 (.A(net651));
 sg13g2_antennanp ANTENNA_597 (.A(net651));
 sg13g2_antennanp ANTENNA_598 (.A(net651));
 sg13g2_antennanp ANTENNA_599 (.A(net651));
 sg13g2_antennanp ANTENNA_600 (.A(net651));
 sg13g2_antennanp ANTENNA_601 (.A(net651));
 sg13g2_antennanp ANTENNA_602 (.A(net651));
 sg13g2_antennanp ANTENNA_603 (.A(net651));
 sg13g2_antennanp ANTENNA_604 (.A(net651));
 sg13g2_antennanp ANTENNA_605 (.A(net651));
 sg13g2_antennanp ANTENNA_606 (.A(net702));
 sg13g2_antennanp ANTENNA_607 (.A(net702));
 sg13g2_antennanp ANTENNA_608 (.A(net702));
 sg13g2_antennanp ANTENNA_609 (.A(net702));
 sg13g2_antennanp ANTENNA_610 (.A(net702));
 sg13g2_antennanp ANTENNA_611 (.A(net702));
 sg13g2_antennanp ANTENNA_612 (.A(net702));
 sg13g2_antennanp ANTENNA_613 (.A(net702));
 sg13g2_antennanp ANTENNA_614 (.A(net704));
 sg13g2_antennanp ANTENNA_615 (.A(net704));
 sg13g2_antennanp ANTENNA_616 (.A(net704));
 sg13g2_antennanp ANTENNA_617 (.A(net704));
 sg13g2_antennanp ANTENNA_618 (.A(net704));
 sg13g2_antennanp ANTENNA_619 (.A(net704));
 sg13g2_antennanp ANTENNA_620 (.A(net704));
 sg13g2_antennanp ANTENNA_621 (.A(net704));
 sg13g2_antennanp ANTENNA_622 (.A(net704));
 sg13g2_antennanp ANTENNA_623 (.A(net704));
 sg13g2_antennanp ANTENNA_624 (.A(net704));
 sg13g2_antennanp ANTENNA_625 (.A(net704));
 sg13g2_antennanp ANTENNA_626 (.A(net704));
 sg13g2_antennanp ANTENNA_627 (.A(net704));
 sg13g2_antennanp ANTENNA_628 (.A(net704));
 sg13g2_antennanp ANTENNA_629 (.A(net704));
 sg13g2_antennanp ANTENNA_630 (.A(net704));
 sg13g2_antennanp ANTENNA_631 (.A(net704));
 sg13g2_antennanp ANTENNA_632 (.A(net704));
 sg13g2_antennanp ANTENNA_633 (.A(net704));
 sg13g2_antennanp ANTENNA_634 (.A(net704));
 sg13g2_antennanp ANTENNA_635 (.A(net780));
 sg13g2_antennanp ANTENNA_636 (.A(net780));
 sg13g2_antennanp ANTENNA_637 (.A(net780));
 sg13g2_antennanp ANTENNA_638 (.A(net780));
 sg13g2_antennanp ANTENNA_639 (.A(net780));
 sg13g2_antennanp ANTENNA_640 (.A(net780));
 sg13g2_antennanp ANTENNA_641 (.A(net780));
 sg13g2_antennanp ANTENNA_642 (.A(net780));
 sg13g2_antennanp ANTENNA_643 (.A(net780));
 sg13g2_antennanp ANTENNA_644 (.A(net860));
 sg13g2_antennanp ANTENNA_645 (.A(net860));
 sg13g2_antennanp ANTENNA_646 (.A(net860));
 sg13g2_antennanp ANTENNA_647 (.A(net860));
 sg13g2_antennanp ANTENNA_648 (.A(net860));
 sg13g2_antennanp ANTENNA_649 (.A(net860));
 sg13g2_antennanp ANTENNA_650 (.A(net860));
 sg13g2_antennanp ANTENNA_651 (.A(net860));
 sg13g2_antennanp ANTENNA_652 (.A(net860));
 sg13g2_antennanp ANTENNA_653 (.A(net891));
 sg13g2_antennanp ANTENNA_654 (.A(net891));
 sg13g2_antennanp ANTENNA_655 (.A(net891));
 sg13g2_antennanp ANTENNA_656 (.A(net891));
 sg13g2_antennanp ANTENNA_657 (.A(net891));
 sg13g2_antennanp ANTENNA_658 (.A(net891));
 sg13g2_antennanp ANTENNA_659 (.A(net891));
 sg13g2_antennanp ANTENNA_660 (.A(net891));
 sg13g2_antennanp ANTENNA_661 (.A(net891));
 sg13g2_antennanp ANTENNA_662 (.A(net891));
 sg13g2_antennanp ANTENNA_663 (.A(net891));
 sg13g2_antennanp ANTENNA_664 (.A(net891));
 sg13g2_antennanp ANTENNA_665 (.A(net891));
 sg13g2_antennanp ANTENNA_666 (.A(net891));
 sg13g2_antennanp ANTENNA_667 (.A(net891));
 sg13g2_antennanp ANTENNA_668 (.A(net891));
 sg13g2_antennanp ANTENNA_669 (.A(net895));
 sg13g2_antennanp ANTENNA_670 (.A(net895));
 sg13g2_antennanp ANTENNA_671 (.A(net895));
 sg13g2_antennanp ANTENNA_672 (.A(net895));
 sg13g2_antennanp ANTENNA_673 (.A(net895));
 sg13g2_antennanp ANTENNA_674 (.A(net895));
 sg13g2_antennanp ANTENNA_675 (.A(net895));
 sg13g2_antennanp ANTENNA_676 (.A(net895));
 sg13g2_antennanp ANTENNA_677 (.A(net895));
 sg13g2_antennanp ANTENNA_678 (.A(net895));
 sg13g2_antennanp ANTENNA_679 (.A(net895));
 sg13g2_antennanp ANTENNA_680 (.A(net895));
 sg13g2_antennanp ANTENNA_681 (.A(net895));
 sg13g2_antennanp ANTENNA_682 (.A(net895));
 sg13g2_antennanp ANTENNA_683 (.A(net895));
 sg13g2_antennanp ANTENNA_684 (.A(net895));
 sg13g2_antennanp ANTENNA_685 (.A(net895));
 sg13g2_antennanp ANTENNA_686 (.A(net895));
 sg13g2_antennanp ANTENNA_687 (.A(net895));
 sg13g2_antennanp ANTENNA_688 (.A(net895));
 sg13g2_antennanp ANTENNA_689 (.A(net899));
 sg13g2_antennanp ANTENNA_690 (.A(net899));
 sg13g2_antennanp ANTENNA_691 (.A(net899));
 sg13g2_antennanp ANTENNA_692 (.A(net899));
 sg13g2_antennanp ANTENNA_693 (.A(net899));
 sg13g2_antennanp ANTENNA_694 (.A(net899));
 sg13g2_antennanp ANTENNA_695 (.A(net899));
 sg13g2_antennanp ANTENNA_696 (.A(net899));
 sg13g2_antennanp ANTENNA_697 (.A(net899));
 sg13g2_antennanp ANTENNA_698 (.A(net899));
 sg13g2_antennanp ANTENNA_699 (.A(net899));
 sg13g2_antennanp ANTENNA_700 (.A(net899));
 sg13g2_antennanp ANTENNA_701 (.A(net899));
 sg13g2_antennanp ANTENNA_702 (.A(net899));
 sg13g2_antennanp ANTENNA_703 (.A(net899));
 sg13g2_antennanp ANTENNA_704 (.A(net899));
 sg13g2_antennanp ANTENNA_705 (.A(net899));
 sg13g2_antennanp ANTENNA_706 (.A(net899));
 sg13g2_antennanp ANTENNA_707 (.A(net899));
 sg13g2_antennanp ANTENNA_708 (.A(net899));
 sg13g2_antennanp ANTENNA_709 (.A(net899));
 sg13g2_antennanp ANTENNA_710 (.A(net899));
 sg13g2_antennanp ANTENNA_711 (.A(net899));
 sg13g2_antennanp ANTENNA_712 (.A(net899));
 sg13g2_antennanp ANTENNA_713 (.A(net899));
 sg13g2_antennanp ANTENNA_714 (.A(net899));
 sg13g2_antennanp ANTENNA_715 (.A(net899));
 sg13g2_antennanp ANTENNA_716 (.A(net899));
 sg13g2_antennanp ANTENNA_717 (.A(net899));
 sg13g2_antennanp ANTENNA_718 (.A(net899));
 sg13g2_antennanp ANTENNA_719 (.A(net899));
 sg13g2_antennanp ANTENNA_720 (.A(net899));
 sg13g2_antennanp ANTENNA_721 (.A(net899));
 sg13g2_antennanp ANTENNA_722 (.A(net899));
 sg13g2_antennanp ANTENNA_723 (.A(net899));
 sg13g2_antennanp ANTENNA_724 (.A(net899));
 sg13g2_antennanp ANTENNA_725 (.A(net899));
 sg13g2_antennanp ANTENNA_726 (.A(net899));
 sg13g2_antennanp ANTENNA_727 (.A(net899));
 sg13g2_antennanp ANTENNA_728 (.A(net899));
 sg13g2_antennanp ANTENNA_729 (.A(net899));
 sg13g2_antennanp ANTENNA_730 (.A(net899));
 sg13g2_antennanp ANTENNA_731 (.A(net899));
 sg13g2_antennanp ANTENNA_732 (.A(net899));
 sg13g2_antennanp ANTENNA_733 (.A(net899));
 sg13g2_antennanp ANTENNA_734 (.A(net899));
 sg13g2_antennanp ANTENNA_735 (.A(net959));
 sg13g2_antennanp ANTENNA_736 (.A(net959));
 sg13g2_antennanp ANTENNA_737 (.A(net959));
 sg13g2_antennanp ANTENNA_738 (.A(net959));
 sg13g2_antennanp ANTENNA_739 (.A(net959));
 sg13g2_antennanp ANTENNA_740 (.A(net959));
 sg13g2_antennanp ANTENNA_741 (.A(net959));
 sg13g2_antennanp ANTENNA_742 (.A(net959));
 sg13g2_antennanp ANTENNA_743 (.A(net959));
 sg13g2_antennanp ANTENNA_744 (.A(net959));
 sg13g2_antennanp ANTENNA_745 (.A(net959));
 sg13g2_antennanp ANTENNA_746 (.A(net959));
 sg13g2_antennanp ANTENNA_747 (.A(net967));
 sg13g2_antennanp ANTENNA_748 (.A(net967));
 sg13g2_antennanp ANTENNA_749 (.A(net967));
 sg13g2_antennanp ANTENNA_750 (.A(net967));
 sg13g2_antennanp ANTENNA_751 (.A(net967));
 sg13g2_antennanp ANTENNA_752 (.A(net967));
 sg13g2_antennanp ANTENNA_753 (.A(net967));
 sg13g2_antennanp ANTENNA_754 (.A(net967));
 sg13g2_antennanp ANTENNA_755 (.A(net967));
 sg13g2_antennanp ANTENNA_756 (.A(net969));
 sg13g2_antennanp ANTENNA_757 (.A(net969));
 sg13g2_antennanp ANTENNA_758 (.A(net969));
 sg13g2_antennanp ANTENNA_759 (.A(net969));
 sg13g2_antennanp ANTENNA_760 (.A(net969));
 sg13g2_antennanp ANTENNA_761 (.A(net969));
 sg13g2_antennanp ANTENNA_762 (.A(net969));
 sg13g2_antennanp ANTENNA_763 (.A(net969));
 sg13g2_antennanp ANTENNA_764 (.A(net969));
 sg13g2_antennanp ANTENNA_765 (.A(net970));
 sg13g2_antennanp ANTENNA_766 (.A(net970));
 sg13g2_antennanp ANTENNA_767 (.A(net970));
 sg13g2_antennanp ANTENNA_768 (.A(net970));
 sg13g2_antennanp ANTENNA_769 (.A(net970));
 sg13g2_antennanp ANTENNA_770 (.A(net970));
 sg13g2_antennanp ANTENNA_771 (.A(net970));
 sg13g2_antennanp ANTENNA_772 (.A(net970));
 sg13g2_antennanp ANTENNA_773 (.A(net970));
 sg13g2_antennanp ANTENNA_774 (.A(net970));
 sg13g2_antennanp ANTENNA_775 (.A(net970));
 sg13g2_antennanp ANTENNA_776 (.A(net970));
 sg13g2_antennanp ANTENNA_777 (.A(net970));
 sg13g2_antennanp ANTENNA_778 (.A(net970));
 sg13g2_antennanp ANTENNA_779 (.A(net971));
 sg13g2_antennanp ANTENNA_780 (.A(net971));
 sg13g2_antennanp ANTENNA_781 (.A(net971));
 sg13g2_antennanp ANTENNA_782 (.A(net971));
 sg13g2_antennanp ANTENNA_783 (.A(net971));
 sg13g2_antennanp ANTENNA_784 (.A(net971));
 sg13g2_antennanp ANTENNA_785 (.A(net971));
 sg13g2_antennanp ANTENNA_786 (.A(net971));
 sg13g2_antennanp ANTENNA_787 (.A(net971));
 sg13g2_antennanp ANTENNA_788 (.A(net971));
 sg13g2_antennanp ANTENNA_789 (.A(net971));
 sg13g2_antennanp ANTENNA_790 (.A(net971));
 sg13g2_antennanp ANTENNA_791 (.A(net971));
 sg13g2_antennanp ANTENNA_792 (.A(net971));
 sg13g2_antennanp ANTENNA_793 (.A(net971));
 sg13g2_antennanp ANTENNA_794 (.A(net971));
 sg13g2_antennanp ANTENNA_795 (.A(net972));
 sg13g2_antennanp ANTENNA_796 (.A(net972));
 sg13g2_antennanp ANTENNA_797 (.A(net972));
 sg13g2_antennanp ANTENNA_798 (.A(net972));
 sg13g2_antennanp ANTENNA_799 (.A(net972));
 sg13g2_antennanp ANTENNA_800 (.A(net972));
 sg13g2_antennanp ANTENNA_801 (.A(net972));
 sg13g2_antennanp ANTENNA_802 (.A(net972));
 sg13g2_antennanp ANTENNA_803 (.A(net995));
 sg13g2_antennanp ANTENNA_804 (.A(net995));
 sg13g2_antennanp ANTENNA_805 (.A(net995));
 sg13g2_antennanp ANTENNA_806 (.A(net995));
 sg13g2_antennanp ANTENNA_807 (.A(net995));
 sg13g2_antennanp ANTENNA_808 (.A(net995));
 sg13g2_antennanp ANTENNA_809 (.A(net995));
 sg13g2_antennanp ANTENNA_810 (.A(net995));
 sg13g2_antennanp ANTENNA_811 (.A(net995));
 sg13g2_antennanp ANTENNA_812 (.A(net995));
 sg13g2_antennanp ANTENNA_813 (.A(net995));
 sg13g2_antennanp ANTENNA_814 (.A(net995));
 sg13g2_antennanp ANTENNA_815 (.A(net995));
 sg13g2_antennanp ANTENNA_816 (.A(net995));
 sg13g2_antennanp ANTENNA_817 (.A(net995));
 sg13g2_antennanp ANTENNA_818 (.A(net995));
 sg13g2_antennanp ANTENNA_819 (.A(net995));
 sg13g2_antennanp ANTENNA_820 (.A(net995));
 sg13g2_antennanp ANTENNA_821 (.A(net995));
 sg13g2_antennanp ANTENNA_822 (.A(net995));
 sg13g2_antennanp ANTENNA_823 (.A(net995));
 sg13g2_antennanp ANTENNA_824 (.A(net995));
 sg13g2_antennanp ANTENNA_825 (.A(net995));
 sg13g2_antennanp ANTENNA_826 (.A(net995));
 sg13g2_antennanp ANTENNA_827 (.A(net995));
 sg13g2_antennanp ANTENNA_828 (.A(net995));
 sg13g2_antennanp ANTENNA_829 (.A(net1000));
 sg13g2_antennanp ANTENNA_830 (.A(net1000));
 sg13g2_antennanp ANTENNA_831 (.A(net1000));
 sg13g2_antennanp ANTENNA_832 (.A(net1000));
 sg13g2_antennanp ANTENNA_833 (.A(net1000));
 sg13g2_antennanp ANTENNA_834 (.A(net1000));
 sg13g2_antennanp ANTENNA_835 (.A(net1000));
 sg13g2_antennanp ANTENNA_836 (.A(net1000));
 sg13g2_antennanp ANTENNA_837 (.A(net1000));
 sg13g2_antennanp ANTENNA_838 (.A(net1000));
 sg13g2_antennanp ANTENNA_839 (.A(net1000));
 sg13g2_antennanp ANTENNA_840 (.A(net1000));
 sg13g2_antennanp ANTENNA_841 (.A(net1000));
 sg13g2_antennanp ANTENNA_842 (.A(net1000));
 sg13g2_antennanp ANTENNA_843 (.A(net1028));
 sg13g2_antennanp ANTENNA_844 (.A(net1028));
 sg13g2_antennanp ANTENNA_845 (.A(net1028));
 sg13g2_antennanp ANTENNA_846 (.A(net1028));
 sg13g2_antennanp ANTENNA_847 (.A(net1028));
 sg13g2_antennanp ANTENNA_848 (.A(net1028));
 sg13g2_antennanp ANTENNA_849 (.A(net1028));
 sg13g2_antennanp ANTENNA_850 (.A(net1028));
 sg13g2_antennanp ANTENNA_851 (.A(net1028));
 sg13g2_antennanp ANTENNA_852 (.A(net1028));
 sg13g2_antennanp ANTENNA_853 (.A(net1028));
 sg13g2_antennanp ANTENNA_854 (.A(net1028));
 sg13g2_antennanp ANTENNA_855 (.A(net1028));
 sg13g2_antennanp ANTENNA_856 (.A(net1028));
 sg13g2_antennanp ANTENNA_857 (.A(net1028));
 sg13g2_antennanp ANTENNA_858 (.A(net1028));
 sg13g2_antennanp ANTENNA_859 (.A(net1028));
 sg13g2_antennanp ANTENNA_860 (.A(net1028));
 sg13g2_antennanp ANTENNA_861 (.A(net1028));
 sg13g2_antennanp ANTENNA_862 (.A(net1028));
 sg13g2_antennanp ANTENNA_863 (.A(net1028));
 sg13g2_antennanp ANTENNA_864 (.A(net1028));
 sg13g2_antennanp ANTENNA_865 (.A(net1028));
 sg13g2_antennanp ANTENNA_866 (.A(net1028));
 sg13g2_antennanp ANTENNA_867 (.A(net1028));
 sg13g2_antennanp ANTENNA_868 (.A(net1028));
 sg13g2_antennanp ANTENNA_869 (.A(net1028));
 sg13g2_antennanp ANTENNA_870 (.A(net1028));
 sg13g2_antennanp ANTENNA_871 (.A(net1028));
 sg13g2_antennanp ANTENNA_872 (.A(net1028));
 sg13g2_antennanp ANTENNA_873 (.A(net1028));
 sg13g2_antennanp ANTENNA_874 (.A(net1028));
 sg13g2_antennanp ANTENNA_875 (.A(net1028));
 sg13g2_antennanp ANTENNA_876 (.A(net1042));
 sg13g2_antennanp ANTENNA_877 (.A(net1042));
 sg13g2_antennanp ANTENNA_878 (.A(net1042));
 sg13g2_antennanp ANTENNA_879 (.A(net1042));
 sg13g2_antennanp ANTENNA_880 (.A(net1042));
 sg13g2_antennanp ANTENNA_881 (.A(net1042));
 sg13g2_antennanp ANTENNA_882 (.A(net1042));
 sg13g2_antennanp ANTENNA_883 (.A(net1042));
 sg13g2_antennanp ANTENNA_884 (.A(net1042));
 sg13g2_antennanp ANTENNA_885 (.A(net1042));
 sg13g2_antennanp ANTENNA_886 (.A(net1042));
 sg13g2_antennanp ANTENNA_887 (.A(net1042));
 sg13g2_antennanp ANTENNA_888 (.A(net1042));
 sg13g2_antennanp ANTENNA_889 (.A(net1042));
 sg13g2_antennanp ANTENNA_890 (.A(net1042));
 sg13g2_antennanp ANTENNA_891 (.A(net1042));
 sg13g2_antennanp ANTENNA_892 (.A(net1042));
 sg13g2_antennanp ANTENNA_893 (.A(net1042));
 sg13g2_antennanp ANTENNA_894 (.A(net1042));
 sg13g2_antennanp ANTENNA_895 (.A(net1042));
 sg13g2_antennanp ANTENNA_896 (.A(net1042));
 sg13g2_antennanp ANTENNA_897 (.A(net1042));
 sg13g2_antennanp ANTENNA_898 (.A(net1042));
 sg13g2_antennanp ANTENNA_899 (.A(net1042));
 sg13g2_antennanp ANTENNA_900 (.A(net1042));
 sg13g2_antennanp ANTENNA_901 (.A(net1042));
 sg13g2_antennanp ANTENNA_902 (.A(net1042));
 sg13g2_antennanp ANTENNA_903 (.A(net1042));
 sg13g2_antennanp ANTENNA_904 (.A(net1043));
 sg13g2_antennanp ANTENNA_905 (.A(net1043));
 sg13g2_antennanp ANTENNA_906 (.A(net1043));
 sg13g2_antennanp ANTENNA_907 (.A(net1043));
 sg13g2_antennanp ANTENNA_908 (.A(net1043));
 sg13g2_antennanp ANTENNA_909 (.A(net1043));
 sg13g2_antennanp ANTENNA_910 (.A(net1043));
 sg13g2_antennanp ANTENNA_911 (.A(net1043));
 sg13g2_antennanp ANTENNA_912 (.A(net1043));
 sg13g2_antennanp ANTENNA_913 (.A(net1043));
 sg13g2_antennanp ANTENNA_914 (.A(net1043));
 sg13g2_antennanp ANTENNA_915 (.A(net1043));
 sg13g2_antennanp ANTENNA_916 (.A(net1043));
 sg13g2_antennanp ANTENNA_917 (.A(net1043));
 sg13g2_antennanp ANTENNA_918 (.A(net1043));
 sg13g2_antennanp ANTENNA_919 (.A(net1043));
 sg13g2_antennanp ANTENNA_920 (.A(net1072));
 sg13g2_antennanp ANTENNA_921 (.A(net1072));
 sg13g2_antennanp ANTENNA_922 (.A(net1072));
 sg13g2_antennanp ANTENNA_923 (.A(net1072));
 sg13g2_antennanp ANTENNA_924 (.A(net1072));
 sg13g2_antennanp ANTENNA_925 (.A(net1072));
 sg13g2_antennanp ANTENNA_926 (.A(net1072));
 sg13g2_antennanp ANTENNA_927 (.A(net1072));
 sg13g2_antennanp ANTENNA_928 (.A(net1072));
 sg13g2_antennanp ANTENNA_929 (.A(net1089));
 sg13g2_antennanp ANTENNA_930 (.A(net1089));
 sg13g2_antennanp ANTENNA_931 (.A(net1089));
 sg13g2_antennanp ANTENNA_932 (.A(net1089));
 sg13g2_antennanp ANTENNA_933 (.A(net1089));
 sg13g2_antennanp ANTENNA_934 (.A(net1089));
 sg13g2_antennanp ANTENNA_935 (.A(net1089));
 sg13g2_antennanp ANTENNA_936 (.A(net1089));
 sg13g2_antennanp ANTENNA_937 (.A(net1104));
 sg13g2_antennanp ANTENNA_938 (.A(net1104));
 sg13g2_antennanp ANTENNA_939 (.A(net1104));
 sg13g2_antennanp ANTENNA_940 (.A(net1104));
 sg13g2_antennanp ANTENNA_941 (.A(net1104));
 sg13g2_antennanp ANTENNA_942 (.A(net1104));
 sg13g2_antennanp ANTENNA_943 (.A(net1104));
 sg13g2_antennanp ANTENNA_944 (.A(net1104));
 sg13g2_antennanp ANTENNA_945 (.A(net1104));
 sg13g2_antennanp ANTENNA_946 (.A(net1104));
 sg13g2_antennanp ANTENNA_947 (.A(net1104));
 sg13g2_antennanp ANTENNA_948 (.A(net1104));
 sg13g2_antennanp ANTENNA_949 (.A(net1104));
 sg13g2_antennanp ANTENNA_950 (.A(net1104));
 sg13g2_antennanp ANTENNA_951 (.A(net1104));
 sg13g2_antennanp ANTENNA_952 (.A(net1104));
 sg13g2_antennanp ANTENNA_953 (.A(net1104));
 sg13g2_antennanp ANTENNA_954 (.A(net1104));
 sg13g2_antennanp ANTENNA_955 (.A(net1104));
 sg13g2_antennanp ANTENNA_956 (.A(_00928_));
 sg13g2_antennanp ANTENNA_957 (.A(_01057_));
 sg13g2_antennanp ANTENNA_958 (.A(_02823_));
 sg13g2_antennanp ANTENNA_959 (.A(_02823_));
 sg13g2_antennanp ANTENNA_960 (.A(_02823_));
 sg13g2_antennanp ANTENNA_961 (.A(_02823_));
 sg13g2_antennanp ANTENNA_962 (.A(_02823_));
 sg13g2_antennanp ANTENNA_963 (.A(_02823_));
 sg13g2_antennanp ANTENNA_964 (.A(_02823_));
 sg13g2_antennanp ANTENNA_965 (.A(_02823_));
 sg13g2_antennanp ANTENNA_966 (.A(_02823_));
 sg13g2_antennanp ANTENNA_967 (.A(_02831_));
 sg13g2_antennanp ANTENNA_968 (.A(_02831_));
 sg13g2_antennanp ANTENNA_969 (.A(_02831_));
 sg13g2_antennanp ANTENNA_970 (.A(_02831_));
 sg13g2_antennanp ANTENNA_971 (.A(_02831_));
 sg13g2_antennanp ANTENNA_972 (.A(_02831_));
 sg13g2_antennanp ANTENNA_973 (.A(_02831_));
 sg13g2_antennanp ANTENNA_974 (.A(_02831_));
 sg13g2_antennanp ANTENNA_975 (.A(_02831_));
 sg13g2_antennanp ANTENNA_976 (.A(_02835_));
 sg13g2_antennanp ANTENNA_977 (.A(_02835_));
 sg13g2_antennanp ANTENNA_978 (.A(_02835_));
 sg13g2_antennanp ANTENNA_979 (.A(_02835_));
 sg13g2_antennanp ANTENNA_980 (.A(_02835_));
 sg13g2_antennanp ANTENNA_981 (.A(_02835_));
 sg13g2_antennanp ANTENNA_982 (.A(_02835_));
 sg13g2_antennanp ANTENNA_983 (.A(_02835_));
 sg13g2_antennanp ANTENNA_984 (.A(_02835_));
 sg13g2_antennanp ANTENNA_985 (.A(_02990_));
 sg13g2_antennanp ANTENNA_986 (.A(_02990_));
 sg13g2_antennanp ANTENNA_987 (.A(_02990_));
 sg13g2_antennanp ANTENNA_988 (.A(_02990_));
 sg13g2_antennanp ANTENNA_989 (.A(_02990_));
 sg13g2_antennanp ANTENNA_990 (.A(_02990_));
 sg13g2_antennanp ANTENNA_991 (.A(_02990_));
 sg13g2_antennanp ANTENNA_992 (.A(_02990_));
 sg13g2_antennanp ANTENNA_993 (.A(_02990_));
 sg13g2_antennanp ANTENNA_994 (.A(_02990_));
 sg13g2_antennanp ANTENNA_995 (.A(_03019_));
 sg13g2_antennanp ANTENNA_996 (.A(_03019_));
 sg13g2_antennanp ANTENNA_997 (.A(_03019_));
 sg13g2_antennanp ANTENNA_998 (.A(_03865_));
 sg13g2_antennanp ANTENNA_999 (.A(_03865_));
 sg13g2_antennanp ANTENNA_1000 (.A(_03865_));
 sg13g2_antennanp ANTENNA_1001 (.A(_03865_));
 sg13g2_antennanp ANTENNA_1002 (.A(_03865_));
 sg13g2_antennanp ANTENNA_1003 (.A(_03865_));
 sg13g2_antennanp ANTENNA_1004 (.A(_04881_));
 sg13g2_antennanp ANTENNA_1005 (.A(_04881_));
 sg13g2_antennanp ANTENNA_1006 (.A(_04881_));
 sg13g2_antennanp ANTENNA_1007 (.A(_04943_));
 sg13g2_antennanp ANTENNA_1008 (.A(_04943_));
 sg13g2_antennanp ANTENNA_1009 (.A(_04943_));
 sg13g2_antennanp ANTENNA_1010 (.A(_04943_));
 sg13g2_antennanp ANTENNA_1011 (.A(_04943_));
 sg13g2_antennanp ANTENNA_1012 (.A(_04943_));
 sg13g2_antennanp ANTENNA_1013 (.A(_04943_));
 sg13g2_antennanp ANTENNA_1014 (.A(_05015_));
 sg13g2_antennanp ANTENNA_1015 (.A(_05189_));
 sg13g2_antennanp ANTENNA_1016 (.A(_05223_));
 sg13g2_antennanp ANTENNA_1017 (.A(_05238_));
 sg13g2_antennanp ANTENNA_1018 (.A(_05278_));
 sg13g2_antennanp ANTENNA_1019 (.A(_05279_));
 sg13g2_antennanp ANTENNA_1020 (.A(_05291_));
 sg13g2_antennanp ANTENNA_1021 (.A(_05306_));
 sg13g2_antennanp ANTENNA_1022 (.A(_05323_));
 sg13g2_antennanp ANTENNA_1023 (.A(_05333_));
 sg13g2_antennanp ANTENNA_1024 (.A(_05406_));
 sg13g2_antennanp ANTENNA_1025 (.A(_05406_));
 sg13g2_antennanp ANTENNA_1026 (.A(_05406_));
 sg13g2_antennanp ANTENNA_1027 (.A(_05478_));
 sg13g2_antennanp ANTENNA_1028 (.A(_05483_));
 sg13g2_antennanp ANTENNA_1029 (.A(_05545_));
 sg13g2_antennanp ANTENNA_1030 (.A(_05551_));
 sg13g2_antennanp ANTENNA_1031 (.A(_05693_));
 sg13g2_antennanp ANTENNA_1032 (.A(_05781_));
 sg13g2_antennanp ANTENNA_1033 (.A(_05797_));
 sg13g2_antennanp ANTENNA_1034 (.A(_05801_));
 sg13g2_antennanp ANTENNA_1035 (.A(_05801_));
 sg13g2_antennanp ANTENNA_1036 (.A(_05815_));
 sg13g2_antennanp ANTENNA_1037 (.A(_05818_));
 sg13g2_antennanp ANTENNA_1038 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1039 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1040 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1041 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1042 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1043 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1044 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1045 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1046 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1047 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1048 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1049 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1050 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1051 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1052 (.A(_06735_));
 sg13g2_antennanp ANTENNA_1053 (.A(_06735_));
 sg13g2_antennanp ANTENNA_1054 (.A(_06735_));
 sg13g2_antennanp ANTENNA_1055 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1056 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1057 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1058 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1059 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1060 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1061 (.A(_07611_));
 sg13g2_antennanp ANTENNA_1062 (.A(_07611_));
 sg13g2_antennanp ANTENNA_1063 (.A(_07611_));
 sg13g2_antennanp ANTENNA_1064 (.A(_07611_));
 sg13g2_antennanp ANTENNA_1065 (.A(_07756_));
 sg13g2_antennanp ANTENNA_1066 (.A(_07756_));
 sg13g2_antennanp ANTENNA_1067 (.A(_07756_));
 sg13g2_antennanp ANTENNA_1068 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1069 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1070 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1071 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1072 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1073 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1074 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1075 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1076 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1077 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1078 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1079 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1080 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1081 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1082 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1083 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1084 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1085 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1086 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1087 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1088 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1089 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1090 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1091 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1092 (.A(_08278_));
 sg13g2_antennanp ANTENNA_1093 (.A(_08278_));
 sg13g2_antennanp ANTENNA_1094 (.A(_08278_));
 sg13g2_antennanp ANTENNA_1095 (.A(_08278_));
 sg13g2_antennanp ANTENNA_1096 (.A(_08648_));
 sg13g2_antennanp ANTENNA_1097 (.A(_08648_));
 sg13g2_antennanp ANTENNA_1098 (.A(_08648_));
 sg13g2_antennanp ANTENNA_1099 (.A(_08648_));
 sg13g2_antennanp ANTENNA_1100 (.A(_08648_));
 sg13g2_antennanp ANTENNA_1101 (.A(_08648_));
 sg13g2_antennanp ANTENNA_1102 (.A(_08681_));
 sg13g2_antennanp ANTENNA_1103 (.A(_08681_));
 sg13g2_antennanp ANTENNA_1104 (.A(_08681_));
 sg13g2_antennanp ANTENNA_1105 (.A(_08681_));
 sg13g2_antennanp ANTENNA_1106 (.A(_08681_));
 sg13g2_antennanp ANTENNA_1107 (.A(_08681_));
 sg13g2_antennanp ANTENNA_1108 (.A(_08712_));
 sg13g2_antennanp ANTENNA_1109 (.A(_08769_));
 sg13g2_antennanp ANTENNA_1110 (.A(_08769_));
 sg13g2_antennanp ANTENNA_1111 (.A(_08769_));
 sg13g2_antennanp ANTENNA_1112 (.A(_08797_));
 sg13g2_antennanp ANTENNA_1113 (.A(_08797_));
 sg13g2_antennanp ANTENNA_1114 (.A(_08797_));
 sg13g2_antennanp ANTENNA_1115 (.A(_08797_));
 sg13g2_antennanp ANTENNA_1116 (.A(_08797_));
 sg13g2_antennanp ANTENNA_1117 (.A(_08817_));
 sg13g2_antennanp ANTENNA_1118 (.A(_08817_));
 sg13g2_antennanp ANTENNA_1119 (.A(_08817_));
 sg13g2_antennanp ANTENNA_1120 (.A(_08817_));
 sg13g2_antennanp ANTENNA_1121 (.A(_08817_));
 sg13g2_antennanp ANTENNA_1122 (.A(_08840_));
 sg13g2_antennanp ANTENNA_1123 (.A(_08855_));
 sg13g2_antennanp ANTENNA_1124 (.A(_08855_));
 sg13g2_antennanp ANTENNA_1125 (.A(_08855_));
 sg13g2_antennanp ANTENNA_1126 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1127 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1128 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1129 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1130 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1131 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1132 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1133 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1134 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1135 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1136 (.A(_08919_));
 sg13g2_antennanp ANTENNA_1137 (.A(_08944_));
 sg13g2_antennanp ANTENNA_1138 (.A(_08944_));
 sg13g2_antennanp ANTENNA_1139 (.A(_08944_));
 sg13g2_antennanp ANTENNA_1140 (.A(_08944_));
 sg13g2_antennanp ANTENNA_1141 (.A(_08944_));
 sg13g2_antennanp ANTENNA_1142 (.A(_08944_));
 sg13g2_antennanp ANTENNA_1143 (.A(_08964_));
 sg13g2_antennanp ANTENNA_1144 (.A(_08965_));
 sg13g2_antennanp ANTENNA_1145 (.A(_08965_));
 sg13g2_antennanp ANTENNA_1146 (.A(_08988_));
 sg13g2_antennanp ANTENNA_1147 (.A(_08988_));
 sg13g2_antennanp ANTENNA_1148 (.A(_08988_));
 sg13g2_antennanp ANTENNA_1149 (.A(_08997_));
 sg13g2_antennanp ANTENNA_1150 (.A(_09012_));
 sg13g2_antennanp ANTENNA_1151 (.A(_09012_));
 sg13g2_antennanp ANTENNA_1152 (.A(_09012_));
 sg13g2_antennanp ANTENNA_1153 (.A(_09012_));
 sg13g2_antennanp ANTENNA_1154 (.A(_09205_));
 sg13g2_antennanp ANTENNA_1155 (.A(_09205_));
 sg13g2_antennanp ANTENNA_1156 (.A(_09205_));
 sg13g2_antennanp ANTENNA_1157 (.A(_09205_));
 sg13g2_antennanp ANTENNA_1158 (.A(_09255_));
 sg13g2_antennanp ANTENNA_1159 (.A(_09255_));
 sg13g2_antennanp ANTENNA_1160 (.A(_09255_));
 sg13g2_antennanp ANTENNA_1161 (.A(_09255_));
 sg13g2_antennanp ANTENNA_1162 (.A(_09258_));
 sg13g2_antennanp ANTENNA_1163 (.A(_09258_));
 sg13g2_antennanp ANTENNA_1164 (.A(_09258_));
 sg13g2_antennanp ANTENNA_1165 (.A(_09258_));
 sg13g2_antennanp ANTENNA_1166 (.A(_09260_));
 sg13g2_antennanp ANTENNA_1167 (.A(_09266_));
 sg13g2_antennanp ANTENNA_1168 (.A(_09266_));
 sg13g2_antennanp ANTENNA_1169 (.A(_09266_));
 sg13g2_antennanp ANTENNA_1170 (.A(_09266_));
 sg13g2_antennanp ANTENNA_1171 (.A(_09294_));
 sg13g2_antennanp ANTENNA_1172 (.A(_09294_));
 sg13g2_antennanp ANTENNA_1173 (.A(_09294_));
 sg13g2_antennanp ANTENNA_1174 (.A(_09294_));
 sg13g2_antennanp ANTENNA_1175 (.A(_09294_));
 sg13g2_antennanp ANTENNA_1176 (.A(_09294_));
 sg13g2_antennanp ANTENNA_1177 (.A(_09294_));
 sg13g2_antennanp ANTENNA_1178 (.A(_09297_));
 sg13g2_antennanp ANTENNA_1179 (.A(_09297_));
 sg13g2_antennanp ANTENNA_1180 (.A(_09297_));
 sg13g2_antennanp ANTENNA_1181 (.A(_09297_));
 sg13g2_antennanp ANTENNA_1182 (.A(_09463_));
 sg13g2_antennanp ANTENNA_1183 (.A(_09488_));
 sg13g2_antennanp ANTENNA_1184 (.A(_09512_));
 sg13g2_antennanp ANTENNA_1185 (.A(_09517_));
 sg13g2_antennanp ANTENNA_1186 (.A(_09517_));
 sg13g2_antennanp ANTENNA_1187 (.A(_09517_));
 sg13g2_antennanp ANTENNA_1188 (.A(_09517_));
 sg13g2_antennanp ANTENNA_1189 (.A(_09517_));
 sg13g2_antennanp ANTENNA_1190 (.A(_09517_));
 sg13g2_antennanp ANTENNA_1191 (.A(_09517_));
 sg13g2_antennanp ANTENNA_1192 (.A(_09524_));
 sg13g2_antennanp ANTENNA_1193 (.A(_09524_));
 sg13g2_antennanp ANTENNA_1194 (.A(_09524_));
 sg13g2_antennanp ANTENNA_1195 (.A(_09544_));
 sg13g2_antennanp ANTENNA_1196 (.A(_09552_));
 sg13g2_antennanp ANTENNA_1197 (.A(_09639_));
 sg13g2_antennanp ANTENNA_1198 (.A(_09664_));
 sg13g2_antennanp ANTENNA_1199 (.A(_09685_));
 sg13g2_antennanp ANTENNA_1200 (.A(_09712_));
 sg13g2_antennanp ANTENNA_1201 (.A(_09727_));
 sg13g2_antennanp ANTENNA_1202 (.A(_09744_));
 sg13g2_antennanp ANTENNA_1203 (.A(_09744_));
 sg13g2_antennanp ANTENNA_1204 (.A(_09744_));
 sg13g2_antennanp ANTENNA_1205 (.A(_09744_));
 sg13g2_antennanp ANTENNA_1206 (.A(_09753_));
 sg13g2_antennanp ANTENNA_1207 (.A(_09775_));
 sg13g2_antennanp ANTENNA_1208 (.A(_09798_));
 sg13g2_antennanp ANTENNA_1209 (.A(_09954_));
 sg13g2_antennanp ANTENNA_1210 (.A(_09954_));
 sg13g2_antennanp ANTENNA_1211 (.A(_09954_));
 sg13g2_antennanp ANTENNA_1212 (.A(_10050_));
 sg13g2_antennanp ANTENNA_1213 (.A(_10050_));
 sg13g2_antennanp ANTENNA_1214 (.A(_10050_));
 sg13g2_antennanp ANTENNA_1215 (.A(_10050_));
 sg13g2_antennanp ANTENNA_1216 (.A(_10050_));
 sg13g2_antennanp ANTENNA_1217 (.A(_10050_));
 sg13g2_antennanp ANTENNA_1218 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1219 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1220 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1221 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1222 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1223 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1224 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1225 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1226 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1227 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1228 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1229 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1230 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1231 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1232 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1233 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1234 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1235 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1236 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1237 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1238 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1239 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1240 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1241 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1242 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1243 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1244 (.A(_10107_));
 sg13g2_antennanp ANTENNA_1245 (.A(_10107_));
 sg13g2_antennanp ANTENNA_1246 (.A(_10107_));
 sg13g2_antennanp ANTENNA_1247 (.A(_10107_));
 sg13g2_antennanp ANTENNA_1248 (.A(_10107_));
 sg13g2_antennanp ANTENNA_1249 (.A(_10107_));
 sg13g2_antennanp ANTENNA_1250 (.A(_10107_));
 sg13g2_antennanp ANTENNA_1251 (.A(_10107_));
 sg13g2_antennanp ANTENNA_1252 (.A(_10107_));
 sg13g2_antennanp ANTENNA_1253 (.A(_10107_));
 sg13g2_antennanp ANTENNA_1254 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1255 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1256 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1257 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1258 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1259 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1260 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1261 (.A(_10191_));
 sg13g2_antennanp ANTENNA_1262 (.A(_10191_));
 sg13g2_antennanp ANTENNA_1263 (.A(_10191_));
 sg13g2_antennanp ANTENNA_1264 (.A(_10191_));
 sg13g2_antennanp ANTENNA_1265 (.A(_10191_));
 sg13g2_antennanp ANTENNA_1266 (.A(_10191_));
 sg13g2_antennanp ANTENNA_1267 (.A(_10191_));
 sg13g2_antennanp ANTENNA_1268 (.A(_10191_));
 sg13g2_antennanp ANTENNA_1269 (.A(_10386_));
 sg13g2_antennanp ANTENNA_1270 (.A(_10386_));
 sg13g2_antennanp ANTENNA_1271 (.A(_10572_));
 sg13g2_antennanp ANTENNA_1272 (.A(_10572_));
 sg13g2_antennanp ANTENNA_1273 (.A(_10572_));
 sg13g2_antennanp ANTENNA_1274 (.A(_10572_));
 sg13g2_antennanp ANTENNA_1275 (.A(_10703_));
 sg13g2_antennanp ANTENNA_1276 (.A(_10703_));
 sg13g2_antennanp ANTENNA_1277 (.A(_10703_));
 sg13g2_antennanp ANTENNA_1278 (.A(_10889_));
 sg13g2_antennanp ANTENNA_1279 (.A(_10889_));
 sg13g2_antennanp ANTENNA_1280 (.A(_10889_));
 sg13g2_antennanp ANTENNA_1281 (.A(_11885_));
 sg13g2_antennanp ANTENNA_1282 (.A(_11885_));
 sg13g2_antennanp ANTENNA_1283 (.A(_11885_));
 sg13g2_antennanp ANTENNA_1284 (.A(_11970_));
 sg13g2_antennanp ANTENNA_1285 (.A(_11970_));
 sg13g2_antennanp ANTENNA_1286 (.A(_11970_));
 sg13g2_antennanp ANTENNA_1287 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1288 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1289 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1290 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1291 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1292 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1293 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1294 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1295 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1296 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1297 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1298 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1299 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1300 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1301 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1302 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1303 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1304 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1305 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1306 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1307 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1308 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1309 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1310 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1311 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1312 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1313 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1314 (.A(_12073_));
 sg13g2_antennanp ANTENNA_1315 (.A(_12073_));
 sg13g2_antennanp ANTENNA_1316 (.A(_12073_));
 sg13g2_antennanp ANTENNA_1317 (.A(_12073_));
 sg13g2_antennanp ANTENNA_1318 (.A(_12073_));
 sg13g2_antennanp ANTENNA_1319 (.A(_12073_));
 sg13g2_antennanp ANTENNA_1320 (.A(_12073_));
 sg13g2_antennanp ANTENNA_1321 (.A(_12073_));
 sg13g2_antennanp ANTENNA_1322 (.A(_12073_));
 sg13g2_antennanp ANTENNA_1323 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1324 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1325 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1326 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1327 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1328 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1329 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1330 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1331 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1332 (.A(_12133_));
 sg13g2_antennanp ANTENNA_1333 (.A(_12133_));
 sg13g2_antennanp ANTENNA_1334 (.A(_12133_));
 sg13g2_antennanp ANTENNA_1335 (.A(_12133_));
 sg13g2_antennanp ANTENNA_1336 (.A(_12133_));
 sg13g2_antennanp ANTENNA_1337 (.A(_12133_));
 sg13g2_antennanp ANTENNA_1338 (.A(_12133_));
 sg13g2_antennanp ANTENNA_1339 (.A(_12133_));
 sg13g2_antennanp ANTENNA_1340 (.A(_12133_));
 sg13g2_antennanp ANTENNA_1341 (.A(_12133_));
 sg13g2_antennanp ANTENNA_1342 (.A(_12156_));
 sg13g2_antennanp ANTENNA_1343 (.A(_12156_));
 sg13g2_antennanp ANTENNA_1344 (.A(_12156_));
 sg13g2_antennanp ANTENNA_1345 (.A(_12156_));
 sg13g2_antennanp ANTENNA_1346 (.A(_12156_));
 sg13g2_antennanp ANTENNA_1347 (.A(_12156_));
 sg13g2_antennanp ANTENNA_1348 (.A(_12156_));
 sg13g2_antennanp ANTENNA_1349 (.A(_12156_));
 sg13g2_antennanp ANTENNA_1350 (.A(_12156_));
 sg13g2_antennanp ANTENNA_1351 (.A(_12156_));
 sg13g2_antennanp ANTENNA_1352 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1353 (.A(r_reset));
 sg13g2_antennanp ANTENNA_1354 (.A(r_reset));
 sg13g2_antennanp ANTENNA_1355 (.A(r_reset));
 sg13g2_antennanp ANTENNA_1356 (.A(net1));
 sg13g2_antennanp ANTENNA_1357 (.A(net1));
 sg13g2_antennanp ANTENNA_1358 (.A(net1));
 sg13g2_antennanp ANTENNA_1359 (.A(net2));
 sg13g2_antennanp ANTENNA_1360 (.A(net2));
 sg13g2_antennanp ANTENNA_1361 (.A(net3));
 sg13g2_antennanp ANTENNA_1362 (.A(net3));
 sg13g2_antennanp ANTENNA_1363 (.A(net3));
 sg13g2_antennanp ANTENNA_1364 (.A(net11));
 sg13g2_antennanp ANTENNA_1365 (.A(net11));
 sg13g2_antennanp ANTENNA_1366 (.A(net11));
 sg13g2_antennanp ANTENNA_1367 (.A(net12));
 sg13g2_antennanp ANTENNA_1368 (.A(net12));
 sg13g2_antennanp ANTENNA_1369 (.A(net12));
 sg13g2_antennanp ANTENNA_1370 (.A(net13));
 sg13g2_antennanp ANTENNA_1371 (.A(net13));
 sg13g2_antennanp ANTENNA_1372 (.A(net13));
 sg13g2_antennanp ANTENNA_1373 (.A(net14));
 sg13g2_antennanp ANTENNA_1374 (.A(net14));
 sg13g2_antennanp ANTENNA_1375 (.A(net14));
 sg13g2_antennanp ANTENNA_1376 (.A(net19));
 sg13g2_antennanp ANTENNA_1377 (.A(net19));
 sg13g2_antennanp ANTENNA_1378 (.A(net19));
 sg13g2_antennanp ANTENNA_1379 (.A(net20));
 sg13g2_antennanp ANTENNA_1380 (.A(net20));
 sg13g2_antennanp ANTENNA_1381 (.A(net153));
 sg13g2_antennanp ANTENNA_1382 (.A(net153));
 sg13g2_antennanp ANTENNA_1383 (.A(net153));
 sg13g2_antennanp ANTENNA_1384 (.A(net153));
 sg13g2_antennanp ANTENNA_1385 (.A(net153));
 sg13g2_antennanp ANTENNA_1386 (.A(net153));
 sg13g2_antennanp ANTENNA_1387 (.A(net153));
 sg13g2_antennanp ANTENNA_1388 (.A(net153));
 sg13g2_antennanp ANTENNA_1389 (.A(net153));
 sg13g2_antennanp ANTENNA_1390 (.A(net153));
 sg13g2_antennanp ANTENNA_1391 (.A(net153));
 sg13g2_antennanp ANTENNA_1392 (.A(net153));
 sg13g2_antennanp ANTENNA_1393 (.A(net153));
 sg13g2_antennanp ANTENNA_1394 (.A(net153));
 sg13g2_antennanp ANTENNA_1395 (.A(net153));
 sg13g2_antennanp ANTENNA_1396 (.A(net153));
 sg13g2_antennanp ANTENNA_1397 (.A(net520));
 sg13g2_antennanp ANTENNA_1398 (.A(net520));
 sg13g2_antennanp ANTENNA_1399 (.A(net520));
 sg13g2_antennanp ANTENNA_1400 (.A(net520));
 sg13g2_antennanp ANTENNA_1401 (.A(net520));
 sg13g2_antennanp ANTENNA_1402 (.A(net520));
 sg13g2_antennanp ANTENNA_1403 (.A(net520));
 sg13g2_antennanp ANTENNA_1404 (.A(net520));
 sg13g2_antennanp ANTENNA_1405 (.A(net520));
 sg13g2_antennanp ANTENNA_1406 (.A(net520));
 sg13g2_antennanp ANTENNA_1407 (.A(net520));
 sg13g2_antennanp ANTENNA_1408 (.A(net520));
 sg13g2_antennanp ANTENNA_1409 (.A(net520));
 sg13g2_antennanp ANTENNA_1410 (.A(net520));
 sg13g2_antennanp ANTENNA_1411 (.A(net520));
 sg13g2_antennanp ANTENNA_1412 (.A(net520));
 sg13g2_antennanp ANTENNA_1413 (.A(net520));
 sg13g2_antennanp ANTENNA_1414 (.A(net520));
 sg13g2_antennanp ANTENNA_1415 (.A(net520));
 sg13g2_antennanp ANTENNA_1416 (.A(net520));
 sg13g2_antennanp ANTENNA_1417 (.A(net520));
 sg13g2_antennanp ANTENNA_1418 (.A(net520));
 sg13g2_antennanp ANTENNA_1419 (.A(net520));
 sg13g2_antennanp ANTENNA_1420 (.A(net520));
 sg13g2_antennanp ANTENNA_1421 (.A(net520));
 sg13g2_antennanp ANTENNA_1422 (.A(net520));
 sg13g2_antennanp ANTENNA_1423 (.A(net520));
 sg13g2_antennanp ANTENNA_1424 (.A(net520));
 sg13g2_antennanp ANTENNA_1425 (.A(net520));
 sg13g2_antennanp ANTENNA_1426 (.A(net520));
 sg13g2_antennanp ANTENNA_1427 (.A(net520));
 sg13g2_antennanp ANTENNA_1428 (.A(net538));
 sg13g2_antennanp ANTENNA_1429 (.A(net538));
 sg13g2_antennanp ANTENNA_1430 (.A(net538));
 sg13g2_antennanp ANTENNA_1431 (.A(net538));
 sg13g2_antennanp ANTENNA_1432 (.A(net538));
 sg13g2_antennanp ANTENNA_1433 (.A(net538));
 sg13g2_antennanp ANTENNA_1434 (.A(net538));
 sg13g2_antennanp ANTENNA_1435 (.A(net538));
 sg13g2_antennanp ANTENNA_1436 (.A(net596));
 sg13g2_antennanp ANTENNA_1437 (.A(net596));
 sg13g2_antennanp ANTENNA_1438 (.A(net596));
 sg13g2_antennanp ANTENNA_1439 (.A(net596));
 sg13g2_antennanp ANTENNA_1440 (.A(net596));
 sg13g2_antennanp ANTENNA_1441 (.A(net596));
 sg13g2_antennanp ANTENNA_1442 (.A(net596));
 sg13g2_antennanp ANTENNA_1443 (.A(net596));
 sg13g2_antennanp ANTENNA_1444 (.A(net618));
 sg13g2_antennanp ANTENNA_1445 (.A(net618));
 sg13g2_antennanp ANTENNA_1446 (.A(net618));
 sg13g2_antennanp ANTENNA_1447 (.A(net618));
 sg13g2_antennanp ANTENNA_1448 (.A(net618));
 sg13g2_antennanp ANTENNA_1449 (.A(net618));
 sg13g2_antennanp ANTENNA_1450 (.A(net618));
 sg13g2_antennanp ANTENNA_1451 (.A(net618));
 sg13g2_antennanp ANTENNA_1452 (.A(net618));
 sg13g2_antennanp ANTENNA_1453 (.A(net618));
 sg13g2_antennanp ANTENNA_1454 (.A(net618));
 sg13g2_antennanp ANTENNA_1455 (.A(net618));
 sg13g2_antennanp ANTENNA_1456 (.A(net618));
 sg13g2_antennanp ANTENNA_1457 (.A(net618));
 sg13g2_antennanp ANTENNA_1458 (.A(net618));
 sg13g2_antennanp ANTENNA_1459 (.A(net618));
 sg13g2_antennanp ANTENNA_1460 (.A(net618));
 sg13g2_antennanp ANTENNA_1461 (.A(net631));
 sg13g2_antennanp ANTENNA_1462 (.A(net631));
 sg13g2_antennanp ANTENNA_1463 (.A(net631));
 sg13g2_antennanp ANTENNA_1464 (.A(net631));
 sg13g2_antennanp ANTENNA_1465 (.A(net631));
 sg13g2_antennanp ANTENNA_1466 (.A(net631));
 sg13g2_antennanp ANTENNA_1467 (.A(net631));
 sg13g2_antennanp ANTENNA_1468 (.A(net631));
 sg13g2_antennanp ANTENNA_1469 (.A(net631));
 sg13g2_antennanp ANTENNA_1470 (.A(net632));
 sg13g2_antennanp ANTENNA_1471 (.A(net632));
 sg13g2_antennanp ANTENNA_1472 (.A(net632));
 sg13g2_antennanp ANTENNA_1473 (.A(net632));
 sg13g2_antennanp ANTENNA_1474 (.A(net632));
 sg13g2_antennanp ANTENNA_1475 (.A(net632));
 sg13g2_antennanp ANTENNA_1476 (.A(net632));
 sg13g2_antennanp ANTENNA_1477 (.A(net632));
 sg13g2_antennanp ANTENNA_1478 (.A(net632));
 sg13g2_antennanp ANTENNA_1479 (.A(net632));
 sg13g2_antennanp ANTENNA_1480 (.A(net632));
 sg13g2_antennanp ANTENNA_1481 (.A(net632));
 sg13g2_antennanp ANTENNA_1482 (.A(net632));
 sg13g2_antennanp ANTENNA_1483 (.A(net651));
 sg13g2_antennanp ANTENNA_1484 (.A(net651));
 sg13g2_antennanp ANTENNA_1485 (.A(net651));
 sg13g2_antennanp ANTENNA_1486 (.A(net651));
 sg13g2_antennanp ANTENNA_1487 (.A(net651));
 sg13g2_antennanp ANTENNA_1488 (.A(net651));
 sg13g2_antennanp ANTENNA_1489 (.A(net651));
 sg13g2_antennanp ANTENNA_1490 (.A(net651));
 sg13g2_antennanp ANTENNA_1491 (.A(net651));
 sg13g2_antennanp ANTENNA_1492 (.A(net651));
 sg13g2_antennanp ANTENNA_1493 (.A(net651));
 sg13g2_antennanp ANTENNA_1494 (.A(net651));
 sg13g2_antennanp ANTENNA_1495 (.A(net651));
 sg13g2_antennanp ANTENNA_1496 (.A(net651));
 sg13g2_antennanp ANTENNA_1497 (.A(net651));
 sg13g2_antennanp ANTENNA_1498 (.A(net651));
 sg13g2_antennanp ANTENNA_1499 (.A(net651));
 sg13g2_antennanp ANTENNA_1500 (.A(net651));
 sg13g2_antennanp ANTENNA_1501 (.A(net651));
 sg13g2_antennanp ANTENNA_1502 (.A(net651));
 sg13g2_antennanp ANTENNA_1503 (.A(net651));
 sg13g2_antennanp ANTENNA_1504 (.A(net651));
 sg13g2_antennanp ANTENNA_1505 (.A(net651));
 sg13g2_antennanp ANTENNA_1506 (.A(net651));
 sg13g2_antennanp ANTENNA_1507 (.A(net651));
 sg13g2_antennanp ANTENNA_1508 (.A(net651));
 sg13g2_antennanp ANTENNA_1509 (.A(net651));
 sg13g2_antennanp ANTENNA_1510 (.A(net651));
 sg13g2_antennanp ANTENNA_1511 (.A(net651));
 sg13g2_antennanp ANTENNA_1512 (.A(net651));
 sg13g2_antennanp ANTENNA_1513 (.A(net704));
 sg13g2_antennanp ANTENNA_1514 (.A(net704));
 sg13g2_antennanp ANTENNA_1515 (.A(net704));
 sg13g2_antennanp ANTENNA_1516 (.A(net704));
 sg13g2_antennanp ANTENNA_1517 (.A(net704));
 sg13g2_antennanp ANTENNA_1518 (.A(net704));
 sg13g2_antennanp ANTENNA_1519 (.A(net704));
 sg13g2_antennanp ANTENNA_1520 (.A(net704));
 sg13g2_antennanp ANTENNA_1521 (.A(net704));
 sg13g2_antennanp ANTENNA_1522 (.A(net860));
 sg13g2_antennanp ANTENNA_1523 (.A(net860));
 sg13g2_antennanp ANTENNA_1524 (.A(net860));
 sg13g2_antennanp ANTENNA_1525 (.A(net860));
 sg13g2_antennanp ANTENNA_1526 (.A(net860));
 sg13g2_antennanp ANTENNA_1527 (.A(net860));
 sg13g2_antennanp ANTENNA_1528 (.A(net860));
 sg13g2_antennanp ANTENNA_1529 (.A(net860));
 sg13g2_antennanp ANTENNA_1530 (.A(net860));
 sg13g2_antennanp ANTENNA_1531 (.A(net860));
 sg13g2_antennanp ANTENNA_1532 (.A(net860));
 sg13g2_antennanp ANTENNA_1533 (.A(net860));
 sg13g2_antennanp ANTENNA_1534 (.A(net860));
 sg13g2_antennanp ANTENNA_1535 (.A(net860));
 sg13g2_antennanp ANTENNA_1536 (.A(net860));
 sg13g2_antennanp ANTENNA_1537 (.A(net860));
 sg13g2_antennanp ANTENNA_1538 (.A(net860));
 sg13g2_antennanp ANTENNA_1539 (.A(net860));
 sg13g2_antennanp ANTENNA_1540 (.A(net860));
 sg13g2_antennanp ANTENNA_1541 (.A(net891));
 sg13g2_antennanp ANTENNA_1542 (.A(net891));
 sg13g2_antennanp ANTENNA_1543 (.A(net891));
 sg13g2_antennanp ANTENNA_1544 (.A(net891));
 sg13g2_antennanp ANTENNA_1545 (.A(net891));
 sg13g2_antennanp ANTENNA_1546 (.A(net891));
 sg13g2_antennanp ANTENNA_1547 (.A(net891));
 sg13g2_antennanp ANTENNA_1548 (.A(net891));
 sg13g2_antennanp ANTENNA_1549 (.A(net891));
 sg13g2_antennanp ANTENNA_1550 (.A(net959));
 sg13g2_antennanp ANTENNA_1551 (.A(net959));
 sg13g2_antennanp ANTENNA_1552 (.A(net959));
 sg13g2_antennanp ANTENNA_1553 (.A(net959));
 sg13g2_antennanp ANTENNA_1554 (.A(net959));
 sg13g2_antennanp ANTENNA_1555 (.A(net959));
 sg13g2_antennanp ANTENNA_1556 (.A(net959));
 sg13g2_antennanp ANTENNA_1557 (.A(net959));
 sg13g2_antennanp ANTENNA_1558 (.A(net959));
 sg13g2_antennanp ANTENNA_1559 (.A(net967));
 sg13g2_antennanp ANTENNA_1560 (.A(net967));
 sg13g2_antennanp ANTENNA_1561 (.A(net967));
 sg13g2_antennanp ANTENNA_1562 (.A(net967));
 sg13g2_antennanp ANTENNA_1563 (.A(net967));
 sg13g2_antennanp ANTENNA_1564 (.A(net967));
 sg13g2_antennanp ANTENNA_1565 (.A(net967));
 sg13g2_antennanp ANTENNA_1566 (.A(net967));
 sg13g2_antennanp ANTENNA_1567 (.A(net967));
 sg13g2_antennanp ANTENNA_1568 (.A(net969));
 sg13g2_antennanp ANTENNA_1569 (.A(net969));
 sg13g2_antennanp ANTENNA_1570 (.A(net969));
 sg13g2_antennanp ANTENNA_1571 (.A(net969));
 sg13g2_antennanp ANTENNA_1572 (.A(net969));
 sg13g2_antennanp ANTENNA_1573 (.A(net969));
 sg13g2_antennanp ANTENNA_1574 (.A(net969));
 sg13g2_antennanp ANTENNA_1575 (.A(net969));
 sg13g2_antennanp ANTENNA_1576 (.A(net969));
 sg13g2_antennanp ANTENNA_1577 (.A(net970));
 sg13g2_antennanp ANTENNA_1578 (.A(net970));
 sg13g2_antennanp ANTENNA_1579 (.A(net970));
 sg13g2_antennanp ANTENNA_1580 (.A(net970));
 sg13g2_antennanp ANTENNA_1581 (.A(net970));
 sg13g2_antennanp ANTENNA_1582 (.A(net970));
 sg13g2_antennanp ANTENNA_1583 (.A(net970));
 sg13g2_antennanp ANTENNA_1584 (.A(net970));
 sg13g2_antennanp ANTENNA_1585 (.A(net970));
 sg13g2_antennanp ANTENNA_1586 (.A(net970));
 sg13g2_antennanp ANTENNA_1587 (.A(net970));
 sg13g2_antennanp ANTENNA_1588 (.A(net970));
 sg13g2_antennanp ANTENNA_1589 (.A(net970));
 sg13g2_antennanp ANTENNA_1590 (.A(net970));
 sg13g2_antennanp ANTENNA_1591 (.A(net970));
 sg13g2_antennanp ANTENNA_1592 (.A(net972));
 sg13g2_antennanp ANTENNA_1593 (.A(net972));
 sg13g2_antennanp ANTENNA_1594 (.A(net972));
 sg13g2_antennanp ANTENNA_1595 (.A(net972));
 sg13g2_antennanp ANTENNA_1596 (.A(net972));
 sg13g2_antennanp ANTENNA_1597 (.A(net972));
 sg13g2_antennanp ANTENNA_1598 (.A(net972));
 sg13g2_antennanp ANTENNA_1599 (.A(net972));
 sg13g2_antennanp ANTENNA_1600 (.A(net972));
 sg13g2_antennanp ANTENNA_1601 (.A(net972));
 sg13g2_antennanp ANTENNA_1602 (.A(net972));
 sg13g2_antennanp ANTENNA_1603 (.A(net972));
 sg13g2_antennanp ANTENNA_1604 (.A(net972));
 sg13g2_antennanp ANTENNA_1605 (.A(net972));
 sg13g2_antennanp ANTENNA_1606 (.A(net972));
 sg13g2_antennanp ANTENNA_1607 (.A(net972));
 sg13g2_antennanp ANTENNA_1608 (.A(net972));
 sg13g2_antennanp ANTENNA_1609 (.A(net972));
 sg13g2_antennanp ANTENNA_1610 (.A(net972));
 sg13g2_antennanp ANTENNA_1611 (.A(net972));
 sg13g2_antennanp ANTENNA_1612 (.A(net972));
 sg13g2_antennanp ANTENNA_1613 (.A(net972));
 sg13g2_antennanp ANTENNA_1614 (.A(net972));
 sg13g2_antennanp ANTENNA_1615 (.A(net972));
 sg13g2_antennanp ANTENNA_1616 (.A(net972));
 sg13g2_antennanp ANTENNA_1617 (.A(net972));
 sg13g2_antennanp ANTENNA_1618 (.A(net972));
 sg13g2_antennanp ANTENNA_1619 (.A(net972));
 sg13g2_antennanp ANTENNA_1620 (.A(net972));
 sg13g2_antennanp ANTENNA_1621 (.A(net1000));
 sg13g2_antennanp ANTENNA_1622 (.A(net1000));
 sg13g2_antennanp ANTENNA_1623 (.A(net1000));
 sg13g2_antennanp ANTENNA_1624 (.A(net1000));
 sg13g2_antennanp ANTENNA_1625 (.A(net1000));
 sg13g2_antennanp ANTENNA_1626 (.A(net1000));
 sg13g2_antennanp ANTENNA_1627 (.A(net1000));
 sg13g2_antennanp ANTENNA_1628 (.A(net1000));
 sg13g2_antennanp ANTENNA_1629 (.A(net1043));
 sg13g2_antennanp ANTENNA_1630 (.A(net1043));
 sg13g2_antennanp ANTENNA_1631 (.A(net1043));
 sg13g2_antennanp ANTENNA_1632 (.A(net1043));
 sg13g2_antennanp ANTENNA_1633 (.A(net1043));
 sg13g2_antennanp ANTENNA_1634 (.A(net1043));
 sg13g2_antennanp ANTENNA_1635 (.A(net1043));
 sg13g2_antennanp ANTENNA_1636 (.A(net1043));
 sg13g2_antennanp ANTENNA_1637 (.A(net1043));
 sg13g2_antennanp ANTENNA_1638 (.A(net1043));
 sg13g2_antennanp ANTENNA_1639 (.A(net1043));
 sg13g2_antennanp ANTENNA_1640 (.A(net1043));
 sg13g2_antennanp ANTENNA_1641 (.A(net1072));
 sg13g2_antennanp ANTENNA_1642 (.A(net1072));
 sg13g2_antennanp ANTENNA_1643 (.A(net1072));
 sg13g2_antennanp ANTENNA_1644 (.A(net1072));
 sg13g2_antennanp ANTENNA_1645 (.A(net1072));
 sg13g2_antennanp ANTENNA_1646 (.A(net1072));
 sg13g2_antennanp ANTENNA_1647 (.A(net1072));
 sg13g2_antennanp ANTENNA_1648 (.A(net1072));
 sg13g2_antennanp ANTENNA_1649 (.A(net1072));
 sg13g2_antennanp ANTENNA_1650 (.A(net1104));
 sg13g2_antennanp ANTENNA_1651 (.A(net1104));
 sg13g2_antennanp ANTENNA_1652 (.A(net1104));
 sg13g2_antennanp ANTENNA_1653 (.A(net1104));
 sg13g2_antennanp ANTENNA_1654 (.A(net1104));
 sg13g2_antennanp ANTENNA_1655 (.A(net1104));
 sg13g2_antennanp ANTENNA_1656 (.A(net1104));
 sg13g2_antennanp ANTENNA_1657 (.A(net1104));
 sg13g2_antennanp ANTENNA_1658 (.A(net1104));
 sg13g2_antennanp ANTENNA_1659 (.A(net1104));
 sg13g2_antennanp ANTENNA_1660 (.A(net1104));
 sg13g2_antennanp ANTENNA_1661 (.A(_00928_));
 sg13g2_antennanp ANTENNA_1662 (.A(_01057_));
 sg13g2_antennanp ANTENNA_1663 (.A(_02823_));
 sg13g2_antennanp ANTENNA_1664 (.A(_02823_));
 sg13g2_antennanp ANTENNA_1665 (.A(_02823_));
 sg13g2_antennanp ANTENNA_1666 (.A(_02823_));
 sg13g2_antennanp ANTENNA_1667 (.A(_02823_));
 sg13g2_antennanp ANTENNA_1668 (.A(_02823_));
 sg13g2_antennanp ANTENNA_1669 (.A(_02823_));
 sg13g2_antennanp ANTENNA_1670 (.A(_02823_));
 sg13g2_antennanp ANTENNA_1671 (.A(_02823_));
 sg13g2_antennanp ANTENNA_1672 (.A(_02831_));
 sg13g2_antennanp ANTENNA_1673 (.A(_02831_));
 sg13g2_antennanp ANTENNA_1674 (.A(_02831_));
 sg13g2_antennanp ANTENNA_1675 (.A(_02831_));
 sg13g2_antennanp ANTENNA_1676 (.A(_02831_));
 sg13g2_antennanp ANTENNA_1677 (.A(_02831_));
 sg13g2_antennanp ANTENNA_1678 (.A(_02831_));
 sg13g2_antennanp ANTENNA_1679 (.A(_02831_));
 sg13g2_antennanp ANTENNA_1680 (.A(_02831_));
 sg13g2_antennanp ANTENNA_1681 (.A(_02835_));
 sg13g2_antennanp ANTENNA_1682 (.A(_02835_));
 sg13g2_antennanp ANTENNA_1683 (.A(_02835_));
 sg13g2_antennanp ANTENNA_1684 (.A(_02835_));
 sg13g2_antennanp ANTENNA_1685 (.A(_02835_));
 sg13g2_antennanp ANTENNA_1686 (.A(_02835_));
 sg13g2_antennanp ANTENNA_1687 (.A(_02835_));
 sg13g2_antennanp ANTENNA_1688 (.A(_02835_));
 sg13g2_antennanp ANTENNA_1689 (.A(_02835_));
 sg13g2_antennanp ANTENNA_1690 (.A(_02990_));
 sg13g2_antennanp ANTENNA_1691 (.A(_02990_));
 sg13g2_antennanp ANTENNA_1692 (.A(_02990_));
 sg13g2_antennanp ANTENNA_1693 (.A(_02990_));
 sg13g2_antennanp ANTENNA_1694 (.A(_02990_));
 sg13g2_antennanp ANTENNA_1695 (.A(_02990_));
 sg13g2_antennanp ANTENNA_1696 (.A(_02990_));
 sg13g2_antennanp ANTENNA_1697 (.A(_02990_));
 sg13g2_antennanp ANTENNA_1698 (.A(_02990_));
 sg13g2_antennanp ANTENNA_1699 (.A(_02990_));
 sg13g2_antennanp ANTENNA_1700 (.A(_03019_));
 sg13g2_antennanp ANTENNA_1701 (.A(_03019_));
 sg13g2_antennanp ANTENNA_1702 (.A(_03019_));
 sg13g2_antennanp ANTENNA_1703 (.A(_03865_));
 sg13g2_antennanp ANTENNA_1704 (.A(_03865_));
 sg13g2_antennanp ANTENNA_1705 (.A(_03865_));
 sg13g2_antennanp ANTENNA_1706 (.A(_03865_));
 sg13g2_antennanp ANTENNA_1707 (.A(_04881_));
 sg13g2_antennanp ANTENNA_1708 (.A(_04881_));
 sg13g2_antennanp ANTENNA_1709 (.A(_04881_));
 sg13g2_antennanp ANTENNA_1710 (.A(_04881_));
 sg13g2_antennanp ANTENNA_1711 (.A(_04881_));
 sg13g2_antennanp ANTENNA_1712 (.A(_05015_));
 sg13g2_antennanp ANTENNA_1713 (.A(_05223_));
 sg13g2_antennanp ANTENNA_1714 (.A(_05238_));
 sg13g2_antennanp ANTENNA_1715 (.A(_05254_));
 sg13g2_antennanp ANTENNA_1716 (.A(_05278_));
 sg13g2_antennanp ANTENNA_1717 (.A(_05291_));
 sg13g2_antennanp ANTENNA_1718 (.A(_05306_));
 sg13g2_antennanp ANTENNA_1719 (.A(_05323_));
 sg13g2_antennanp ANTENNA_1720 (.A(_05333_));
 sg13g2_antennanp ANTENNA_1721 (.A(_05406_));
 sg13g2_antennanp ANTENNA_1722 (.A(_05406_));
 sg13g2_antennanp ANTENNA_1723 (.A(_05406_));
 sg13g2_antennanp ANTENNA_1724 (.A(_05478_));
 sg13g2_antennanp ANTENNA_1725 (.A(_05478_));
 sg13g2_antennanp ANTENNA_1726 (.A(_05483_));
 sg13g2_antennanp ANTENNA_1727 (.A(_05545_));
 sg13g2_antennanp ANTENNA_1728 (.A(_05551_));
 sg13g2_antennanp ANTENNA_1729 (.A(_05781_));
 sg13g2_antennanp ANTENNA_1730 (.A(_05797_));
 sg13g2_antennanp ANTENNA_1731 (.A(_05801_));
 sg13g2_antennanp ANTENNA_1732 (.A(_05801_));
 sg13g2_antennanp ANTENNA_1733 (.A(_05801_));
 sg13g2_antennanp ANTENNA_1734 (.A(_05801_));
 sg13g2_antennanp ANTENNA_1735 (.A(_05815_));
 sg13g2_antennanp ANTENNA_1736 (.A(_05818_));
 sg13g2_antennanp ANTENNA_1737 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1738 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1739 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1740 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1741 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1742 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1743 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1744 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1745 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1746 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1747 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1748 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1749 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1750 (.A(_06734_));
 sg13g2_antennanp ANTENNA_1751 (.A(_06735_));
 sg13g2_antennanp ANTENNA_1752 (.A(_06735_));
 sg13g2_antennanp ANTENNA_1753 (.A(_06735_));
 sg13g2_antennanp ANTENNA_1754 (.A(_06735_));
 sg13g2_antennanp ANTENNA_1755 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1756 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1757 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1758 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1759 (.A(_07611_));
 sg13g2_antennanp ANTENNA_1760 (.A(_07611_));
 sg13g2_antennanp ANTENNA_1761 (.A(_07611_));
 sg13g2_antennanp ANTENNA_1762 (.A(_07611_));
 sg13g2_antennanp ANTENNA_1763 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1764 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1765 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1766 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1767 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1768 (.A(_08265_));
 sg13g2_antennanp ANTENNA_1769 (.A(_08278_));
 sg13g2_antennanp ANTENNA_1770 (.A(_08278_));
 sg13g2_antennanp ANTENNA_1771 (.A(_08278_));
 sg13g2_antennanp ANTENNA_1772 (.A(_08278_));
 sg13g2_antennanp ANTENNA_1773 (.A(_08648_));
 sg13g2_antennanp ANTENNA_1774 (.A(_08648_));
 sg13g2_antennanp ANTENNA_1775 (.A(_08648_));
 sg13g2_antennanp ANTENNA_1776 (.A(_08648_));
 sg13g2_antennanp ANTENNA_1777 (.A(_08648_));
 sg13g2_antennanp ANTENNA_1778 (.A(_08648_));
 sg13g2_antennanp ANTENNA_1779 (.A(_08681_));
 sg13g2_antennanp ANTENNA_1780 (.A(_08681_));
 sg13g2_antennanp ANTENNA_1781 (.A(_08681_));
 sg13g2_antennanp ANTENNA_1782 (.A(_08681_));
 sg13g2_antennanp ANTENNA_1783 (.A(_08712_));
 sg13g2_antennanp ANTENNA_1784 (.A(_08758_));
 sg13g2_antennanp ANTENNA_1785 (.A(_08758_));
 sg13g2_antennanp ANTENNA_1786 (.A(_08758_));
 sg13g2_antennanp ANTENNA_1787 (.A(_08758_));
 sg13g2_antennanp ANTENNA_1788 (.A(_08758_));
 sg13g2_antennanp ANTENNA_1789 (.A(_08758_));
 sg13g2_antennanp ANTENNA_1790 (.A(_08758_));
 sg13g2_antennanp ANTENNA_1791 (.A(_08758_));
 sg13g2_antennanp ANTENNA_1792 (.A(_08758_));
 sg13g2_antennanp ANTENNA_1793 (.A(_08758_));
 sg13g2_antennanp ANTENNA_1794 (.A(_08769_));
 sg13g2_antennanp ANTENNA_1795 (.A(_08769_));
 sg13g2_antennanp ANTENNA_1796 (.A(_08769_));
 sg13g2_antennanp ANTENNA_1797 (.A(_08797_));
 sg13g2_antennanp ANTENNA_1798 (.A(_08797_));
 sg13g2_antennanp ANTENNA_1799 (.A(_08797_));
 sg13g2_antennanp ANTENNA_1800 (.A(_08797_));
 sg13g2_antennanp ANTENNA_1801 (.A(_08797_));
 sg13g2_antennanp ANTENNA_1802 (.A(_08817_));
 sg13g2_antennanp ANTENNA_1803 (.A(_08817_));
 sg13g2_antennanp ANTENNA_1804 (.A(_08817_));
 sg13g2_antennanp ANTENNA_1805 (.A(_08817_));
 sg13g2_antennanp ANTENNA_1806 (.A(_08817_));
 sg13g2_antennanp ANTENNA_1807 (.A(_08840_));
 sg13g2_antennanp ANTENNA_1808 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1809 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1810 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1811 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1812 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1813 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1814 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1815 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1816 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1817 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1818 (.A(_08879_));
 sg13g2_antennanp ANTENNA_1819 (.A(_08919_));
 sg13g2_antennanp ANTENNA_1820 (.A(_08944_));
 sg13g2_antennanp ANTENNA_1821 (.A(_08944_));
 sg13g2_antennanp ANTENNA_1822 (.A(_08944_));
 sg13g2_antennanp ANTENNA_1823 (.A(_08964_));
 sg13g2_antennanp ANTENNA_1824 (.A(_08965_));
 sg13g2_antennanp ANTENNA_1825 (.A(_08965_));
 sg13g2_antennanp ANTENNA_1826 (.A(_08988_));
 sg13g2_antennanp ANTENNA_1827 (.A(_08988_));
 sg13g2_antennanp ANTENNA_1828 (.A(_08988_));
 sg13g2_antennanp ANTENNA_1829 (.A(_08997_));
 sg13g2_antennanp ANTENNA_1830 (.A(_09012_));
 sg13g2_antennanp ANTENNA_1831 (.A(_09012_));
 sg13g2_antennanp ANTENNA_1832 (.A(_09012_));
 sg13g2_antennanp ANTENNA_1833 (.A(_09012_));
 sg13g2_antennanp ANTENNA_1834 (.A(_09205_));
 sg13g2_antennanp ANTENNA_1835 (.A(_09205_));
 sg13g2_antennanp ANTENNA_1836 (.A(_09205_));
 sg13g2_antennanp ANTENNA_1837 (.A(_09205_));
 sg13g2_antennanp ANTENNA_1838 (.A(_09255_));
 sg13g2_antennanp ANTENNA_1839 (.A(_09255_));
 sg13g2_antennanp ANTENNA_1840 (.A(_09255_));
 sg13g2_antennanp ANTENNA_1841 (.A(_09255_));
 sg13g2_antennanp ANTENNA_1842 (.A(_09258_));
 sg13g2_antennanp ANTENNA_1843 (.A(_09258_));
 sg13g2_antennanp ANTENNA_1844 (.A(_09258_));
 sg13g2_antennanp ANTENNA_1845 (.A(_09258_));
 sg13g2_antennanp ANTENNA_1846 (.A(_09260_));
 sg13g2_antennanp ANTENNA_1847 (.A(_09266_));
 sg13g2_antennanp ANTENNA_1848 (.A(_09266_));
 sg13g2_antennanp ANTENNA_1849 (.A(_09266_));
 sg13g2_antennanp ANTENNA_1850 (.A(_09266_));
 sg13g2_antennanp ANTENNA_1851 (.A(_09294_));
 sg13g2_antennanp ANTENNA_1852 (.A(_09294_));
 sg13g2_antennanp ANTENNA_1853 (.A(_09294_));
 sg13g2_antennanp ANTENNA_1854 (.A(_09294_));
 sg13g2_antennanp ANTENNA_1855 (.A(_09297_));
 sg13g2_antennanp ANTENNA_1856 (.A(_09297_));
 sg13g2_antennanp ANTENNA_1857 (.A(_09297_));
 sg13g2_antennanp ANTENNA_1858 (.A(_09297_));
 sg13g2_antennanp ANTENNA_1859 (.A(_09463_));
 sg13g2_antennanp ANTENNA_1860 (.A(_09488_));
 sg13g2_antennanp ANTENNA_1861 (.A(_09512_));
 sg13g2_antennanp ANTENNA_1862 (.A(_09524_));
 sg13g2_antennanp ANTENNA_1863 (.A(_09524_));
 sg13g2_antennanp ANTENNA_1864 (.A(_09524_));
 sg13g2_antennanp ANTENNA_1865 (.A(_09544_));
 sg13g2_antennanp ANTENNA_1866 (.A(_09552_));
 sg13g2_antennanp ANTENNA_1867 (.A(_09639_));
 sg13g2_antennanp ANTENNA_1868 (.A(_09664_));
 sg13g2_antennanp ANTENNA_1869 (.A(_09685_));
 sg13g2_antennanp ANTENNA_1870 (.A(_09712_));
 sg13g2_antennanp ANTENNA_1871 (.A(_09727_));
 sg13g2_antennanp ANTENNA_1872 (.A(_09744_));
 sg13g2_antennanp ANTENNA_1873 (.A(_09744_));
 sg13g2_antennanp ANTENNA_1874 (.A(_09744_));
 sg13g2_antennanp ANTENNA_1875 (.A(_09744_));
 sg13g2_antennanp ANTENNA_1876 (.A(_09753_));
 sg13g2_antennanp ANTENNA_1877 (.A(_09798_));
 sg13g2_antennanp ANTENNA_1878 (.A(_09954_));
 sg13g2_antennanp ANTENNA_1879 (.A(_09954_));
 sg13g2_antennanp ANTENNA_1880 (.A(_09954_));
 sg13g2_antennanp ANTENNA_1881 (.A(_09954_));
 sg13g2_antennanp ANTENNA_1882 (.A(_09954_));
 sg13g2_antennanp ANTENNA_1883 (.A(_09954_));
 sg13g2_antennanp ANTENNA_1884 (.A(_10050_));
 sg13g2_antennanp ANTENNA_1885 (.A(_10050_));
 sg13g2_antennanp ANTENNA_1886 (.A(_10050_));
 sg13g2_antennanp ANTENNA_1887 (.A(_10050_));
 sg13g2_antennanp ANTENNA_1888 (.A(_10050_));
 sg13g2_antennanp ANTENNA_1889 (.A(_10050_));
 sg13g2_antennanp ANTENNA_1890 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1891 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1892 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1893 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1894 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1895 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1896 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1897 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1898 (.A(_10054_));
 sg13g2_antennanp ANTENNA_1899 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1900 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1901 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1902 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1903 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1904 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1905 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1906 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1907 (.A(_10057_));
 sg13g2_antennanp ANTENNA_1908 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1909 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1910 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1911 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1912 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1913 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1914 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1915 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1916 (.A(_10107_));
 sg13g2_antennanp ANTENNA_1917 (.A(_10107_));
 sg13g2_antennanp ANTENNA_1918 (.A(_10107_));
 sg13g2_antennanp ANTENNA_1919 (.A(_10110_));
 sg13g2_antennanp ANTENNA_1920 (.A(_10110_));
 sg13g2_antennanp ANTENNA_1921 (.A(_10110_));
 sg13g2_antennanp ANTENNA_1922 (.A(_10110_));
 sg13g2_antennanp ANTENNA_1923 (.A(_10110_));
 sg13g2_antennanp ANTENNA_1924 (.A(_10110_));
 sg13g2_antennanp ANTENNA_1925 (.A(_10110_));
 sg13g2_antennanp ANTENNA_1926 (.A(_10110_));
 sg13g2_antennanp ANTENNA_1927 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1928 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1929 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1930 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1931 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1932 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1933 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1934 (.A(_10181_));
 sg13g2_antennanp ANTENNA_1935 (.A(_10386_));
 sg13g2_antennanp ANTENNA_1936 (.A(_10386_));
 sg13g2_antennanp ANTENNA_1937 (.A(_10572_));
 sg13g2_antennanp ANTENNA_1938 (.A(_10572_));
 sg13g2_antennanp ANTENNA_1939 (.A(_10572_));
 sg13g2_antennanp ANTENNA_1940 (.A(_10572_));
 sg13g2_antennanp ANTENNA_1941 (.A(_10703_));
 sg13g2_antennanp ANTENNA_1942 (.A(_10703_));
 sg13g2_antennanp ANTENNA_1943 (.A(_10703_));
 sg13g2_antennanp ANTENNA_1944 (.A(_10889_));
 sg13g2_antennanp ANTENNA_1945 (.A(_10889_));
 sg13g2_antennanp ANTENNA_1946 (.A(_10889_));
 sg13g2_antennanp ANTENNA_1947 (.A(_11885_));
 sg13g2_antennanp ANTENNA_1948 (.A(_11885_));
 sg13g2_antennanp ANTENNA_1949 (.A(_11885_));
 sg13g2_antennanp ANTENNA_1950 (.A(_11970_));
 sg13g2_antennanp ANTENNA_1951 (.A(_11970_));
 sg13g2_antennanp ANTENNA_1952 (.A(_11970_));
 sg13g2_antennanp ANTENNA_1953 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1954 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1955 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1956 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1957 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1958 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1959 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1960 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1961 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1962 (.A(_12023_));
 sg13g2_antennanp ANTENNA_1963 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1964 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1965 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1966 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1967 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1968 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1969 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1970 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1971 (.A(_12046_));
 sg13g2_antennanp ANTENNA_1972 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1973 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1974 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1975 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1976 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1977 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1978 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1979 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1980 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1981 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1982 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1983 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1984 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1985 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1986 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1987 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1988 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1989 (.A(_12063_));
 sg13g2_antennanp ANTENNA_1990 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1991 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1992 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1993 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1994 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1995 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1996 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1997 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1998 (.A(_12096_));
 sg13g2_antennanp ANTENNA_1999 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2000 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2001 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2002 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2003 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2004 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2005 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2006 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2007 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2008 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2009 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2010 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2011 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2012 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2013 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2014 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2015 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2016 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2017 (.A(_12156_));
 sg13g2_antennanp ANTENNA_2018 (.A(_12156_));
 sg13g2_antennanp ANTENNA_2019 (.A(_12156_));
 sg13g2_antennanp ANTENNA_2020 (.A(_12156_));
 sg13g2_antennanp ANTENNA_2021 (.A(_12156_));
 sg13g2_antennanp ANTENNA_2022 (.A(_12156_));
 sg13g2_antennanp ANTENNA_2023 (.A(_12156_));
 sg13g2_antennanp ANTENNA_2024 (.A(_12156_));
 sg13g2_antennanp ANTENNA_2025 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2026 (.A(r_reset));
 sg13g2_antennanp ANTENNA_2027 (.A(r_reset));
 sg13g2_antennanp ANTENNA_2028 (.A(r_reset));
 sg13g2_antennanp ANTENNA_2029 (.A(net1));
 sg13g2_antennanp ANTENNA_2030 (.A(net1));
 sg13g2_antennanp ANTENNA_2031 (.A(net1));
 sg13g2_antennanp ANTENNA_2032 (.A(net2));
 sg13g2_antennanp ANTENNA_2033 (.A(net2));
 sg13g2_antennanp ANTENNA_2034 (.A(net11));
 sg13g2_antennanp ANTENNA_2035 (.A(net11));
 sg13g2_antennanp ANTENNA_2036 (.A(net11));
 sg13g2_antennanp ANTENNA_2037 (.A(net12));
 sg13g2_antennanp ANTENNA_2038 (.A(net12));
 sg13g2_antennanp ANTENNA_2039 (.A(net12));
 sg13g2_antennanp ANTENNA_2040 (.A(net13));
 sg13g2_antennanp ANTENNA_2041 (.A(net13));
 sg13g2_antennanp ANTENNA_2042 (.A(net13));
 sg13g2_antennanp ANTENNA_2043 (.A(net14));
 sg13g2_antennanp ANTENNA_2044 (.A(net14));
 sg13g2_antennanp ANTENNA_2045 (.A(net14));
 sg13g2_antennanp ANTENNA_2046 (.A(net19));
 sg13g2_antennanp ANTENNA_2047 (.A(net19));
 sg13g2_antennanp ANTENNA_2048 (.A(net20));
 sg13g2_antennanp ANTENNA_2049 (.A(net20));
 sg13g2_antennanp ANTENNA_2050 (.A(net596));
 sg13g2_antennanp ANTENNA_2051 (.A(net596));
 sg13g2_antennanp ANTENNA_2052 (.A(net596));
 sg13g2_antennanp ANTENNA_2053 (.A(net596));
 sg13g2_antennanp ANTENNA_2054 (.A(net596));
 sg13g2_antennanp ANTENNA_2055 (.A(net596));
 sg13g2_antennanp ANTENNA_2056 (.A(net596));
 sg13g2_antennanp ANTENNA_2057 (.A(net596));
 sg13g2_antennanp ANTENNA_2058 (.A(net596));
 sg13g2_antennanp ANTENNA_2059 (.A(net618));
 sg13g2_antennanp ANTENNA_2060 (.A(net618));
 sg13g2_antennanp ANTENNA_2061 (.A(net618));
 sg13g2_antennanp ANTENNA_2062 (.A(net618));
 sg13g2_antennanp ANTENNA_2063 (.A(net618));
 sg13g2_antennanp ANTENNA_2064 (.A(net618));
 sg13g2_antennanp ANTENNA_2065 (.A(net618));
 sg13g2_antennanp ANTENNA_2066 (.A(net618));
 sg13g2_antennanp ANTENNA_2067 (.A(net618));
 sg13g2_antennanp ANTENNA_2068 (.A(net618));
 sg13g2_antennanp ANTENNA_2069 (.A(net618));
 sg13g2_antennanp ANTENNA_2070 (.A(net618));
 sg13g2_antennanp ANTENNA_2071 (.A(net631));
 sg13g2_antennanp ANTENNA_2072 (.A(net631));
 sg13g2_antennanp ANTENNA_2073 (.A(net631));
 sg13g2_antennanp ANTENNA_2074 (.A(net631));
 sg13g2_antennanp ANTENNA_2075 (.A(net631));
 sg13g2_antennanp ANTENNA_2076 (.A(net631));
 sg13g2_antennanp ANTENNA_2077 (.A(net631));
 sg13g2_antennanp ANTENNA_2078 (.A(net631));
 sg13g2_antennanp ANTENNA_2079 (.A(net651));
 sg13g2_antennanp ANTENNA_2080 (.A(net651));
 sg13g2_antennanp ANTENNA_2081 (.A(net651));
 sg13g2_antennanp ANTENNA_2082 (.A(net651));
 sg13g2_antennanp ANTENNA_2083 (.A(net651));
 sg13g2_antennanp ANTENNA_2084 (.A(net651));
 sg13g2_antennanp ANTENNA_2085 (.A(net651));
 sg13g2_antennanp ANTENNA_2086 (.A(net651));
 sg13g2_antennanp ANTENNA_2087 (.A(net651));
 sg13g2_antennanp ANTENNA_2088 (.A(net651));
 sg13g2_antennanp ANTENNA_2089 (.A(net651));
 sg13g2_antennanp ANTENNA_2090 (.A(net651));
 sg13g2_antennanp ANTENNA_2091 (.A(net651));
 sg13g2_antennanp ANTENNA_2092 (.A(net651));
 sg13g2_antennanp ANTENNA_2093 (.A(net651));
 sg13g2_antennanp ANTENNA_2094 (.A(net651));
 sg13g2_antennanp ANTENNA_2095 (.A(net651));
 sg13g2_antennanp ANTENNA_2096 (.A(net651));
 sg13g2_antennanp ANTENNA_2097 (.A(net651));
 sg13g2_antennanp ANTENNA_2098 (.A(net651));
 sg13g2_antennanp ANTENNA_2099 (.A(net651));
 sg13g2_antennanp ANTENNA_2100 (.A(net651));
 sg13g2_antennanp ANTENNA_2101 (.A(net704));
 sg13g2_antennanp ANTENNA_2102 (.A(net704));
 sg13g2_antennanp ANTENNA_2103 (.A(net704));
 sg13g2_antennanp ANTENNA_2104 (.A(net704));
 sg13g2_antennanp ANTENNA_2105 (.A(net704));
 sg13g2_antennanp ANTENNA_2106 (.A(net704));
 sg13g2_antennanp ANTENNA_2107 (.A(net704));
 sg13g2_antennanp ANTENNA_2108 (.A(net704));
 sg13g2_antennanp ANTENNA_2109 (.A(net704));
 sg13g2_antennanp ANTENNA_2110 (.A(net860));
 sg13g2_antennanp ANTENNA_2111 (.A(net860));
 sg13g2_antennanp ANTENNA_2112 (.A(net860));
 sg13g2_antennanp ANTENNA_2113 (.A(net860));
 sg13g2_antennanp ANTENNA_2114 (.A(net860));
 sg13g2_antennanp ANTENNA_2115 (.A(net860));
 sg13g2_antennanp ANTENNA_2116 (.A(net860));
 sg13g2_antennanp ANTENNA_2117 (.A(net860));
 sg13g2_antennanp ANTENNA_2118 (.A(net860));
 sg13g2_antennanp ANTENNA_2119 (.A(net891));
 sg13g2_antennanp ANTENNA_2120 (.A(net891));
 sg13g2_antennanp ANTENNA_2121 (.A(net891));
 sg13g2_antennanp ANTENNA_2122 (.A(net891));
 sg13g2_antennanp ANTENNA_2123 (.A(net891));
 sg13g2_antennanp ANTENNA_2124 (.A(net891));
 sg13g2_antennanp ANTENNA_2125 (.A(net891));
 sg13g2_antennanp ANTENNA_2126 (.A(net891));
 sg13g2_antennanp ANTENNA_2127 (.A(net891));
 sg13g2_antennanp ANTENNA_2128 (.A(net959));
 sg13g2_antennanp ANTENNA_2129 (.A(net959));
 sg13g2_antennanp ANTENNA_2130 (.A(net959));
 sg13g2_antennanp ANTENNA_2131 (.A(net959));
 sg13g2_antennanp ANTENNA_2132 (.A(net959));
 sg13g2_antennanp ANTENNA_2133 (.A(net959));
 sg13g2_antennanp ANTENNA_2134 (.A(net959));
 sg13g2_antennanp ANTENNA_2135 (.A(net959));
 sg13g2_antennanp ANTENNA_2136 (.A(net959));
 sg13g2_antennanp ANTENNA_2137 (.A(net967));
 sg13g2_antennanp ANTENNA_2138 (.A(net967));
 sg13g2_antennanp ANTENNA_2139 (.A(net967));
 sg13g2_antennanp ANTENNA_2140 (.A(net967));
 sg13g2_antennanp ANTENNA_2141 (.A(net967));
 sg13g2_antennanp ANTENNA_2142 (.A(net967));
 sg13g2_antennanp ANTENNA_2143 (.A(net967));
 sg13g2_antennanp ANTENNA_2144 (.A(net967));
 sg13g2_antennanp ANTENNA_2145 (.A(net967));
 sg13g2_antennanp ANTENNA_2146 (.A(net972));
 sg13g2_antennanp ANTENNA_2147 (.A(net972));
 sg13g2_antennanp ANTENNA_2148 (.A(net972));
 sg13g2_antennanp ANTENNA_2149 (.A(net972));
 sg13g2_antennanp ANTENNA_2150 (.A(net972));
 sg13g2_antennanp ANTENNA_2151 (.A(net972));
 sg13g2_antennanp ANTENNA_2152 (.A(net972));
 sg13g2_antennanp ANTENNA_2153 (.A(net972));
 sg13g2_antennanp ANTENNA_2154 (.A(net972));
 sg13g2_antennanp ANTENNA_2155 (.A(net972));
 sg13g2_antennanp ANTENNA_2156 (.A(net972));
 sg13g2_antennanp ANTENNA_2157 (.A(net972));
 sg13g2_antennanp ANTENNA_2158 (.A(net972));
 sg13g2_antennanp ANTENNA_2159 (.A(net972));
 sg13g2_antennanp ANTENNA_2160 (.A(net972));
 sg13g2_antennanp ANTENNA_2161 (.A(net972));
 sg13g2_antennanp ANTENNA_2162 (.A(net1000));
 sg13g2_antennanp ANTENNA_2163 (.A(net1000));
 sg13g2_antennanp ANTENNA_2164 (.A(net1000));
 sg13g2_antennanp ANTENNA_2165 (.A(net1000));
 sg13g2_antennanp ANTENNA_2166 (.A(net1000));
 sg13g2_antennanp ANTENNA_2167 (.A(net1000));
 sg13g2_antennanp ANTENNA_2168 (.A(net1000));
 sg13g2_antennanp ANTENNA_2169 (.A(net1000));
 sg13g2_antennanp ANTENNA_2170 (.A(net1043));
 sg13g2_antennanp ANTENNA_2171 (.A(net1043));
 sg13g2_antennanp ANTENNA_2172 (.A(net1043));
 sg13g2_antennanp ANTENNA_2173 (.A(net1043));
 sg13g2_antennanp ANTENNA_2174 (.A(net1043));
 sg13g2_antennanp ANTENNA_2175 (.A(net1043));
 sg13g2_antennanp ANTENNA_2176 (.A(net1043));
 sg13g2_antennanp ANTENNA_2177 (.A(net1043));
 sg13g2_antennanp ANTENNA_2178 (.A(net1043));
 sg13g2_antennanp ANTENNA_2179 (.A(net1043));
 sg13g2_antennanp ANTENNA_2180 (.A(net1043));
 sg13g2_antennanp ANTENNA_2181 (.A(net1043));
 sg13g2_antennanp ANTENNA_2182 (.A(net1043));
 sg13g2_antennanp ANTENNA_2183 (.A(net1043));
 sg13g2_antennanp ANTENNA_2184 (.A(net1043));
 sg13g2_antennanp ANTENNA_2185 (.A(net1043));
 sg13g2_antennanp ANTENNA_2186 (.A(net1043));
 sg13g2_antennanp ANTENNA_2187 (.A(net1043));
 sg13g2_antennanp ANTENNA_2188 (.A(net1043));
 sg13g2_antennanp ANTENNA_2189 (.A(net1043));
 sg13g2_antennanp ANTENNA_2190 (.A(net1043));
 sg13g2_antennanp ANTENNA_2191 (.A(net1043));
 sg13g2_antennanp ANTENNA_2192 (.A(net1043));
 sg13g2_antennanp ANTENNA_2193 (.A(net1043));
 sg13g2_antennanp ANTENNA_2194 (.A(net1043));
 sg13g2_antennanp ANTENNA_2195 (.A(net1043));
 sg13g2_antennanp ANTENNA_2196 (.A(net1043));
 sg13g2_antennanp ANTENNA_2197 (.A(net1043));
 sg13g2_antennanp ANTENNA_2198 (.A(net1043));
 sg13g2_antennanp ANTENNA_2199 (.A(net1043));
 sg13g2_antennanp ANTENNA_2200 (.A(net1053));
 sg13g2_antennanp ANTENNA_2201 (.A(net1053));
 sg13g2_antennanp ANTENNA_2202 (.A(net1053));
 sg13g2_antennanp ANTENNA_2203 (.A(net1053));
 sg13g2_antennanp ANTENNA_2204 (.A(net1053));
 sg13g2_antennanp ANTENNA_2205 (.A(net1053));
 sg13g2_antennanp ANTENNA_2206 (.A(net1053));
 sg13g2_antennanp ANTENNA_2207 (.A(net1053));
 sg13g2_antennanp ANTENNA_2208 (.A(net1072));
 sg13g2_antennanp ANTENNA_2209 (.A(net1072));
 sg13g2_antennanp ANTENNA_2210 (.A(net1072));
 sg13g2_antennanp ANTENNA_2211 (.A(net1072));
 sg13g2_antennanp ANTENNA_2212 (.A(net1072));
 sg13g2_antennanp ANTENNA_2213 (.A(net1072));
 sg13g2_antennanp ANTENNA_2214 (.A(net1072));
 sg13g2_antennanp ANTENNA_2215 (.A(net1072));
 sg13g2_antennanp ANTENNA_2216 (.A(net1072));
 sg13g2_antennanp ANTENNA_2217 (.A(net1104));
 sg13g2_antennanp ANTENNA_2218 (.A(net1104));
 sg13g2_antennanp ANTENNA_2219 (.A(net1104));
 sg13g2_antennanp ANTENNA_2220 (.A(net1104));
 sg13g2_antennanp ANTENNA_2221 (.A(net1104));
 sg13g2_antennanp ANTENNA_2222 (.A(net1104));
 sg13g2_antennanp ANTENNA_2223 (.A(net1104));
 sg13g2_antennanp ANTENNA_2224 (.A(net1104));
 sg13g2_antennanp ANTENNA_2225 (.A(net1104));
 sg13g2_antennanp ANTENNA_2226 (.A(net1104));
 sg13g2_antennanp ANTENNA_2227 (.A(net1104));
 sg13g2_antennanp ANTENNA_2228 (.A(_00928_));
 sg13g2_antennanp ANTENNA_2229 (.A(_01057_));
 sg13g2_antennanp ANTENNA_2230 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2231 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2232 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2233 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2234 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2235 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2236 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2237 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2238 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2239 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2240 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2241 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2242 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2243 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2244 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2245 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2246 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2247 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2248 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2249 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2250 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2251 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2252 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2253 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2254 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2255 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2256 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2257 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2258 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2259 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2260 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2261 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2262 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2263 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2264 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2265 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2266 (.A(_03019_));
 sg13g2_antennanp ANTENNA_2267 (.A(_03019_));
 sg13g2_antennanp ANTENNA_2268 (.A(_03019_));
 sg13g2_antennanp ANTENNA_2269 (.A(_03865_));
 sg13g2_antennanp ANTENNA_2270 (.A(_03865_));
 sg13g2_antennanp ANTENNA_2271 (.A(_03865_));
 sg13g2_antennanp ANTENNA_2272 (.A(_03865_));
 sg13g2_antennanp ANTENNA_2273 (.A(_05015_));
 sg13g2_antennanp ANTENNA_2274 (.A(_05223_));
 sg13g2_antennanp ANTENNA_2275 (.A(_05238_));
 sg13g2_antennanp ANTENNA_2276 (.A(_05278_));
 sg13g2_antennanp ANTENNA_2277 (.A(_05291_));
 sg13g2_antennanp ANTENNA_2278 (.A(_05306_));
 sg13g2_antennanp ANTENNA_2279 (.A(_05323_));
 sg13g2_antennanp ANTENNA_2280 (.A(_05333_));
 sg13g2_antennanp ANTENNA_2281 (.A(_05406_));
 sg13g2_antennanp ANTENNA_2282 (.A(_05406_));
 sg13g2_antennanp ANTENNA_2283 (.A(_05406_));
 sg13g2_antennanp ANTENNA_2284 (.A(_05478_));
 sg13g2_antennanp ANTENNA_2285 (.A(_05483_));
 sg13g2_antennanp ANTENNA_2286 (.A(_05545_));
 sg13g2_antennanp ANTENNA_2287 (.A(_05551_));
 sg13g2_antennanp ANTENNA_2288 (.A(_05781_));
 sg13g2_antennanp ANTENNA_2289 (.A(_05797_));
 sg13g2_antennanp ANTENNA_2290 (.A(_05798_));
 sg13g2_antennanp ANTENNA_2291 (.A(_05798_));
 sg13g2_antennanp ANTENNA_2292 (.A(_05798_));
 sg13g2_antennanp ANTENNA_2293 (.A(_05801_));
 sg13g2_antennanp ANTENNA_2294 (.A(_05801_));
 sg13g2_antennanp ANTENNA_2295 (.A(_05801_));
 sg13g2_antennanp ANTENNA_2296 (.A(_05801_));
 sg13g2_antennanp ANTENNA_2297 (.A(_05815_));
 sg13g2_antennanp ANTENNA_2298 (.A(_05818_));
 sg13g2_antennanp ANTENNA_2299 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2300 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2301 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2302 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2303 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2304 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2305 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2306 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2307 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2308 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2309 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2310 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2311 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2312 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2313 (.A(_06735_));
 sg13g2_antennanp ANTENNA_2314 (.A(_06735_));
 sg13g2_antennanp ANTENNA_2315 (.A(_06735_));
 sg13g2_antennanp ANTENNA_2316 (.A(_06735_));
 sg13g2_antennanp ANTENNA_2317 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2318 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2319 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2320 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2321 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2322 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2323 (.A(_07611_));
 sg13g2_antennanp ANTENNA_2324 (.A(_07611_));
 sg13g2_antennanp ANTENNA_2325 (.A(_07611_));
 sg13g2_antennanp ANTENNA_2326 (.A(_07611_));
 sg13g2_antennanp ANTENNA_2327 (.A(_08265_));
 sg13g2_antennanp ANTENNA_2328 (.A(_08265_));
 sg13g2_antennanp ANTENNA_2329 (.A(_08265_));
 sg13g2_antennanp ANTENNA_2330 (.A(_08265_));
 sg13g2_antennanp ANTENNA_2331 (.A(_08265_));
 sg13g2_antennanp ANTENNA_2332 (.A(_08265_));
 sg13g2_antennanp ANTENNA_2333 (.A(_08278_));
 sg13g2_antennanp ANTENNA_2334 (.A(_08278_));
 sg13g2_antennanp ANTENNA_2335 (.A(_08278_));
 sg13g2_antennanp ANTENNA_2336 (.A(_08278_));
 sg13g2_antennanp ANTENNA_2337 (.A(_08648_));
 sg13g2_antennanp ANTENNA_2338 (.A(_08648_));
 sg13g2_antennanp ANTENNA_2339 (.A(_08648_));
 sg13g2_antennanp ANTENNA_2340 (.A(_08648_));
 sg13g2_antennanp ANTENNA_2341 (.A(_08648_));
 sg13g2_antennanp ANTENNA_2342 (.A(_08648_));
 sg13g2_antennanp ANTENNA_2343 (.A(_08681_));
 sg13g2_antennanp ANTENNA_2344 (.A(_08681_));
 sg13g2_antennanp ANTENNA_2345 (.A(_08681_));
 sg13g2_antennanp ANTENNA_2346 (.A(_08681_));
 sg13g2_antennanp ANTENNA_2347 (.A(_08712_));
 sg13g2_antennanp ANTENNA_2348 (.A(_08712_));
 sg13g2_antennanp ANTENNA_2349 (.A(_08758_));
 sg13g2_antennanp ANTENNA_2350 (.A(_08758_));
 sg13g2_antennanp ANTENNA_2351 (.A(_08758_));
 sg13g2_antennanp ANTENNA_2352 (.A(_08758_));
 sg13g2_antennanp ANTENNA_2353 (.A(_08758_));
 sg13g2_antennanp ANTENNA_2354 (.A(_08758_));
 sg13g2_antennanp ANTENNA_2355 (.A(_08758_));
 sg13g2_antennanp ANTENNA_2356 (.A(_08758_));
 sg13g2_antennanp ANTENNA_2357 (.A(_08758_));
 sg13g2_antennanp ANTENNA_2358 (.A(_08758_));
 sg13g2_antennanp ANTENNA_2359 (.A(_08797_));
 sg13g2_antennanp ANTENNA_2360 (.A(_08797_));
 sg13g2_antennanp ANTENNA_2361 (.A(_08797_));
 sg13g2_antennanp ANTENNA_2362 (.A(_08797_));
 sg13g2_antennanp ANTENNA_2363 (.A(_08797_));
 sg13g2_antennanp ANTENNA_2364 (.A(_08817_));
 sg13g2_antennanp ANTENNA_2365 (.A(_08817_));
 sg13g2_antennanp ANTENNA_2366 (.A(_08817_));
 sg13g2_antennanp ANTENNA_2367 (.A(_08817_));
 sg13g2_antennanp ANTENNA_2368 (.A(_08817_));
 sg13g2_antennanp ANTENNA_2369 (.A(_08840_));
 sg13g2_antennanp ANTENNA_2370 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2371 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2372 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2373 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2374 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2375 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2376 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2377 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2378 (.A(_08919_));
 sg13g2_antennanp ANTENNA_2379 (.A(_08944_));
 sg13g2_antennanp ANTENNA_2380 (.A(_08944_));
 sg13g2_antennanp ANTENNA_2381 (.A(_08944_));
 sg13g2_antennanp ANTENNA_2382 (.A(_08964_));
 sg13g2_antennanp ANTENNA_2383 (.A(_08965_));
 sg13g2_antennanp ANTENNA_2384 (.A(_08965_));
 sg13g2_antennanp ANTENNA_2385 (.A(_08988_));
 sg13g2_antennanp ANTENNA_2386 (.A(_08988_));
 sg13g2_antennanp ANTENNA_2387 (.A(_08988_));
 sg13g2_antennanp ANTENNA_2388 (.A(_08997_));
 sg13g2_antennanp ANTENNA_2389 (.A(_09012_));
 sg13g2_antennanp ANTENNA_2390 (.A(_09012_));
 sg13g2_antennanp ANTENNA_2391 (.A(_09012_));
 sg13g2_antennanp ANTENNA_2392 (.A(_09012_));
 sg13g2_antennanp ANTENNA_2393 (.A(_09205_));
 sg13g2_antennanp ANTENNA_2394 (.A(_09205_));
 sg13g2_antennanp ANTENNA_2395 (.A(_09205_));
 sg13g2_antennanp ANTENNA_2396 (.A(_09205_));
 sg13g2_antennanp ANTENNA_2397 (.A(_09255_));
 sg13g2_antennanp ANTENNA_2398 (.A(_09255_));
 sg13g2_antennanp ANTENNA_2399 (.A(_09255_));
 sg13g2_antennanp ANTENNA_2400 (.A(_09255_));
 sg13g2_antennanp ANTENNA_2401 (.A(_09258_));
 sg13g2_antennanp ANTENNA_2402 (.A(_09258_));
 sg13g2_antennanp ANTENNA_2403 (.A(_09258_));
 sg13g2_antennanp ANTENNA_2404 (.A(_09258_));
 sg13g2_antennanp ANTENNA_2405 (.A(_09260_));
 sg13g2_antennanp ANTENNA_2406 (.A(_09294_));
 sg13g2_antennanp ANTENNA_2407 (.A(_09294_));
 sg13g2_antennanp ANTENNA_2408 (.A(_09294_));
 sg13g2_antennanp ANTENNA_2409 (.A(_09294_));
 sg13g2_antennanp ANTENNA_2410 (.A(_09297_));
 sg13g2_antennanp ANTENNA_2411 (.A(_09297_));
 sg13g2_antennanp ANTENNA_2412 (.A(_09297_));
 sg13g2_antennanp ANTENNA_2413 (.A(_09297_));
 sg13g2_antennanp ANTENNA_2414 (.A(_09463_));
 sg13g2_antennanp ANTENNA_2415 (.A(_09488_));
 sg13g2_antennanp ANTENNA_2416 (.A(_09512_));
 sg13g2_antennanp ANTENNA_2417 (.A(_09524_));
 sg13g2_antennanp ANTENNA_2418 (.A(_09524_));
 sg13g2_antennanp ANTENNA_2419 (.A(_09524_));
 sg13g2_antennanp ANTENNA_2420 (.A(_09544_));
 sg13g2_antennanp ANTENNA_2421 (.A(_09552_));
 sg13g2_antennanp ANTENNA_2422 (.A(_09639_));
 sg13g2_antennanp ANTENNA_2423 (.A(_09664_));
 sg13g2_antennanp ANTENNA_2424 (.A(_09685_));
 sg13g2_antennanp ANTENNA_2425 (.A(_09712_));
 sg13g2_antennanp ANTENNA_2426 (.A(_09727_));
 sg13g2_antennanp ANTENNA_2427 (.A(_09744_));
 sg13g2_antennanp ANTENNA_2428 (.A(_09744_));
 sg13g2_antennanp ANTENNA_2429 (.A(_09744_));
 sg13g2_antennanp ANTENNA_2430 (.A(_09744_));
 sg13g2_antennanp ANTENNA_2431 (.A(_09753_));
 sg13g2_antennanp ANTENNA_2432 (.A(_09798_));
 sg13g2_antennanp ANTENNA_2433 (.A(_09798_));
 sg13g2_antennanp ANTENNA_2434 (.A(_09954_));
 sg13g2_antennanp ANTENNA_2435 (.A(_09954_));
 sg13g2_antennanp ANTENNA_2436 (.A(_09954_));
 sg13g2_antennanp ANTENNA_2437 (.A(_09954_));
 sg13g2_antennanp ANTENNA_2438 (.A(_09954_));
 sg13g2_antennanp ANTENNA_2439 (.A(_09954_));
 sg13g2_antennanp ANTENNA_2440 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2441 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2442 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2443 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2444 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2445 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2446 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2447 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2448 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2449 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2450 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2451 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2452 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2453 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2454 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2455 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2456 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2457 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2458 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2459 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2460 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2461 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2462 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2463 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2464 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2465 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2466 (.A(_10107_));
 sg13g2_antennanp ANTENNA_2467 (.A(_10107_));
 sg13g2_antennanp ANTENNA_2468 (.A(_10107_));
 sg13g2_antennanp ANTENNA_2469 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2470 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2471 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2472 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2473 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2474 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2475 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2476 (.A(_10386_));
 sg13g2_antennanp ANTENNA_2477 (.A(_10386_));
 sg13g2_antennanp ANTENNA_2478 (.A(_10572_));
 sg13g2_antennanp ANTENNA_2479 (.A(_10572_));
 sg13g2_antennanp ANTENNA_2480 (.A(_10572_));
 sg13g2_antennanp ANTENNA_2481 (.A(_10572_));
 sg13g2_antennanp ANTENNA_2482 (.A(_10703_));
 sg13g2_antennanp ANTENNA_2483 (.A(_10703_));
 sg13g2_antennanp ANTENNA_2484 (.A(_10703_));
 sg13g2_antennanp ANTENNA_2485 (.A(_10889_));
 sg13g2_antennanp ANTENNA_2486 (.A(_10889_));
 sg13g2_antennanp ANTENNA_2487 (.A(_10889_));
 sg13g2_antennanp ANTENNA_2488 (.A(_10889_));
 sg13g2_antennanp ANTENNA_2489 (.A(_10889_));
 sg13g2_antennanp ANTENNA_2490 (.A(_10889_));
 sg13g2_antennanp ANTENNA_2491 (.A(_11885_));
 sg13g2_antennanp ANTENNA_2492 (.A(_11885_));
 sg13g2_antennanp ANTENNA_2493 (.A(_11885_));
 sg13g2_antennanp ANTENNA_2494 (.A(_11970_));
 sg13g2_antennanp ANTENNA_2495 (.A(_11970_));
 sg13g2_antennanp ANTENNA_2496 (.A(_11970_));
 sg13g2_antennanp ANTENNA_2497 (.A(_12023_));
 sg13g2_antennanp ANTENNA_2498 (.A(_12023_));
 sg13g2_antennanp ANTENNA_2499 (.A(_12023_));
 sg13g2_antennanp ANTENNA_2500 (.A(_12023_));
 sg13g2_antennanp ANTENNA_2501 (.A(_12023_));
 sg13g2_antennanp ANTENNA_2502 (.A(_12023_));
 sg13g2_antennanp ANTENNA_2503 (.A(_12023_));
 sg13g2_antennanp ANTENNA_2504 (.A(_12023_));
 sg13g2_antennanp ANTENNA_2505 (.A(_12023_));
 sg13g2_antennanp ANTENNA_2506 (.A(_12046_));
 sg13g2_antennanp ANTENNA_2507 (.A(_12046_));
 sg13g2_antennanp ANTENNA_2508 (.A(_12046_));
 sg13g2_antennanp ANTENNA_2509 (.A(_12046_));
 sg13g2_antennanp ANTENNA_2510 (.A(_12046_));
 sg13g2_antennanp ANTENNA_2511 (.A(_12046_));
 sg13g2_antennanp ANTENNA_2512 (.A(_12046_));
 sg13g2_antennanp ANTENNA_2513 (.A(_12046_));
 sg13g2_antennanp ANTENNA_2514 (.A(_12046_));
 sg13g2_antennanp ANTENNA_2515 (.A(_12063_));
 sg13g2_antennanp ANTENNA_2516 (.A(_12063_));
 sg13g2_antennanp ANTENNA_2517 (.A(_12063_));
 sg13g2_antennanp ANTENNA_2518 (.A(_12063_));
 sg13g2_antennanp ANTENNA_2519 (.A(_12063_));
 sg13g2_antennanp ANTENNA_2520 (.A(_12063_));
 sg13g2_antennanp ANTENNA_2521 (.A(_12063_));
 sg13g2_antennanp ANTENNA_2522 (.A(_12063_));
 sg13g2_antennanp ANTENNA_2523 (.A(_12063_));
 sg13g2_antennanp ANTENNA_2524 (.A(_12084_));
 sg13g2_antennanp ANTENNA_2525 (.A(_12084_));
 sg13g2_antennanp ANTENNA_2526 (.A(_12084_));
 sg13g2_antennanp ANTENNA_2527 (.A(_12096_));
 sg13g2_antennanp ANTENNA_2528 (.A(_12096_));
 sg13g2_antennanp ANTENNA_2529 (.A(_12096_));
 sg13g2_antennanp ANTENNA_2530 (.A(_12096_));
 sg13g2_antennanp ANTENNA_2531 (.A(_12096_));
 sg13g2_antennanp ANTENNA_2532 (.A(_12096_));
 sg13g2_antennanp ANTENNA_2533 (.A(_12096_));
 sg13g2_antennanp ANTENNA_2534 (.A(_12096_));
 sg13g2_antennanp ANTENNA_2535 (.A(_12096_));
 sg13g2_antennanp ANTENNA_2536 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2537 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2538 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2539 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2540 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2541 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2542 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2543 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2544 (.A(_12133_));
 sg13g2_antennanp ANTENNA_2545 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2546 (.A(r_reset));
 sg13g2_antennanp ANTENNA_2547 (.A(r_reset));
 sg13g2_antennanp ANTENNA_2548 (.A(r_reset));
 sg13g2_antennanp ANTENNA_2549 (.A(net1));
 sg13g2_antennanp ANTENNA_2550 (.A(net1));
 sg13g2_antennanp ANTENNA_2551 (.A(net1));
 sg13g2_antennanp ANTENNA_2552 (.A(net2));
 sg13g2_antennanp ANTENNA_2553 (.A(net2));
 sg13g2_antennanp ANTENNA_2554 (.A(net12));
 sg13g2_antennanp ANTENNA_2555 (.A(net12));
 sg13g2_antennanp ANTENNA_2556 (.A(net12));
 sg13g2_antennanp ANTENNA_2557 (.A(net13));
 sg13g2_antennanp ANTENNA_2558 (.A(net13));
 sg13g2_antennanp ANTENNA_2559 (.A(net13));
 sg13g2_antennanp ANTENNA_2560 (.A(net19));
 sg13g2_antennanp ANTENNA_2561 (.A(net19));
 sg13g2_antennanp ANTENNA_2562 (.A(net20));
 sg13g2_antennanp ANTENNA_2563 (.A(net20));
 sg13g2_antennanp ANTENNA_2564 (.A(net596));
 sg13g2_antennanp ANTENNA_2565 (.A(net596));
 sg13g2_antennanp ANTENNA_2566 (.A(net596));
 sg13g2_antennanp ANTENNA_2567 (.A(net596));
 sg13g2_antennanp ANTENNA_2568 (.A(net596));
 sg13g2_antennanp ANTENNA_2569 (.A(net596));
 sg13g2_antennanp ANTENNA_2570 (.A(net596));
 sg13g2_antennanp ANTENNA_2571 (.A(net596));
 sg13g2_antennanp ANTENNA_2572 (.A(net596));
 sg13g2_antennanp ANTENNA_2573 (.A(net618));
 sg13g2_antennanp ANTENNA_2574 (.A(net618));
 sg13g2_antennanp ANTENNA_2575 (.A(net618));
 sg13g2_antennanp ANTENNA_2576 (.A(net618));
 sg13g2_antennanp ANTENNA_2577 (.A(net618));
 sg13g2_antennanp ANTENNA_2578 (.A(net618));
 sg13g2_antennanp ANTENNA_2579 (.A(net618));
 sg13g2_antennanp ANTENNA_2580 (.A(net618));
 sg13g2_antennanp ANTENNA_2581 (.A(net618));
 sg13g2_antennanp ANTENNA_2582 (.A(net618));
 sg13g2_antennanp ANTENNA_2583 (.A(net618));
 sg13g2_antennanp ANTENNA_2584 (.A(net618));
 sg13g2_antennanp ANTENNA_2585 (.A(net631));
 sg13g2_antennanp ANTENNA_2586 (.A(net631));
 sg13g2_antennanp ANTENNA_2587 (.A(net631));
 sg13g2_antennanp ANTENNA_2588 (.A(net631));
 sg13g2_antennanp ANTENNA_2589 (.A(net631));
 sg13g2_antennanp ANTENNA_2590 (.A(net631));
 sg13g2_antennanp ANTENNA_2591 (.A(net631));
 sg13g2_antennanp ANTENNA_2592 (.A(net631));
 sg13g2_antennanp ANTENNA_2593 (.A(net651));
 sg13g2_antennanp ANTENNA_2594 (.A(net651));
 sg13g2_antennanp ANTENNA_2595 (.A(net651));
 sg13g2_antennanp ANTENNA_2596 (.A(net651));
 sg13g2_antennanp ANTENNA_2597 (.A(net651));
 sg13g2_antennanp ANTENNA_2598 (.A(net651));
 sg13g2_antennanp ANTENNA_2599 (.A(net651));
 sg13g2_antennanp ANTENNA_2600 (.A(net651));
 sg13g2_antennanp ANTENNA_2601 (.A(net651));
 sg13g2_antennanp ANTENNA_2602 (.A(net651));
 sg13g2_antennanp ANTENNA_2603 (.A(net651));
 sg13g2_antennanp ANTENNA_2604 (.A(net651));
 sg13g2_antennanp ANTENNA_2605 (.A(net651));
 sg13g2_antennanp ANTENNA_2606 (.A(net651));
 sg13g2_antennanp ANTENNA_2607 (.A(net651));
 sg13g2_antennanp ANTENNA_2608 (.A(net651));
 sg13g2_antennanp ANTENNA_2609 (.A(net651));
 sg13g2_antennanp ANTENNA_2610 (.A(net651));
 sg13g2_antennanp ANTENNA_2611 (.A(net651));
 sg13g2_antennanp ANTENNA_2612 (.A(net651));
 sg13g2_antennanp ANTENNA_2613 (.A(net651));
 sg13g2_antennanp ANTENNA_2614 (.A(net651));
 sg13g2_antennanp ANTENNA_2615 (.A(net860));
 sg13g2_antennanp ANTENNA_2616 (.A(net860));
 sg13g2_antennanp ANTENNA_2617 (.A(net860));
 sg13g2_antennanp ANTENNA_2618 (.A(net860));
 sg13g2_antennanp ANTENNA_2619 (.A(net860));
 sg13g2_antennanp ANTENNA_2620 (.A(net860));
 sg13g2_antennanp ANTENNA_2621 (.A(net860));
 sg13g2_antennanp ANTENNA_2622 (.A(net860));
 sg13g2_antennanp ANTENNA_2623 (.A(net860));
 sg13g2_antennanp ANTENNA_2624 (.A(net891));
 sg13g2_antennanp ANTENNA_2625 (.A(net891));
 sg13g2_antennanp ANTENNA_2626 (.A(net891));
 sg13g2_antennanp ANTENNA_2627 (.A(net891));
 sg13g2_antennanp ANTENNA_2628 (.A(net891));
 sg13g2_antennanp ANTENNA_2629 (.A(net891));
 sg13g2_antennanp ANTENNA_2630 (.A(net891));
 sg13g2_antennanp ANTENNA_2631 (.A(net891));
 sg13g2_antennanp ANTENNA_2632 (.A(net891));
 sg13g2_antennanp ANTENNA_2633 (.A(net899));
 sg13g2_antennanp ANTENNA_2634 (.A(net899));
 sg13g2_antennanp ANTENNA_2635 (.A(net899));
 sg13g2_antennanp ANTENNA_2636 (.A(net899));
 sg13g2_antennanp ANTENNA_2637 (.A(net899));
 sg13g2_antennanp ANTENNA_2638 (.A(net899));
 sg13g2_antennanp ANTENNA_2639 (.A(net899));
 sg13g2_antennanp ANTENNA_2640 (.A(net899));
 sg13g2_antennanp ANTENNA_2641 (.A(net899));
 sg13g2_antennanp ANTENNA_2642 (.A(net899));
 sg13g2_antennanp ANTENNA_2643 (.A(net899));
 sg13g2_antennanp ANTENNA_2644 (.A(net899));
 sg13g2_antennanp ANTENNA_2645 (.A(net899));
 sg13g2_antennanp ANTENNA_2646 (.A(net899));
 sg13g2_antennanp ANTENNA_2647 (.A(net899));
 sg13g2_antennanp ANTENNA_2648 (.A(net899));
 sg13g2_antennanp ANTENNA_2649 (.A(net899));
 sg13g2_antennanp ANTENNA_2650 (.A(net899));
 sg13g2_antennanp ANTENNA_2651 (.A(net899));
 sg13g2_antennanp ANTENNA_2652 (.A(net899));
 sg13g2_antennanp ANTENNA_2653 (.A(net959));
 sg13g2_antennanp ANTENNA_2654 (.A(net959));
 sg13g2_antennanp ANTENNA_2655 (.A(net959));
 sg13g2_antennanp ANTENNA_2656 (.A(net959));
 sg13g2_antennanp ANTENNA_2657 (.A(net959));
 sg13g2_antennanp ANTENNA_2658 (.A(net959));
 sg13g2_antennanp ANTENNA_2659 (.A(net959));
 sg13g2_antennanp ANTENNA_2660 (.A(net959));
 sg13g2_antennanp ANTENNA_2661 (.A(net959));
 sg13g2_antennanp ANTENNA_2662 (.A(net970));
 sg13g2_antennanp ANTENNA_2663 (.A(net970));
 sg13g2_antennanp ANTENNA_2664 (.A(net970));
 sg13g2_antennanp ANTENNA_2665 (.A(net970));
 sg13g2_antennanp ANTENNA_2666 (.A(net970));
 sg13g2_antennanp ANTENNA_2667 (.A(net970));
 sg13g2_antennanp ANTENNA_2668 (.A(net970));
 sg13g2_antennanp ANTENNA_2669 (.A(net970));
 sg13g2_antennanp ANTENNA_2670 (.A(net971));
 sg13g2_antennanp ANTENNA_2671 (.A(net971));
 sg13g2_antennanp ANTENNA_2672 (.A(net971));
 sg13g2_antennanp ANTENNA_2673 (.A(net971));
 sg13g2_antennanp ANTENNA_2674 (.A(net971));
 sg13g2_antennanp ANTENNA_2675 (.A(net971));
 sg13g2_antennanp ANTENNA_2676 (.A(net971));
 sg13g2_antennanp ANTENNA_2677 (.A(net971));
 sg13g2_antennanp ANTENNA_2678 (.A(net971));
 sg13g2_antennanp ANTENNA_2679 (.A(net971));
 sg13g2_antennanp ANTENNA_2680 (.A(net971));
 sg13g2_antennanp ANTENNA_2681 (.A(net971));
 sg13g2_antennanp ANTENNA_2682 (.A(net971));
 sg13g2_antennanp ANTENNA_2683 (.A(net971));
 sg13g2_antennanp ANTENNA_2684 (.A(net971));
 sg13g2_antennanp ANTENNA_2685 (.A(net972));
 sg13g2_antennanp ANTENNA_2686 (.A(net972));
 sg13g2_antennanp ANTENNA_2687 (.A(net972));
 sg13g2_antennanp ANTENNA_2688 (.A(net972));
 sg13g2_antennanp ANTENNA_2689 (.A(net972));
 sg13g2_antennanp ANTENNA_2690 (.A(net972));
 sg13g2_antennanp ANTENNA_2691 (.A(net972));
 sg13g2_antennanp ANTENNA_2692 (.A(net972));
 sg13g2_antennanp ANTENNA_2693 (.A(net972));
 sg13g2_antennanp ANTENNA_2694 (.A(net972));
 sg13g2_antennanp ANTENNA_2695 (.A(net972));
 sg13g2_antennanp ANTENNA_2696 (.A(net1000));
 sg13g2_antennanp ANTENNA_2697 (.A(net1000));
 sg13g2_antennanp ANTENNA_2698 (.A(net1000));
 sg13g2_antennanp ANTENNA_2699 (.A(net1000));
 sg13g2_antennanp ANTENNA_2700 (.A(net1000));
 sg13g2_antennanp ANTENNA_2701 (.A(net1000));
 sg13g2_antennanp ANTENNA_2702 (.A(net1000));
 sg13g2_antennanp ANTENNA_2703 (.A(net1000));
 sg13g2_antennanp ANTENNA_2704 (.A(net1043));
 sg13g2_antennanp ANTENNA_2705 (.A(net1043));
 sg13g2_antennanp ANTENNA_2706 (.A(net1043));
 sg13g2_antennanp ANTENNA_2707 (.A(net1043));
 sg13g2_antennanp ANTENNA_2708 (.A(net1043));
 sg13g2_antennanp ANTENNA_2709 (.A(net1043));
 sg13g2_antennanp ANTENNA_2710 (.A(net1043));
 sg13g2_antennanp ANTENNA_2711 (.A(net1043));
 sg13g2_antennanp ANTENNA_2712 (.A(net1043));
 sg13g2_antennanp ANTENNA_2713 (.A(net1043));
 sg13g2_antennanp ANTENNA_2714 (.A(net1043));
 sg13g2_antennanp ANTENNA_2715 (.A(net1043));
 sg13g2_antennanp ANTENNA_2716 (.A(net1053));
 sg13g2_antennanp ANTENNA_2717 (.A(net1053));
 sg13g2_antennanp ANTENNA_2718 (.A(net1053));
 sg13g2_antennanp ANTENNA_2719 (.A(net1053));
 sg13g2_antennanp ANTENNA_2720 (.A(net1053));
 sg13g2_antennanp ANTENNA_2721 (.A(net1053));
 sg13g2_antennanp ANTENNA_2722 (.A(net1053));
 sg13g2_antennanp ANTENNA_2723 (.A(net1053));
 sg13g2_antennanp ANTENNA_2724 (.A(net1072));
 sg13g2_antennanp ANTENNA_2725 (.A(net1072));
 sg13g2_antennanp ANTENNA_2726 (.A(net1072));
 sg13g2_antennanp ANTENNA_2727 (.A(net1072));
 sg13g2_antennanp ANTENNA_2728 (.A(net1072));
 sg13g2_antennanp ANTENNA_2729 (.A(net1072));
 sg13g2_antennanp ANTENNA_2730 (.A(net1072));
 sg13g2_antennanp ANTENNA_2731 (.A(net1072));
 sg13g2_antennanp ANTENNA_2732 (.A(net1072));
 sg13g2_antennanp ANTENNA_2733 (.A(net1104));
 sg13g2_antennanp ANTENNA_2734 (.A(net1104));
 sg13g2_antennanp ANTENNA_2735 (.A(net1104));
 sg13g2_antennanp ANTENNA_2736 (.A(net1104));
 sg13g2_antennanp ANTENNA_2737 (.A(net1104));
 sg13g2_antennanp ANTENNA_2738 (.A(net1104));
 sg13g2_antennanp ANTENNA_2739 (.A(net1104));
 sg13g2_antennanp ANTENNA_2740 (.A(net1104));
 sg13g2_antennanp ANTENNA_2741 (.A(net1104));
 sg13g2_antennanp ANTENNA_2742 (.A(net1104));
 sg13g2_antennanp ANTENNA_2743 (.A(net1104));
 sg13g2_antennanp ANTENNA_2744 (.A(_00928_));
 sg13g2_antennanp ANTENNA_2745 (.A(_01057_));
 sg13g2_antennanp ANTENNA_2746 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2747 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2748 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2749 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2750 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2751 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2752 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2753 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2754 (.A(_02823_));
 sg13g2_antennanp ANTENNA_2755 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2756 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2757 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2758 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2759 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2760 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2761 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2762 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2763 (.A(_02831_));
 sg13g2_antennanp ANTENNA_2764 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2765 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2766 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2767 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2768 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2769 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2770 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2771 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2772 (.A(_02835_));
 sg13g2_antennanp ANTENNA_2773 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2774 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2775 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2776 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2777 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2778 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2779 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2780 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2781 (.A(_02990_));
 sg13g2_antennanp ANTENNA_2782 (.A(_03865_));
 sg13g2_antennanp ANTENNA_2783 (.A(_03865_));
 sg13g2_antennanp ANTENNA_2784 (.A(_03865_));
 sg13g2_antennanp ANTENNA_2785 (.A(_03865_));
 sg13g2_antennanp ANTENNA_2786 (.A(_05015_));
 sg13g2_antennanp ANTENNA_2787 (.A(_05223_));
 sg13g2_antennanp ANTENNA_2788 (.A(_05238_));
 sg13g2_antennanp ANTENNA_2789 (.A(_05278_));
 sg13g2_antennanp ANTENNA_2790 (.A(_05279_));
 sg13g2_antennanp ANTENNA_2791 (.A(_05291_));
 sg13g2_antennanp ANTENNA_2792 (.A(_05306_));
 sg13g2_antennanp ANTENNA_2793 (.A(_05323_));
 sg13g2_antennanp ANTENNA_2794 (.A(_05333_));
 sg13g2_antennanp ANTENNA_2795 (.A(_05406_));
 sg13g2_antennanp ANTENNA_2796 (.A(_05406_));
 sg13g2_antennanp ANTENNA_2797 (.A(_05406_));
 sg13g2_antennanp ANTENNA_2798 (.A(_05406_));
 sg13g2_antennanp ANTENNA_2799 (.A(_05478_));
 sg13g2_antennanp ANTENNA_2800 (.A(_05483_));
 sg13g2_antennanp ANTENNA_2801 (.A(_05545_));
 sg13g2_antennanp ANTENNA_2802 (.A(_05551_));
 sg13g2_antennanp ANTENNA_2803 (.A(_05781_));
 sg13g2_antennanp ANTENNA_2804 (.A(_05797_));
 sg13g2_antennanp ANTENNA_2805 (.A(_05801_));
 sg13g2_antennanp ANTENNA_2806 (.A(_05801_));
 sg13g2_antennanp ANTENNA_2807 (.A(_05801_));
 sg13g2_antennanp ANTENNA_2808 (.A(_05801_));
 sg13g2_antennanp ANTENNA_2809 (.A(_05815_));
 sg13g2_antennanp ANTENNA_2810 (.A(_05818_));
 sg13g2_antennanp ANTENNA_2811 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2812 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2813 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2814 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2815 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2816 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2817 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2818 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2819 (.A(_06734_));
 sg13g2_antennanp ANTENNA_2820 (.A(_06735_));
 sg13g2_antennanp ANTENNA_2821 (.A(_06735_));
 sg13g2_antennanp ANTENNA_2822 (.A(_06735_));
 sg13g2_antennanp ANTENNA_2823 (.A(_06735_));
 sg13g2_antennanp ANTENNA_2824 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2825 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2826 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2827 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2828 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2829 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2830 (.A(_07611_));
 sg13g2_antennanp ANTENNA_2831 (.A(_07611_));
 sg13g2_antennanp ANTENNA_2832 (.A(_07611_));
 sg13g2_antennanp ANTENNA_2833 (.A(_07611_));
 sg13g2_antennanp ANTENNA_2834 (.A(_07756_));
 sg13g2_antennanp ANTENNA_2835 (.A(_07756_));
 sg13g2_antennanp ANTENNA_2836 (.A(_07756_));
 sg13g2_antennanp ANTENNA_2837 (.A(_08265_));
 sg13g2_antennanp ANTENNA_2838 (.A(_08265_));
 sg13g2_antennanp ANTENNA_2839 (.A(_08265_));
 sg13g2_antennanp ANTENNA_2840 (.A(_08265_));
 sg13g2_antennanp ANTENNA_2841 (.A(_08265_));
 sg13g2_antennanp ANTENNA_2842 (.A(_08265_));
 sg13g2_antennanp ANTENNA_2843 (.A(_08278_));
 sg13g2_antennanp ANTENNA_2844 (.A(_08278_));
 sg13g2_antennanp ANTENNA_2845 (.A(_08278_));
 sg13g2_antennanp ANTENNA_2846 (.A(_08278_));
 sg13g2_antennanp ANTENNA_2847 (.A(_08648_));
 sg13g2_antennanp ANTENNA_2848 (.A(_08648_));
 sg13g2_antennanp ANTENNA_2849 (.A(_08648_));
 sg13g2_antennanp ANTENNA_2850 (.A(_08648_));
 sg13g2_antennanp ANTENNA_2851 (.A(_08648_));
 sg13g2_antennanp ANTENNA_2852 (.A(_08648_));
 sg13g2_antennanp ANTENNA_2853 (.A(_08681_));
 sg13g2_antennanp ANTENNA_2854 (.A(_08681_));
 sg13g2_antennanp ANTENNA_2855 (.A(_08681_));
 sg13g2_antennanp ANTENNA_2856 (.A(_08681_));
 sg13g2_antennanp ANTENNA_2857 (.A(_08712_));
 sg13g2_antennanp ANTENNA_2858 (.A(_08712_));
 sg13g2_antennanp ANTENNA_2859 (.A(_08788_));
 sg13g2_antennanp ANTENNA_2860 (.A(_08788_));
 sg13g2_antennanp ANTENNA_2861 (.A(_08788_));
 sg13g2_antennanp ANTENNA_2862 (.A(_08788_));
 sg13g2_antennanp ANTENNA_2863 (.A(_08797_));
 sg13g2_antennanp ANTENNA_2864 (.A(_08797_));
 sg13g2_antennanp ANTENNA_2865 (.A(_08797_));
 sg13g2_antennanp ANTENNA_2866 (.A(_08797_));
 sg13g2_antennanp ANTENNA_2867 (.A(_08797_));
 sg13g2_antennanp ANTENNA_2868 (.A(_08817_));
 sg13g2_antennanp ANTENNA_2869 (.A(_08817_));
 sg13g2_antennanp ANTENNA_2870 (.A(_08817_));
 sg13g2_antennanp ANTENNA_2871 (.A(_08817_));
 sg13g2_antennanp ANTENNA_2872 (.A(_08817_));
 sg13g2_antennanp ANTENNA_2873 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2874 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2875 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2876 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2877 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2878 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2879 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2880 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2881 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2882 (.A(_08879_));
 sg13g2_antennanp ANTENNA_2883 (.A(_08919_));
 sg13g2_antennanp ANTENNA_2884 (.A(_08944_));
 sg13g2_antennanp ANTENNA_2885 (.A(_08944_));
 sg13g2_antennanp ANTENNA_2886 (.A(_08944_));
 sg13g2_antennanp ANTENNA_2887 (.A(_08964_));
 sg13g2_antennanp ANTENNA_2888 (.A(_08965_));
 sg13g2_antennanp ANTENNA_2889 (.A(_08965_));
 sg13g2_antennanp ANTENNA_2890 (.A(_08988_));
 sg13g2_antennanp ANTENNA_2891 (.A(_08988_));
 sg13g2_antennanp ANTENNA_2892 (.A(_08988_));
 sg13g2_antennanp ANTENNA_2893 (.A(_08997_));
 sg13g2_antennanp ANTENNA_2894 (.A(_09012_));
 sg13g2_antennanp ANTENNA_2895 (.A(_09012_));
 sg13g2_antennanp ANTENNA_2896 (.A(_09012_));
 sg13g2_antennanp ANTENNA_2897 (.A(_09012_));
 sg13g2_antennanp ANTENNA_2898 (.A(_09205_));
 sg13g2_antennanp ANTENNA_2899 (.A(_09205_));
 sg13g2_antennanp ANTENNA_2900 (.A(_09205_));
 sg13g2_antennanp ANTENNA_2901 (.A(_09205_));
 sg13g2_antennanp ANTENNA_2902 (.A(_09255_));
 sg13g2_antennanp ANTENNA_2903 (.A(_09255_));
 sg13g2_antennanp ANTENNA_2904 (.A(_09255_));
 sg13g2_antennanp ANTENNA_2905 (.A(_09255_));
 sg13g2_antennanp ANTENNA_2906 (.A(_09258_));
 sg13g2_antennanp ANTENNA_2907 (.A(_09258_));
 sg13g2_antennanp ANTENNA_2908 (.A(_09258_));
 sg13g2_antennanp ANTENNA_2909 (.A(_09258_));
 sg13g2_antennanp ANTENNA_2910 (.A(_09294_));
 sg13g2_antennanp ANTENNA_2911 (.A(_09294_));
 sg13g2_antennanp ANTENNA_2912 (.A(_09294_));
 sg13g2_antennanp ANTENNA_2913 (.A(_09294_));
 sg13g2_antennanp ANTENNA_2914 (.A(_09294_));
 sg13g2_antennanp ANTENNA_2915 (.A(_09294_));
 sg13g2_antennanp ANTENNA_2916 (.A(_09294_));
 sg13g2_antennanp ANTENNA_2917 (.A(_09294_));
 sg13g2_antennanp ANTENNA_2918 (.A(_09294_));
 sg13g2_antennanp ANTENNA_2919 (.A(_09297_));
 sg13g2_antennanp ANTENNA_2920 (.A(_09297_));
 sg13g2_antennanp ANTENNA_2921 (.A(_09297_));
 sg13g2_antennanp ANTENNA_2922 (.A(_09297_));
 sg13g2_antennanp ANTENNA_2923 (.A(_09463_));
 sg13g2_antennanp ANTENNA_2924 (.A(_09488_));
 sg13g2_antennanp ANTENNA_2925 (.A(_09512_));
 sg13g2_antennanp ANTENNA_2926 (.A(_09544_));
 sg13g2_antennanp ANTENNA_2927 (.A(_09552_));
 sg13g2_antennanp ANTENNA_2928 (.A(_09639_));
 sg13g2_antennanp ANTENNA_2929 (.A(_09664_));
 sg13g2_antennanp ANTENNA_2930 (.A(_09685_));
 sg13g2_antennanp ANTENNA_2931 (.A(_09712_));
 sg13g2_antennanp ANTENNA_2932 (.A(_09727_));
 sg13g2_antennanp ANTENNA_2933 (.A(_09727_));
 sg13g2_antennanp ANTENNA_2934 (.A(_09744_));
 sg13g2_antennanp ANTENNA_2935 (.A(_09744_));
 sg13g2_antennanp ANTENNA_2936 (.A(_09744_));
 sg13g2_antennanp ANTENNA_2937 (.A(_09744_));
 sg13g2_antennanp ANTENNA_2938 (.A(_09753_));
 sg13g2_antennanp ANTENNA_2939 (.A(_09798_));
 sg13g2_antennanp ANTENNA_2940 (.A(_09798_));
 sg13g2_antennanp ANTENNA_2941 (.A(_09954_));
 sg13g2_antennanp ANTENNA_2942 (.A(_09954_));
 sg13g2_antennanp ANTENNA_2943 (.A(_09954_));
 sg13g2_antennanp ANTENNA_2944 (.A(_09954_));
 sg13g2_antennanp ANTENNA_2945 (.A(_09954_));
 sg13g2_antennanp ANTENNA_2946 (.A(_09954_));
 sg13g2_antennanp ANTENNA_2947 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2948 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2949 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2950 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2951 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2952 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2953 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2954 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2955 (.A(_10054_));
 sg13g2_antennanp ANTENNA_2956 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2957 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2958 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2959 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2960 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2961 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2962 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2963 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2964 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2965 (.A(_10057_));
 sg13g2_antennanp ANTENNA_2966 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2967 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2968 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2969 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2970 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2971 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2972 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2973 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2974 (.A(_10107_));
 sg13g2_antennanp ANTENNA_2975 (.A(_10107_));
 sg13g2_antennanp ANTENNA_2976 (.A(_10107_));
 sg13g2_antennanp ANTENNA_2977 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2978 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2979 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2980 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2981 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2982 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2983 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2984 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2985 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2986 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2987 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2988 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2989 (.A(_10181_));
 sg13g2_antennanp ANTENNA_2990 (.A(_10386_));
 sg13g2_antennanp ANTENNA_2991 (.A(_10386_));
 sg13g2_antennanp ANTENNA_2992 (.A(_10572_));
 sg13g2_antennanp ANTENNA_2993 (.A(_10572_));
 sg13g2_antennanp ANTENNA_2994 (.A(_10572_));
 sg13g2_antennanp ANTENNA_2995 (.A(_10572_));
 sg13g2_antennanp ANTENNA_2996 (.A(_10703_));
 sg13g2_antennanp ANTENNA_2997 (.A(_10703_));
 sg13g2_antennanp ANTENNA_2998 (.A(_10703_));
 sg13g2_antennanp ANTENNA_2999 (.A(_10889_));
 sg13g2_antennanp ANTENNA_3000 (.A(_10889_));
 sg13g2_antennanp ANTENNA_3001 (.A(_10889_));
 sg13g2_antennanp ANTENNA_3002 (.A(_10889_));
 sg13g2_antennanp ANTENNA_3003 (.A(_10889_));
 sg13g2_antennanp ANTENNA_3004 (.A(_10889_));
 sg13g2_antennanp ANTENNA_3005 (.A(_11885_));
 sg13g2_antennanp ANTENNA_3006 (.A(_11885_));
 sg13g2_antennanp ANTENNA_3007 (.A(_11885_));
 sg13g2_antennanp ANTENNA_3008 (.A(_11970_));
 sg13g2_antennanp ANTENNA_3009 (.A(_11970_));
 sg13g2_antennanp ANTENNA_3010 (.A(_11970_));
 sg13g2_antennanp ANTENNA_3011 (.A(_12023_));
 sg13g2_antennanp ANTENNA_3012 (.A(_12023_));
 sg13g2_antennanp ANTENNA_3013 (.A(_12023_));
 sg13g2_antennanp ANTENNA_3014 (.A(_12023_));
 sg13g2_antennanp ANTENNA_3015 (.A(_12023_));
 sg13g2_antennanp ANTENNA_3016 (.A(_12023_));
 sg13g2_antennanp ANTENNA_3017 (.A(_12023_));
 sg13g2_antennanp ANTENNA_3018 (.A(_12023_));
 sg13g2_antennanp ANTENNA_3019 (.A(_12023_));
 sg13g2_antennanp ANTENNA_3020 (.A(_12046_));
 sg13g2_antennanp ANTENNA_3021 (.A(_12046_));
 sg13g2_antennanp ANTENNA_3022 (.A(_12046_));
 sg13g2_antennanp ANTENNA_3023 (.A(_12046_));
 sg13g2_antennanp ANTENNA_3024 (.A(_12046_));
 sg13g2_antennanp ANTENNA_3025 (.A(_12046_));
 sg13g2_antennanp ANTENNA_3026 (.A(_12046_));
 sg13g2_antennanp ANTENNA_3027 (.A(_12046_));
 sg13g2_antennanp ANTENNA_3028 (.A(_12046_));
 sg13g2_antennanp ANTENNA_3029 (.A(_12063_));
 sg13g2_antennanp ANTENNA_3030 (.A(_12063_));
 sg13g2_antennanp ANTENNA_3031 (.A(_12063_));
 sg13g2_antennanp ANTENNA_3032 (.A(_12063_));
 sg13g2_antennanp ANTENNA_3033 (.A(_12063_));
 sg13g2_antennanp ANTENNA_3034 (.A(_12063_));
 sg13g2_antennanp ANTENNA_3035 (.A(_12063_));
 sg13g2_antennanp ANTENNA_3036 (.A(_12063_));
 sg13g2_antennanp ANTENNA_3037 (.A(_12063_));
 sg13g2_antennanp ANTENNA_3038 (.A(_12096_));
 sg13g2_antennanp ANTENNA_3039 (.A(_12096_));
 sg13g2_antennanp ANTENNA_3040 (.A(_12096_));
 sg13g2_antennanp ANTENNA_3041 (.A(_12096_));
 sg13g2_antennanp ANTENNA_3042 (.A(_12096_));
 sg13g2_antennanp ANTENNA_3043 (.A(_12096_));
 sg13g2_antennanp ANTENNA_3044 (.A(_12096_));
 sg13g2_antennanp ANTENNA_3045 (.A(_12096_));
 sg13g2_antennanp ANTENNA_3046 (.A(_12096_));
 sg13g2_antennanp ANTENNA_3047 (.A(_12133_));
 sg13g2_antennanp ANTENNA_3048 (.A(_12133_));
 sg13g2_antennanp ANTENNA_3049 (.A(_12133_));
 sg13g2_antennanp ANTENNA_3050 (.A(_12133_));
 sg13g2_antennanp ANTENNA_3051 (.A(_12133_));
 sg13g2_antennanp ANTENNA_3052 (.A(_12133_));
 sg13g2_antennanp ANTENNA_3053 (.A(_12133_));
 sg13g2_antennanp ANTENNA_3054 (.A(_12133_));
 sg13g2_antennanp ANTENNA_3055 (.A(_12133_));
 sg13g2_antennanp ANTENNA_3056 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3057 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3058 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3059 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3060 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3061 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3062 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3063 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3064 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3065 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3066 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3067 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3068 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3069 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3070 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3071 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3072 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3073 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3074 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3075 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3076 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3077 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3078 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3079 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3080 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3081 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3082 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3083 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3084 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3085 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3086 (.A(_12156_));
 sg13g2_antennanp ANTENNA_3087 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_3088 (.A(r_reset));
 sg13g2_antennanp ANTENNA_3089 (.A(r_reset));
 sg13g2_antennanp ANTENNA_3090 (.A(r_reset));
 sg13g2_antennanp ANTENNA_3091 (.A(net1));
 sg13g2_antennanp ANTENNA_3092 (.A(net1));
 sg13g2_antennanp ANTENNA_3093 (.A(net1));
 sg13g2_antennanp ANTENNA_3094 (.A(net2));
 sg13g2_antennanp ANTENNA_3095 (.A(net2));
 sg13g2_antennanp ANTENNA_3096 (.A(net12));
 sg13g2_antennanp ANTENNA_3097 (.A(net12));
 sg13g2_antennanp ANTENNA_3098 (.A(net12));
 sg13g2_antennanp ANTENNA_3099 (.A(net19));
 sg13g2_antennanp ANTENNA_3100 (.A(net19));
 sg13g2_antennanp ANTENNA_3101 (.A(net20));
 sg13g2_antennanp ANTENNA_3102 (.A(net20));
 sg13g2_antennanp ANTENNA_3103 (.A(net153));
 sg13g2_antennanp ANTENNA_3104 (.A(net153));
 sg13g2_antennanp ANTENNA_3105 (.A(net153));
 sg13g2_antennanp ANTENNA_3106 (.A(net153));
 sg13g2_antennanp ANTENNA_3107 (.A(net153));
 sg13g2_antennanp ANTENNA_3108 (.A(net153));
 sg13g2_antennanp ANTENNA_3109 (.A(net153));
 sg13g2_antennanp ANTENNA_3110 (.A(net153));
 sg13g2_antennanp ANTENNA_3111 (.A(net153));
 sg13g2_antennanp ANTENNA_3112 (.A(net596));
 sg13g2_antennanp ANTENNA_3113 (.A(net596));
 sg13g2_antennanp ANTENNA_3114 (.A(net596));
 sg13g2_antennanp ANTENNA_3115 (.A(net596));
 sg13g2_antennanp ANTENNA_3116 (.A(net596));
 sg13g2_antennanp ANTENNA_3117 (.A(net596));
 sg13g2_antennanp ANTENNA_3118 (.A(net596));
 sg13g2_antennanp ANTENNA_3119 (.A(net596));
 sg13g2_antennanp ANTENNA_3120 (.A(net596));
 sg13g2_antennanp ANTENNA_3121 (.A(net618));
 sg13g2_antennanp ANTENNA_3122 (.A(net618));
 sg13g2_antennanp ANTENNA_3123 (.A(net618));
 sg13g2_antennanp ANTENNA_3124 (.A(net618));
 sg13g2_antennanp ANTENNA_3125 (.A(net618));
 sg13g2_antennanp ANTENNA_3126 (.A(net618));
 sg13g2_antennanp ANTENNA_3127 (.A(net618));
 sg13g2_antennanp ANTENNA_3128 (.A(net618));
 sg13g2_antennanp ANTENNA_3129 (.A(net618));
 sg13g2_antennanp ANTENNA_3130 (.A(net618));
 sg13g2_antennanp ANTENNA_3131 (.A(net618));
 sg13g2_antennanp ANTENNA_3132 (.A(net618));
 sg13g2_antennanp ANTENNA_3133 (.A(net618));
 sg13g2_antennanp ANTENNA_3134 (.A(net618));
 sg13g2_antennanp ANTENNA_3135 (.A(net618));
 sg13g2_antennanp ANTENNA_3136 (.A(net618));
 sg13g2_antennanp ANTENNA_3137 (.A(net618));
 sg13g2_antennanp ANTENNA_3138 (.A(net618));
 sg13g2_antennanp ANTENNA_3139 (.A(net618));
 sg13g2_antennanp ANTENNA_3140 (.A(net618));
 sg13g2_antennanp ANTENNA_3141 (.A(net618));
 sg13g2_antennanp ANTENNA_3142 (.A(net618));
 sg13g2_antennanp ANTENNA_3143 (.A(net618));
 sg13g2_antennanp ANTENNA_3144 (.A(net618));
 sg13g2_antennanp ANTENNA_3145 (.A(net618));
 sg13g2_antennanp ANTENNA_3146 (.A(net618));
 sg13g2_antennanp ANTENNA_3147 (.A(net618));
 sg13g2_antennanp ANTENNA_3148 (.A(net618));
 sg13g2_antennanp ANTENNA_3149 (.A(net618));
 sg13g2_antennanp ANTENNA_3150 (.A(net618));
 sg13g2_antennanp ANTENNA_3151 (.A(net618));
 sg13g2_antennanp ANTENNA_3152 (.A(net618));
 sg13g2_antennanp ANTENNA_3153 (.A(net618));
 sg13g2_antennanp ANTENNA_3154 (.A(net618));
 sg13g2_antennanp ANTENNA_3155 (.A(net618));
 sg13g2_antennanp ANTENNA_3156 (.A(net618));
 sg13g2_antennanp ANTENNA_3157 (.A(net618));
 sg13g2_antennanp ANTENNA_3158 (.A(net618));
 sg13g2_antennanp ANTENNA_3159 (.A(net618));
 sg13g2_antennanp ANTENNA_3160 (.A(net618));
 sg13g2_antennanp ANTENNA_3161 (.A(net618));
 sg13g2_antennanp ANTENNA_3162 (.A(net618));
 sg13g2_antennanp ANTENNA_3163 (.A(net618));
 sg13g2_antennanp ANTENNA_3164 (.A(net618));
 sg13g2_antennanp ANTENNA_3165 (.A(net618));
 sg13g2_antennanp ANTENNA_3166 (.A(net651));
 sg13g2_antennanp ANTENNA_3167 (.A(net651));
 sg13g2_antennanp ANTENNA_3168 (.A(net651));
 sg13g2_antennanp ANTENNA_3169 (.A(net651));
 sg13g2_antennanp ANTENNA_3170 (.A(net651));
 sg13g2_antennanp ANTENNA_3171 (.A(net651));
 sg13g2_antennanp ANTENNA_3172 (.A(net651));
 sg13g2_antennanp ANTENNA_3173 (.A(net651));
 sg13g2_antennanp ANTENNA_3174 (.A(net651));
 sg13g2_antennanp ANTENNA_3175 (.A(net651));
 sg13g2_antennanp ANTENNA_3176 (.A(net651));
 sg13g2_antennanp ANTENNA_3177 (.A(net651));
 sg13g2_antennanp ANTENNA_3178 (.A(net651));
 sg13g2_antennanp ANTENNA_3179 (.A(net651));
 sg13g2_antennanp ANTENNA_3180 (.A(net651));
 sg13g2_antennanp ANTENNA_3181 (.A(net651));
 sg13g2_antennanp ANTENNA_3182 (.A(net651));
 sg13g2_antennanp ANTENNA_3183 (.A(net651));
 sg13g2_antennanp ANTENNA_3184 (.A(net651));
 sg13g2_antennanp ANTENNA_3185 (.A(net651));
 sg13g2_antennanp ANTENNA_3186 (.A(net704));
 sg13g2_antennanp ANTENNA_3187 (.A(net704));
 sg13g2_antennanp ANTENNA_3188 (.A(net704));
 sg13g2_antennanp ANTENNA_3189 (.A(net704));
 sg13g2_antennanp ANTENNA_3190 (.A(net704));
 sg13g2_antennanp ANTENNA_3191 (.A(net704));
 sg13g2_antennanp ANTENNA_3192 (.A(net704));
 sg13g2_antennanp ANTENNA_3193 (.A(net704));
 sg13g2_antennanp ANTENNA_3194 (.A(net704));
 sg13g2_antennanp ANTENNA_3195 (.A(net860));
 sg13g2_antennanp ANTENNA_3196 (.A(net860));
 sg13g2_antennanp ANTENNA_3197 (.A(net860));
 sg13g2_antennanp ANTENNA_3198 (.A(net860));
 sg13g2_antennanp ANTENNA_3199 (.A(net860));
 sg13g2_antennanp ANTENNA_3200 (.A(net860));
 sg13g2_antennanp ANTENNA_3201 (.A(net860));
 sg13g2_antennanp ANTENNA_3202 (.A(net860));
 sg13g2_antennanp ANTENNA_3203 (.A(net860));
 sg13g2_antennanp ANTENNA_3204 (.A(net891));
 sg13g2_antennanp ANTENNA_3205 (.A(net891));
 sg13g2_antennanp ANTENNA_3206 (.A(net891));
 sg13g2_antennanp ANTENNA_3207 (.A(net891));
 sg13g2_antennanp ANTENNA_3208 (.A(net891));
 sg13g2_antennanp ANTENNA_3209 (.A(net891));
 sg13g2_antennanp ANTENNA_3210 (.A(net891));
 sg13g2_antennanp ANTENNA_3211 (.A(net891));
 sg13g2_antennanp ANTENNA_3212 (.A(net891));
 sg13g2_antennanp ANTENNA_3213 (.A(net899));
 sg13g2_antennanp ANTENNA_3214 (.A(net899));
 sg13g2_antennanp ANTENNA_3215 (.A(net899));
 sg13g2_antennanp ANTENNA_3216 (.A(net899));
 sg13g2_antennanp ANTENNA_3217 (.A(net899));
 sg13g2_antennanp ANTENNA_3218 (.A(net899));
 sg13g2_antennanp ANTENNA_3219 (.A(net899));
 sg13g2_antennanp ANTENNA_3220 (.A(net899));
 sg13g2_antennanp ANTENNA_3221 (.A(net899));
 sg13g2_antennanp ANTENNA_3222 (.A(net899));
 sg13g2_antennanp ANTENNA_3223 (.A(net899));
 sg13g2_antennanp ANTENNA_3224 (.A(net899));
 sg13g2_antennanp ANTENNA_3225 (.A(net899));
 sg13g2_antennanp ANTENNA_3226 (.A(net959));
 sg13g2_antennanp ANTENNA_3227 (.A(net959));
 sg13g2_antennanp ANTENNA_3228 (.A(net959));
 sg13g2_antennanp ANTENNA_3229 (.A(net959));
 sg13g2_antennanp ANTENNA_3230 (.A(net959));
 sg13g2_antennanp ANTENNA_3231 (.A(net959));
 sg13g2_antennanp ANTENNA_3232 (.A(net959));
 sg13g2_antennanp ANTENNA_3233 (.A(net959));
 sg13g2_antennanp ANTENNA_3234 (.A(net959));
 sg13g2_antennanp ANTENNA_3235 (.A(net970));
 sg13g2_antennanp ANTENNA_3236 (.A(net970));
 sg13g2_antennanp ANTENNA_3237 (.A(net970));
 sg13g2_antennanp ANTENNA_3238 (.A(net970));
 sg13g2_antennanp ANTENNA_3239 (.A(net970));
 sg13g2_antennanp ANTENNA_3240 (.A(net970));
 sg13g2_antennanp ANTENNA_3241 (.A(net970));
 sg13g2_antennanp ANTENNA_3242 (.A(net970));
 sg13g2_antennanp ANTENNA_3243 (.A(net971));
 sg13g2_antennanp ANTENNA_3244 (.A(net971));
 sg13g2_antennanp ANTENNA_3245 (.A(net971));
 sg13g2_antennanp ANTENNA_3246 (.A(net971));
 sg13g2_antennanp ANTENNA_3247 (.A(net971));
 sg13g2_antennanp ANTENNA_3248 (.A(net971));
 sg13g2_antennanp ANTENNA_3249 (.A(net971));
 sg13g2_antennanp ANTENNA_3250 (.A(net971));
 sg13g2_antennanp ANTENNA_3251 (.A(net971));
 sg13g2_antennanp ANTENNA_3252 (.A(net971));
 sg13g2_antennanp ANTENNA_3253 (.A(net971));
 sg13g2_antennanp ANTENNA_3254 (.A(net971));
 sg13g2_antennanp ANTENNA_3255 (.A(net971));
 sg13g2_antennanp ANTENNA_3256 (.A(net971));
 sg13g2_antennanp ANTENNA_3257 (.A(net971));
 sg13g2_antennanp ANTENNA_3258 (.A(net971));
 sg13g2_antennanp ANTENNA_3259 (.A(net971));
 sg13g2_antennanp ANTENNA_3260 (.A(net971));
 sg13g2_antennanp ANTENNA_3261 (.A(net971));
 sg13g2_antennanp ANTENNA_3262 (.A(net971));
 sg13g2_antennanp ANTENNA_3263 (.A(net972));
 sg13g2_antennanp ANTENNA_3264 (.A(net972));
 sg13g2_antennanp ANTENNA_3265 (.A(net972));
 sg13g2_antennanp ANTENNA_3266 (.A(net972));
 sg13g2_antennanp ANTENNA_3267 (.A(net972));
 sg13g2_antennanp ANTENNA_3268 (.A(net972));
 sg13g2_antennanp ANTENNA_3269 (.A(net972));
 sg13g2_antennanp ANTENNA_3270 (.A(net972));
 sg13g2_antennanp ANTENNA_3271 (.A(net972));
 sg13g2_antennanp ANTENNA_3272 (.A(net972));
 sg13g2_antennanp ANTENNA_3273 (.A(net972));
 sg13g2_antennanp ANTENNA_3274 (.A(net1000));
 sg13g2_antennanp ANTENNA_3275 (.A(net1000));
 sg13g2_antennanp ANTENNA_3276 (.A(net1000));
 sg13g2_antennanp ANTENNA_3277 (.A(net1000));
 sg13g2_antennanp ANTENNA_3278 (.A(net1000));
 sg13g2_antennanp ANTENNA_3279 (.A(net1000));
 sg13g2_antennanp ANTENNA_3280 (.A(net1000));
 sg13g2_antennanp ANTENNA_3281 (.A(net1000));
 sg13g2_antennanp ANTENNA_3282 (.A(net1043));
 sg13g2_antennanp ANTENNA_3283 (.A(net1043));
 sg13g2_antennanp ANTENNA_3284 (.A(net1043));
 sg13g2_antennanp ANTENNA_3285 (.A(net1043));
 sg13g2_antennanp ANTENNA_3286 (.A(net1043));
 sg13g2_antennanp ANTENNA_3287 (.A(net1043));
 sg13g2_antennanp ANTENNA_3288 (.A(net1043));
 sg13g2_antennanp ANTENNA_3289 (.A(net1043));
 sg13g2_antennanp ANTENNA_3290 (.A(net1043));
 sg13g2_antennanp ANTENNA_3291 (.A(net1043));
 sg13g2_antennanp ANTENNA_3292 (.A(net1043));
 sg13g2_antennanp ANTENNA_3293 (.A(net1043));
 sg13g2_antennanp ANTENNA_3294 (.A(net1053));
 sg13g2_antennanp ANTENNA_3295 (.A(net1053));
 sg13g2_antennanp ANTENNA_3296 (.A(net1053));
 sg13g2_antennanp ANTENNA_3297 (.A(net1053));
 sg13g2_antennanp ANTENNA_3298 (.A(net1053));
 sg13g2_antennanp ANTENNA_3299 (.A(net1053));
 sg13g2_antennanp ANTENNA_3300 (.A(net1053));
 sg13g2_antennanp ANTENNA_3301 (.A(net1053));
 sg13g2_antennanp ANTENNA_3302 (.A(net1053));
 sg13g2_antennanp ANTENNA_3303 (.A(net1053));
 sg13g2_antennanp ANTENNA_3304 (.A(net1053));
 sg13g2_antennanp ANTENNA_3305 (.A(net1053));
 sg13g2_antennanp ANTENNA_3306 (.A(net1053));
 sg13g2_antennanp ANTENNA_3307 (.A(net1053));
 sg13g2_antennanp ANTENNA_3308 (.A(net1053));
 sg13g2_antennanp ANTENNA_3309 (.A(net1072));
 sg13g2_antennanp ANTENNA_3310 (.A(net1072));
 sg13g2_antennanp ANTENNA_3311 (.A(net1072));
 sg13g2_antennanp ANTENNA_3312 (.A(net1072));
 sg13g2_antennanp ANTENNA_3313 (.A(net1072));
 sg13g2_antennanp ANTENNA_3314 (.A(net1072));
 sg13g2_antennanp ANTENNA_3315 (.A(net1072));
 sg13g2_antennanp ANTENNA_3316 (.A(net1072));
 sg13g2_antennanp ANTENNA_3317 (.A(net1072));
 sg13g2_antennanp ANTENNA_3318 (.A(net1104));
 sg13g2_antennanp ANTENNA_3319 (.A(net1104));
 sg13g2_antennanp ANTENNA_3320 (.A(net1104));
 sg13g2_antennanp ANTENNA_3321 (.A(net1104));
 sg13g2_antennanp ANTENNA_3322 (.A(net1104));
 sg13g2_antennanp ANTENNA_3323 (.A(net1104));
 sg13g2_antennanp ANTENNA_3324 (.A(net1104));
 sg13g2_antennanp ANTENNA_3325 (.A(net1104));
 sg13g2_antennanp ANTENNA_3326 (.A(net1104));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_4 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_85 ();
 sg13g2_decap_8 FILLER_0_92 ();
 sg13g2_decap_8 FILLER_0_99 ();
 sg13g2_decap_8 FILLER_0_106 ();
 sg13g2_decap_8 FILLER_0_113 ();
 sg13g2_decap_8 FILLER_0_120 ();
 sg13g2_decap_8 FILLER_0_127 ();
 sg13g2_decap_8 FILLER_0_134 ();
 sg13g2_decap_8 FILLER_0_141 ();
 sg13g2_decap_8 FILLER_0_148 ();
 sg13g2_decap_4 FILLER_0_155 ();
 sg13g2_fill_2 FILLER_0_159 ();
 sg13g2_decap_8 FILLER_0_187 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_decap_8 FILLER_0_208 ();
 sg13g2_decap_8 FILLER_0_215 ();
 sg13g2_decap_8 FILLER_0_222 ();
 sg13g2_decap_8 FILLER_0_255 ();
 sg13g2_decap_8 FILLER_0_262 ();
 sg13g2_decap_8 FILLER_0_269 ();
 sg13g2_decap_8 FILLER_0_276 ();
 sg13g2_decap_8 FILLER_0_283 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_decap_8 FILLER_0_297 ();
 sg13g2_decap_8 FILLER_0_304 ();
 sg13g2_fill_1 FILLER_0_311 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_4 FILLER_0_372 ();
 sg13g2_fill_2 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_4 FILLER_0_396 ();
 sg13g2_decap_8 FILLER_0_404 ();
 sg13g2_fill_2 FILLER_0_411 ();
 sg13g2_fill_1 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_418 ();
 sg13g2_decap_8 FILLER_0_425 ();
 sg13g2_decap_8 FILLER_0_432 ();
 sg13g2_decap_8 FILLER_0_439 ();
 sg13g2_decap_8 FILLER_0_446 ();
 sg13g2_decap_8 FILLER_0_453 ();
 sg13g2_fill_1 FILLER_0_460 ();
 sg13g2_decap_8 FILLER_0_487 ();
 sg13g2_decap_8 FILLER_0_494 ();
 sg13g2_decap_8 FILLER_0_501 ();
 sg13g2_decap_4 FILLER_0_508 ();
 sg13g2_fill_2 FILLER_0_512 ();
 sg13g2_decap_8 FILLER_0_540 ();
 sg13g2_decap_8 FILLER_0_547 ();
 sg13g2_decap_8 FILLER_0_554 ();
 sg13g2_decap_8 FILLER_0_561 ();
 sg13g2_decap_8 FILLER_0_568 ();
 sg13g2_decap_8 FILLER_0_575 ();
 sg13g2_decap_8 FILLER_0_582 ();
 sg13g2_decap_8 FILLER_0_589 ();
 sg13g2_decap_8 FILLER_0_596 ();
 sg13g2_fill_1 FILLER_0_603 ();
 sg13g2_decap_4 FILLER_0_614 ();
 sg13g2_decap_8 FILLER_0_628 ();
 sg13g2_decap_8 FILLER_0_635 ();
 sg13g2_decap_8 FILLER_0_642 ();
 sg13g2_decap_8 FILLER_0_649 ();
 sg13g2_decap_4 FILLER_0_656 ();
 sg13g2_decap_8 FILLER_0_670 ();
 sg13g2_decap_8 FILLER_0_677 ();
 sg13g2_decap_8 FILLER_0_684 ();
 sg13g2_decap_4 FILLER_0_691 ();
 sg13g2_fill_1 FILLER_0_695 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_fill_2 FILLER_0_707 ();
 sg13g2_fill_1 FILLER_0_709 ();
 sg13g2_decap_8 FILLER_0_724 ();
 sg13g2_decap_4 FILLER_0_731 ();
 sg13g2_fill_1 FILLER_0_735 ();
 sg13g2_decap_4 FILLER_0_740 ();
 sg13g2_fill_1 FILLER_0_744 ();
 sg13g2_decap_8 FILLER_0_765 ();
 sg13g2_decap_4 FILLER_0_772 ();
 sg13g2_decap_8 FILLER_0_786 ();
 sg13g2_fill_2 FILLER_0_793 ();
 sg13g2_fill_1 FILLER_0_795 ();
 sg13g2_decap_8 FILLER_0_806 ();
 sg13g2_decap_8 FILLER_0_813 ();
 sg13g2_decap_8 FILLER_0_820 ();
 sg13g2_decap_8 FILLER_0_827 ();
 sg13g2_decap_8 FILLER_0_834 ();
 sg13g2_decap_8 FILLER_0_841 ();
 sg13g2_decap_4 FILLER_0_848 ();
 sg13g2_fill_1 FILLER_0_862 ();
 sg13g2_decap_4 FILLER_0_889 ();
 sg13g2_fill_2 FILLER_0_893 ();
 sg13g2_decap_4 FILLER_0_921 ();
 sg13g2_fill_2 FILLER_0_925 ();
 sg13g2_decap_8 FILLER_0_953 ();
 sg13g2_decap_8 FILLER_0_960 ();
 sg13g2_decap_8 FILLER_0_967 ();
 sg13g2_decap_8 FILLER_0_974 ();
 sg13g2_fill_2 FILLER_0_981 ();
 sg13g2_fill_1 FILLER_0_983 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_decap_4 FILLER_0_1001 ();
 sg13g2_fill_1 FILLER_0_1005 ();
 sg13g2_decap_8 FILLER_0_1036 ();
 sg13g2_decap_4 FILLER_0_1043 ();
 sg13g2_fill_2 FILLER_0_1047 ();
 sg13g2_fill_2 FILLER_0_1053 ();
 sg13g2_fill_1 FILLER_0_1055 ();
 sg13g2_decap_8 FILLER_0_1064 ();
 sg13g2_decap_8 FILLER_0_1071 ();
 sg13g2_decap_8 FILLER_0_1078 ();
 sg13g2_decap_8 FILLER_0_1085 ();
 sg13g2_decap_8 FILLER_0_1092 ();
 sg13g2_decap_8 FILLER_0_1099 ();
 sg13g2_fill_2 FILLER_0_1106 ();
 sg13g2_decap_8 FILLER_0_1146 ();
 sg13g2_decap_8 FILLER_0_1153 ();
 sg13g2_fill_2 FILLER_0_1160 ();
 sg13g2_fill_1 FILLER_0_1162 ();
 sg13g2_decap_8 FILLER_0_1189 ();
 sg13g2_decap_8 FILLER_0_1222 ();
 sg13g2_decap_8 FILLER_0_1229 ();
 sg13g2_decap_8 FILLER_0_1262 ();
 sg13g2_decap_8 FILLER_0_1269 ();
 sg13g2_decap_4 FILLER_0_1276 ();
 sg13g2_fill_1 FILLER_0_1280 ();
 sg13g2_decap_8 FILLER_0_1311 ();
 sg13g2_decap_8 FILLER_0_1318 ();
 sg13g2_decap_8 FILLER_0_1351 ();
 sg13g2_decap_8 FILLER_0_1358 ();
 sg13g2_decap_8 FILLER_0_1365 ();
 sg13g2_fill_2 FILLER_0_1372 ();
 sg13g2_fill_1 FILLER_0_1410 ();
 sg13g2_decap_8 FILLER_0_1415 ();
 sg13g2_decap_8 FILLER_0_1422 ();
 sg13g2_decap_8 FILLER_0_1429 ();
 sg13g2_fill_1 FILLER_0_1436 ();
 sg13g2_decap_8 FILLER_0_1441 ();
 sg13g2_decap_8 FILLER_0_1448 ();
 sg13g2_decap_8 FILLER_0_1455 ();
 sg13g2_decap_8 FILLER_0_1462 ();
 sg13g2_decap_8 FILLER_0_1469 ();
 sg13g2_decap_8 FILLER_0_1476 ();
 sg13g2_fill_2 FILLER_0_1483 ();
 sg13g2_decap_8 FILLER_0_1511 ();
 sg13g2_decap_8 FILLER_0_1518 ();
 sg13g2_fill_2 FILLER_0_1525 ();
 sg13g2_fill_1 FILLER_0_1527 ();
 sg13g2_fill_2 FILLER_0_1532 ();
 sg13g2_decap_8 FILLER_0_1544 ();
 sg13g2_decap_8 FILLER_0_1551 ();
 sg13g2_decap_8 FILLER_0_1571 ();
 sg13g2_decap_8 FILLER_0_1578 ();
 sg13g2_decap_8 FILLER_0_1611 ();
 sg13g2_decap_4 FILLER_0_1618 ();
 sg13g2_fill_1 FILLER_0_1622 ();
 sg13g2_decap_8 FILLER_0_1653 ();
 sg13g2_decap_8 FILLER_0_1660 ();
 sg13g2_fill_2 FILLER_0_1667 ();
 sg13g2_fill_2 FILLER_0_1677 ();
 sg13g2_decap_8 FILLER_0_1683 ();
 sg13g2_decap_4 FILLER_0_1690 ();
 sg13g2_fill_1 FILLER_0_1698 ();
 sg13g2_decap_8 FILLER_0_1725 ();
 sg13g2_decap_8 FILLER_0_1732 ();
 sg13g2_decap_8 FILLER_0_1739 ();
 sg13g2_decap_4 FILLER_0_1746 ();
 sg13g2_fill_1 FILLER_0_1750 ();
 sg13g2_decap_8 FILLER_0_1755 ();
 sg13g2_decap_8 FILLER_0_1772 ();
 sg13g2_decap_4 FILLER_0_1779 ();
 sg13g2_fill_2 FILLER_0_1783 ();
 sg13g2_decap_8 FILLER_0_1811 ();
 sg13g2_decap_4 FILLER_0_1818 ();
 sg13g2_fill_2 FILLER_0_1822 ();
 sg13g2_decap_8 FILLER_0_1850 ();
 sg13g2_decap_8 FILLER_0_1857 ();
 sg13g2_fill_2 FILLER_0_1864 ();
 sg13g2_fill_1 FILLER_0_1866 ();
 sg13g2_decap_4 FILLER_0_1877 ();
 sg13g2_fill_2 FILLER_0_1911 ();
 sg13g2_fill_1 FILLER_0_1913 ();
 sg13g2_decap_8 FILLER_0_1927 ();
 sg13g2_decap_8 FILLER_0_1934 ();
 sg13g2_decap_8 FILLER_0_1941 ();
 sg13g2_decap_8 FILLER_0_1948 ();
 sg13g2_decap_8 FILLER_0_1955 ();
 sg13g2_decap_8 FILLER_0_1962 ();
 sg13g2_decap_8 FILLER_0_1973 ();
 sg13g2_fill_1 FILLER_0_1980 ();
 sg13g2_decap_8 FILLER_0_1991 ();
 sg13g2_decap_8 FILLER_0_1998 ();
 sg13g2_decap_8 FILLER_0_2005 ();
 sg13g2_decap_4 FILLER_0_2012 ();
 sg13g2_fill_2 FILLER_0_2016 ();
 sg13g2_decap_8 FILLER_0_2044 ();
 sg13g2_decap_4 FILLER_0_2051 ();
 sg13g2_fill_2 FILLER_0_2055 ();
 sg13g2_decap_4 FILLER_0_2061 ();
 sg13g2_fill_2 FILLER_0_2065 ();
 sg13g2_decap_8 FILLER_0_2080 ();
 sg13g2_decap_8 FILLER_0_2087 ();
 sg13g2_decap_4 FILLER_0_2094 ();
 sg13g2_fill_1 FILLER_0_2098 ();
 sg13g2_decap_8 FILLER_0_2103 ();
 sg13g2_decap_8 FILLER_0_2114 ();
 sg13g2_decap_8 FILLER_0_2121 ();
 sg13g2_fill_2 FILLER_0_2128 ();
 sg13g2_decap_4 FILLER_0_2170 ();
 sg13g2_decap_8 FILLER_0_2178 ();
 sg13g2_decap_8 FILLER_0_2185 ();
 sg13g2_decap_4 FILLER_0_2192 ();
 sg13g2_fill_1 FILLER_0_2196 ();
 sg13g2_decap_4 FILLER_0_2205 ();
 sg13g2_fill_2 FILLER_0_2209 ();
 sg13g2_decap_8 FILLER_0_2235 ();
 sg13g2_decap_8 FILLER_0_2242 ();
 sg13g2_decap_8 FILLER_0_2249 ();
 sg13g2_decap_8 FILLER_0_2256 ();
 sg13g2_decap_8 FILLER_0_2263 ();
 sg13g2_decap_8 FILLER_0_2270 ();
 sg13g2_decap_8 FILLER_0_2277 ();
 sg13g2_decap_8 FILLER_0_2284 ();
 sg13g2_decap_8 FILLER_0_2291 ();
 sg13g2_decap_8 FILLER_0_2298 ();
 sg13g2_decap_8 FILLER_0_2305 ();
 sg13g2_decap_8 FILLER_0_2312 ();
 sg13g2_decap_8 FILLER_0_2319 ();
 sg13g2_decap_8 FILLER_0_2326 ();
 sg13g2_decap_8 FILLER_0_2333 ();
 sg13g2_decap_8 FILLER_0_2340 ();
 sg13g2_decap_8 FILLER_0_2347 ();
 sg13g2_decap_8 FILLER_0_2354 ();
 sg13g2_decap_8 FILLER_0_2361 ();
 sg13g2_decap_8 FILLER_0_2368 ();
 sg13g2_decap_8 FILLER_0_2375 ();
 sg13g2_decap_8 FILLER_0_2382 ();
 sg13g2_decap_8 FILLER_0_2389 ();
 sg13g2_decap_8 FILLER_0_2396 ();
 sg13g2_decap_8 FILLER_0_2403 ();
 sg13g2_decap_8 FILLER_0_2410 ();
 sg13g2_decap_8 FILLER_0_2417 ();
 sg13g2_decap_8 FILLER_0_2424 ();
 sg13g2_decap_8 FILLER_0_2431 ();
 sg13g2_decap_8 FILLER_0_2438 ();
 sg13g2_decap_8 FILLER_0_2445 ();
 sg13g2_decap_8 FILLER_0_2452 ();
 sg13g2_decap_8 FILLER_0_2459 ();
 sg13g2_decap_8 FILLER_0_2466 ();
 sg13g2_decap_8 FILLER_0_2473 ();
 sg13g2_decap_8 FILLER_0_2480 ();
 sg13g2_decap_8 FILLER_0_2487 ();
 sg13g2_decap_8 FILLER_0_2494 ();
 sg13g2_decap_8 FILLER_0_2501 ();
 sg13g2_decap_8 FILLER_0_2508 ();
 sg13g2_decap_8 FILLER_0_2515 ();
 sg13g2_decap_8 FILLER_0_2522 ();
 sg13g2_decap_8 FILLER_0_2529 ();
 sg13g2_decap_8 FILLER_0_2536 ();
 sg13g2_decap_8 FILLER_0_2543 ();
 sg13g2_decap_8 FILLER_0_2550 ();
 sg13g2_decap_8 FILLER_0_2557 ();
 sg13g2_decap_8 FILLER_0_2564 ();
 sg13g2_decap_8 FILLER_0_2571 ();
 sg13g2_decap_8 FILLER_0_2578 ();
 sg13g2_decap_8 FILLER_0_2585 ();
 sg13g2_decap_8 FILLER_0_2592 ();
 sg13g2_decap_8 FILLER_0_2599 ();
 sg13g2_decap_8 FILLER_0_2606 ();
 sg13g2_decap_8 FILLER_0_2613 ();
 sg13g2_decap_8 FILLER_0_2620 ();
 sg13g2_decap_8 FILLER_0_2627 ();
 sg13g2_decap_8 FILLER_0_2634 ();
 sg13g2_decap_8 FILLER_0_2641 ();
 sg13g2_decap_8 FILLER_0_2648 ();
 sg13g2_decap_8 FILLER_0_2655 ();
 sg13g2_decap_8 FILLER_0_2662 ();
 sg13g2_fill_1 FILLER_0_2669 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_4 FILLER_1_70 ();
 sg13g2_fill_2 FILLER_1_104 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_fill_2 FILLER_1_126 ();
 sg13g2_fill_1 FILLER_1_128 ();
 sg13g2_decap_8 FILLER_1_159 ();
 sg13g2_fill_2 FILLER_1_166 ();
 sg13g2_decap_8 FILLER_1_209 ();
 sg13g2_decap_8 FILLER_1_216 ();
 sg13g2_fill_2 FILLER_1_223 ();
 sg13g2_decap_8 FILLER_1_263 ();
 sg13g2_decap_8 FILLER_1_270 ();
 sg13g2_decap_8 FILLER_1_277 ();
 sg13g2_decap_8 FILLER_1_284 ();
 sg13g2_decap_8 FILLER_1_291 ();
 sg13g2_decap_8 FILLER_1_298 ();
 sg13g2_fill_1 FILLER_1_344 ();
 sg13g2_fill_2 FILLER_1_391 ();
 sg13g2_fill_2 FILLER_1_398 ();
 sg13g2_fill_1 FILLER_1_404 ();
 sg13g2_fill_1 FILLER_1_457 ();
 sg13g2_decap_4 FILLER_1_462 ();
 sg13g2_fill_1 FILLER_1_475 ();
 sg13g2_decap_4 FILLER_1_502 ();
 sg13g2_fill_2 FILLER_1_506 ();
 sg13g2_decap_4 FILLER_1_538 ();
 sg13g2_fill_1 FILLER_1_542 ();
 sg13g2_decap_8 FILLER_1_547 ();
 sg13g2_decap_8 FILLER_1_554 ();
 sg13g2_decap_4 FILLER_1_561 ();
 sg13g2_fill_2 FILLER_1_578 ();
 sg13g2_decap_8 FILLER_1_584 ();
 sg13g2_fill_2 FILLER_1_591 ();
 sg13g2_fill_1 FILLER_1_593 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_fill_2 FILLER_1_637 ();
 sg13g2_fill_1 FILLER_1_639 ();
 sg13g2_fill_2 FILLER_1_676 ();
 sg13g2_decap_4 FILLER_1_724 ();
 sg13g2_fill_1 FILLER_1_728 ();
 sg13g2_fill_1 FILLER_1_765 ();
 sg13g2_fill_2 FILLER_1_770 ();
 sg13g2_fill_1 FILLER_1_802 ();
 sg13g2_fill_1 FILLER_1_829 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_4 FILLER_1_847 ();
 sg13g2_fill_2 FILLER_1_851 ();
 sg13g2_decap_4 FILLER_1_863 ();
 sg13g2_fill_2 FILLER_1_867 ();
 sg13g2_decap_4 FILLER_1_873 ();
 sg13g2_fill_2 FILLER_1_923 ();
 sg13g2_decap_4 FILLER_1_939 ();
 sg13g2_fill_1 FILLER_1_969 ();
 sg13g2_fill_1 FILLER_1_980 ();
 sg13g2_fill_1 FILLER_1_1033 ();
 sg13g2_fill_2 FILLER_1_1038 ();
 sg13g2_fill_1 FILLER_1_1040 ();
 sg13g2_decap_4 FILLER_1_1076 ();
 sg13g2_fill_2 FILLER_1_1088 ();
 sg13g2_fill_1 FILLER_1_1090 ();
 sg13g2_fill_1 FILLER_1_1126 ();
 sg13g2_decap_8 FILLER_1_1157 ();
 sg13g2_decap_4 FILLER_1_1164 ();
 sg13g2_fill_1 FILLER_1_1168 ();
 sg13g2_decap_4 FILLER_1_1173 ();
 sg13g2_fill_1 FILLER_1_1203 ();
 sg13g2_decap_4 FILLER_1_1234 ();
 sg13g2_fill_2 FILLER_1_1238 ();
 sg13g2_decap_8 FILLER_1_1275 ();
 sg13g2_fill_1 FILLER_1_1318 ();
 sg13g2_decap_8 FILLER_1_1355 ();
 sg13g2_fill_2 FILLER_1_1362 ();
 sg13g2_fill_1 FILLER_1_1364 ();
 sg13g2_decap_8 FILLER_1_1369 ();
 sg13g2_fill_2 FILLER_1_1376 ();
 sg13g2_fill_1 FILLER_1_1378 ();
 sg13g2_decap_8 FILLER_1_1461 ();
 sg13g2_decap_4 FILLER_1_1468 ();
 sg13g2_fill_2 FILLER_1_1498 ();
 sg13g2_fill_1 FILLER_1_1552 ();
 sg13g2_fill_1 FILLER_1_1566 ();
 sg13g2_fill_1 FILLER_1_1571 ();
 sg13g2_fill_1 FILLER_1_1598 ();
 sg13g2_decap_8 FILLER_1_1603 ();
 sg13g2_fill_2 FILLER_1_1610 ();
 sg13g2_fill_1 FILLER_1_1612 ();
 sg13g2_decap_8 FILLER_1_1617 ();
 sg13g2_decap_8 FILLER_1_1624 ();
 sg13g2_fill_2 FILLER_1_1631 ();
 sg13g2_decap_4 FILLER_1_1637 ();
 sg13g2_fill_2 FILLER_1_1641 ();
 sg13g2_decap_4 FILLER_1_1647 ();
 sg13g2_fill_2 FILLER_1_1655 ();
 sg13g2_fill_2 FILLER_1_1665 ();
 sg13g2_fill_1 FILLER_1_1667 ();
 sg13g2_decap_8 FILLER_1_1724 ();
 sg13g2_decap_8 FILLER_1_1731 ();
 sg13g2_decap_4 FILLER_1_1738 ();
 sg13g2_fill_2 FILLER_1_1742 ();
 sg13g2_fill_1 FILLER_1_1831 ();
 sg13g2_decap_8 FILLER_1_1836 ();
 sg13g2_fill_1 FILLER_1_1879 ();
 sg13g2_fill_1 FILLER_1_1901 ();
 sg13g2_fill_1 FILLER_1_1906 ();
 sg13g2_decap_8 FILLER_1_1928 ();
 sg13g2_fill_2 FILLER_1_1961 ();
 sg13g2_decap_8 FILLER_1_1997 ();
 sg13g2_decap_8 FILLER_1_2004 ();
 sg13g2_decap_8 FILLER_1_2011 ();
 sg13g2_decap_8 FILLER_1_2032 ();
 sg13g2_fill_2 FILLER_1_2039 ();
 sg13g2_decap_4 FILLER_1_2077 ();
 sg13g2_fill_1 FILLER_1_2081 ();
 sg13g2_decap_8 FILLER_1_2118 ();
 sg13g2_decap_8 FILLER_1_2125 ();
 sg13g2_decap_4 FILLER_1_2132 ();
 sg13g2_fill_1 FILLER_1_2136 ();
 sg13g2_decap_4 FILLER_1_2151 ();
 sg13g2_fill_2 FILLER_1_2155 ();
 sg13g2_decap_4 FILLER_1_2219 ();
 sg13g2_fill_1 FILLER_1_2223 ();
 sg13g2_decap_8 FILLER_1_2250 ();
 sg13g2_decap_8 FILLER_1_2257 ();
 sg13g2_decap_8 FILLER_1_2264 ();
 sg13g2_decap_8 FILLER_1_2271 ();
 sg13g2_decap_8 FILLER_1_2278 ();
 sg13g2_decap_8 FILLER_1_2285 ();
 sg13g2_decap_8 FILLER_1_2292 ();
 sg13g2_decap_8 FILLER_1_2299 ();
 sg13g2_decap_8 FILLER_1_2306 ();
 sg13g2_decap_8 FILLER_1_2313 ();
 sg13g2_decap_8 FILLER_1_2320 ();
 sg13g2_decap_8 FILLER_1_2327 ();
 sg13g2_decap_8 FILLER_1_2334 ();
 sg13g2_decap_8 FILLER_1_2341 ();
 sg13g2_decap_8 FILLER_1_2348 ();
 sg13g2_decap_8 FILLER_1_2355 ();
 sg13g2_decap_8 FILLER_1_2362 ();
 sg13g2_decap_8 FILLER_1_2369 ();
 sg13g2_decap_8 FILLER_1_2376 ();
 sg13g2_decap_8 FILLER_1_2383 ();
 sg13g2_decap_8 FILLER_1_2390 ();
 sg13g2_decap_8 FILLER_1_2397 ();
 sg13g2_decap_8 FILLER_1_2404 ();
 sg13g2_decap_8 FILLER_1_2411 ();
 sg13g2_decap_8 FILLER_1_2418 ();
 sg13g2_decap_8 FILLER_1_2425 ();
 sg13g2_decap_8 FILLER_1_2432 ();
 sg13g2_decap_8 FILLER_1_2439 ();
 sg13g2_decap_8 FILLER_1_2446 ();
 sg13g2_decap_8 FILLER_1_2453 ();
 sg13g2_decap_8 FILLER_1_2460 ();
 sg13g2_decap_8 FILLER_1_2467 ();
 sg13g2_decap_8 FILLER_1_2474 ();
 sg13g2_decap_8 FILLER_1_2481 ();
 sg13g2_decap_8 FILLER_1_2488 ();
 sg13g2_decap_8 FILLER_1_2495 ();
 sg13g2_decap_8 FILLER_1_2502 ();
 sg13g2_decap_8 FILLER_1_2509 ();
 sg13g2_decap_8 FILLER_1_2516 ();
 sg13g2_decap_8 FILLER_1_2523 ();
 sg13g2_decap_8 FILLER_1_2530 ();
 sg13g2_decap_8 FILLER_1_2537 ();
 sg13g2_decap_8 FILLER_1_2544 ();
 sg13g2_decap_8 FILLER_1_2551 ();
 sg13g2_decap_8 FILLER_1_2558 ();
 sg13g2_decap_8 FILLER_1_2565 ();
 sg13g2_decap_8 FILLER_1_2572 ();
 sg13g2_decap_8 FILLER_1_2579 ();
 sg13g2_decap_8 FILLER_1_2586 ();
 sg13g2_decap_8 FILLER_1_2593 ();
 sg13g2_decap_8 FILLER_1_2600 ();
 sg13g2_decap_8 FILLER_1_2607 ();
 sg13g2_decap_8 FILLER_1_2614 ();
 sg13g2_decap_8 FILLER_1_2621 ();
 sg13g2_decap_8 FILLER_1_2628 ();
 sg13g2_decap_8 FILLER_1_2635 ();
 sg13g2_decap_8 FILLER_1_2642 ();
 sg13g2_decap_8 FILLER_1_2649 ();
 sg13g2_decap_8 FILLER_1_2656 ();
 sg13g2_decap_8 FILLER_1_2663 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_fill_1 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_fill_2 FILLER_2_126 ();
 sg13g2_fill_2 FILLER_2_177 ();
 sg13g2_fill_1 FILLER_2_185 ();
 sg13g2_fill_2 FILLER_2_216 ();
 sg13g2_fill_1 FILLER_2_218 ();
 sg13g2_decap_8 FILLER_2_290 ();
 sg13g2_fill_2 FILLER_2_297 ();
 sg13g2_fill_1 FILLER_2_299 ();
 sg13g2_fill_1 FILLER_2_331 ();
 sg13g2_fill_2 FILLER_2_373 ();
 sg13g2_fill_1 FILLER_2_375 ();
 sg13g2_fill_1 FILLER_2_407 ();
 sg13g2_fill_1 FILLER_2_413 ();
 sg13g2_fill_2 FILLER_2_436 ();
 sg13g2_fill_1 FILLER_2_438 ();
 sg13g2_decap_8 FILLER_2_447 ();
 sg13g2_fill_2 FILLER_2_454 ();
 sg13g2_fill_1 FILLER_2_456 ();
 sg13g2_fill_1 FILLER_2_462 ();
 sg13g2_fill_2 FILLER_2_484 ();
 sg13g2_fill_2 FILLER_2_494 ();
 sg13g2_fill_1 FILLER_2_496 ();
 sg13g2_decap_4 FILLER_2_501 ();
 sg13g2_fill_1 FILLER_2_505 ();
 sg13g2_decap_8 FILLER_2_510 ();
 sg13g2_fill_1 FILLER_2_517 ();
 sg13g2_fill_2 FILLER_2_544 ();
 sg13g2_fill_1 FILLER_2_546 ();
 sg13g2_fill_2 FILLER_2_755 ();
 sg13g2_fill_1 FILLER_2_757 ();
 sg13g2_fill_1 FILLER_2_797 ();
 sg13g2_fill_1 FILLER_2_802 ();
 sg13g2_fill_2 FILLER_2_829 ();
 sg13g2_fill_1 FILLER_2_926 ();
 sg13g2_fill_2 FILLER_2_948 ();
 sg13g2_decap_8 FILLER_2_954 ();
 sg13g2_fill_2 FILLER_2_961 ();
 sg13g2_fill_1 FILLER_2_999 ();
 sg13g2_fill_1 FILLER_2_1009 ();
 sg13g2_fill_1 FILLER_2_1040 ();
 sg13g2_fill_1 FILLER_2_1046 ();
 sg13g2_fill_1 FILLER_2_1096 ();
 sg13g2_decap_4 FILLER_2_1123 ();
 sg13g2_fill_2 FILLER_2_1127 ();
 sg13g2_fill_2 FILLER_2_1134 ();
 sg13g2_fill_1 FILLER_2_1162 ();
 sg13g2_decap_4 FILLER_2_1190 ();
 sg13g2_fill_2 FILLER_2_1212 ();
 sg13g2_decap_8 FILLER_2_1218 ();
 sg13g2_fill_2 FILLER_2_1225 ();
 sg13g2_fill_1 FILLER_2_1227 ();
 sg13g2_fill_1 FILLER_2_1233 ();
 sg13g2_fill_1 FILLER_2_1238 ();
 sg13g2_fill_1 FILLER_2_1265 ();
 sg13g2_fill_1 FILLER_2_1287 ();
 sg13g2_fill_1 FILLER_2_1298 ();
 sg13g2_decap_8 FILLER_2_1303 ();
 sg13g2_fill_1 FILLER_2_1310 ();
 sg13g2_fill_2 FILLER_2_1357 ();
 sg13g2_fill_2 FILLER_2_1389 ();
 sg13g2_fill_1 FILLER_2_1401 ();
 sg13g2_fill_2 FILLER_2_1464 ();
 sg13g2_fill_1 FILLER_2_1496 ();
 sg13g2_fill_2 FILLER_2_1501 ();
 sg13g2_fill_1 FILLER_2_1521 ();
 sg13g2_fill_1 FILLER_2_1532 ();
 sg13g2_fill_1 FILLER_2_1536 ();
 sg13g2_fill_1 FILLER_2_1571 ();
 sg13g2_decap_8 FILLER_2_1594 ();
 sg13g2_fill_2 FILLER_2_1601 ();
 sg13g2_fill_1 FILLER_2_1603 ();
 sg13g2_fill_1 FILLER_2_1634 ();
 sg13g2_fill_2 FILLER_2_1661 ();
 sg13g2_fill_1 FILLER_2_1689 ();
 sg13g2_fill_2 FILLER_2_1695 ();
 sg13g2_fill_1 FILLER_2_1697 ();
 sg13g2_decap_8 FILLER_2_1725 ();
 sg13g2_fill_1 FILLER_2_1732 ();
 sg13g2_decap_8 FILLER_2_1769 ();
 sg13g2_decap_4 FILLER_2_1776 ();
 sg13g2_fill_2 FILLER_2_1780 ();
 sg13g2_decap_8 FILLER_2_1796 ();
 sg13g2_decap_4 FILLER_2_1803 ();
 sg13g2_fill_1 FILLER_2_1807 ();
 sg13g2_fill_2 FILLER_2_1844 ();
 sg13g2_fill_2 FILLER_2_1928 ();
 sg13g2_fill_1 FILLER_2_1930 ();
 sg13g2_fill_1 FILLER_2_1957 ();
 sg13g2_fill_2 FILLER_2_1984 ();
 sg13g2_fill_2 FILLER_2_2012 ();
 sg13g2_fill_1 FILLER_2_2014 ();
 sg13g2_fill_2 FILLER_2_2041 ();
 sg13g2_fill_1 FILLER_2_2043 ();
 sg13g2_fill_2 FILLER_2_2070 ();
 sg13g2_fill_2 FILLER_2_2098 ();
 sg13g2_fill_1 FILLER_2_2100 ();
 sg13g2_fill_1 FILLER_2_2127 ();
 sg13g2_fill_2 FILLER_2_2154 ();
 sg13g2_fill_1 FILLER_2_2156 ();
 sg13g2_decap_4 FILLER_2_2178 ();
 sg13g2_fill_1 FILLER_2_2182 ();
 sg13g2_fill_1 FILLER_2_2193 ();
 sg13g2_fill_2 FILLER_2_2204 ();
 sg13g2_decap_4 FILLER_2_2216 ();
 sg13g2_fill_1 FILLER_2_2220 ();
 sg13g2_decap_8 FILLER_2_2251 ();
 sg13g2_decap_8 FILLER_2_2258 ();
 sg13g2_decap_8 FILLER_2_2265 ();
 sg13g2_decap_8 FILLER_2_2272 ();
 sg13g2_decap_8 FILLER_2_2279 ();
 sg13g2_decap_8 FILLER_2_2286 ();
 sg13g2_decap_8 FILLER_2_2293 ();
 sg13g2_decap_8 FILLER_2_2300 ();
 sg13g2_decap_8 FILLER_2_2307 ();
 sg13g2_decap_8 FILLER_2_2314 ();
 sg13g2_decap_8 FILLER_2_2321 ();
 sg13g2_decap_8 FILLER_2_2328 ();
 sg13g2_decap_8 FILLER_2_2335 ();
 sg13g2_decap_8 FILLER_2_2342 ();
 sg13g2_decap_8 FILLER_2_2349 ();
 sg13g2_decap_8 FILLER_2_2356 ();
 sg13g2_decap_8 FILLER_2_2363 ();
 sg13g2_decap_8 FILLER_2_2370 ();
 sg13g2_decap_8 FILLER_2_2377 ();
 sg13g2_decap_8 FILLER_2_2384 ();
 sg13g2_decap_8 FILLER_2_2391 ();
 sg13g2_decap_8 FILLER_2_2398 ();
 sg13g2_decap_8 FILLER_2_2405 ();
 sg13g2_decap_8 FILLER_2_2412 ();
 sg13g2_decap_8 FILLER_2_2419 ();
 sg13g2_decap_8 FILLER_2_2426 ();
 sg13g2_decap_8 FILLER_2_2433 ();
 sg13g2_decap_8 FILLER_2_2440 ();
 sg13g2_decap_8 FILLER_2_2447 ();
 sg13g2_decap_8 FILLER_2_2454 ();
 sg13g2_decap_8 FILLER_2_2461 ();
 sg13g2_decap_8 FILLER_2_2468 ();
 sg13g2_decap_8 FILLER_2_2475 ();
 sg13g2_decap_8 FILLER_2_2482 ();
 sg13g2_decap_8 FILLER_2_2489 ();
 sg13g2_decap_8 FILLER_2_2496 ();
 sg13g2_decap_8 FILLER_2_2503 ();
 sg13g2_decap_8 FILLER_2_2510 ();
 sg13g2_decap_8 FILLER_2_2517 ();
 sg13g2_decap_8 FILLER_2_2524 ();
 sg13g2_decap_8 FILLER_2_2531 ();
 sg13g2_decap_8 FILLER_2_2538 ();
 sg13g2_decap_8 FILLER_2_2545 ();
 sg13g2_decap_8 FILLER_2_2552 ();
 sg13g2_decap_8 FILLER_2_2559 ();
 sg13g2_decap_8 FILLER_2_2566 ();
 sg13g2_decap_8 FILLER_2_2573 ();
 sg13g2_decap_8 FILLER_2_2580 ();
 sg13g2_decap_8 FILLER_2_2587 ();
 sg13g2_decap_8 FILLER_2_2594 ();
 sg13g2_decap_8 FILLER_2_2601 ();
 sg13g2_decap_8 FILLER_2_2608 ();
 sg13g2_decap_8 FILLER_2_2615 ();
 sg13g2_decap_8 FILLER_2_2622 ();
 sg13g2_decap_8 FILLER_2_2629 ();
 sg13g2_decap_8 FILLER_2_2636 ();
 sg13g2_decap_8 FILLER_2_2643 ();
 sg13g2_decap_8 FILLER_2_2650 ();
 sg13g2_decap_8 FILLER_2_2657 ();
 sg13g2_decap_4 FILLER_2_2664 ();
 sg13g2_fill_2 FILLER_2_2668 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_4 FILLER_3_56 ();
 sg13g2_fill_2 FILLER_3_60 ();
 sg13g2_fill_2 FILLER_3_74 ();
 sg13g2_fill_1 FILLER_3_80 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_decap_8 FILLER_3_123 ();
 sg13g2_decap_8 FILLER_3_130 ();
 sg13g2_decap_8 FILLER_3_137 ();
 sg13g2_fill_2 FILLER_3_172 ();
 sg13g2_fill_2 FILLER_3_182 ();
 sg13g2_fill_1 FILLER_3_187 ();
 sg13g2_fill_1 FILLER_3_192 ();
 sg13g2_fill_2 FILLER_3_197 ();
 sg13g2_decap_8 FILLER_3_206 ();
 sg13g2_fill_2 FILLER_3_217 ();
 sg13g2_fill_2 FILLER_3_248 ();
 sg13g2_fill_1 FILLER_3_263 ();
 sg13g2_fill_1 FILLER_3_339 ();
 sg13g2_fill_2 FILLER_3_353 ();
 sg13g2_fill_2 FILLER_3_401 ();
 sg13g2_fill_1 FILLER_3_413 ();
 sg13g2_fill_1 FILLER_3_444 ();
 sg13g2_fill_1 FILLER_3_463 ();
 sg13g2_fill_2 FILLER_3_472 ();
 sg13g2_decap_4 FILLER_3_500 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_fill_1 FILLER_3_547 ();
 sg13g2_decap_8 FILLER_3_582 ();
 sg13g2_fill_2 FILLER_3_589 ();
 sg13g2_fill_1 FILLER_3_591 ();
 sg13g2_decap_8 FILLER_3_675 ();
 sg13g2_fill_1 FILLER_3_682 ();
 sg13g2_decap_4 FILLER_3_687 ();
 sg13g2_fill_2 FILLER_3_727 ();
 sg13g2_decap_4 FILLER_3_816 ();
 sg13g2_fill_1 FILLER_3_820 ();
 sg13g2_fill_2 FILLER_3_857 ();
 sg13g2_decap_8 FILLER_3_880 ();
 sg13g2_decap_4 FILLER_3_887 ();
 sg13g2_fill_1 FILLER_3_891 ();
 sg13g2_decap_8 FILLER_3_914 ();
 sg13g2_decap_4 FILLER_3_921 ();
 sg13g2_decap_4 FILLER_3_946 ();
 sg13g2_fill_2 FILLER_3_950 ();
 sg13g2_fill_1 FILLER_3_962 ();
 sg13g2_fill_2 FILLER_3_1001 ();
 sg13g2_fill_1 FILLER_3_1003 ();
 sg13g2_fill_1 FILLER_3_1017 ();
 sg13g2_fill_2 FILLER_3_1070 ();
 sg13g2_fill_2 FILLER_3_1076 ();
 sg13g2_fill_2 FILLER_3_1082 ();
 sg13g2_fill_1 FILLER_3_1084 ();
 sg13g2_fill_2 FILLER_3_1125 ();
 sg13g2_fill_1 FILLER_3_1127 ();
 sg13g2_decap_8 FILLER_3_1163 ();
 sg13g2_decap_8 FILLER_3_1170 ();
 sg13g2_fill_2 FILLER_3_1177 ();
 sg13g2_fill_1 FILLER_3_1179 ();
 sg13g2_fill_2 FILLER_3_1184 ();
 sg13g2_fill_1 FILLER_3_1194 ();
 sg13g2_fill_1 FILLER_3_1200 ();
 sg13g2_decap_4 FILLER_3_1227 ();
 sg13g2_fill_1 FILLER_3_1231 ();
 sg13g2_fill_2 FILLER_3_1237 ();
 sg13g2_fill_1 FILLER_3_1239 ();
 sg13g2_decap_4 FILLER_3_1248 ();
 sg13g2_fill_2 FILLER_3_1313 ();
 sg13g2_fill_1 FILLER_3_1344 ();
 sg13g2_decap_8 FILLER_3_1349 ();
 sg13g2_fill_1 FILLER_3_1356 ();
 sg13g2_decap_8 FILLER_3_1367 ();
 sg13g2_decap_4 FILLER_3_1374 ();
 sg13g2_fill_2 FILLER_3_1378 ();
 sg13g2_fill_2 FILLER_3_1421 ();
 sg13g2_fill_2 FILLER_3_1433 ();
 sg13g2_fill_2 FILLER_3_1478 ();
 sg13g2_decap_8 FILLER_3_1484 ();
 sg13g2_fill_1 FILLER_3_1495 ();
 sg13g2_fill_2 FILLER_3_1500 ();
 sg13g2_fill_2 FILLER_3_1513 ();
 sg13g2_fill_2 FILLER_3_1526 ();
 sg13g2_fill_2 FILLER_3_1537 ();
 sg13g2_fill_1 FILLER_3_1585 ();
 sg13g2_fill_2 FILLER_3_1590 ();
 sg13g2_decap_4 FILLER_3_1598 ();
 sg13g2_fill_2 FILLER_3_1602 ();
 sg13g2_decap_8 FILLER_3_1607 ();
 sg13g2_fill_1 FILLER_3_1614 ();
 sg13g2_fill_1 FILLER_3_1630 ();
 sg13g2_fill_2 FILLER_3_1643 ();
 sg13g2_fill_2 FILLER_3_1692 ();
 sg13g2_fill_1 FILLER_3_1694 ();
 sg13g2_fill_1 FILLER_3_1732 ();
 sg13g2_fill_2 FILLER_3_1737 ();
 sg13g2_fill_1 FILLER_3_1739 ();
 sg13g2_fill_1 FILLER_3_1748 ();
 sg13g2_decap_8 FILLER_3_1785 ();
 sg13g2_fill_1 FILLER_3_1792 ();
 sg13g2_decap_4 FILLER_3_1807 ();
 sg13g2_fill_1 FILLER_3_1811 ();
 sg13g2_fill_1 FILLER_3_1822 ();
 sg13g2_fill_1 FILLER_3_1849 ();
 sg13g2_fill_1 FILLER_3_1854 ();
 sg13g2_fill_1 FILLER_3_1865 ();
 sg13g2_fill_2 FILLER_3_1892 ();
 sg13g2_fill_1 FILLER_3_1894 ();
 sg13g2_fill_1 FILLER_3_1909 ();
 sg13g2_fill_1 FILLER_3_1936 ();
 sg13g2_fill_2 FILLER_3_1951 ();
 sg13g2_fill_1 FILLER_3_1963 ();
 sg13g2_fill_1 FILLER_3_1968 ();
 sg13g2_fill_2 FILLER_3_1979 ();
 sg13g2_decap_4 FILLER_3_2033 ();
 sg13g2_fill_1 FILLER_3_2051 ();
 sg13g2_fill_1 FILLER_3_2078 ();
 sg13g2_decap_4 FILLER_3_2083 ();
 sg13g2_fill_1 FILLER_3_2087 ();
 sg13g2_fill_1 FILLER_3_2128 ();
 sg13g2_decap_4 FILLER_3_2193 ();
 sg13g2_fill_2 FILLER_3_2227 ();
 sg13g2_decap_8 FILLER_3_2255 ();
 sg13g2_decap_8 FILLER_3_2262 ();
 sg13g2_decap_8 FILLER_3_2269 ();
 sg13g2_decap_8 FILLER_3_2276 ();
 sg13g2_decap_8 FILLER_3_2283 ();
 sg13g2_decap_8 FILLER_3_2290 ();
 sg13g2_decap_8 FILLER_3_2297 ();
 sg13g2_decap_8 FILLER_3_2304 ();
 sg13g2_decap_8 FILLER_3_2311 ();
 sg13g2_decap_8 FILLER_3_2318 ();
 sg13g2_decap_8 FILLER_3_2325 ();
 sg13g2_decap_8 FILLER_3_2332 ();
 sg13g2_decap_8 FILLER_3_2339 ();
 sg13g2_decap_8 FILLER_3_2346 ();
 sg13g2_decap_8 FILLER_3_2353 ();
 sg13g2_decap_8 FILLER_3_2360 ();
 sg13g2_decap_8 FILLER_3_2367 ();
 sg13g2_decap_8 FILLER_3_2374 ();
 sg13g2_decap_8 FILLER_3_2381 ();
 sg13g2_decap_8 FILLER_3_2388 ();
 sg13g2_decap_8 FILLER_3_2395 ();
 sg13g2_decap_8 FILLER_3_2402 ();
 sg13g2_decap_8 FILLER_3_2409 ();
 sg13g2_decap_8 FILLER_3_2416 ();
 sg13g2_decap_8 FILLER_3_2423 ();
 sg13g2_decap_8 FILLER_3_2430 ();
 sg13g2_decap_8 FILLER_3_2437 ();
 sg13g2_decap_8 FILLER_3_2444 ();
 sg13g2_decap_8 FILLER_3_2451 ();
 sg13g2_decap_8 FILLER_3_2458 ();
 sg13g2_decap_8 FILLER_3_2465 ();
 sg13g2_decap_8 FILLER_3_2472 ();
 sg13g2_decap_8 FILLER_3_2479 ();
 sg13g2_decap_8 FILLER_3_2486 ();
 sg13g2_decap_8 FILLER_3_2493 ();
 sg13g2_decap_8 FILLER_3_2500 ();
 sg13g2_decap_8 FILLER_3_2507 ();
 sg13g2_decap_8 FILLER_3_2514 ();
 sg13g2_decap_8 FILLER_3_2521 ();
 sg13g2_decap_8 FILLER_3_2528 ();
 sg13g2_decap_8 FILLER_3_2535 ();
 sg13g2_decap_8 FILLER_3_2542 ();
 sg13g2_decap_8 FILLER_3_2549 ();
 sg13g2_decap_8 FILLER_3_2556 ();
 sg13g2_decap_8 FILLER_3_2563 ();
 sg13g2_decap_8 FILLER_3_2570 ();
 sg13g2_decap_8 FILLER_3_2577 ();
 sg13g2_decap_8 FILLER_3_2584 ();
 sg13g2_decap_8 FILLER_3_2591 ();
 sg13g2_decap_8 FILLER_3_2598 ();
 sg13g2_decap_8 FILLER_3_2605 ();
 sg13g2_decap_8 FILLER_3_2612 ();
 sg13g2_decap_8 FILLER_3_2619 ();
 sg13g2_decap_8 FILLER_3_2626 ();
 sg13g2_decap_8 FILLER_3_2633 ();
 sg13g2_decap_8 FILLER_3_2640 ();
 sg13g2_decap_8 FILLER_3_2647 ();
 sg13g2_decap_8 FILLER_3_2654 ();
 sg13g2_decap_8 FILLER_3_2661 ();
 sg13g2_fill_2 FILLER_3_2668 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_fill_2 FILLER_4_49 ();
 sg13g2_fill_1 FILLER_4_51 ();
 sg13g2_fill_2 FILLER_4_66 ();
 sg13g2_fill_2 FILLER_4_89 ();
 sg13g2_fill_1 FILLER_4_120 ();
 sg13g2_fill_2 FILLER_4_128 ();
 sg13g2_fill_1 FILLER_4_130 ();
 sg13g2_decap_8 FILLER_4_137 ();
 sg13g2_fill_2 FILLER_4_144 ();
 sg13g2_fill_1 FILLER_4_210 ();
 sg13g2_fill_1 FILLER_4_227 ();
 sg13g2_fill_1 FILLER_4_269 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_fill_2 FILLER_4_341 ();
 sg13g2_fill_1 FILLER_4_363 ();
 sg13g2_fill_2 FILLER_4_379 ();
 sg13g2_fill_1 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_444 ();
 sg13g2_fill_1 FILLER_4_453 ();
 sg13g2_fill_1 FILLER_4_480 ();
 sg13g2_decap_8 FILLER_4_485 ();
 sg13g2_decap_8 FILLER_4_492 ();
 sg13g2_decap_4 FILLER_4_499 ();
 sg13g2_fill_1 FILLER_4_523 ();
 sg13g2_decap_4 FILLER_4_529 ();
 sg13g2_fill_2 FILLER_4_533 ();
 sg13g2_fill_1 FILLER_4_554 ();
 sg13g2_fill_2 FILLER_4_560 ();
 sg13g2_fill_1 FILLER_4_562 ();
 sg13g2_fill_2 FILLER_4_593 ();
 sg13g2_fill_2 FILLER_4_612 ();
 sg13g2_fill_1 FILLER_4_614 ();
 sg13g2_decap_8 FILLER_4_625 ();
 sg13g2_fill_2 FILLER_4_632 ();
 sg13g2_fill_1 FILLER_4_638 ();
 sg13g2_fill_2 FILLER_4_657 ();
 sg13g2_fill_1 FILLER_4_659 ();
 sg13g2_decap_8 FILLER_4_664 ();
 sg13g2_fill_2 FILLER_4_671 ();
 sg13g2_decap_4 FILLER_4_694 ();
 sg13g2_fill_1 FILLER_4_698 ();
 sg13g2_fill_2 FILLER_4_703 ();
 sg13g2_fill_2 FILLER_4_726 ();
 sg13g2_decap_8 FILLER_4_766 ();
 sg13g2_decap_8 FILLER_4_773 ();
 sg13g2_fill_2 FILLER_4_780 ();
 sg13g2_decap_8 FILLER_4_786 ();
 sg13g2_decap_4 FILLER_4_793 ();
 sg13g2_fill_1 FILLER_4_797 ();
 sg13g2_decap_4 FILLER_4_808 ();
 sg13g2_fill_1 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_817 ();
 sg13g2_fill_2 FILLER_4_824 ();
 sg13g2_fill_1 FILLER_4_826 ();
 sg13g2_fill_1 FILLER_4_841 ();
 sg13g2_decap_8 FILLER_4_876 ();
 sg13g2_decap_4 FILLER_4_883 ();
 sg13g2_fill_2 FILLER_4_887 ();
 sg13g2_fill_1 FILLER_4_925 ();
 sg13g2_decap_4 FILLER_4_965 ();
 sg13g2_fill_1 FILLER_4_969 ();
 sg13g2_decap_8 FILLER_4_1001 ();
 sg13g2_decap_8 FILLER_4_1008 ();
 sg13g2_decap_4 FILLER_4_1015 ();
 sg13g2_fill_1 FILLER_4_1019 ();
 sg13g2_fill_2 FILLER_4_1025 ();
 sg13g2_decap_8 FILLER_4_1040 ();
 sg13g2_decap_4 FILLER_4_1047 ();
 sg13g2_fill_2 FILLER_4_1060 ();
 sg13g2_fill_2 FILLER_4_1124 ();
 sg13g2_fill_1 FILLER_4_1139 ();
 sg13g2_fill_2 FILLER_4_1169 ();
 sg13g2_fill_1 FILLER_4_1171 ();
 sg13g2_fill_2 FILLER_4_1193 ();
 sg13g2_fill_1 FILLER_4_1208 ();
 sg13g2_fill_1 FILLER_4_1240 ();
 sg13g2_fill_1 FILLER_4_1245 ();
 sg13g2_fill_1 FILLER_4_1250 ();
 sg13g2_fill_2 FILLER_4_1287 ();
 sg13g2_fill_1 FILLER_4_1289 ();
 sg13g2_decap_8 FILLER_4_1321 ();
 sg13g2_decap_8 FILLER_4_1328 ();
 sg13g2_decap_8 FILLER_4_1335 ();
 sg13g2_decap_8 FILLER_4_1342 ();
 sg13g2_decap_8 FILLER_4_1349 ();
 sg13g2_decap_8 FILLER_4_1356 ();
 sg13g2_fill_1 FILLER_4_1363 ();
 sg13g2_decap_4 FILLER_4_1421 ();
 sg13g2_fill_2 FILLER_4_1425 ();
 sg13g2_decap_8 FILLER_4_1473 ();
 sg13g2_decap_4 FILLER_4_1480 ();
 sg13g2_fill_2 FILLER_4_1484 ();
 sg13g2_fill_2 FILLER_4_1503 ();
 sg13g2_fill_1 FILLER_4_1515 ();
 sg13g2_fill_1 FILLER_4_1609 ();
 sg13g2_decap_8 FILLER_4_1644 ();
 sg13g2_decap_8 FILLER_4_1651 ();
 sg13g2_fill_1 FILLER_4_1673 ();
 sg13g2_fill_2 FILLER_4_1689 ();
 sg13g2_fill_1 FILLER_4_1691 ();
 sg13g2_decap_8 FILLER_4_1718 ();
 sg13g2_decap_8 FILLER_4_1725 ();
 sg13g2_decap_8 FILLER_4_1732 ();
 sg13g2_decap_8 FILLER_4_1739 ();
 sg13g2_fill_2 FILLER_4_1746 ();
 sg13g2_fill_1 FILLER_4_1748 ();
 sg13g2_fill_1 FILLER_4_1759 ();
 sg13g2_decap_4 FILLER_4_1786 ();
 sg13g2_decap_8 FILLER_4_1795 ();
 sg13g2_fill_2 FILLER_4_1802 ();
 sg13g2_fill_2 FILLER_4_1809 ();
 sg13g2_fill_1 FILLER_4_1811 ();
 sg13g2_decap_8 FILLER_4_1852 ();
 sg13g2_fill_2 FILLER_4_1859 ();
 sg13g2_decap_8 FILLER_4_1865 ();
 sg13g2_fill_2 FILLER_4_1872 ();
 sg13g2_decap_4 FILLER_4_1878 ();
 sg13g2_fill_2 FILLER_4_1882 ();
 sg13g2_fill_2 FILLER_4_1894 ();
 sg13g2_decap_4 FILLER_4_1906 ();
 sg13g2_fill_1 FILLER_4_1910 ();
 sg13g2_decap_4 FILLER_4_1921 ();
 sg13g2_decap_4 FILLER_4_1952 ();
 sg13g2_fill_2 FILLER_4_1956 ();
 sg13g2_decap_8 FILLER_4_1962 ();
 sg13g2_decap_8 FILLER_4_1969 ();
 sg13g2_fill_2 FILLER_4_1976 ();
 sg13g2_fill_2 FILLER_4_2019 ();
 sg13g2_decap_4 FILLER_4_2039 ();
 sg13g2_fill_1 FILLER_4_2043 ();
 sg13g2_decap_4 FILLER_4_2087 ();
 sg13g2_fill_1 FILLER_4_2091 ();
 sg13g2_decap_4 FILLER_4_2179 ();
 sg13g2_decap_8 FILLER_4_2199 ();
 sg13g2_fill_1 FILLER_4_2206 ();
 sg13g2_fill_2 FILLER_4_2232 ();
 sg13g2_fill_1 FILLER_4_2234 ();
 sg13g2_decap_4 FILLER_4_2239 ();
 sg13g2_decap_8 FILLER_4_2256 ();
 sg13g2_decap_8 FILLER_4_2263 ();
 sg13g2_decap_8 FILLER_4_2270 ();
 sg13g2_decap_8 FILLER_4_2277 ();
 sg13g2_decap_8 FILLER_4_2284 ();
 sg13g2_decap_8 FILLER_4_2291 ();
 sg13g2_decap_8 FILLER_4_2298 ();
 sg13g2_decap_8 FILLER_4_2305 ();
 sg13g2_decap_8 FILLER_4_2312 ();
 sg13g2_decap_8 FILLER_4_2319 ();
 sg13g2_decap_8 FILLER_4_2326 ();
 sg13g2_decap_8 FILLER_4_2333 ();
 sg13g2_decap_8 FILLER_4_2340 ();
 sg13g2_decap_8 FILLER_4_2347 ();
 sg13g2_decap_8 FILLER_4_2354 ();
 sg13g2_decap_8 FILLER_4_2361 ();
 sg13g2_decap_8 FILLER_4_2368 ();
 sg13g2_decap_8 FILLER_4_2375 ();
 sg13g2_decap_8 FILLER_4_2382 ();
 sg13g2_decap_8 FILLER_4_2389 ();
 sg13g2_decap_8 FILLER_4_2396 ();
 sg13g2_decap_8 FILLER_4_2403 ();
 sg13g2_decap_8 FILLER_4_2410 ();
 sg13g2_decap_8 FILLER_4_2417 ();
 sg13g2_decap_8 FILLER_4_2424 ();
 sg13g2_decap_8 FILLER_4_2431 ();
 sg13g2_decap_8 FILLER_4_2438 ();
 sg13g2_decap_8 FILLER_4_2445 ();
 sg13g2_decap_8 FILLER_4_2452 ();
 sg13g2_decap_8 FILLER_4_2459 ();
 sg13g2_decap_8 FILLER_4_2466 ();
 sg13g2_decap_8 FILLER_4_2473 ();
 sg13g2_decap_8 FILLER_4_2480 ();
 sg13g2_decap_8 FILLER_4_2487 ();
 sg13g2_decap_8 FILLER_4_2494 ();
 sg13g2_decap_8 FILLER_4_2501 ();
 sg13g2_decap_8 FILLER_4_2508 ();
 sg13g2_decap_8 FILLER_4_2515 ();
 sg13g2_decap_8 FILLER_4_2522 ();
 sg13g2_decap_8 FILLER_4_2529 ();
 sg13g2_decap_8 FILLER_4_2536 ();
 sg13g2_decap_8 FILLER_4_2543 ();
 sg13g2_decap_8 FILLER_4_2550 ();
 sg13g2_decap_8 FILLER_4_2557 ();
 sg13g2_decap_8 FILLER_4_2564 ();
 sg13g2_decap_8 FILLER_4_2571 ();
 sg13g2_decap_8 FILLER_4_2578 ();
 sg13g2_decap_8 FILLER_4_2585 ();
 sg13g2_decap_8 FILLER_4_2592 ();
 sg13g2_decap_8 FILLER_4_2599 ();
 sg13g2_decap_8 FILLER_4_2606 ();
 sg13g2_decap_8 FILLER_4_2613 ();
 sg13g2_decap_8 FILLER_4_2620 ();
 sg13g2_decap_8 FILLER_4_2627 ();
 sg13g2_decap_8 FILLER_4_2634 ();
 sg13g2_decap_8 FILLER_4_2641 ();
 sg13g2_decap_8 FILLER_4_2648 ();
 sg13g2_decap_8 FILLER_4_2655 ();
 sg13g2_decap_8 FILLER_4_2662 ();
 sg13g2_fill_1 FILLER_4_2669 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_fill_2 FILLER_5_42 ();
 sg13g2_fill_1 FILLER_5_44 ();
 sg13g2_fill_1 FILLER_5_82 ();
 sg13g2_fill_2 FILLER_5_91 ();
 sg13g2_fill_1 FILLER_5_186 ();
 sg13g2_fill_1 FILLER_5_200 ();
 sg13g2_fill_1 FILLER_5_205 ();
 sg13g2_fill_2 FILLER_5_214 ();
 sg13g2_fill_1 FILLER_5_225 ();
 sg13g2_fill_2 FILLER_5_234 ();
 sg13g2_fill_1 FILLER_5_236 ();
 sg13g2_fill_2 FILLER_5_250 ();
 sg13g2_decap_8 FILLER_5_257 ();
 sg13g2_fill_2 FILLER_5_264 ();
 sg13g2_fill_1 FILLER_5_275 ();
 sg13g2_decap_4 FILLER_5_281 ();
 sg13g2_fill_2 FILLER_5_285 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_4 FILLER_5_321 ();
 sg13g2_decap_4 FILLER_5_343 ();
 sg13g2_fill_1 FILLER_5_347 ();
 sg13g2_fill_1 FILLER_5_357 ();
 sg13g2_fill_2 FILLER_5_362 ();
 sg13g2_fill_2 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_fill_2 FILLER_5_393 ();
 sg13g2_fill_1 FILLER_5_395 ();
 sg13g2_fill_2 FILLER_5_409 ();
 sg13g2_fill_1 FILLER_5_425 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_fill_2 FILLER_5_514 ();
 sg13g2_fill_1 FILLER_5_516 ();
 sg13g2_fill_2 FILLER_5_534 ();
 sg13g2_fill_2 FILLER_5_540 ();
 sg13g2_decap_8 FILLER_5_582 ();
 sg13g2_decap_8 FILLER_5_589 ();
 sg13g2_fill_1 FILLER_5_596 ();
 sg13g2_decap_4 FILLER_5_601 ();
 sg13g2_fill_2 FILLER_5_605 ();
 sg13g2_decap_8 FILLER_5_611 ();
 sg13g2_decap_4 FILLER_5_618 ();
 sg13g2_fill_2 FILLER_5_622 ();
 sg13g2_decap_8 FILLER_5_650 ();
 sg13g2_decap_8 FILLER_5_657 ();
 sg13g2_decap_8 FILLER_5_664 ();
 sg13g2_decap_8 FILLER_5_671 ();
 sg13g2_decap_8 FILLER_5_678 ();
 sg13g2_decap_8 FILLER_5_685 ();
 sg13g2_decap_8 FILLER_5_692 ();
 sg13g2_decap_8 FILLER_5_699 ();
 sg13g2_decap_8 FILLER_5_706 ();
 sg13g2_decap_8 FILLER_5_713 ();
 sg13g2_decap_4 FILLER_5_720 ();
 sg13g2_fill_2 FILLER_5_724 ();
 sg13g2_decap_8 FILLER_5_766 ();
 sg13g2_fill_1 FILLER_5_773 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_4 FILLER_5_805 ();
 sg13g2_fill_1 FILLER_5_843 ();
 sg13g2_fill_2 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_856 ();
 sg13g2_decap_8 FILLER_5_883 ();
 sg13g2_decap_8 FILLER_5_890 ();
 sg13g2_decap_8 FILLER_5_897 ();
 sg13g2_fill_2 FILLER_5_904 ();
 sg13g2_fill_1 FILLER_5_906 ();
 sg13g2_decap_4 FILLER_5_911 ();
 sg13g2_fill_2 FILLER_5_915 ();
 sg13g2_decap_8 FILLER_5_957 ();
 sg13g2_decap_8 FILLER_5_964 ();
 sg13g2_decap_8 FILLER_5_971 ();
 sg13g2_fill_2 FILLER_5_978 ();
 sg13g2_fill_1 FILLER_5_980 ();
 sg13g2_decap_8 FILLER_5_991 ();
 sg13g2_decap_8 FILLER_5_998 ();
 sg13g2_decap_8 FILLER_5_1005 ();
 sg13g2_decap_8 FILLER_5_1012 ();
 sg13g2_decap_8 FILLER_5_1019 ();
 sg13g2_decap_8 FILLER_5_1026 ();
 sg13g2_fill_2 FILLER_5_1080 ();
 sg13g2_decap_8 FILLER_5_1087 ();
 sg13g2_fill_1 FILLER_5_1098 ();
 sg13g2_fill_2 FILLER_5_1103 ();
 sg13g2_fill_2 FILLER_5_1109 ();
 sg13g2_decap_8 FILLER_5_1132 ();
 sg13g2_decap_4 FILLER_5_1139 ();
 sg13g2_fill_1 FILLER_5_1143 ();
 sg13g2_decap_8 FILLER_5_1148 ();
 sg13g2_decap_8 FILLER_5_1155 ();
 sg13g2_decap_8 FILLER_5_1192 ();
 sg13g2_fill_1 FILLER_5_1199 ();
 sg13g2_fill_2 FILLER_5_1229 ();
 sg13g2_decap_4 FILLER_5_1235 ();
 sg13g2_decap_8 FILLER_5_1251 ();
 sg13g2_decap_4 FILLER_5_1262 ();
 sg13g2_fill_1 FILLER_5_1266 ();
 sg13g2_fill_2 FILLER_5_1281 ();
 sg13g2_fill_1 FILLER_5_1283 ();
 sg13g2_fill_2 FILLER_5_1288 ();
 sg13g2_fill_1 FILLER_5_1290 ();
 sg13g2_decap_8 FILLER_5_1320 ();
 sg13g2_fill_1 FILLER_5_1327 ();
 sg13g2_decap_8 FILLER_5_1338 ();
 sg13g2_fill_2 FILLER_5_1345 ();
 sg13g2_fill_1 FILLER_5_1347 ();
 sg13g2_decap_8 FILLER_5_1405 ();
 sg13g2_decap_8 FILLER_5_1412 ();
 sg13g2_decap_4 FILLER_5_1419 ();
 sg13g2_decap_4 FILLER_5_1427 ();
 sg13g2_fill_2 FILLER_5_1431 ();
 sg13g2_fill_2 FILLER_5_1438 ();
 sg13g2_fill_1 FILLER_5_1440 ();
 sg13g2_decap_8 FILLER_5_1466 ();
 sg13g2_fill_2 FILLER_5_1473 ();
 sg13g2_decap_8 FILLER_5_1479 ();
 sg13g2_decap_4 FILLER_5_1486 ();
 sg13g2_fill_1 FILLER_5_1598 ();
 sg13g2_fill_2 FILLER_5_1633 ();
 sg13g2_fill_1 FILLER_5_1635 ();
 sg13g2_decap_8 FILLER_5_1646 ();
 sg13g2_fill_2 FILLER_5_1653 ();
 sg13g2_fill_1 FILLER_5_1655 ();
 sg13g2_fill_1 FILLER_5_1666 ();
 sg13g2_fill_1 FILLER_5_1671 ();
 sg13g2_decap_4 FILLER_5_1693 ();
 sg13g2_fill_1 FILLER_5_1697 ();
 sg13g2_decap_8 FILLER_5_1702 ();
 sg13g2_decap_4 FILLER_5_1709 ();
 sg13g2_fill_1 FILLER_5_1713 ();
 sg13g2_decap_8 FILLER_5_1719 ();
 sg13g2_decap_8 FILLER_5_1730 ();
 sg13g2_decap_8 FILLER_5_1737 ();
 sg13g2_fill_2 FILLER_5_1760 ();
 sg13g2_fill_2 FILLER_5_1812 ();
 sg13g2_fill_1 FILLER_5_1814 ();
 sg13g2_decap_8 FILLER_5_1825 ();
 sg13g2_fill_2 FILLER_5_1832 ();
 sg13g2_fill_1 FILLER_5_1834 ();
 sg13g2_decap_8 FILLER_5_1839 ();
 sg13g2_decap_8 FILLER_5_1846 ();
 sg13g2_decap_8 FILLER_5_1853 ();
 sg13g2_decap_8 FILLER_5_1860 ();
 sg13g2_decap_4 FILLER_5_1867 ();
 sg13g2_fill_2 FILLER_5_1881 ();
 sg13g2_fill_1 FILLER_5_1883 ();
 sg13g2_decap_8 FILLER_5_1908 ();
 sg13g2_decap_8 FILLER_5_1915 ();
 sg13g2_decap_8 FILLER_5_1922 ();
 sg13g2_decap_8 FILLER_5_1929 ();
 sg13g2_fill_2 FILLER_5_1936 ();
 sg13g2_fill_1 FILLER_5_1938 ();
 sg13g2_decap_8 FILLER_5_1965 ();
 sg13g2_decap_8 FILLER_5_1972 ();
 sg13g2_decap_4 FILLER_5_1979 ();
 sg13g2_fill_2 FILLER_5_1991 ();
 sg13g2_fill_1 FILLER_5_2003 ();
 sg13g2_decap_8 FILLER_5_2008 ();
 sg13g2_decap_8 FILLER_5_2015 ();
 sg13g2_decap_4 FILLER_5_2022 ();
 sg13g2_fill_1 FILLER_5_2056 ();
 sg13g2_fill_1 FILLER_5_2061 ();
 sg13g2_fill_2 FILLER_5_2076 ();
 sg13g2_decap_8 FILLER_5_2086 ();
 sg13g2_decap_8 FILLER_5_2093 ();
 sg13g2_decap_4 FILLER_5_2110 ();
 sg13g2_decap_8 FILLER_5_2196 ();
 sg13g2_decap_8 FILLER_5_2203 ();
 sg13g2_decap_8 FILLER_5_2210 ();
 sg13g2_decap_8 FILLER_5_2217 ();
 sg13g2_decap_8 FILLER_5_2224 ();
 sg13g2_decap_8 FILLER_5_2231 ();
 sg13g2_decap_8 FILLER_5_2238 ();
 sg13g2_fill_1 FILLER_5_2245 ();
 sg13g2_decap_8 FILLER_5_2272 ();
 sg13g2_decap_8 FILLER_5_2279 ();
 sg13g2_decap_8 FILLER_5_2286 ();
 sg13g2_decap_8 FILLER_5_2293 ();
 sg13g2_decap_8 FILLER_5_2300 ();
 sg13g2_decap_8 FILLER_5_2307 ();
 sg13g2_decap_8 FILLER_5_2314 ();
 sg13g2_decap_8 FILLER_5_2321 ();
 sg13g2_decap_8 FILLER_5_2328 ();
 sg13g2_decap_8 FILLER_5_2335 ();
 sg13g2_decap_8 FILLER_5_2342 ();
 sg13g2_decap_8 FILLER_5_2349 ();
 sg13g2_decap_8 FILLER_5_2356 ();
 sg13g2_decap_8 FILLER_5_2363 ();
 sg13g2_decap_8 FILLER_5_2370 ();
 sg13g2_decap_8 FILLER_5_2377 ();
 sg13g2_decap_8 FILLER_5_2384 ();
 sg13g2_decap_8 FILLER_5_2391 ();
 sg13g2_decap_8 FILLER_5_2398 ();
 sg13g2_decap_8 FILLER_5_2405 ();
 sg13g2_decap_8 FILLER_5_2412 ();
 sg13g2_decap_8 FILLER_5_2419 ();
 sg13g2_decap_8 FILLER_5_2426 ();
 sg13g2_decap_8 FILLER_5_2433 ();
 sg13g2_decap_4 FILLER_5_2440 ();
 sg13g2_fill_1 FILLER_5_2444 ();
 sg13g2_decap_8 FILLER_5_2475 ();
 sg13g2_decap_8 FILLER_5_2482 ();
 sg13g2_decap_8 FILLER_5_2489 ();
 sg13g2_decap_8 FILLER_5_2496 ();
 sg13g2_decap_8 FILLER_5_2503 ();
 sg13g2_decap_8 FILLER_5_2510 ();
 sg13g2_decap_8 FILLER_5_2517 ();
 sg13g2_decap_8 FILLER_5_2524 ();
 sg13g2_decap_8 FILLER_5_2531 ();
 sg13g2_decap_8 FILLER_5_2538 ();
 sg13g2_decap_8 FILLER_5_2545 ();
 sg13g2_decap_8 FILLER_5_2552 ();
 sg13g2_decap_8 FILLER_5_2559 ();
 sg13g2_decap_8 FILLER_5_2566 ();
 sg13g2_decap_8 FILLER_5_2573 ();
 sg13g2_decap_8 FILLER_5_2580 ();
 sg13g2_decap_8 FILLER_5_2587 ();
 sg13g2_decap_8 FILLER_5_2594 ();
 sg13g2_decap_8 FILLER_5_2601 ();
 sg13g2_decap_8 FILLER_5_2608 ();
 sg13g2_decap_8 FILLER_5_2615 ();
 sg13g2_decap_8 FILLER_5_2622 ();
 sg13g2_decap_8 FILLER_5_2629 ();
 sg13g2_decap_8 FILLER_5_2636 ();
 sg13g2_decap_8 FILLER_5_2643 ();
 sg13g2_decap_8 FILLER_5_2650 ();
 sg13g2_decap_8 FILLER_5_2657 ();
 sg13g2_decap_4 FILLER_5_2664 ();
 sg13g2_fill_2 FILLER_5_2668 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_fill_1 FILLER_6_35 ();
 sg13g2_fill_2 FILLER_6_107 ();
 sg13g2_fill_1 FILLER_6_115 ();
 sg13g2_fill_2 FILLER_6_120 ();
 sg13g2_fill_1 FILLER_6_148 ();
 sg13g2_fill_1 FILLER_6_156 ();
 sg13g2_fill_1 FILLER_6_163 ();
 sg13g2_fill_1 FILLER_6_169 ();
 sg13g2_fill_1 FILLER_6_200 ();
 sg13g2_fill_1 FILLER_6_224 ();
 sg13g2_fill_2 FILLER_6_230 ();
 sg13g2_fill_1 FILLER_6_270 ();
 sg13g2_decap_8 FILLER_6_281 ();
 sg13g2_decap_8 FILLER_6_288 ();
 sg13g2_decap_8 FILLER_6_295 ();
 sg13g2_decap_8 FILLER_6_302 ();
 sg13g2_decap_8 FILLER_6_309 ();
 sg13g2_decap_8 FILLER_6_316 ();
 sg13g2_decap_8 FILLER_6_323 ();
 sg13g2_fill_2 FILLER_6_330 ();
 sg13g2_decap_8 FILLER_6_358 ();
 sg13g2_decap_8 FILLER_6_365 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_fill_2 FILLER_6_386 ();
 sg13g2_fill_1 FILLER_6_418 ();
 sg13g2_fill_2 FILLER_6_424 ();
 sg13g2_fill_2 FILLER_6_431 ();
 sg13g2_fill_2 FILLER_6_439 ();
 sg13g2_fill_1 FILLER_6_449 ();
 sg13g2_fill_1 FILLER_6_466 ();
 sg13g2_decap_4 FILLER_6_475 ();
 sg13g2_decap_8 FILLER_6_493 ();
 sg13g2_fill_2 FILLER_6_511 ();
 sg13g2_fill_1 FILLER_6_513 ();
 sg13g2_decap_4 FILLER_6_559 ();
 sg13g2_fill_1 FILLER_6_572 ();
 sg13g2_fill_2 FILLER_6_583 ();
 sg13g2_decap_8 FILLER_6_589 ();
 sg13g2_decap_8 FILLER_6_596 ();
 sg13g2_decap_8 FILLER_6_603 ();
 sg13g2_fill_1 FILLER_6_610 ();
 sg13g2_fill_2 FILLER_6_621 ();
 sg13g2_decap_4 FILLER_6_633 ();
 sg13g2_fill_2 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_649 ();
 sg13g2_decap_8 FILLER_6_656 ();
 sg13g2_decap_8 FILLER_6_663 ();
 sg13g2_fill_1 FILLER_6_670 ();
 sg13g2_fill_1 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_decap_8 FILLER_6_725 ();
 sg13g2_decap_4 FILLER_6_732 ();
 sg13g2_decap_4 FILLER_6_746 ();
 sg13g2_fill_2 FILLER_6_776 ();
 sg13g2_decap_4 FILLER_6_816 ();
 sg13g2_fill_1 FILLER_6_820 ();
 sg13g2_fill_1 FILLER_6_825 ();
 sg13g2_decap_8 FILLER_6_898 ();
 sg13g2_decap_8 FILLER_6_905 ();
 sg13g2_decap_4 FILLER_6_912 ();
 sg13g2_decap_4 FILLER_6_952 ();
 sg13g2_decap_4 FILLER_6_960 ();
 sg13g2_decap_8 FILLER_6_998 ();
 sg13g2_decap_8 FILLER_6_1005 ();
 sg13g2_decap_8 FILLER_6_1012 ();
 sg13g2_decap_8 FILLER_6_1019 ();
 sg13g2_decap_4 FILLER_6_1043 ();
 sg13g2_fill_1 FILLER_6_1047 ();
 sg13g2_decap_8 FILLER_6_1078 ();
 sg13g2_decap_8 FILLER_6_1110 ();
 sg13g2_fill_2 FILLER_6_1117 ();
 sg13g2_fill_1 FILLER_6_1119 ();
 sg13g2_decap_4 FILLER_6_1124 ();
 sg13g2_fill_2 FILLER_6_1128 ();
 sg13g2_fill_1 FILLER_6_1143 ();
 sg13g2_decap_8 FILLER_6_1149 ();
 sg13g2_decap_8 FILLER_6_1207 ();
 sg13g2_fill_2 FILLER_6_1214 ();
 sg13g2_fill_2 FILLER_6_1224 ();
 sg13g2_decap_8 FILLER_6_1230 ();
 sg13g2_fill_2 FILLER_6_1237 ();
 sg13g2_fill_1 FILLER_6_1239 ();
 sg13g2_fill_2 FILLER_6_1245 ();
 sg13g2_fill_1 FILLER_6_1247 ();
 sg13g2_fill_1 FILLER_6_1253 ();
 sg13g2_fill_2 FILLER_6_1258 ();
 sg13g2_decap_4 FILLER_6_1264 ();
 sg13g2_fill_1 FILLER_6_1268 ();
 sg13g2_decap_8 FILLER_6_1295 ();
 sg13g2_fill_1 FILLER_6_1302 ();
 sg13g2_decap_4 FILLER_6_1308 ();
 sg13g2_fill_1 FILLER_6_1312 ();
 sg13g2_fill_2 FILLER_6_1323 ();
 sg13g2_fill_2 FILLER_6_1335 ();
 sg13g2_fill_1 FILLER_6_1337 ();
 sg13g2_fill_1 FILLER_6_1364 ();
 sg13g2_fill_2 FILLER_6_1369 ();
 sg13g2_fill_1 FILLER_6_1371 ();
 sg13g2_decap_8 FILLER_6_1398 ();
 sg13g2_decap_8 FILLER_6_1405 ();
 sg13g2_fill_2 FILLER_6_1412 ();
 sg13g2_decap_8 FILLER_6_1435 ();
 sg13g2_decap_8 FILLER_6_1442 ();
 sg13g2_decap_8 FILLER_6_1449 ();
 sg13g2_decap_8 FILLER_6_1456 ();
 sg13g2_decap_4 FILLER_6_1463 ();
 sg13g2_fill_1 FILLER_6_1467 ();
 sg13g2_decap_4 FILLER_6_1494 ();
 sg13g2_fill_2 FILLER_6_1498 ();
 sg13g2_fill_1 FILLER_6_1508 ();
 sg13g2_fill_1 FILLER_6_1516 ();
 sg13g2_fill_1 FILLER_6_1536 ();
 sg13g2_fill_1 FILLER_6_1542 ();
 sg13g2_fill_1 FILLER_6_1547 ();
 sg13g2_fill_2 FILLER_6_1555 ();
 sg13g2_fill_1 FILLER_6_1561 ();
 sg13g2_fill_1 FILLER_6_1576 ();
 sg13g2_fill_1 FILLER_6_1582 ();
 sg13g2_fill_1 FILLER_6_1588 ();
 sg13g2_fill_2 FILLER_6_1598 ();
 sg13g2_fill_1 FILLER_6_1635 ();
 sg13g2_fill_2 FILLER_6_1641 ();
 sg13g2_fill_1 FILLER_6_1643 ();
 sg13g2_fill_2 FILLER_6_1654 ();
 sg13g2_fill_2 FILLER_6_1662 ();
 sg13g2_decap_4 FILLER_6_1683 ();
 sg13g2_decap_8 FILLER_6_1691 ();
 sg13g2_decap_8 FILLER_6_1698 ();
 sg13g2_decap_8 FILLER_6_1705 ();
 sg13g2_decap_8 FILLER_6_1712 ();
 sg13g2_fill_2 FILLER_6_1719 ();
 sg13g2_fill_1 FILLER_6_1721 ();
 sg13g2_fill_1 FILLER_6_1726 ();
 sg13g2_fill_2 FILLER_6_1753 ();
 sg13g2_fill_1 FILLER_6_1800 ();
 sg13g2_decap_8 FILLER_6_1806 ();
 sg13g2_fill_2 FILLER_6_1813 ();
 sg13g2_decap_8 FILLER_6_1820 ();
 sg13g2_decap_4 FILLER_6_1827 ();
 sg13g2_decap_4 FILLER_6_1857 ();
 sg13g2_decap_8 FILLER_6_1917 ();
 sg13g2_fill_2 FILLER_6_1960 ();
 sg13g2_fill_1 FILLER_6_1962 ();
 sg13g2_decap_4 FILLER_6_1985 ();
 sg13g2_fill_2 FILLER_6_2019 ();
 sg13g2_decap_4 FILLER_6_2031 ();
 sg13g2_fill_2 FILLER_6_2035 ();
 sg13g2_fill_2 FILLER_6_2058 ();
 sg13g2_fill_1 FILLER_6_2089 ();
 sg13g2_fill_1 FILLER_6_2094 ();
 sg13g2_decap_4 FILLER_6_2103 ();
 sg13g2_decap_4 FILLER_6_2167 ();
 sg13g2_decap_8 FILLER_6_2197 ();
 sg13g2_decap_8 FILLER_6_2204 ();
 sg13g2_decap_8 FILLER_6_2211 ();
 sg13g2_decap_8 FILLER_6_2218 ();
 sg13g2_fill_2 FILLER_6_2225 ();
 sg13g2_fill_1 FILLER_6_2237 ();
 sg13g2_fill_1 FILLER_6_2273 ();
 sg13g2_decap_8 FILLER_6_2278 ();
 sg13g2_decap_8 FILLER_6_2285 ();
 sg13g2_decap_8 FILLER_6_2292 ();
 sg13g2_decap_8 FILLER_6_2299 ();
 sg13g2_decap_8 FILLER_6_2306 ();
 sg13g2_decap_8 FILLER_6_2313 ();
 sg13g2_decap_8 FILLER_6_2320 ();
 sg13g2_decap_8 FILLER_6_2327 ();
 sg13g2_decap_8 FILLER_6_2334 ();
 sg13g2_decap_8 FILLER_6_2341 ();
 sg13g2_decap_8 FILLER_6_2348 ();
 sg13g2_decap_8 FILLER_6_2355 ();
 sg13g2_decap_8 FILLER_6_2362 ();
 sg13g2_decap_8 FILLER_6_2369 ();
 sg13g2_decap_8 FILLER_6_2376 ();
 sg13g2_decap_8 FILLER_6_2383 ();
 sg13g2_decap_8 FILLER_6_2390 ();
 sg13g2_fill_2 FILLER_6_2397 ();
 sg13g2_decap_4 FILLER_6_2425 ();
 sg13g2_fill_1 FILLER_6_2429 ();
 sg13g2_decap_4 FILLER_6_2434 ();
 sg13g2_fill_2 FILLER_6_2442 ();
 sg13g2_decap_8 FILLER_6_2483 ();
 sg13g2_decap_8 FILLER_6_2490 ();
 sg13g2_decap_4 FILLER_6_2497 ();
 sg13g2_fill_2 FILLER_6_2501 ();
 sg13g2_fill_2 FILLER_6_2533 ();
 sg13g2_decap_8 FILLER_6_2545 ();
 sg13g2_decap_8 FILLER_6_2552 ();
 sg13g2_decap_8 FILLER_6_2559 ();
 sg13g2_decap_8 FILLER_6_2566 ();
 sg13g2_decap_8 FILLER_6_2573 ();
 sg13g2_decap_8 FILLER_6_2580 ();
 sg13g2_decap_8 FILLER_6_2587 ();
 sg13g2_decap_8 FILLER_6_2594 ();
 sg13g2_decap_8 FILLER_6_2601 ();
 sg13g2_decap_8 FILLER_6_2608 ();
 sg13g2_decap_8 FILLER_6_2615 ();
 sg13g2_decap_8 FILLER_6_2622 ();
 sg13g2_decap_8 FILLER_6_2629 ();
 sg13g2_decap_8 FILLER_6_2636 ();
 sg13g2_decap_8 FILLER_6_2643 ();
 sg13g2_decap_8 FILLER_6_2650 ();
 sg13g2_decap_8 FILLER_6_2657 ();
 sg13g2_decap_4 FILLER_6_2664 ();
 sg13g2_fill_2 FILLER_6_2668 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_fill_1 FILLER_7_35 ();
 sg13g2_fill_2 FILLER_7_88 ();
 sg13g2_fill_1 FILLER_7_124 ();
 sg13g2_fill_1 FILLER_7_131 ();
 sg13g2_fill_1 FILLER_7_136 ();
 sg13g2_fill_1 FILLER_7_166 ();
 sg13g2_fill_1 FILLER_7_181 ();
 sg13g2_fill_1 FILLER_7_194 ();
 sg13g2_fill_1 FILLER_7_200 ();
 sg13g2_fill_1 FILLER_7_206 ();
 sg13g2_fill_2 FILLER_7_214 ();
 sg13g2_fill_1 FILLER_7_224 ();
 sg13g2_fill_1 FILLER_7_230 ();
 sg13g2_fill_1 FILLER_7_235 ();
 sg13g2_fill_2 FILLER_7_266 ();
 sg13g2_fill_1 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_279 ();
 sg13g2_decap_4 FILLER_7_286 ();
 sg13g2_decap_8 FILLER_7_320 ();
 sg13g2_decap_4 FILLER_7_327 ();
 sg13g2_fill_2 FILLER_7_396 ();
 sg13g2_fill_1 FILLER_7_398 ();
 sg13g2_fill_2 FILLER_7_429 ();
 sg13g2_fill_2 FILLER_7_448 ();
 sg13g2_fill_1 FILLER_7_467 ();
 sg13g2_fill_2 FILLER_7_542 ();
 sg13g2_fill_1 FILLER_7_544 ();
 sg13g2_decap_4 FILLER_7_549 ();
 sg13g2_fill_2 FILLER_7_566 ();
 sg13g2_fill_1 FILLER_7_604 ();
 sg13g2_fill_2 FILLER_7_661 ();
 sg13g2_fill_1 FILLER_7_663 ();
 sg13g2_fill_1 FILLER_7_674 ();
 sg13g2_fill_2 FILLER_7_726 ();
 sg13g2_fill_1 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_764 ();
 sg13g2_fill_1 FILLER_7_771 ();
 sg13g2_decap_8 FILLER_7_793 ();
 sg13g2_decap_4 FILLER_7_800 ();
 sg13g2_fill_1 FILLER_7_804 ();
 sg13g2_fill_2 FILLER_7_841 ();
 sg13g2_fill_1 FILLER_7_864 ();
 sg13g2_fill_1 FILLER_7_873 ();
 sg13g2_fill_1 FILLER_7_878 ();
 sg13g2_fill_2 FILLER_7_905 ();
 sg13g2_fill_2 FILLER_7_912 ();
 sg13g2_fill_2 FILLER_7_927 ();
 sg13g2_fill_1 FILLER_7_929 ();
 sg13g2_decap_8 FILLER_7_944 ();
 sg13g2_decap_8 FILLER_7_951 ();
 sg13g2_decap_8 FILLER_7_958 ();
 sg13g2_fill_2 FILLER_7_965 ();
 sg13g2_fill_1 FILLER_7_985 ();
 sg13g2_fill_2 FILLER_7_1012 ();
 sg13g2_fill_1 FILLER_7_1019 ();
 sg13g2_fill_2 FILLER_7_1046 ();
 sg13g2_fill_1 FILLER_7_1074 ();
 sg13g2_decap_4 FILLER_7_1101 ();
 sg13g2_decap_8 FILLER_7_1109 ();
 sg13g2_fill_2 FILLER_7_1116 ();
 sg13g2_fill_1 FILLER_7_1118 ();
 sg13g2_fill_2 FILLER_7_1124 ();
 sg13g2_fill_1 FILLER_7_1126 ();
 sg13g2_fill_1 FILLER_7_1153 ();
 sg13g2_decap_8 FILLER_7_1158 ();
 sg13g2_fill_2 FILLER_7_1165 ();
 sg13g2_fill_2 FILLER_7_1171 ();
 sg13g2_fill_1 FILLER_7_1178 ();
 sg13g2_decap_8 FILLER_7_1226 ();
 sg13g2_fill_1 FILLER_7_1233 ();
 sg13g2_decap_8 FILLER_7_1273 ();
 sg13g2_decap_8 FILLER_7_1280 ();
 sg13g2_decap_4 FILLER_7_1287 ();
 sg13g2_decap_8 FILLER_7_1295 ();
 sg13g2_fill_1 FILLER_7_1302 ();
 sg13g2_fill_2 FILLER_7_1334 ();
 sg13g2_fill_1 FILLER_7_1336 ();
 sg13g2_decap_4 FILLER_7_1363 ();
 sg13g2_fill_1 FILLER_7_1367 ();
 sg13g2_fill_2 FILLER_7_1378 ();
 sg13g2_fill_1 FILLER_7_1384 ();
 sg13g2_fill_2 FILLER_7_1389 ();
 sg13g2_fill_1 FILLER_7_1391 ();
 sg13g2_fill_2 FILLER_7_1431 ();
 sg13g2_decap_8 FILLER_7_1437 ();
 sg13g2_decap_8 FILLER_7_1444 ();
 sg13g2_decap_8 FILLER_7_1451 ();
 sg13g2_decap_4 FILLER_7_1458 ();
 sg13g2_fill_1 FILLER_7_1462 ();
 sg13g2_decap_8 FILLER_7_1467 ();
 sg13g2_decap_8 FILLER_7_1474 ();
 sg13g2_decap_8 FILLER_7_1481 ();
 sg13g2_fill_2 FILLER_7_1488 ();
 sg13g2_fill_1 FILLER_7_1501 ();
 sg13g2_fill_2 FILLER_7_1508 ();
 sg13g2_fill_1 FILLER_7_1520 ();
 sg13g2_fill_1 FILLER_7_1527 ();
 sg13g2_fill_1 FILLER_7_1534 ();
 sg13g2_fill_2 FILLER_7_1550 ();
 sg13g2_fill_1 FILLER_7_1556 ();
 sg13g2_fill_1 FILLER_7_1581 ();
 sg13g2_fill_1 FILLER_7_1591 ();
 sg13g2_fill_2 FILLER_7_1622 ();
 sg13g2_fill_2 FILLER_7_1697 ();
 sg13g2_decap_4 FILLER_7_1720 ();
 sg13g2_fill_1 FILLER_7_1724 ();
 sg13g2_fill_1 FILLER_7_1754 ();
 sg13g2_decap_8 FILLER_7_1785 ();
 sg13g2_decap_8 FILLER_7_1792 ();
 sg13g2_fill_1 FILLER_7_1799 ();
 sg13g2_decap_4 FILLER_7_1804 ();
 sg13g2_fill_2 FILLER_7_1808 ();
 sg13g2_fill_2 FILLER_7_1814 ();
 sg13g2_decap_4 FILLER_7_1820 ();
 sg13g2_fill_2 FILLER_7_1838 ();
 sg13g2_fill_1 FILLER_7_1840 ();
 sg13g2_fill_2 FILLER_7_1893 ();
 sg13g2_fill_1 FILLER_7_1895 ();
 sg13g2_decap_4 FILLER_7_1922 ();
 sg13g2_fill_1 FILLER_7_1926 ();
 sg13g2_decap_8 FILLER_7_1957 ();
 sg13g2_fill_2 FILLER_7_1964 ();
 sg13g2_fill_1 FILLER_7_1992 ();
 sg13g2_fill_1 FILLER_7_2014 ();
 sg13g2_fill_1 FILLER_7_2019 ();
 sg13g2_fill_2 FILLER_7_2046 ();
 sg13g2_fill_2 FILLER_7_2084 ();
 sg13g2_fill_1 FILLER_7_2090 ();
 sg13g2_decap_8 FILLER_7_2188 ();
 sg13g2_fill_1 FILLER_7_2195 ();
 sg13g2_decap_8 FILLER_7_2284 ();
 sg13g2_decap_8 FILLER_7_2291 ();
 sg13g2_decap_8 FILLER_7_2298 ();
 sg13g2_decap_8 FILLER_7_2305 ();
 sg13g2_decap_8 FILLER_7_2312 ();
 sg13g2_decap_8 FILLER_7_2319 ();
 sg13g2_decap_8 FILLER_7_2326 ();
 sg13g2_decap_8 FILLER_7_2333 ();
 sg13g2_decap_8 FILLER_7_2340 ();
 sg13g2_decap_8 FILLER_7_2347 ();
 sg13g2_decap_8 FILLER_7_2354 ();
 sg13g2_decap_8 FILLER_7_2361 ();
 sg13g2_decap_8 FILLER_7_2368 ();
 sg13g2_decap_8 FILLER_7_2375 ();
 sg13g2_decap_8 FILLER_7_2382 ();
 sg13g2_decap_8 FILLER_7_2389 ();
 sg13g2_fill_2 FILLER_7_2396 ();
 sg13g2_fill_2 FILLER_7_2456 ();
 sg13g2_fill_1 FILLER_7_2458 ();
 sg13g2_decap_8 FILLER_7_2485 ();
 sg13g2_decap_8 FILLER_7_2492 ();
 sg13g2_decap_8 FILLER_7_2499 ();
 sg13g2_fill_2 FILLER_7_2506 ();
 sg13g2_fill_1 FILLER_7_2508 ();
 sg13g2_decap_8 FILLER_7_2552 ();
 sg13g2_fill_2 FILLER_7_2559 ();
 sg13g2_fill_1 FILLER_7_2561 ();
 sg13g2_decap_4 FILLER_7_2588 ();
 sg13g2_decap_8 FILLER_7_2596 ();
 sg13g2_decap_8 FILLER_7_2603 ();
 sg13g2_decap_8 FILLER_7_2610 ();
 sg13g2_decap_8 FILLER_7_2617 ();
 sg13g2_decap_8 FILLER_7_2624 ();
 sg13g2_decap_8 FILLER_7_2631 ();
 sg13g2_decap_8 FILLER_7_2638 ();
 sg13g2_decap_8 FILLER_7_2645 ();
 sg13g2_decap_8 FILLER_7_2652 ();
 sg13g2_decap_8 FILLER_7_2659 ();
 sg13g2_decap_4 FILLER_7_2666 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_fill_1 FILLER_8_35 ();
 sg13g2_fill_1 FILLER_8_48 ();
 sg13g2_fill_2 FILLER_8_53 ();
 sg13g2_fill_2 FILLER_8_70 ();
 sg13g2_fill_1 FILLER_8_94 ();
 sg13g2_fill_1 FILLER_8_130 ();
 sg13g2_fill_2 FILLER_8_149 ();
 sg13g2_fill_2 FILLER_8_159 ();
 sg13g2_fill_1 FILLER_8_212 ();
 sg13g2_fill_2 FILLER_8_227 ();
 sg13g2_fill_2 FILLER_8_233 ();
 sg13g2_fill_1 FILLER_8_235 ();
 sg13g2_fill_2 FILLER_8_241 ();
 sg13g2_fill_1 FILLER_8_243 ();
 sg13g2_fill_1 FILLER_8_290 ();
 sg13g2_fill_1 FILLER_8_295 ();
 sg13g2_fill_2 FILLER_8_300 ();
 sg13g2_decap_4 FILLER_8_307 ();
 sg13g2_fill_1 FILLER_8_345 ();
 sg13g2_fill_2 FILLER_8_350 ();
 sg13g2_fill_1 FILLER_8_352 ();
 sg13g2_fill_2 FILLER_8_378 ();
 sg13g2_fill_1 FILLER_8_380 ();
 sg13g2_fill_2 FILLER_8_391 ();
 sg13g2_decap_4 FILLER_8_398 ();
 sg13g2_fill_2 FILLER_8_402 ();
 sg13g2_fill_2 FILLER_8_443 ();
 sg13g2_fill_2 FILLER_8_521 ();
 sg13g2_fill_1 FILLER_8_527 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_fill_2 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_552 ();
 sg13g2_fill_1 FILLER_8_559 ();
 sg13g2_fill_2 FILLER_8_568 ();
 sg13g2_decap_4 FILLER_8_596 ();
 sg13g2_fill_2 FILLER_8_600 ();
 sg13g2_fill_2 FILLER_8_628 ();
 sg13g2_fill_2 FILLER_8_655 ();
 sg13g2_fill_2 FILLER_8_687 ();
 sg13g2_fill_1 FILLER_8_689 ();
 sg13g2_fill_2 FILLER_8_747 ();
 sg13g2_fill_1 FILLER_8_749 ();
 sg13g2_fill_2 FILLER_8_754 ();
 sg13g2_fill_2 FILLER_8_792 ();
 sg13g2_fill_1 FILLER_8_794 ();
 sg13g2_decap_4 FILLER_8_816 ();
 sg13g2_fill_2 FILLER_8_820 ();
 sg13g2_decap_4 FILLER_8_861 ();
 sg13g2_fill_2 FILLER_8_865 ();
 sg13g2_decap_8 FILLER_8_888 ();
 sg13g2_decap_8 FILLER_8_895 ();
 sg13g2_decap_4 FILLER_8_902 ();
 sg13g2_fill_2 FILLER_8_906 ();
 sg13g2_decap_4 FILLER_8_955 ();
 sg13g2_fill_2 FILLER_8_959 ();
 sg13g2_fill_2 FILLER_8_1062 ();
 sg13g2_decap_4 FILLER_8_1068 ();
 sg13g2_fill_2 FILLER_8_1072 ();
 sg13g2_fill_1 FILLER_8_1105 ();
 sg13g2_fill_1 FILLER_8_1140 ();
 sg13g2_fill_1 FILLER_8_1171 ();
 sg13g2_decap_4 FILLER_8_1218 ();
 sg13g2_fill_2 FILLER_8_1252 ();
 sg13g2_fill_1 FILLER_8_1254 ();
 sg13g2_fill_1 FILLER_8_1294 ();
 sg13g2_decap_8 FILLER_8_1355 ();
 sg13g2_fill_2 FILLER_8_1362 ();
 sg13g2_fill_1 FILLER_8_1364 ();
 sg13g2_decap_4 FILLER_8_1370 ();
 sg13g2_fill_1 FILLER_8_1374 ();
 sg13g2_decap_8 FILLER_8_1380 ();
 sg13g2_decap_4 FILLER_8_1387 ();
 sg13g2_fill_1 FILLER_8_1391 ();
 sg13g2_fill_1 FILLER_8_1422 ();
 sg13g2_decap_4 FILLER_8_1480 ();
 sg13g2_fill_1 FILLER_8_1484 ();
 sg13g2_fill_1 FILLER_8_1499 ();
 sg13g2_fill_2 FILLER_8_1577 ();
 sg13g2_fill_1 FILLER_8_1608 ();
 sg13g2_fill_1 FILLER_8_1643 ();
 sg13g2_fill_1 FILLER_8_1653 ();
 sg13g2_fill_1 FILLER_8_1658 ();
 sg13g2_fill_2 FILLER_8_1685 ();
 sg13g2_decap_8 FILLER_8_1719 ();
 sg13g2_fill_2 FILLER_8_1757 ();
 sg13g2_decap_8 FILLER_8_1859 ();
 sg13g2_fill_1 FILLER_8_1866 ();
 sg13g2_fill_1 FILLER_8_1871 ();
 sg13g2_fill_1 FILLER_8_1882 ();
 sg13g2_fill_1 FILLER_8_1904 ();
 sg13g2_fill_1 FILLER_8_1909 ();
 sg13g2_fill_1 FILLER_8_1915 ();
 sg13g2_fill_2 FILLER_8_1926 ();
 sg13g2_fill_2 FILLER_8_1938 ();
 sg13g2_fill_1 FILLER_8_1940 ();
 sg13g2_fill_2 FILLER_8_1945 ();
 sg13g2_fill_1 FILLER_8_1947 ();
 sg13g2_fill_2 FILLER_8_1969 ();
 sg13g2_fill_1 FILLER_8_1971 ();
 sg13g2_fill_1 FILLER_8_2012 ();
 sg13g2_fill_1 FILLER_8_2023 ();
 sg13g2_decap_4 FILLER_8_2063 ();
 sg13g2_fill_2 FILLER_8_2073 ();
 sg13g2_fill_1 FILLER_8_2101 ();
 sg13g2_fill_1 FILLER_8_2106 ();
 sg13g2_fill_1 FILLER_8_2117 ();
 sg13g2_fill_2 FILLER_8_2180 ();
 sg13g2_decap_8 FILLER_8_2222 ();
 sg13g2_decap_8 FILLER_8_2229 ();
 sg13g2_decap_4 FILLER_8_2240 ();
 sg13g2_fill_2 FILLER_8_2244 ();
 sg13g2_fill_1 FILLER_8_2260 ();
 sg13g2_decap_8 FILLER_8_2291 ();
 sg13g2_decap_8 FILLER_8_2298 ();
 sg13g2_decap_8 FILLER_8_2305 ();
 sg13g2_decap_8 FILLER_8_2312 ();
 sg13g2_decap_8 FILLER_8_2319 ();
 sg13g2_decap_8 FILLER_8_2326 ();
 sg13g2_decap_8 FILLER_8_2333 ();
 sg13g2_decap_8 FILLER_8_2340 ();
 sg13g2_decap_8 FILLER_8_2347 ();
 sg13g2_decap_8 FILLER_8_2354 ();
 sg13g2_decap_4 FILLER_8_2361 ();
 sg13g2_decap_8 FILLER_8_2391 ();
 sg13g2_fill_2 FILLER_8_2398 ();
 sg13g2_fill_2 FILLER_8_2472 ();
 sg13g2_fill_1 FILLER_8_2500 ();
 sg13g2_fill_1 FILLER_8_2505 ();
 sg13g2_fill_1 FILLER_8_2558 ();
 sg13g2_decap_8 FILLER_8_2611 ();
 sg13g2_decap_8 FILLER_8_2618 ();
 sg13g2_decap_8 FILLER_8_2625 ();
 sg13g2_decap_8 FILLER_8_2632 ();
 sg13g2_decap_8 FILLER_8_2639 ();
 sg13g2_decap_8 FILLER_8_2646 ();
 sg13g2_decap_8 FILLER_8_2653 ();
 sg13g2_decap_8 FILLER_8_2660 ();
 sg13g2_fill_2 FILLER_8_2667 ();
 sg13g2_fill_1 FILLER_8_2669 ();
 sg13g2_fill_1 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_51 ();
 sg13g2_decap_4 FILLER_9_58 ();
 sg13g2_fill_2 FILLER_9_82 ();
 sg13g2_fill_1 FILLER_9_97 ();
 sg13g2_fill_2 FILLER_9_119 ();
 sg13g2_fill_2 FILLER_9_155 ();
 sg13g2_decap_4 FILLER_9_245 ();
 sg13g2_fill_1 FILLER_9_254 ();
 sg13g2_decap_4 FILLER_9_259 ();
 sg13g2_fill_1 FILLER_9_263 ();
 sg13g2_fill_2 FILLER_9_303 ();
 sg13g2_fill_2 FILLER_9_309 ();
 sg13g2_fill_1 FILLER_9_311 ();
 sg13g2_fill_1 FILLER_9_343 ();
 sg13g2_fill_1 FILLER_9_348 ();
 sg13g2_fill_2 FILLER_9_379 ();
 sg13g2_fill_2 FILLER_9_394 ();
 sg13g2_fill_1 FILLER_9_396 ();
 sg13g2_fill_1 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_471 ();
 sg13g2_fill_2 FILLER_9_483 ();
 sg13g2_fill_1 FILLER_9_485 ();
 sg13g2_fill_2 FILLER_9_495 ();
 sg13g2_fill_1 FILLER_9_506 ();
 sg13g2_fill_2 FILLER_9_579 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_4 FILLER_9_602 ();
 sg13g2_fill_2 FILLER_9_606 ();
 sg13g2_decap_8 FILLER_9_639 ();
 sg13g2_fill_2 FILLER_9_646 ();
 sg13g2_decap_8 FILLER_9_652 ();
 sg13g2_fill_2 FILLER_9_659 ();
 sg13g2_fill_1 FILLER_9_661 ();
 sg13g2_fill_2 FILLER_9_672 ();
 sg13g2_fill_1 FILLER_9_674 ();
 sg13g2_fill_1 FILLER_9_679 ();
 sg13g2_fill_1 FILLER_9_705 ();
 sg13g2_decap_4 FILLER_9_729 ();
 sg13g2_decap_8 FILLER_9_764 ();
 sg13g2_decap_4 FILLER_9_771 ();
 sg13g2_decap_8 FILLER_9_815 ();
 sg13g2_fill_2 FILLER_9_832 ();
 sg13g2_decap_4 FILLER_9_838 ();
 sg13g2_decap_8 FILLER_9_856 ();
 sg13g2_fill_2 FILLER_9_863 ();
 sg13g2_fill_1 FILLER_9_865 ();
 sg13g2_fill_1 FILLER_9_897 ();
 sg13g2_fill_1 FILLER_9_924 ();
 sg13g2_fill_1 FILLER_9_935 ();
 sg13g2_decap_4 FILLER_9_967 ();
 sg13g2_decap_8 FILLER_9_1007 ();
 sg13g2_fill_1 FILLER_9_1053 ();
 sg13g2_decap_4 FILLER_9_1058 ();
 sg13g2_fill_1 FILLER_9_1062 ();
 sg13g2_fill_2 FILLER_9_1067 ();
 sg13g2_decap_8 FILLER_9_1073 ();
 sg13g2_fill_1 FILLER_9_1080 ();
 sg13g2_fill_1 FILLER_9_1115 ();
 sg13g2_fill_1 FILLER_9_1121 ();
 sg13g2_fill_1 FILLER_9_1126 ();
 sg13g2_decap_8 FILLER_9_1157 ();
 sg13g2_decap_4 FILLER_9_1164 ();
 sg13g2_fill_2 FILLER_9_1168 ();
 sg13g2_fill_2 FILLER_9_1222 ();
 sg13g2_decap_4 FILLER_9_1232 ();
 sg13g2_decap_8 FILLER_9_1274 ();
 sg13g2_decap_8 FILLER_9_1281 ();
 sg13g2_fill_2 FILLER_9_1288 ();
 sg13g2_fill_1 FILLER_9_1290 ();
 sg13g2_fill_2 FILLER_9_1295 ();
 sg13g2_fill_1 FILLER_9_1297 ();
 sg13g2_fill_2 FILLER_9_1308 ();
 sg13g2_fill_1 FILLER_9_1310 ();
 sg13g2_decap_8 FILLER_9_1315 ();
 sg13g2_decap_8 FILLER_9_1322 ();
 sg13g2_fill_1 FILLER_9_1329 ();
 sg13g2_decap_8 FILLER_9_1334 ();
 sg13g2_decap_8 FILLER_9_1341 ();
 sg13g2_decap_4 FILLER_9_1357 ();
 sg13g2_fill_2 FILLER_9_1361 ();
 sg13g2_decap_4 FILLER_9_1368 ();
 sg13g2_fill_1 FILLER_9_1385 ();
 sg13g2_fill_1 FILLER_9_1390 ();
 sg13g2_fill_2 FILLER_9_1396 ();
 sg13g2_fill_2 FILLER_9_1408 ();
 sg13g2_fill_2 FILLER_9_1431 ();
 sg13g2_fill_2 FILLER_9_1461 ();
 sg13g2_fill_1 FILLER_9_1484 ();
 sg13g2_fill_2 FILLER_9_1518 ();
 sg13g2_fill_1 FILLER_9_1524 ();
 sg13g2_fill_1 FILLER_9_1556 ();
 sg13g2_fill_1 FILLER_9_1598 ();
 sg13g2_fill_2 FILLER_9_1616 ();
 sg13g2_fill_2 FILLER_9_1626 ();
 sg13g2_decap_4 FILLER_9_1643 ();
 sg13g2_fill_2 FILLER_9_1647 ();
 sg13g2_decap_4 FILLER_9_1654 ();
 sg13g2_fill_2 FILLER_9_1658 ();
 sg13g2_fill_2 FILLER_9_1671 ();
 sg13g2_fill_2 FILLER_9_1699 ();
 sg13g2_decap_8 FILLER_9_1705 ();
 sg13g2_decap_8 FILLER_9_1712 ();
 sg13g2_decap_4 FILLER_9_1719 ();
 sg13g2_fill_1 FILLER_9_1723 ();
 sg13g2_fill_2 FILLER_9_1733 ();
 sg13g2_fill_1 FILLER_9_1735 ();
 sg13g2_fill_2 FILLER_9_1751 ();
 sg13g2_fill_2 FILLER_9_1756 ();
 sg13g2_fill_1 FILLER_9_1767 ();
 sg13g2_fill_2 FILLER_9_1778 ();
 sg13g2_fill_2 FILLER_9_1802 ();
 sg13g2_fill_1 FILLER_9_1804 ();
 sg13g2_decap_8 FILLER_9_1859 ();
 sg13g2_decap_4 FILLER_9_1866 ();
 sg13g2_fill_2 FILLER_9_1870 ();
 sg13g2_decap_8 FILLER_9_1876 ();
 sg13g2_fill_2 FILLER_9_1887 ();
 sg13g2_decap_8 FILLER_9_1925 ();
 sg13g2_decap_8 FILLER_9_1942 ();
 sg13g2_fill_2 FILLER_9_1949 ();
 sg13g2_fill_1 FILLER_9_1964 ();
 sg13g2_decap_4 FILLER_9_2031 ();
 sg13g2_fill_2 FILLER_9_2043 ();
 sg13g2_fill_1 FILLER_9_2045 ();
 sg13g2_fill_1 FILLER_9_2050 ();
 sg13g2_fill_2 FILLER_9_2055 ();
 sg13g2_decap_4 FILLER_9_2140 ();
 sg13g2_fill_2 FILLER_9_2152 ();
 sg13g2_fill_1 FILLER_9_2154 ();
 sg13g2_fill_1 FILLER_9_2165 ();
 sg13g2_decap_8 FILLER_9_2204 ();
 sg13g2_decap_8 FILLER_9_2211 ();
 sg13g2_fill_1 FILLER_9_2218 ();
 sg13g2_fill_2 FILLER_9_2255 ();
 sg13g2_decap_8 FILLER_9_2267 ();
 sg13g2_decap_8 FILLER_9_2274 ();
 sg13g2_decap_8 FILLER_9_2281 ();
 sg13g2_decap_8 FILLER_9_2288 ();
 sg13g2_decap_8 FILLER_9_2295 ();
 sg13g2_decap_8 FILLER_9_2302 ();
 sg13g2_decap_8 FILLER_9_2309 ();
 sg13g2_decap_8 FILLER_9_2316 ();
 sg13g2_decap_8 FILLER_9_2323 ();
 sg13g2_decap_8 FILLER_9_2330 ();
 sg13g2_decap_8 FILLER_9_2337 ();
 sg13g2_decap_8 FILLER_9_2344 ();
 sg13g2_decap_8 FILLER_9_2351 ();
 sg13g2_decap_8 FILLER_9_2358 ();
 sg13g2_decap_8 FILLER_9_2365 ();
 sg13g2_fill_1 FILLER_9_2372 ();
 sg13g2_decap_8 FILLER_9_2381 ();
 sg13g2_fill_1 FILLER_9_2414 ();
 sg13g2_fill_2 FILLER_9_2444 ();
 sg13g2_decap_4 FILLER_9_2450 ();
 sg13g2_fill_1 FILLER_9_2500 ();
 sg13g2_fill_2 FILLER_9_2531 ();
 sg13g2_fill_2 FILLER_9_2573 ();
 sg13g2_decap_4 FILLER_9_2579 ();
 sg13g2_decap_8 FILLER_9_2593 ();
 sg13g2_decap_8 FILLER_9_2610 ();
 sg13g2_decap_8 FILLER_9_2617 ();
 sg13g2_decap_8 FILLER_9_2624 ();
 sg13g2_decap_8 FILLER_9_2631 ();
 sg13g2_decap_8 FILLER_9_2638 ();
 sg13g2_decap_8 FILLER_9_2645 ();
 sg13g2_decap_8 FILLER_9_2652 ();
 sg13g2_decap_8 FILLER_9_2659 ();
 sg13g2_decap_4 FILLER_9_2666 ();
 sg13g2_fill_1 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_5 ();
 sg13g2_decap_4 FILLER_10_12 ();
 sg13g2_fill_2 FILLER_10_16 ();
 sg13g2_decap_4 FILLER_10_28 ();
 sg13g2_fill_2 FILLER_10_42 ();
 sg13g2_fill_2 FILLER_10_93 ();
 sg13g2_fill_2 FILLER_10_98 ();
 sg13g2_fill_1 FILLER_10_151 ();
 sg13g2_fill_2 FILLER_10_190 ();
 sg13g2_fill_1 FILLER_10_224 ();
 sg13g2_fill_1 FILLER_10_241 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_4 FILLER_10_266 ();
 sg13g2_decap_4 FILLER_10_274 ();
 sg13g2_fill_1 FILLER_10_278 ();
 sg13g2_fill_1 FILLER_10_314 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_decap_8 FILLER_10_327 ();
 sg13g2_fill_2 FILLER_10_334 ();
 sg13g2_decap_4 FILLER_10_341 ();
 sg13g2_fill_2 FILLER_10_357 ();
 sg13g2_fill_1 FILLER_10_377 ();
 sg13g2_fill_1 FILLER_10_383 ();
 sg13g2_fill_2 FILLER_10_398 ();
 sg13g2_fill_1 FILLER_10_400 ();
 sg13g2_fill_1 FILLER_10_426 ();
 sg13g2_fill_1 FILLER_10_434 ();
 sg13g2_fill_2 FILLER_10_448 ();
 sg13g2_fill_1 FILLER_10_460 ();
 sg13g2_fill_1 FILLER_10_466 ();
 sg13g2_decap_4 FILLER_10_475 ();
 sg13g2_fill_1 FILLER_10_479 ();
 sg13g2_fill_2 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_530 ();
 sg13g2_decap_4 FILLER_10_583 ();
 sg13g2_fill_1 FILLER_10_587 ();
 sg13g2_decap_8 FILLER_10_631 ();
 sg13g2_decap_4 FILLER_10_638 ();
 sg13g2_decap_4 FILLER_10_694 ();
 sg13g2_fill_1 FILLER_10_698 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_fill_2 FILLER_10_840 ();
 sg13g2_decap_4 FILLER_10_850 ();
 sg13g2_fill_2 FILLER_10_858 ();
 sg13g2_fill_1 FILLER_10_860 ();
 sg13g2_decap_8 FILLER_10_882 ();
 sg13g2_decap_8 FILLER_10_889 ();
 sg13g2_fill_2 FILLER_10_896 ();
 sg13g2_fill_2 FILLER_10_914 ();
 sg13g2_fill_1 FILLER_10_946 ();
 sg13g2_fill_1 FILLER_10_973 ();
 sg13g2_fill_1 FILLER_10_978 ();
 sg13g2_decap_4 FILLER_10_1008 ();
 sg13g2_fill_2 FILLER_10_1016 ();
 sg13g2_fill_1 FILLER_10_1018 ();
 sg13g2_fill_2 FILLER_10_1027 ();
 sg13g2_fill_1 FILLER_10_1029 ();
 sg13g2_decap_4 FILLER_10_1034 ();
 sg13g2_fill_2 FILLER_10_1048 ();
 sg13g2_fill_1 FILLER_10_1050 ();
 sg13g2_fill_2 FILLER_10_1060 ();
 sg13g2_fill_1 FILLER_10_1062 ();
 sg13g2_fill_2 FILLER_10_1084 ();
 sg13g2_fill_1 FILLER_10_1086 ();
 sg13g2_fill_1 FILLER_10_1126 ();
 sg13g2_fill_1 FILLER_10_1132 ();
 sg13g2_fill_2 FILLER_10_1137 ();
 sg13g2_fill_1 FILLER_10_1160 ();
 sg13g2_fill_1 FILLER_10_1187 ();
 sg13g2_fill_1 FILLER_10_1193 ();
 sg13g2_fill_2 FILLER_10_1228 ();
 sg13g2_fill_1 FILLER_10_1230 ();
 sg13g2_decap_4 FILLER_10_1235 ();
 sg13g2_fill_2 FILLER_10_1239 ();
 sg13g2_decap_8 FILLER_10_1262 ();
 sg13g2_fill_2 FILLER_10_1269 ();
 sg13g2_fill_1 FILLER_10_1271 ();
 sg13g2_decap_8 FILLER_10_1343 ();
 sg13g2_decap_8 FILLER_10_1350 ();
 sg13g2_decap_8 FILLER_10_1357 ();
 sg13g2_fill_1 FILLER_10_1364 ();
 sg13g2_fill_1 FILLER_10_1373 ();
 sg13g2_fill_1 FILLER_10_1388 ();
 sg13g2_fill_1 FILLER_10_1394 ();
 sg13g2_fill_1 FILLER_10_1400 ();
 sg13g2_fill_1 FILLER_10_1411 ();
 sg13g2_fill_2 FILLER_10_1417 ();
 sg13g2_decap_4 FILLER_10_1429 ();
 sg13g2_fill_1 FILLER_10_1433 ();
 sg13g2_decap_4 FILLER_10_1437 ();
 sg13g2_fill_1 FILLER_10_1441 ();
 sg13g2_fill_2 FILLER_10_1470 ();
 sg13g2_fill_1 FILLER_10_1472 ();
 sg13g2_fill_2 FILLER_10_1509 ();
 sg13g2_fill_1 FILLER_10_1537 ();
 sg13g2_fill_2 FILLER_10_1566 ();
 sg13g2_fill_2 FILLER_10_1572 ();
 sg13g2_fill_2 FILLER_10_1582 ();
 sg13g2_fill_1 FILLER_10_1612 ();
 sg13g2_fill_2 FILLER_10_1630 ();
 sg13g2_decap_8 FILLER_10_1643 ();
 sg13g2_decap_8 FILLER_10_1650 ();
 sg13g2_decap_8 FILLER_10_1657 ();
 sg13g2_decap_4 FILLER_10_1664 ();
 sg13g2_fill_2 FILLER_10_1668 ();
 sg13g2_decap_4 FILLER_10_1674 ();
 sg13g2_fill_2 FILLER_10_1678 ();
 sg13g2_decap_8 FILLER_10_1705 ();
 sg13g2_decap_4 FILLER_10_1712 ();
 sg13g2_fill_2 FILLER_10_1716 ();
 sg13g2_decap_8 FILLER_10_1792 ();
 sg13g2_fill_1 FILLER_10_1799 ();
 sg13g2_fill_2 FILLER_10_1836 ();
 sg13g2_decap_8 FILLER_10_1842 ();
 sg13g2_decap_8 FILLER_10_1849 ();
 sg13g2_decap_8 FILLER_10_1856 ();
 sg13g2_fill_2 FILLER_10_1889 ();
 sg13g2_fill_1 FILLER_10_1891 ();
 sg13g2_fill_1 FILLER_10_1913 ();
 sg13g2_fill_2 FILLER_10_1935 ();
 sg13g2_fill_1 FILLER_10_1963 ();
 sg13g2_fill_1 FILLER_10_1968 ();
 sg13g2_decap_8 FILLER_10_1979 ();
 sg13g2_fill_1 FILLER_10_1986 ();
 sg13g2_fill_1 FILLER_10_1999 ();
 sg13g2_decap_8 FILLER_10_2004 ();
 sg13g2_decap_8 FILLER_10_2011 ();
 sg13g2_decap_8 FILLER_10_2018 ();
 sg13g2_decap_4 FILLER_10_2025 ();
 sg13g2_fill_1 FILLER_10_2029 ();
 sg13g2_fill_1 FILLER_10_2058 ();
 sg13g2_fill_1 FILLER_10_2066 ();
 sg13g2_decap_8 FILLER_10_2105 ();
 sg13g2_fill_2 FILLER_10_2112 ();
 sg13g2_fill_1 FILLER_10_2114 ();
 sg13g2_fill_1 FILLER_10_2131 ();
 sg13g2_fill_1 FILLER_10_2144 ();
 sg13g2_fill_2 FILLER_10_2166 ();
 sg13g2_fill_2 FILLER_10_2208 ();
 sg13g2_fill_1 FILLER_10_2231 ();
 sg13g2_decap_8 FILLER_10_2278 ();
 sg13g2_decap_8 FILLER_10_2285 ();
 sg13g2_decap_8 FILLER_10_2292 ();
 sg13g2_decap_8 FILLER_10_2299 ();
 sg13g2_decap_8 FILLER_10_2306 ();
 sg13g2_fill_1 FILLER_10_2313 ();
 sg13g2_decap_8 FILLER_10_2324 ();
 sg13g2_decap_8 FILLER_10_2331 ();
 sg13g2_decap_8 FILLER_10_2338 ();
 sg13g2_decap_8 FILLER_10_2397 ();
 sg13g2_decap_4 FILLER_10_2404 ();
 sg13g2_fill_2 FILLER_10_2434 ();
 sg13g2_fill_1 FILLER_10_2436 ();
 sg13g2_decap_4 FILLER_10_2463 ();
 sg13g2_fill_1 FILLER_10_2467 ();
 sg13g2_fill_2 FILLER_10_2478 ();
 sg13g2_fill_1 FILLER_10_2484 ();
 sg13g2_fill_1 FILLER_10_2489 ();
 sg13g2_decap_8 FILLER_10_2494 ();
 sg13g2_decap_8 FILLER_10_2501 ();
 sg13g2_fill_2 FILLER_10_2522 ();
 sg13g2_fill_1 FILLER_10_2524 ();
 sg13g2_fill_1 FILLER_10_2535 ();
 sg13g2_decap_8 FILLER_10_2544 ();
 sg13g2_decap_8 FILLER_10_2551 ();
 sg13g2_decap_8 FILLER_10_2558 ();
 sg13g2_decap_4 FILLER_10_2565 ();
 sg13g2_fill_1 FILLER_10_2569 ();
 sg13g2_decap_8 FILLER_10_2580 ();
 sg13g2_decap_8 FILLER_10_2623 ();
 sg13g2_decap_8 FILLER_10_2630 ();
 sg13g2_decap_8 FILLER_10_2637 ();
 sg13g2_decap_8 FILLER_10_2644 ();
 sg13g2_decap_8 FILLER_10_2651 ();
 sg13g2_decap_8 FILLER_10_2658 ();
 sg13g2_decap_4 FILLER_10_2665 ();
 sg13g2_fill_1 FILLER_10_2669 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_58 ();
 sg13g2_decap_4 FILLER_11_86 ();
 sg13g2_fill_2 FILLER_11_116 ();
 sg13g2_fill_2 FILLER_11_148 ();
 sg13g2_fill_1 FILLER_11_159 ();
 sg13g2_fill_2 FILLER_11_175 ();
 sg13g2_fill_1 FILLER_11_185 ();
 sg13g2_fill_2 FILLER_11_209 ();
 sg13g2_fill_1 FILLER_11_211 ();
 sg13g2_fill_2 FILLER_11_216 ();
 sg13g2_fill_1 FILLER_11_249 ();
 sg13g2_fill_1 FILLER_11_285 ();
 sg13g2_fill_1 FILLER_11_328 ();
 sg13g2_decap_8 FILLER_11_337 ();
 sg13g2_decap_4 FILLER_11_344 ();
 sg13g2_fill_2 FILLER_11_348 ();
 sg13g2_fill_2 FILLER_11_386 ();
 sg13g2_fill_2 FILLER_11_393 ();
 sg13g2_fill_1 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_408 ();
 sg13g2_fill_1 FILLER_11_423 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_fill_1 FILLER_11_444 ();
 sg13g2_fill_1 FILLER_11_454 ();
 sg13g2_fill_1 FILLER_11_460 ();
 sg13g2_fill_2 FILLER_11_472 ();
 sg13g2_decap_4 FILLER_11_484 ();
 sg13g2_fill_1 FILLER_11_492 ();
 sg13g2_fill_2 FILLER_11_497 ();
 sg13g2_fill_2 FILLER_11_514 ();
 sg13g2_decap_8 FILLER_11_526 ();
 sg13g2_decap_4 FILLER_11_533 ();
 sg13g2_fill_1 FILLER_11_537 ();
 sg13g2_fill_1 FILLER_11_550 ();
 sg13g2_fill_1 FILLER_11_556 ();
 sg13g2_decap_4 FILLER_11_569 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_4 FILLER_11_651 ();
 sg13g2_fill_1 FILLER_11_655 ();
 sg13g2_decap_8 FILLER_11_660 ();
 sg13g2_fill_2 FILLER_11_667 ();
 sg13g2_fill_2 FILLER_11_699 ();
 sg13g2_fill_2 FILLER_11_705 ();
 sg13g2_fill_1 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_800 ();
 sg13g2_decap_8 FILLER_11_807 ();
 sg13g2_decap_4 FILLER_11_814 ();
 sg13g2_fill_2 FILLER_11_818 ();
 sg13g2_fill_1 FILLER_11_840 ();
 sg13g2_fill_2 FILLER_11_867 ();
 sg13g2_fill_1 FILLER_11_869 ();
 sg13g2_decap_8 FILLER_11_896 ();
 sg13g2_fill_2 FILLER_11_903 ();
 sg13g2_fill_2 FILLER_11_954 ();
 sg13g2_fill_1 FILLER_11_956 ();
 sg13g2_fill_2 FILLER_11_983 ();
 sg13g2_fill_1 FILLER_11_985 ();
 sg13g2_fill_2 FILLER_11_1027 ();
 sg13g2_fill_2 FILLER_11_1033 ();
 sg13g2_fill_1 FILLER_11_1061 ();
 sg13g2_fill_2 FILLER_11_1088 ();
 sg13g2_fill_2 FILLER_11_1095 ();
 sg13g2_fill_2 FILLER_11_1101 ();
 sg13g2_decap_8 FILLER_11_1107 ();
 sg13g2_fill_2 FILLER_11_1114 ();
 sg13g2_fill_1 FILLER_11_1116 ();
 sg13g2_decap_8 FILLER_11_1143 ();
 sg13g2_decap_4 FILLER_11_1150 ();
 sg13g2_fill_2 FILLER_11_1154 ();
 sg13g2_fill_1 FILLER_11_1177 ();
 sg13g2_fill_2 FILLER_11_1191 ();
 sg13g2_fill_1 FILLER_11_1193 ();
 sg13g2_fill_2 FILLER_11_1199 ();
 sg13g2_fill_1 FILLER_11_1201 ();
 sg13g2_fill_1 FILLER_11_1219 ();
 sg13g2_decap_8 FILLER_11_1331 ();
 sg13g2_decap_8 FILLER_11_1338 ();
 sg13g2_decap_4 FILLER_11_1345 ();
 sg13g2_fill_1 FILLER_11_1349 ();
 sg13g2_fill_2 FILLER_11_1386 ();
 sg13g2_fill_1 FILLER_11_1388 ();
 sg13g2_decap_8 FILLER_11_1394 ();
 sg13g2_decap_4 FILLER_11_1401 ();
 sg13g2_fill_1 FILLER_11_1405 ();
 sg13g2_fill_2 FILLER_11_1429 ();
 sg13g2_fill_1 FILLER_11_1436 ();
 sg13g2_fill_1 FILLER_11_1445 ();
 sg13g2_fill_1 FILLER_11_1477 ();
 sg13g2_fill_1 FILLER_11_1483 ();
 sg13g2_fill_2 FILLER_11_1489 ();
 sg13g2_fill_2 FILLER_11_1511 ();
 sg13g2_fill_1 FILLER_11_1556 ();
 sg13g2_fill_2 FILLER_11_1591 ();
 sg13g2_fill_1 FILLER_11_1601 ();
 sg13g2_fill_2 FILLER_11_1635 ();
 sg13g2_fill_1 FILLER_11_1652 ();
 sg13g2_decap_8 FILLER_11_1683 ();
 sg13g2_fill_2 FILLER_11_1690 ();
 sg13g2_fill_2 FILLER_11_1696 ();
 sg13g2_fill_1 FILLER_11_1698 ();
 sg13g2_decap_8 FILLER_11_1708 ();
 sg13g2_fill_1 FILLER_11_1715 ();
 sg13g2_fill_2 FILLER_11_1724 ();
 sg13g2_fill_1 FILLER_11_1726 ();
 sg13g2_fill_1 FILLER_11_1737 ();
 sg13g2_fill_2 FILLER_11_1754 ();
 sg13g2_fill_2 FILLER_11_1760 ();
 sg13g2_fill_1 FILLER_11_1762 ();
 sg13g2_fill_1 FILLER_11_1767 ();
 sg13g2_fill_2 FILLER_11_1772 ();
 sg13g2_fill_1 FILLER_11_1774 ();
 sg13g2_fill_2 FILLER_11_1792 ();
 sg13g2_fill_1 FILLER_11_1794 ();
 sg13g2_fill_2 FILLER_11_1811 ();
 sg13g2_decap_8 FILLER_11_1821 ();
 sg13g2_decap_8 FILLER_11_1828 ();
 sg13g2_decap_8 FILLER_11_1835 ();
 sg13g2_decap_4 FILLER_11_1842 ();
 sg13g2_fill_2 FILLER_11_1846 ();
 sg13g2_fill_2 FILLER_11_1894 ();
 sg13g2_fill_2 FILLER_11_1904 ();
 sg13g2_decap_8 FILLER_11_1910 ();
 sg13g2_decap_4 FILLER_11_1917 ();
 sg13g2_fill_2 FILLER_11_1921 ();
 sg13g2_decap_4 FILLER_11_1959 ();
 sg13g2_decap_8 FILLER_11_1967 ();
 sg13g2_fill_2 FILLER_11_1974 ();
 sg13g2_decap_8 FILLER_11_2006 ();
 sg13g2_fill_1 FILLER_11_2013 ();
 sg13g2_decap_8 FILLER_11_2018 ();
 sg13g2_fill_2 FILLER_11_2035 ();
 sg13g2_fill_1 FILLER_11_2037 ();
 sg13g2_decap_4 FILLER_11_2096 ();
 sg13g2_fill_2 FILLER_11_2116 ();
 sg13g2_fill_2 FILLER_11_2144 ();
 sg13g2_decap_8 FILLER_11_2182 ();
 sg13g2_decap_4 FILLER_11_2189 ();
 sg13g2_fill_2 FILLER_11_2193 ();
 sg13g2_decap_8 FILLER_11_2280 ();
 sg13g2_decap_8 FILLER_11_2287 ();
 sg13g2_decap_4 FILLER_11_2294 ();
 sg13g2_fill_2 FILLER_11_2324 ();
 sg13g2_fill_2 FILLER_11_2330 ();
 sg13g2_fill_2 FILLER_11_2342 ();
 sg13g2_decap_4 FILLER_11_2348 ();
 sg13g2_fill_2 FILLER_11_2356 ();
 sg13g2_fill_2 FILLER_11_2368 ();
 sg13g2_fill_2 FILLER_11_2380 ();
 sg13g2_fill_1 FILLER_11_2382 ();
 sg13g2_fill_1 FILLER_11_2393 ();
 sg13g2_fill_2 FILLER_11_2420 ();
 sg13g2_fill_1 FILLER_11_2422 ();
 sg13g2_decap_8 FILLER_11_2469 ();
 sg13g2_decap_8 FILLER_11_2476 ();
 sg13g2_fill_2 FILLER_11_2483 ();
 sg13g2_fill_1 FILLER_11_2485 ();
 sg13g2_decap_8 FILLER_11_2512 ();
 sg13g2_decap_8 FILLER_11_2519 ();
 sg13g2_fill_2 FILLER_11_2526 ();
 sg13g2_fill_1 FILLER_11_2528 ();
 sg13g2_fill_2 FILLER_11_2555 ();
 sg13g2_decap_4 FILLER_11_2567 ();
 sg13g2_fill_2 FILLER_11_2571 ();
 sg13g2_decap_8 FILLER_11_2617 ();
 sg13g2_fill_1 FILLER_11_2624 ();
 sg13g2_decap_8 FILLER_11_2629 ();
 sg13g2_decap_8 FILLER_11_2636 ();
 sg13g2_decap_8 FILLER_11_2643 ();
 sg13g2_decap_8 FILLER_11_2650 ();
 sg13g2_decap_8 FILLER_11_2657 ();
 sg13g2_decap_4 FILLER_11_2664 ();
 sg13g2_fill_2 FILLER_11_2668 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_12 ();
 sg13g2_fill_2 FILLER_12_129 ();
 sg13g2_fill_2 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_147 ();
 sg13g2_fill_2 FILLER_12_155 ();
 sg13g2_fill_2 FILLER_12_177 ();
 sg13g2_fill_1 FILLER_12_188 ();
 sg13g2_fill_1 FILLER_12_231 ();
 sg13g2_fill_2 FILLER_12_279 ();
 sg13g2_fill_2 FILLER_12_285 ();
 sg13g2_fill_1 FILLER_12_325 ();
 sg13g2_decap_4 FILLER_12_331 ();
 sg13g2_fill_1 FILLER_12_335 ();
 sg13g2_fill_1 FILLER_12_350 ();
 sg13g2_fill_2 FILLER_12_374 ();
 sg13g2_decap_4 FILLER_12_381 ();
 sg13g2_fill_2 FILLER_12_385 ();
 sg13g2_fill_1 FILLER_12_391 ();
 sg13g2_fill_2 FILLER_12_397 ();
 sg13g2_fill_1 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_fill_1 FILLER_12_444 ();
 sg13g2_fill_1 FILLER_12_450 ();
 sg13g2_decap_4 FILLER_12_507 ();
 sg13g2_fill_2 FILLER_12_511 ();
 sg13g2_decap_4 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_540 ();
 sg13g2_fill_2 FILLER_12_573 ();
 sg13g2_fill_1 FILLER_12_575 ();
 sg13g2_fill_1 FILLER_12_585 ();
 sg13g2_fill_2 FILLER_12_609 ();
 sg13g2_fill_2 FILLER_12_621 ();
 sg13g2_fill_2 FILLER_12_646 ();
 sg13g2_decap_8 FILLER_12_684 ();
 sg13g2_decap_4 FILLER_12_731 ();
 sg13g2_fill_2 FILLER_12_745 ();
 sg13g2_fill_1 FILLER_12_747 ();
 sg13g2_fill_2 FILLER_12_752 ();
 sg13g2_decap_8 FILLER_12_758 ();
 sg13g2_decap_4 FILLER_12_770 ();
 sg13g2_fill_1 FILLER_12_774 ();
 sg13g2_decap_8 FILLER_12_815 ();
 sg13g2_fill_1 FILLER_12_822 ();
 sg13g2_fill_2 FILLER_12_875 ();
 sg13g2_decap_4 FILLER_12_881 ();
 sg13g2_fill_2 FILLER_12_885 ();
 sg13g2_decap_8 FILLER_12_913 ();
 sg13g2_decap_4 FILLER_12_920 ();
 sg13g2_decap_8 FILLER_12_949 ();
 sg13g2_decap_4 FILLER_12_956 ();
 sg13g2_fill_1 FILLER_12_960 ();
 sg13g2_decap_8 FILLER_12_971 ();
 sg13g2_decap_8 FILLER_12_1025 ();
 sg13g2_decap_4 FILLER_12_1032 ();
 sg13g2_fill_1 FILLER_12_1036 ();
 sg13g2_decap_8 FILLER_12_1077 ();
 sg13g2_decap_8 FILLER_12_1084 ();
 sg13g2_decap_4 FILLER_12_1091 ();
 sg13g2_fill_1 FILLER_12_1095 ();
 sg13g2_fill_1 FILLER_12_1113 ();
 sg13g2_fill_1 FILLER_12_1127 ();
 sg13g2_decap_8 FILLER_12_1140 ();
 sg13g2_fill_2 FILLER_12_1147 ();
 sg13g2_fill_1 FILLER_12_1149 ();
 sg13g2_fill_1 FILLER_12_1163 ();
 sg13g2_fill_2 FILLER_12_1202 ();
 sg13g2_fill_2 FILLER_12_1234 ();
 sg13g2_fill_1 FILLER_12_1339 ();
 sg13g2_fill_1 FILLER_12_1344 ();
 sg13g2_fill_2 FILLER_12_1349 ();
 sg13g2_fill_2 FILLER_12_1356 ();
 sg13g2_fill_2 FILLER_12_1368 ();
 sg13g2_fill_1 FILLER_12_1370 ();
 sg13g2_fill_2 FILLER_12_1381 ();
 sg13g2_fill_1 FILLER_12_1433 ();
 sg13g2_decap_4 FILLER_12_1439 ();
 sg13g2_fill_2 FILLER_12_1447 ();
 sg13g2_decap_4 FILLER_12_1459 ();
 sg13g2_fill_1 FILLER_12_1463 ();
 sg13g2_fill_1 FILLER_12_1480 ();
 sg13g2_fill_1 FILLER_12_1486 ();
 sg13g2_fill_1 FILLER_12_1491 ();
 sg13g2_fill_1 FILLER_12_1496 ();
 sg13g2_fill_1 FILLER_12_1506 ();
 sg13g2_fill_1 FILLER_12_1533 ();
 sg13g2_fill_1 FILLER_12_1560 ();
 sg13g2_fill_1 FILLER_12_1571 ();
 sg13g2_fill_1 FILLER_12_1598 ();
 sg13g2_fill_2 FILLER_12_1608 ();
 sg13g2_fill_1 FILLER_12_1645 ();
 sg13g2_fill_1 FILLER_12_1677 ();
 sg13g2_decap_8 FILLER_12_1715 ();
 sg13g2_fill_2 FILLER_12_1735 ();
 sg13g2_fill_2 FILLER_12_1749 ();
 sg13g2_fill_2 FILLER_12_1755 ();
 sg13g2_fill_2 FILLER_12_1762 ();
 sg13g2_fill_1 FILLER_12_1768 ();
 sg13g2_fill_1 FILLER_12_1803 ();
 sg13g2_fill_2 FILLER_12_1809 ();
 sg13g2_decap_8 FILLER_12_1847 ();
 sg13g2_decap_4 FILLER_12_1854 ();
 sg13g2_fill_2 FILLER_12_1858 ();
 sg13g2_decap_8 FILLER_12_1874 ();
 sg13g2_fill_2 FILLER_12_1881 ();
 sg13g2_fill_1 FILLER_12_1919 ();
 sg13g2_decap_8 FILLER_12_1965 ();
 sg13g2_decap_8 FILLER_12_1998 ();
 sg13g2_fill_2 FILLER_12_2005 ();
 sg13g2_fill_1 FILLER_12_2015 ();
 sg13g2_fill_1 FILLER_12_2052 ();
 sg13g2_fill_2 FILLER_12_2085 ();
 sg13g2_fill_1 FILLER_12_2156 ();
 sg13g2_fill_1 FILLER_12_2170 ();
 sg13g2_decap_4 FILLER_12_2194 ();
 sg13g2_fill_2 FILLER_12_2198 ();
 sg13g2_fill_2 FILLER_12_2230 ();
 sg13g2_fill_1 FILLER_12_2232 ();
 sg13g2_fill_1 FILLER_12_2311 ();
 sg13g2_decap_8 FILLER_12_2352 ();
 sg13g2_decap_8 FILLER_12_2359 ();
 sg13g2_fill_1 FILLER_12_2418 ();
 sg13g2_decap_8 FILLER_12_2423 ();
 sg13g2_fill_2 FILLER_12_2430 ();
 sg13g2_fill_1 FILLER_12_2432 ();
 sg13g2_fill_2 FILLER_12_2469 ();
 sg13g2_fill_1 FILLER_12_2471 ();
 sg13g2_fill_1 FILLER_12_2484 ();
 sg13g2_fill_2 FILLER_12_2490 ();
 sg13g2_fill_1 FILLER_12_2492 ();
 sg13g2_decap_4 FILLER_12_2516 ();
 sg13g2_fill_1 FILLER_12_2520 ();
 sg13g2_decap_8 FILLER_12_2635 ();
 sg13g2_decap_8 FILLER_12_2642 ();
 sg13g2_decap_8 FILLER_12_2649 ();
 sg13g2_decap_8 FILLER_12_2656 ();
 sg13g2_decap_8 FILLER_12_2663 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_4 FILLER_13_14 ();
 sg13g2_fill_2 FILLER_13_18 ();
 sg13g2_decap_8 FILLER_13_81 ();
 sg13g2_decap_8 FILLER_13_88 ();
 sg13g2_fill_1 FILLER_13_132 ();
 sg13g2_fill_1 FILLER_13_164 ();
 sg13g2_fill_2 FILLER_13_194 ();
 sg13g2_fill_2 FILLER_13_205 ();
 sg13g2_fill_1 FILLER_13_211 ();
 sg13g2_fill_1 FILLER_13_216 ();
 sg13g2_fill_2 FILLER_13_236 ();
 sg13g2_fill_1 FILLER_13_264 ();
 sg13g2_fill_1 FILLER_13_268 ();
 sg13g2_fill_2 FILLER_13_283 ();
 sg13g2_fill_1 FILLER_13_290 ();
 sg13g2_fill_2 FILLER_13_296 ();
 sg13g2_fill_1 FILLER_13_308 ();
 sg13g2_fill_1 FILLER_13_315 ();
 sg13g2_fill_1 FILLER_13_326 ();
 sg13g2_decap_4 FILLER_13_332 ();
 sg13g2_fill_2 FILLER_13_336 ();
 sg13g2_fill_1 FILLER_13_366 ();
 sg13g2_fill_2 FILLER_13_370 ();
 sg13g2_fill_1 FILLER_13_381 ();
 sg13g2_fill_1 FILLER_13_387 ();
 sg13g2_fill_1 FILLER_13_440 ();
 sg13g2_fill_2 FILLER_13_445 ();
 sg13g2_decap_8 FILLER_13_452 ();
 sg13g2_fill_1 FILLER_13_459 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_fill_2 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_537 ();
 sg13g2_decap_8 FILLER_13_544 ();
 sg13g2_fill_2 FILLER_13_551 ();
 sg13g2_fill_1 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_558 ();
 sg13g2_decap_4 FILLER_13_565 ();
 sg13g2_fill_1 FILLER_13_569 ();
 sg13g2_fill_2 FILLER_13_619 ();
 sg13g2_fill_1 FILLER_13_621 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_682 ();
 sg13g2_decap_4 FILLER_13_699 ();
 sg13g2_fill_2 FILLER_13_707 ();
 sg13g2_fill_2 FILLER_13_722 ();
 sg13g2_decap_8 FILLER_13_732 ();
 sg13g2_decap_8 FILLER_13_739 ();
 sg13g2_decap_8 FILLER_13_746 ();
 sg13g2_fill_2 FILLER_13_753 ();
 sg13g2_decap_4 FILLER_13_759 ();
 sg13g2_fill_2 FILLER_13_763 ();
 sg13g2_decap_4 FILLER_13_774 ();
 sg13g2_fill_1 FILLER_13_778 ();
 sg13g2_decap_8 FILLER_13_810 ();
 sg13g2_fill_2 FILLER_13_817 ();
 sg13g2_fill_1 FILLER_13_819 ();
 sg13g2_fill_1 FILLER_13_828 ();
 sg13g2_fill_1 FILLER_13_843 ();
 sg13g2_fill_1 FILLER_13_854 ();
 sg13g2_fill_2 FILLER_13_859 ();
 sg13g2_fill_1 FILLER_13_866 ();
 sg13g2_decap_8 FILLER_13_877 ();
 sg13g2_fill_1 FILLER_13_884 ();
 sg13g2_decap_8 FILLER_13_941 ();
 sg13g2_fill_2 FILLER_13_948 ();
 sg13g2_fill_1 FILLER_13_950 ();
 sg13g2_fill_1 FILLER_13_977 ();
 sg13g2_fill_2 FILLER_13_1018 ();
 sg13g2_decap_8 FILLER_13_1025 ();
 sg13g2_decap_4 FILLER_13_1032 ();
 sg13g2_fill_2 FILLER_13_1062 ();
 sg13g2_fill_1 FILLER_13_1064 ();
 sg13g2_fill_2 FILLER_13_1082 ();
 sg13g2_fill_1 FILLER_13_1084 ();
 sg13g2_fill_2 FILLER_13_1115 ();
 sg13g2_fill_1 FILLER_13_1117 ();
 sg13g2_fill_1 FILLER_13_1122 ();
 sg13g2_fill_2 FILLER_13_1149 ();
 sg13g2_fill_1 FILLER_13_1151 ();
 sg13g2_fill_2 FILLER_13_1222 ();
 sg13g2_decap_8 FILLER_13_1253 ();
 sg13g2_fill_2 FILLER_13_1260 ();
 sg13g2_fill_2 FILLER_13_1288 ();
 sg13g2_decap_4 FILLER_13_1294 ();
 sg13g2_fill_1 FILLER_13_1298 ();
 sg13g2_fill_1 FILLER_13_1309 ();
 sg13g2_fill_1 FILLER_13_1331 ();
 sg13g2_fill_1 FILLER_13_1384 ();
 sg13g2_decap_4 FILLER_13_1406 ();
 sg13g2_fill_2 FILLER_13_1418 ();
 sg13g2_fill_1 FILLER_13_1425 ();
 sg13g2_fill_1 FILLER_13_1431 ();
 sg13g2_fill_1 FILLER_13_1436 ();
 sg13g2_fill_1 FILLER_13_1441 ();
 sg13g2_fill_2 FILLER_13_1446 ();
 sg13g2_fill_2 FILLER_13_1453 ();
 sg13g2_fill_2 FILLER_13_1460 ();
 sg13g2_fill_1 FILLER_13_1462 ();
 sg13g2_fill_1 FILLER_13_1480 ();
 sg13g2_fill_2 FILLER_13_1513 ();
 sg13g2_fill_1 FILLER_13_1525 ();
 sg13g2_fill_1 FILLER_13_1531 ();
 sg13g2_fill_1 FILLER_13_1541 ();
 sg13g2_fill_1 FILLER_13_1553 ();
 sg13g2_fill_2 FILLER_13_1558 ();
 sg13g2_fill_1 FILLER_13_1564 ();
 sg13g2_fill_1 FILLER_13_1570 ();
 sg13g2_fill_1 FILLER_13_1575 ();
 sg13g2_fill_1 FILLER_13_1580 ();
 sg13g2_fill_1 FILLER_13_1585 ();
 sg13g2_decap_4 FILLER_13_1720 ();
 sg13g2_fill_1 FILLER_13_1724 ();
 sg13g2_fill_1 FILLER_13_1752 ();
 sg13g2_decap_8 FILLER_13_1758 ();
 sg13g2_fill_1 FILLER_13_1765 ();
 sg13g2_decap_4 FILLER_13_1776 ();
 sg13g2_fill_1 FILLER_13_1780 ();
 sg13g2_decap_4 FILLER_13_1807 ();
 sg13g2_fill_2 FILLER_13_1811 ();
 sg13g2_fill_1 FILLER_13_1818 ();
 sg13g2_fill_2 FILLER_13_1845 ();
 sg13g2_decap_8 FILLER_13_1904 ();
 sg13g2_decap_8 FILLER_13_1911 ();
 sg13g2_fill_2 FILLER_13_1943 ();
 sg13g2_fill_2 FILLER_13_1949 ();
 sg13g2_fill_1 FILLER_13_1951 ();
 sg13g2_fill_2 FILLER_13_1962 ();
 sg13g2_fill_1 FILLER_13_1964 ();
 sg13g2_decap_4 FILLER_13_1975 ();
 sg13g2_fill_2 FILLER_13_1979 ();
 sg13g2_decap_8 FILLER_13_1985 ();
 sg13g2_decap_8 FILLER_13_1992 ();
 sg13g2_fill_1 FILLER_13_2016 ();
 sg13g2_fill_1 FILLER_13_2021 ();
 sg13g2_fill_1 FILLER_13_2069 ();
 sg13g2_fill_1 FILLER_13_2096 ();
 sg13g2_fill_2 FILLER_13_2101 ();
 sg13g2_fill_2 FILLER_13_2160 ();
 sg13g2_fill_1 FILLER_13_2162 ();
 sg13g2_decap_4 FILLER_13_2184 ();
 sg13g2_fill_2 FILLER_13_2192 ();
 sg13g2_decap_4 FILLER_13_2204 ();
 sg13g2_decap_8 FILLER_13_2218 ();
 sg13g2_decap_8 FILLER_13_2225 ();
 sg13g2_decap_8 FILLER_13_2232 ();
 sg13g2_fill_1 FILLER_13_2239 ();
 sg13g2_fill_1 FILLER_13_2273 ();
 sg13g2_decap_8 FILLER_13_2278 ();
 sg13g2_decap_8 FILLER_13_2285 ();
 sg13g2_decap_4 FILLER_13_2309 ();
 sg13g2_fill_2 FILLER_13_2313 ();
 sg13g2_fill_2 FILLER_13_2323 ();
 sg13g2_fill_1 FILLER_13_2325 ();
 sg13g2_fill_2 FILLER_13_2331 ();
 sg13g2_fill_1 FILLER_13_2359 ();
 sg13g2_fill_1 FILLER_13_2364 ();
 sg13g2_fill_1 FILLER_13_2397 ();
 sg13g2_decap_8 FILLER_13_2416 ();
 sg13g2_decap_8 FILLER_13_2429 ();
 sg13g2_decap_4 FILLER_13_2436 ();
 sg13g2_fill_1 FILLER_13_2440 ();
 sg13g2_fill_2 FILLER_13_2491 ();
 sg13g2_fill_1 FILLER_13_2493 ();
 sg13g2_fill_2 FILLER_13_2506 ();
 sg13g2_fill_1 FILLER_13_2514 ();
 sg13g2_fill_1 FILLER_13_2541 ();
 sg13g2_fill_1 FILLER_13_2569 ();
 sg13g2_fill_2 FILLER_13_2574 ();
 sg13g2_fill_1 FILLER_13_2600 ();
 sg13g2_fill_2 FILLER_13_2604 ();
 sg13g2_fill_1 FILLER_13_2630 ();
 sg13g2_decap_8 FILLER_13_2657 ();
 sg13g2_decap_4 FILLER_13_2664 ();
 sg13g2_fill_2 FILLER_13_2668 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_1 FILLER_14_18 ();
 sg13g2_decap_4 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_53 ();
 sg13g2_decap_4 FILLER_14_59 ();
 sg13g2_fill_1 FILLER_14_63 ();
 sg13g2_decap_4 FILLER_14_72 ();
 sg13g2_decap_8 FILLER_14_85 ();
 sg13g2_fill_1 FILLER_14_92 ();
 sg13g2_fill_2 FILLER_14_183 ();
 sg13g2_fill_1 FILLER_14_288 ();
 sg13g2_fill_2 FILLER_14_298 ();
 sg13g2_fill_1 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_332 ();
 sg13g2_fill_2 FILLER_14_339 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_fill_2 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_decap_8 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_decap_4 FILLER_14_388 ();
 sg13g2_fill_1 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_fill_1 FILLER_14_409 ();
 sg13g2_fill_1 FILLER_14_414 ();
 sg13g2_fill_1 FILLER_14_420 ();
 sg13g2_fill_1 FILLER_14_451 ();
 sg13g2_decap_8 FILLER_14_457 ();
 sg13g2_fill_2 FILLER_14_464 ();
 sg13g2_fill_2 FILLER_14_470 ();
 sg13g2_decap_8 FILLER_14_488 ();
 sg13g2_decap_8 FILLER_14_495 ();
 sg13g2_decap_8 FILLER_14_502 ();
 sg13g2_decap_4 FILLER_14_509 ();
 sg13g2_fill_2 FILLER_14_513 ();
 sg13g2_fill_2 FILLER_14_554 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_4 FILLER_14_581 ();
 sg13g2_fill_2 FILLER_14_585 ();
 sg13g2_fill_2 FILLER_14_609 ();
 sg13g2_fill_1 FILLER_14_611 ();
 sg13g2_fill_2 FILLER_14_623 ();
 sg13g2_fill_2 FILLER_14_639 ();
 sg13g2_fill_2 FILLER_14_645 ();
 sg13g2_fill_1 FILLER_14_647 ();
 sg13g2_fill_1 FILLER_14_674 ();
 sg13g2_fill_1 FILLER_14_701 ();
 sg13g2_fill_2 FILLER_14_726 ();
 sg13g2_fill_1 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_775 ();
 sg13g2_fill_1 FILLER_14_782 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_4 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_867 ();
 sg13g2_decap_4 FILLER_14_874 ();
 sg13g2_fill_1 FILLER_14_878 ();
 sg13g2_decap_8 FILLER_14_883 ();
 sg13g2_decap_4 FILLER_14_890 ();
 sg13g2_fill_2 FILLER_14_898 ();
 sg13g2_fill_2 FILLER_14_905 ();
 sg13g2_decap_4 FILLER_14_943 ();
 sg13g2_fill_2 FILLER_14_947 ();
 sg13g2_fill_1 FILLER_14_975 ();
 sg13g2_fill_2 FILLER_14_986 ();
 sg13g2_fill_2 FILLER_14_998 ();
 sg13g2_fill_2 FILLER_14_1004 ();
 sg13g2_fill_1 FILLER_14_1006 ();
 sg13g2_decap_8 FILLER_14_1011 ();
 sg13g2_decap_8 FILLER_14_1018 ();
 sg13g2_decap_8 FILLER_14_1025 ();
 sg13g2_decap_8 FILLER_14_1032 ();
 sg13g2_decap_4 FILLER_14_1039 ();
 sg13g2_fill_1 FILLER_14_1043 ();
 sg13g2_fill_2 FILLER_14_1048 ();
 sg13g2_decap_8 FILLER_14_1085 ();
 sg13g2_fill_1 FILLER_14_1126 ();
 sg13g2_decap_8 FILLER_14_1136 ();
 sg13g2_decap_8 FILLER_14_1143 ();
 sg13g2_fill_2 FILLER_14_1150 ();
 sg13g2_fill_1 FILLER_14_1152 ();
 sg13g2_decap_4 FILLER_14_1193 ();
 sg13g2_decap_8 FILLER_14_1245 ();
 sg13g2_decap_8 FILLER_14_1252 ();
 sg13g2_decap_8 FILLER_14_1259 ();
 sg13g2_decap_4 FILLER_14_1266 ();
 sg13g2_fill_1 FILLER_14_1270 ();
 sg13g2_fill_2 FILLER_14_1275 ();
 sg13g2_fill_1 FILLER_14_1290 ();
 sg13g2_decap_8 FILLER_14_1341 ();
 sg13g2_fill_2 FILLER_14_1409 ();
 sg13g2_fill_1 FILLER_14_1429 ();
 sg13g2_fill_2 FILLER_14_1439 ();
 sg13g2_fill_1 FILLER_14_1452 ();
 sg13g2_fill_1 FILLER_14_1457 ();
 sg13g2_fill_1 FILLER_14_1462 ();
 sg13g2_fill_1 FILLER_14_1468 ();
 sg13g2_fill_1 FILLER_14_1473 ();
 sg13g2_fill_1 FILLER_14_1479 ();
 sg13g2_fill_1 FILLER_14_1484 ();
 sg13g2_fill_1 FILLER_14_1490 ();
 sg13g2_fill_1 FILLER_14_1519 ();
 sg13g2_fill_2 FILLER_14_1537 ();
 sg13g2_fill_2 FILLER_14_1545 ();
 sg13g2_fill_1 FILLER_14_1599 ();
 sg13g2_fill_2 FILLER_14_1609 ();
 sg13g2_fill_1 FILLER_14_1618 ();
 sg13g2_fill_2 FILLER_14_1719 ();
 sg13g2_fill_2 FILLER_14_1731 ();
 sg13g2_fill_1 FILLER_14_1733 ();
 sg13g2_fill_2 FILLER_14_1776 ();
 sg13g2_fill_1 FILLER_14_1778 ();
 sg13g2_fill_2 FILLER_14_1793 ();
 sg13g2_fill_2 FILLER_14_1807 ();
 sg13g2_fill_1 FILLER_14_1813 ();
 sg13g2_fill_1 FILLER_14_1824 ();
 sg13g2_decap_8 FILLER_14_1884 ();
 sg13g2_fill_2 FILLER_14_1891 ();
 sg13g2_fill_1 FILLER_14_1893 ();
 sg13g2_decap_4 FILLER_14_1904 ();
 sg13g2_fill_2 FILLER_14_1934 ();
 sg13g2_fill_2 FILLER_14_1975 ();
 sg13g2_fill_1 FILLER_14_1977 ();
 sg13g2_fill_2 FILLER_14_1988 ();
 sg13g2_fill_1 FILLER_14_1990 ();
 sg13g2_fill_1 FILLER_14_2016 ();
 sg13g2_fill_2 FILLER_14_2021 ();
 sg13g2_fill_1 FILLER_14_2053 ();
 sg13g2_fill_2 FILLER_14_2061 ();
 sg13g2_fill_1 FILLER_14_2083 ();
 sg13g2_fill_2 FILLER_14_2179 ();
 sg13g2_fill_1 FILLER_14_2228 ();
 sg13g2_decap_8 FILLER_14_2233 ();
 sg13g2_decap_8 FILLER_14_2289 ();
 sg13g2_decap_4 FILLER_14_2296 ();
 sg13g2_fill_2 FILLER_14_2300 ();
 sg13g2_decap_4 FILLER_14_2317 ();
 sg13g2_decap_8 FILLER_14_2357 ();
 sg13g2_fill_2 FILLER_14_2364 ();
 sg13g2_fill_1 FILLER_14_2366 ();
 sg13g2_fill_1 FILLER_14_2381 ();
 sg13g2_fill_1 FILLER_14_2387 ();
 sg13g2_decap_8 FILLER_14_2401 ();
 sg13g2_decap_4 FILLER_14_2408 ();
 sg13g2_fill_1 FILLER_14_2412 ();
 sg13g2_decap_4 FILLER_14_2439 ();
 sg13g2_fill_2 FILLER_14_2443 ();
 sg13g2_fill_1 FILLER_14_2462 ();
 sg13g2_fill_1 FILLER_14_2473 ();
 sg13g2_fill_1 FILLER_14_2484 ();
 sg13g2_decap_4 FILLER_14_2491 ();
 sg13g2_fill_2 FILLER_14_2506 ();
 sg13g2_fill_1 FILLER_14_2508 ();
 sg13g2_fill_1 FILLER_14_2519 ();
 sg13g2_decap_8 FILLER_14_2557 ();
 sg13g2_fill_1 FILLER_14_2564 ();
 sg13g2_fill_2 FILLER_14_2591 ();
 sg13g2_decap_4 FILLER_14_2616 ();
 sg13g2_decap_8 FILLER_14_2650 ();
 sg13g2_decap_8 FILLER_14_2657 ();
 sg13g2_decap_4 FILLER_14_2664 ();
 sg13g2_fill_2 FILLER_14_2668 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_14 ();
 sg13g2_fill_2 FILLER_15_52 ();
 sg13g2_fill_1 FILLER_15_54 ();
 sg13g2_fill_2 FILLER_15_81 ();
 sg13g2_fill_1 FILLER_15_83 ();
 sg13g2_fill_1 FILLER_15_117 ();
 sg13g2_fill_2 FILLER_15_139 ();
 sg13g2_fill_2 FILLER_15_148 ();
 sg13g2_fill_1 FILLER_15_164 ();
 sg13g2_fill_1 FILLER_15_214 ();
 sg13g2_fill_2 FILLER_15_223 ();
 sg13g2_fill_1 FILLER_15_251 ();
 sg13g2_fill_2 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_314 ();
 sg13g2_decap_8 FILLER_15_321 ();
 sg13g2_decap_8 FILLER_15_328 ();
 sg13g2_decap_8 FILLER_15_335 ();
 sg13g2_fill_2 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_fill_2 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_416 ();
 sg13g2_fill_1 FILLER_15_462 ();
 sg13g2_decap_4 FILLER_15_468 ();
 sg13g2_fill_2 FILLER_15_475 ();
 sg13g2_fill_1 FILLER_15_477 ();
 sg13g2_fill_2 FILLER_15_538 ();
 sg13g2_decap_8 FILLER_15_571 ();
 sg13g2_decap_8 FILLER_15_578 ();
 sg13g2_fill_2 FILLER_15_585 ();
 sg13g2_fill_1 FILLER_15_587 ();
 sg13g2_fill_2 FILLER_15_592 ();
 sg13g2_fill_1 FILLER_15_599 ();
 sg13g2_fill_2 FILLER_15_634 ();
 sg13g2_fill_1 FILLER_15_636 ();
 sg13g2_fill_2 FILLER_15_642 ();
 sg13g2_fill_1 FILLER_15_644 ();
 sg13g2_fill_1 FILLER_15_649 ();
 sg13g2_decap_4 FILLER_15_680 ();
 sg13g2_fill_1 FILLER_15_684 ();
 sg13g2_decap_8 FILLER_15_722 ();
 sg13g2_fill_2 FILLER_15_765 ();
 sg13g2_fill_1 FILLER_15_767 ();
 sg13g2_decap_8 FILLER_15_776 ();
 sg13g2_decap_4 FILLER_15_783 ();
 sg13g2_fill_1 FILLER_15_787 ();
 sg13g2_decap_4 FILLER_15_835 ();
 sg13g2_fill_1 FILLER_15_839 ();
 sg13g2_decap_4 FILLER_15_844 ();
 sg13g2_decap_8 FILLER_15_858 ();
 sg13g2_decap_4 FILLER_15_902 ();
 sg13g2_fill_2 FILLER_15_906 ();
 sg13g2_fill_2 FILLER_15_921 ();
 sg13g2_fill_1 FILLER_15_923 ();
 sg13g2_fill_1 FILLER_15_928 ();
 sg13g2_fill_1 FILLER_15_938 ();
 sg13g2_fill_1 FILLER_15_978 ();
 sg13g2_fill_1 FILLER_15_983 ();
 sg13g2_decap_4 FILLER_15_1040 ();
 sg13g2_decap_8 FILLER_15_1083 ();
 sg13g2_fill_1 FILLER_15_1090 ();
 sg13g2_decap_8 FILLER_15_1127 ();
 sg13g2_fill_2 FILLER_15_1134 ();
 sg13g2_fill_1 FILLER_15_1136 ();
 sg13g2_decap_4 FILLER_15_1177 ();
 sg13g2_fill_2 FILLER_15_1181 ();
 sg13g2_decap_4 FILLER_15_1188 ();
 sg13g2_fill_1 FILLER_15_1192 ();
 sg13g2_decap_4 FILLER_15_1198 ();
 sg13g2_fill_2 FILLER_15_1202 ();
 sg13g2_fill_2 FILLER_15_1216 ();
 sg13g2_fill_1 FILLER_15_1218 ();
 sg13g2_fill_2 FILLER_15_1257 ();
 sg13g2_fill_1 FILLER_15_1259 ();
 sg13g2_decap_8 FILLER_15_1296 ();
 sg13g2_fill_2 FILLER_15_1303 ();
 sg13g2_fill_1 FILLER_15_1305 ();
 sg13g2_decap_8 FILLER_15_1310 ();
 sg13g2_decap_8 FILLER_15_1317 ();
 sg13g2_decap_4 FILLER_15_1324 ();
 sg13g2_decap_8 FILLER_15_1338 ();
 sg13g2_decap_8 FILLER_15_1345 ();
 sg13g2_fill_1 FILLER_15_1352 ();
 sg13g2_fill_1 FILLER_15_1362 ();
 sg13g2_decap_8 FILLER_15_1371 ();
 sg13g2_fill_2 FILLER_15_1378 ();
 sg13g2_fill_1 FILLER_15_1385 ();
 sg13g2_fill_2 FILLER_15_1423 ();
 sg13g2_decap_4 FILLER_15_1435 ();
 sg13g2_decap_8 FILLER_15_1447 ();
 sg13g2_fill_2 FILLER_15_1454 ();
 sg13g2_fill_2 FILLER_15_1463 ();
 sg13g2_fill_1 FILLER_15_1470 ();
 sg13g2_fill_1 FILLER_15_1502 ();
 sg13g2_fill_1 FILLER_15_1508 ();
 sg13g2_fill_1 FILLER_15_1545 ();
 sg13g2_fill_1 FILLER_15_1592 ();
 sg13g2_fill_1 FILLER_15_1601 ();
 sg13g2_fill_1 FILLER_15_1672 ();
 sg13g2_decap_8 FILLER_15_1677 ();
 sg13g2_fill_2 FILLER_15_1715 ();
 sg13g2_fill_1 FILLER_15_1717 ();
 sg13g2_fill_1 FILLER_15_1769 ();
 sg13g2_fill_2 FILLER_15_1787 ();
 sg13g2_fill_1 FILLER_15_1789 ();
 sg13g2_decap_4 FILLER_15_1798 ();
 sg13g2_fill_2 FILLER_15_1802 ();
 sg13g2_decap_4 FILLER_15_1808 ();
 sg13g2_decap_8 FILLER_15_1816 ();
 sg13g2_decap_8 FILLER_15_1823 ();
 sg13g2_decap_4 FILLER_15_1830 ();
 sg13g2_fill_1 FILLER_15_1834 ();
 sg13g2_fill_2 FILLER_15_1839 ();
 sg13g2_decap_8 FILLER_15_1845 ();
 sg13g2_decap_4 FILLER_15_1852 ();
 sg13g2_decap_4 FILLER_15_1860 ();
 sg13g2_fill_2 FILLER_15_1864 ();
 sg13g2_fill_2 FILLER_15_1939 ();
 sg13g2_fill_1 FILLER_15_1941 ();
 sg13g2_decap_8 FILLER_15_1946 ();
 sg13g2_fill_2 FILLER_15_1953 ();
 sg13g2_decap_8 FILLER_15_1959 ();
 sg13g2_decap_8 FILLER_15_1966 ();
 sg13g2_fill_2 FILLER_15_2003 ();
 sg13g2_fill_1 FILLER_15_2062 ();
 sg13g2_fill_2 FILLER_15_2106 ();
 sg13g2_fill_2 FILLER_15_2122 ();
 sg13g2_fill_1 FILLER_15_2153 ();
 sg13g2_fill_2 FILLER_15_2195 ();
 sg13g2_decap_4 FILLER_15_2213 ();
 sg13g2_fill_1 FILLER_15_2217 ();
 sg13g2_decap_8 FILLER_15_2244 ();
 sg13g2_decap_4 FILLER_15_2251 ();
 sg13g2_fill_1 FILLER_15_2255 ();
 sg13g2_decap_4 FILLER_15_2281 ();
 sg13g2_fill_2 FILLER_15_2285 ();
 sg13g2_decap_8 FILLER_15_2317 ();
 sg13g2_decap_4 FILLER_15_2324 ();
 sg13g2_fill_2 FILLER_15_2328 ();
 sg13g2_decap_4 FILLER_15_2334 ();
 sg13g2_decap_8 FILLER_15_2352 ();
 sg13g2_decap_8 FILLER_15_2359 ();
 sg13g2_decap_8 FILLER_15_2366 ();
 sg13g2_fill_2 FILLER_15_2373 ();
 sg13g2_fill_2 FILLER_15_2381 ();
 sg13g2_fill_1 FILLER_15_2383 ();
 sg13g2_fill_2 FILLER_15_2394 ();
 sg13g2_fill_1 FILLER_15_2396 ();
 sg13g2_fill_1 FILLER_15_2401 ();
 sg13g2_fill_2 FILLER_15_2412 ();
 sg13g2_fill_2 FILLER_15_2420 ();
 sg13g2_fill_1 FILLER_15_2422 ();
 sg13g2_fill_1 FILLER_15_2433 ();
 sg13g2_fill_2 FILLER_15_2460 ();
 sg13g2_fill_2 FILLER_15_2466 ();
 sg13g2_fill_1 FILLER_15_2468 ();
 sg13g2_fill_1 FILLER_15_2495 ();
 sg13g2_fill_2 FILLER_15_2522 ();
 sg13g2_fill_1 FILLER_15_2524 ();
 sg13g2_fill_1 FILLER_15_2550 ();
 sg13g2_fill_1 FILLER_15_2587 ();
 sg13g2_fill_1 FILLER_15_2598 ();
 sg13g2_fill_2 FILLER_15_2605 ();
 sg13g2_decap_4 FILLER_15_2633 ();
 sg13g2_decap_8 FILLER_15_2663 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_fill_1 FILLER_16_72 ();
 sg13g2_fill_1 FILLER_16_86 ();
 sg13g2_fill_1 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_96 ();
 sg13g2_fill_1 FILLER_16_102 ();
 sg13g2_fill_2 FILLER_16_108 ();
 sg13g2_fill_1 FILLER_16_115 ();
 sg13g2_fill_1 FILLER_16_136 ();
 sg13g2_fill_1 FILLER_16_156 ();
 sg13g2_fill_2 FILLER_16_168 ();
 sg13g2_fill_2 FILLER_16_175 ();
 sg13g2_fill_1 FILLER_16_181 ();
 sg13g2_fill_1 FILLER_16_213 ();
 sg13g2_fill_2 FILLER_16_218 ();
 sg13g2_fill_2 FILLER_16_224 ();
 sg13g2_decap_4 FILLER_16_235 ();
 sg13g2_fill_1 FILLER_16_239 ();
 sg13g2_fill_1 FILLER_16_255 ();
 sg13g2_decap_4 FILLER_16_322 ();
 sg13g2_fill_1 FILLER_16_368 ();
 sg13g2_fill_1 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_412 ();
 sg13g2_fill_1 FILLER_16_422 ();
 sg13g2_fill_1 FILLER_16_431 ();
 sg13g2_fill_1 FILLER_16_439 ();
 sg13g2_fill_1 FILLER_16_461 ();
 sg13g2_decap_8 FILLER_16_488 ();
 sg13g2_decap_8 FILLER_16_495 ();
 sg13g2_decap_8 FILLER_16_506 ();
 sg13g2_fill_2 FILLER_16_513 ();
 sg13g2_fill_1 FILLER_16_515 ();
 sg13g2_decap_4 FILLER_16_520 ();
 sg13g2_fill_2 FILLER_16_528 ();
 sg13g2_fill_1 FILLER_16_539 ();
 sg13g2_fill_1 FILLER_16_544 ();
 sg13g2_decap_8 FILLER_16_580 ();
 sg13g2_fill_1 FILLER_16_629 ();
 sg13g2_decap_8 FILLER_16_641 ();
 sg13g2_decap_8 FILLER_16_648 ();
 sg13g2_decap_8 FILLER_16_659 ();
 sg13g2_decap_4 FILLER_16_676 ();
 sg13g2_fill_2 FILLER_16_765 ();
 sg13g2_decap_8 FILLER_16_799 ();
 sg13g2_fill_1 FILLER_16_806 ();
 sg13g2_decap_8 FILLER_16_828 ();
 sg13g2_fill_2 FILLER_16_835 ();
 sg13g2_fill_1 FILLER_16_837 ();
 sg13g2_decap_4 FILLER_16_864 ();
 sg13g2_fill_2 FILLER_16_898 ();
 sg13g2_fill_1 FILLER_16_900 ();
 sg13g2_fill_1 FILLER_16_911 ();
 sg13g2_fill_2 FILLER_16_916 ();
 sg13g2_fill_1 FILLER_16_918 ();
 sg13g2_fill_1 FILLER_16_933 ();
 sg13g2_decap_8 FILLER_16_997 ();
 sg13g2_fill_2 FILLER_16_1004 ();
 sg13g2_fill_1 FILLER_16_1006 ();
 sg13g2_fill_2 FILLER_16_1042 ();
 sg13g2_fill_1 FILLER_16_1048 ();
 sg13g2_decap_8 FILLER_16_1089 ();
 sg13g2_fill_2 FILLER_16_1096 ();
 sg13g2_decap_4 FILLER_16_1103 ();
 sg13g2_fill_1 FILLER_16_1107 ();
 sg13g2_fill_2 FILLER_16_1137 ();
 sg13g2_fill_1 FILLER_16_1139 ();
 sg13g2_fill_1 FILLER_16_1145 ();
 sg13g2_decap_8 FILLER_16_1172 ();
 sg13g2_decap_8 FILLER_16_1179 ();
 sg13g2_fill_1 FILLER_16_1194 ();
 sg13g2_fill_1 FILLER_16_1221 ();
 sg13g2_fill_2 FILLER_16_1226 ();
 sg13g2_fill_1 FILLER_16_1228 ();
 sg13g2_fill_2 FILLER_16_1259 ();
 sg13g2_fill_1 FILLER_16_1261 ();
 sg13g2_decap_4 FILLER_16_1272 ();
 sg13g2_fill_1 FILLER_16_1276 ();
 sg13g2_decap_8 FILLER_16_1281 ();
 sg13g2_decap_8 FILLER_16_1298 ();
 sg13g2_decap_8 FILLER_16_1305 ();
 sg13g2_decap_4 FILLER_16_1357 ();
 sg13g2_decap_4 FILLER_16_1366 ();
 sg13g2_fill_1 FILLER_16_1370 ();
 sg13g2_decap_4 FILLER_16_1375 ();
 sg13g2_fill_1 FILLER_16_1379 ();
 sg13g2_fill_1 FILLER_16_1390 ();
 sg13g2_fill_1 FILLER_16_1396 ();
 sg13g2_fill_1 FILLER_16_1401 ();
 sg13g2_fill_1 FILLER_16_1428 ();
 sg13g2_fill_2 FILLER_16_1434 ();
 sg13g2_fill_1 FILLER_16_1445 ();
 sg13g2_fill_2 FILLER_16_1497 ();
 sg13g2_fill_1 FILLER_16_1591 ();
 sg13g2_fill_1 FILLER_16_1597 ();
 sg13g2_fill_2 FILLER_16_1637 ();
 sg13g2_fill_1 FILLER_16_1668 ();
 sg13g2_fill_2 FILLER_16_1684 ();
 sg13g2_fill_1 FILLER_16_1686 ();
 sg13g2_decap_8 FILLER_16_1733 ();
 sg13g2_decap_8 FILLER_16_1740 ();
 sg13g2_fill_1 FILLER_16_1747 ();
 sg13g2_fill_2 FILLER_16_1760 ();
 sg13g2_fill_1 FILLER_16_1767 ();
 sg13g2_fill_2 FILLER_16_1774 ();
 sg13g2_fill_2 FILLER_16_1799 ();
 sg13g2_fill_1 FILLER_16_1801 ();
 sg13g2_decap_8 FILLER_16_1825 ();
 sg13g2_fill_2 FILLER_16_1832 ();
 sg13g2_fill_1 FILLER_16_1834 ();
 sg13g2_fill_1 FILLER_16_1849 ();
 sg13g2_fill_2 FILLER_16_1876 ();
 sg13g2_fill_1 FILLER_16_1995 ();
 sg13g2_decap_4 FILLER_16_2000 ();
 sg13g2_fill_1 FILLER_16_2004 ();
 sg13g2_fill_2 FILLER_16_2031 ();
 sg13g2_fill_2 FILLER_16_2061 ();
 sg13g2_fill_1 FILLER_16_2102 ();
 sg13g2_fill_1 FILLER_16_2124 ();
 sg13g2_fill_2 FILLER_16_2135 ();
 sg13g2_decap_8 FILLER_16_2239 ();
 sg13g2_fill_2 FILLER_16_2246 ();
 sg13g2_decap_4 FILLER_16_2258 ();
 sg13g2_fill_1 FILLER_16_2292 ();
 sg13g2_fill_2 FILLER_16_2323 ();
 sg13g2_fill_1 FILLER_16_2325 ();
 sg13g2_decap_8 FILLER_16_2343 ();
 sg13g2_fill_1 FILLER_16_2350 ();
 sg13g2_fill_1 FILLER_16_2377 ();
 sg13g2_fill_2 FILLER_16_2388 ();
 sg13g2_fill_2 FILLER_16_2421 ();
 sg13g2_fill_1 FILLER_16_2423 ();
 sg13g2_decap_4 FILLER_16_2484 ();
 sg13g2_fill_1 FILLER_16_2488 ();
 sg13g2_fill_1 FILLER_16_2495 ();
 sg13g2_decap_4 FILLER_16_2502 ();
 sg13g2_fill_2 FILLER_16_2506 ();
 sg13g2_fill_1 FILLER_16_2512 ();
 sg13g2_fill_1 FILLER_16_2521 ();
 sg13g2_decap_8 FILLER_16_2527 ();
 sg13g2_decap_8 FILLER_16_2573 ();
 sg13g2_decap_4 FILLER_16_2580 ();
 sg13g2_fill_2 FILLER_16_2584 ();
 sg13g2_fill_1 FILLER_16_2598 ();
 sg13g2_fill_2 FILLER_16_2668 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_4 ();
 sg13g2_fill_2 FILLER_17_68 ();
 sg13g2_decap_8 FILLER_17_104 ();
 sg13g2_decap_4 FILLER_17_116 ();
 sg13g2_fill_2 FILLER_17_120 ();
 sg13g2_decap_4 FILLER_17_127 ();
 sg13g2_fill_1 FILLER_17_131 ();
 sg13g2_fill_1 FILLER_17_192 ();
 sg13g2_fill_2 FILLER_17_215 ();
 sg13g2_fill_1 FILLER_17_217 ();
 sg13g2_fill_2 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_238 ();
 sg13g2_decap_4 FILLER_17_243 ();
 sg13g2_fill_1 FILLER_17_247 ();
 sg13g2_fill_1 FILLER_17_253 ();
 sg13g2_fill_2 FILLER_17_318 ();
 sg13g2_fill_1 FILLER_17_320 ();
 sg13g2_decap_4 FILLER_17_326 ();
 sg13g2_fill_1 FILLER_17_330 ();
 sg13g2_decap_4 FILLER_17_335 ();
 sg13g2_fill_1 FILLER_17_353 ();
 sg13g2_fill_1 FILLER_17_369 ();
 sg13g2_fill_2 FILLER_17_374 ();
 sg13g2_fill_2 FILLER_17_385 ();
 sg13g2_fill_1 FILLER_17_391 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_2 FILLER_17_480 ();
 sg13g2_fill_1 FILLER_17_482 ();
 sg13g2_decap_4 FILLER_17_491 ();
 sg13g2_decap_8 FILLER_17_499 ();
 sg13g2_decap_4 FILLER_17_506 ();
 sg13g2_decap_8 FILLER_17_514 ();
 sg13g2_fill_1 FILLER_17_521 ();
 sg13g2_fill_2 FILLER_17_526 ();
 sg13g2_fill_1 FILLER_17_528 ();
 sg13g2_fill_2 FILLER_17_573 ();
 sg13g2_fill_2 FILLER_17_595 ();
 sg13g2_fill_1 FILLER_17_597 ();
 sg13g2_fill_2 FILLER_17_620 ();
 sg13g2_fill_1 FILLER_17_648 ();
 sg13g2_fill_1 FILLER_17_685 ();
 sg13g2_decap_4 FILLER_17_726 ();
 sg13g2_fill_2 FILLER_17_770 ();
 sg13g2_fill_2 FILLER_17_798 ();
 sg13g2_fill_1 FILLER_17_800 ();
 sg13g2_fill_2 FILLER_17_827 ();
 sg13g2_fill_1 FILLER_17_829 ();
 sg13g2_fill_2 FILLER_17_866 ();
 sg13g2_fill_1 FILLER_17_868 ();
 sg13g2_fill_2 FILLER_17_886 ();
 sg13g2_fill_2 FILLER_17_922 ();
 sg13g2_fill_1 FILLER_17_950 ();
 sg13g2_fill_1 FILLER_17_956 ();
 sg13g2_fill_2 FILLER_17_961 ();
 sg13g2_fill_2 FILLER_17_973 ();
 sg13g2_decap_8 FILLER_17_1000 ();
 sg13g2_decap_8 FILLER_17_1007 ();
 sg13g2_fill_1 FILLER_17_1014 ();
 sg13g2_fill_2 FILLER_17_1074 ();
 sg13g2_fill_1 FILLER_17_1097 ();
 sg13g2_decap_8 FILLER_17_1178 ();
 sg13g2_decap_8 FILLER_17_1234 ();
 sg13g2_fill_1 FILLER_17_1245 ();
 sg13g2_fill_2 FILLER_17_1276 ();
 sg13g2_fill_1 FILLER_17_1278 ();
 sg13g2_fill_2 FILLER_17_1334 ();
 sg13g2_decap_4 FILLER_17_1362 ();
 sg13g2_fill_2 FILLER_17_1392 ();
 sg13g2_decap_4 FILLER_17_1420 ();
 sg13g2_fill_1 FILLER_17_1453 ();
 sg13g2_fill_1 FILLER_17_1466 ();
 sg13g2_fill_1 FILLER_17_1483 ();
 sg13g2_fill_2 FILLER_17_1494 ();
 sg13g2_fill_2 FILLER_17_1506 ();
 sg13g2_fill_2 FILLER_17_1572 ();
 sg13g2_fill_1 FILLER_17_1591 ();
 sg13g2_fill_1 FILLER_17_1600 ();
 sg13g2_fill_2 FILLER_17_1606 ();
 sg13g2_fill_2 FILLER_17_1616 ();
 sg13g2_fill_2 FILLER_17_1632 ();
 sg13g2_decap_8 FILLER_17_1663 ();
 sg13g2_fill_1 FILLER_17_1670 ();
 sg13g2_decap_4 FILLER_17_1680 ();
 sg13g2_fill_1 FILLER_17_1706 ();
 sg13g2_decap_8 FILLER_17_1725 ();
 sg13g2_decap_4 FILLER_17_1732 ();
 sg13g2_fill_2 FILLER_17_1736 ();
 sg13g2_decap_4 FILLER_17_1742 ();
 sg13g2_fill_1 FILLER_17_1746 ();
 sg13g2_fill_2 FILLER_17_1751 ();
 sg13g2_fill_1 FILLER_17_1753 ();
 sg13g2_decap_4 FILLER_17_1758 ();
 sg13g2_fill_1 FILLER_17_1762 ();
 sg13g2_fill_1 FILLER_17_1773 ();
 sg13g2_fill_2 FILLER_17_1779 ();
 sg13g2_fill_1 FILLER_17_1786 ();
 sg13g2_fill_1 FILLER_17_1813 ();
 sg13g2_fill_2 FILLER_17_1840 ();
 sg13g2_fill_1 FILLER_17_1868 ();
 sg13g2_fill_1 FILLER_17_1895 ();
 sg13g2_fill_1 FILLER_17_1906 ();
 sg13g2_fill_2 FILLER_17_1911 ();
 sg13g2_fill_1 FILLER_17_1975 ();
 sg13g2_fill_1 FILLER_17_2028 ();
 sg13g2_fill_2 FILLER_17_2041 ();
 sg13g2_fill_1 FILLER_17_2073 ();
 sg13g2_fill_1 FILLER_17_2078 ();
 sg13g2_fill_1 FILLER_17_2094 ();
 sg13g2_fill_2 FILLER_17_2170 ();
 sg13g2_fill_1 FILLER_17_2172 ();
 sg13g2_fill_1 FILLER_17_2177 ();
 sg13g2_fill_1 FILLER_17_2182 ();
 sg13g2_fill_1 FILLER_17_2209 ();
 sg13g2_fill_1 FILLER_17_2246 ();
 sg13g2_decap_8 FILLER_17_2287 ();
 sg13g2_decap_4 FILLER_17_2294 ();
 sg13g2_decap_4 FILLER_17_2331 ();
 sg13g2_decap_4 FILLER_17_2365 ();
 sg13g2_fill_1 FILLER_17_2399 ();
 sg13g2_fill_1 FILLER_17_2426 ();
 sg13g2_fill_1 FILLER_17_2437 ();
 sg13g2_fill_1 FILLER_17_2442 ();
 sg13g2_decap_8 FILLER_17_2447 ();
 sg13g2_decap_8 FILLER_17_2454 ();
 sg13g2_decap_8 FILLER_17_2461 ();
 sg13g2_fill_1 FILLER_17_2468 ();
 sg13g2_decap_8 FILLER_17_2479 ();
 sg13g2_fill_1 FILLER_17_2486 ();
 sg13g2_fill_2 FILLER_17_2501 ();
 sg13g2_decap_4 FILLER_17_2529 ();
 sg13g2_fill_2 FILLER_17_2543 ();
 sg13g2_fill_1 FILLER_17_2554 ();
 sg13g2_fill_1 FILLER_17_2568 ();
 sg13g2_decap_4 FILLER_17_2582 ();
 sg13g2_fill_1 FILLER_17_2595 ();
 sg13g2_decap_8 FILLER_17_2631 ();
 sg13g2_fill_1 FILLER_17_2669 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_19 ();
 sg13g2_fill_1 FILLER_18_25 ();
 sg13g2_fill_2 FILLER_18_39 ();
 sg13g2_fill_2 FILLER_18_58 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_fill_1 FILLER_18_69 ();
 sg13g2_fill_2 FILLER_18_86 ();
 sg13g2_fill_1 FILLER_18_97 ();
 sg13g2_fill_2 FILLER_18_108 ();
 sg13g2_fill_1 FILLER_18_110 ();
 sg13g2_fill_1 FILLER_18_159 ();
 sg13g2_fill_2 FILLER_18_173 ();
 sg13g2_fill_1 FILLER_18_175 ();
 sg13g2_fill_1 FILLER_18_186 ();
 sg13g2_fill_1 FILLER_18_192 ();
 sg13g2_decap_4 FILLER_18_231 ();
 sg13g2_fill_1 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_240 ();
 sg13g2_decap_8 FILLER_18_247 ();
 sg13g2_fill_2 FILLER_18_254 ();
 sg13g2_fill_2 FILLER_18_271 ();
 sg13g2_fill_1 FILLER_18_281 ();
 sg13g2_fill_1 FILLER_18_286 ();
 sg13g2_decap_4 FILLER_18_322 ();
 sg13g2_fill_1 FILLER_18_326 ();
 sg13g2_fill_2 FILLER_18_369 ();
 sg13g2_fill_2 FILLER_18_383 ();
 sg13g2_fill_1 FILLER_18_385 ();
 sg13g2_fill_1 FILLER_18_391 ();
 sg13g2_fill_2 FILLER_18_397 ();
 sg13g2_fill_1 FILLER_18_419 ();
 sg13g2_fill_1 FILLER_18_424 ();
 sg13g2_fill_2 FILLER_18_430 ();
 sg13g2_fill_2 FILLER_18_436 ();
 sg13g2_fill_2 FILLER_18_456 ();
 sg13g2_fill_2 FILLER_18_463 ();
 sg13g2_fill_1 FILLER_18_465 ();
 sg13g2_fill_1 FILLER_18_470 ();
 sg13g2_fill_1 FILLER_18_475 ();
 sg13g2_fill_1 FILLER_18_480 ();
 sg13g2_fill_2 FILLER_18_486 ();
 sg13g2_fill_2 FILLER_18_492 ();
 sg13g2_decap_8 FILLER_18_520 ();
 sg13g2_fill_2 FILLER_18_539 ();
 sg13g2_fill_1 FILLER_18_541 ();
 sg13g2_decap_8 FILLER_18_550 ();
 sg13g2_decap_8 FILLER_18_557 ();
 sg13g2_decap_4 FILLER_18_564 ();
 sg13g2_fill_1 FILLER_18_568 ();
 sg13g2_fill_1 FILLER_18_580 ();
 sg13g2_fill_2 FILLER_18_587 ();
 sg13g2_fill_1 FILLER_18_670 ();
 sg13g2_decap_8 FILLER_18_675 ();
 sg13g2_decap_8 FILLER_18_682 ();
 sg13g2_decap_8 FILLER_18_689 ();
 sg13g2_decap_8 FILLER_18_696 ();
 sg13g2_fill_2 FILLER_18_703 ();
 sg13g2_fill_1 FILLER_18_719 ();
 sg13g2_decap_8 FILLER_18_730 ();
 sg13g2_fill_2 FILLER_18_737 ();
 sg13g2_fill_1 FILLER_18_743 ();
 sg13g2_decap_8 FILLER_18_800 ();
 sg13g2_fill_2 FILLER_18_807 ();
 sg13g2_fill_2 FILLER_18_856 ();
 sg13g2_fill_1 FILLER_18_868 ();
 sg13g2_decap_8 FILLER_18_875 ();
 sg13g2_fill_1 FILLER_18_887 ();
 sg13g2_fill_1 FILLER_18_893 ();
 sg13g2_fill_2 FILLER_18_899 ();
 sg13g2_fill_1 FILLER_18_937 ();
 sg13g2_fill_1 FILLER_18_943 ();
 sg13g2_fill_2 FILLER_18_948 ();
 sg13g2_decap_4 FILLER_18_991 ();
 sg13g2_fill_1 FILLER_18_995 ();
 sg13g2_decap_8 FILLER_18_1000 ();
 sg13g2_decap_8 FILLER_18_1007 ();
 sg13g2_decap_4 FILLER_18_1014 ();
 sg13g2_fill_2 FILLER_18_1018 ();
 sg13g2_decap_4 FILLER_18_1024 ();
 sg13g2_fill_1 FILLER_18_1032 ();
 sg13g2_fill_2 FILLER_18_1065 ();
 sg13g2_fill_1 FILLER_18_1067 ();
 sg13g2_decap_8 FILLER_18_1076 ();
 sg13g2_fill_1 FILLER_18_1083 ();
 sg13g2_fill_1 FILLER_18_1092 ();
 sg13g2_fill_2 FILLER_18_1128 ();
 sg13g2_fill_1 FILLER_18_1130 ();
 sg13g2_fill_2 FILLER_18_1157 ();
 sg13g2_decap_4 FILLER_18_1184 ();
 sg13g2_fill_2 FILLER_18_1188 ();
 sg13g2_decap_4 FILLER_18_1263 ();
 sg13g2_fill_2 FILLER_18_1293 ();
 sg13g2_fill_2 FILLER_18_1342 ();
 sg13g2_fill_2 FILLER_18_1348 ();
 sg13g2_fill_1 FILLER_18_1350 ();
 sg13g2_decap_8 FILLER_18_1355 ();
 sg13g2_decap_8 FILLER_18_1362 ();
 sg13g2_decap_8 FILLER_18_1369 ();
 sg13g2_fill_1 FILLER_18_1430 ();
 sg13g2_fill_2 FILLER_18_1434 ();
 sg13g2_fill_1 FILLER_18_1496 ();
 sg13g2_fill_1 FILLER_18_1510 ();
 sg13g2_fill_1 FILLER_18_1525 ();
 sg13g2_fill_1 FILLER_18_1555 ();
 sg13g2_fill_1 FILLER_18_1616 ();
 sg13g2_fill_1 FILLER_18_1622 ();
 sg13g2_fill_1 FILLER_18_1635 ();
 sg13g2_fill_1 FILLER_18_1643 ();
 sg13g2_decap_8 FILLER_18_1658 ();
 sg13g2_decap_4 FILLER_18_1665 ();
 sg13g2_fill_1 FILLER_18_1669 ();
 sg13g2_decap_8 FILLER_18_1686 ();
 sg13g2_fill_2 FILLER_18_1693 ();
 sg13g2_fill_1 FILLER_18_1695 ();
 sg13g2_fill_1 FILLER_18_1708 ();
 sg13g2_decap_8 FILLER_18_1714 ();
 sg13g2_decap_4 FILLER_18_1811 ();
 sg13g2_fill_1 FILLER_18_1815 ();
 sg13g2_fill_2 FILLER_18_1847 ();
 sg13g2_fill_1 FILLER_18_1849 ();
 sg13g2_fill_2 FILLER_18_1860 ();
 sg13g2_fill_1 FILLER_18_1876 ();
 sg13g2_decap_8 FILLER_18_1881 ();
 sg13g2_decap_8 FILLER_18_1888 ();
 sg13g2_decap_8 FILLER_18_1895 ();
 sg13g2_fill_2 FILLER_18_1902 ();
 sg13g2_fill_1 FILLER_18_1904 ();
 sg13g2_decap_4 FILLER_18_1915 ();
 sg13g2_fill_1 FILLER_18_1919 ();
 sg13g2_decap_8 FILLER_18_1924 ();
 sg13g2_fill_2 FILLER_18_1931 ();
 sg13g2_fill_2 FILLER_18_1950 ();
 sg13g2_fill_2 FILLER_18_1956 ();
 sg13g2_fill_2 FILLER_18_1994 ();
 sg13g2_fill_1 FILLER_18_2012 ();
 sg13g2_fill_1 FILLER_18_2016 ();
 sg13g2_fill_1 FILLER_18_2025 ();
 sg13g2_fill_1 FILLER_18_2112 ();
 sg13g2_decap_4 FILLER_18_2175 ();
 sg13g2_fill_1 FILLER_18_2198 ();
 sg13g2_decap_4 FILLER_18_2234 ();
 sg13g2_fill_2 FILLER_18_2238 ();
 sg13g2_decap_8 FILLER_18_2276 ();
 sg13g2_decap_8 FILLER_18_2283 ();
 sg13g2_decap_8 FILLER_18_2290 ();
 sg13g2_decap_8 FILLER_18_2297 ();
 sg13g2_decap_4 FILLER_18_2304 ();
 sg13g2_decap_8 FILLER_18_2347 ();
 sg13g2_decap_4 FILLER_18_2354 ();
 sg13g2_fill_2 FILLER_18_2358 ();
 sg13g2_decap_4 FILLER_18_2364 ();
 sg13g2_fill_1 FILLER_18_2373 ();
 sg13g2_fill_1 FILLER_18_2419 ();
 sg13g2_decap_8 FILLER_18_2444 ();
 sg13g2_fill_1 FILLER_18_2451 ();
 sg13g2_decap_8 FILLER_18_2457 ();
 sg13g2_decap_8 FILLER_18_2464 ();
 sg13g2_decap_4 FILLER_18_2471 ();
 sg13g2_fill_2 FILLER_18_2534 ();
 sg13g2_decap_4 FILLER_18_2585 ();
 sg13g2_decap_8 FILLER_18_2592 ();
 sg13g2_fill_2 FILLER_18_2620 ();
 sg13g2_fill_1 FILLER_18_2622 ();
 sg13g2_decap_4 FILLER_18_2633 ();
 sg13g2_fill_1 FILLER_18_2637 ();
 sg13g2_fill_2 FILLER_18_2668 ();
 sg13g2_decap_8 FILLER_19_45 ();
 sg13g2_decap_8 FILLER_19_52 ();
 sg13g2_decap_4 FILLER_19_59 ();
 sg13g2_fill_2 FILLER_19_63 ();
 sg13g2_fill_1 FILLER_19_78 ();
 sg13g2_fill_1 FILLER_19_92 ();
 sg13g2_fill_2 FILLER_19_175 ();
 sg13g2_fill_1 FILLER_19_182 ();
 sg13g2_fill_1 FILLER_19_231 ();
 sg13g2_fill_1 FILLER_19_304 ();
 sg13g2_fill_1 FILLER_19_329 ();
 sg13g2_fill_1 FILLER_19_369 ();
 sg13g2_fill_1 FILLER_19_389 ();
 sg13g2_fill_2 FILLER_19_395 ();
 sg13g2_fill_2 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_413 ();
 sg13g2_fill_2 FILLER_19_422 ();
 sg13g2_fill_2 FILLER_19_458 ();
 sg13g2_fill_1 FILLER_19_460 ();
 sg13g2_fill_2 FILLER_19_465 ();
 sg13g2_fill_1 FILLER_19_467 ();
 sg13g2_fill_1 FILLER_19_568 ();
 sg13g2_fill_1 FILLER_19_574 ();
 sg13g2_fill_2 FILLER_19_596 ();
 sg13g2_fill_1 FILLER_19_598 ();
 sg13g2_fill_2 FILLER_19_604 ();
 sg13g2_fill_1 FILLER_19_617 ();
 sg13g2_fill_1 FILLER_19_622 ();
 sg13g2_fill_1 FILLER_19_637 ();
 sg13g2_fill_1 FILLER_19_646 ();
 sg13g2_fill_2 FILLER_19_667 ();
 sg13g2_fill_1 FILLER_19_669 ();
 sg13g2_decap_8 FILLER_19_674 ();
 sg13g2_decap_4 FILLER_19_681 ();
 sg13g2_fill_1 FILLER_19_685 ();
 sg13g2_decap_4 FILLER_19_695 ();
 sg13g2_fill_2 FILLER_19_699 ();
 sg13g2_fill_2 FILLER_19_727 ();
 sg13g2_fill_2 FILLER_19_739 ();
 sg13g2_fill_1 FILLER_19_741 ();
 sg13g2_fill_2 FILLER_19_752 ();
 sg13g2_fill_1 FILLER_19_754 ();
 sg13g2_fill_2 FILLER_19_765 ();
 sg13g2_decap_4 FILLER_19_813 ();
 sg13g2_decap_4 FILLER_19_827 ();
 sg13g2_fill_1 FILLER_19_831 ();
 sg13g2_fill_1 FILLER_19_842 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_fill_2 FILLER_19_854 ();
 sg13g2_fill_2 FILLER_19_882 ();
 sg13g2_fill_1 FILLER_19_884 ();
 sg13g2_fill_1 FILLER_19_893 ();
 sg13g2_fill_1 FILLER_19_920 ();
 sg13g2_fill_2 FILLER_19_925 ();
 sg13g2_fill_2 FILLER_19_948 ();
 sg13g2_decap_4 FILLER_19_1014 ();
 sg13g2_fill_2 FILLER_19_1018 ();
 sg13g2_fill_2 FILLER_19_1146 ();
 sg13g2_fill_1 FILLER_19_1148 ();
 sg13g2_fill_1 FILLER_19_1161 ();
 sg13g2_decap_8 FILLER_19_1170 ();
 sg13g2_decap_8 FILLER_19_1177 ();
 sg13g2_decap_8 FILLER_19_1184 ();
 sg13g2_decap_8 FILLER_19_1191 ();
 sg13g2_fill_2 FILLER_19_1198 ();
 sg13g2_fill_2 FILLER_19_1204 ();
 sg13g2_fill_2 FILLER_19_1210 ();
 sg13g2_fill_1 FILLER_19_1212 ();
 sg13g2_fill_2 FILLER_19_1217 ();
 sg13g2_fill_1 FILLER_19_1219 ();
 sg13g2_fill_2 FILLER_19_1225 ();
 sg13g2_fill_1 FILLER_19_1227 ();
 sg13g2_decap_8 FILLER_19_1254 ();
 sg13g2_fill_2 FILLER_19_1261 ();
 sg13g2_fill_1 FILLER_19_1263 ();
 sg13g2_decap_4 FILLER_19_1277 ();
 sg13g2_fill_2 FILLER_19_1281 ();
 sg13g2_fill_2 FILLER_19_1287 ();
 sg13g2_fill_1 FILLER_19_1289 ();
 sg13g2_fill_2 FILLER_19_1300 ();
 sg13g2_decap_4 FILLER_19_1306 ();
 sg13g2_decap_8 FILLER_19_1359 ();
 sg13g2_decap_4 FILLER_19_1366 ();
 sg13g2_fill_1 FILLER_19_1370 ();
 sg13g2_fill_1 FILLER_19_1375 ();
 sg13g2_fill_1 FILLER_19_1402 ();
 sg13g2_fill_2 FILLER_19_1454 ();
 sg13g2_fill_1 FILLER_19_1459 ();
 sg13g2_fill_1 FILLER_19_1463 ();
 sg13g2_fill_2 FILLER_19_1495 ();
 sg13g2_fill_2 FILLER_19_1554 ();
 sg13g2_fill_2 FILLER_19_1559 ();
 sg13g2_fill_1 FILLER_19_1565 ();
 sg13g2_fill_1 FILLER_19_1602 ();
 sg13g2_fill_1 FILLER_19_1685 ();
 sg13g2_decap_4 FILLER_19_1694 ();
 sg13g2_fill_2 FILLER_19_1698 ();
 sg13g2_fill_2 FILLER_19_1726 ();
 sg13g2_fill_1 FILLER_19_1728 ();
 sg13g2_decap_4 FILLER_19_1787 ();
 sg13g2_decap_8 FILLER_19_1840 ();
 sg13g2_decap_8 FILLER_19_1847 ();
 sg13g2_decap_8 FILLER_19_1854 ();
 sg13g2_decap_8 FILLER_19_1861 ();
 sg13g2_decap_8 FILLER_19_1868 ();
 sg13g2_decap_8 FILLER_19_1875 ();
 sg13g2_decap_8 FILLER_19_1882 ();
 sg13g2_decap_4 FILLER_19_1889 ();
 sg13g2_fill_1 FILLER_19_1893 ();
 sg13g2_fill_2 FILLER_19_1897 ();
 sg13g2_decap_8 FILLER_19_1916 ();
 sg13g2_decap_8 FILLER_19_1923 ();
 sg13g2_decap_4 FILLER_19_1930 ();
 sg13g2_decap_8 FILLER_19_1939 ();
 sg13g2_decap_4 FILLER_19_1950 ();
 sg13g2_fill_1 FILLER_19_1954 ();
 sg13g2_decap_8 FILLER_19_1969 ();
 sg13g2_decap_8 FILLER_19_1986 ();
 sg13g2_fill_2 FILLER_19_1993 ();
 sg13g2_fill_1 FILLER_19_2005 ();
 sg13g2_fill_2 FILLER_19_2027 ();
 sg13g2_fill_1 FILLER_19_2036 ();
 sg13g2_fill_2 FILLER_19_2051 ();
 sg13g2_decap_4 FILLER_19_2081 ();
 sg13g2_fill_2 FILLER_19_2159 ();
 sg13g2_fill_1 FILLER_19_2161 ();
 sg13g2_fill_2 FILLER_19_2172 ();
 sg13g2_fill_1 FILLER_19_2174 ();
 sg13g2_decap_4 FILLER_19_2211 ();
 sg13g2_fill_2 FILLER_19_2215 ();
 sg13g2_decap_8 FILLER_19_2243 ();
 sg13g2_decap_4 FILLER_19_2250 ();
 sg13g2_fill_2 FILLER_19_2254 ();
 sg13g2_decap_8 FILLER_19_2260 ();
 sg13g2_decap_8 FILLER_19_2267 ();
 sg13g2_fill_2 FILLER_19_2274 ();
 sg13g2_decap_4 FILLER_19_2329 ();
 sg13g2_fill_2 FILLER_19_2333 ();
 sg13g2_decap_8 FILLER_19_2339 ();
 sg13g2_decap_4 FILLER_19_2346 ();
 sg13g2_fill_1 FILLER_19_2350 ();
 sg13g2_decap_8 FILLER_19_2360 ();
 sg13g2_fill_1 FILLER_19_2367 ();
 sg13g2_decap_4 FILLER_19_2378 ();
 sg13g2_fill_1 FILLER_19_2382 ();
 sg13g2_decap_8 FILLER_19_2396 ();
 sg13g2_decap_4 FILLER_19_2403 ();
 sg13g2_fill_1 FILLER_19_2407 ();
 sg13g2_decap_8 FILLER_19_2413 ();
 sg13g2_decap_4 FILLER_19_2420 ();
 sg13g2_fill_2 FILLER_19_2424 ();
 sg13g2_decap_8 FILLER_19_2430 ();
 sg13g2_fill_2 FILLER_19_2437 ();
 sg13g2_fill_1 FILLER_19_2439 ();
 sg13g2_fill_2 FILLER_19_2450 ();
 sg13g2_fill_2 FILLER_19_2456 ();
 sg13g2_fill_2 FILLER_19_2468 ();
 sg13g2_fill_1 FILLER_19_2470 ();
 sg13g2_fill_2 FILLER_19_2480 ();
 sg13g2_fill_1 FILLER_19_2482 ();
 sg13g2_fill_2 FILLER_19_2493 ();
 sg13g2_fill_1 FILLER_19_2495 ();
 sg13g2_fill_1 FILLER_19_2506 ();
 sg13g2_fill_2 FILLER_19_2517 ();
 sg13g2_fill_2 FILLER_19_2544 ();
 sg13g2_decap_8 FILLER_19_2604 ();
 sg13g2_fill_1 FILLER_19_2617 ();
 sg13g2_fill_1 FILLER_19_2622 ();
 sg13g2_fill_2 FILLER_19_2633 ();
 sg13g2_decap_8 FILLER_19_2661 ();
 sg13g2_fill_2 FILLER_19_2668 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_9 ();
 sg13g2_fill_2 FILLER_20_44 ();
 sg13g2_decap_4 FILLER_20_56 ();
 sg13g2_fill_2 FILLER_20_60 ();
 sg13g2_fill_2 FILLER_20_96 ();
 sg13g2_fill_2 FILLER_20_119 ();
 sg13g2_fill_1 FILLER_20_134 ();
 sg13g2_fill_1 FILLER_20_143 ();
 sg13g2_fill_1 FILLER_20_152 ();
 sg13g2_fill_1 FILLER_20_157 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_178 ();
 sg13g2_decap_4 FILLER_20_185 ();
 sg13g2_fill_2 FILLER_20_189 ();
 sg13g2_fill_1 FILLER_20_195 ();
 sg13g2_fill_2 FILLER_20_276 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_294 ();
 sg13g2_fill_2 FILLER_20_309 ();
 sg13g2_fill_1 FILLER_20_311 ();
 sg13g2_decap_8 FILLER_20_320 ();
 sg13g2_fill_2 FILLER_20_336 ();
 sg13g2_fill_1 FILLER_20_342 ();
 sg13g2_fill_1 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_409 ();
 sg13g2_decap_8 FILLER_20_478 ();
 sg13g2_fill_1 FILLER_20_485 ();
 sg13g2_fill_2 FILLER_20_499 ();
 sg13g2_fill_1 FILLER_20_514 ();
 sg13g2_fill_1 FILLER_20_539 ();
 sg13g2_fill_2 FILLER_20_544 ();
 sg13g2_fill_2 FILLER_20_551 ();
 sg13g2_decap_4 FILLER_20_613 ();
 sg13g2_fill_1 FILLER_20_617 ();
 sg13g2_fill_2 FILLER_20_650 ();
 sg13g2_fill_1 FILLER_20_659 ();
 sg13g2_decap_8 FILLER_20_696 ();
 sg13g2_fill_1 FILLER_20_703 ();
 sg13g2_fill_2 FILLER_20_802 ();
 sg13g2_decap_8 FILLER_20_830 ();
 sg13g2_decap_8 FILLER_20_837 ();
 sg13g2_decap_8 FILLER_20_844 ();
 sg13g2_fill_2 FILLER_20_851 ();
 sg13g2_decap_8 FILLER_20_887 ();
 sg13g2_fill_1 FILLER_20_894 ();
 sg13g2_decap_8 FILLER_20_909 ();
 sg13g2_fill_1 FILLER_20_930 ();
 sg13g2_decap_4 FILLER_20_936 ();
 sg13g2_fill_1 FILLER_20_940 ();
 sg13g2_fill_2 FILLER_20_972 ();
 sg13g2_fill_2 FILLER_20_984 ();
 sg13g2_fill_2 FILLER_20_1012 ();
 sg13g2_fill_1 FILLER_20_1014 ();
 sg13g2_fill_2 FILLER_20_1024 ();
 sg13g2_fill_2 FILLER_20_1031 ();
 sg13g2_fill_2 FILLER_20_1037 ();
 sg13g2_fill_2 FILLER_20_1043 ();
 sg13g2_fill_2 FILLER_20_1050 ();
 sg13g2_fill_2 FILLER_20_1056 ();
 sg13g2_decap_4 FILLER_20_1062 ();
 sg13g2_fill_1 FILLER_20_1066 ();
 sg13g2_fill_2 FILLER_20_1072 ();
 sg13g2_fill_1 FILLER_20_1088 ();
 sg13g2_decap_4 FILLER_20_1172 ();
 sg13g2_fill_1 FILLER_20_1176 ();
 sg13g2_decap_8 FILLER_20_1181 ();
 sg13g2_decap_8 FILLER_20_1188 ();
 sg13g2_decap_8 FILLER_20_1195 ();
 sg13g2_decap_8 FILLER_20_1202 ();
 sg13g2_decap_8 FILLER_20_1209 ();
 sg13g2_decap_8 FILLER_20_1216 ();
 sg13g2_decap_8 FILLER_20_1223 ();
 sg13g2_decap_4 FILLER_20_1230 ();
 sg13g2_fill_2 FILLER_20_1234 ();
 sg13g2_decap_8 FILLER_20_1240 ();
 sg13g2_decap_8 FILLER_20_1247 ();
 sg13g2_decap_8 FILLER_20_1254 ();
 sg13g2_fill_1 FILLER_20_1261 ();
 sg13g2_fill_2 FILLER_20_1272 ();
 sg13g2_decap_4 FILLER_20_1313 ();
 sg13g2_fill_1 FILLER_20_1317 ();
 sg13g2_decap_4 FILLER_20_1322 ();
 sg13g2_fill_2 FILLER_20_1336 ();
 sg13g2_decap_4 FILLER_20_1348 ();
 sg13g2_fill_1 FILLER_20_1352 ();
 sg13g2_decap_8 FILLER_20_1410 ();
 sg13g2_fill_1 FILLER_20_1455 ();
 sg13g2_fill_1 FILLER_20_1459 ();
 sg13g2_fill_1 FILLER_20_1463 ();
 sg13g2_fill_2 FILLER_20_1484 ();
 sg13g2_fill_1 FILLER_20_1494 ();
 sg13g2_decap_4 FILLER_20_1555 ();
 sg13g2_fill_2 FILLER_20_1633 ();
 sg13g2_fill_1 FILLER_20_1716 ();
 sg13g2_decap_4 FILLER_20_1757 ();
 sg13g2_fill_1 FILLER_20_1761 ();
 sg13g2_fill_1 FILLER_20_1792 ();
 sg13g2_fill_2 FILLER_20_1797 ();
 sg13g2_decap_8 FILLER_20_1804 ();
 sg13g2_decap_8 FILLER_20_1811 ();
 sg13g2_decap_4 FILLER_20_1818 ();
 sg13g2_fill_2 FILLER_20_1822 ();
 sg13g2_fill_1 FILLER_20_1832 ();
 sg13g2_decap_8 FILLER_20_1837 ();
 sg13g2_decap_8 FILLER_20_1844 ();
 sg13g2_decap_4 FILLER_20_1851 ();
 sg13g2_fill_1 FILLER_20_1855 ();
 sg13g2_fill_2 FILLER_20_1860 ();
 sg13g2_fill_1 FILLER_20_1862 ();
 sg13g2_fill_2 FILLER_20_1867 ();
 sg13g2_fill_1 FILLER_20_1869 ();
 sg13g2_decap_8 FILLER_20_1874 ();
 sg13g2_decap_4 FILLER_20_1881 ();
 sg13g2_fill_1 FILLER_20_1885 ();
 sg13g2_fill_1 FILLER_20_1894 ();
 sg13g2_fill_2 FILLER_20_1923 ();
 sg13g2_decap_4 FILLER_20_1929 ();
 sg13g2_fill_1 FILLER_20_1933 ();
 sg13g2_decap_4 FILLER_20_1938 ();
 sg13g2_decap_8 FILLER_20_1951 ();
 sg13g2_decap_4 FILLER_20_1967 ();
 sg13g2_fill_1 FILLER_20_1971 ();
 sg13g2_fill_2 FILLER_20_2007 ();
 sg13g2_fill_1 FILLER_20_2021 ();
 sg13g2_fill_2 FILLER_20_2053 ();
 sg13g2_fill_1 FILLER_20_2055 ();
 sg13g2_fill_1 FILLER_20_2090 ();
 sg13g2_fill_2 FILLER_20_2094 ();
 sg13g2_fill_2 FILLER_20_2112 ();
 sg13g2_decap_8 FILLER_20_2140 ();
 sg13g2_decap_4 FILLER_20_2147 ();
 sg13g2_decap_4 FILLER_20_2159 ();
 sg13g2_decap_8 FILLER_20_2173 ();
 sg13g2_decap_8 FILLER_20_2180 ();
 sg13g2_decap_4 FILLER_20_2187 ();
 sg13g2_fill_1 FILLER_20_2191 ();
 sg13g2_decap_8 FILLER_20_2196 ();
 sg13g2_decap_8 FILLER_20_2203 ();
 sg13g2_fill_2 FILLER_20_2210 ();
 sg13g2_fill_1 FILLER_20_2212 ();
 sg13g2_decap_8 FILLER_20_2223 ();
 sg13g2_decap_4 FILLER_20_2266 ();
 sg13g2_fill_2 FILLER_20_2270 ();
 sg13g2_fill_2 FILLER_20_2316 ();
 sg13g2_fill_1 FILLER_20_2318 ();
 sg13g2_fill_1 FILLER_20_2324 ();
 sg13g2_decap_4 FILLER_20_2330 ();
 sg13g2_fill_1 FILLER_20_2334 ();
 sg13g2_fill_1 FILLER_20_2347 ();
 sg13g2_fill_2 FILLER_20_2354 ();
 sg13g2_decap_4 FILLER_20_2398 ();
 sg13g2_fill_2 FILLER_20_2402 ();
 sg13g2_fill_1 FILLER_20_2408 ();
 sg13g2_fill_1 FILLER_20_2419 ();
 sg13g2_fill_1 FILLER_20_2436 ();
 sg13g2_fill_1 FILLER_20_2469 ();
 sg13g2_fill_1 FILLER_20_2551 ();
 sg13g2_fill_1 FILLER_20_2563 ();
 sg13g2_fill_1 FILLER_20_2576 ();
 sg13g2_fill_2 FILLER_20_2615 ();
 sg13g2_fill_1 FILLER_20_2617 ();
 sg13g2_fill_2 FILLER_20_2623 ();
 sg13g2_fill_1 FILLER_20_2625 ();
 sg13g2_fill_2 FILLER_20_2636 ();
 sg13g2_fill_2 FILLER_20_2668 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_decap_8 FILLER_21_34 ();
 sg13g2_fill_2 FILLER_21_51 ();
 sg13g2_decap_4 FILLER_21_57 ();
 sg13g2_fill_1 FILLER_21_61 ();
 sg13g2_decap_4 FILLER_21_97 ();
 sg13g2_fill_2 FILLER_21_101 ();
 sg13g2_decap_8 FILLER_21_111 ();
 sg13g2_decap_8 FILLER_21_118 ();
 sg13g2_fill_1 FILLER_21_125 ();
 sg13g2_decap_8 FILLER_21_130 ();
 sg13g2_decap_8 FILLER_21_137 ();
 sg13g2_decap_8 FILLER_21_144 ();
 sg13g2_decap_4 FILLER_21_151 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_fill_2 FILLER_21_185 ();
 sg13g2_fill_1 FILLER_21_187 ();
 sg13g2_fill_1 FILLER_21_193 ();
 sg13g2_decap_4 FILLER_21_228 ();
 sg13g2_fill_1 FILLER_21_232 ();
 sg13g2_decap_4 FILLER_21_238 ();
 sg13g2_fill_2 FILLER_21_290 ();
 sg13g2_fill_1 FILLER_21_304 ();
 sg13g2_fill_1 FILLER_21_309 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_fill_2 FILLER_21_322 ();
 sg13g2_fill_1 FILLER_21_344 ();
 sg13g2_fill_2 FILLER_21_364 ();
 sg13g2_decap_4 FILLER_21_397 ();
 sg13g2_fill_1 FILLER_21_401 ();
 sg13g2_fill_2 FILLER_21_420 ();
 sg13g2_fill_1 FILLER_21_426 ();
 sg13g2_fill_2 FILLER_21_469 ();
 sg13g2_fill_1 FILLER_21_471 ();
 sg13g2_fill_2 FILLER_21_511 ();
 sg13g2_fill_1 FILLER_21_578 ();
 sg13g2_fill_2 FILLER_21_586 ();
 sg13g2_fill_2 FILLER_21_599 ();
 sg13g2_fill_1 FILLER_21_601 ();
 sg13g2_decap_8 FILLER_21_606 ();
 sg13g2_decap_4 FILLER_21_613 ();
 sg13g2_fill_2 FILLER_21_617 ();
 sg13g2_decap_8 FILLER_21_694 ();
 sg13g2_decap_8 FILLER_21_701 ();
 sg13g2_fill_1 FILLER_21_708 ();
 sg13g2_fill_1 FILLER_21_719 ();
 sg13g2_fill_2 FILLER_21_741 ();
 sg13g2_fill_1 FILLER_21_743 ();
 sg13g2_fill_2 FILLER_21_776 ();
 sg13g2_fill_2 FILLER_21_782 ();
 sg13g2_fill_1 FILLER_21_784 ();
 sg13g2_fill_2 FILLER_21_815 ();
 sg13g2_decap_4 FILLER_21_853 ();
 sg13g2_fill_1 FILLER_21_857 ();
 sg13g2_fill_2 FILLER_21_868 ();
 sg13g2_fill_1 FILLER_21_870 ();
 sg13g2_decap_8 FILLER_21_897 ();
 sg13g2_fill_2 FILLER_21_904 ();
 sg13g2_decap_8 FILLER_21_940 ();
 sg13g2_decap_4 FILLER_21_947 ();
 sg13g2_fill_1 FILLER_21_951 ();
 sg13g2_decap_4 FILLER_21_988 ();
 sg13g2_fill_1 FILLER_21_992 ();
 sg13g2_decap_8 FILLER_21_997 ();
 sg13g2_fill_2 FILLER_21_1004 ();
 sg13g2_fill_1 FILLER_21_1009 ();
 sg13g2_fill_1 FILLER_21_1044 ();
 sg13g2_decap_4 FILLER_21_1071 ();
 sg13g2_fill_1 FILLER_21_1075 ();
 sg13g2_fill_1 FILLER_21_1094 ();
 sg13g2_fill_1 FILLER_21_1103 ();
 sg13g2_fill_1 FILLER_21_1122 ();
 sg13g2_fill_1 FILLER_21_1129 ();
 sg13g2_fill_2 FILLER_21_1134 ();
 sg13g2_decap_4 FILLER_21_1203 ();
 sg13g2_fill_1 FILLER_21_1211 ();
 sg13g2_fill_2 FILLER_21_1217 ();
 sg13g2_fill_1 FILLER_21_1219 ();
 sg13g2_decap_8 FILLER_21_1228 ();
 sg13g2_decap_8 FILLER_21_1235 ();
 sg13g2_decap_8 FILLER_21_1242 ();
 sg13g2_fill_2 FILLER_21_1249 ();
 sg13g2_decap_4 FILLER_21_1255 ();
 sg13g2_fill_1 FILLER_21_1259 ();
 sg13g2_decap_8 FILLER_21_1270 ();
 sg13g2_decap_8 FILLER_21_1277 ();
 sg13g2_fill_2 FILLER_21_1284 ();
 sg13g2_decap_8 FILLER_21_1290 ();
 sg13g2_fill_2 FILLER_21_1297 ();
 sg13g2_decap_8 FILLER_21_1308 ();
 sg13g2_decap_8 FILLER_21_1315 ();
 sg13g2_decap_8 FILLER_21_1322 ();
 sg13g2_decap_4 FILLER_21_1329 ();
 sg13g2_fill_2 FILLER_21_1333 ();
 sg13g2_decap_8 FILLER_21_1395 ();
 sg13g2_decap_8 FILLER_21_1402 ();
 sg13g2_fill_2 FILLER_21_1409 ();
 sg13g2_fill_2 FILLER_21_1421 ();
 sg13g2_fill_2 FILLER_21_1428 ();
 sg13g2_fill_1 FILLER_21_1430 ();
 sg13g2_fill_1 FILLER_21_1441 ();
 sg13g2_fill_1 FILLER_21_1494 ();
 sg13g2_fill_2 FILLER_21_1509 ();
 sg13g2_fill_1 FILLER_21_1516 ();
 sg13g2_fill_1 FILLER_21_1556 ();
 sg13g2_fill_2 FILLER_21_1578 ();
 sg13g2_fill_1 FILLER_21_1580 ();
 sg13g2_fill_2 FILLER_21_1586 ();
 sg13g2_fill_1 FILLER_21_1630 ();
 sg13g2_fill_2 FILLER_21_1636 ();
 sg13g2_fill_2 FILLER_21_1643 ();
 sg13g2_fill_1 FILLER_21_1711 ();
 sg13g2_decap_4 FILLER_21_1717 ();
 sg13g2_fill_2 FILLER_21_1721 ();
 sg13g2_decap_8 FILLER_21_1727 ();
 sg13g2_decap_8 FILLER_21_1734 ();
 sg13g2_decap_8 FILLER_21_1741 ();
 sg13g2_decap_8 FILLER_21_1748 ();
 sg13g2_decap_8 FILLER_21_1755 ();
 sg13g2_decap_8 FILLER_21_1762 ();
 sg13g2_decap_4 FILLER_21_1769 ();
 sg13g2_fill_1 FILLER_21_1773 ();
 sg13g2_decap_8 FILLER_21_1778 ();
 sg13g2_fill_2 FILLER_21_1785 ();
 sg13g2_fill_1 FILLER_21_1787 ();
 sg13g2_fill_1 FILLER_21_1800 ();
 sg13g2_decap_4 FILLER_21_1805 ();
 sg13g2_fill_1 FILLER_21_1856 ();
 sg13g2_fill_2 FILLER_21_1871 ();
 sg13g2_fill_1 FILLER_21_1873 ();
 sg13g2_fill_1 FILLER_21_1902 ();
 sg13g2_fill_1 FILLER_21_1944 ();
 sg13g2_fill_1 FILLER_21_1954 ();
 sg13g2_decap_8 FILLER_21_1964 ();
 sg13g2_decap_4 FILLER_21_1971 ();
 sg13g2_fill_2 FILLER_21_1982 ();
 sg13g2_decap_8 FILLER_21_2056 ();
 sg13g2_fill_1 FILLER_21_2063 ();
 sg13g2_fill_2 FILLER_21_2074 ();
 sg13g2_fill_1 FILLER_21_2090 ();
 sg13g2_fill_2 FILLER_21_2104 ();
 sg13g2_fill_1 FILLER_21_2116 ();
 sg13g2_fill_2 FILLER_21_2125 ();
 sg13g2_decap_8 FILLER_21_2131 ();
 sg13g2_fill_2 FILLER_21_2138 ();
 sg13g2_fill_1 FILLER_21_2140 ();
 sg13g2_decap_8 FILLER_21_2177 ();
 sg13g2_fill_2 FILLER_21_2184 ();
 sg13g2_fill_2 FILLER_21_2252 ();
 sg13g2_fill_1 FILLER_21_2254 ();
 sg13g2_fill_1 FILLER_21_2281 ();
 sg13g2_fill_1 FILLER_21_2287 ();
 sg13g2_fill_1 FILLER_21_2294 ();
 sg13g2_decap_8 FILLER_21_2311 ();
 sg13g2_fill_1 FILLER_21_2318 ();
 sg13g2_fill_1 FILLER_21_2329 ();
 sg13g2_fill_1 FILLER_21_2340 ();
 sg13g2_fill_1 FILLER_21_2347 ();
 sg13g2_fill_1 FILLER_21_2353 ();
 sg13g2_fill_2 FILLER_21_2364 ();
 sg13g2_fill_1 FILLER_21_2370 ();
 sg13g2_fill_2 FILLER_21_2481 ();
 sg13g2_fill_2 FILLER_21_2515 ();
 sg13g2_fill_1 FILLER_21_2584 ();
 sg13g2_decap_8 FILLER_21_2663 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_9 ();
 sg13g2_decap_4 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_22 ();
 sg13g2_decap_8 FILLER_22_29 ();
 sg13g2_fill_2 FILLER_22_36 ();
 sg13g2_fill_1 FILLER_22_69 ();
 sg13g2_fill_2 FILLER_22_74 ();
 sg13g2_fill_1 FILLER_22_76 ();
 sg13g2_decap_4 FILLER_22_82 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_decap_4 FILLER_22_116 ();
 sg13g2_fill_2 FILLER_22_120 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_fill_1 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_152 ();
 sg13g2_decap_4 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_163 ();
 sg13g2_decap_4 FILLER_22_231 ();
 sg13g2_fill_1 FILLER_22_235 ();
 sg13g2_decap_4 FILLER_22_241 ();
 sg13g2_fill_1 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_276 ();
 sg13g2_fill_2 FILLER_22_283 ();
 sg13g2_fill_1 FILLER_22_285 ();
 sg13g2_fill_1 FILLER_22_294 ();
 sg13g2_fill_1 FILLER_22_303 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_fill_1 FILLER_22_351 ();
 sg13g2_fill_2 FILLER_22_356 ();
 sg13g2_fill_1 FILLER_22_364 ();
 sg13g2_fill_1 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_399 ();
 sg13g2_fill_1 FILLER_22_405 ();
 sg13g2_fill_1 FILLER_22_416 ();
 sg13g2_fill_1 FILLER_22_427 ();
 sg13g2_fill_2 FILLER_22_440 ();
 sg13g2_fill_1 FILLER_22_442 ();
 sg13g2_decap_4 FILLER_22_457 ();
 sg13g2_decap_4 FILLER_22_465 ();
 sg13g2_fill_1 FILLER_22_479 ();
 sg13g2_fill_2 FILLER_22_484 ();
 sg13g2_fill_2 FILLER_22_512 ();
 sg13g2_fill_2 FILLER_22_518 ();
 sg13g2_decap_4 FILLER_22_524 ();
 sg13g2_fill_1 FILLER_22_528 ();
 sg13g2_fill_1 FILLER_22_583 ();
 sg13g2_fill_2 FILLER_22_591 ();
 sg13g2_fill_2 FILLER_22_604 ();
 sg13g2_fill_1 FILLER_22_685 ();
 sg13g2_fill_2 FILLER_22_716 ();
 sg13g2_fill_2 FILLER_22_744 ();
 sg13g2_fill_1 FILLER_22_782 ();
 sg13g2_fill_1 FILLER_22_787 ();
 sg13g2_fill_1 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_820 ();
 sg13g2_decap_4 FILLER_22_827 ();
 sg13g2_fill_2 FILLER_22_831 ();
 sg13g2_decap_4 FILLER_22_837 ();
 sg13g2_fill_1 FILLER_22_841 ();
 sg13g2_decap_4 FILLER_22_889 ();
 sg13g2_fill_2 FILLER_22_893 ();
 sg13g2_fill_2 FILLER_22_905 ();
 sg13g2_fill_1 FILLER_22_907 ();
 sg13g2_decap_4 FILLER_22_918 ();
 sg13g2_fill_2 FILLER_22_922 ();
 sg13g2_decap_8 FILLER_22_945 ();
 sg13g2_decap_8 FILLER_22_952 ();
 sg13g2_decap_4 FILLER_22_959 ();
 sg13g2_fill_2 FILLER_22_994 ();
 sg13g2_fill_2 FILLER_22_1020 ();
 sg13g2_fill_1 FILLER_22_1022 ();
 sg13g2_fill_2 FILLER_22_1035 ();
 sg13g2_fill_2 FILLER_22_1042 ();
 sg13g2_fill_1 FILLER_22_1044 ();
 sg13g2_decap_4 FILLER_22_1085 ();
 sg13g2_fill_2 FILLER_22_1089 ();
 sg13g2_fill_1 FILLER_22_1108 ();
 sg13g2_fill_2 FILLER_22_1117 ();
 sg13g2_fill_2 FILLER_22_1165 ();
 sg13g2_fill_2 FILLER_22_1176 ();
 sg13g2_fill_1 FILLER_22_1212 ();
 sg13g2_fill_2 FILLER_22_1239 ();
 sg13g2_fill_2 FILLER_22_1267 ();
 sg13g2_fill_2 FILLER_22_1295 ();
 sg13g2_fill_1 FILLER_22_1297 ();
 sg13g2_fill_2 FILLER_22_1308 ();
 sg13g2_fill_1 FILLER_22_1310 ();
 sg13g2_fill_2 FILLER_22_1321 ();
 sg13g2_fill_1 FILLER_22_1323 ();
 sg13g2_fill_1 FILLER_22_1358 ();
 sg13g2_decap_4 FILLER_22_1369 ();
 sg13g2_decap_8 FILLER_22_1377 ();
 sg13g2_decap_4 FILLER_22_1384 ();
 sg13g2_fill_2 FILLER_22_1388 ();
 sg13g2_decap_8 FILLER_22_1400 ();
 sg13g2_fill_1 FILLER_22_1459 ();
 sg13g2_fill_2 FILLER_22_1473 ();
 sg13g2_fill_2 FILLER_22_1486 ();
 sg13g2_fill_1 FILLER_22_1517 ();
 sg13g2_decap_4 FILLER_22_1551 ();
 sg13g2_fill_2 FILLER_22_1555 ();
 sg13g2_decap_8 FILLER_22_1567 ();
 sg13g2_decap_4 FILLER_22_1574 ();
 sg13g2_fill_2 FILLER_22_1578 ();
 sg13g2_decap_8 FILLER_22_1611 ();
 sg13g2_decap_8 FILLER_22_1618 ();
 sg13g2_fill_1 FILLER_22_1625 ();
 sg13g2_decap_8 FILLER_22_1671 ();
 sg13g2_decap_8 FILLER_22_1678 ();
 sg13g2_decap_8 FILLER_22_1685 ();
 sg13g2_fill_2 FILLER_22_1692 ();
 sg13g2_fill_1 FILLER_22_1694 ();
 sg13g2_decap_8 FILLER_22_1699 ();
 sg13g2_decap_8 FILLER_22_1706 ();
 sg13g2_decap_4 FILLER_22_1713 ();
 sg13g2_fill_2 FILLER_22_1717 ();
 sg13g2_fill_1 FILLER_22_1733 ();
 sg13g2_decap_8 FILLER_22_1739 ();
 sg13g2_decap_4 FILLER_22_1746 ();
 sg13g2_decap_8 FILLER_22_1755 ();
 sg13g2_decap_8 FILLER_22_1762 ();
 sg13g2_decap_8 FILLER_22_1769 ();
 sg13g2_decap_8 FILLER_22_1776 ();
 sg13g2_fill_2 FILLER_22_1783 ();
 sg13g2_fill_1 FILLER_22_1785 ();
 sg13g2_fill_1 FILLER_22_1817 ();
 sg13g2_fill_2 FILLER_22_1827 ();
 sg13g2_fill_2 FILLER_22_1851 ();
 sg13g2_fill_2 FILLER_22_1878 ();
 sg13g2_decap_4 FILLER_22_1965 ();
 sg13g2_fill_2 FILLER_22_1978 ();
 sg13g2_fill_1 FILLER_22_1984 ();
 sg13g2_decap_4 FILLER_22_1993 ();
 sg13g2_fill_2 FILLER_22_1997 ();
 sg13g2_fill_1 FILLER_22_2017 ();
 sg13g2_decap_8 FILLER_22_2054 ();
 sg13g2_fill_1 FILLER_22_2098 ();
 sg13g2_fill_2 FILLER_22_2198 ();
 sg13g2_fill_1 FILLER_22_2200 ();
 sg13g2_fill_1 FILLER_22_2231 ();
 sg13g2_decap_8 FILLER_22_2257 ();
 sg13g2_decap_8 FILLER_22_2268 ();
 sg13g2_decap_8 FILLER_22_2275 ();
 sg13g2_fill_2 FILLER_22_2286 ();
 sg13g2_fill_2 FILLER_22_2294 ();
 sg13g2_fill_1 FILLER_22_2305 ();
 sg13g2_fill_2 FILLER_22_2366 ();
 sg13g2_fill_1 FILLER_22_2368 ();
 sg13g2_fill_1 FILLER_22_2373 ();
 sg13g2_decap_4 FILLER_22_2400 ();
 sg13g2_fill_1 FILLER_22_2424 ();
 sg13g2_fill_1 FILLER_22_2434 ();
 sg13g2_decap_8 FILLER_22_2479 ();
 sg13g2_decap_4 FILLER_22_2486 ();
 sg13g2_fill_1 FILLER_22_2490 ();
 sg13g2_fill_2 FILLER_22_2505 ();
 sg13g2_decap_8 FILLER_22_2515 ();
 sg13g2_decap_8 FILLER_22_2522 ();
 sg13g2_decap_8 FILLER_22_2529 ();
 sg13g2_fill_1 FILLER_22_2536 ();
 sg13g2_fill_1 FILLER_22_2577 ();
 sg13g2_fill_1 FILLER_22_2588 ();
 sg13g2_fill_1 FILLER_22_2623 ();
 sg13g2_fill_1 FILLER_22_2638 ();
 sg13g2_decap_8 FILLER_22_2657 ();
 sg13g2_decap_4 FILLER_22_2664 ();
 sg13g2_fill_2 FILLER_22_2668 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_fill_1 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_52 ();
 sg13g2_fill_1 FILLER_23_59 ();
 sg13g2_fill_2 FILLER_23_64 ();
 sg13g2_decap_8 FILLER_23_74 ();
 sg13g2_decap_4 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_85 ();
 sg13g2_fill_1 FILLER_23_89 ();
 sg13g2_fill_1 FILLER_23_94 ();
 sg13g2_fill_1 FILLER_23_100 ();
 sg13g2_fill_2 FILLER_23_105 ();
 sg13g2_fill_2 FILLER_23_111 ();
 sg13g2_fill_1 FILLER_23_113 ();
 sg13g2_decap_8 FILLER_23_174 ();
 sg13g2_decap_4 FILLER_23_181 ();
 sg13g2_fill_1 FILLER_23_185 ();
 sg13g2_decap_8 FILLER_23_191 ();
 sg13g2_fill_2 FILLER_23_198 ();
 sg13g2_fill_1 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_205 ();
 sg13g2_decap_4 FILLER_23_212 ();
 sg13g2_fill_2 FILLER_23_220 ();
 sg13g2_fill_1 FILLER_23_222 ();
 sg13g2_decap_4 FILLER_23_227 ();
 sg13g2_fill_2 FILLER_23_231 ();
 sg13g2_fill_2 FILLER_23_238 ();
 sg13g2_fill_1 FILLER_23_240 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_fill_2 FILLER_23_250 ();
 sg13g2_fill_1 FILLER_23_252 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_fill_2 FILLER_23_300 ();
 sg13g2_fill_2 FILLER_23_307 ();
 sg13g2_fill_2 FILLER_23_314 ();
 sg13g2_fill_1 FILLER_23_371 ();
 sg13g2_fill_2 FILLER_23_413 ();
 sg13g2_fill_1 FILLER_23_419 ();
 sg13g2_fill_2 FILLER_23_438 ();
 sg13g2_fill_1 FILLER_23_449 ();
 sg13g2_decap_8 FILLER_23_458 ();
 sg13g2_decap_4 FILLER_23_465 ();
 sg13g2_fill_2 FILLER_23_469 ();
 sg13g2_fill_1 FILLER_23_480 ();
 sg13g2_fill_1 FILLER_23_486 ();
 sg13g2_fill_1 FILLER_23_491 ();
 sg13g2_fill_2 FILLER_23_496 ();
 sg13g2_fill_2 FILLER_23_528 ();
 sg13g2_fill_2 FILLER_23_559 ();
 sg13g2_fill_1 FILLER_23_574 ();
 sg13g2_fill_2 FILLER_23_586 ();
 sg13g2_fill_1 FILLER_23_618 ();
 sg13g2_fill_1 FILLER_23_645 ();
 sg13g2_fill_2 FILLER_23_653 ();
 sg13g2_fill_2 FILLER_23_667 ();
 sg13g2_decap_8 FILLER_23_685 ();
 sg13g2_decap_4 FILLER_23_692 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_4 FILLER_23_707 ();
 sg13g2_fill_1 FILLER_23_725 ();
 sg13g2_decap_4 FILLER_23_736 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_fill_2 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_828 ();
 sg13g2_decap_4 FILLER_23_835 ();
 sg13g2_decap_4 FILLER_23_853 ();
 sg13g2_fill_1 FILLER_23_857 ();
 sg13g2_fill_1 FILLER_23_867 ();
 sg13g2_fill_2 FILLER_23_899 ();
 sg13g2_decap_8 FILLER_23_974 ();
 sg13g2_fill_2 FILLER_23_981 ();
 sg13g2_fill_2 FILLER_23_1022 ();
 sg13g2_fill_1 FILLER_23_1029 ();
 sg13g2_fill_1 FILLER_23_1034 ();
 sg13g2_fill_2 FILLER_23_1040 ();
 sg13g2_fill_1 FILLER_23_1046 ();
 sg13g2_fill_1 FILLER_23_1051 ();
 sg13g2_fill_2 FILLER_23_1078 ();
 sg13g2_fill_1 FILLER_23_1080 ();
 sg13g2_decap_4 FILLER_23_1145 ();
 sg13g2_fill_1 FILLER_23_1149 ();
 sg13g2_decap_8 FILLER_23_1158 ();
 sg13g2_fill_1 FILLER_23_1165 ();
 sg13g2_decap_8 FILLER_23_1223 ();
 sg13g2_decap_4 FILLER_23_1230 ();
 sg13g2_fill_2 FILLER_23_1234 ();
 sg13g2_fill_1 FILLER_23_1289 ();
 sg13g2_fill_2 FILLER_23_1311 ();
 sg13g2_decap_8 FILLER_23_1343 ();
 sg13g2_decap_8 FILLER_23_1354 ();
 sg13g2_decap_8 FILLER_23_1361 ();
 sg13g2_decap_8 FILLER_23_1368 ();
 sg13g2_decap_8 FILLER_23_1375 ();
 sg13g2_fill_1 FILLER_23_1382 ();
 sg13g2_fill_2 FILLER_23_1386 ();
 sg13g2_decap_4 FILLER_23_1414 ();
 sg13g2_fill_1 FILLER_23_1444 ();
 sg13g2_fill_2 FILLER_23_1448 ();
 sg13g2_fill_1 FILLER_23_1459 ();
 sg13g2_fill_1 FILLER_23_1477 ();
 sg13g2_fill_1 FILLER_23_1492 ();
 sg13g2_fill_2 FILLER_23_1513 ();
 sg13g2_fill_2 FILLER_23_1520 ();
 sg13g2_fill_2 FILLER_23_1529 ();
 sg13g2_decap_8 FILLER_23_1555 ();
 sg13g2_decap_8 FILLER_23_1562 ();
 sg13g2_fill_1 FILLER_23_1569 ();
 sg13g2_decap_4 FILLER_23_1574 ();
 sg13g2_fill_2 FILLER_23_1578 ();
 sg13g2_decap_4 FILLER_23_1621 ();
 sg13g2_fill_1 FILLER_23_1629 ();
 sg13g2_fill_2 FILLER_23_1638 ();
 sg13g2_fill_1 FILLER_23_1640 ();
 sg13g2_fill_2 FILLER_23_1655 ();
 sg13g2_fill_1 FILLER_23_1657 ();
 sg13g2_fill_1 FILLER_23_1662 ();
 sg13g2_fill_2 FILLER_23_1689 ();
 sg13g2_fill_1 FILLER_23_1691 ();
 sg13g2_decap_8 FILLER_23_1697 ();
 sg13g2_decap_8 FILLER_23_1704 ();
 sg13g2_fill_1 FILLER_23_1722 ();
 sg13g2_decap_4 FILLER_23_1736 ();
 sg13g2_fill_2 FILLER_23_1740 ();
 sg13g2_fill_2 FILLER_23_1772 ();
 sg13g2_fill_1 FILLER_23_1774 ();
 sg13g2_fill_1 FILLER_23_1837 ();
 sg13g2_fill_2 FILLER_23_1867 ();
 sg13g2_fill_1 FILLER_23_1884 ();
 sg13g2_fill_1 FILLER_23_1896 ();
 sg13g2_fill_1 FILLER_23_1901 ();
 sg13g2_fill_1 FILLER_23_1927 ();
 sg13g2_fill_2 FILLER_23_1931 ();
 sg13g2_fill_1 FILLER_23_1943 ();
 sg13g2_fill_1 FILLER_23_1966 ();
 sg13g2_decap_8 FILLER_23_1972 ();
 sg13g2_decap_4 FILLER_23_1991 ();
 sg13g2_fill_1 FILLER_23_1995 ();
 sg13g2_fill_2 FILLER_23_2039 ();
 sg13g2_fill_1 FILLER_23_2041 ();
 sg13g2_fill_1 FILLER_23_2068 ();
 sg13g2_fill_1 FILLER_23_2079 ();
 sg13g2_decap_4 FILLER_23_2106 ();
 sg13g2_fill_2 FILLER_23_2114 ();
 sg13g2_fill_2 FILLER_23_2190 ();
 sg13g2_fill_1 FILLER_23_2192 ();
 sg13g2_decap_8 FILLER_23_2197 ();
 sg13g2_decap_8 FILLER_23_2204 ();
 sg13g2_decap_4 FILLER_23_2211 ();
 sg13g2_fill_2 FILLER_23_2225 ();
 sg13g2_decap_4 FILLER_23_2251 ();
 sg13g2_fill_1 FILLER_23_2255 ();
 sg13g2_decap_8 FILLER_23_2260 ();
 sg13g2_fill_1 FILLER_23_2267 ();
 sg13g2_decap_4 FILLER_23_2273 ();
 sg13g2_fill_2 FILLER_23_2277 ();
 sg13g2_decap_4 FILLER_23_2283 ();
 sg13g2_fill_1 FILLER_23_2287 ();
 sg13g2_fill_2 FILLER_23_2297 ();
 sg13g2_fill_2 FILLER_23_2303 ();
 sg13g2_fill_1 FILLER_23_2340 ();
 sg13g2_decap_8 FILLER_23_2356 ();
 sg13g2_decap_4 FILLER_23_2363 ();
 sg13g2_fill_2 FILLER_23_2367 ();
 sg13g2_fill_2 FILLER_23_2379 ();
 sg13g2_fill_1 FILLER_23_2381 ();
 sg13g2_fill_2 FILLER_23_2388 ();
 sg13g2_fill_1 FILLER_23_2395 ();
 sg13g2_decap_8 FILLER_23_2402 ();
 sg13g2_decap_8 FILLER_23_2409 ();
 sg13g2_fill_2 FILLER_23_2431 ();
 sg13g2_decap_4 FILLER_23_2536 ();
 sg13g2_fill_2 FILLER_23_2551 ();
 sg13g2_fill_1 FILLER_23_2553 ();
 sg13g2_fill_2 FILLER_23_2558 ();
 sg13g2_decap_4 FILLER_23_2570 ();
 sg13g2_fill_1 FILLER_23_2574 ();
 sg13g2_fill_2 FILLER_23_2581 ();
 sg13g2_fill_2 FILLER_23_2602 ();
 sg13g2_fill_1 FILLER_23_2604 ();
 sg13g2_decap_8 FILLER_23_2610 ();
 sg13g2_decap_8 FILLER_23_2617 ();
 sg13g2_decap_8 FILLER_23_2624 ();
 sg13g2_decap_8 FILLER_23_2631 ();
 sg13g2_decap_8 FILLER_23_2638 ();
 sg13g2_decap_8 FILLER_23_2645 ();
 sg13g2_decap_8 FILLER_23_2652 ();
 sg13g2_decap_8 FILLER_23_2659 ();
 sg13g2_decap_4 FILLER_23_2666 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_2 ();
 sg13g2_fill_2 FILLER_24_33 ();
 sg13g2_fill_1 FILLER_24_35 ();
 sg13g2_decap_4 FILLER_24_41 ();
 sg13g2_fill_1 FILLER_24_45 ();
 sg13g2_fill_1 FILLER_24_51 ();
 sg13g2_decap_4 FILLER_24_134 ();
 sg13g2_fill_1 FILLER_24_138 ();
 sg13g2_fill_1 FILLER_24_169 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_210 ();
 sg13g2_fill_1 FILLER_24_212 ();
 sg13g2_decap_4 FILLER_24_217 ();
 sg13g2_fill_2 FILLER_24_221 ();
 sg13g2_decap_4 FILLER_24_227 ();
 sg13g2_fill_1 FILLER_24_236 ();
 sg13g2_fill_1 FILLER_24_246 ();
 sg13g2_fill_2 FILLER_24_252 ();
 sg13g2_fill_1 FILLER_24_254 ();
 sg13g2_fill_1 FILLER_24_260 ();
 sg13g2_fill_2 FILLER_24_275 ();
 sg13g2_fill_2 FILLER_24_285 ();
 sg13g2_fill_2 FILLER_24_354 ();
 sg13g2_fill_1 FILLER_24_361 ();
 sg13g2_fill_1 FILLER_24_366 ();
 sg13g2_fill_2 FILLER_24_371 ();
 sg13g2_fill_1 FILLER_24_396 ();
 sg13g2_fill_1 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_fill_2 FILLER_24_465 ();
 sg13g2_decap_4 FILLER_24_471 ();
 sg13g2_fill_2 FILLER_24_475 ();
 sg13g2_decap_8 FILLER_24_487 ();
 sg13g2_decap_4 FILLER_24_494 ();
 sg13g2_fill_2 FILLER_24_498 ();
 sg13g2_fill_2 FILLER_24_509 ();
 sg13g2_decap_8 FILLER_24_514 ();
 sg13g2_decap_8 FILLER_24_521 ();
 sg13g2_decap_8 FILLER_24_528 ();
 sg13g2_fill_2 FILLER_24_535 ();
 sg13g2_fill_1 FILLER_24_537 ();
 sg13g2_fill_1 FILLER_24_541 ();
 sg13g2_fill_2 FILLER_24_569 ();
 sg13g2_fill_1 FILLER_24_571 ();
 sg13g2_fill_2 FILLER_24_611 ();
 sg13g2_fill_2 FILLER_24_626 ();
 sg13g2_fill_2 FILLER_24_632 ();
 sg13g2_fill_1 FILLER_24_663 ();
 sg13g2_fill_1 FILLER_24_684 ();
 sg13g2_decap_8 FILLER_24_715 ();
 sg13g2_fill_2 FILLER_24_732 ();
 sg13g2_fill_1 FILLER_24_734 ();
 sg13g2_decap_8 FILLER_24_772 ();
 sg13g2_fill_1 FILLER_24_779 ();
 sg13g2_decap_8 FILLER_24_806 ();
 sg13g2_fill_2 FILLER_24_813 ();
 sg13g2_decap_8 FILLER_24_835 ();
 sg13g2_decap_8 FILLER_24_842 ();
 sg13g2_decap_8 FILLER_24_849 ();
 sg13g2_decap_8 FILLER_24_856 ();
 sg13g2_decap_8 FILLER_24_863 ();
 sg13g2_decap_4 FILLER_24_870 ();
 sg13g2_decap_8 FILLER_24_884 ();
 sg13g2_decap_8 FILLER_24_891 ();
 sg13g2_fill_1 FILLER_24_898 ();
 sg13g2_fill_1 FILLER_24_939 ();
 sg13g2_fill_2 FILLER_24_1004 ();
 sg13g2_fill_1 FILLER_24_1012 ();
 sg13g2_fill_1 FILLER_24_1016 ();
 sg13g2_fill_2 FILLER_24_1068 ();
 sg13g2_fill_1 FILLER_24_1070 ();
 sg13g2_fill_2 FILLER_24_1092 ();
 sg13g2_fill_2 FILLER_24_1119 ();
 sg13g2_fill_1 FILLER_24_1121 ();
 sg13g2_fill_2 FILLER_24_1148 ();
 sg13g2_fill_1 FILLER_24_1150 ();
 sg13g2_fill_1 FILLER_24_1172 ();
 sg13g2_fill_1 FILLER_24_1178 ();
 sg13g2_fill_1 FILLER_24_1188 ();
 sg13g2_fill_1 FILLER_24_1197 ();
 sg13g2_fill_2 FILLER_24_1215 ();
 sg13g2_decap_8 FILLER_24_1230 ();
 sg13g2_fill_2 FILLER_24_1242 ();
 sg13g2_fill_1 FILLER_24_1244 ();
 sg13g2_fill_1 FILLER_24_1250 ();
 sg13g2_fill_1 FILLER_24_1256 ();
 sg13g2_fill_2 FILLER_24_1261 ();
 sg13g2_decap_4 FILLER_24_1289 ();
 sg13g2_fill_1 FILLER_24_1293 ();
 sg13g2_decap_8 FILLER_24_1307 ();
 sg13g2_fill_2 FILLER_24_1314 ();
 sg13g2_decap_8 FILLER_24_1330 ();
 sg13g2_decap_8 FILLER_24_1337 ();
 sg13g2_decap_8 FILLER_24_1362 ();
 sg13g2_fill_2 FILLER_24_1369 ();
 sg13g2_fill_2 FILLER_24_1407 ();
 sg13g2_decap_4 FILLER_24_1422 ();
 sg13g2_decap_8 FILLER_24_1442 ();
 sg13g2_decap_8 FILLER_24_1449 ();
 sg13g2_decap_4 FILLER_24_1456 ();
 sg13g2_decap_4 FILLER_24_1470 ();
 sg13g2_decap_4 FILLER_24_1492 ();
 sg13g2_fill_2 FILLER_24_1505 ();
 sg13g2_decap_8 FILLER_24_1551 ();
 sg13g2_decap_8 FILLER_24_1558 ();
 sg13g2_fill_2 FILLER_24_1565 ();
 sg13g2_decap_4 FILLER_24_1572 ();
 sg13g2_fill_1 FILLER_24_1576 ();
 sg13g2_fill_2 FILLER_24_1587 ();
 sg13g2_decap_4 FILLER_24_1599 ();
 sg13g2_fill_1 FILLER_24_1603 ();
 sg13g2_decap_8 FILLER_24_1613 ();
 sg13g2_fill_1 FILLER_24_1620 ();
 sg13g2_fill_2 FILLER_24_1631 ();
 sg13g2_decap_8 FILLER_24_1638 ();
 sg13g2_decap_8 FILLER_24_1645 ();
 sg13g2_fill_1 FILLER_24_1652 ();
 sg13g2_decap_4 FILLER_24_1666 ();
 sg13g2_decap_4 FILLER_24_1674 ();
 sg13g2_fill_2 FILLER_24_1678 ();
 sg13g2_decap_8 FILLER_24_1697 ();
 sg13g2_fill_1 FILLER_24_1704 ();
 sg13g2_fill_2 FILLER_24_1721 ();
 sg13g2_decap_8 FILLER_24_1760 ();
 sg13g2_fill_1 FILLER_24_1767 ();
 sg13g2_decap_4 FILLER_24_1772 ();
 sg13g2_fill_1 FILLER_24_1789 ();
 sg13g2_fill_1 FILLER_24_1811 ();
 sg13g2_fill_2 FILLER_24_1817 ();
 sg13g2_fill_1 FILLER_24_1819 ();
 sg13g2_fill_2 FILLER_24_1826 ();
 sg13g2_fill_2 FILLER_24_1873 ();
 sg13g2_fill_1 FILLER_24_1901 ();
 sg13g2_fill_1 FILLER_24_1907 ();
 sg13g2_fill_1 FILLER_24_1922 ();
 sg13g2_fill_2 FILLER_24_1937 ();
 sg13g2_fill_1 FILLER_24_1963 ();
 sg13g2_decap_8 FILLER_24_1971 ();
 sg13g2_fill_2 FILLER_24_1978 ();
 sg13g2_fill_1 FILLER_24_2040 ();
 sg13g2_fill_2 FILLER_24_2062 ();
 sg13g2_fill_1 FILLER_24_2074 ();
 sg13g2_fill_1 FILLER_24_2101 ();
 sg13g2_fill_1 FILLER_24_2128 ();
 sg13g2_fill_2 FILLER_24_2164 ();
 sg13g2_decap_8 FILLER_24_2196 ();
 sg13g2_decap_8 FILLER_24_2203 ();
 sg13g2_decap_8 FILLER_24_2210 ();
 sg13g2_decap_4 FILLER_24_2217 ();
 sg13g2_fill_2 FILLER_24_2221 ();
 sg13g2_fill_2 FILLER_24_2233 ();
 sg13g2_fill_2 FILLER_24_2300 ();
 sg13g2_fill_1 FILLER_24_2302 ();
 sg13g2_decap_8 FILLER_24_2317 ();
 sg13g2_fill_1 FILLER_24_2324 ();
 sg13g2_decap_4 FILLER_24_2330 ();
 sg13g2_fill_2 FILLER_24_2334 ();
 sg13g2_decap_8 FILLER_24_2352 ();
 sg13g2_decap_8 FILLER_24_2359 ();
 sg13g2_decap_4 FILLER_24_2366 ();
 sg13g2_fill_1 FILLER_24_2370 ();
 sg13g2_decap_4 FILLER_24_2375 ();
 sg13g2_fill_2 FILLER_24_2379 ();
 sg13g2_decap_8 FILLER_24_2385 ();
 sg13g2_decap_8 FILLER_24_2392 ();
 sg13g2_decap_4 FILLER_24_2399 ();
 sg13g2_decap_4 FILLER_24_2429 ();
 sg13g2_fill_1 FILLER_24_2433 ();
 sg13g2_decap_4 FILLER_24_2438 ();
 sg13g2_fill_1 FILLER_24_2442 ();
 sg13g2_fill_2 FILLER_24_2451 ();
 sg13g2_fill_1 FILLER_24_2453 ();
 sg13g2_decap_4 FILLER_24_2463 ();
 sg13g2_fill_1 FILLER_24_2467 ();
 sg13g2_decap_8 FILLER_24_2477 ();
 sg13g2_fill_2 FILLER_24_2484 ();
 sg13g2_decap_8 FILLER_24_2490 ();
 sg13g2_decap_8 FILLER_24_2497 ();
 sg13g2_decap_8 FILLER_24_2504 ();
 sg13g2_decap_8 FILLER_24_2511 ();
 sg13g2_fill_1 FILLER_24_2518 ();
 sg13g2_decap_8 FILLER_24_2523 ();
 sg13g2_decap_4 FILLER_24_2530 ();
 sg13g2_fill_1 FILLER_24_2534 ();
 sg13g2_decap_8 FILLER_24_2544 ();
 sg13g2_decap_8 FILLER_24_2551 ();
 sg13g2_decap_8 FILLER_24_2573 ();
 sg13g2_decap_8 FILLER_24_2580 ();
 sg13g2_decap_4 FILLER_24_2587 ();
 sg13g2_fill_2 FILLER_24_2591 ();
 sg13g2_decap_4 FILLER_24_2597 ();
 sg13g2_decap_8 FILLER_24_2618 ();
 sg13g2_decap_8 FILLER_24_2625 ();
 sg13g2_fill_2 FILLER_24_2668 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_5 ();
 sg13g2_fill_1 FILLER_25_32 ();
 sg13g2_decap_4 FILLER_25_37 ();
 sg13g2_fill_2 FILLER_25_41 ();
 sg13g2_fill_2 FILLER_25_73 ();
 sg13g2_fill_1 FILLER_25_75 ();
 sg13g2_fill_1 FILLER_25_101 ();
 sg13g2_decap_4 FILLER_25_121 ();
 sg13g2_decap_4 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_163 ();
 sg13g2_fill_1 FILLER_25_194 ();
 sg13g2_fill_1 FILLER_25_199 ();
 sg13g2_fill_2 FILLER_25_230 ();
 sg13g2_fill_1 FILLER_25_232 ();
 sg13g2_fill_2 FILLER_25_282 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_fill_1 FILLER_25_355 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_fill_1 FILLER_25_409 ();
 sg13g2_fill_2 FILLER_25_413 ();
 sg13g2_fill_1 FILLER_25_415 ();
 sg13g2_decap_8 FILLER_25_490 ();
 sg13g2_decap_8 FILLER_25_497 ();
 sg13g2_fill_2 FILLER_25_504 ();
 sg13g2_fill_1 FILLER_25_608 ();
 sg13g2_fill_1 FILLER_25_619 ();
 sg13g2_decap_8 FILLER_25_688 ();
 sg13g2_fill_1 FILLER_25_695 ();
 sg13g2_fill_2 FILLER_25_743 ();
 sg13g2_fill_2 FILLER_25_807 ();
 sg13g2_fill_1 FILLER_25_809 ();
 sg13g2_decap_4 FILLER_25_887 ();
 sg13g2_fill_2 FILLER_25_891 ();
 sg13g2_fill_1 FILLER_25_933 ();
 sg13g2_fill_1 FILLER_25_938 ();
 sg13g2_decap_8 FILLER_25_943 ();
 sg13g2_decap_8 FILLER_25_950 ();
 sg13g2_fill_1 FILLER_25_1065 ();
 sg13g2_fill_2 FILLER_25_1097 ();
 sg13g2_decap_4 FILLER_25_1130 ();
 sg13g2_fill_2 FILLER_25_1176 ();
 sg13g2_fill_2 FILLER_25_1182 ();
 sg13g2_fill_2 FILLER_25_1193 ();
 sg13g2_fill_1 FILLER_25_1195 ();
 sg13g2_fill_2 FILLER_25_1235 ();
 sg13g2_decap_4 FILLER_25_1267 ();
 sg13g2_decap_8 FILLER_25_1279 ();
 sg13g2_fill_2 FILLER_25_1322 ();
 sg13g2_fill_1 FILLER_25_1324 ();
 sg13g2_fill_2 FILLER_25_1329 ();
 sg13g2_fill_1 FILLER_25_1357 ();
 sg13g2_fill_1 FILLER_25_1384 ();
 sg13g2_fill_2 FILLER_25_1390 ();
 sg13g2_decap_8 FILLER_25_1430 ();
 sg13g2_decap_8 FILLER_25_1437 ();
 sg13g2_decap_8 FILLER_25_1444 ();
 sg13g2_decap_8 FILLER_25_1451 ();
 sg13g2_decap_8 FILLER_25_1458 ();
 sg13g2_decap_8 FILLER_25_1465 ();
 sg13g2_fill_2 FILLER_25_1472 ();
 sg13g2_fill_2 FILLER_25_1478 ();
 sg13g2_fill_1 FILLER_25_1480 ();
 sg13g2_fill_2 FILLER_25_1510 ();
 sg13g2_fill_2 FILLER_25_1537 ();
 sg13g2_decap_8 FILLER_25_1557 ();
 sg13g2_decap_8 FILLER_25_1564 ();
 sg13g2_fill_1 FILLER_25_1571 ();
 sg13g2_fill_2 FILLER_25_1577 ();
 sg13g2_fill_1 FILLER_25_1579 ();
 sg13g2_fill_1 FILLER_25_1597 ();
 sg13g2_decap_8 FILLER_25_1606 ();
 sg13g2_fill_2 FILLER_25_1613 ();
 sg13g2_fill_1 FILLER_25_1634 ();
 sg13g2_decap_4 FILLER_25_1639 ();
 sg13g2_fill_1 FILLER_25_1643 ();
 sg13g2_decap_8 FILLER_25_1657 ();
 sg13g2_decap_8 FILLER_25_1664 ();
 sg13g2_fill_1 FILLER_25_1705 ();
 sg13g2_decap_4 FILLER_25_1710 ();
 sg13g2_decap_4 FILLER_25_1717 ();
 sg13g2_fill_1 FILLER_25_1721 ();
 sg13g2_decap_4 FILLER_25_1748 ();
 sg13g2_decap_8 FILLER_25_1756 ();
 sg13g2_decap_4 FILLER_25_1763 ();
 sg13g2_fill_1 FILLER_25_1767 ();
 sg13g2_decap_8 FILLER_25_1773 ();
 sg13g2_fill_2 FILLER_25_1780 ();
 sg13g2_fill_2 FILLER_25_1832 ();
 sg13g2_fill_1 FILLER_25_1844 ();
 sg13g2_fill_2 FILLER_25_1851 ();
 sg13g2_fill_1 FILLER_25_1853 ();
 sg13g2_fill_2 FILLER_25_1865 ();
 sg13g2_fill_2 FILLER_25_1871 ();
 sg13g2_fill_2 FILLER_25_1887 ();
 sg13g2_fill_1 FILLER_25_1944 ();
 sg13g2_fill_2 FILLER_25_1960 ();
 sg13g2_fill_1 FILLER_25_1962 ();
 sg13g2_decap_8 FILLER_25_1968 ();
 sg13g2_decap_4 FILLER_25_1975 ();
 sg13g2_fill_2 FILLER_25_2015 ();
 sg13g2_fill_1 FILLER_25_2017 ();
 sg13g2_fill_2 FILLER_25_2044 ();
 sg13g2_fill_1 FILLER_25_2050 ();
 sg13g2_fill_1 FILLER_25_2055 ();
 sg13g2_fill_2 FILLER_25_2096 ();
 sg13g2_fill_1 FILLER_25_2126 ();
 sg13g2_decap_4 FILLER_25_2166 ();
 sg13g2_decap_8 FILLER_25_2196 ();
 sg13g2_decap_8 FILLER_25_2203 ();
 sg13g2_fill_2 FILLER_25_2210 ();
 sg13g2_fill_1 FILLER_25_2212 ();
 sg13g2_decap_4 FILLER_25_2270 ();
 sg13g2_fill_1 FILLER_25_2316 ();
 sg13g2_fill_2 FILLER_25_2357 ();
 sg13g2_fill_1 FILLER_25_2359 ();
 sg13g2_fill_1 FILLER_25_2416 ();
 sg13g2_fill_1 FILLER_25_2444 ();
 sg13g2_decap_8 FILLER_25_2494 ();
 sg13g2_decap_8 FILLER_25_2501 ();
 sg13g2_decap_8 FILLER_25_2508 ();
 sg13g2_fill_1 FILLER_25_2557 ();
 sg13g2_fill_2 FILLER_25_2584 ();
 sg13g2_fill_1 FILLER_25_2586 ();
 sg13g2_fill_1 FILLER_25_2637 ();
 sg13g2_fill_2 FILLER_25_2668 ();
 sg13g2_fill_1 FILLER_26_38 ();
 sg13g2_fill_1 FILLER_26_82 ();
 sg13g2_fill_1 FILLER_26_91 ();
 sg13g2_fill_1 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_139 ();
 sg13g2_fill_1 FILLER_26_148 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_decap_4 FILLER_26_160 ();
 sg13g2_fill_2 FILLER_26_164 ();
 sg13g2_fill_1 FILLER_26_171 ();
 sg13g2_fill_1 FILLER_26_176 ();
 sg13g2_decap_4 FILLER_26_203 ();
 sg13g2_fill_2 FILLER_26_207 ();
 sg13g2_fill_1 FILLER_26_243 ();
 sg13g2_fill_2 FILLER_26_248 ();
 sg13g2_decap_8 FILLER_26_254 ();
 sg13g2_fill_1 FILLER_26_261 ();
 sg13g2_fill_2 FILLER_26_292 ();
 sg13g2_fill_1 FILLER_26_325 ();
 sg13g2_fill_2 FILLER_26_338 ();
 sg13g2_fill_2 FILLER_26_349 ();
 sg13g2_fill_1 FILLER_26_364 ();
 sg13g2_fill_2 FILLER_26_374 ();
 sg13g2_fill_1 FILLER_26_384 ();
 sg13g2_fill_1 FILLER_26_406 ();
 sg13g2_fill_2 FILLER_26_417 ();
 sg13g2_decap_4 FILLER_26_456 ();
 sg13g2_fill_2 FILLER_26_460 ();
 sg13g2_fill_2 FILLER_26_467 ();
 sg13g2_decap_8 FILLER_26_495 ();
 sg13g2_decap_8 FILLER_26_502 ();
 sg13g2_decap_4 FILLER_26_509 ();
 sg13g2_fill_1 FILLER_26_513 ();
 sg13g2_decap_8 FILLER_26_518 ();
 sg13g2_fill_1 FILLER_26_525 ();
 sg13g2_fill_1 FILLER_26_566 ();
 sg13g2_fill_2 FILLER_26_603 ();
 sg13g2_fill_2 FILLER_26_626 ();
 sg13g2_fill_2 FILLER_26_653 ();
 sg13g2_fill_2 FILLER_26_715 ();
 sg13g2_fill_1 FILLER_26_717 ();
 sg13g2_decap_8 FILLER_26_728 ();
 sg13g2_fill_2 FILLER_26_735 ();
 sg13g2_fill_2 FILLER_26_747 ();
 sg13g2_fill_1 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_754 ();
 sg13g2_decap_8 FILLER_26_761 ();
 sg13g2_decap_8 FILLER_26_768 ();
 sg13g2_decap_8 FILLER_26_775 ();
 sg13g2_decap_4 FILLER_26_827 ();
 sg13g2_decap_4 FILLER_26_841 ();
 sg13g2_decap_8 FILLER_26_875 ();
 sg13g2_fill_1 FILLER_26_882 ();
 sg13g2_decap_8 FILLER_26_909 ();
 sg13g2_decap_8 FILLER_26_916 ();
 sg13g2_fill_1 FILLER_26_923 ();
 sg13g2_fill_2 FILLER_26_934 ();
 sg13g2_fill_1 FILLER_26_936 ();
 sg13g2_decap_8 FILLER_26_950 ();
 sg13g2_fill_2 FILLER_26_957 ();
 sg13g2_fill_2 FILLER_26_967 ();
 sg13g2_fill_1 FILLER_26_969 ();
 sg13g2_fill_2 FILLER_26_992 ();
 sg13g2_fill_2 FILLER_26_998 ();
 sg13g2_fill_1 FILLER_26_1016 ();
 sg13g2_fill_2 FILLER_26_1022 ();
 sg13g2_fill_1 FILLER_26_1054 ();
 sg13g2_decap_4 FILLER_26_1105 ();
 sg13g2_fill_2 FILLER_26_1126 ();
 sg13g2_fill_2 FILLER_26_1142 ();
 sg13g2_fill_2 FILLER_26_1179 ();
 sg13g2_fill_1 FILLER_26_1181 ();
 sg13g2_fill_2 FILLER_26_1187 ();
 sg13g2_fill_1 FILLER_26_1189 ();
 sg13g2_fill_1 FILLER_26_1216 ();
 sg13g2_fill_1 FILLER_26_1238 ();
 sg13g2_fill_2 FILLER_26_1244 ();
 sg13g2_decap_4 FILLER_26_1251 ();
 sg13g2_decap_8 FILLER_26_1259 ();
 sg13g2_fill_2 FILLER_26_1266 ();
 sg13g2_decap_4 FILLER_26_1330 ();
 sg13g2_fill_2 FILLER_26_1334 ();
 sg13g2_decap_4 FILLER_26_1362 ();
 sg13g2_fill_1 FILLER_26_1366 ();
 sg13g2_fill_2 FILLER_26_1376 ();
 sg13g2_fill_1 FILLER_26_1378 ();
 sg13g2_decap_8 FILLER_26_1383 ();
 sg13g2_decap_8 FILLER_26_1390 ();
 sg13g2_decap_8 FILLER_26_1401 ();
 sg13g2_decap_8 FILLER_26_1408 ();
 sg13g2_decap_8 FILLER_26_1415 ();
 sg13g2_decap_4 FILLER_26_1427 ();
 sg13g2_decap_8 FILLER_26_1457 ();
 sg13g2_fill_1 FILLER_26_1464 ();
 sg13g2_fill_2 FILLER_26_1505 ();
 sg13g2_fill_1 FILLER_26_1519 ();
 sg13g2_fill_1 FILLER_26_1555 ();
 sg13g2_decap_4 FILLER_26_1601 ();
 sg13g2_fill_2 FILLER_26_1605 ();
 sg13g2_fill_2 FILLER_26_1612 ();
 sg13g2_fill_2 FILLER_26_1628 ();
 sg13g2_fill_1 FILLER_26_1637 ();
 sg13g2_decap_8 FILLER_26_1643 ();
 sg13g2_decap_4 FILLER_26_1650 ();
 sg13g2_fill_2 FILLER_26_1654 ();
 sg13g2_decap_8 FILLER_26_1682 ();
 sg13g2_fill_2 FILLER_26_1689 ();
 sg13g2_decap_4 FILLER_26_1698 ();
 sg13g2_fill_2 FILLER_26_1702 ();
 sg13g2_decap_4 FILLER_26_1709 ();
 sg13g2_fill_1 FILLER_26_1713 ();
 sg13g2_fill_2 FILLER_26_1724 ();
 sg13g2_fill_2 FILLER_26_1733 ();
 sg13g2_fill_1 FILLER_26_1735 ();
 sg13g2_decap_8 FILLER_26_1746 ();
 sg13g2_decap_8 FILLER_26_1753 ();
 sg13g2_decap_8 FILLER_26_1760 ();
 sg13g2_fill_1 FILLER_26_1767 ();
 sg13g2_decap_4 FILLER_26_1777 ();
 sg13g2_fill_2 FILLER_26_1781 ();
 sg13g2_fill_1 FILLER_26_1787 ();
 sg13g2_decap_4 FILLER_26_1800 ();
 sg13g2_fill_1 FILLER_26_1804 ();
 sg13g2_fill_1 FILLER_26_1817 ();
 sg13g2_fill_2 FILLER_26_1827 ();
 sg13g2_fill_1 FILLER_26_1829 ();
 sg13g2_fill_2 FILLER_26_1844 ();
 sg13g2_fill_1 FILLER_26_1846 ();
 sg13g2_fill_1 FILLER_26_1856 ();
 sg13g2_fill_1 FILLER_26_1862 ();
 sg13g2_fill_1 FILLER_26_1883 ();
 sg13g2_fill_1 FILLER_26_1909 ();
 sg13g2_fill_1 FILLER_26_1918 ();
 sg13g2_fill_1 FILLER_26_1944 ();
 sg13g2_fill_2 FILLER_26_1949 ();
 sg13g2_fill_1 FILLER_26_1951 ();
 sg13g2_decap_8 FILLER_26_1973 ();
 sg13g2_decap_8 FILLER_26_1980 ();
 sg13g2_fill_2 FILLER_26_1987 ();
 sg13g2_decap_8 FILLER_26_2003 ();
 sg13g2_fill_2 FILLER_26_2010 ();
 sg13g2_fill_1 FILLER_26_2012 ();
 sg13g2_fill_2 FILLER_26_2023 ();
 sg13g2_fill_1 FILLER_26_2025 ();
 sg13g2_decap_8 FILLER_26_2058 ();
 sg13g2_fill_2 FILLER_26_2082 ();
 sg13g2_fill_1 FILLER_26_2084 ();
 sg13g2_fill_1 FILLER_26_2098 ();
 sg13g2_decap_8 FILLER_26_2107 ();
 sg13g2_decap_8 FILLER_26_2114 ();
 sg13g2_decap_4 FILLER_26_2121 ();
 sg13g2_fill_1 FILLER_26_2125 ();
 sg13g2_decap_4 FILLER_26_2136 ();
 sg13g2_decap_8 FILLER_26_2144 ();
 sg13g2_fill_2 FILLER_26_2151 ();
 sg13g2_decap_8 FILLER_26_2183 ();
 sg13g2_fill_2 FILLER_26_2190 ();
 sg13g2_fill_1 FILLER_26_2192 ();
 sg13g2_decap_4 FILLER_26_2203 ();
 sg13g2_fill_1 FILLER_26_2211 ();
 sg13g2_fill_1 FILLER_26_2217 ();
 sg13g2_decap_8 FILLER_26_2244 ();
 sg13g2_decap_8 FILLER_26_2251 ();
 sg13g2_fill_1 FILLER_26_2258 ();
 sg13g2_fill_2 FILLER_26_2309 ();
 sg13g2_fill_2 FILLER_26_2359 ();
 sg13g2_fill_1 FILLER_26_2361 ();
 sg13g2_fill_1 FILLER_26_2394 ();
 sg13g2_decap_4 FILLER_26_2422 ();
 sg13g2_fill_1 FILLER_26_2426 ();
 sg13g2_fill_2 FILLER_26_2453 ();
 sg13g2_fill_2 FILLER_26_2465 ();
 sg13g2_fill_2 FILLER_26_2493 ();
 sg13g2_fill_2 FILLER_26_2501 ();
 sg13g2_fill_2 FILLER_26_2533 ();
 sg13g2_fill_1 FILLER_26_2535 ();
 sg13g2_fill_2 FILLER_26_2542 ();
 sg13g2_fill_2 FILLER_26_2580 ();
 sg13g2_fill_1 FILLER_26_2644 ();
 sg13g2_decap_8 FILLER_26_2659 ();
 sg13g2_decap_4 FILLER_26_2666 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_19 ();
 sg13g2_decap_8 FILLER_27_26 ();
 sg13g2_decap_8 FILLER_27_33 ();
 sg13g2_fill_1 FILLER_27_50 ();
 sg13g2_fill_1 FILLER_27_74 ();
 sg13g2_decap_4 FILLER_27_88 ();
 sg13g2_fill_2 FILLER_27_92 ();
 sg13g2_fill_2 FILLER_27_125 ();
 sg13g2_decap_4 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_140 ();
 sg13g2_decap_4 FILLER_27_146 ();
 sg13g2_fill_1 FILLER_27_155 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_4 FILLER_27_175 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_fill_2 FILLER_27_289 ();
 sg13g2_fill_2 FILLER_27_303 ();
 sg13g2_fill_1 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_315 ();
 sg13g2_fill_1 FILLER_27_356 ();
 sg13g2_fill_1 FILLER_27_370 ();
 sg13g2_fill_1 FILLER_27_380 ();
 sg13g2_fill_2 FILLER_27_412 ();
 sg13g2_fill_1 FILLER_27_417 ();
 sg13g2_decap_4 FILLER_27_436 ();
 sg13g2_fill_1 FILLER_27_440 ();
 sg13g2_decap_8 FILLER_27_446 ();
 sg13g2_fill_2 FILLER_27_453 ();
 sg13g2_fill_1 FILLER_27_455 ();
 sg13g2_decap_8 FILLER_27_466 ();
 sg13g2_fill_2 FILLER_27_478 ();
 sg13g2_fill_2 FILLER_27_484 ();
 sg13g2_fill_1 FILLER_27_489 ();
 sg13g2_fill_1 FILLER_27_509 ();
 sg13g2_decap_8 FILLER_27_514 ();
 sg13g2_fill_2 FILLER_27_521 ();
 sg13g2_fill_1 FILLER_27_561 ();
 sg13g2_fill_2 FILLER_27_609 ();
 sg13g2_fill_1 FILLER_27_611 ();
 sg13g2_fill_2 FILLER_27_631 ();
 sg13g2_fill_1 FILLER_27_646 ();
 sg13g2_fill_1 FILLER_27_653 ();
 sg13g2_fill_1 FILLER_27_664 ();
 sg13g2_fill_1 FILLER_27_669 ();
 sg13g2_fill_1 FILLER_27_685 ();
 sg13g2_decap_8 FILLER_27_702 ();
 sg13g2_decap_8 FILLER_27_709 ();
 sg13g2_decap_8 FILLER_27_769 ();
 sg13g2_decap_4 FILLER_27_776 ();
 sg13g2_fill_1 FILLER_27_780 ();
 sg13g2_decap_8 FILLER_27_818 ();
 sg13g2_decap_8 FILLER_27_825 ();
 sg13g2_decap_8 FILLER_27_832 ();
 sg13g2_decap_8 FILLER_27_839 ();
 sg13g2_fill_1 FILLER_27_846 ();
 sg13g2_fill_2 FILLER_27_857 ();
 sg13g2_fill_1 FILLER_27_863 ();
 sg13g2_fill_2 FILLER_27_890 ();
 sg13g2_decap_8 FILLER_27_896 ();
 sg13g2_fill_2 FILLER_27_903 ();
 sg13g2_decap_8 FILLER_27_951 ();
 sg13g2_fill_2 FILLER_27_958 ();
 sg13g2_fill_1 FILLER_27_960 ();
 sg13g2_decap_4 FILLER_27_978 ();
 sg13g2_fill_1 FILLER_27_1011 ();
 sg13g2_fill_2 FILLER_27_1017 ();
 sg13g2_fill_2 FILLER_27_1032 ();
 sg13g2_fill_1 FILLER_27_1038 ();
 sg13g2_decap_8 FILLER_27_1047 ();
 sg13g2_decap_4 FILLER_27_1062 ();
 sg13g2_fill_1 FILLER_27_1066 ();
 sg13g2_fill_1 FILLER_27_1093 ();
 sg13g2_fill_2 FILLER_27_1120 ();
 sg13g2_fill_1 FILLER_27_1122 ();
 sg13g2_fill_1 FILLER_27_1148 ();
 sg13g2_fill_2 FILLER_27_1158 ();
 sg13g2_fill_1 FILLER_27_1160 ();
 sg13g2_fill_2 FILLER_27_1221 ();
 sg13g2_decap_4 FILLER_27_1258 ();
 sg13g2_fill_1 FILLER_27_1262 ();
 sg13g2_decap_8 FILLER_27_1267 ();
 sg13g2_fill_2 FILLER_27_1321 ();
 sg13g2_fill_1 FILLER_27_1323 ();
 sg13g2_decap_8 FILLER_27_1348 ();
 sg13g2_fill_2 FILLER_27_1359 ();
 sg13g2_fill_1 FILLER_27_1371 ();
 sg13g2_fill_1 FILLER_27_1411 ();
 sg13g2_decap_8 FILLER_27_1417 ();
 sg13g2_fill_2 FILLER_27_1424 ();
 sg13g2_fill_1 FILLER_27_1426 ();
 sg13g2_decap_4 FILLER_27_1470 ();
 sg13g2_fill_2 FILLER_27_1474 ();
 sg13g2_fill_2 FILLER_27_1480 ();
 sg13g2_fill_1 FILLER_27_1482 ();
 sg13g2_fill_2 FILLER_27_1487 ();
 sg13g2_fill_1 FILLER_27_1489 ();
 sg13g2_decap_8 FILLER_27_1597 ();
 sg13g2_decap_8 FILLER_27_1604 ();
 sg13g2_decap_4 FILLER_27_1611 ();
 sg13g2_fill_1 FILLER_27_1615 ();
 sg13g2_decap_4 FILLER_27_1624 ();
 sg13g2_fill_1 FILLER_27_1632 ();
 sg13g2_fill_1 FILLER_27_1676 ();
 sg13g2_decap_8 FILLER_27_1681 ();
 sg13g2_decap_4 FILLER_27_1688 ();
 sg13g2_fill_1 FILLER_27_1692 ();
 sg13g2_fill_1 FILLER_27_1697 ();
 sg13g2_decap_8 FILLER_27_1738 ();
 sg13g2_decap_8 FILLER_27_1749 ();
 sg13g2_decap_8 FILLER_27_1756 ();
 sg13g2_decap_8 FILLER_27_1763 ();
 sg13g2_fill_1 FILLER_27_1788 ();
 sg13g2_fill_1 FILLER_27_1816 ();
 sg13g2_fill_2 FILLER_27_1836 ();
 sg13g2_fill_1 FILLER_27_1838 ();
 sg13g2_fill_2 FILLER_27_1843 ();
 sg13g2_fill_1 FILLER_27_1845 ();
 sg13g2_fill_2 FILLER_27_1859 ();
 sg13g2_decap_4 FILLER_27_1870 ();
 sg13g2_fill_2 FILLER_27_1883 ();
 sg13g2_fill_2 FILLER_27_1899 ();
 sg13g2_fill_1 FILLER_27_1901 ();
 sg13g2_fill_1 FILLER_27_1945 ();
 sg13g2_fill_1 FILLER_27_1953 ();
 sg13g2_fill_2 FILLER_27_1968 ();
 sg13g2_decap_8 FILLER_27_1974 ();
 sg13g2_decap_8 FILLER_27_1981 ();
 sg13g2_decap_8 FILLER_27_1988 ();
 sg13g2_decap_4 FILLER_27_1995 ();
 sg13g2_decap_4 FILLER_27_2009 ();
 sg13g2_fill_1 FILLER_27_2013 ();
 sg13g2_decap_8 FILLER_27_2019 ();
 sg13g2_decap_8 FILLER_27_2026 ();
 sg13g2_decap_8 FILLER_27_2033 ();
 sg13g2_decap_4 FILLER_27_2070 ();
 sg13g2_decap_8 FILLER_27_2120 ();
 sg13g2_decap_4 FILLER_27_2127 ();
 sg13g2_fill_1 FILLER_27_2131 ();
 sg13g2_decap_8 FILLER_27_2137 ();
 sg13g2_decap_8 FILLER_27_2144 ();
 sg13g2_fill_2 FILLER_27_2151 ();
 sg13g2_fill_1 FILLER_27_2153 ();
 sg13g2_decap_8 FILLER_27_2244 ();
 sg13g2_fill_1 FILLER_27_2251 ();
 sg13g2_fill_2 FILLER_27_2260 ();
 sg13g2_fill_1 FILLER_27_2262 ();
 sg13g2_fill_1 FILLER_27_2267 ();
 sg13g2_fill_2 FILLER_27_2271 ();
 sg13g2_fill_1 FILLER_27_2273 ();
 sg13g2_decap_8 FILLER_27_2283 ();
 sg13g2_decap_8 FILLER_27_2290 ();
 sg13g2_fill_2 FILLER_27_2297 ();
 sg13g2_fill_1 FILLER_27_2299 ();
 sg13g2_fill_1 FILLER_27_2338 ();
 sg13g2_fill_2 FILLER_27_2349 ();
 sg13g2_decap_4 FILLER_27_2356 ();
 sg13g2_decap_4 FILLER_27_2370 ();
 sg13g2_decap_4 FILLER_27_2384 ();
 sg13g2_fill_2 FILLER_27_2407 ();
 sg13g2_fill_1 FILLER_27_2409 ();
 sg13g2_decap_4 FILLER_27_2426 ();
 sg13g2_fill_1 FILLER_27_2462 ();
 sg13g2_fill_1 FILLER_27_2468 ();
 sg13g2_fill_1 FILLER_27_2473 ();
 sg13g2_fill_1 FILLER_27_2500 ();
 sg13g2_fill_1 FILLER_27_2511 ();
 sg13g2_fill_1 FILLER_27_2518 ();
 sg13g2_fill_2 FILLER_27_2525 ();
 sg13g2_fill_1 FILLER_27_2527 ();
 sg13g2_fill_2 FILLER_27_2536 ();
 sg13g2_fill_1 FILLER_27_2538 ();
 sg13g2_fill_2 FILLER_27_2549 ();
 sg13g2_decap_4 FILLER_27_2569 ();
 sg13g2_fill_2 FILLER_27_2583 ();
 sg13g2_fill_1 FILLER_27_2585 ();
 sg13g2_decap_4 FILLER_27_2596 ();
 sg13g2_fill_1 FILLER_27_2600 ();
 sg13g2_decap_8 FILLER_27_2652 ();
 sg13g2_decap_8 FILLER_27_2659 ();
 sg13g2_decap_4 FILLER_27_2666 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_4 ();
 sg13g2_fill_2 FILLER_28_31 ();
 sg13g2_fill_1 FILLER_28_33 ();
 sg13g2_fill_1 FILLER_28_62 ();
 sg13g2_fill_1 FILLER_28_81 ();
 sg13g2_fill_1 FILLER_28_95 ();
 sg13g2_fill_2 FILLER_28_138 ();
 sg13g2_decap_4 FILLER_28_148 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_decap_8 FILLER_28_157 ();
 sg13g2_decap_8 FILLER_28_164 ();
 sg13g2_decap_4 FILLER_28_171 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_decap_8 FILLER_28_226 ();
 sg13g2_decap_8 FILLER_28_233 ();
 sg13g2_decap_8 FILLER_28_244 ();
 sg13g2_decap_8 FILLER_28_251 ();
 sg13g2_decap_8 FILLER_28_258 ();
 sg13g2_fill_2 FILLER_28_265 ();
 sg13g2_fill_1 FILLER_28_272 ();
 sg13g2_fill_1 FILLER_28_277 ();
 sg13g2_fill_1 FILLER_28_287 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_fill_2 FILLER_28_336 ();
 sg13g2_fill_1 FILLER_28_348 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_fill_1 FILLER_28_359 ();
 sg13g2_fill_1 FILLER_28_369 ();
 sg13g2_fill_1 FILLER_28_386 ();
 sg13g2_fill_2 FILLER_28_397 ();
 sg13g2_fill_1 FILLER_28_423 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_fill_1 FILLER_28_430 ();
 sg13g2_decap_8 FILLER_28_434 ();
 sg13g2_fill_1 FILLER_28_441 ();
 sg13g2_decap_4 FILLER_28_453 ();
 sg13g2_decap_4 FILLER_28_469 ();
 sg13g2_fill_1 FILLER_28_473 ();
 sg13g2_fill_2 FILLER_28_500 ();
 sg13g2_fill_2 FILLER_28_517 ();
 sg13g2_fill_2 FILLER_28_527 ();
 sg13g2_fill_1 FILLER_28_529 ();
 sg13g2_fill_2 FILLER_28_540 ();
 sg13g2_fill_1 FILLER_28_555 ();
 sg13g2_decap_4 FILLER_28_562 ();
 sg13g2_fill_2 FILLER_28_598 ();
 sg13g2_fill_1 FILLER_28_600 ();
 sg13g2_fill_2 FILLER_28_614 ();
 sg13g2_fill_1 FILLER_28_616 ();
 sg13g2_fill_1 FILLER_28_621 ();
 sg13g2_fill_1 FILLER_28_632 ();
 sg13g2_fill_1 FILLER_28_665 ();
 sg13g2_fill_1 FILLER_28_685 ();
 sg13g2_decap_4 FILLER_28_701 ();
 sg13g2_fill_1 FILLER_28_705 ();
 sg13g2_decap_8 FILLER_28_710 ();
 sg13g2_fill_1 FILLER_28_717 ();
 sg13g2_decap_8 FILLER_28_774 ();
 sg13g2_decap_4 FILLER_28_781 ();
 sg13g2_fill_2 FILLER_28_785 ();
 sg13g2_fill_2 FILLER_28_816 ();
 sg13g2_fill_1 FILLER_28_818 ();
 sg13g2_decap_4 FILLER_28_842 ();
 sg13g2_fill_2 FILLER_28_846 ();
 sg13g2_fill_2 FILLER_28_874 ();
 sg13g2_fill_2 FILLER_28_890 ();
 sg13g2_fill_2 FILLER_28_1004 ();
 sg13g2_decap_8 FILLER_28_1032 ();
 sg13g2_decap_8 FILLER_28_1039 ();
 sg13g2_fill_2 FILLER_28_1046 ();
 sg13g2_fill_1 FILLER_28_1048 ();
 sg13g2_decap_4 FILLER_28_1053 ();
 sg13g2_fill_1 FILLER_28_1066 ();
 sg13g2_fill_2 FILLER_28_1076 ();
 sg13g2_fill_1 FILLER_28_1078 ();
 sg13g2_fill_2 FILLER_28_1100 ();
 sg13g2_decap_8 FILLER_28_1133 ();
 sg13g2_fill_1 FILLER_28_1140 ();
 sg13g2_fill_2 FILLER_28_1180 ();
 sg13g2_fill_1 FILLER_28_1182 ();
 sg13g2_fill_2 FILLER_28_1204 ();
 sg13g2_fill_1 FILLER_28_1206 ();
 sg13g2_fill_2 FILLER_28_1212 ();
 sg13g2_decap_4 FILLER_28_1239 ();
 sg13g2_decap_8 FILLER_28_1248 ();
 sg13g2_fill_2 FILLER_28_1255 ();
 sg13g2_decap_4 FILLER_28_1261 ();
 sg13g2_fill_2 FILLER_28_1275 ();
 sg13g2_fill_2 FILLER_28_1281 ();
 sg13g2_fill_1 FILLER_28_1283 ();
 sg13g2_decap_4 FILLER_28_1294 ();
 sg13g2_fill_1 FILLER_28_1328 ();
 sg13g2_decap_4 FILLER_28_1337 ();
 sg13g2_decap_8 FILLER_28_1351 ();
 sg13g2_fill_2 FILLER_28_1449 ();
 sg13g2_fill_2 FILLER_28_1506 ();
 sg13g2_fill_1 FILLER_28_1515 ();
 sg13g2_fill_1 FILLER_28_1529 ();
 sg13g2_fill_2 FILLER_28_1545 ();
 sg13g2_fill_1 FILLER_28_1567 ();
 sg13g2_fill_1 FILLER_28_1572 ();
 sg13g2_fill_1 FILLER_28_1581 ();
 sg13g2_fill_1 FILLER_28_1616 ();
 sg13g2_decap_4 FILLER_28_1627 ();
 sg13g2_fill_2 FILLER_28_1631 ();
 sg13g2_decap_8 FILLER_28_1645 ();
 sg13g2_decap_8 FILLER_28_1652 ();
 sg13g2_decap_8 FILLER_28_1659 ();
 sg13g2_decap_4 FILLER_28_1666 ();
 sg13g2_fill_2 FILLER_28_1703 ();
 sg13g2_fill_1 FILLER_28_1705 ();
 sg13g2_decap_8 FILLER_28_1720 ();
 sg13g2_decap_4 FILLER_28_1727 ();
 sg13g2_fill_1 FILLER_28_1735 ();
 sg13g2_fill_1 FILLER_28_1766 ();
 sg13g2_fill_1 FILLER_28_1772 ();
 sg13g2_fill_1 FILLER_28_1782 ();
 sg13g2_fill_2 FILLER_28_1806 ();
 sg13g2_fill_1 FILLER_28_1808 ();
 sg13g2_fill_2 FILLER_28_1819 ();
 sg13g2_fill_1 FILLER_28_1821 ();
 sg13g2_fill_2 FILLER_28_1827 ();
 sg13g2_fill_1 FILLER_28_1834 ();
 sg13g2_fill_1 FILLER_28_1840 ();
 sg13g2_fill_1 FILLER_28_1850 ();
 sg13g2_decap_4 FILLER_28_1855 ();
 sg13g2_fill_1 FILLER_28_1864 ();
 sg13g2_fill_1 FILLER_28_1871 ();
 sg13g2_fill_1 FILLER_28_1878 ();
 sg13g2_fill_1 FILLER_28_1889 ();
 sg13g2_fill_2 FILLER_28_1899 ();
 sg13g2_fill_1 FILLER_28_1901 ();
 sg13g2_fill_1 FILLER_28_1908 ();
 sg13g2_fill_2 FILLER_28_1916 ();
 sg13g2_fill_2 FILLER_28_1967 ();
 sg13g2_decap_8 FILLER_28_1974 ();
 sg13g2_decap_4 FILLER_28_2011 ();
 sg13g2_fill_2 FILLER_28_2015 ();
 sg13g2_decap_4 FILLER_28_2027 ();
 sg13g2_fill_1 FILLER_28_2031 ();
 sg13g2_decap_4 FILLER_28_2046 ();
 sg13g2_fill_1 FILLER_28_2050 ();
 sg13g2_fill_2 FILLER_28_2076 ();
 sg13g2_fill_1 FILLER_28_2102 ();
 sg13g2_decap_4 FILLER_28_2111 ();
 sg13g2_fill_1 FILLER_28_2115 ();
 sg13g2_decap_8 FILLER_28_2129 ();
 sg13g2_decap_4 FILLER_28_2136 ();
 sg13g2_fill_2 FILLER_28_2145 ();
 sg13g2_fill_2 FILLER_28_2160 ();
 sg13g2_fill_1 FILLER_28_2162 ();
 sg13g2_fill_1 FILLER_28_2181 ();
 sg13g2_decap_8 FILLER_28_2203 ();
 sg13g2_decap_4 FILLER_28_2210 ();
 sg13g2_fill_1 FILLER_28_2214 ();
 sg13g2_decap_8 FILLER_28_2266 ();
 sg13g2_decap_4 FILLER_28_2273 ();
 sg13g2_fill_2 FILLER_28_2277 ();
 sg13g2_decap_8 FILLER_28_2315 ();
 sg13g2_fill_2 FILLER_28_2322 ();
 sg13g2_fill_1 FILLER_28_2324 ();
 sg13g2_fill_1 FILLER_28_2339 ();
 sg13g2_fill_1 FILLER_28_2345 ();
 sg13g2_decap_8 FILLER_28_2351 ();
 sg13g2_decap_4 FILLER_28_2358 ();
 sg13g2_fill_2 FILLER_28_2362 ();
 sg13g2_fill_2 FILLER_28_2383 ();
 sg13g2_decap_8 FILLER_28_2425 ();
 sg13g2_fill_1 FILLER_28_2432 ();
 sg13g2_fill_1 FILLER_28_2437 ();
 sg13g2_decap_8 FILLER_28_2446 ();
 sg13g2_decap_8 FILLER_28_2453 ();
 sg13g2_fill_2 FILLER_28_2460 ();
 sg13g2_fill_1 FILLER_28_2462 ();
 sg13g2_fill_1 FILLER_28_2473 ();
 sg13g2_fill_1 FILLER_28_2484 ();
 sg13g2_decap_4 FILLER_28_2511 ();
 sg13g2_fill_1 FILLER_28_2515 ();
 sg13g2_fill_1 FILLER_28_2542 ();
 sg13g2_decap_4 FILLER_28_2569 ();
 sg13g2_decap_8 FILLER_28_2583 ();
 sg13g2_decap_4 FILLER_28_2590 ();
 sg13g2_decap_8 FILLER_28_2609 ();
 sg13g2_fill_1 FILLER_28_2620 ();
 sg13g2_fill_1 FILLER_28_2625 ();
 sg13g2_decap_8 FILLER_28_2662 ();
 sg13g2_fill_1 FILLER_28_2669 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_1 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_40 ();
 sg13g2_fill_2 FILLER_29_61 ();
 sg13g2_fill_1 FILLER_29_72 ();
 sg13g2_decap_8 FILLER_29_219 ();
 sg13g2_decap_4 FILLER_29_229 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_decap_8 FILLER_29_255 ();
 sg13g2_decap_8 FILLER_29_262 ();
 sg13g2_fill_1 FILLER_29_269 ();
 sg13g2_decap_4 FILLER_29_274 ();
 sg13g2_fill_2 FILLER_29_331 ();
 sg13g2_fill_1 FILLER_29_359 ();
 sg13g2_fill_1 FILLER_29_368 ();
 sg13g2_fill_2 FILLER_29_380 ();
 sg13g2_fill_1 FILLER_29_452 ();
 sg13g2_fill_1 FILLER_29_484 ();
 sg13g2_fill_1 FILLER_29_547 ();
 sg13g2_fill_1 FILLER_29_564 ();
 sg13g2_decap_4 FILLER_29_616 ();
 sg13g2_fill_2 FILLER_29_669 ();
 sg13g2_fill_1 FILLER_29_671 ();
 sg13g2_fill_2 FILLER_29_702 ();
 sg13g2_fill_1 FILLER_29_704 ();
 sg13g2_decap_8 FILLER_29_770 ();
 sg13g2_decap_4 FILLER_29_777 ();
 sg13g2_decap_4 FILLER_29_827 ();
 sg13g2_decap_4 FILLER_29_857 ();
 sg13g2_fill_1 FILLER_29_861 ();
 sg13g2_decap_4 FILLER_29_947 ();
 sg13g2_fill_1 FILLER_29_1000 ();
 sg13g2_fill_1 FILLER_29_1011 ();
 sg13g2_decap_8 FILLER_29_1016 ();
 sg13g2_decap_8 FILLER_29_1023 ();
 sg13g2_decap_8 FILLER_29_1030 ();
 sg13g2_fill_2 FILLER_29_1037 ();
 sg13g2_fill_1 FILLER_29_1096 ();
 sg13g2_decap_4 FILLER_29_1149 ();
 sg13g2_decap_4 FILLER_29_1183 ();
 sg13g2_fill_1 FILLER_29_1191 ();
 sg13g2_fill_1 FILLER_29_1201 ();
 sg13g2_fill_2 FILLER_29_1236 ();
 sg13g2_fill_1 FILLER_29_1238 ();
 sg13g2_decap_4 FILLER_29_1275 ();
 sg13g2_fill_1 FILLER_29_1279 ();
 sg13g2_decap_4 FILLER_29_1284 ();
 sg13g2_fill_2 FILLER_29_1298 ();
 sg13g2_decap_4 FILLER_29_1304 ();
 sg13g2_fill_2 FILLER_29_1354 ();
 sg13g2_decap_4 FILLER_29_1386 ();
 sg13g2_fill_2 FILLER_29_1390 ();
 sg13g2_decap_8 FILLER_29_1406 ();
 sg13g2_decap_8 FILLER_29_1413 ();
 sg13g2_fill_1 FILLER_29_1434 ();
 sg13g2_fill_1 FILLER_29_1440 ();
 sg13g2_fill_1 FILLER_29_1445 ();
 sg13g2_decap_4 FILLER_29_1498 ();
 sg13g2_fill_1 FILLER_29_1502 ();
 sg13g2_decap_4 FILLER_29_1507 ();
 sg13g2_fill_1 FILLER_29_1511 ();
 sg13g2_fill_1 FILLER_29_1515 ();
 sg13g2_fill_2 FILLER_29_1522 ();
 sg13g2_fill_2 FILLER_29_1543 ();
 sg13g2_fill_1 FILLER_29_1583 ();
 sg13g2_fill_1 FILLER_29_1589 ();
 sg13g2_fill_2 FILLER_29_1594 ();
 sg13g2_decap_8 FILLER_29_1611 ();
 sg13g2_decap_8 FILLER_29_1618 ();
 sg13g2_fill_1 FILLER_29_1625 ();
 sg13g2_decap_8 FILLER_29_1630 ();
 sg13g2_decap_8 FILLER_29_1637 ();
 sg13g2_decap_8 FILLER_29_1644 ();
 sg13g2_decap_8 FILLER_29_1655 ();
 sg13g2_fill_2 FILLER_29_1662 ();
 sg13g2_fill_1 FILLER_29_1664 ();
 sg13g2_fill_2 FILLER_29_1673 ();
 sg13g2_fill_1 FILLER_29_1701 ();
 sg13g2_decap_8 FILLER_29_1728 ();
 sg13g2_decap_4 FILLER_29_1735 ();
 sg13g2_fill_2 FILLER_29_1743 ();
 sg13g2_fill_1 FILLER_29_1745 ();
 sg13g2_decap_8 FILLER_29_1751 ();
 sg13g2_decap_8 FILLER_29_1758 ();
 sg13g2_decap_8 FILLER_29_1765 ();
 sg13g2_fill_2 FILLER_29_1830 ();
 sg13g2_fill_1 FILLER_29_1852 ();
 sg13g2_fill_1 FILLER_29_1861 ();
 sg13g2_fill_2 FILLER_29_1867 ();
 sg13g2_fill_1 FILLER_29_1874 ();
 sg13g2_fill_1 FILLER_29_1888 ();
 sg13g2_fill_1 FILLER_29_1893 ();
 sg13g2_fill_1 FILLER_29_1899 ();
 sg13g2_fill_1 FILLER_29_1905 ();
 sg13g2_fill_2 FILLER_29_1911 ();
 sg13g2_decap_8 FILLER_29_1918 ();
 sg13g2_fill_2 FILLER_29_1935 ();
 sg13g2_fill_1 FILLER_29_1967 ();
 sg13g2_decap_8 FILLER_29_1973 ();
 sg13g2_decap_8 FILLER_29_1980 ();
 sg13g2_decap_8 FILLER_29_1991 ();
 sg13g2_fill_2 FILLER_29_1998 ();
 sg13g2_fill_2 FILLER_29_2119 ();
 sg13g2_fill_1 FILLER_29_2121 ();
 sg13g2_fill_2 FILLER_29_2127 ();
 sg13g2_fill_1 FILLER_29_2129 ();
 sg13g2_decap_4 FILLER_29_2134 ();
 sg13g2_fill_1 FILLER_29_2138 ();
 sg13g2_decap_8 FILLER_29_2152 ();
 sg13g2_decap_8 FILLER_29_2185 ();
 sg13g2_decap_8 FILLER_29_2196 ();
 sg13g2_decap_8 FILLER_29_2203 ();
 sg13g2_decap_8 FILLER_29_2210 ();
 sg13g2_decap_4 FILLER_29_2217 ();
 sg13g2_fill_2 FILLER_29_2221 ();
 sg13g2_decap_4 FILLER_29_2263 ();
 sg13g2_fill_2 FILLER_29_2309 ();
 sg13g2_fill_2 FILLER_29_2333 ();
 sg13g2_decap_8 FILLER_29_2347 ();
 sg13g2_fill_1 FILLER_29_2354 ();
 sg13g2_fill_1 FILLER_29_2381 ();
 sg13g2_fill_1 FILLER_29_2392 ();
 sg13g2_fill_1 FILLER_29_2419 ();
 sg13g2_fill_1 FILLER_29_2430 ();
 sg13g2_fill_2 FILLER_29_2463 ();
 sg13g2_fill_1 FILLER_29_2465 ();
 sg13g2_fill_1 FILLER_29_2475 ();
 sg13g2_fill_1 FILLER_29_2480 ();
 sg13g2_fill_1 FILLER_29_2485 ();
 sg13g2_fill_1 FILLER_29_2491 ();
 sg13g2_fill_2 FILLER_29_2496 ();
 sg13g2_fill_2 FILLER_29_2502 ();
 sg13g2_decap_4 FILLER_29_2520 ();
 sg13g2_fill_1 FILLER_29_2524 ();
 sg13g2_fill_1 FILLER_29_2538 ();
 sg13g2_decap_4 FILLER_29_2545 ();
 sg13g2_fill_1 FILLER_29_2549 ();
 sg13g2_fill_2 FILLER_29_2554 ();
 sg13g2_fill_1 FILLER_29_2556 ();
 sg13g2_decap_4 FILLER_29_2567 ();
 sg13g2_fill_2 FILLER_29_2571 ();
 sg13g2_decap_4 FILLER_29_2609 ();
 sg13g2_fill_2 FILLER_29_2618 ();
 sg13g2_fill_2 FILLER_29_2630 ();
 sg13g2_fill_2 FILLER_29_2668 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_17 ();
 sg13g2_decap_4 FILLER_30_24 ();
 sg13g2_fill_1 FILLER_30_35 ();
 sg13g2_fill_2 FILLER_30_51 ();
 sg13g2_fill_1 FILLER_30_53 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_fill_1 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_fill_1 FILLER_30_178 ();
 sg13g2_fill_1 FILLER_30_186 ();
 sg13g2_fill_1 FILLER_30_194 ();
 sg13g2_fill_1 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_219 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_decap_4 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_279 ();
 sg13g2_fill_2 FILLER_30_305 ();
 sg13g2_fill_1 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_341 ();
 sg13g2_fill_2 FILLER_30_380 ();
 sg13g2_fill_1 FILLER_30_449 ();
 sg13g2_fill_2 FILLER_30_476 ();
 sg13g2_fill_1 FILLER_30_496 ();
 sg13g2_fill_2 FILLER_30_531 ();
 sg13g2_fill_2 FILLER_30_559 ();
 sg13g2_fill_2 FILLER_30_587 ();
 sg13g2_fill_1 FILLER_30_589 ();
 sg13g2_fill_1 FILLER_30_605 ();
 sg13g2_fill_1 FILLER_30_615 ();
 sg13g2_decap_4 FILLER_30_631 ();
 sg13g2_fill_2 FILLER_30_647 ();
 sg13g2_fill_1 FILLER_30_649 ();
 sg13g2_decap_4 FILLER_30_657 ();
 sg13g2_fill_2 FILLER_30_661 ();
 sg13g2_fill_2 FILLER_30_693 ();
 sg13g2_fill_2 FILLER_30_782 ();
 sg13g2_fill_1 FILLER_30_784 ();
 sg13g2_fill_2 FILLER_30_825 ();
 sg13g2_decap_4 FILLER_30_848 ();
 sg13g2_fill_2 FILLER_30_852 ();
 sg13g2_fill_2 FILLER_30_887 ();
 sg13g2_fill_1 FILLER_30_949 ();
 sg13g2_fill_1 FILLER_30_974 ();
 sg13g2_fill_1 FILLER_30_991 ();
 sg13g2_decap_8 FILLER_30_1025 ();
 sg13g2_decap_4 FILLER_30_1032 ();
 sg13g2_fill_2 FILLER_30_1036 ();
 sg13g2_fill_1 FILLER_30_1076 ();
 sg13g2_fill_1 FILLER_30_1081 ();
 sg13g2_fill_2 FILLER_30_1122 ();
 sg13g2_fill_2 FILLER_30_1137 ();
 sg13g2_fill_1 FILLER_30_1139 ();
 sg13g2_decap_4 FILLER_30_1148 ();
 sg13g2_fill_1 FILLER_30_1152 ();
 sg13g2_fill_2 FILLER_30_1166 ();
 sg13g2_fill_1 FILLER_30_1168 ();
 sg13g2_decap_8 FILLER_30_1233 ();
 sg13g2_decap_8 FILLER_30_1240 ();
 sg13g2_fill_1 FILLER_30_1247 ();
 sg13g2_decap_8 FILLER_30_1278 ();
 sg13g2_fill_2 FILLER_30_1285 ();
 sg13g2_fill_1 FILLER_30_1287 ();
 sg13g2_decap_4 FILLER_30_1314 ();
 sg13g2_fill_1 FILLER_30_1318 ();
 sg13g2_decap_8 FILLER_30_1349 ();
 sg13g2_decap_4 FILLER_30_1356 ();
 sg13g2_fill_2 FILLER_30_1360 ();
 sg13g2_fill_2 FILLER_30_1380 ();
 sg13g2_decap_8 FILLER_30_1392 ();
 sg13g2_fill_1 FILLER_30_1399 ();
 sg13g2_fill_2 FILLER_30_1426 ();
 sg13g2_fill_1 FILLER_30_1443 ();
 sg13g2_decap_4 FILLER_30_1448 ();
 sg13g2_fill_2 FILLER_30_1452 ();
 sg13g2_fill_1 FILLER_30_1460 ();
 sg13g2_fill_2 FILLER_30_1468 ();
 sg13g2_fill_1 FILLER_30_1484 ();
 sg13g2_fill_2 FILLER_30_1490 ();
 sg13g2_fill_1 FILLER_30_1535 ();
 sg13g2_fill_2 FILLER_30_1540 ();
 sg13g2_fill_2 FILLER_30_1590 ();
 sg13g2_fill_2 FILLER_30_1602 ();
 sg13g2_fill_2 FILLER_30_1648 ();
 sg13g2_decap_4 FILLER_30_1655 ();
 sg13g2_decap_8 FILLER_30_1663 ();
 sg13g2_fill_2 FILLER_30_1670 ();
 sg13g2_fill_1 FILLER_30_1672 ();
 sg13g2_fill_1 FILLER_30_1681 ();
 sg13g2_decap_4 FILLER_30_1686 ();
 sg13g2_decap_8 FILLER_30_1694 ();
 sg13g2_fill_2 FILLER_30_1701 ();
 sg13g2_decap_4 FILLER_30_1715 ();
 sg13g2_decap_4 FILLER_30_1753 ();
 sg13g2_fill_2 FILLER_30_1757 ();
 sg13g2_fill_2 FILLER_30_1773 ();
 sg13g2_fill_1 FILLER_30_1775 ();
 sg13g2_fill_1 FILLER_30_1786 ();
 sg13g2_fill_2 FILLER_30_1800 ();
 sg13g2_fill_2 FILLER_30_1824 ();
 sg13g2_fill_2 FILLER_30_1832 ();
 sg13g2_fill_1 FILLER_30_1834 ();
 sg13g2_fill_2 FILLER_30_1841 ();
 sg13g2_fill_1 FILLER_30_1843 ();
 sg13g2_fill_1 FILLER_30_1860 ();
 sg13g2_fill_1 FILLER_30_1868 ();
 sg13g2_fill_2 FILLER_30_1874 ();
 sg13g2_fill_2 FILLER_30_1880 ();
 sg13g2_fill_1 FILLER_30_1887 ();
 sg13g2_fill_2 FILLER_30_1893 ();
 sg13g2_fill_1 FILLER_30_1904 ();
 sg13g2_fill_2 FILLER_30_1909 ();
 sg13g2_decap_8 FILLER_30_1927 ();
 sg13g2_decap_4 FILLER_30_1934 ();
 sg13g2_fill_2 FILLER_30_1970 ();
 sg13g2_decap_8 FILLER_30_1976 ();
 sg13g2_fill_1 FILLER_30_1983 ();
 sg13g2_fill_2 FILLER_30_1988 ();
 sg13g2_decap_8 FILLER_30_2028 ();
 sg13g2_fill_2 FILLER_30_2035 ();
 sg13g2_fill_2 FILLER_30_2057 ();
 sg13g2_fill_1 FILLER_30_2059 ();
 sg13g2_fill_1 FILLER_30_2089 ();
 sg13g2_fill_2 FILLER_30_2118 ();
 sg13g2_fill_1 FILLER_30_2120 ();
 sg13g2_decap_8 FILLER_30_2156 ();
 sg13g2_decap_4 FILLER_30_2163 ();
 sg13g2_fill_1 FILLER_30_2193 ();
 sg13g2_fill_1 FILLER_30_2240 ();
 sg13g2_fill_2 FILLER_30_2251 ();
 sg13g2_decap_8 FILLER_30_2266 ();
 sg13g2_decap_4 FILLER_30_2273 ();
 sg13g2_fill_1 FILLER_30_2277 ();
 sg13g2_fill_1 FILLER_30_2290 ();
 sg13g2_decap_8 FILLER_30_2316 ();
 sg13g2_fill_2 FILLER_30_2349 ();
 sg13g2_decap_4 FILLER_30_2396 ();
 sg13g2_decap_8 FILLER_30_2446 ();
 sg13g2_decap_4 FILLER_30_2453 ();
 sg13g2_fill_1 FILLER_30_2457 ();
 sg13g2_fill_1 FILLER_30_2473 ();
 sg13g2_decap_8 FILLER_30_2487 ();
 sg13g2_decap_8 FILLER_30_2498 ();
 sg13g2_decap_8 FILLER_30_2505 ();
 sg13g2_fill_2 FILLER_30_2512 ();
 sg13g2_fill_1 FILLER_30_2514 ();
 sg13g2_fill_2 FILLER_30_2587 ();
 sg13g2_decap_8 FILLER_30_2625 ();
 sg13g2_decap_8 FILLER_30_2662 ();
 sg13g2_fill_1 FILLER_30_2669 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_34 ();
 sg13g2_fill_1 FILLER_31_36 ();
 sg13g2_fill_1 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_69 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_fill_2 FILLER_31_107 ();
 sg13g2_decap_4 FILLER_31_147 ();
 sg13g2_fill_1 FILLER_31_214 ();
 sg13g2_fill_1 FILLER_31_275 ();
 sg13g2_fill_2 FILLER_31_355 ();
 sg13g2_fill_1 FILLER_31_410 ();
 sg13g2_fill_1 FILLER_31_454 ();
 sg13g2_fill_2 FILLER_31_471 ();
 sg13g2_fill_2 FILLER_31_484 ();
 sg13g2_fill_1 FILLER_31_493 ();
 sg13g2_fill_1 FILLER_31_498 ();
 sg13g2_fill_1 FILLER_31_527 ();
 sg13g2_fill_2 FILLER_31_534 ();
 sg13g2_fill_1 FILLER_31_572 ();
 sg13g2_fill_1 FILLER_31_634 ();
 sg13g2_decap_8 FILLER_31_651 ();
 sg13g2_fill_1 FILLER_31_658 ();
 sg13g2_fill_1 FILLER_31_667 ();
 sg13g2_fill_1 FILLER_31_671 ();
 sg13g2_decap_8 FILLER_31_677 ();
 sg13g2_decap_8 FILLER_31_684 ();
 sg13g2_decap_8 FILLER_31_691 ();
 sg13g2_decap_4 FILLER_31_698 ();
 sg13g2_fill_2 FILLER_31_702 ();
 sg13g2_decap_8 FILLER_31_708 ();
 sg13g2_decap_8 FILLER_31_715 ();
 sg13g2_decap_8 FILLER_31_722 ();
 sg13g2_fill_2 FILLER_31_729 ();
 sg13g2_decap_8 FILLER_31_735 ();
 sg13g2_decap_8 FILLER_31_742 ();
 sg13g2_decap_4 FILLER_31_749 ();
 sg13g2_fill_2 FILLER_31_761 ();
 sg13g2_fill_1 FILLER_31_763 ();
 sg13g2_fill_1 FILLER_31_768 ();
 sg13g2_fill_2 FILLER_31_795 ();
 sg13g2_fill_1 FILLER_31_915 ();
 sg13g2_fill_1 FILLER_31_965 ();
 sg13g2_fill_2 FILLER_31_1038 ();
 sg13g2_fill_1 FILLER_31_1040 ();
 sg13g2_fill_2 FILLER_31_1050 ();
 sg13g2_fill_1 FILLER_31_1052 ();
 sg13g2_fill_2 FILLER_31_1063 ();
 sg13g2_fill_2 FILLER_31_1070 ();
 sg13g2_fill_1 FILLER_31_1072 ();
 sg13g2_fill_1 FILLER_31_1081 ();
 sg13g2_decap_8 FILLER_31_1086 ();
 sg13g2_decap_4 FILLER_31_1093 ();
 sg13g2_fill_1 FILLER_31_1101 ();
 sg13g2_fill_1 FILLER_31_1106 ();
 sg13g2_decap_8 FILLER_31_1115 ();
 sg13g2_decap_8 FILLER_31_1135 ();
 sg13g2_fill_1 FILLER_31_1142 ();
 sg13g2_fill_2 FILLER_31_1146 ();
 sg13g2_fill_1 FILLER_31_1148 ();
 sg13g2_fill_1 FILLER_31_1188 ();
 sg13g2_fill_2 FILLER_31_1193 ();
 sg13g2_fill_2 FILLER_31_1198 ();
 sg13g2_fill_1 FILLER_31_1200 ();
 sg13g2_decap_4 FILLER_31_1205 ();
 sg13g2_fill_1 FILLER_31_1209 ();
 sg13g2_decap_4 FILLER_31_1222 ();
 sg13g2_fill_2 FILLER_31_1226 ();
 sg13g2_fill_2 FILLER_31_1232 ();
 sg13g2_fill_2 FILLER_31_1244 ();
 sg13g2_fill_2 FILLER_31_1256 ();
 sg13g2_decap_4 FILLER_31_1268 ();
 sg13g2_decap_4 FILLER_31_1298 ();
 sg13g2_decap_8 FILLER_31_1306 ();
 sg13g2_fill_2 FILLER_31_1313 ();
 sg13g2_fill_1 FILLER_31_1315 ();
 sg13g2_fill_2 FILLER_31_1407 ();
 sg13g2_fill_1 FILLER_31_1409 ();
 sg13g2_decap_4 FILLER_31_1414 ();
 sg13g2_fill_1 FILLER_31_1418 ();
 sg13g2_fill_2 FILLER_31_1463 ();
 sg13g2_decap_8 FILLER_31_1629 ();
 sg13g2_fill_2 FILLER_31_1636 ();
 sg13g2_fill_1 FILLER_31_1643 ();
 sg13g2_decap_4 FILLER_31_1725 ();
 sg13g2_fill_2 FILLER_31_1729 ();
 sg13g2_decap_8 FILLER_31_1766 ();
 sg13g2_decap_8 FILLER_31_1773 ();
 sg13g2_fill_2 FILLER_31_1780 ();
 sg13g2_fill_1 FILLER_31_1795 ();
 sg13g2_fill_2 FILLER_31_1824 ();
 sg13g2_fill_1 FILLER_31_1826 ();
 sg13g2_fill_1 FILLER_31_1847 ();
 sg13g2_fill_2 FILLER_31_1853 ();
 sg13g2_fill_2 FILLER_31_1872 ();
 sg13g2_fill_1 FILLER_31_1874 ();
 sg13g2_fill_1 FILLER_31_1879 ();
 sg13g2_fill_1 FILLER_31_1885 ();
 sg13g2_fill_1 FILLER_31_1891 ();
 sg13g2_fill_2 FILLER_31_1901 ();
 sg13g2_fill_1 FILLER_31_1903 ();
 sg13g2_fill_2 FILLER_31_1912 ();
 sg13g2_fill_1 FILLER_31_1914 ();
 sg13g2_decap_4 FILLER_31_1921 ();
 sg13g2_fill_1 FILLER_31_1925 ();
 sg13g2_decap_8 FILLER_31_1973 ();
 sg13g2_fill_1 FILLER_31_1980 ();
 sg13g2_fill_1 FILLER_31_2011 ();
 sg13g2_decap_8 FILLER_31_2038 ();
 sg13g2_decap_4 FILLER_31_2045 ();
 sg13g2_fill_1 FILLER_31_2049 ();
 sg13g2_fill_2 FILLER_31_2126 ();
 sg13g2_fill_2 FILLER_31_2146 ();
 sg13g2_decap_8 FILLER_31_2184 ();
 sg13g2_decap_8 FILLER_31_2272 ();
 sg13g2_fill_2 FILLER_31_2291 ();
 sg13g2_fill_1 FILLER_31_2293 ();
 sg13g2_fill_1 FILLER_31_2299 ();
 sg13g2_fill_1 FILLER_31_2305 ();
 sg13g2_decap_8 FILLER_31_2350 ();
 sg13g2_decap_8 FILLER_31_2381 ();
 sg13g2_fill_2 FILLER_31_2388 ();
 sg13g2_decap_8 FILLER_31_2395 ();
 sg13g2_decap_8 FILLER_31_2402 ();
 sg13g2_decap_4 FILLER_31_2409 ();
 sg13g2_fill_1 FILLER_31_2413 ();
 sg13g2_fill_1 FILLER_31_2443 ();
 sg13g2_fill_2 FILLER_31_2484 ();
 sg13g2_decap_4 FILLER_31_2490 ();
 sg13g2_fill_2 FILLER_31_2494 ();
 sg13g2_fill_2 FILLER_31_2502 ();
 sg13g2_fill_2 FILLER_31_2520 ();
 sg13g2_fill_1 FILLER_31_2522 ();
 sg13g2_fill_2 FILLER_31_2543 ();
 sg13g2_fill_1 FILLER_31_2581 ();
 sg13g2_decap_8 FILLER_31_2596 ();
 sg13g2_fill_2 FILLER_31_2603 ();
 sg13g2_decap_8 FILLER_31_2625 ();
 sg13g2_fill_2 FILLER_31_2668 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_2 ();
 sg13g2_fill_2 FILLER_32_29 ();
 sg13g2_fill_2 FILLER_32_35 ();
 sg13g2_fill_1 FILLER_32_46 ();
 sg13g2_fill_1 FILLER_32_50 ();
 sg13g2_fill_1 FILLER_32_68 ();
 sg13g2_fill_2 FILLER_32_73 ();
 sg13g2_fill_1 FILLER_32_90 ();
 sg13g2_fill_1 FILLER_32_105 ();
 sg13g2_decap_4 FILLER_32_137 ();
 sg13g2_fill_2 FILLER_32_141 ();
 sg13g2_decap_8 FILLER_32_151 ();
 sg13g2_decap_8 FILLER_32_158 ();
 sg13g2_decap_4 FILLER_32_165 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_fill_2 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_197 ();
 sg13g2_fill_1 FILLER_32_203 ();
 sg13g2_fill_1 FILLER_32_211 ();
 sg13g2_fill_1 FILLER_32_255 ();
 sg13g2_fill_2 FILLER_32_282 ();
 sg13g2_fill_2 FILLER_32_366 ();
 sg13g2_fill_2 FILLER_32_432 ();
 sg13g2_fill_2 FILLER_32_438 ();
 sg13g2_fill_1 FILLER_32_444 ();
 sg13g2_fill_2 FILLER_32_461 ();
 sg13g2_fill_1 FILLER_32_493 ();
 sg13g2_fill_2 FILLER_32_506 ();
 sg13g2_fill_1 FILLER_32_524 ();
 sg13g2_fill_2 FILLER_32_538 ();
 sg13g2_fill_2 FILLER_32_560 ();
 sg13g2_fill_1 FILLER_32_568 ();
 sg13g2_fill_1 FILLER_32_572 ();
 sg13g2_fill_2 FILLER_32_579 ();
 sg13g2_fill_1 FILLER_32_585 ();
 sg13g2_fill_1 FILLER_32_612 ();
 sg13g2_decap_8 FILLER_32_661 ();
 sg13g2_fill_1 FILLER_32_668 ();
 sg13g2_fill_1 FILLER_32_684 ();
 sg13g2_decap_4 FILLER_32_701 ();
 sg13g2_fill_2 FILLER_32_705 ();
 sg13g2_decap_8 FILLER_32_724 ();
 sg13g2_decap_8 FILLER_32_731 ();
 sg13g2_decap_8 FILLER_32_738 ();
 sg13g2_decap_8 FILLER_32_745 ();
 sg13g2_decap_4 FILLER_32_752 ();
 sg13g2_fill_2 FILLER_32_756 ();
 sg13g2_decap_8 FILLER_32_763 ();
 sg13g2_decap_4 FILLER_32_770 ();
 sg13g2_fill_2 FILLER_32_778 ();
 sg13g2_decap_4 FILLER_32_815 ();
 sg13g2_fill_2 FILLER_32_853 ();
 sg13g2_fill_2 FILLER_32_973 ();
 sg13g2_fill_1 FILLER_32_1011 ();
 sg13g2_fill_1 FILLER_32_1038 ();
 sg13g2_fill_2 FILLER_32_1070 ();
 sg13g2_fill_1 FILLER_32_1077 ();
 sg13g2_fill_1 FILLER_32_1083 ();
 sg13g2_decap_8 FILLER_32_1088 ();
 sg13g2_decap_4 FILLER_32_1095 ();
 sg13g2_fill_2 FILLER_32_1099 ();
 sg13g2_fill_1 FILLER_32_1105 ();
 sg13g2_fill_1 FILLER_32_1111 ();
 sg13g2_fill_1 FILLER_32_1116 ();
 sg13g2_fill_1 FILLER_32_1138 ();
 sg13g2_fill_2 FILLER_32_1146 ();
 sg13g2_decap_8 FILLER_32_1196 ();
 sg13g2_decap_8 FILLER_32_1203 ();
 sg13g2_fill_2 FILLER_32_1210 ();
 sg13g2_decap_4 FILLER_32_1217 ();
 sg13g2_fill_1 FILLER_32_1221 ();
 sg13g2_fill_2 FILLER_32_1282 ();
 sg13g2_fill_1 FILLER_32_1284 ();
 sg13g2_decap_8 FILLER_32_1321 ();
 sg13g2_decap_8 FILLER_32_1352 ();
 sg13g2_decap_8 FILLER_32_1359 ();
 sg13g2_fill_2 FILLER_32_1366 ();
 sg13g2_fill_1 FILLER_32_1368 ();
 sg13g2_decap_4 FILLER_32_1374 ();
 sg13g2_fill_2 FILLER_32_1378 ();
 sg13g2_fill_2 FILLER_32_1393 ();
 sg13g2_fill_1 FILLER_32_1395 ();
 sg13g2_fill_1 FILLER_32_1422 ();
 sg13g2_fill_2 FILLER_32_1449 ();
 sg13g2_fill_2 FILLER_32_1455 ();
 sg13g2_fill_1 FILLER_32_1480 ();
 sg13g2_fill_2 FILLER_32_1486 ();
 sg13g2_fill_1 FILLER_32_1488 ();
 sg13g2_fill_2 FILLER_32_1494 ();
 sg13g2_fill_1 FILLER_32_1501 ();
 sg13g2_fill_1 FILLER_32_1506 ();
 sg13g2_fill_2 FILLER_32_1515 ();
 sg13g2_fill_1 FILLER_32_1522 ();
 sg13g2_fill_1 FILLER_32_1532 ();
 sg13g2_fill_2 FILLER_32_1549 ();
 sg13g2_fill_2 FILLER_32_1559 ();
 sg13g2_fill_2 FILLER_32_1617 ();
 sg13g2_decap_8 FILLER_32_1688 ();
 sg13g2_decap_8 FILLER_32_1699 ();
 sg13g2_decap_8 FILLER_32_1706 ();
 sg13g2_decap_4 FILLER_32_1718 ();
 sg13g2_fill_2 FILLER_32_1722 ();
 sg13g2_decap_4 FILLER_32_1754 ();
 sg13g2_fill_1 FILLER_32_1758 ();
 sg13g2_decap_8 FILLER_32_1762 ();
 sg13g2_decap_8 FILLER_32_1769 ();
 sg13g2_decap_8 FILLER_32_1776 ();
 sg13g2_fill_2 FILLER_32_1783 ();
 sg13g2_fill_1 FILLER_32_1785 ();
 sg13g2_decap_8 FILLER_32_1849 ();
 sg13g2_fill_1 FILLER_32_1856 ();
 sg13g2_fill_1 FILLER_32_1871 ();
 sg13g2_fill_1 FILLER_32_1913 ();
 sg13g2_fill_1 FILLER_32_1920 ();
 sg13g2_fill_2 FILLER_32_1925 ();
 sg13g2_fill_1 FILLER_32_1931 ();
 sg13g2_fill_1 FILLER_32_1963 ();
 sg13g2_decap_8 FILLER_32_1978 ();
 sg13g2_decap_8 FILLER_32_1985 ();
 sg13g2_decap_8 FILLER_32_1992 ();
 sg13g2_fill_1 FILLER_32_1999 ();
 sg13g2_decap_8 FILLER_32_2024 ();
 sg13g2_decap_8 FILLER_32_2031 ();
 sg13g2_fill_1 FILLER_32_2079 ();
 sg13g2_fill_2 FILLER_32_2105 ();
 sg13g2_fill_2 FILLER_32_2182 ();
 sg13g2_fill_1 FILLER_32_2184 ();
 sg13g2_decap_4 FILLER_32_2206 ();
 sg13g2_fill_1 FILLER_32_2210 ();
 sg13g2_decap_8 FILLER_32_2228 ();
 sg13g2_decap_8 FILLER_32_2235 ();
 sg13g2_fill_2 FILLER_32_2242 ();
 sg13g2_fill_2 FILLER_32_2270 ();
 sg13g2_fill_1 FILLER_32_2272 ();
 sg13g2_fill_2 FILLER_32_2299 ();
 sg13g2_fill_1 FILLER_32_2301 ();
 sg13g2_fill_2 FILLER_32_2312 ();
 sg13g2_fill_2 FILLER_32_2326 ();
 sg13g2_fill_1 FILLER_32_2328 ();
 sg13g2_fill_2 FILLER_32_2334 ();
 sg13g2_fill_2 FILLER_32_2341 ();
 sg13g2_fill_2 FILLER_32_2351 ();
 sg13g2_fill_1 FILLER_32_2353 ();
 sg13g2_fill_1 FILLER_32_2380 ();
 sg13g2_fill_1 FILLER_32_2407 ();
 sg13g2_fill_1 FILLER_32_2412 ();
 sg13g2_fill_2 FILLER_32_2423 ();
 sg13g2_fill_1 FILLER_32_2459 ();
 sg13g2_decap_8 FILLER_32_2495 ();
 sg13g2_fill_1 FILLER_32_2502 ();
 sg13g2_decap_4 FILLER_32_2529 ();
 sg13g2_decap_8 FILLER_32_2567 ();
 sg13g2_decap_8 FILLER_32_2610 ();
 sg13g2_decap_8 FILLER_32_2617 ();
 sg13g2_decap_4 FILLER_32_2624 ();
 sg13g2_fill_1 FILLER_32_2628 ();
 sg13g2_decap_8 FILLER_32_2633 ();
 sg13g2_decap_4 FILLER_32_2644 ();
 sg13g2_fill_1 FILLER_32_2648 ();
 sg13g2_decap_8 FILLER_32_2653 ();
 sg13g2_decap_8 FILLER_32_2660 ();
 sg13g2_fill_2 FILLER_32_2667 ();
 sg13g2_fill_1 FILLER_32_2669 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_8 ();
 sg13g2_fill_1 FILLER_33_35 ();
 sg13g2_fill_2 FILLER_33_40 ();
 sg13g2_fill_1 FILLER_33_42 ();
 sg13g2_fill_2 FILLER_33_48 ();
 sg13g2_fill_2 FILLER_33_59 ();
 sg13g2_fill_1 FILLER_33_61 ();
 sg13g2_fill_2 FILLER_33_75 ();
 sg13g2_fill_1 FILLER_33_85 ();
 sg13g2_fill_2 FILLER_33_117 ();
 sg13g2_decap_4 FILLER_33_130 ();
 sg13g2_fill_2 FILLER_33_134 ();
 sg13g2_fill_2 FILLER_33_167 ();
 sg13g2_fill_1 FILLER_33_169 ();
 sg13g2_decap_8 FILLER_33_227 ();
 sg13g2_decap_4 FILLER_33_238 ();
 sg13g2_fill_1 FILLER_33_247 ();
 sg13g2_fill_1 FILLER_33_296 ();
 sg13g2_fill_2 FILLER_33_343 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_fill_2 FILLER_33_415 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_fill_1 FILLER_33_477 ();
 sg13g2_fill_2 FILLER_33_512 ();
 sg13g2_fill_1 FILLER_33_527 ();
 sg13g2_fill_2 FILLER_33_531 ();
 sg13g2_fill_2 FILLER_33_549 ();
 sg13g2_fill_1 FILLER_33_639 ();
 sg13g2_decap_4 FILLER_33_650 ();
 sg13g2_fill_2 FILLER_33_654 ();
 sg13g2_decap_8 FILLER_33_662 ();
 sg13g2_fill_1 FILLER_33_669 ();
 sg13g2_fill_1 FILLER_33_679 ();
 sg13g2_fill_2 FILLER_33_696 ();
 sg13g2_fill_1 FILLER_33_698 ();
 sg13g2_decap_4 FILLER_33_733 ();
 sg13g2_fill_1 FILLER_33_737 ();
 sg13g2_decap_8 FILLER_33_742 ();
 sg13g2_decap_4 FILLER_33_762 ();
 sg13g2_fill_2 FILLER_33_792 ();
 sg13g2_fill_1 FILLER_33_794 ();
 sg13g2_decap_4 FILLER_33_818 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_fill_1 FILLER_33_875 ();
 sg13g2_fill_2 FILLER_33_896 ();
 sg13g2_fill_1 FILLER_33_975 ();
 sg13g2_fill_1 FILLER_33_993 ();
 sg13g2_fill_1 FILLER_33_998 ();
 sg13g2_fill_2 FILLER_33_1020 ();
 sg13g2_fill_2 FILLER_33_1029 ();
 sg13g2_fill_2 FILLER_33_1100 ();
 sg13g2_fill_1 FILLER_33_1133 ();
 sg13g2_decap_4 FILLER_33_1165 ();
 sg13g2_fill_2 FILLER_33_1169 ();
 sg13g2_decap_8 FILLER_33_1183 ();
 sg13g2_decap_8 FILLER_33_1190 ();
 sg13g2_decap_8 FILLER_33_1197 ();
 sg13g2_decap_8 FILLER_33_1204 ();
 sg13g2_decap_8 FILLER_33_1211 ();
 sg13g2_decap_4 FILLER_33_1218 ();
 sg13g2_fill_1 FILLER_33_1222 ();
 sg13g2_decap_8 FILLER_33_1231 ();
 sg13g2_fill_2 FILLER_33_1243 ();
 sg13g2_fill_2 FILLER_33_1255 ();
 sg13g2_fill_2 FILLER_33_1261 ();
 sg13g2_decap_8 FILLER_33_1289 ();
 sg13g2_decap_8 FILLER_33_1296 ();
 sg13g2_decap_8 FILLER_33_1303 ();
 sg13g2_fill_1 FILLER_33_1310 ();
 sg13g2_decap_4 FILLER_33_1316 ();
 sg13g2_decap_4 FILLER_33_1334 ();
 sg13g2_decap_4 FILLER_33_1360 ();
 sg13g2_fill_1 FILLER_33_1390 ();
 sg13g2_fill_1 FILLER_33_1401 ();
 sg13g2_fill_1 FILLER_33_1406 ();
 sg13g2_fill_1 FILLER_33_1468 ();
 sg13g2_fill_2 FILLER_33_1474 ();
 sg13g2_fill_1 FILLER_33_1506 ();
 sg13g2_fill_1 FILLER_33_1538 ();
 sg13g2_fill_1 FILLER_33_1547 ();
 sg13g2_fill_2 FILLER_33_1604 ();
 sg13g2_decap_8 FILLER_33_1632 ();
 sg13g2_decap_8 FILLER_33_1639 ();
 sg13g2_fill_2 FILLER_33_1646 ();
 sg13g2_fill_1 FILLER_33_1648 ();
 sg13g2_decap_8 FILLER_33_1701 ();
 sg13g2_decap_8 FILLER_33_1708 ();
 sg13g2_decap_8 FILLER_33_1715 ();
 sg13g2_decap_4 FILLER_33_1722 ();
 sg13g2_fill_1 FILLER_33_1726 ();
 sg13g2_fill_1 FILLER_33_1749 ();
 sg13g2_fill_2 FILLER_33_1776 ();
 sg13g2_decap_8 FILLER_33_1781 ();
 sg13g2_fill_1 FILLER_33_1793 ();
 sg13g2_fill_1 FILLER_33_1803 ();
 sg13g2_fill_1 FILLER_33_1808 ();
 sg13g2_fill_2 FILLER_33_1819 ();
 sg13g2_fill_1 FILLER_33_1826 ();
 sg13g2_decap_4 FILLER_33_1833 ();
 sg13g2_fill_1 FILLER_33_1837 ();
 sg13g2_decap_4 FILLER_33_1851 ();
 sg13g2_fill_1 FILLER_33_1855 ();
 sg13g2_fill_1 FILLER_33_1865 ();
 sg13g2_fill_2 FILLER_33_1879 ();
 sg13g2_fill_1 FILLER_33_1881 ();
 sg13g2_fill_1 FILLER_33_1946 ();
 sg13g2_fill_2 FILLER_33_1961 ();
 sg13g2_fill_1 FILLER_33_1971 ();
 sg13g2_fill_2 FILLER_33_1980 ();
 sg13g2_decap_8 FILLER_33_2027 ();
 sg13g2_fill_2 FILLER_33_2034 ();
 sg13g2_decap_4 FILLER_33_2066 ();
 sg13g2_fill_2 FILLER_33_2070 ();
 sg13g2_fill_1 FILLER_33_2101 ();
 sg13g2_fill_1 FILLER_33_2158 ();
 sg13g2_decap_8 FILLER_33_2169 ();
 sg13g2_fill_2 FILLER_33_2176 ();
 sg13g2_decap_4 FILLER_33_2208 ();
 sg13g2_decap_8 FILLER_33_2258 ();
 sg13g2_decap_8 FILLER_33_2265 ();
 sg13g2_decap_8 FILLER_33_2272 ();
 sg13g2_fill_1 FILLER_33_2279 ();
 sg13g2_decap_4 FILLER_33_2284 ();
 sg13g2_fill_1 FILLER_33_2288 ();
 sg13g2_decap_8 FILLER_33_2299 ();
 sg13g2_decap_8 FILLER_33_2306 ();
 sg13g2_decap_8 FILLER_33_2313 ();
 sg13g2_decap_8 FILLER_33_2323 ();
 sg13g2_decap_8 FILLER_33_2330 ();
 sg13g2_fill_2 FILLER_33_2337 ();
 sg13g2_fill_1 FILLER_33_2339 ();
 sg13g2_fill_2 FILLER_33_2344 ();
 sg13g2_decap_8 FILLER_33_2352 ();
 sg13g2_fill_2 FILLER_33_2359 ();
 sg13g2_decap_8 FILLER_33_2365 ();
 sg13g2_decap_8 FILLER_33_2372 ();
 sg13g2_decap_8 FILLER_33_2379 ();
 sg13g2_fill_1 FILLER_33_2386 ();
 sg13g2_fill_2 FILLER_33_2400 ();
 sg13g2_fill_2 FILLER_33_2458 ();
 sg13g2_fill_2 FILLER_33_2477 ();
 sg13g2_decap_4 FILLER_33_2531 ();
 sg13g2_fill_1 FILLER_33_2535 ();
 sg13g2_decap_8 FILLER_33_2562 ();
 sg13g2_fill_1 FILLER_33_2569 ();
 sg13g2_decap_4 FILLER_33_2580 ();
 sg13g2_fill_1 FILLER_33_2584 ();
 sg13g2_fill_2 FILLER_33_2632 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_18 ();
 sg13g2_decap_8 FILLER_34_25 ();
 sg13g2_decap_8 FILLER_34_32 ();
 sg13g2_decap_8 FILLER_34_39 ();
 sg13g2_fill_2 FILLER_34_57 ();
 sg13g2_fill_1 FILLER_34_64 ();
 sg13g2_decap_4 FILLER_34_73 ();
 sg13g2_fill_1 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_97 ();
 sg13g2_fill_1 FILLER_34_111 ();
 sg13g2_decap_8 FILLER_34_141 ();
 sg13g2_fill_1 FILLER_34_181 ();
 sg13g2_fill_1 FILLER_34_187 ();
 sg13g2_fill_1 FILLER_34_193 ();
 sg13g2_fill_2 FILLER_34_202 ();
 sg13g2_fill_1 FILLER_34_204 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_decap_8 FILLER_34_227 ();
 sg13g2_fill_2 FILLER_34_237 ();
 sg13g2_decap_8 FILLER_34_242 ();
 sg13g2_decap_4 FILLER_34_249 ();
 sg13g2_fill_2 FILLER_34_253 ();
 sg13g2_fill_2 FILLER_34_260 ();
 sg13g2_fill_1 FILLER_34_274 ();
 sg13g2_fill_1 FILLER_34_293 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_fill_2 FILLER_34_377 ();
 sg13g2_fill_1 FILLER_34_432 ();
 sg13g2_fill_2 FILLER_34_452 ();
 sg13g2_fill_2 FILLER_34_459 ();
 sg13g2_fill_1 FILLER_34_473 ();
 sg13g2_fill_2 FILLER_34_544 ();
 sg13g2_fill_1 FILLER_34_572 ();
 sg13g2_fill_2 FILLER_34_606 ();
 sg13g2_fill_1 FILLER_34_632 ();
 sg13g2_fill_1 FILLER_34_643 ();
 sg13g2_fill_1 FILLER_34_650 ();
 sg13g2_fill_2 FILLER_34_659 ();
 sg13g2_fill_2 FILLER_34_680 ();
 sg13g2_fill_1 FILLER_34_693 ();
 sg13g2_decap_8 FILLER_34_777 ();
 sg13g2_fill_2 FILLER_34_784 ();
 sg13g2_fill_1 FILLER_34_880 ();
 sg13g2_fill_1 FILLER_34_902 ();
 sg13g2_fill_2 FILLER_34_908 ();
 sg13g2_fill_2 FILLER_34_926 ();
 sg13g2_fill_2 FILLER_34_966 ();
 sg13g2_fill_2 FILLER_34_1020 ();
 sg13g2_fill_1 FILLER_34_1139 ();
 sg13g2_fill_1 FILLER_34_1152 ();
 sg13g2_decap_8 FILLER_34_1166 ();
 sg13g2_decap_8 FILLER_34_1173 ();
 sg13g2_decap_8 FILLER_34_1180 ();
 sg13g2_decap_4 FILLER_34_1187 ();
 sg13g2_fill_2 FILLER_34_1191 ();
 sg13g2_fill_2 FILLER_34_1203 ();
 sg13g2_fill_1 FILLER_34_1205 ();
 sg13g2_decap_4 FILLER_34_1232 ();
 sg13g2_fill_2 FILLER_34_1236 ();
 sg13g2_decap_8 FILLER_34_1243 ();
 sg13g2_decap_4 FILLER_34_1250 ();
 sg13g2_fill_1 FILLER_34_1282 ();
 sg13g2_decap_4 FILLER_34_1309 ();
 sg13g2_fill_2 FILLER_34_1313 ();
 sg13g2_fill_2 FILLER_34_1348 ();
 sg13g2_decap_8 FILLER_34_1360 ();
 sg13g2_fill_1 FILLER_34_1367 ();
 sg13g2_fill_2 FILLER_34_1373 ();
 sg13g2_fill_1 FILLER_34_1375 ();
 sg13g2_decap_8 FILLER_34_1389 ();
 sg13g2_decap_8 FILLER_34_1396 ();
 sg13g2_fill_2 FILLER_34_1403 ();
 sg13g2_fill_1 FILLER_34_1405 ();
 sg13g2_fill_1 FILLER_34_1410 ();
 sg13g2_fill_2 FILLER_34_1424 ();
 sg13g2_fill_1 FILLER_34_1444 ();
 sg13g2_fill_2 FILLER_34_1450 ();
 sg13g2_fill_2 FILLER_34_1498 ();
 sg13g2_fill_1 FILLER_34_1546 ();
 sg13g2_fill_1 FILLER_34_1559 ();
 sg13g2_decap_4 FILLER_34_1623 ();
 sg13g2_fill_2 FILLER_34_1627 ();
 sg13g2_fill_1 FILLER_34_1689 ();
 sg13g2_decap_8 FILLER_34_1782 ();
 sg13g2_decap_4 FILLER_34_1789 ();
 sg13g2_decap_4 FILLER_34_1810 ();
 sg13g2_fill_2 FILLER_34_1823 ();
 sg13g2_fill_1 FILLER_34_1829 ();
 sg13g2_fill_1 FILLER_34_1854 ();
 sg13g2_fill_2 FILLER_34_1860 ();
 sg13g2_fill_1 FILLER_34_1870 ();
 sg13g2_fill_2 FILLER_34_1891 ();
 sg13g2_fill_1 FILLER_34_1902 ();
 sg13g2_fill_2 FILLER_34_1912 ();
 sg13g2_fill_1 FILLER_34_1931 ();
 sg13g2_decap_8 FILLER_34_1965 ();
 sg13g2_decap_8 FILLER_34_1972 ();
 sg13g2_decap_8 FILLER_34_1979 ();
 sg13g2_decap_4 FILLER_34_1986 ();
 sg13g2_fill_1 FILLER_34_1990 ();
 sg13g2_decap_4 FILLER_34_1996 ();
 sg13g2_fill_2 FILLER_34_2000 ();
 sg13g2_fill_1 FILLER_34_2093 ();
 sg13g2_fill_1 FILLER_34_2134 ();
 sg13g2_decap_8 FILLER_34_2161 ();
 sg13g2_decap_8 FILLER_34_2168 ();
 sg13g2_decap_4 FILLER_34_2175 ();
 sg13g2_fill_1 FILLER_34_2242 ();
 sg13g2_decap_8 FILLER_34_2260 ();
 sg13g2_decap_8 FILLER_34_2267 ();
 sg13g2_decap_8 FILLER_34_2274 ();
 sg13g2_fill_1 FILLER_34_2281 ();
 sg13g2_decap_8 FILLER_34_2362 ();
 sg13g2_decap_4 FILLER_34_2369 ();
 sg13g2_fill_1 FILLER_34_2373 ();
 sg13g2_decap_4 FILLER_34_2386 ();
 sg13g2_fill_1 FILLER_34_2429 ();
 sg13g2_fill_1 FILLER_34_2524 ();
 sg13g2_fill_1 FILLER_34_2534 ();
 sg13g2_fill_2 FILLER_34_2557 ();
 sg13g2_fill_2 FILLER_34_2570 ();
 sg13g2_decap_8 FILLER_34_2608 ();
 sg13g2_fill_2 FILLER_34_2615 ();
 sg13g2_fill_1 FILLER_34_2617 ();
 sg13g2_fill_2 FILLER_34_2644 ();
 sg13g2_fill_1 FILLER_34_2646 ();
 sg13g2_decap_8 FILLER_34_2655 ();
 sg13g2_decap_8 FILLER_34_2662 ();
 sg13g2_fill_1 FILLER_34_2669 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_37 ();
 sg13g2_fill_1 FILLER_35_98 ();
 sg13g2_fill_1 FILLER_35_142 ();
 sg13g2_fill_2 FILLER_35_153 ();
 sg13g2_fill_1 FILLER_35_155 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_fill_2 FILLER_35_172 ();
 sg13g2_decap_8 FILLER_35_178 ();
 sg13g2_decap_8 FILLER_35_185 ();
 sg13g2_decap_8 FILLER_35_192 ();
 sg13g2_decap_8 FILLER_35_199 ();
 sg13g2_decap_8 FILLER_35_206 ();
 sg13g2_decap_4 FILLER_35_213 ();
 sg13g2_fill_1 FILLER_35_221 ();
 sg13g2_decap_8 FILLER_35_227 ();
 sg13g2_decap_8 FILLER_35_243 ();
 sg13g2_decap_4 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_259 ();
 sg13g2_fill_1 FILLER_35_265 ();
 sg13g2_fill_2 FILLER_35_289 ();
 sg13g2_fill_1 FILLER_35_319 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_fill_1 FILLER_35_362 ();
 sg13g2_fill_1 FILLER_35_384 ();
 sg13g2_fill_1 FILLER_35_427 ();
 sg13g2_fill_2 FILLER_35_443 ();
 sg13g2_fill_1 FILLER_35_539 ();
 sg13g2_fill_1 FILLER_35_551 ();
 sg13g2_fill_2 FILLER_35_565 ();
 sg13g2_fill_2 FILLER_35_571 ();
 sg13g2_fill_2 FILLER_35_586 ();
 sg13g2_fill_1 FILLER_35_596 ();
 sg13g2_fill_2 FILLER_35_614 ();
 sg13g2_fill_1 FILLER_35_637 ();
 sg13g2_fill_1 FILLER_35_651 ();
 sg13g2_fill_2 FILLER_35_722 ();
 sg13g2_fill_2 FILLER_35_729 ();
 sg13g2_fill_2 FILLER_35_811 ();
 sg13g2_fill_2 FILLER_35_821 ();
 sg13g2_fill_1 FILLER_35_831 ();
 sg13g2_fill_2 FILLER_35_898 ();
 sg13g2_fill_2 FILLER_35_908 ();
 sg13g2_fill_1 FILLER_35_914 ();
 sg13g2_fill_2 FILLER_35_959 ();
 sg13g2_fill_1 FILLER_35_984 ();
 sg13g2_fill_1 FILLER_35_996 ();
 sg13g2_fill_1 FILLER_35_1003 ();
 sg13g2_fill_2 FILLER_35_1059 ();
 sg13g2_fill_2 FILLER_35_1068 ();
 sg13g2_fill_2 FILLER_35_1080 ();
 sg13g2_fill_1 FILLER_35_1125 ();
 sg13g2_fill_2 FILLER_35_1144 ();
 sg13g2_fill_2 FILLER_35_1210 ();
 sg13g2_decap_8 FILLER_35_1221 ();
 sg13g2_fill_1 FILLER_35_1228 ();
 sg13g2_decap_4 FILLER_35_1255 ();
 sg13g2_fill_1 FILLER_35_1259 ();
 sg13g2_fill_1 FILLER_35_1270 ();
 sg13g2_fill_1 FILLER_35_1285 ();
 sg13g2_fill_1 FILLER_35_1313 ();
 sg13g2_decap_4 FILLER_35_1368 ();
 sg13g2_fill_1 FILLER_35_1376 ();
 sg13g2_decap_4 FILLER_35_1387 ();
 sg13g2_fill_2 FILLER_35_1391 ();
 sg13g2_decap_4 FILLER_35_1437 ();
 sg13g2_fill_1 FILLER_35_1441 ();
 sg13g2_decap_8 FILLER_35_1451 ();
 sg13g2_fill_2 FILLER_35_1458 ();
 sg13g2_decap_4 FILLER_35_1463 ();
 sg13g2_fill_1 FILLER_35_1467 ();
 sg13g2_fill_2 FILLER_35_1486 ();
 sg13g2_fill_1 FILLER_35_1488 ();
 sg13g2_fill_1 FILLER_35_1495 ();
 sg13g2_fill_1 FILLER_35_1502 ();
 sg13g2_fill_1 FILLER_35_1506 ();
 sg13g2_fill_2 FILLER_35_1510 ();
 sg13g2_fill_1 FILLER_35_1602 ();
 sg13g2_decap_4 FILLER_35_1622 ();
 sg13g2_decap_4 FILLER_35_1638 ();
 sg13g2_fill_2 FILLER_35_1642 ();
 sg13g2_decap_4 FILLER_35_1651 ();
 sg13g2_fill_2 FILLER_35_1655 ();
 sg13g2_fill_2 FILLER_35_1666 ();
 sg13g2_fill_1 FILLER_35_1668 ();
 sg13g2_decap_4 FILLER_35_1673 ();
 sg13g2_fill_2 FILLER_35_1677 ();
 sg13g2_decap_4 FILLER_35_1689 ();
 sg13g2_fill_2 FILLER_35_1693 ();
 sg13g2_decap_4 FILLER_35_1705 ();
 sg13g2_decap_4 FILLER_35_1713 ();
 sg13g2_fill_1 FILLER_35_1722 ();
 sg13g2_decap_8 FILLER_35_1791 ();
 sg13g2_decap_8 FILLER_35_1798 ();
 sg13g2_fill_2 FILLER_35_1817 ();
 sg13g2_fill_1 FILLER_35_1824 ();
 sg13g2_fill_1 FILLER_35_1830 ();
 sg13g2_fill_2 FILLER_35_1836 ();
 sg13g2_fill_1 FILLER_35_1860 ();
 sg13g2_fill_2 FILLER_35_1874 ();
 sg13g2_fill_2 FILLER_35_1911 ();
 sg13g2_fill_1 FILLER_35_1913 ();
 sg13g2_fill_1 FILLER_35_1924 ();
 sg13g2_fill_2 FILLER_35_1945 ();
 sg13g2_fill_2 FILLER_35_1951 ();
 sg13g2_fill_1 FILLER_35_1953 ();
 sg13g2_decap_8 FILLER_35_1958 ();
 sg13g2_fill_2 FILLER_35_1965 ();
 sg13g2_decap_8 FILLER_35_1971 ();
 sg13g2_decap_8 FILLER_35_1978 ();
 sg13g2_fill_1 FILLER_35_1994 ();
 sg13g2_fill_2 FILLER_35_2025 ();
 sg13g2_fill_2 FILLER_35_2057 ();
 sg13g2_fill_2 FILLER_35_2098 ();
 sg13g2_fill_1 FILLER_35_2100 ();
 sg13g2_fill_1 FILLER_35_2108 ();
 sg13g2_decap_4 FILLER_35_2113 ();
 sg13g2_fill_1 FILLER_35_2117 ();
 sg13g2_decap_8 FILLER_35_2149 ();
 sg13g2_fill_2 FILLER_35_2156 ();
 sg13g2_fill_1 FILLER_35_2158 ();
 sg13g2_fill_2 FILLER_35_2163 ();
 sg13g2_decap_4 FILLER_35_2191 ();
 sg13g2_fill_1 FILLER_35_2195 ();
 sg13g2_fill_1 FILLER_35_2200 ();
 sg13g2_fill_2 FILLER_35_2227 ();
 sg13g2_fill_1 FILLER_35_2239 ();
 sg13g2_fill_2 FILLER_35_2266 ();
 sg13g2_fill_1 FILLER_35_2319 ();
 sg13g2_fill_2 FILLER_35_2363 ();
 sg13g2_decap_8 FILLER_35_2372 ();
 sg13g2_decap_8 FILLER_35_2379 ();
 sg13g2_fill_1 FILLER_35_2386 ();
 sg13g2_fill_2 FILLER_35_2477 ();
 sg13g2_fill_1 FILLER_35_2484 ();
 sg13g2_fill_2 FILLER_35_2497 ();
 sg13g2_fill_1 FILLER_35_2519 ();
 sg13g2_decap_8 FILLER_35_2579 ();
 sg13g2_decap_8 FILLER_35_2586 ();
 sg13g2_fill_1 FILLER_35_2593 ();
 sg13g2_fill_2 FILLER_35_2606 ();
 sg13g2_decap_4 FILLER_35_2664 ();
 sg13g2_fill_2 FILLER_35_2668 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_65 ();
 sg13g2_fill_2 FILLER_36_72 ();
 sg13g2_fill_1 FILLER_36_111 ();
 sg13g2_fill_1 FILLER_36_115 ();
 sg13g2_fill_1 FILLER_36_123 ();
 sg13g2_fill_1 FILLER_36_129 ();
 sg13g2_decap_8 FILLER_36_134 ();
 sg13g2_fill_2 FILLER_36_141 ();
 sg13g2_fill_1 FILLER_36_143 ();
 sg13g2_decap_4 FILLER_36_238 ();
 sg13g2_fill_1 FILLER_36_242 ();
 sg13g2_fill_2 FILLER_36_269 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_fill_2 FILLER_36_306 ();
 sg13g2_fill_1 FILLER_36_320 ();
 sg13g2_fill_2 FILLER_36_347 ();
 sg13g2_fill_1 FILLER_36_352 ();
 sg13g2_fill_1 FILLER_36_362 ();
 sg13g2_fill_2 FILLER_36_374 ();
 sg13g2_fill_1 FILLER_36_392 ();
 sg13g2_fill_2 FILLER_36_432 ();
 sg13g2_fill_1 FILLER_36_439 ();
 sg13g2_fill_1 FILLER_36_448 ();
 sg13g2_fill_2 FILLER_36_479 ();
 sg13g2_fill_2 FILLER_36_506 ();
 sg13g2_fill_1 FILLER_36_518 ();
 sg13g2_fill_1 FILLER_36_529 ();
 sg13g2_fill_1 FILLER_36_544 ();
 sg13g2_fill_2 FILLER_36_558 ();
 sg13g2_fill_1 FILLER_36_582 ();
 sg13g2_fill_2 FILLER_36_593 ();
 sg13g2_fill_2 FILLER_36_624 ();
 sg13g2_fill_2 FILLER_36_632 ();
 sg13g2_fill_2 FILLER_36_698 ();
 sg13g2_fill_1 FILLER_36_700 ();
 sg13g2_fill_1 FILLER_36_715 ();
 sg13g2_fill_2 FILLER_36_732 ();
 sg13g2_fill_2 FILLER_36_739 ();
 sg13g2_fill_1 FILLER_36_745 ();
 sg13g2_fill_1 FILLER_36_751 ();
 sg13g2_decap_8 FILLER_36_781 ();
 sg13g2_decap_8 FILLER_36_792 ();
 sg13g2_decap_8 FILLER_36_799 ();
 sg13g2_decap_8 FILLER_36_806 ();
 sg13g2_fill_1 FILLER_36_813 ();
 sg13g2_fill_1 FILLER_36_844 ();
 sg13g2_fill_2 FILLER_36_862 ();
 sg13g2_fill_1 FILLER_36_867 ();
 sg13g2_fill_1 FILLER_36_880 ();
 sg13g2_fill_1 FILLER_36_885 ();
 sg13g2_fill_2 FILLER_36_919 ();
 sg13g2_fill_2 FILLER_36_935 ();
 sg13g2_fill_2 FILLER_36_944 ();
 sg13g2_fill_1 FILLER_36_997 ();
 sg13g2_fill_2 FILLER_36_1068 ();
 sg13g2_fill_2 FILLER_36_1073 ();
 sg13g2_fill_1 FILLER_36_1087 ();
 sg13g2_fill_2 FILLER_36_1092 ();
 sg13g2_fill_2 FILLER_36_1115 ();
 sg13g2_fill_1 FILLER_36_1117 ();
 sg13g2_fill_2 FILLER_36_1171 ();
 sg13g2_fill_2 FILLER_36_1191 ();
 sg13g2_decap_8 FILLER_36_1219 ();
 sg13g2_fill_1 FILLER_36_1226 ();
 sg13g2_fill_2 FILLER_36_1231 ();
 sg13g2_fill_1 FILLER_36_1233 ();
 sg13g2_fill_1 FILLER_36_1238 ();
 sg13g2_fill_2 FILLER_36_1285 ();
 sg13g2_fill_2 FILLER_36_1321 ();
 sg13g2_fill_1 FILLER_36_1331 ();
 sg13g2_fill_2 FILLER_36_1345 ();
 sg13g2_fill_1 FILLER_36_1353 ();
 sg13g2_fill_1 FILLER_36_1359 ();
 sg13g2_fill_1 FILLER_36_1367 ();
 sg13g2_decap_4 FILLER_36_1386 ();
 sg13g2_fill_1 FILLER_36_1390 ();
 sg13g2_decap_8 FILLER_36_1431 ();
 sg13g2_fill_1 FILLER_36_1438 ();
 sg13g2_decap_8 FILLER_36_1443 ();
 sg13g2_fill_1 FILLER_36_1450 ();
 sg13g2_decap_8 FILLER_36_1460 ();
 sg13g2_decap_8 FILLER_36_1467 ();
 sg13g2_fill_1 FILLER_36_1474 ();
 sg13g2_fill_1 FILLER_36_1506 ();
 sg13g2_fill_2 FILLER_36_1515 ();
 sg13g2_fill_1 FILLER_36_1536 ();
 sg13g2_fill_2 FILLER_36_1569 ();
 sg13g2_fill_2 FILLER_36_1624 ();
 sg13g2_fill_2 FILLER_36_1631 ();
 sg13g2_fill_1 FILLER_36_1638 ();
 sg13g2_fill_2 FILLER_36_1665 ();
 sg13g2_decap_4 FILLER_36_1671 ();
 sg13g2_decap_8 FILLER_36_1680 ();
 sg13g2_decap_4 FILLER_36_1687 ();
 sg13g2_fill_1 FILLER_36_1691 ();
 sg13g2_decap_4 FILLER_36_1696 ();
 sg13g2_fill_1 FILLER_36_1726 ();
 sg13g2_fill_2 FILLER_36_1799 ();
 sg13g2_fill_2 FILLER_36_1869 ();
 sg13g2_fill_2 FILLER_36_1890 ();
 sg13g2_fill_1 FILLER_36_1906 ();
 sg13g2_fill_1 FILLER_36_1921 ();
 sg13g2_decap_8 FILLER_36_1957 ();
 sg13g2_decap_8 FILLER_36_1964 ();
 sg13g2_decap_4 FILLER_36_1971 ();
 sg13g2_fill_2 FILLER_36_1975 ();
 sg13g2_decap_8 FILLER_36_2038 ();
 sg13g2_fill_2 FILLER_36_2045 ();
 sg13g2_fill_1 FILLER_36_2061 ();
 sg13g2_decap_8 FILLER_36_2098 ();
 sg13g2_decap_8 FILLER_36_2105 ();
 sg13g2_decap_8 FILLER_36_2112 ();
 sg13g2_decap_8 FILLER_36_2137 ();
 sg13g2_fill_2 FILLER_36_2190 ();
 sg13g2_fill_1 FILLER_36_2192 ();
 sg13g2_decap_8 FILLER_36_2242 ();
 sg13g2_decap_8 FILLER_36_2249 ();
 sg13g2_decap_8 FILLER_36_2256 ();
 sg13g2_decap_4 FILLER_36_2263 ();
 sg13g2_fill_2 FILLER_36_2267 ();
 sg13g2_fill_2 FILLER_36_2276 ();
 sg13g2_fill_2 FILLER_36_2296 ();
 sg13g2_fill_1 FILLER_36_2312 ();
 sg13g2_fill_1 FILLER_36_2325 ();
 sg13g2_fill_1 FILLER_36_2330 ();
 sg13g2_fill_1 FILLER_36_2336 ();
 sg13g2_fill_1 FILLER_36_2363 ();
 sg13g2_fill_1 FILLER_36_2408 ();
 sg13g2_fill_1 FILLER_36_2484 ();
 sg13g2_fill_2 FILLER_36_2489 ();
 sg13g2_fill_1 FILLER_36_2491 ();
 sg13g2_fill_2 FILLER_36_2515 ();
 sg13g2_fill_1 FILLER_36_2590 ();
 sg13g2_decap_4 FILLER_36_2609 ();
 sg13g2_fill_2 FILLER_36_2613 ();
 sg13g2_fill_2 FILLER_36_2630 ();
 sg13g2_fill_2 FILLER_36_2668 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_15 ();
 sg13g2_decap_4 FILLER_37_47 ();
 sg13g2_fill_2 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_83 ();
 sg13g2_fill_2 FILLER_37_90 ();
 sg13g2_fill_2 FILLER_37_100 ();
 sg13g2_fill_1 FILLER_37_152 ();
 sg13g2_fill_2 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_223 ();
 sg13g2_fill_2 FILLER_37_230 ();
 sg13g2_fill_1 FILLER_37_232 ();
 sg13g2_decap_8 FILLER_37_243 ();
 sg13g2_fill_1 FILLER_37_250 ();
 sg13g2_fill_1 FILLER_37_259 ();
 sg13g2_fill_2 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_291 ();
 sg13g2_fill_1 FILLER_37_347 ();
 sg13g2_fill_1 FILLER_37_359 ();
 sg13g2_fill_2 FILLER_37_390 ();
 sg13g2_fill_2 FILLER_37_425 ();
 sg13g2_fill_2 FILLER_37_443 ();
 sg13g2_fill_1 FILLER_37_518 ();
 sg13g2_fill_2 FILLER_37_522 ();
 sg13g2_fill_1 FILLER_37_609 ();
 sg13g2_fill_1 FILLER_37_613 ();
 sg13g2_fill_1 FILLER_37_644 ();
 sg13g2_fill_1 FILLER_37_649 ();
 sg13g2_fill_1 FILLER_37_655 ();
 sg13g2_fill_2 FILLER_37_692 ();
 sg13g2_fill_1 FILLER_37_694 ();
 sg13g2_fill_1 FILLER_37_740 ();
 sg13g2_decap_8 FILLER_37_779 ();
 sg13g2_decap_8 FILLER_37_786 ();
 sg13g2_decap_8 FILLER_37_793 ();
 sg13g2_decap_8 FILLER_37_800 ();
 sg13g2_decap_8 FILLER_37_807 ();
 sg13g2_fill_2 FILLER_37_814 ();
 sg13g2_fill_1 FILLER_37_821 ();
 sg13g2_fill_1 FILLER_37_827 ();
 sg13g2_fill_1 FILLER_37_836 ();
 sg13g2_decap_8 FILLER_37_846 ();
 sg13g2_fill_2 FILLER_37_853 ();
 sg13g2_fill_2 FILLER_37_877 ();
 sg13g2_fill_2 FILLER_37_927 ();
 sg13g2_fill_1 FILLER_37_945 ();
 sg13g2_fill_2 FILLER_37_971 ();
 sg13g2_fill_2 FILLER_37_1006 ();
 sg13g2_fill_1 FILLER_37_1021 ();
 sg13g2_fill_1 FILLER_37_1032 ();
 sg13g2_fill_1 FILLER_37_1088 ();
 sg13g2_fill_2 FILLER_37_1105 ();
 sg13g2_fill_1 FILLER_37_1149 ();
 sg13g2_fill_1 FILLER_37_1172 ();
 sg13g2_fill_2 FILLER_37_1183 ();
 sg13g2_fill_1 FILLER_37_1185 ();
 sg13g2_fill_2 FILLER_37_1210 ();
 sg13g2_fill_1 FILLER_37_1212 ();
 sg13g2_fill_2 FILLER_37_1217 ();
 sg13g2_fill_1 FILLER_37_1219 ();
 sg13g2_decap_4 FILLER_37_1246 ();
 sg13g2_fill_1 FILLER_37_1276 ();
 sg13g2_fill_1 FILLER_37_1290 ();
 sg13g2_fill_1 FILLER_37_1309 ();
 sg13g2_fill_1 FILLER_37_1317 ();
 sg13g2_fill_2 FILLER_37_1325 ();
 sg13g2_fill_2 FILLER_37_1354 ();
 sg13g2_fill_1 FILLER_37_1356 ();
 sg13g2_fill_1 FILLER_37_1375 ();
 sg13g2_decap_8 FILLER_37_1381 ();
 sg13g2_decap_8 FILLER_37_1388 ();
 sg13g2_decap_8 FILLER_37_1395 ();
 sg13g2_fill_2 FILLER_37_1402 ();
 sg13g2_fill_1 FILLER_37_1409 ();
 sg13g2_fill_1 FILLER_37_1419 ();
 sg13g2_fill_2 FILLER_37_1433 ();
 sg13g2_fill_1 FILLER_37_1435 ();
 sg13g2_fill_2 FILLER_37_1449 ();
 sg13g2_fill_2 FILLER_37_1454 ();
 sg13g2_fill_2 FILLER_37_1461 ();
 sg13g2_fill_1 FILLER_37_1486 ();
 sg13g2_fill_1 FILLER_37_1491 ();
 sg13g2_fill_1 FILLER_37_1499 ();
 sg13g2_fill_2 FILLER_37_1510 ();
 sg13g2_fill_1 FILLER_37_1528 ();
 sg13g2_fill_1 FILLER_37_1554 ();
 sg13g2_fill_2 FILLER_37_1594 ();
 sg13g2_decap_8 FILLER_37_1634 ();
 sg13g2_fill_2 FILLER_37_1654 ();
 sg13g2_fill_1 FILLER_37_1656 ();
 sg13g2_fill_2 FILLER_37_1683 ();
 sg13g2_fill_1 FILLER_37_1685 ();
 sg13g2_decap_8 FILLER_37_1690 ();
 sg13g2_fill_1 FILLER_37_1697 ();
 sg13g2_fill_1 FILLER_37_1711 ();
 sg13g2_fill_2 FILLER_37_1717 ();
 sg13g2_fill_1 FILLER_37_1723 ();
 sg13g2_fill_1 FILLER_37_1739 ();
 sg13g2_fill_1 FILLER_37_1770 ();
 sg13g2_fill_2 FILLER_37_1809 ();
 sg13g2_fill_2 FILLER_37_1855 ();
 sg13g2_fill_1 FILLER_37_1866 ();
 sg13g2_fill_2 FILLER_37_1873 ();
 sg13g2_fill_2 FILLER_37_1885 ();
 sg13g2_fill_2 FILLER_37_1891 ();
 sg13g2_fill_2 FILLER_37_1902 ();
 sg13g2_fill_2 FILLER_37_1909 ();
 sg13g2_fill_1 FILLER_37_1921 ();
 sg13g2_fill_1 FILLER_37_1927 ();
 sg13g2_fill_1 FILLER_37_1933 ();
 sg13g2_decap_8 FILLER_37_1956 ();
 sg13g2_decap_8 FILLER_37_1963 ();
 sg13g2_fill_2 FILLER_37_1970 ();
 sg13g2_fill_2 FILLER_37_1998 ();
 sg13g2_fill_1 FILLER_37_2000 ();
 sg13g2_decap_4 FILLER_37_2027 ();
 sg13g2_fill_2 FILLER_37_2031 ();
 sg13g2_decap_4 FILLER_37_2043 ();
 sg13g2_fill_2 FILLER_37_2047 ();
 sg13g2_decap_4 FILLER_37_2059 ();
 sg13g2_fill_1 FILLER_37_2089 ();
 sg13g2_decap_4 FILLER_37_2094 ();
 sg13g2_fill_1 FILLER_37_2098 ();
 sg13g2_decap_4 FILLER_37_2109 ();
 sg13g2_fill_1 FILLER_37_2139 ();
 sg13g2_decap_8 FILLER_37_2248 ();
 sg13g2_decap_4 FILLER_37_2255 ();
 sg13g2_decap_8 FILLER_37_2263 ();
 sg13g2_decap_8 FILLER_37_2270 ();
 sg13g2_fill_1 FILLER_37_2277 ();
 sg13g2_fill_2 FILLER_37_2282 ();
 sg13g2_fill_1 FILLER_37_2383 ();
 sg13g2_fill_1 FILLER_37_2414 ();
 sg13g2_fill_2 FILLER_37_2509 ();
 sg13g2_fill_1 FILLER_37_2540 ();
 sg13g2_fill_2 FILLER_37_2547 ();
 sg13g2_fill_1 FILLER_37_2549 ();
 sg13g2_fill_2 FILLER_37_2556 ();
 sg13g2_fill_1 FILLER_37_2558 ();
 sg13g2_fill_2 FILLER_37_2563 ();
 sg13g2_fill_1 FILLER_37_2565 ();
 sg13g2_decap_4 FILLER_37_2597 ();
 sg13g2_fill_2 FILLER_37_2601 ();
 sg13g2_fill_1 FILLER_37_2611 ();
 sg13g2_decap_8 FILLER_37_2616 ();
 sg13g2_fill_1 FILLER_37_2623 ();
 sg13g2_fill_1 FILLER_37_2638 ();
 sg13g2_decap_4 FILLER_37_2665 ();
 sg13g2_fill_1 FILLER_37_2669 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_9 ();
 sg13g2_decap_8 FILLER_38_50 ();
 sg13g2_decap_8 FILLER_38_57 ();
 sg13g2_decap_8 FILLER_38_64 ();
 sg13g2_fill_2 FILLER_38_71 ();
 sg13g2_fill_1 FILLER_38_73 ();
 sg13g2_decap_8 FILLER_38_85 ();
 sg13g2_fill_2 FILLER_38_92 ();
 sg13g2_fill_2 FILLER_38_115 ();
 sg13g2_fill_1 FILLER_38_117 ();
 sg13g2_fill_2 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_173 ();
 sg13g2_fill_1 FILLER_38_180 ();
 sg13g2_fill_1 FILLER_38_209 ();
 sg13g2_fill_1 FILLER_38_218 ();
 sg13g2_fill_1 FILLER_38_231 ();
 sg13g2_decap_4 FILLER_38_242 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_fill_2 FILLER_38_257 ();
 sg13g2_fill_2 FILLER_38_267 ();
 sg13g2_fill_1 FILLER_38_281 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_296 ();
 sg13g2_fill_2 FILLER_38_369 ();
 sg13g2_fill_1 FILLER_38_378 ();
 sg13g2_fill_1 FILLER_38_397 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_fill_2 FILLER_38_414 ();
 sg13g2_fill_2 FILLER_38_421 ();
 sg13g2_fill_1 FILLER_38_433 ();
 sg13g2_fill_1 FILLER_38_495 ();
 sg13g2_fill_2 FILLER_38_584 ();
 sg13g2_fill_2 FILLER_38_638 ();
 sg13g2_fill_2 FILLER_38_648 ();
 sg13g2_fill_2 FILLER_38_660 ();
 sg13g2_fill_1 FILLER_38_680 ();
 sg13g2_fill_1 FILLER_38_712 ();
 sg13g2_fill_2 FILLER_38_717 ();
 sg13g2_fill_1 FILLER_38_727 ();
 sg13g2_fill_2 FILLER_38_732 ();
 sg13g2_fill_2 FILLER_38_742 ();
 sg13g2_fill_2 FILLER_38_755 ();
 sg13g2_fill_1 FILLER_38_762 ();
 sg13g2_decap_4 FILLER_38_810 ();
 sg13g2_fill_1 FILLER_38_814 ();
 sg13g2_fill_1 FILLER_38_833 ();
 sg13g2_fill_1 FILLER_38_839 ();
 sg13g2_fill_1 FILLER_38_850 ();
 sg13g2_fill_1 FILLER_38_870 ();
 sg13g2_fill_1 FILLER_38_906 ();
 sg13g2_fill_2 FILLER_38_986 ();
 sg13g2_fill_2 FILLER_38_1013 ();
 sg13g2_fill_2 FILLER_38_1023 ();
 sg13g2_fill_2 FILLER_38_1031 ();
 sg13g2_fill_1 FILLER_38_1041 ();
 sg13g2_fill_1 FILLER_38_1128 ();
 sg13g2_fill_2 FILLER_38_1141 ();
 sg13g2_fill_2 FILLER_38_1157 ();
 sg13g2_decap_4 FILLER_38_1194 ();
 sg13g2_fill_1 FILLER_38_1198 ();
 sg13g2_fill_2 FILLER_38_1279 ();
 sg13g2_fill_2 FILLER_38_1299 ();
 sg13g2_fill_1 FILLER_38_1316 ();
 sg13g2_fill_1 FILLER_38_1334 ();
 sg13g2_fill_1 FILLER_38_1358 ();
 sg13g2_fill_2 FILLER_38_1364 ();
 sg13g2_decap_4 FILLER_38_1375 ();
 sg13g2_fill_1 FILLER_38_1384 ();
 sg13g2_fill_2 FILLER_38_1412 ();
 sg13g2_fill_2 FILLER_38_1495 ();
 sg13g2_fill_2 FILLER_38_1502 ();
 sg13g2_fill_2 FILLER_38_1551 ();
 sg13g2_fill_1 FILLER_38_1559 ();
 sg13g2_fill_2 FILLER_38_1599 ();
 sg13g2_fill_1 FILLER_38_1620 ();
 sg13g2_fill_2 FILLER_38_1631 ();
 sg13g2_decap_8 FILLER_38_1652 ();
 sg13g2_fill_2 FILLER_38_1669 ();
 sg13g2_fill_1 FILLER_38_1671 ();
 sg13g2_decap_4 FILLER_38_1677 ();
 sg13g2_fill_1 FILLER_38_1681 ();
 sg13g2_decap_4 FILLER_38_1686 ();
 sg13g2_fill_1 FILLER_38_1690 ();
 sg13g2_fill_1 FILLER_38_1704 ();
 sg13g2_fill_2 FILLER_38_1731 ();
 sg13g2_fill_2 FILLER_38_1756 ();
 sg13g2_fill_2 FILLER_38_1784 ();
 sg13g2_fill_1 FILLER_38_1806 ();
 sg13g2_fill_1 FILLER_38_1821 ();
 sg13g2_fill_2 FILLER_38_1827 ();
 sg13g2_fill_1 FILLER_38_1866 ();
 sg13g2_fill_2 FILLER_38_1886 ();
 sg13g2_fill_2 FILLER_38_1905 ();
 sg13g2_fill_1 FILLER_38_1924 ();
 sg13g2_decap_8 FILLER_38_1961 ();
 sg13g2_decap_8 FILLER_38_1968 ();
 sg13g2_decap_4 FILLER_38_1975 ();
 sg13g2_fill_1 FILLER_38_1993 ();
 sg13g2_fill_1 FILLER_38_2008 ();
 sg13g2_fill_1 FILLER_38_2019 ();
 sg13g2_fill_2 FILLER_38_2093 ();
 sg13g2_fill_1 FILLER_38_2095 ();
 sg13g2_decap_8 FILLER_38_2136 ();
 sg13g2_fill_2 FILLER_38_2143 ();
 sg13g2_fill_2 FILLER_38_2212 ();
 sg13g2_decap_4 FILLER_38_2236 ();
 sg13g2_decap_4 FILLER_38_2244 ();
 sg13g2_fill_2 FILLER_38_2248 ();
 sg13g2_decap_8 FILLER_38_2286 ();
 sg13g2_decap_8 FILLER_38_2301 ();
 sg13g2_decap_8 FILLER_38_2308 ();
 sg13g2_fill_2 FILLER_38_2408 ();
 sg13g2_fill_2 FILLER_38_2455 ();
 sg13g2_fill_1 FILLER_38_2468 ();
 sg13g2_fill_1 FILLER_38_2535 ();
 sg13g2_decap_4 FILLER_38_2562 ();
 sg13g2_fill_1 FILLER_38_2571 ();
 sg13g2_decap_4 FILLER_38_2576 ();
 sg13g2_fill_2 FILLER_38_2580 ();
 sg13g2_decap_4 FILLER_38_2592 ();
 sg13g2_fill_1 FILLER_38_2596 ();
 sg13g2_decap_8 FILLER_38_2601 ();
 sg13g2_decap_8 FILLER_38_2608 ();
 sg13g2_fill_1 FILLER_38_2615 ();
 sg13g2_fill_2 FILLER_38_2626 ();
 sg13g2_decap_4 FILLER_38_2655 ();
 sg13g2_decap_8 FILLER_38_2662 ();
 sg13g2_fill_1 FILLER_38_2669 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_4 FILLER_39_14 ();
 sg13g2_fill_2 FILLER_39_22 ();
 sg13g2_fill_1 FILLER_39_24 ();
 sg13g2_decap_4 FILLER_39_63 ();
 sg13g2_fill_2 FILLER_39_67 ();
 sg13g2_fill_2 FILLER_39_75 ();
 sg13g2_fill_2 FILLER_39_155 ();
 sg13g2_decap_8 FILLER_39_183 ();
 sg13g2_fill_1 FILLER_39_196 ();
 sg13g2_fill_1 FILLER_39_207 ();
 sg13g2_fill_1 FILLER_39_234 ();
 sg13g2_fill_2 FILLER_39_241 ();
 sg13g2_fill_1 FILLER_39_261 ();
 sg13g2_fill_1 FILLER_39_268 ();
 sg13g2_fill_2 FILLER_39_280 ();
 sg13g2_fill_1 FILLER_39_297 ();
 sg13g2_fill_2 FILLER_39_347 ();
 sg13g2_fill_2 FILLER_39_377 ();
 sg13g2_fill_1 FILLER_39_382 ();
 sg13g2_fill_1 FILLER_39_388 ();
 sg13g2_fill_1 FILLER_39_423 ();
 sg13g2_fill_2 FILLER_39_455 ();
 sg13g2_fill_1 FILLER_39_465 ();
 sg13g2_fill_2 FILLER_39_532 ();
 sg13g2_fill_2 FILLER_39_543 ();
 sg13g2_fill_1 FILLER_39_563 ();
 sg13g2_fill_1 FILLER_39_568 ();
 sg13g2_fill_2 FILLER_39_582 ();
 sg13g2_fill_1 FILLER_39_589 ();
 sg13g2_fill_1 FILLER_39_603 ();
 sg13g2_fill_1 FILLER_39_617 ();
 sg13g2_fill_2 FILLER_39_629 ();
 sg13g2_fill_1 FILLER_39_649 ();
 sg13g2_fill_1 FILLER_39_660 ();
 sg13g2_fill_2 FILLER_39_668 ();
 sg13g2_fill_2 FILLER_39_688 ();
 sg13g2_fill_1 FILLER_39_690 ();
 sg13g2_fill_2 FILLER_39_721 ();
 sg13g2_fill_2 FILLER_39_773 ();
 sg13g2_fill_2 FILLER_39_779 ();
 sg13g2_fill_2 FILLER_39_807 ();
 sg13g2_fill_2 FILLER_39_819 ();
 sg13g2_fill_2 FILLER_39_847 ();
 sg13g2_fill_1 FILLER_39_849 ();
 sg13g2_fill_2 FILLER_39_855 ();
 sg13g2_fill_1 FILLER_39_857 ();
 sg13g2_fill_1 FILLER_39_862 ();
 sg13g2_fill_2 FILLER_39_868 ();
 sg13g2_fill_1 FILLER_39_881 ();
 sg13g2_decap_8 FILLER_39_898 ();
 sg13g2_fill_2 FILLER_39_909 ();
 sg13g2_fill_2 FILLER_39_916 ();
 sg13g2_fill_2 FILLER_39_945 ();
 sg13g2_fill_1 FILLER_39_957 ();
 sg13g2_fill_2 FILLER_39_962 ();
 sg13g2_fill_2 FILLER_39_981 ();
 sg13g2_fill_2 FILLER_39_1000 ();
 sg13g2_fill_1 FILLER_39_1054 ();
 sg13g2_fill_1 FILLER_39_1074 ();
 sg13g2_fill_1 FILLER_39_1104 ();
 sg13g2_fill_2 FILLER_39_1112 ();
 sg13g2_fill_1 FILLER_39_1127 ();
 sg13g2_fill_1 FILLER_39_1158 ();
 sg13g2_decap_4 FILLER_39_1231 ();
 sg13g2_fill_1 FILLER_39_1271 ();
 sg13g2_fill_1 FILLER_39_1288 ();
 sg13g2_fill_1 FILLER_39_1381 ();
 sg13g2_decap_4 FILLER_39_1407 ();
 sg13g2_fill_2 FILLER_39_1416 ();
 sg13g2_fill_1 FILLER_39_1418 ();
 sg13g2_fill_1 FILLER_39_1450 ();
 sg13g2_fill_2 FILLER_39_1467 ();
 sg13g2_fill_1 FILLER_39_1495 ();
 sg13g2_fill_1 FILLER_39_1505 ();
 sg13g2_fill_1 FILLER_39_1599 ();
 sg13g2_fill_1 FILLER_39_1608 ();
 sg13g2_fill_1 FILLER_39_1635 ();
 sg13g2_fill_1 FILLER_39_1662 ();
 sg13g2_fill_1 FILLER_39_1669 ();
 sg13g2_fill_1 FILLER_39_1675 ();
 sg13g2_fill_2 FILLER_39_1681 ();
 sg13g2_fill_2 FILLER_39_1722 ();
 sg13g2_fill_2 FILLER_39_1731 ();
 sg13g2_fill_2 FILLER_39_1759 ();
 sg13g2_fill_2 FILLER_39_1774 ();
 sg13g2_fill_1 FILLER_39_1776 ();
 sg13g2_fill_2 FILLER_39_1781 ();
 sg13g2_fill_2 FILLER_39_1791 ();
 sg13g2_decap_4 FILLER_39_1822 ();
 sg13g2_fill_1 FILLER_39_1826 ();
 sg13g2_fill_2 FILLER_39_1833 ();
 sg13g2_fill_2 FILLER_39_1846 ();
 sg13g2_fill_2 FILLER_39_1853 ();
 sg13g2_fill_1 FILLER_39_1855 ();
 sg13g2_fill_2 FILLER_39_1861 ();
 sg13g2_fill_1 FILLER_39_1863 ();
 sg13g2_decap_4 FILLER_39_1870 ();
 sg13g2_fill_1 FILLER_39_1874 ();
 sg13g2_fill_2 FILLER_39_1880 ();
 sg13g2_fill_1 FILLER_39_1882 ();
 sg13g2_decap_8 FILLER_39_1888 ();
 sg13g2_fill_2 FILLER_39_1905 ();
 sg13g2_fill_2 FILLER_39_1913 ();
 sg13g2_fill_1 FILLER_39_1915 ();
 sg13g2_fill_1 FILLER_39_1921 ();
 sg13g2_fill_2 FILLER_39_1927 ();
 sg13g2_fill_2 FILLER_39_1933 ();
 sg13g2_fill_2 FILLER_39_1940 ();
 sg13g2_decap_8 FILLER_39_1968 ();
 sg13g2_decap_8 FILLER_39_1975 ();
 sg13g2_decap_4 FILLER_39_1982 ();
 sg13g2_fill_2 FILLER_39_1986 ();
 sg13g2_decap_8 FILLER_39_1992 ();
 sg13g2_fill_2 FILLER_39_1999 ();
 sg13g2_fill_1 FILLER_39_2016 ();
 sg13g2_fill_2 FILLER_39_2059 ();
 sg13g2_fill_1 FILLER_39_2061 ();
 sg13g2_fill_2 FILLER_39_2072 ();
 sg13g2_fill_2 FILLER_39_2087 ();
 sg13g2_fill_1 FILLER_39_2161 ();
 sg13g2_fill_2 FILLER_39_2198 ();
 sg13g2_fill_1 FILLER_39_2200 ();
 sg13g2_fill_2 FILLER_39_2283 ();
 sg13g2_fill_1 FILLER_39_2285 ();
 sg13g2_fill_1 FILLER_39_2325 ();
 sg13g2_fill_2 FILLER_39_2339 ();
 sg13g2_fill_2 FILLER_39_2386 ();
 sg13g2_fill_1 FILLER_39_2401 ();
 sg13g2_fill_1 FILLER_39_2489 ();
 sg13g2_fill_1 FILLER_39_2506 ();
 sg13g2_fill_2 FILLER_39_2542 ();
 sg13g2_fill_2 FILLER_39_2548 ();
 sg13g2_fill_1 FILLER_39_2550 ();
 sg13g2_decap_4 FILLER_39_2571 ();
 sg13g2_fill_1 FILLER_39_2575 ();
 sg13g2_fill_2 FILLER_39_2616 ();
 sg13g2_fill_1 FILLER_39_2618 ();
 sg13g2_fill_2 FILLER_39_2668 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_4 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_11 ();
 sg13g2_fill_2 FILLER_40_58 ();
 sg13g2_fill_2 FILLER_40_76 ();
 sg13g2_decap_4 FILLER_40_86 ();
 sg13g2_decap_4 FILLER_40_95 ();
 sg13g2_decap_4 FILLER_40_103 ();
 sg13g2_decap_8 FILLER_40_150 ();
 sg13g2_decap_4 FILLER_40_157 ();
 sg13g2_fill_2 FILLER_40_161 ();
 sg13g2_decap_4 FILLER_40_171 ();
 sg13g2_fill_2 FILLER_40_175 ();
 sg13g2_fill_2 FILLER_40_185 ();
 sg13g2_fill_1 FILLER_40_187 ();
 sg13g2_decap_4 FILLER_40_200 ();
 sg13g2_decap_4 FILLER_40_212 ();
 sg13g2_fill_1 FILLER_40_216 ();
 sg13g2_decap_4 FILLER_40_221 ();
 sg13g2_fill_1 FILLER_40_225 ();
 sg13g2_fill_1 FILLER_40_261 ();
 sg13g2_fill_1 FILLER_40_311 ();
 sg13g2_fill_2 FILLER_40_316 ();
 sg13g2_fill_2 FILLER_40_373 ();
 sg13g2_fill_2 FILLER_40_382 ();
 sg13g2_fill_2 FILLER_40_388 ();
 sg13g2_fill_1 FILLER_40_437 ();
 sg13g2_fill_2 FILLER_40_452 ();
 sg13g2_fill_1 FILLER_40_470 ();
 sg13g2_fill_2 FILLER_40_476 ();
 sg13g2_fill_1 FILLER_40_503 ();
 sg13g2_fill_1 FILLER_40_519 ();
 sg13g2_decap_8 FILLER_40_524 ();
 sg13g2_decap_8 FILLER_40_531 ();
 sg13g2_fill_2 FILLER_40_538 ();
 sg13g2_fill_1 FILLER_40_540 ();
 sg13g2_fill_1 FILLER_40_555 ();
 sg13g2_fill_1 FILLER_40_580 ();
 sg13g2_fill_1 FILLER_40_604 ();
 sg13g2_fill_1 FILLER_40_610 ();
 sg13g2_fill_1 FILLER_40_639 ();
 sg13g2_fill_1 FILLER_40_659 ();
 sg13g2_fill_1 FILLER_40_684 ();
 sg13g2_fill_1 FILLER_40_713 ();
 sg13g2_decap_8 FILLER_40_760 ();
 sg13g2_decap_4 FILLER_40_791 ();
 sg13g2_fill_2 FILLER_40_795 ();
 sg13g2_decap_4 FILLER_40_806 ();
 sg13g2_fill_1 FILLER_40_846 ();
 sg13g2_fill_2 FILLER_40_873 ();
 sg13g2_fill_2 FILLER_40_891 ();
 sg13g2_fill_1 FILLER_40_922 ();
 sg13g2_decap_4 FILLER_40_938 ();
 sg13g2_decap_4 FILLER_40_949 ();
 sg13g2_fill_2 FILLER_40_953 ();
 sg13g2_decap_4 FILLER_40_980 ();
 sg13g2_fill_1 FILLER_40_984 ();
 sg13g2_fill_2 FILLER_40_990 ();
 sg13g2_fill_1 FILLER_40_997 ();
 sg13g2_fill_2 FILLER_40_1005 ();
 sg13g2_fill_1 FILLER_40_1019 ();
 sg13g2_fill_1 FILLER_40_1028 ();
 sg13g2_fill_2 FILLER_40_1033 ();
 sg13g2_fill_1 FILLER_40_1045 ();
 sg13g2_fill_1 FILLER_40_1082 ();
 sg13g2_fill_1 FILLER_40_1088 ();
 sg13g2_fill_1 FILLER_40_1105 ();
 sg13g2_fill_2 FILLER_40_1110 ();
 sg13g2_decap_8 FILLER_40_1168 ();
 sg13g2_decap_8 FILLER_40_1175 ();
 sg13g2_decap_8 FILLER_40_1182 ();
 sg13g2_decap_4 FILLER_40_1199 ();
 sg13g2_fill_2 FILLER_40_1220 ();
 sg13g2_decap_8 FILLER_40_1234 ();
 sg13g2_decap_4 FILLER_40_1241 ();
 sg13g2_fill_1 FILLER_40_1245 ();
 sg13g2_fill_1 FILLER_40_1255 ();
 sg13g2_fill_1 FILLER_40_1267 ();
 sg13g2_fill_2 FILLER_40_1321 ();
 sg13g2_fill_1 FILLER_40_1329 ();
 sg13g2_fill_2 FILLER_40_1351 ();
 sg13g2_fill_1 FILLER_40_1380 ();
 sg13g2_fill_2 FILLER_40_1392 ();
 sg13g2_fill_1 FILLER_40_1402 ();
 sg13g2_decap_4 FILLER_40_1428 ();
 sg13g2_decap_4 FILLER_40_1437 ();
 sg13g2_fill_1 FILLER_40_1462 ();
 sg13g2_fill_1 FILLER_40_1485 ();
 sg13g2_fill_1 FILLER_40_1491 ();
 sg13g2_fill_1 FILLER_40_1497 ();
 sg13g2_fill_1 FILLER_40_1541 ();
 sg13g2_fill_2 FILLER_40_1551 ();
 sg13g2_fill_1 FILLER_40_1587 ();
 sg13g2_fill_2 FILLER_40_1595 ();
 sg13g2_fill_2 FILLER_40_1619 ();
 sg13g2_fill_2 FILLER_40_1626 ();
 sg13g2_fill_2 FILLER_40_1691 ();
 sg13g2_fill_1 FILLER_40_1693 ();
 sg13g2_fill_2 FILLER_40_1711 ();
 sg13g2_fill_1 FILLER_40_1713 ();
 sg13g2_decap_8 FILLER_40_1723 ();
 sg13g2_fill_2 FILLER_40_1730 ();
 sg13g2_fill_1 FILLER_40_1732 ();
 sg13g2_decap_8 FILLER_40_1762 ();
 sg13g2_decap_8 FILLER_40_1769 ();
 sg13g2_decap_8 FILLER_40_1776 ();
 sg13g2_fill_2 FILLER_40_1783 ();
 sg13g2_fill_1 FILLER_40_1785 ();
 sg13g2_decap_8 FILLER_40_1815 ();
 sg13g2_decap_8 FILLER_40_1822 ();
 sg13g2_decap_8 FILLER_40_1829 ();
 sg13g2_decap_8 FILLER_40_1836 ();
 sg13g2_decap_8 FILLER_40_1843 ();
 sg13g2_decap_8 FILLER_40_1850 ();
 sg13g2_decap_8 FILLER_40_1857 ();
 sg13g2_decap_8 FILLER_40_1864 ();
 sg13g2_decap_8 FILLER_40_1871 ();
 sg13g2_decap_4 FILLER_40_1878 ();
 sg13g2_decap_8 FILLER_40_1886 ();
 sg13g2_fill_1 FILLER_40_1928 ();
 sg13g2_decap_8 FILLER_40_1938 ();
 sg13g2_decap_8 FILLER_40_1945 ();
 sg13g2_decap_8 FILLER_40_1952 ();
 sg13g2_decap_4 FILLER_40_1959 ();
 sg13g2_fill_1 FILLER_40_1963 ();
 sg13g2_decap_8 FILLER_40_2000 ();
 sg13g2_fill_1 FILLER_40_2007 ();
 sg13g2_fill_2 FILLER_40_2027 ();
 sg13g2_fill_1 FILLER_40_2029 ();
 sg13g2_decap_8 FILLER_40_2034 ();
 sg13g2_decap_8 FILLER_40_2041 ();
 sg13g2_decap_4 FILLER_40_2048 ();
 sg13g2_fill_1 FILLER_40_2052 ();
 sg13g2_fill_1 FILLER_40_2057 ();
 sg13g2_decap_4 FILLER_40_2063 ();
 sg13g2_fill_1 FILLER_40_2067 ();
 sg13g2_decap_4 FILLER_40_2090 ();
 sg13g2_fill_2 FILLER_40_2094 ();
 sg13g2_decap_8 FILLER_40_2100 ();
 sg13g2_fill_1 FILLER_40_2107 ();
 sg13g2_fill_2 FILLER_40_2139 ();
 sg13g2_decap_4 FILLER_40_2145 ();
 sg13g2_fill_2 FILLER_40_2149 ();
 sg13g2_decap_4 FILLER_40_2161 ();
 sg13g2_fill_1 FILLER_40_2165 ();
 sg13g2_fill_2 FILLER_40_2192 ();
 sg13g2_decap_4 FILLER_40_2220 ();
 sg13g2_fill_2 FILLER_40_2224 ();
 sg13g2_fill_2 FILLER_40_2255 ();
 sg13g2_decap_4 FILLER_40_2267 ();
 sg13g2_fill_1 FILLER_40_2271 ();
 sg13g2_fill_2 FILLER_40_2347 ();
 sg13g2_fill_2 FILLER_40_2377 ();
 sg13g2_fill_2 FILLER_40_2487 ();
 sg13g2_fill_2 FILLER_40_2559 ();
 sg13g2_fill_1 FILLER_40_2561 ();
 sg13g2_fill_2 FILLER_40_2625 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_9 ();
 sg13g2_fill_1 FILLER_41_69 ();
 sg13g2_fill_1 FILLER_41_76 ();
 sg13g2_fill_1 FILLER_41_85 ();
 sg13g2_fill_2 FILLER_41_94 ();
 sg13g2_decap_8 FILLER_41_101 ();
 sg13g2_fill_1 FILLER_41_108 ();
 sg13g2_decap_8 FILLER_41_115 ();
 sg13g2_fill_2 FILLER_41_122 ();
 sg13g2_decap_8 FILLER_41_129 ();
 sg13g2_decap_4 FILLER_41_136 ();
 sg13g2_fill_1 FILLER_41_140 ();
 sg13g2_decap_4 FILLER_41_156 ();
 sg13g2_fill_1 FILLER_41_177 ();
 sg13g2_fill_1 FILLER_41_186 ();
 sg13g2_fill_2 FILLER_41_200 ();
 sg13g2_fill_1 FILLER_41_202 ();
 sg13g2_decap_8 FILLER_41_208 ();
 sg13g2_decap_8 FILLER_41_215 ();
 sg13g2_fill_2 FILLER_41_227 ();
 sg13g2_fill_1 FILLER_41_229 ();
 sg13g2_fill_1 FILLER_41_268 ();
 sg13g2_fill_1 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_317 ();
 sg13g2_fill_2 FILLER_41_332 ();
 sg13g2_fill_1 FILLER_41_360 ();
 sg13g2_fill_1 FILLER_41_373 ();
 sg13g2_fill_2 FILLER_41_418 ();
 sg13g2_fill_2 FILLER_41_464 ();
 sg13g2_fill_1 FILLER_41_466 ();
 sg13g2_fill_1 FILLER_41_475 ();
 sg13g2_fill_2 FILLER_41_493 ();
 sg13g2_decap_8 FILLER_41_515 ();
 sg13g2_decap_4 FILLER_41_522 ();
 sg13g2_decap_8 FILLER_41_530 ();
 sg13g2_decap_4 FILLER_41_537 ();
 sg13g2_fill_1 FILLER_41_549 ();
 sg13g2_fill_2 FILLER_41_598 ();
 sg13g2_fill_1 FILLER_41_612 ();
 sg13g2_fill_1 FILLER_41_620 ();
 sg13g2_fill_2 FILLER_41_631 ();
 sg13g2_fill_1 FILLER_41_695 ();
 sg13g2_decap_8 FILLER_41_706 ();
 sg13g2_fill_1 FILLER_41_728 ();
 sg13g2_fill_1 FILLER_41_750 ();
 sg13g2_decap_8 FILLER_41_760 ();
 sg13g2_fill_2 FILLER_41_767 ();
 sg13g2_fill_1 FILLER_41_795 ();
 sg13g2_fill_1 FILLER_41_817 ();
 sg13g2_decap_4 FILLER_41_869 ();
 sg13g2_fill_2 FILLER_41_873 ();
 sg13g2_fill_2 FILLER_41_889 ();
 sg13g2_fill_1 FILLER_41_891 ();
 sg13g2_fill_2 FILLER_41_902 ();
 sg13g2_fill_1 FILLER_41_923 ();
 sg13g2_decap_4 FILLER_41_950 ();
 sg13g2_decap_8 FILLER_41_959 ();
 sg13g2_fill_1 FILLER_41_966 ();
 sg13g2_decap_8 FILLER_41_992 ();
 sg13g2_fill_2 FILLER_41_999 ();
 sg13g2_fill_2 FILLER_41_1006 ();
 sg13g2_fill_1 FILLER_41_1008 ();
 sg13g2_fill_2 FILLER_41_1014 ();
 sg13g2_fill_2 FILLER_41_1063 ();
 sg13g2_fill_1 FILLER_41_1065 ();
 sg13g2_fill_2 FILLER_41_1092 ();
 sg13g2_fill_2 FILLER_41_1118 ();
 sg13g2_fill_1 FILLER_41_1130 ();
 sg13g2_decap_8 FILLER_41_1176 ();
 sg13g2_decap_8 FILLER_41_1183 ();
 sg13g2_decap_8 FILLER_41_1190 ();
 sg13g2_fill_2 FILLER_41_1207 ();
 sg13g2_fill_1 FILLER_41_1209 ();
 sg13g2_fill_2 FILLER_41_1214 ();
 sg13g2_decap_8 FILLER_41_1229 ();
 sg13g2_decap_4 FILLER_41_1236 ();
 sg13g2_fill_2 FILLER_41_1244 ();
 sg13g2_fill_1 FILLER_41_1261 ();
 sg13g2_fill_1 FILLER_41_1268 ();
 sg13g2_fill_1 FILLER_41_1273 ();
 sg13g2_fill_1 FILLER_41_1310 ();
 sg13g2_fill_1 FILLER_41_1332 ();
 sg13g2_fill_1 FILLER_41_1355 ();
 sg13g2_fill_2 FILLER_41_1363 ();
 sg13g2_fill_1 FILLER_41_1372 ();
 sg13g2_fill_1 FILLER_41_1378 ();
 sg13g2_fill_2 FILLER_41_1384 ();
 sg13g2_fill_1 FILLER_41_1386 ();
 sg13g2_fill_2 FILLER_41_1394 ();
 sg13g2_decap_4 FILLER_41_1423 ();
 sg13g2_fill_1 FILLER_41_1427 ();
 sg13g2_fill_2 FILLER_41_1432 ();
 sg13g2_fill_2 FILLER_41_1439 ();
 sg13g2_fill_1 FILLER_41_1455 ();
 sg13g2_fill_1 FILLER_41_1465 ();
 sg13g2_fill_1 FILLER_41_1471 ();
 sg13g2_fill_2 FILLER_41_1495 ();
 sg13g2_fill_1 FILLER_41_1553 ();
 sg13g2_fill_1 FILLER_41_1561 ();
 sg13g2_fill_1 FILLER_41_1574 ();
 sg13g2_fill_2 FILLER_41_1593 ();
 sg13g2_fill_2 FILLER_41_1607 ();
 sg13g2_fill_2 FILLER_41_1618 ();
 sg13g2_fill_1 FILLER_41_1636 ();
 sg13g2_fill_2 FILLER_41_1642 ();
 sg13g2_fill_1 FILLER_41_1652 ();
 sg13g2_decap_8 FILLER_41_1658 ();
 sg13g2_fill_2 FILLER_41_1665 ();
 sg13g2_decap_8 FILLER_41_1677 ();
 sg13g2_fill_1 FILLER_41_1694 ();
 sg13g2_decap_8 FILLER_41_1722 ();
 sg13g2_decap_8 FILLER_41_1729 ();
 sg13g2_decap_4 FILLER_41_1740 ();
 sg13g2_decap_8 FILLER_41_1774 ();
 sg13g2_decap_8 FILLER_41_1781 ();
 sg13g2_fill_2 FILLER_41_1793 ();
 sg13g2_fill_1 FILLER_41_1795 ();
 sg13g2_fill_2 FILLER_41_1832 ();
 sg13g2_decap_4 FILLER_41_1860 ();
 sg13g2_fill_1 FILLER_41_1864 ();
 sg13g2_fill_1 FILLER_41_1869 ();
 sg13g2_decap_4 FILLER_41_1877 ();
 sg13g2_fill_2 FILLER_41_1881 ();
 sg13g2_fill_1 FILLER_41_1888 ();
 sg13g2_fill_1 FILLER_41_1915 ();
 sg13g2_fill_1 FILLER_41_1929 ();
 sg13g2_decap_4 FILLER_41_1968 ();
 sg13g2_fill_1 FILLER_41_1972 ();
 sg13g2_fill_2 FILLER_41_2009 ();
 sg13g2_fill_1 FILLER_41_2017 ();
 sg13g2_decap_4 FILLER_41_2048 ();
 sg13g2_fill_2 FILLER_41_2052 ();
 sg13g2_decap_8 FILLER_41_2090 ();
 sg13g2_decap_8 FILLER_41_2097 ();
 sg13g2_decap_8 FILLER_41_2104 ();
 sg13g2_fill_1 FILLER_41_2111 ();
 sg13g2_decap_8 FILLER_41_2139 ();
 sg13g2_fill_2 FILLER_41_2146 ();
 sg13g2_fill_2 FILLER_41_2178 ();
 sg13g2_decap_8 FILLER_41_2205 ();
 sg13g2_decap_8 FILLER_41_2212 ();
 sg13g2_decap_8 FILLER_41_2219 ();
 sg13g2_fill_2 FILLER_41_2240 ();
 sg13g2_fill_2 FILLER_41_2263 ();
 sg13g2_fill_1 FILLER_41_2280 ();
 sg13g2_fill_1 FILLER_41_2314 ();
 sg13g2_fill_1 FILLER_41_2322 ();
 sg13g2_fill_1 FILLER_41_2366 ();
 sg13g2_fill_1 FILLER_41_2387 ();
 sg13g2_decap_4 FILLER_41_2401 ();
 sg13g2_fill_1 FILLER_41_2405 ();
 sg13g2_fill_2 FILLER_41_2445 ();
 sg13g2_fill_1 FILLER_41_2462 ();
 sg13g2_fill_1 FILLER_41_2499 ();
 sg13g2_fill_1 FILLER_41_2507 ();
 sg13g2_fill_2 FILLER_41_2537 ();
 sg13g2_decap_4 FILLER_41_2546 ();
 sg13g2_fill_2 FILLER_41_2550 ();
 sg13g2_fill_2 FILLER_41_2578 ();
 sg13g2_fill_1 FILLER_41_2612 ();
 sg13g2_fill_1 FILLER_41_2623 ();
 sg13g2_fill_1 FILLER_41_2628 ();
 sg13g2_fill_2 FILLER_41_2638 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_34 ();
 sg13g2_fill_1 FILLER_42_36 ();
 sg13g2_decap_8 FILLER_42_47 ();
 sg13g2_decap_4 FILLER_42_60 ();
 sg13g2_fill_1 FILLER_42_69 ();
 sg13g2_fill_1 FILLER_42_76 ();
 sg13g2_fill_1 FILLER_42_82 ();
 sg13g2_fill_1 FILLER_42_89 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_fill_1 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_114 ();
 sg13g2_fill_1 FILLER_42_121 ();
 sg13g2_decap_8 FILLER_42_127 ();
 sg13g2_fill_2 FILLER_42_134 ();
 sg13g2_fill_1 FILLER_42_174 ();
 sg13g2_fill_1 FILLER_42_201 ();
 sg13g2_decap_8 FILLER_42_219 ();
 sg13g2_fill_2 FILLER_42_226 ();
 sg13g2_fill_1 FILLER_42_239 ();
 sg13g2_decap_4 FILLER_42_244 ();
 sg13g2_fill_1 FILLER_42_261 ();
 sg13g2_decap_8 FILLER_42_282 ();
 sg13g2_fill_2 FILLER_42_293 ();
 sg13g2_decap_8 FILLER_42_300 ();
 sg13g2_decap_8 FILLER_42_307 ();
 sg13g2_decap_4 FILLER_42_314 ();
 sg13g2_decap_4 FILLER_42_328 ();
 sg13g2_fill_2 FILLER_42_336 ();
 sg13g2_fill_1 FILLER_42_338 ();
 sg13g2_fill_2 FILLER_42_360 ();
 sg13g2_fill_1 FILLER_42_380 ();
 sg13g2_fill_1 FILLER_42_401 ();
 sg13g2_fill_2 FILLER_42_427 ();
 sg13g2_fill_2 FILLER_42_438 ();
 sg13g2_fill_1 FILLER_42_440 ();
 sg13g2_fill_2 FILLER_42_501 ();
 sg13g2_fill_2 FILLER_42_511 ();
 sg13g2_fill_2 FILLER_42_547 ();
 sg13g2_decap_8 FILLER_42_566 ();
 sg13g2_decap_8 FILLER_42_592 ();
 sg13g2_decap_8 FILLER_42_599 ();
 sg13g2_fill_2 FILLER_42_606 ();
 sg13g2_fill_1 FILLER_42_608 ();
 sg13g2_fill_1 FILLER_42_634 ();
 sg13g2_fill_1 FILLER_42_676 ();
 sg13g2_fill_1 FILLER_42_689 ();
 sg13g2_fill_2 FILLER_42_700 ();
 sg13g2_fill_1 FILLER_42_702 ();
 sg13g2_decap_8 FILLER_42_711 ();
 sg13g2_decap_4 FILLER_42_718 ();
 sg13g2_fill_1 FILLER_42_722 ();
 sg13g2_decap_4 FILLER_42_735 ();
 sg13g2_fill_1 FILLER_42_739 ();
 sg13g2_fill_1 FILLER_42_766 ();
 sg13g2_fill_1 FILLER_42_777 ();
 sg13g2_fill_1 FILLER_42_808 ();
 sg13g2_decap_8 FILLER_42_839 ();
 sg13g2_decap_4 FILLER_42_846 ();
 sg13g2_fill_2 FILLER_42_881 ();
 sg13g2_fill_2 FILLER_42_887 ();
 sg13g2_decap_8 FILLER_42_919 ();
 sg13g2_fill_1 FILLER_42_926 ();
 sg13g2_decap_8 FILLER_42_934 ();
 sg13g2_decap_4 FILLER_42_941 ();
 sg13g2_fill_1 FILLER_42_945 ();
 sg13g2_decap_8 FILLER_42_951 ();
 sg13g2_decap_4 FILLER_42_958 ();
 sg13g2_fill_1 FILLER_42_975 ();
 sg13g2_fill_2 FILLER_42_992 ();
 sg13g2_fill_2 FILLER_42_1018 ();
 sg13g2_fill_2 FILLER_42_1040 ();
 sg13g2_fill_1 FILLER_42_1042 ();
 sg13g2_fill_1 FILLER_42_1052 ();
 sg13g2_decap_4 FILLER_42_1061 ();
 sg13g2_fill_1 FILLER_42_1065 ();
 sg13g2_decap_8 FILLER_42_1070 ();
 sg13g2_fill_1 FILLER_42_1077 ();
 sg13g2_decap_4 FILLER_42_1097 ();
 sg13g2_decap_4 FILLER_42_1160 ();
 sg13g2_fill_2 FILLER_42_1164 ();
 sg13g2_fill_1 FILLER_42_1225 ();
 sg13g2_decap_8 FILLER_42_1230 ();
 sg13g2_decap_8 FILLER_42_1237 ();
 sg13g2_decap_4 FILLER_42_1244 ();
 sg13g2_fill_1 FILLER_42_1248 ();
 sg13g2_decap_8 FILLER_42_1252 ();
 sg13g2_fill_2 FILLER_42_1259 ();
 sg13g2_fill_1 FILLER_42_1261 ();
 sg13g2_decap_8 FILLER_42_1266 ();
 sg13g2_fill_1 FILLER_42_1273 ();
 sg13g2_fill_2 FILLER_42_1291 ();
 sg13g2_fill_1 FILLER_42_1313 ();
 sg13g2_fill_2 FILLER_42_1338 ();
 sg13g2_fill_1 FILLER_42_1351 ();
 sg13g2_fill_1 FILLER_42_1360 ();
 sg13g2_fill_2 FILLER_42_1365 ();
 sg13g2_fill_2 FILLER_42_1377 ();
 sg13g2_fill_2 FILLER_42_1382 ();
 sg13g2_fill_1 FILLER_42_1391 ();
 sg13g2_fill_2 FILLER_42_1397 ();
 sg13g2_decap_4 FILLER_42_1420 ();
 sg13g2_fill_1 FILLER_42_1449 ();
 sg13g2_fill_1 FILLER_42_1457 ();
 sg13g2_fill_2 FILLER_42_1468 ();
 sg13g2_fill_1 FILLER_42_1502 ();
 sg13g2_fill_2 FILLER_42_1511 ();
 sg13g2_fill_1 FILLER_42_1513 ();
 sg13g2_fill_2 FILLER_42_1557 ();
 sg13g2_fill_2 FILLER_42_1571 ();
 sg13g2_fill_1 FILLER_42_1593 ();
 sg13g2_decap_4 FILLER_42_1649 ();
 sg13g2_fill_1 FILLER_42_1658 ();
 sg13g2_decap_8 FILLER_42_1662 ();
 sg13g2_fill_1 FILLER_42_1702 ();
 sg13g2_fill_2 FILLER_42_1712 ();
 sg13g2_decap_4 FILLER_42_1718 ();
 sg13g2_fill_1 FILLER_42_1722 ();
 sg13g2_fill_2 FILLER_42_1735 ();
 sg13g2_fill_1 FILLER_42_1737 ();
 sg13g2_fill_1 FILLER_42_1746 ();
 sg13g2_fill_2 FILLER_42_1753 ();
 sg13g2_fill_1 FILLER_42_1755 ();
 sg13g2_fill_2 FILLER_42_1812 ();
 sg13g2_fill_1 FILLER_42_1814 ();
 sg13g2_fill_2 FILLER_42_1851 ();
 sg13g2_fill_1 FILLER_42_1853 ();
 sg13g2_fill_1 FILLER_42_1885 ();
 sg13g2_decap_4 FILLER_42_1891 ();
 sg13g2_fill_2 FILLER_42_1895 ();
 sg13g2_fill_2 FILLER_42_1905 ();
 sg13g2_fill_1 FILLER_42_1907 ();
 sg13g2_decap_4 FILLER_42_1921 ();
 sg13g2_fill_2 FILLER_42_1925 ();
 sg13g2_fill_1 FILLER_42_1956 ();
 sg13g2_decap_8 FILLER_42_2038 ();
 sg13g2_decap_8 FILLER_42_2045 ();
 sg13g2_fill_1 FILLER_42_2052 ();
 sg13g2_fill_1 FILLER_42_2079 ();
 sg13g2_fill_2 FILLER_42_2116 ();
 sg13g2_fill_2 FILLER_42_2152 ();
 sg13g2_decap_8 FILLER_42_2158 ();
 sg13g2_decap_8 FILLER_42_2165 ();
 sg13g2_decap_4 FILLER_42_2172 ();
 sg13g2_fill_2 FILLER_42_2176 ();
 sg13g2_decap_8 FILLER_42_2199 ();
 sg13g2_decap_8 FILLER_42_2206 ();
 sg13g2_decap_8 FILLER_42_2213 ();
 sg13g2_decap_8 FILLER_42_2220 ();
 sg13g2_fill_1 FILLER_42_2227 ();
 sg13g2_fill_2 FILLER_42_2232 ();
 sg13g2_fill_1 FILLER_42_2278 ();
 sg13g2_fill_2 FILLER_42_2312 ();
 sg13g2_fill_1 FILLER_42_2314 ();
 sg13g2_fill_1 FILLER_42_2322 ();
 sg13g2_fill_2 FILLER_42_2326 ();
 sg13g2_fill_2 FILLER_42_2341 ();
 sg13g2_fill_2 FILLER_42_2355 ();
 sg13g2_fill_2 FILLER_42_2451 ();
 sg13g2_fill_2 FILLER_42_2505 ();
 sg13g2_fill_2 FILLER_42_2554 ();
 sg13g2_fill_1 FILLER_42_2573 ();
 sg13g2_fill_2 FILLER_42_2609 ();
 sg13g2_fill_1 FILLER_42_2611 ();
 sg13g2_fill_2 FILLER_42_2615 ();
 sg13g2_fill_2 FILLER_42_2620 ();
 sg13g2_fill_1 FILLER_42_2641 ();
 sg13g2_fill_2 FILLER_42_2668 ();
 sg13g2_fill_2 FILLER_43_10 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_4 FILLER_43_49 ();
 sg13g2_fill_2 FILLER_43_53 ();
 sg13g2_fill_1 FILLER_43_61 ();
 sg13g2_fill_1 FILLER_43_87 ();
 sg13g2_fill_2 FILLER_43_131 ();
 sg13g2_decap_4 FILLER_43_137 ();
 sg13g2_fill_1 FILLER_43_141 ();
 sg13g2_fill_2 FILLER_43_159 ();
 sg13g2_fill_2 FILLER_43_166 ();
 sg13g2_fill_1 FILLER_43_168 ();
 sg13g2_decap_4 FILLER_43_181 ();
 sg13g2_fill_2 FILLER_43_185 ();
 sg13g2_decap_4 FILLER_43_193 ();
 sg13g2_fill_1 FILLER_43_197 ();
 sg13g2_fill_2 FILLER_43_211 ();
 sg13g2_fill_1 FILLER_43_213 ();
 sg13g2_fill_2 FILLER_43_228 ();
 sg13g2_fill_2 FILLER_43_248 ();
 sg13g2_decap_8 FILLER_43_302 ();
 sg13g2_fill_2 FILLER_43_313 ();
 sg13g2_fill_2 FILLER_43_324 ();
 sg13g2_fill_1 FILLER_43_326 ();
 sg13g2_fill_2 FILLER_43_331 ();
 sg13g2_decap_4 FILLER_43_337 ();
 sg13g2_fill_1 FILLER_43_341 ();
 sg13g2_fill_1 FILLER_43_352 ();
 sg13g2_fill_1 FILLER_43_366 ();
 sg13g2_fill_1 FILLER_43_379 ();
 sg13g2_fill_1 FILLER_43_384 ();
 sg13g2_decap_4 FILLER_43_396 ();
 sg13g2_fill_2 FILLER_43_400 ();
 sg13g2_decap_4 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_413 ();
 sg13g2_fill_1 FILLER_43_427 ();
 sg13g2_fill_1 FILLER_43_449 ();
 sg13g2_decap_4 FILLER_43_476 ();
 sg13g2_fill_2 FILLER_43_480 ();
 sg13g2_fill_2 FILLER_43_507 ();
 sg13g2_fill_1 FILLER_43_514 ();
 sg13g2_fill_1 FILLER_43_519 ();
 sg13g2_fill_1 FILLER_43_530 ();
 sg13g2_fill_1 FILLER_43_536 ();
 sg13g2_fill_1 FILLER_43_554 ();
 sg13g2_fill_2 FILLER_43_570 ();
 sg13g2_fill_1 FILLER_43_579 ();
 sg13g2_fill_2 FILLER_43_652 ();
 sg13g2_fill_1 FILLER_43_695 ();
 sg13g2_fill_2 FILLER_43_722 ();
 sg13g2_fill_1 FILLER_43_724 ();
 sg13g2_decap_4 FILLER_43_737 ();
 sg13g2_fill_2 FILLER_43_741 ();
 sg13g2_decap_8 FILLER_43_747 ();
 sg13g2_fill_2 FILLER_43_754 ();
 sg13g2_fill_2 FILLER_43_761 ();
 sg13g2_fill_1 FILLER_43_763 ();
 sg13g2_fill_2 FILLER_43_789 ();
 sg13g2_fill_1 FILLER_43_791 ();
 sg13g2_fill_2 FILLER_43_828 ();
 sg13g2_fill_2 FILLER_43_834 ();
 sg13g2_fill_1 FILLER_43_836 ();
 sg13g2_fill_2 FILLER_43_842 ();
 sg13g2_fill_1 FILLER_43_844 ();
 sg13g2_fill_2 FILLER_43_849 ();
 sg13g2_fill_1 FILLER_43_855 ();
 sg13g2_decap_8 FILLER_43_957 ();
 sg13g2_fill_1 FILLER_43_998 ();
 sg13g2_decap_4 FILLER_43_1025 ();
 sg13g2_fill_1 FILLER_43_1029 ();
 sg13g2_decap_4 FILLER_43_1035 ();
 sg13g2_fill_2 FILLER_43_1049 ();
 sg13g2_fill_1 FILLER_43_1051 ();
 sg13g2_fill_2 FILLER_43_1057 ();
 sg13g2_fill_1 FILLER_43_1059 ();
 sg13g2_decap_4 FILLER_43_1078 ();
 sg13g2_fill_2 FILLER_43_1082 ();
 sg13g2_decap_8 FILLER_43_1088 ();
 sg13g2_fill_1 FILLER_43_1095 ();
 sg13g2_fill_2 FILLER_43_1182 ();
 sg13g2_fill_1 FILLER_43_1184 ();
 sg13g2_fill_1 FILLER_43_1211 ();
 sg13g2_fill_2 FILLER_43_1238 ();
 sg13g2_fill_1 FILLER_43_1240 ();
 sg13g2_fill_2 FILLER_43_1273 ();
 sg13g2_fill_1 FILLER_43_1285 ();
 sg13g2_fill_1 FILLER_43_1311 ();
 sg13g2_fill_2 FILLER_43_1317 ();
 sg13g2_fill_2 FILLER_43_1327 ();
 sg13g2_decap_4 FILLER_43_1343 ();
 sg13g2_decap_8 FILLER_43_1354 ();
 sg13g2_fill_2 FILLER_43_1361 ();
 sg13g2_fill_1 FILLER_43_1363 ();
 sg13g2_fill_2 FILLER_43_1377 ();
 sg13g2_fill_1 FILLER_43_1379 ();
 sg13g2_fill_2 FILLER_43_1385 ();
 sg13g2_fill_1 FILLER_43_1387 ();
 sg13g2_fill_2 FILLER_43_1395 ();
 sg13g2_fill_1 FILLER_43_1397 ();
 sg13g2_decap_8 FILLER_43_1403 ();
 sg13g2_fill_2 FILLER_43_1410 ();
 sg13g2_fill_2 FILLER_43_1425 ();
 sg13g2_fill_1 FILLER_43_1427 ();
 sg13g2_decap_4 FILLER_43_1438 ();
 sg13g2_fill_1 FILLER_43_1442 ();
 sg13g2_fill_2 FILLER_43_1451 ();
 sg13g2_fill_1 FILLER_43_1453 ();
 sg13g2_decap_8 FILLER_43_1457 ();
 sg13g2_decap_8 FILLER_43_1464 ();
 sg13g2_decap_8 FILLER_43_1471 ();
 sg13g2_fill_2 FILLER_43_1478 ();
 sg13g2_decap_8 FILLER_43_1489 ();
 sg13g2_decap_8 FILLER_43_1496 ();
 sg13g2_fill_2 FILLER_43_1520 ();
 sg13g2_decap_8 FILLER_43_1526 ();
 sg13g2_fill_2 FILLER_43_1533 ();
 sg13g2_decap_8 FILLER_43_1539 ();
 sg13g2_decap_8 FILLER_43_1546 ();
 sg13g2_decap_8 FILLER_43_1553 ();
 sg13g2_decap_8 FILLER_43_1560 ();
 sg13g2_decap_8 FILLER_43_1567 ();
 sg13g2_fill_1 FILLER_43_1574 ();
 sg13g2_fill_1 FILLER_43_1609 ();
 sg13g2_decap_8 FILLER_43_1660 ();
 sg13g2_fill_2 FILLER_43_1667 ();
 sg13g2_fill_2 FILLER_43_1682 ();
 sg13g2_decap_4 FILLER_43_1725 ();
 sg13g2_fill_2 FILLER_43_1729 ();
 sg13g2_fill_2 FILLER_43_1755 ();
 sg13g2_fill_1 FILLER_43_1757 ();
 sg13g2_fill_1 FILLER_43_1788 ();
 sg13g2_fill_1 FILLER_43_1794 ();
 sg13g2_fill_2 FILLER_43_1808 ();
 sg13g2_fill_1 FILLER_43_1810 ();
 sg13g2_fill_2 FILLER_43_1822 ();
 sg13g2_decap_4 FILLER_43_1827 ();
 sg13g2_fill_1 FILLER_43_1867 ();
 sg13g2_fill_1 FILLER_43_1898 ();
 sg13g2_fill_2 FILLER_43_1903 ();
 sg13g2_decap_4 FILLER_43_1909 ();
 sg13g2_fill_2 FILLER_43_1925 ();
 sg13g2_fill_2 FILLER_43_1930 ();
 sg13g2_decap_8 FILLER_43_1941 ();
 sg13g2_decap_4 FILLER_43_1948 ();
 sg13g2_fill_1 FILLER_43_1952 ();
 sg13g2_decap_4 FILLER_43_1979 ();
 sg13g2_decap_4 FILLER_43_2001 ();
 sg13g2_decap_8 FILLER_43_2024 ();
 sg13g2_decap_4 FILLER_43_2031 ();
 sg13g2_fill_2 FILLER_43_2035 ();
 sg13g2_fill_1 FILLER_43_2125 ();
 sg13g2_decap_8 FILLER_43_2162 ();
 sg13g2_decap_8 FILLER_43_2169 ();
 sg13g2_decap_4 FILLER_43_2176 ();
 sg13g2_fill_1 FILLER_43_2180 ();
 sg13g2_decap_8 FILLER_43_2207 ();
 sg13g2_decap_4 FILLER_43_2214 ();
 sg13g2_fill_2 FILLER_43_2286 ();
 sg13g2_fill_1 FILLER_43_2301 ();
 sg13g2_fill_2 FILLER_43_2328 ();
 sg13g2_fill_1 FILLER_43_2330 ();
 sg13g2_fill_2 FILLER_43_2383 ();
 sg13g2_fill_2 FILLER_43_2423 ();
 sg13g2_fill_1 FILLER_43_2454 ();
 sg13g2_fill_1 FILLER_43_2461 ();
 sg13g2_fill_1 FILLER_43_2493 ();
 sg13g2_fill_2 FILLER_43_2505 ();
 sg13g2_fill_2 FILLER_43_2560 ();
 sg13g2_fill_1 FILLER_43_2584 ();
 sg13g2_fill_2 FILLER_43_2598 ();
 sg13g2_fill_2 FILLER_43_2621 ();
 sg13g2_fill_1 FILLER_43_2660 ();
 sg13g2_fill_2 FILLER_43_2668 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_decap_4 FILLER_44_28 ();
 sg13g2_fill_2 FILLER_44_32 ();
 sg13g2_fill_1 FILLER_44_71 ();
 sg13g2_fill_2 FILLER_44_91 ();
 sg13g2_decap_4 FILLER_44_142 ();
 sg13g2_fill_2 FILLER_44_160 ();
 sg13g2_fill_2 FILLER_44_170 ();
 sg13g2_decap_4 FILLER_44_180 ();
 sg13g2_decap_8 FILLER_44_199 ();
 sg13g2_fill_2 FILLER_44_206 ();
 sg13g2_decap_4 FILLER_44_222 ();
 sg13g2_fill_2 FILLER_44_230 ();
 sg13g2_fill_1 FILLER_44_232 ();
 sg13g2_decap_8 FILLER_44_241 ();
 sg13g2_decap_8 FILLER_44_248 ();
 sg13g2_fill_1 FILLER_44_255 ();
 sg13g2_fill_2 FILLER_44_276 ();
 sg13g2_fill_2 FILLER_44_323 ();
 sg13g2_fill_2 FILLER_44_335 ();
 sg13g2_fill_1 FILLER_44_365 ();
 sg13g2_fill_1 FILLER_44_377 ();
 sg13g2_decap_8 FILLER_44_386 ();
 sg13g2_decap_8 FILLER_44_393 ();
 sg13g2_decap_8 FILLER_44_400 ();
 sg13g2_decap_8 FILLER_44_407 ();
 sg13g2_decap_4 FILLER_44_414 ();
 sg13g2_fill_2 FILLER_44_447 ();
 sg13g2_fill_1 FILLER_44_449 ();
 sg13g2_fill_1 FILLER_44_456 ();
 sg13g2_fill_2 FILLER_44_463 ();
 sg13g2_fill_1 FILLER_44_471 ();
 sg13g2_fill_2 FILLER_44_501 ();
 sg13g2_fill_2 FILLER_44_529 ();
 sg13g2_fill_1 FILLER_44_531 ();
 sg13g2_decap_4 FILLER_44_586 ();
 sg13g2_fill_2 FILLER_44_590 ();
 sg13g2_fill_1 FILLER_44_638 ();
 sg13g2_fill_2 FILLER_44_659 ();
 sg13g2_fill_1 FILLER_44_688 ();
 sg13g2_fill_1 FILLER_44_699 ();
 sg13g2_decap_8 FILLER_44_705 ();
 sg13g2_fill_1 FILLER_44_712 ();
 sg13g2_decap_4 FILLER_44_716 ();
 sg13g2_fill_1 FILLER_44_720 ();
 sg13g2_fill_2 FILLER_44_729 ();
 sg13g2_fill_1 FILLER_44_731 ();
 sg13g2_decap_8 FILLER_44_742 ();
 sg13g2_decap_4 FILLER_44_749 ();
 sg13g2_fill_1 FILLER_44_753 ();
 sg13g2_fill_1 FILLER_44_768 ();
 sg13g2_decap_8 FILLER_44_796 ();
 sg13g2_fill_1 FILLER_44_807 ();
 sg13g2_decap_8 FILLER_44_848 ();
 sg13g2_decap_8 FILLER_44_855 ();
 sg13g2_decap_4 FILLER_44_862 ();
 sg13g2_fill_2 FILLER_44_866 ();
 sg13g2_decap_8 FILLER_44_872 ();
 sg13g2_decap_4 FILLER_44_879 ();
 sg13g2_fill_2 FILLER_44_883 ();
 sg13g2_decap_8 FILLER_44_921 ();
 sg13g2_fill_2 FILLER_44_928 ();
 sg13g2_fill_1 FILLER_44_930 ();
 sg13g2_decap_8 FILLER_44_944 ();
 sg13g2_fill_2 FILLER_44_951 ();
 sg13g2_fill_2 FILLER_44_958 ();
 sg13g2_fill_2 FILLER_44_965 ();
 sg13g2_fill_1 FILLER_44_971 ();
 sg13g2_fill_2 FILLER_44_1025 ();
 sg13g2_fill_2 FILLER_44_1041 ();
 sg13g2_fill_1 FILLER_44_1043 ();
 sg13g2_fill_1 FILLER_44_1084 ();
 sg13g2_fill_1 FILLER_44_1224 ();
 sg13g2_fill_2 FILLER_44_1239 ();
 sg13g2_fill_2 FILLER_44_1253 ();
 sg13g2_fill_2 FILLER_44_1292 ();
 sg13g2_fill_1 FILLER_44_1305 ();
 sg13g2_fill_1 FILLER_44_1311 ();
 sg13g2_fill_1 FILLER_44_1318 ();
 sg13g2_fill_1 FILLER_44_1327 ();
 sg13g2_fill_1 FILLER_44_1333 ();
 sg13g2_decap_8 FILLER_44_1343 ();
 sg13g2_decap_8 FILLER_44_1350 ();
 sg13g2_fill_2 FILLER_44_1357 ();
 sg13g2_fill_1 FILLER_44_1359 ();
 sg13g2_fill_1 FILLER_44_1365 ();
 sg13g2_decap_4 FILLER_44_1387 ();
 sg13g2_fill_2 FILLER_44_1391 ();
 sg13g2_fill_2 FILLER_44_1398 ();
 sg13g2_fill_1 FILLER_44_1400 ();
 sg13g2_decap_4 FILLER_44_1411 ();
 sg13g2_fill_1 FILLER_44_1415 ();
 sg13g2_fill_2 FILLER_44_1431 ();
 sg13g2_fill_1 FILLER_44_1437 ();
 sg13g2_decap_8 FILLER_44_1455 ();
 sg13g2_fill_1 FILLER_44_1462 ();
 sg13g2_fill_2 FILLER_44_1467 ();
 sg13g2_fill_1 FILLER_44_1469 ();
 sg13g2_fill_2 FILLER_44_1482 ();
 sg13g2_fill_2 FILLER_44_1497 ();
 sg13g2_fill_2 FILLER_44_1511 ();
 sg13g2_decap_4 FILLER_44_1551 ();
 sg13g2_fill_2 FILLER_44_1592 ();
 sg13g2_fill_2 FILLER_44_1641 ();
 sg13g2_fill_1 FILLER_44_1648 ();
 sg13g2_fill_2 FILLER_44_1656 ();
 sg13g2_fill_1 FILLER_44_1658 ();
 sg13g2_fill_2 FILLER_44_1667 ();
 sg13g2_fill_1 FILLER_44_1672 ();
 sg13g2_fill_1 FILLER_44_1678 ();
 sg13g2_fill_1 FILLER_44_1689 ();
 sg13g2_decap_4 FILLER_44_1695 ();
 sg13g2_fill_1 FILLER_44_1699 ();
 sg13g2_fill_1 FILLER_44_1715 ();
 sg13g2_fill_1 FILLER_44_1722 ();
 sg13g2_fill_1 FILLER_44_1751 ();
 sg13g2_fill_2 FILLER_44_1772 ();
 sg13g2_fill_1 FILLER_44_1774 ();
 sg13g2_fill_1 FILLER_44_1791 ();
 sg13g2_fill_2 FILLER_44_1810 ();
 sg13g2_decap_4 FILLER_44_1829 ();
 sg13g2_fill_1 FILLER_44_1833 ();
 sg13g2_fill_2 FILLER_44_1843 ();
 sg13g2_fill_1 FILLER_44_1845 ();
 sg13g2_fill_2 FILLER_44_1854 ();
 sg13g2_decap_4 FILLER_44_1860 ();
 sg13g2_fill_1 FILLER_44_1864 ();
 sg13g2_fill_2 FILLER_44_1869 ();
 sg13g2_fill_1 FILLER_44_1871 ();
 sg13g2_fill_2 FILLER_44_1876 ();
 sg13g2_fill_2 FILLER_44_1882 ();
 sg13g2_fill_1 FILLER_44_1910 ();
 sg13g2_decap_8 FILLER_44_1918 ();
 sg13g2_fill_2 FILLER_44_1925 ();
 sg13g2_fill_2 FILLER_44_1957 ();
 sg13g2_fill_2 FILLER_44_1963 ();
 sg13g2_fill_1 FILLER_44_1965 ();
 sg13g2_decap_4 FILLER_44_1976 ();
 sg13g2_fill_1 FILLER_44_1980 ();
 sg13g2_decap_8 FILLER_44_1989 ();
 sg13g2_fill_2 FILLER_44_1996 ();
 sg13g2_fill_1 FILLER_44_1998 ();
 sg13g2_fill_1 FILLER_44_2057 ();
 sg13g2_decap_8 FILLER_44_2071 ();
 sg13g2_decap_4 FILLER_44_2078 ();
 sg13g2_decap_8 FILLER_44_2099 ();
 sg13g2_fill_2 FILLER_44_2106 ();
 sg13g2_fill_1 FILLER_44_2108 ();
 sg13g2_fill_1 FILLER_44_2160 ();
 sg13g2_fill_2 FILLER_44_2171 ();
 sg13g2_decap_8 FILLER_44_2183 ();
 sg13g2_fill_2 FILLER_44_2190 ();
 sg13g2_decap_8 FILLER_44_2279 ();
 sg13g2_fill_2 FILLER_44_2286 ();
 sg13g2_decap_8 FILLER_44_2321 ();
 sg13g2_decap_4 FILLER_44_2328 ();
 sg13g2_fill_2 FILLER_44_2342 ();
 sg13g2_fill_2 FILLER_44_2443 ();
 sg13g2_fill_2 FILLER_44_2517 ();
 sg13g2_fill_2 FILLER_44_2551 ();
 sg13g2_fill_2 FILLER_44_2579 ();
 sg13g2_fill_2 FILLER_44_2640 ();
 sg13g2_fill_2 FILLER_44_2668 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_79 ();
 sg13g2_fill_1 FILLER_45_81 ();
 sg13g2_decap_8 FILLER_45_87 ();
 sg13g2_decap_4 FILLER_45_94 ();
 sg13g2_fill_1 FILLER_45_138 ();
 sg13g2_decap_4 FILLER_45_184 ();
 sg13g2_decap_8 FILLER_45_218 ();
 sg13g2_decap_8 FILLER_45_251 ();
 sg13g2_fill_2 FILLER_45_258 ();
 sg13g2_fill_1 FILLER_45_275 ();
 sg13g2_fill_2 FILLER_45_290 ();
 sg13g2_fill_1 FILLER_45_292 ();
 sg13g2_fill_1 FILLER_45_297 ();
 sg13g2_fill_1 FILLER_45_311 ();
 sg13g2_decap_4 FILLER_45_357 ();
 sg13g2_fill_1 FILLER_45_361 ();
 sg13g2_fill_1 FILLER_45_372 ();
 sg13g2_fill_1 FILLER_45_381 ();
 sg13g2_fill_1 FILLER_45_446 ();
 sg13g2_fill_2 FILLER_45_452 ();
 sg13g2_fill_1 FILLER_45_454 ();
 sg13g2_decap_4 FILLER_45_460 ();
 sg13g2_fill_2 FILLER_45_464 ();
 sg13g2_fill_2 FILLER_45_481 ();
 sg13g2_fill_1 FILLER_45_483 ();
 sg13g2_fill_2 FILLER_45_503 ();
 sg13g2_fill_1 FILLER_45_509 ();
 sg13g2_fill_2 FILLER_45_518 ();
 sg13g2_fill_1 FILLER_45_520 ();
 sg13g2_fill_1 FILLER_45_542 ();
 sg13g2_fill_1 FILLER_45_572 ();
 sg13g2_fill_2 FILLER_45_583 ();
 sg13g2_fill_1 FILLER_45_585 ();
 sg13g2_fill_2 FILLER_45_601 ();
 sg13g2_fill_1 FILLER_45_639 ();
 sg13g2_fill_1 FILLER_45_645 ();
 sg13g2_fill_2 FILLER_45_673 ();
 sg13g2_fill_1 FILLER_45_700 ();
 sg13g2_fill_1 FILLER_45_712 ();
 sg13g2_fill_1 FILLER_45_728 ();
 sg13g2_decap_8 FILLER_45_742 ();
 sg13g2_fill_1 FILLER_45_749 ();
 sg13g2_decap_4 FILLER_45_754 ();
 sg13g2_fill_1 FILLER_45_773 ();
 sg13g2_decap_8 FILLER_45_786 ();
 sg13g2_decap_8 FILLER_45_793 ();
 sg13g2_decap_4 FILLER_45_804 ();
 sg13g2_fill_1 FILLER_45_811 ();
 sg13g2_fill_2 FILLER_45_877 ();
 sg13g2_fill_1 FILLER_45_883 ();
 sg13g2_fill_2 FILLER_45_888 ();
 sg13g2_fill_1 FILLER_45_890 ();
 sg13g2_fill_2 FILLER_45_901 ();
 sg13g2_decap_8 FILLER_45_907 ();
 sg13g2_fill_2 FILLER_45_914 ();
 sg13g2_fill_1 FILLER_45_916 ();
 sg13g2_decap_8 FILLER_45_932 ();
 sg13g2_fill_1 FILLER_45_943 ();
 sg13g2_fill_1 FILLER_45_950 ();
 sg13g2_decap_8 FILLER_45_977 ();
 sg13g2_fill_2 FILLER_45_984 ();
 sg13g2_fill_1 FILLER_45_986 ();
 sg13g2_fill_1 FILLER_45_992 ();
 sg13g2_decap_4 FILLER_45_997 ();
 sg13g2_fill_2 FILLER_45_1001 ();
 sg13g2_decap_8 FILLER_45_1008 ();
 sg13g2_decap_4 FILLER_45_1015 ();
 sg13g2_fill_1 FILLER_45_1019 ();
 sg13g2_fill_2 FILLER_45_1026 ();
 sg13g2_fill_1 FILLER_45_1028 ();
 sg13g2_decap_8 FILLER_45_1101 ();
 sg13g2_fill_1 FILLER_45_1108 ();
 sg13g2_fill_2 FILLER_45_1115 ();
 sg13g2_fill_1 FILLER_45_1129 ();
 sg13g2_fill_2 FILLER_45_1140 ();
 sg13g2_fill_1 FILLER_45_1164 ();
 sg13g2_fill_2 FILLER_45_1189 ();
 sg13g2_fill_1 FILLER_45_1191 ();
 sg13g2_fill_1 FILLER_45_1218 ();
 sg13g2_fill_2 FILLER_45_1238 ();
 sg13g2_fill_1 FILLER_45_1255 ();
 sg13g2_fill_1 FILLER_45_1264 ();
 sg13g2_fill_1 FILLER_45_1270 ();
 sg13g2_fill_2 FILLER_45_1276 ();
 sg13g2_fill_1 FILLER_45_1292 ();
 sg13g2_fill_2 FILLER_45_1299 ();
 sg13g2_fill_2 FILLER_45_1306 ();
 sg13g2_fill_2 FILLER_45_1329 ();
 sg13g2_fill_2 FILLER_45_1336 ();
 sg13g2_fill_1 FILLER_45_1338 ();
 sg13g2_decap_8 FILLER_45_1348 ();
 sg13g2_fill_2 FILLER_45_1355 ();
 sg13g2_fill_1 FILLER_45_1357 ();
 sg13g2_decap_4 FILLER_45_1368 ();
 sg13g2_decap_4 FILLER_45_1389 ();
 sg13g2_fill_2 FILLER_45_1393 ();
 sg13g2_decap_4 FILLER_45_1432 ();
 sg13g2_decap_8 FILLER_45_1440 ();
 sg13g2_fill_2 FILLER_45_1447 ();
 sg13g2_decap_8 FILLER_45_1454 ();
 sg13g2_fill_2 FILLER_45_1461 ();
 sg13g2_fill_2 FILLER_45_1501 ();
 sg13g2_decap_4 FILLER_45_1541 ();
 sg13g2_fill_1 FILLER_45_1545 ();
 sg13g2_decap_8 FILLER_45_1550 ();
 sg13g2_decap_4 FILLER_45_1557 ();
 sg13g2_fill_1 FILLER_45_1561 ();
 sg13g2_decap_4 FILLER_45_1566 ();
 sg13g2_fill_1 FILLER_45_1570 ();
 sg13g2_fill_1 FILLER_45_1576 ();
 sg13g2_decap_8 FILLER_45_1582 ();
 sg13g2_decap_4 FILLER_45_1589 ();
 sg13g2_fill_1 FILLER_45_1593 ();
 sg13g2_decap_8 FILLER_45_1599 ();
 sg13g2_decap_8 FILLER_45_1610 ();
 sg13g2_decap_4 FILLER_45_1617 ();
 sg13g2_fill_2 FILLER_45_1639 ();
 sg13g2_fill_2 FILLER_45_1667 ();
 sg13g2_decap_4 FILLER_45_1684 ();
 sg13g2_fill_2 FILLER_45_1688 ();
 sg13g2_fill_2 FILLER_45_1695 ();
 sg13g2_fill_1 FILLER_45_1697 ();
 sg13g2_fill_2 FILLER_45_1718 ();
 sg13g2_fill_1 FILLER_45_1730 ();
 sg13g2_fill_1 FILLER_45_1741 ();
 sg13g2_fill_1 FILLER_45_1751 ();
 sg13g2_fill_2 FILLER_45_1757 ();
 sg13g2_fill_2 FILLER_45_1821 ();
 sg13g2_fill_2 FILLER_45_1849 ();
 sg13g2_fill_2 FILLER_45_1856 ();
 sg13g2_fill_2 FILLER_45_1899 ();
 sg13g2_decap_8 FILLER_45_1919 ();
 sg13g2_fill_1 FILLER_45_1926 ();
 sg13g2_decap_8 FILLER_45_1953 ();
 sg13g2_decap_8 FILLER_45_1960 ();
 sg13g2_decap_4 FILLER_45_1967 ();
 sg13g2_fill_1 FILLER_45_1971 ();
 sg13g2_decap_8 FILLER_45_1977 ();
 sg13g2_fill_2 FILLER_45_1988 ();
 sg13g2_fill_1 FILLER_45_1990 ();
 sg13g2_fill_2 FILLER_45_2001 ();
 sg13g2_fill_1 FILLER_45_2003 ();
 sg13g2_decap_8 FILLER_45_2040 ();
 sg13g2_fill_2 FILLER_45_2047 ();
 sg13g2_fill_1 FILLER_45_2049 ();
 sg13g2_fill_2 FILLER_45_2055 ();
 sg13g2_fill_1 FILLER_45_2057 ();
 sg13g2_fill_2 FILLER_45_2066 ();
 sg13g2_fill_1 FILLER_45_2068 ();
 sg13g2_decap_8 FILLER_45_2113 ();
 sg13g2_fill_1 FILLER_45_2120 ();
 sg13g2_fill_1 FILLER_45_2197 ();
 sg13g2_fill_1 FILLER_45_2224 ();
 sg13g2_fill_2 FILLER_45_2261 ();
 sg13g2_decap_8 FILLER_45_2276 ();
 sg13g2_fill_2 FILLER_45_2283 ();
 sg13g2_fill_2 FILLER_45_2295 ();
 sg13g2_fill_1 FILLER_45_2297 ();
 sg13g2_fill_2 FILLER_45_2301 ();
 sg13g2_fill_2 FILLER_45_2342 ();
 sg13g2_fill_2 FILLER_45_2355 ();
 sg13g2_fill_1 FILLER_45_2408 ();
 sg13g2_fill_2 FILLER_45_2442 ();
 sg13g2_fill_1 FILLER_45_2451 ();
 sg13g2_fill_1 FILLER_45_2471 ();
 sg13g2_fill_1 FILLER_45_2494 ();
 sg13g2_fill_1 FILLER_45_2508 ();
 sg13g2_fill_2 FILLER_45_2534 ();
 sg13g2_fill_1 FILLER_45_2546 ();
 sg13g2_fill_1 FILLER_45_2553 ();
 sg13g2_fill_1 FILLER_45_2580 ();
 sg13g2_fill_2 FILLER_45_2633 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_12 ();
 sg13g2_decap_4 FILLER_46_19 ();
 sg13g2_fill_1 FILLER_46_23 ();
 sg13g2_fill_2 FILLER_46_42 ();
 sg13g2_fill_1 FILLER_46_44 ();
 sg13g2_decap_8 FILLER_46_90 ();
 sg13g2_decap_8 FILLER_46_97 ();
 sg13g2_fill_2 FILLER_46_104 ();
 sg13g2_fill_1 FILLER_46_106 ();
 sg13g2_decap_8 FILLER_46_116 ();
 sg13g2_fill_1 FILLER_46_123 ();
 sg13g2_fill_1 FILLER_46_132 ();
 sg13g2_fill_1 FILLER_46_141 ();
 sg13g2_fill_1 FILLER_46_147 ();
 sg13g2_fill_1 FILLER_46_154 ();
 sg13g2_fill_2 FILLER_46_254 ();
 sg13g2_decap_8 FILLER_46_270 ();
 sg13g2_fill_2 FILLER_46_277 ();
 sg13g2_fill_1 FILLER_46_279 ();
 sg13g2_decap_4 FILLER_46_283 ();
 sg13g2_fill_2 FILLER_46_287 ();
 sg13g2_decap_4 FILLER_46_294 ();
 sg13g2_fill_2 FILLER_46_298 ();
 sg13g2_fill_2 FILLER_46_309 ();
 sg13g2_fill_1 FILLER_46_391 ();
 sg13g2_fill_1 FILLER_46_396 ();
 sg13g2_decap_4 FILLER_46_428 ();
 sg13g2_decap_4 FILLER_46_438 ();
 sg13g2_fill_2 FILLER_46_442 ();
 sg13g2_decap_4 FILLER_46_470 ();
 sg13g2_fill_2 FILLER_46_474 ();
 sg13g2_fill_1 FILLER_46_482 ();
 sg13g2_decap_8 FILLER_46_498 ();
 sg13g2_decap_4 FILLER_46_514 ();
 sg13g2_decap_8 FILLER_46_528 ();
 sg13g2_decap_8 FILLER_46_535 ();
 sg13g2_decap_4 FILLER_46_542 ();
 sg13g2_fill_1 FILLER_46_546 ();
 sg13g2_fill_2 FILLER_46_656 ();
 sg13g2_fill_2 FILLER_46_698 ();
 sg13g2_fill_2 FILLER_46_710 ();
 sg13g2_fill_1 FILLER_46_730 ();
 sg13g2_fill_2 FILLER_46_741 ();
 sg13g2_fill_2 FILLER_46_781 ();
 sg13g2_decap_4 FILLER_46_800 ();
 sg13g2_fill_1 FILLER_46_804 ();
 sg13g2_decap_8 FILLER_46_809 ();
 sg13g2_decap_8 FILLER_46_816 ();
 sg13g2_fill_1 FILLER_46_823 ();
 sg13g2_fill_2 FILLER_46_828 ();
 sg13g2_fill_1 FILLER_46_856 ();
 sg13g2_decap_4 FILLER_46_871 ();
 sg13g2_decap_8 FILLER_46_905 ();
 sg13g2_fill_2 FILLER_46_912 ();
 sg13g2_fill_1 FILLER_46_914 ();
 sg13g2_fill_1 FILLER_46_921 ();
 sg13g2_fill_1 FILLER_46_944 ();
 sg13g2_fill_1 FILLER_46_955 ();
 sg13g2_decap_4 FILLER_46_965 ();
 sg13g2_fill_2 FILLER_46_969 ();
 sg13g2_decap_4 FILLER_46_975 ();
 sg13g2_fill_2 FILLER_46_979 ();
 sg13g2_decap_4 FILLER_46_995 ();
 sg13g2_decap_8 FILLER_46_1035 ();
 sg13g2_fill_2 FILLER_46_1042 ();
 sg13g2_fill_2 FILLER_46_1070 ();
 sg13g2_decap_8 FILLER_46_1112 ();
 sg13g2_decap_8 FILLER_46_1119 ();
 sg13g2_decap_8 FILLER_46_1126 ();
 sg13g2_fill_1 FILLER_46_1133 ();
 sg13g2_decap_8 FILLER_46_1137 ();
 sg13g2_decap_4 FILLER_46_1144 ();
 sg13g2_fill_2 FILLER_46_1148 ();
 sg13g2_decap_8 FILLER_46_1154 ();
 sg13g2_decap_8 FILLER_46_1175 ();
 sg13g2_decap_8 FILLER_46_1182 ();
 sg13g2_fill_1 FILLER_46_1189 ();
 sg13g2_fill_2 FILLER_46_1204 ();
 sg13g2_fill_1 FILLER_46_1206 ();
 sg13g2_fill_2 FILLER_46_1243 ();
 sg13g2_fill_1 FILLER_46_1264 ();
 sg13g2_fill_1 FILLER_46_1270 ();
 sg13g2_fill_1 FILLER_46_1287 ();
 sg13g2_fill_1 FILLER_46_1295 ();
 sg13g2_fill_1 FILLER_46_1301 ();
 sg13g2_decap_4 FILLER_46_1336 ();
 sg13g2_fill_2 FILLER_46_1345 ();
 sg13g2_decap_8 FILLER_46_1356 ();
 sg13g2_fill_2 FILLER_46_1363 ();
 sg13g2_fill_2 FILLER_46_1376 ();
 sg13g2_fill_1 FILLER_46_1378 ();
 sg13g2_decap_4 FILLER_46_1410 ();
 sg13g2_fill_1 FILLER_46_1414 ();
 sg13g2_fill_2 FILLER_46_1433 ();
 sg13g2_decap_8 FILLER_46_1449 ();
 sg13g2_fill_2 FILLER_46_1456 ();
 sg13g2_fill_2 FILLER_46_1466 ();
 sg13g2_fill_1 FILLER_46_1487 ();
 sg13g2_decap_4 FILLER_46_1548 ();
 sg13g2_fill_2 FILLER_46_1552 ();
 sg13g2_fill_1 FILLER_46_1567 ();
 sg13g2_decap_8 FILLER_46_1601 ();
 sg13g2_decap_8 FILLER_46_1608 ();
 sg13g2_decap_8 FILLER_46_1615 ();
 sg13g2_decap_8 FILLER_46_1691 ();
 sg13g2_fill_1 FILLER_46_1698 ();
 sg13g2_decap_4 FILLER_46_1709 ();
 sg13g2_fill_2 FILLER_46_1724 ();
 sg13g2_fill_1 FILLER_46_1740 ();
 sg13g2_fill_2 FILLER_46_1768 ();
 sg13g2_fill_1 FILLER_46_1777 ();
 sg13g2_fill_2 FILLER_46_1804 ();
 sg13g2_fill_2 FILLER_46_1810 ();
 sg13g2_decap_4 FILLER_46_1815 ();
 sg13g2_decap_4 FILLER_46_1849 ();
 sg13g2_fill_1 FILLER_46_1931 ();
 sg13g2_decap_8 FILLER_46_1958 ();
 sg13g2_decap_8 FILLER_46_1965 ();
 sg13g2_fill_1 FILLER_46_1972 ();
 sg13g2_fill_1 FILLER_46_1977 ();
 sg13g2_fill_1 FILLER_46_2004 ();
 sg13g2_decap_8 FILLER_46_2030 ();
 sg13g2_decap_8 FILLER_46_2037 ();
 sg13g2_decap_8 FILLER_46_2044 ();
 sg13g2_decap_8 FILLER_46_2051 ();
 sg13g2_decap_8 FILLER_46_2058 ();
 sg13g2_decap_4 FILLER_46_2065 ();
 sg13g2_decap_4 FILLER_46_2095 ();
 sg13g2_decap_8 FILLER_46_2103 ();
 sg13g2_fill_1 FILLER_46_2110 ();
 sg13g2_fill_2 FILLER_46_2116 ();
 sg13g2_fill_1 FILLER_46_2118 ();
 sg13g2_decap_4 FILLER_46_2123 ();
 sg13g2_fill_1 FILLER_46_2163 ();
 sg13g2_fill_1 FILLER_46_2222 ();
 sg13g2_decap_8 FILLER_46_2227 ();
 sg13g2_fill_1 FILLER_46_2261 ();
 sg13g2_decap_8 FILLER_46_2266 ();
 sg13g2_decap_8 FILLER_46_2273 ();
 sg13g2_fill_2 FILLER_46_2311 ();
 sg13g2_fill_1 FILLER_46_2317 ();
 sg13g2_fill_1 FILLER_46_2344 ();
 sg13g2_fill_2 FILLER_46_2351 ();
 sg13g2_fill_2 FILLER_46_2478 ();
 sg13g2_fill_2 FILLER_46_2483 ();
 sg13g2_fill_1 FILLER_46_2490 ();
 sg13g2_fill_1 FILLER_46_2587 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_11 ();
 sg13g2_fill_2 FILLER_47_60 ();
 sg13g2_fill_1 FILLER_47_62 ();
 sg13g2_fill_2 FILLER_47_101 ();
 sg13g2_fill_1 FILLER_47_103 ();
 sg13g2_decap_4 FILLER_47_130 ();
 sg13g2_fill_2 FILLER_47_134 ();
 sg13g2_decap_8 FILLER_47_146 ();
 sg13g2_fill_1 FILLER_47_153 ();
 sg13g2_decap_8 FILLER_47_158 ();
 sg13g2_fill_2 FILLER_47_165 ();
 sg13g2_fill_1 FILLER_47_167 ();
 sg13g2_fill_2 FILLER_47_222 ();
 sg13g2_decap_4 FILLER_47_243 ();
 sg13g2_fill_1 FILLER_47_247 ();
 sg13g2_fill_2 FILLER_47_302 ();
 sg13g2_fill_1 FILLER_47_304 ();
 sg13g2_fill_2 FILLER_47_316 ();
 sg13g2_fill_1 FILLER_47_318 ();
 sg13g2_decap_8 FILLER_47_324 ();
 sg13g2_fill_2 FILLER_47_335 ();
 sg13g2_fill_2 FILLER_47_347 ();
 sg13g2_fill_1 FILLER_47_349 ();
 sg13g2_fill_2 FILLER_47_388 ();
 sg13g2_fill_1 FILLER_47_404 ();
 sg13g2_decap_8 FILLER_47_430 ();
 sg13g2_decap_8 FILLER_47_437 ();
 sg13g2_decap_4 FILLER_47_444 ();
 sg13g2_decap_4 FILLER_47_478 ();
 sg13g2_fill_1 FILLER_47_482 ();
 sg13g2_decap_8 FILLER_47_489 ();
 sg13g2_fill_1 FILLER_47_496 ();
 sg13g2_decap_4 FILLER_47_535 ();
 sg13g2_fill_2 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_546 ();
 sg13g2_fill_2 FILLER_47_553 ();
 sg13g2_fill_1 FILLER_47_568 ();
 sg13g2_fill_2 FILLER_47_625 ();
 sg13g2_fill_2 FILLER_47_632 ();
 sg13g2_fill_1 FILLER_47_638 ();
 sg13g2_fill_2 FILLER_47_681 ();
 sg13g2_fill_1 FILLER_47_688 ();
 sg13g2_fill_2 FILLER_47_724 ();
 sg13g2_fill_1 FILLER_47_726 ();
 sg13g2_fill_1 FILLER_47_750 ();
 sg13g2_fill_2 FILLER_47_756 ();
 sg13g2_fill_2 FILLER_47_763 ();
 sg13g2_fill_2 FILLER_47_773 ();
 sg13g2_fill_1 FILLER_47_775 ();
 sg13g2_decap_8 FILLER_47_807 ();
 sg13g2_decap_8 FILLER_47_814 ();
 sg13g2_fill_1 FILLER_47_821 ();
 sg13g2_decap_8 FILLER_47_878 ();
 sg13g2_decap_8 FILLER_47_885 ();
 sg13g2_decap_8 FILLER_47_892 ();
 sg13g2_decap_8 FILLER_47_899 ();
 sg13g2_decap_4 FILLER_47_906 ();
 sg13g2_fill_1 FILLER_47_910 ();
 sg13g2_decap_8 FILLER_47_916 ();
 sg13g2_decap_8 FILLER_47_923 ();
 sg13g2_fill_1 FILLER_47_944 ();
 sg13g2_fill_1 FILLER_47_958 ();
 sg13g2_fill_2 FILLER_47_969 ();
 sg13g2_fill_1 FILLER_47_975 ();
 sg13g2_fill_1 FILLER_47_982 ();
 sg13g2_fill_2 FILLER_47_1038 ();
 sg13g2_fill_1 FILLER_47_1050 ();
 sg13g2_decap_4 FILLER_47_1055 ();
 sg13g2_fill_1 FILLER_47_1059 ();
 sg13g2_decap_8 FILLER_47_1121 ();
 sg13g2_fill_2 FILLER_47_1128 ();
 sg13g2_decap_8 FILLER_47_1135 ();
 sg13g2_fill_1 FILLER_47_1142 ();
 sg13g2_fill_2 FILLER_47_1169 ();
 sg13g2_fill_1 FILLER_47_1171 ();
 sg13g2_decap_4 FILLER_47_1208 ();
 sg13g2_fill_1 FILLER_47_1212 ();
 sg13g2_decap_8 FILLER_47_1221 ();
 sg13g2_decap_4 FILLER_47_1228 ();
 sg13g2_decap_4 FILLER_47_1236 ();
 sg13g2_fill_1 FILLER_47_1258 ();
 sg13g2_decap_4 FILLER_47_1265 ();
 sg13g2_fill_2 FILLER_47_1269 ();
 sg13g2_fill_1 FILLER_47_1295 ();
 sg13g2_decap_8 FILLER_47_1301 ();
 sg13g2_fill_2 FILLER_47_1308 ();
 sg13g2_fill_1 FILLER_47_1310 ();
 sg13g2_fill_2 FILLER_47_1329 ();
 sg13g2_fill_1 FILLER_47_1331 ();
 sg13g2_decap_4 FILLER_47_1337 ();
 sg13g2_fill_1 FILLER_47_1341 ();
 sg13g2_decap_8 FILLER_47_1348 ();
 sg13g2_decap_4 FILLER_47_1355 ();
 sg13g2_fill_2 FILLER_47_1359 ();
 sg13g2_fill_2 FILLER_47_1371 ();
 sg13g2_fill_1 FILLER_47_1373 ();
 sg13g2_fill_2 FILLER_47_1378 ();
 sg13g2_fill_2 FILLER_47_1404 ();
 sg13g2_fill_2 FILLER_47_1410 ();
 sg13g2_fill_1 FILLER_47_1451 ();
 sg13g2_fill_1 FILLER_47_1461 ();
 sg13g2_fill_2 FILLER_47_1520 ();
 sg13g2_decap_4 FILLER_47_1533 ();
 sg13g2_fill_2 FILLER_47_1546 ();
 sg13g2_fill_1 FILLER_47_1548 ();
 sg13g2_fill_1 FILLER_47_1553 ();
 sg13g2_fill_2 FILLER_47_1567 ();
 sg13g2_fill_2 FILLER_47_1574 ();
 sg13g2_fill_2 FILLER_47_1584 ();
 sg13g2_decap_8 FILLER_47_1608 ();
 sg13g2_decap_8 FILLER_47_1615 ();
 sg13g2_decap_8 FILLER_47_1622 ();
 sg13g2_decap_4 FILLER_47_1629 ();
 sg13g2_decap_4 FILLER_47_1694 ();
 sg13g2_decap_4 FILLER_47_1703 ();
 sg13g2_decap_4 FILLER_47_1711 ();
 sg13g2_fill_2 FILLER_47_1715 ();
 sg13g2_decap_8 FILLER_47_1721 ();
 sg13g2_fill_1 FILLER_47_1763 ();
 sg13g2_fill_2 FILLER_47_1785 ();
 sg13g2_fill_2 FILLER_47_1790 ();
 sg13g2_decap_4 FILLER_47_1823 ();
 sg13g2_fill_1 FILLER_47_1827 ();
 sg13g2_decap_8 FILLER_47_1836 ();
 sg13g2_fill_2 FILLER_47_1843 ();
 sg13g2_fill_1 FILLER_47_1845 ();
 sg13g2_fill_2 FILLER_47_1850 ();
 sg13g2_fill_2 FILLER_47_1856 ();
 sg13g2_fill_1 FILLER_47_1858 ();
 sg13g2_fill_2 FILLER_47_1864 ();
 sg13g2_fill_1 FILLER_47_1866 ();
 sg13g2_fill_1 FILLER_47_1879 ();
 sg13g2_decap_4 FILLER_47_1894 ();
 sg13g2_fill_1 FILLER_47_1898 ();
 sg13g2_fill_1 FILLER_47_1903 ();
 sg13g2_fill_2 FILLER_47_1911 ();
 sg13g2_decap_4 FILLER_47_1917 ();
 sg13g2_fill_1 FILLER_47_1921 ();
 sg13g2_fill_2 FILLER_47_1927 ();
 sg13g2_fill_1 FILLER_47_1929 ();
 sg13g2_decap_8 FILLER_47_1964 ();
 sg13g2_decap_8 FILLER_47_1971 ();
 sg13g2_fill_1 FILLER_47_1978 ();
 sg13g2_fill_2 FILLER_47_2019 ();
 sg13g2_fill_1 FILLER_47_2021 ();
 sg13g2_fill_1 FILLER_47_2036 ();
 sg13g2_fill_2 FILLER_47_2063 ();
 sg13g2_decap_8 FILLER_47_2117 ();
 sg13g2_decap_8 FILLER_47_2124 ();
 sg13g2_decap_8 FILLER_47_2131 ();
 sg13g2_fill_2 FILLER_47_2138 ();
 sg13g2_fill_2 FILLER_47_2144 ();
 sg13g2_fill_1 FILLER_47_2150 ();
 sg13g2_fill_2 FILLER_47_2182 ();
 sg13g2_fill_1 FILLER_47_2198 ();
 sg13g2_decap_4 FILLER_47_2206 ();
 sg13g2_fill_1 FILLER_47_2210 ();
 sg13g2_decap_8 FILLER_47_2216 ();
 sg13g2_decap_8 FILLER_47_2223 ();
 sg13g2_decap_8 FILLER_47_2230 ();
 sg13g2_decap_4 FILLER_47_2237 ();
 sg13g2_fill_2 FILLER_47_2241 ();
 sg13g2_decap_8 FILLER_47_2256 ();
 sg13g2_decap_8 FILLER_47_2263 ();
 sg13g2_decap_8 FILLER_47_2270 ();
 sg13g2_decap_8 FILLER_47_2277 ();
 sg13g2_decap_4 FILLER_47_2284 ();
 sg13g2_decap_8 FILLER_47_2292 ();
 sg13g2_decap_8 FILLER_47_2299 ();
 sg13g2_decap_4 FILLER_47_2306 ();
 sg13g2_fill_2 FILLER_47_2310 ();
 sg13g2_fill_2 FILLER_47_2316 ();
 sg13g2_fill_2 FILLER_47_2356 ();
 sg13g2_fill_2 FILLER_47_2365 ();
 sg13g2_fill_1 FILLER_47_2444 ();
 sg13g2_fill_1 FILLER_47_2462 ();
 sg13g2_fill_2 FILLER_47_2475 ();
 sg13g2_fill_1 FILLER_47_2520 ();
 sg13g2_fill_1 FILLER_47_2527 ();
 sg13g2_fill_2 FILLER_47_2544 ();
 sg13g2_fill_1 FILLER_47_2567 ();
 sg13g2_fill_1 FILLER_47_2574 ();
 sg13g2_fill_1 FILLER_47_2608 ();
 sg13g2_fill_2 FILLER_47_2668 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_7 ();
 sg13g2_fill_2 FILLER_48_21 ();
 sg13g2_fill_2 FILLER_48_66 ();
 sg13g2_fill_1 FILLER_48_68 ();
 sg13g2_fill_1 FILLER_48_79 ();
 sg13g2_fill_2 FILLER_48_87 ();
 sg13g2_fill_1 FILLER_48_93 ();
 sg13g2_fill_1 FILLER_48_104 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_fill_1 FILLER_48_196 ();
 sg13g2_decap_4 FILLER_48_206 ();
 sg13g2_decap_4 FILLER_48_215 ();
 sg13g2_fill_1 FILLER_48_232 ();
 sg13g2_decap_8 FILLER_48_237 ();
 sg13g2_fill_1 FILLER_48_244 ();
 sg13g2_decap_8 FILLER_48_254 ();
 sg13g2_fill_2 FILLER_48_261 ();
 sg13g2_fill_1 FILLER_48_269 ();
 sg13g2_decap_8 FILLER_48_302 ();
 sg13g2_fill_2 FILLER_48_309 ();
 sg13g2_fill_1 FILLER_48_311 ();
 sg13g2_decap_8 FILLER_48_316 ();
 sg13g2_decap_4 FILLER_48_323 ();
 sg13g2_decap_8 FILLER_48_335 ();
 sg13g2_decap_8 FILLER_48_342 ();
 sg13g2_fill_2 FILLER_48_349 ();
 sg13g2_fill_1 FILLER_48_351 ();
 sg13g2_fill_2 FILLER_48_385 ();
 sg13g2_fill_1 FILLER_48_387 ();
 sg13g2_fill_1 FILLER_48_392 ();
 sg13g2_fill_1 FILLER_48_401 ();
 sg13g2_decap_8 FILLER_48_439 ();
 sg13g2_decap_8 FILLER_48_446 ();
 sg13g2_decap_8 FILLER_48_485 ();
 sg13g2_decap_8 FILLER_48_492 ();
 sg13g2_fill_1 FILLER_48_512 ();
 sg13g2_fill_1 FILLER_48_518 ();
 sg13g2_fill_1 FILLER_48_524 ();
 sg13g2_fill_1 FILLER_48_530 ();
 sg13g2_fill_1 FILLER_48_571 ();
 sg13g2_fill_1 FILLER_48_588 ();
 sg13g2_fill_2 FILLER_48_605 ();
 sg13g2_fill_2 FILLER_48_618 ();
 sg13g2_fill_1 FILLER_48_625 ();
 sg13g2_fill_1 FILLER_48_630 ();
 sg13g2_fill_1 FILLER_48_665 ();
 sg13g2_fill_1 FILLER_48_674 ();
 sg13g2_fill_1 FILLER_48_680 ();
 sg13g2_decap_4 FILLER_48_711 ();
 sg13g2_fill_2 FILLER_48_759 ();
 sg13g2_decap_8 FILLER_48_816 ();
 sg13g2_fill_2 FILLER_48_823 ();
 sg13g2_fill_1 FILLER_48_829 ();
 sg13g2_fill_1 FILLER_48_836 ();
 sg13g2_fill_1 FILLER_48_841 ();
 sg13g2_fill_1 FILLER_48_846 ();
 sg13g2_fill_1 FILLER_48_932 ();
 sg13g2_fill_1 FILLER_48_937 ();
 sg13g2_fill_1 FILLER_48_943 ();
 sg13g2_fill_2 FILLER_48_949 ();
 sg13g2_fill_2 FILLER_48_962 ();
 sg13g2_fill_1 FILLER_48_994 ();
 sg13g2_decap_8 FILLER_48_1031 ();
 sg13g2_decap_8 FILLER_48_1038 ();
 sg13g2_decap_8 FILLER_48_1045 ();
 sg13g2_fill_2 FILLER_48_1052 ();
 sg13g2_fill_1 FILLER_48_1054 ();
 sg13g2_decap_4 FILLER_48_1065 ();
 sg13g2_decap_8 FILLER_48_1073 ();
 sg13g2_fill_2 FILLER_48_1080 ();
 sg13g2_decap_4 FILLER_48_1088 ();
 sg13g2_fill_1 FILLER_48_1092 ();
 sg13g2_decap_4 FILLER_48_1097 ();
 sg13g2_fill_2 FILLER_48_1101 ();
 sg13g2_decap_4 FILLER_48_1113 ();
 sg13g2_fill_1 FILLER_48_1117 ();
 sg13g2_fill_2 FILLER_48_1123 ();
 sg13g2_fill_1 FILLER_48_1125 ();
 sg13g2_fill_2 FILLER_48_1130 ();
 sg13g2_fill_2 FILLER_48_1136 ();
 sg13g2_fill_1 FILLER_48_1138 ();
 sg13g2_fill_1 FILLER_48_1188 ();
 sg13g2_fill_1 FILLER_48_1193 ();
 sg13g2_decap_8 FILLER_48_1204 ();
 sg13g2_decap_8 FILLER_48_1211 ();
 sg13g2_decap_8 FILLER_48_1218 ();
 sg13g2_decap_8 FILLER_48_1279 ();
 sg13g2_fill_2 FILLER_48_1286 ();
 sg13g2_decap_4 FILLER_48_1296 ();
 sg13g2_fill_2 FILLER_48_1322 ();
 sg13g2_decap_4 FILLER_48_1329 ();
 sg13g2_fill_1 FILLER_48_1333 ();
 sg13g2_decap_4 FILLER_48_1339 ();
 sg13g2_decap_4 FILLER_48_1347 ();
 sg13g2_fill_1 FILLER_48_1351 ();
 sg13g2_decap_4 FILLER_48_1361 ();
 sg13g2_fill_2 FILLER_48_1365 ();
 sg13g2_decap_4 FILLER_48_1376 ();
 sg13g2_decap_8 FILLER_48_1393 ();
 sg13g2_fill_2 FILLER_48_1400 ();
 sg13g2_decap_8 FILLER_48_1415 ();
 sg13g2_decap_8 FILLER_48_1422 ();
 sg13g2_fill_2 FILLER_48_1429 ();
 sg13g2_fill_2 FILLER_48_1436 ();
 sg13g2_fill_2 FILLER_48_1443 ();
 sg13g2_fill_1 FILLER_48_1445 ();
 sg13g2_fill_2 FILLER_48_1454 ();
 sg13g2_fill_1 FILLER_48_1456 ();
 sg13g2_fill_1 FILLER_48_1473 ();
 sg13g2_fill_1 FILLER_48_1483 ();
 sg13g2_fill_1 FILLER_48_1489 ();
 sg13g2_fill_2 FILLER_48_1499 ();
 sg13g2_decap_8 FILLER_48_1546 ();
 sg13g2_fill_1 FILLER_48_1553 ();
 sg13g2_fill_1 FILLER_48_1563 ();
 sg13g2_fill_2 FILLER_48_1584 ();
 sg13g2_fill_2 FILLER_48_1598 ();
 sg13g2_fill_1 FILLER_48_1608 ();
 sg13g2_fill_1 FILLER_48_1614 ();
 sg13g2_decap_8 FILLER_48_1628 ();
 sg13g2_decap_8 FILLER_48_1635 ();
 sg13g2_decap_4 FILLER_48_1642 ();
 sg13g2_fill_1 FILLER_48_1646 ();
 sg13g2_fill_2 FILLER_48_1651 ();
 sg13g2_fill_2 FILLER_48_1657 ();
 sg13g2_fill_1 FILLER_48_1659 ();
 sg13g2_fill_2 FILLER_48_1663 ();
 sg13g2_fill_1 FILLER_48_1665 ();
 sg13g2_decap_4 FILLER_48_1670 ();
 sg13g2_fill_2 FILLER_48_1674 ();
 sg13g2_fill_1 FILLER_48_1685 ();
 sg13g2_fill_1 FILLER_48_1690 ();
 sg13g2_fill_2 FILLER_48_1696 ();
 sg13g2_fill_2 FILLER_48_1703 ();
 sg13g2_fill_1 FILLER_48_1739 ();
 sg13g2_fill_2 FILLER_48_1761 ();
 sg13g2_fill_1 FILLER_48_1782 ();
 sg13g2_fill_1 FILLER_48_1788 ();
 sg13g2_fill_2 FILLER_48_1817 ();
 sg13g2_decap_8 FILLER_48_1842 ();
 sg13g2_decap_8 FILLER_48_1849 ();
 sg13g2_decap_8 FILLER_48_1856 ();
 sg13g2_decap_8 FILLER_48_1863 ();
 sg13g2_decap_8 FILLER_48_1870 ();
 sg13g2_fill_2 FILLER_48_1877 ();
 sg13g2_fill_1 FILLER_48_1893 ();
 sg13g2_decap_8 FILLER_48_1922 ();
 sg13g2_decap_8 FILLER_48_1932 ();
 sg13g2_fill_1 FILLER_48_1943 ();
 sg13g2_fill_1 FILLER_48_1975 ();
 sg13g2_decap_8 FILLER_48_1981 ();
 sg13g2_decap_8 FILLER_48_1988 ();
 sg13g2_decap_8 FILLER_48_1995 ();
 sg13g2_fill_2 FILLER_48_2067 ();
 sg13g2_fill_1 FILLER_48_2069 ();
 sg13g2_decap_8 FILLER_48_2136 ();
 sg13g2_decap_4 FILLER_48_2143 ();
 sg13g2_fill_2 FILLER_48_2147 ();
 sg13g2_decap_8 FILLER_48_2201 ();
 sg13g2_decap_8 FILLER_48_2208 ();
 sg13g2_fill_1 FILLER_48_2215 ();
 sg13g2_fill_2 FILLER_48_2224 ();
 sg13g2_fill_2 FILLER_48_2236 ();
 sg13g2_fill_1 FILLER_48_2238 ();
 sg13g2_fill_1 FILLER_48_2249 ();
 sg13g2_decap_4 FILLER_48_2276 ();
 sg13g2_fill_2 FILLER_48_2318 ();
 sg13g2_fill_1 FILLER_48_2320 ();
 sg13g2_fill_2 FILLER_48_2325 ();
 sg13g2_fill_1 FILLER_48_2429 ();
 sg13g2_fill_1 FILLER_48_2519 ();
 sg13g2_fill_2 FILLER_48_2533 ();
 sg13g2_fill_1 FILLER_48_2551 ();
 sg13g2_fill_1 FILLER_48_2581 ();
 sg13g2_fill_1 FILLER_49_30 ();
 sg13g2_decap_4 FILLER_49_36 ();
 sg13g2_fill_1 FILLER_49_40 ();
 sg13g2_fill_2 FILLER_49_49 ();
 sg13g2_fill_1 FILLER_49_51 ();
 sg13g2_fill_1 FILLER_49_99 ();
 sg13g2_fill_2 FILLER_49_106 ();
 sg13g2_fill_2 FILLER_49_118 ();
 sg13g2_fill_2 FILLER_49_124 ();
 sg13g2_fill_2 FILLER_49_131 ();
 sg13g2_fill_1 FILLER_49_133 ();
 sg13g2_fill_2 FILLER_49_139 ();
 sg13g2_fill_1 FILLER_49_141 ();
 sg13g2_fill_2 FILLER_49_146 ();
 sg13g2_fill_1 FILLER_49_148 ();
 sg13g2_fill_1 FILLER_49_154 ();
 sg13g2_fill_2 FILLER_49_168 ();
 sg13g2_decap_4 FILLER_49_174 ();
 sg13g2_decap_8 FILLER_49_218 ();
 sg13g2_decap_8 FILLER_49_225 ();
 sg13g2_decap_4 FILLER_49_237 ();
 sg13g2_fill_1 FILLER_49_241 ();
 sg13g2_decap_4 FILLER_49_253 ();
 sg13g2_fill_1 FILLER_49_277 ();
 sg13g2_fill_2 FILLER_49_286 ();
 sg13g2_fill_2 FILLER_49_316 ();
 sg13g2_fill_1 FILLER_49_354 ();
 sg13g2_fill_2 FILLER_49_364 ();
 sg13g2_decap_4 FILLER_49_387 ();
 sg13g2_fill_2 FILLER_49_391 ();
 sg13g2_fill_1 FILLER_49_397 ();
 sg13g2_fill_1 FILLER_49_402 ();
 sg13g2_fill_1 FILLER_49_412 ();
 sg13g2_fill_2 FILLER_49_417 ();
 sg13g2_fill_1 FILLER_49_449 ();
 sg13g2_fill_1 FILLER_49_455 ();
 sg13g2_fill_2 FILLER_49_461 ();
 sg13g2_fill_1 FILLER_49_463 ();
 sg13g2_decap_4 FILLER_49_468 ();
 sg13g2_fill_1 FILLER_49_472 ();
 sg13g2_fill_2 FILLER_49_478 ();
 sg13g2_fill_1 FILLER_49_480 ();
 sg13g2_fill_2 FILLER_49_496 ();
 sg13g2_fill_1 FILLER_49_498 ();
 sg13g2_fill_2 FILLER_49_513 ();
 sg13g2_fill_2 FILLER_49_526 ();
 sg13g2_fill_2 FILLER_49_564 ();
 sg13g2_fill_1 FILLER_49_612 ();
 sg13g2_fill_1 FILLER_49_617 ();
 sg13g2_fill_2 FILLER_49_628 ();
 sg13g2_fill_2 FILLER_49_710 ();
 sg13g2_fill_1 FILLER_49_712 ();
 sg13g2_fill_2 FILLER_49_717 ();
 sg13g2_fill_1 FILLER_49_719 ();
 sg13g2_fill_1 FILLER_49_724 ();
 sg13g2_fill_2 FILLER_49_788 ();
 sg13g2_fill_2 FILLER_49_805 ();
 sg13g2_fill_1 FILLER_49_823 ();
 sg13g2_fill_2 FILLER_49_837 ();
 sg13g2_fill_2 FILLER_49_865 ();
 sg13g2_fill_1 FILLER_49_920 ();
 sg13g2_fill_1 FILLER_49_925 ();
 sg13g2_fill_2 FILLER_49_931 ();
 sg13g2_fill_1 FILLER_49_933 ();
 sg13g2_fill_1 FILLER_49_944 ();
 sg13g2_fill_1 FILLER_49_958 ();
 sg13g2_fill_1 FILLER_49_964 ();
 sg13g2_fill_1 FILLER_49_970 ();
 sg13g2_fill_2 FILLER_49_975 ();
 sg13g2_fill_1 FILLER_49_982 ();
 sg13g2_fill_2 FILLER_49_993 ();
 sg13g2_fill_1 FILLER_49_1000 ();
 sg13g2_fill_2 FILLER_49_1010 ();
 sg13g2_fill_1 FILLER_49_1012 ();
 sg13g2_fill_2 FILLER_49_1017 ();
 sg13g2_decap_8 FILLER_49_1028 ();
 sg13g2_fill_2 FILLER_49_1035 ();
 sg13g2_fill_1 FILLER_49_1037 ();
 sg13g2_decap_4 FILLER_49_1042 ();
 sg13g2_fill_1 FILLER_49_1056 ();
 sg13g2_fill_1 FILLER_49_1060 ();
 sg13g2_decap_4 FILLER_49_1066 ();
 sg13g2_fill_2 FILLER_49_1076 ();
 sg13g2_fill_1 FILLER_49_1078 ();
 sg13g2_fill_2 FILLER_49_1091 ();
 sg13g2_fill_1 FILLER_49_1153 ();
 sg13g2_fill_2 FILLER_49_1158 ();
 sg13g2_fill_2 FILLER_49_1170 ();
 sg13g2_fill_1 FILLER_49_1172 ();
 sg13g2_fill_2 FILLER_49_1199 ();
 sg13g2_fill_1 FILLER_49_1201 ();
 sg13g2_fill_2 FILLER_49_1228 ();
 sg13g2_decap_8 FILLER_49_1234 ();
 sg13g2_decap_8 FILLER_49_1241 ();
 sg13g2_fill_2 FILLER_49_1248 ();
 sg13g2_decap_8 FILLER_49_1254 ();
 sg13g2_decap_4 FILLER_49_1261 ();
 sg13g2_decap_4 FILLER_49_1275 ();
 sg13g2_fill_1 FILLER_49_1279 ();
 sg13g2_fill_1 FILLER_49_1290 ();
 sg13g2_fill_1 FILLER_49_1295 ();
 sg13g2_fill_2 FILLER_49_1301 ();
 sg13g2_fill_1 FILLER_49_1307 ();
 sg13g2_fill_1 FILLER_49_1312 ();
 sg13g2_fill_2 FILLER_49_1318 ();
 sg13g2_decap_8 FILLER_49_1325 ();
 sg13g2_decap_8 FILLER_49_1352 ();
 sg13g2_fill_1 FILLER_49_1359 ();
 sg13g2_fill_2 FILLER_49_1373 ();
 sg13g2_fill_1 FILLER_49_1385 ();
 sg13g2_decap_8 FILLER_49_1391 ();
 sg13g2_fill_2 FILLER_49_1398 ();
 sg13g2_fill_1 FILLER_49_1412 ();
 sg13g2_fill_2 FILLER_49_1418 ();
 sg13g2_decap_4 FILLER_49_1424 ();
 sg13g2_decap_8 FILLER_49_1442 ();
 sg13g2_decap_8 FILLER_49_1449 ();
 sg13g2_decap_4 FILLER_49_1456 ();
 sg13g2_fill_2 FILLER_49_1460 ();
 sg13g2_fill_1 FILLER_49_1470 ();
 sg13g2_decap_4 FILLER_49_1501 ();
 sg13g2_fill_2 FILLER_49_1505 ();
 sg13g2_fill_2 FILLER_49_1516 ();
 sg13g2_decap_4 FILLER_49_1535 ();
 sg13g2_fill_2 FILLER_49_1539 ();
 sg13g2_fill_1 FILLER_49_1560 ();
 sg13g2_decap_8 FILLER_49_1571 ();
 sg13g2_fill_1 FILLER_49_1578 ();
 sg13g2_decap_8 FILLER_49_1585 ();
 sg13g2_fill_1 FILLER_49_1611 ();
 sg13g2_decap_8 FILLER_49_1616 ();
 sg13g2_decap_4 FILLER_49_1623 ();
 sg13g2_fill_2 FILLER_49_1627 ();
 sg13g2_fill_2 FILLER_49_1655 ();
 sg13g2_decap_8 FILLER_49_1678 ();
 sg13g2_fill_1 FILLER_49_1685 ();
 sg13g2_fill_1 FILLER_49_1690 ();
 sg13g2_fill_2 FILLER_49_1695 ();
 sg13g2_fill_2 FILLER_49_1706 ();
 sg13g2_fill_2 FILLER_49_1721 ();
 sg13g2_fill_2 FILLER_49_1732 ();
 sg13g2_fill_2 FILLER_49_1756 ();
 sg13g2_fill_1 FILLER_49_1793 ();
 sg13g2_fill_1 FILLER_49_1802 ();
 sg13g2_fill_2 FILLER_49_1827 ();
 sg13g2_fill_1 FILLER_49_1829 ();
 sg13g2_decap_4 FILLER_49_1835 ();
 sg13g2_decap_8 FILLER_49_1850 ();
 sg13g2_decap_8 FILLER_49_1857 ();
 sg13g2_decap_8 FILLER_49_1864 ();
 sg13g2_decap_8 FILLER_49_1871 ();
 sg13g2_decap_4 FILLER_49_1878 ();
 sg13g2_fill_1 FILLER_49_1882 ();
 sg13g2_fill_2 FILLER_49_1922 ();
 sg13g2_decap_4 FILLER_49_1929 ();
 sg13g2_fill_1 FILLER_49_1933 ();
 sg13g2_fill_1 FILLER_49_1946 ();
 sg13g2_fill_1 FILLER_49_1951 ();
 sg13g2_fill_1 FILLER_49_1956 ();
 sg13g2_decap_8 FILLER_49_1961 ();
 sg13g2_decap_8 FILLER_49_1968 ();
 sg13g2_decap_4 FILLER_49_1975 ();
 sg13g2_fill_2 FILLER_49_1983 ();
 sg13g2_fill_2 FILLER_49_2056 ();
 sg13g2_fill_1 FILLER_49_2071 ();
 sg13g2_fill_2 FILLER_49_2080 ();
 sg13g2_decap_4 FILLER_49_2092 ();
 sg13g2_decap_4 FILLER_49_2117 ();
 sg13g2_decap_8 FILLER_49_2147 ();
 sg13g2_decap_4 FILLER_49_2154 ();
 sg13g2_fill_1 FILLER_49_2158 ();
 sg13g2_fill_2 FILLER_49_2183 ();
 sg13g2_fill_1 FILLER_49_2200 ();
 sg13g2_fill_2 FILLER_49_2245 ();
 sg13g2_fill_2 FILLER_49_2273 ();
 sg13g2_fill_1 FILLER_49_2275 ();
 sg13g2_fill_1 FILLER_49_2327 ();
 sg13g2_fill_2 FILLER_49_2333 ();
 sg13g2_fill_1 FILLER_49_2359 ();
 sg13g2_fill_1 FILLER_49_2393 ();
 sg13g2_fill_2 FILLER_49_2400 ();
 sg13g2_fill_2 FILLER_49_2450 ();
 sg13g2_fill_2 FILLER_49_2478 ();
 sg13g2_fill_1 FILLER_49_2499 ();
 sg13g2_fill_1 FILLER_49_2538 ();
 sg13g2_fill_2 FILLER_49_2556 ();
 sg13g2_fill_2 FILLER_49_2618 ();
 sg13g2_fill_2 FILLER_49_2640 ();
 sg13g2_fill_2 FILLER_49_2668 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_41 ();
 sg13g2_fill_2 FILLER_50_73 ();
 sg13g2_decap_8 FILLER_50_111 ();
 sg13g2_decap_8 FILLER_50_118 ();
 sg13g2_decap_4 FILLER_50_125 ();
 sg13g2_fill_1 FILLER_50_129 ();
 sg13g2_decap_8 FILLER_50_138 ();
 sg13g2_fill_2 FILLER_50_145 ();
 sg13g2_decap_4 FILLER_50_155 ();
 sg13g2_decap_8 FILLER_50_166 ();
 sg13g2_fill_2 FILLER_50_173 ();
 sg13g2_fill_2 FILLER_50_188 ();
 sg13g2_fill_1 FILLER_50_190 ();
 sg13g2_decap_8 FILLER_50_217 ();
 sg13g2_fill_1 FILLER_50_224 ();
 sg13g2_fill_1 FILLER_50_274 ();
 sg13g2_fill_2 FILLER_50_315 ();
 sg13g2_fill_1 FILLER_50_317 ();
 sg13g2_fill_1 FILLER_50_344 ();
 sg13g2_fill_1 FILLER_50_379 ();
 sg13g2_fill_1 FILLER_50_385 ();
 sg13g2_fill_2 FILLER_50_403 ();
 sg13g2_fill_1 FILLER_50_405 ();
 sg13g2_decap_4 FILLER_50_415 ();
 sg13g2_fill_1 FILLER_50_419 ();
 sg13g2_decap_4 FILLER_50_424 ();
 sg13g2_fill_2 FILLER_50_450 ();
 sg13g2_fill_1 FILLER_50_470 ();
 sg13g2_fill_1 FILLER_50_480 ();
 sg13g2_decap_8 FILLER_50_490 ();
 sg13g2_decap_8 FILLER_50_497 ();
 sg13g2_fill_1 FILLER_50_513 ();
 sg13g2_fill_1 FILLER_50_528 ();
 sg13g2_fill_2 FILLER_50_542 ();
 sg13g2_fill_1 FILLER_50_544 ();
 sg13g2_fill_1 FILLER_50_554 ();
 sg13g2_fill_2 FILLER_50_559 ();
 sg13g2_fill_1 FILLER_50_592 ();
 sg13g2_fill_2 FILLER_50_617 ();
 sg13g2_fill_2 FILLER_50_650 ();
 sg13g2_decap_8 FILLER_50_699 ();
 sg13g2_decap_8 FILLER_50_706 ();
 sg13g2_fill_1 FILLER_50_718 ();
 sg13g2_fill_2 FILLER_50_723 ();
 sg13g2_fill_1 FILLER_50_725 ();
 sg13g2_fill_2 FILLER_50_743 ();
 sg13g2_decap_4 FILLER_50_823 ();
 sg13g2_fill_2 FILLER_50_827 ();
 sg13g2_decap_8 FILLER_50_914 ();
 sg13g2_fill_1 FILLER_50_931 ();
 sg13g2_fill_2 FILLER_50_942 ();
 sg13g2_fill_1 FILLER_50_944 ();
 sg13g2_fill_2 FILLER_50_950 ();
 sg13g2_fill_1 FILLER_50_952 ();
 sg13g2_fill_2 FILLER_50_963 ();
 sg13g2_decap_8 FILLER_50_1005 ();
 sg13g2_decap_8 FILLER_50_1012 ();
 sg13g2_fill_2 FILLER_50_1029 ();
 sg13g2_fill_2 FILLER_50_1063 ();
 sg13g2_fill_1 FILLER_50_1124 ();
 sg13g2_fill_2 FILLER_50_1129 ();
 sg13g2_fill_1 FILLER_50_1169 ();
 sg13g2_fill_1 FILLER_50_1184 ();
 sg13g2_decap_8 FILLER_50_1220 ();
 sg13g2_fill_2 FILLER_50_1227 ();
 sg13g2_fill_1 FILLER_50_1229 ();
 sg13g2_decap_8 FILLER_50_1235 ();
 sg13g2_decap_4 FILLER_50_1242 ();
 sg13g2_fill_2 FILLER_50_1246 ();
 sg13g2_decap_8 FILLER_50_1252 ();
 sg13g2_decap_4 FILLER_50_1259 ();
 sg13g2_fill_2 FILLER_50_1263 ();
 sg13g2_fill_1 FILLER_50_1270 ();
 sg13g2_fill_1 FILLER_50_1275 ();
 sg13g2_fill_1 FILLER_50_1288 ();
 sg13g2_fill_1 FILLER_50_1318 ();
 sg13g2_decap_8 FILLER_50_1332 ();
 sg13g2_fill_1 FILLER_50_1339 ();
 sg13g2_decap_8 FILLER_50_1344 ();
 sg13g2_decap_8 FILLER_50_1351 ();
 sg13g2_fill_1 FILLER_50_1358 ();
 sg13g2_fill_2 FILLER_50_1376 ();
 sg13g2_fill_1 FILLER_50_1378 ();
 sg13g2_fill_1 FILLER_50_1384 ();
 sg13g2_fill_1 FILLER_50_1393 ();
 sg13g2_fill_2 FILLER_50_1415 ();
 sg13g2_decap_8 FILLER_50_1421 ();
 sg13g2_decap_8 FILLER_50_1443 ();
 sg13g2_fill_2 FILLER_50_1450 ();
 sg13g2_decap_8 FILLER_50_1456 ();
 sg13g2_fill_2 FILLER_50_1496 ();
 sg13g2_fill_2 FILLER_50_1537 ();
 sg13g2_fill_1 FILLER_50_1554 ();
 sg13g2_fill_1 FILLER_50_1577 ();
 sg13g2_decap_8 FILLER_50_1583 ();
 sg13g2_decap_8 FILLER_50_1590 ();
 sg13g2_fill_2 FILLER_50_1597 ();
 sg13g2_fill_1 FILLER_50_1599 ();
 sg13g2_decap_4 FILLER_50_1608 ();
 sg13g2_fill_2 FILLER_50_1612 ();
 sg13g2_decap_8 FILLER_50_1618 ();
 sg13g2_decap_8 FILLER_50_1625 ();
 sg13g2_fill_1 FILLER_50_1632 ();
 sg13g2_fill_1 FILLER_50_1641 ();
 sg13g2_fill_1 FILLER_50_1647 ();
 sg13g2_decap_4 FILLER_50_1653 ();
 sg13g2_decap_4 FILLER_50_1681 ();
 sg13g2_fill_2 FILLER_50_1697 ();
 sg13g2_fill_1 FILLER_50_1699 ();
 sg13g2_decap_8 FILLER_50_1704 ();
 sg13g2_fill_1 FILLER_50_1711 ();
 sg13g2_decap_8 FILLER_50_1726 ();
 sg13g2_decap_4 FILLER_50_1733 ();
 sg13g2_fill_1 FILLER_50_1737 ();
 sg13g2_fill_1 FILLER_50_1742 ();
 sg13g2_fill_2 FILLER_50_1763 ();
 sg13g2_fill_1 FILLER_50_1809 ();
 sg13g2_fill_2 FILLER_50_1842 ();
 sg13g2_fill_1 FILLER_50_1853 ();
 sg13g2_fill_2 FILLER_50_1859 ();
 sg13g2_fill_1 FILLER_50_1871 ();
 sg13g2_fill_1 FILLER_50_1876 ();
 sg13g2_fill_2 FILLER_50_1882 ();
 sg13g2_fill_1 FILLER_50_1884 ();
 sg13g2_fill_2 FILLER_50_1943 ();
 sg13g2_fill_1 FILLER_50_1963 ();
 sg13g2_fill_1 FILLER_50_1967 ();
 sg13g2_decap_8 FILLER_50_1972 ();
 sg13g2_decap_8 FILLER_50_1979 ();
 sg13g2_decap_8 FILLER_50_1986 ();
 sg13g2_decap_4 FILLER_50_1993 ();
 sg13g2_fill_1 FILLER_50_1997 ();
 sg13g2_decap_4 FILLER_50_2029 ();
 sg13g2_decap_8 FILLER_50_2062 ();
 sg13g2_fill_1 FILLER_50_2069 ();
 sg13g2_decap_8 FILLER_50_2096 ();
 sg13g2_fill_1 FILLER_50_2103 ();
 sg13g2_decap_4 FILLER_50_2186 ();
 sg13g2_fill_1 FILLER_50_2190 ();
 sg13g2_fill_1 FILLER_50_2252 ();
 sg13g2_decap_8 FILLER_50_2261 ();
 sg13g2_decap_8 FILLER_50_2272 ();
 sg13g2_fill_2 FILLER_50_2279 ();
 sg13g2_fill_1 FILLER_50_2288 ();
 sg13g2_fill_2 FILLER_50_2315 ();
 sg13g2_fill_2 FILLER_50_2347 ();
 sg13g2_fill_2 FILLER_50_2360 ();
 sg13g2_fill_2 FILLER_50_2450 ();
 sg13g2_fill_2 FILLER_50_2468 ();
 sg13g2_fill_1 FILLER_50_2487 ();
 sg13g2_fill_2 FILLER_50_2572 ();
 sg13g2_fill_1 FILLER_50_2581 ();
 sg13g2_fill_2 FILLER_50_2668 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_4 ();
 sg13g2_fill_1 FILLER_51_10 ();
 sg13g2_fill_1 FILLER_51_21 ();
 sg13g2_fill_1 FILLER_51_35 ();
 sg13g2_decap_4 FILLER_51_41 ();
 sg13g2_fill_1 FILLER_51_45 ();
 sg13g2_fill_2 FILLER_51_64 ();
 sg13g2_fill_2 FILLER_51_73 ();
 sg13g2_fill_2 FILLER_51_85 ();
 sg13g2_fill_1 FILLER_51_91 ();
 sg13g2_fill_1 FILLER_51_103 ();
 sg13g2_decap_8 FILLER_51_108 ();
 sg13g2_decap_8 FILLER_51_115 ();
 sg13g2_decap_8 FILLER_51_151 ();
 sg13g2_fill_1 FILLER_51_158 ();
 sg13g2_fill_2 FILLER_51_179 ();
 sg13g2_fill_2 FILLER_51_212 ();
 sg13g2_decap_4 FILLER_51_227 ();
 sg13g2_fill_2 FILLER_51_269 ();
 sg13g2_fill_2 FILLER_51_317 ();
 sg13g2_fill_2 FILLER_51_333 ();
 sg13g2_decap_4 FILLER_51_355 ();
 sg13g2_fill_2 FILLER_51_359 ();
 sg13g2_fill_2 FILLER_51_396 ();
 sg13g2_fill_2 FILLER_51_438 ();
 sg13g2_fill_1 FILLER_51_440 ();
 sg13g2_decap_8 FILLER_51_445 ();
 sg13g2_decap_4 FILLER_51_462 ();
 sg13g2_decap_4 FILLER_51_501 ();
 sg13g2_decap_4 FILLER_51_540 ();
 sg13g2_fill_1 FILLER_51_544 ();
 sg13g2_fill_1 FILLER_51_591 ();
 sg13g2_fill_2 FILLER_51_673 ();
 sg13g2_fill_2 FILLER_51_685 ();
 sg13g2_decap_8 FILLER_51_697 ();
 sg13g2_fill_2 FILLER_51_704 ();
 sg13g2_fill_1 FILLER_51_706 ();
 sg13g2_fill_2 FILLER_51_711 ();
 sg13g2_fill_1 FILLER_51_713 ();
 sg13g2_fill_2 FILLER_51_719 ();
 sg13g2_fill_1 FILLER_51_721 ();
 sg13g2_fill_1 FILLER_51_736 ();
 sg13g2_fill_2 FILLER_51_755 ();
 sg13g2_decap_8 FILLER_51_825 ();
 sg13g2_fill_1 FILLER_51_832 ();
 sg13g2_decap_8 FILLER_51_837 ();
 sg13g2_decap_8 FILLER_51_844 ();
 sg13g2_decap_8 FILLER_51_851 ();
 sg13g2_decap_4 FILLER_51_862 ();
 sg13g2_fill_1 FILLER_51_866 ();
 sg13g2_decap_4 FILLER_51_903 ();
 sg13g2_fill_1 FILLER_51_958 ();
 sg13g2_fill_2 FILLER_51_985 ();
 sg13g2_fill_1 FILLER_51_992 ();
 sg13g2_decap_8 FILLER_51_997 ();
 sg13g2_decap_4 FILLER_51_1004 ();
 sg13g2_fill_2 FILLER_51_1008 ();
 sg13g2_fill_1 FILLER_51_1046 ();
 sg13g2_fill_1 FILLER_51_1131 ();
 sg13g2_fill_1 FILLER_51_1158 ();
 sg13g2_fill_2 FILLER_51_1194 ();
 sg13g2_decap_8 FILLER_51_1257 ();
 sg13g2_fill_1 FILLER_51_1264 ();
 sg13g2_fill_2 FILLER_51_1303 ();
 sg13g2_fill_1 FILLER_51_1305 ();
 sg13g2_fill_2 FILLER_51_1329 ();
 sg13g2_fill_1 FILLER_51_1331 ();
 sg13g2_decap_8 FILLER_51_1337 ();
 sg13g2_decap_8 FILLER_51_1348 ();
 sg13g2_fill_1 FILLER_51_1355 ();
 sg13g2_fill_2 FILLER_51_1376 ();
 sg13g2_fill_1 FILLER_51_1404 ();
 sg13g2_fill_2 FILLER_51_1410 ();
 sg13g2_fill_1 FILLER_51_1447 ();
 sg13g2_decap_8 FILLER_51_1453 ();
 sg13g2_decap_4 FILLER_51_1460 ();
 sg13g2_fill_1 FILLER_51_1469 ();
 sg13g2_fill_2 FILLER_51_1502 ();
 sg13g2_fill_2 FILLER_51_1507 ();
 sg13g2_fill_1 FILLER_51_1509 ();
 sg13g2_decap_8 FILLER_51_1516 ();
 sg13g2_fill_1 FILLER_51_1523 ();
 sg13g2_fill_1 FILLER_51_1529 ();
 sg13g2_fill_2 FILLER_51_1542 ();
 sg13g2_fill_1 FILLER_51_1560 ();
 sg13g2_fill_1 FILLER_51_1571 ();
 sg13g2_fill_2 FILLER_51_1585 ();
 sg13g2_fill_2 FILLER_51_1591 ();
 sg13g2_fill_2 FILLER_51_1597 ();
 sg13g2_fill_1 FILLER_51_1604 ();
 sg13g2_fill_2 FILLER_51_1616 ();
 sg13g2_fill_2 FILLER_51_1644 ();
 sg13g2_fill_1 FILLER_51_1651 ();
 sg13g2_decap_8 FILLER_51_1656 ();
 sg13g2_decap_8 FILLER_51_1690 ();
 sg13g2_decap_8 FILLER_51_1697 ();
 sg13g2_decap_8 FILLER_51_1704 ();
 sg13g2_decap_8 FILLER_51_1711 ();
 sg13g2_decap_8 FILLER_51_1724 ();
 sg13g2_decap_4 FILLER_51_1731 ();
 sg13g2_decap_8 FILLER_51_1740 ();
 sg13g2_fill_1 FILLER_51_1747 ();
 sg13g2_decap_4 FILLER_51_1752 ();
 sg13g2_fill_1 FILLER_51_1756 ();
 sg13g2_fill_1 FILLER_51_1775 ();
 sg13g2_fill_1 FILLER_51_1783 ();
 sg13g2_fill_1 FILLER_51_1789 ();
 sg13g2_fill_2 FILLER_51_1831 ();
 sg13g2_fill_1 FILLER_51_1849 ();
 sg13g2_decap_4 FILLER_51_1854 ();
 sg13g2_fill_1 FILLER_51_1858 ();
 sg13g2_fill_2 FILLER_51_1871 ();
 sg13g2_fill_1 FILLER_51_1902 ();
 sg13g2_fill_2 FILLER_51_1920 ();
 sg13g2_fill_1 FILLER_51_1945 ();
 sg13g2_fill_1 FILLER_51_1958 ();
 sg13g2_decap_4 FILLER_51_2003 ();
 sg13g2_decap_4 FILLER_51_2011 ();
 sg13g2_fill_2 FILLER_51_2015 ();
 sg13g2_fill_2 FILLER_51_2046 ();
 sg13g2_fill_1 FILLER_51_2058 ();
 sg13g2_decap_8 FILLER_51_2099 ();
 sg13g2_decap_8 FILLER_51_2106 ();
 sg13g2_fill_2 FILLER_51_2113 ();
 sg13g2_fill_2 FILLER_51_2151 ();
 sg13g2_decap_4 FILLER_51_2157 ();
 sg13g2_fill_2 FILLER_51_2161 ();
 sg13g2_decap_8 FILLER_51_2171 ();
 sg13g2_decap_4 FILLER_51_2178 ();
 sg13g2_fill_2 FILLER_51_2182 ();
 sg13g2_fill_2 FILLER_51_2215 ();
 sg13g2_fill_2 FILLER_51_2243 ();
 sg13g2_fill_1 FILLER_51_2245 ();
 sg13g2_decap_8 FILLER_51_2293 ();
 sg13g2_fill_2 FILLER_51_2533 ();
 sg13g2_fill_1 FILLER_51_2608 ();
 sg13g2_fill_1 FILLER_51_2663 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_4 FILLER_52_56 ();
 sg13g2_fill_1 FILLER_52_60 ();
 sg13g2_fill_2 FILLER_52_65 ();
 sg13g2_fill_2 FILLER_52_101 ();
 sg13g2_fill_1 FILLER_52_133 ();
 sg13g2_fill_2 FILLER_52_190 ();
 sg13g2_fill_1 FILLER_52_196 ();
 sg13g2_fill_1 FILLER_52_201 ();
 sg13g2_decap_4 FILLER_52_206 ();
 sg13g2_decap_8 FILLER_52_227 ();
 sg13g2_fill_2 FILLER_52_257 ();
 sg13g2_fill_2 FILLER_52_283 ();
 sg13g2_fill_2 FILLER_52_307 ();
 sg13g2_fill_1 FILLER_52_309 ();
 sg13g2_decap_8 FILLER_52_330 ();
 sg13g2_decap_8 FILLER_52_337 ();
 sg13g2_decap_4 FILLER_52_344 ();
 sg13g2_fill_2 FILLER_52_348 ();
 sg13g2_decap_8 FILLER_52_360 ();
 sg13g2_fill_2 FILLER_52_367 ();
 sg13g2_decap_4 FILLER_52_378 ();
 sg13g2_fill_1 FILLER_52_387 ();
 sg13g2_fill_1 FILLER_52_393 ();
 sg13g2_decap_4 FILLER_52_398 ();
 sg13g2_fill_1 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_52_469 ();
 sg13g2_decap_8 FILLER_52_476 ();
 sg13g2_decap_8 FILLER_52_483 ();
 sg13g2_decap_8 FILLER_52_490 ();
 sg13g2_fill_2 FILLER_52_497 ();
 sg13g2_fill_1 FILLER_52_499 ();
 sg13g2_decap_4 FILLER_52_511 ();
 sg13g2_fill_1 FILLER_52_520 ();
 sg13g2_fill_1 FILLER_52_527 ();
 sg13g2_decap_4 FILLER_52_537 ();
 sg13g2_fill_2 FILLER_52_541 ();
 sg13g2_fill_2 FILLER_52_582 ();
 sg13g2_fill_1 FILLER_52_597 ();
 sg13g2_fill_2 FILLER_52_635 ();
 sg13g2_fill_1 FILLER_52_667 ();
 sg13g2_fill_1 FILLER_52_699 ();
 sg13g2_fill_2 FILLER_52_704 ();
 sg13g2_fill_1 FILLER_52_706 ();
 sg13g2_fill_1 FILLER_52_733 ();
 sg13g2_fill_2 FILLER_52_757 ();
 sg13g2_fill_1 FILLER_52_805 ();
 sg13g2_decap_4 FILLER_52_845 ();
 sg13g2_fill_2 FILLER_52_849 ();
 sg13g2_fill_1 FILLER_52_889 ();
 sg13g2_decap_8 FILLER_52_939 ();
 sg13g2_fill_2 FILLER_52_1033 ();
 sg13g2_fill_2 FILLER_52_1066 ();
 sg13g2_decap_8 FILLER_52_1072 ();
 sg13g2_decap_8 FILLER_52_1079 ();
 sg13g2_fill_2 FILLER_52_1086 ();
 sg13g2_fill_2 FILLER_52_1098 ();
 sg13g2_fill_1 FILLER_52_1100 ();
 sg13g2_fill_2 FILLER_52_1105 ();
 sg13g2_fill_1 FILLER_52_1107 ();
 sg13g2_decap_8 FILLER_52_1112 ();
 sg13g2_fill_1 FILLER_52_1119 ();
 sg13g2_fill_2 FILLER_52_1131 ();
 sg13g2_fill_1 FILLER_52_1149 ();
 sg13g2_fill_1 FILLER_52_1182 ();
 sg13g2_decap_8 FILLER_52_1214 ();
 sg13g2_fill_2 FILLER_52_1221 ();
 sg13g2_fill_2 FILLER_52_1232 ();
 sg13g2_decap_8 FILLER_52_1242 ();
 sg13g2_fill_2 FILLER_52_1249 ();
 sg13g2_fill_1 FILLER_52_1251 ();
 sg13g2_decap_4 FILLER_52_1264 ();
 sg13g2_fill_1 FILLER_52_1278 ();
 sg13g2_fill_1 FILLER_52_1283 ();
 sg13g2_fill_1 FILLER_52_1289 ();
 sg13g2_fill_1 FILLER_52_1304 ();
 sg13g2_fill_2 FILLER_52_1315 ();
 sg13g2_decap_8 FILLER_52_1333 ();
 sg13g2_fill_2 FILLER_52_1340 ();
 sg13g2_fill_2 FILLER_52_1364 ();
 sg13g2_fill_1 FILLER_52_1366 ();
 sg13g2_fill_1 FILLER_52_1372 ();
 sg13g2_fill_1 FILLER_52_1421 ();
 sg13g2_fill_1 FILLER_52_1428 ();
 sg13g2_fill_2 FILLER_52_1448 ();
 sg13g2_fill_1 FILLER_52_1499 ();
 sg13g2_fill_1 FILLER_52_1523 ();
 sg13g2_fill_2 FILLER_52_1532 ();
 sg13g2_fill_1 FILLER_52_1552 ();
 sg13g2_fill_1 FILLER_52_1561 ();
 sg13g2_fill_1 FILLER_52_1603 ();
 sg13g2_decap_8 FILLER_52_1609 ();
 sg13g2_decap_4 FILLER_52_1616 ();
 sg13g2_fill_2 FILLER_52_1620 ();
 sg13g2_fill_2 FILLER_52_1685 ();
 sg13g2_decap_8 FILLER_52_1692 ();
 sg13g2_decap_4 FILLER_52_1760 ();
 sg13g2_fill_2 FILLER_52_1764 ();
 sg13g2_fill_2 FILLER_52_1776 ();
 sg13g2_fill_1 FILLER_52_1811 ();
 sg13g2_fill_2 FILLER_52_1819 ();
 sg13g2_fill_2 FILLER_52_1825 ();
 sg13g2_fill_1 FILLER_52_1831 ();
 sg13g2_fill_1 FILLER_52_1860 ();
 sg13g2_fill_2 FILLER_52_1869 ();
 sg13g2_fill_2 FILLER_52_1875 ();
 sg13g2_fill_2 FILLER_52_1882 ();
 sg13g2_fill_1 FILLER_52_1894 ();
 sg13g2_fill_1 FILLER_52_1927 ();
 sg13g2_fill_1 FILLER_52_1942 ();
 sg13g2_decap_4 FILLER_52_1952 ();
 sg13g2_fill_1 FILLER_52_1956 ();
 sg13g2_decap_4 FILLER_52_1962 ();
 sg13g2_decap_8 FILLER_52_1977 ();
 sg13g2_fill_2 FILLER_52_1984 ();
 sg13g2_fill_1 FILLER_52_1986 ();
 sg13g2_decap_8 FILLER_52_1991 ();
 sg13g2_fill_2 FILLER_52_1998 ();
 sg13g2_fill_1 FILLER_52_2000 ();
 sg13g2_fill_1 FILLER_52_2037 ();
 sg13g2_fill_1 FILLER_52_2042 ();
 sg13g2_decap_8 FILLER_52_2053 ();
 sg13g2_decap_4 FILLER_52_2070 ();
 sg13g2_fill_2 FILLER_52_2078 ();
 sg13g2_fill_2 FILLER_52_2101 ();
 sg13g2_fill_2 FILLER_52_2129 ();
 sg13g2_fill_1 FILLER_52_2131 ();
 sg13g2_fill_1 FILLER_52_2136 ();
 sg13g2_decap_4 FILLER_52_2141 ();
 sg13g2_fill_2 FILLER_52_2145 ();
 sg13g2_decap_8 FILLER_52_2173 ();
 sg13g2_fill_1 FILLER_52_2180 ();
 sg13g2_fill_2 FILLER_52_2191 ();
 sg13g2_fill_1 FILLER_52_2224 ();
 sg13g2_decap_8 FILLER_52_2229 ();
 sg13g2_fill_2 FILLER_52_2236 ();
 sg13g2_decap_8 FILLER_52_2251 ();
 sg13g2_decap_8 FILLER_52_2258 ();
 sg13g2_decap_8 FILLER_52_2265 ();
 sg13g2_fill_1 FILLER_52_2272 ();
 sg13g2_fill_1 FILLER_52_2299 ();
 sg13g2_fill_1 FILLER_52_2310 ();
 sg13g2_decap_8 FILLER_52_2314 ();
 sg13g2_fill_1 FILLER_52_2321 ();
 sg13g2_fill_1 FILLER_52_2326 ();
 sg13g2_fill_1 FILLER_52_2331 ();
 sg13g2_fill_1 FILLER_52_2337 ();
 sg13g2_fill_1 FILLER_52_2342 ();
 sg13g2_fill_2 FILLER_52_2373 ();
 sg13g2_fill_2 FILLER_52_2382 ();
 sg13g2_fill_2 FILLER_52_2387 ();
 sg13g2_fill_2 FILLER_52_2403 ();
 sg13g2_fill_2 FILLER_52_2485 ();
 sg13g2_fill_1 FILLER_52_2516 ();
 sg13g2_fill_2 FILLER_52_2530 ();
 sg13g2_fill_2 FILLER_52_2537 ();
 sg13g2_fill_2 FILLER_52_2575 ();
 sg13g2_fill_1 FILLER_52_2669 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_13 ();
 sg13g2_decap_8 FILLER_53_18 ();
 sg13g2_decap_4 FILLER_53_25 ();
 sg13g2_fill_2 FILLER_53_46 ();
 sg13g2_fill_1 FILLER_53_48 ();
 sg13g2_fill_1 FILLER_53_79 ();
 sg13g2_fill_2 FILLER_53_111 ();
 sg13g2_fill_1 FILLER_53_113 ();
 sg13g2_decap_8 FILLER_53_118 ();
 sg13g2_fill_2 FILLER_53_125 ();
 sg13g2_fill_1 FILLER_53_131 ();
 sg13g2_fill_2 FILLER_53_136 ();
 sg13g2_fill_2 FILLER_53_143 ();
 sg13g2_fill_2 FILLER_53_150 ();
 sg13g2_fill_1 FILLER_53_156 ();
 sg13g2_fill_2 FILLER_53_160 ();
 sg13g2_fill_2 FILLER_53_166 ();
 sg13g2_fill_1 FILLER_53_168 ();
 sg13g2_fill_2 FILLER_53_174 ();
 sg13g2_fill_1 FILLER_53_176 ();
 sg13g2_fill_2 FILLER_53_181 ();
 sg13g2_decap_4 FILLER_53_188 ();
 sg13g2_fill_1 FILLER_53_192 ();
 sg13g2_fill_1 FILLER_53_201 ();
 sg13g2_decap_8 FILLER_53_206 ();
 sg13g2_fill_1 FILLER_53_213 ();
 sg13g2_fill_1 FILLER_53_229 ();
 sg13g2_decap_8 FILLER_53_256 ();
 sg13g2_decap_8 FILLER_53_263 ();
 sg13g2_fill_2 FILLER_53_302 ();
 sg13g2_fill_1 FILLER_53_304 ();
 sg13g2_fill_2 FILLER_53_315 ();
 sg13g2_fill_2 FILLER_53_321 ();
 sg13g2_fill_1 FILLER_53_323 ();
 sg13g2_fill_2 FILLER_53_334 ();
 sg13g2_fill_1 FILLER_53_336 ();
 sg13g2_fill_2 FILLER_53_363 ();
 sg13g2_fill_2 FILLER_53_401 ();
 sg13g2_fill_1 FILLER_53_403 ();
 sg13g2_fill_1 FILLER_53_430 ();
 sg13g2_fill_2 FILLER_53_454 ();
 sg13g2_fill_1 FILLER_53_461 ();
 sg13g2_decap_4 FILLER_53_467 ();
 sg13g2_fill_1 FILLER_53_471 ();
 sg13g2_decap_4 FILLER_53_478 ();
 sg13g2_fill_2 FILLER_53_482 ();
 sg13g2_fill_1 FILLER_53_493 ();
 sg13g2_fill_2 FILLER_53_552 ();
 sg13g2_fill_2 FILLER_53_580 ();
 sg13g2_fill_2 FILLER_53_603 ();
 sg13g2_fill_1 FILLER_53_614 ();
 sg13g2_fill_1 FILLER_53_623 ();
 sg13g2_fill_2 FILLER_53_636 ();
 sg13g2_fill_1 FILLER_53_648 ();
 sg13g2_fill_1 FILLER_53_658 ();
 sg13g2_fill_2 FILLER_53_663 ();
 sg13g2_fill_1 FILLER_53_678 ();
 sg13g2_fill_1 FILLER_53_695 ();
 sg13g2_fill_2 FILLER_53_706 ();
 sg13g2_fill_1 FILLER_53_713 ();
 sg13g2_fill_1 FILLER_53_718 ();
 sg13g2_fill_2 FILLER_53_739 ();
 sg13g2_fill_1 FILLER_53_751 ();
 sg13g2_fill_2 FILLER_53_808 ();
 sg13g2_fill_1 FILLER_53_884 ();
 sg13g2_decap_8 FILLER_53_893 ();
 sg13g2_decap_4 FILLER_53_900 ();
 sg13g2_fill_2 FILLER_53_928 ();
 sg13g2_decap_4 FILLER_53_940 ();
 sg13g2_fill_1 FILLER_53_948 ();
 sg13g2_fill_2 FILLER_53_965 ();
 sg13g2_fill_1 FILLER_53_967 ();
 sg13g2_decap_8 FILLER_53_991 ();
 sg13g2_decap_8 FILLER_53_998 ();
 sg13g2_decap_4 FILLER_53_1005 ();
 sg13g2_fill_1 FILLER_53_1009 ();
 sg13g2_decap_8 FILLER_53_1014 ();
 sg13g2_decap_8 FILLER_53_1021 ();
 sg13g2_fill_2 FILLER_53_1028 ();
 sg13g2_fill_2 FILLER_53_1057 ();
 sg13g2_fill_2 FILLER_53_1091 ();
 sg13g2_fill_1 FILLER_53_1093 ();
 sg13g2_fill_2 FILLER_53_1132 ();
 sg13g2_fill_1 FILLER_53_1142 ();
 sg13g2_decap_4 FILLER_53_1206 ();
 sg13g2_decap_8 FILLER_53_1240 ();
 sg13g2_fill_1 FILLER_53_1247 ();
 sg13g2_fill_2 FILLER_53_1279 ();
 sg13g2_fill_1 FILLER_53_1288 ();
 sg13g2_decap_4 FILLER_53_1300 ();
 sg13g2_decap_8 FILLER_53_1309 ();
 sg13g2_decap_8 FILLER_53_1316 ();
 sg13g2_fill_2 FILLER_53_1323 ();
 sg13g2_fill_2 FILLER_53_1334 ();
 sg13g2_decap_4 FILLER_53_1349 ();
 sg13g2_fill_1 FILLER_53_1353 ();
 sg13g2_fill_2 FILLER_53_1363 ();
 sg13g2_fill_1 FILLER_53_1365 ();
 sg13g2_fill_1 FILLER_53_1389 ();
 sg13g2_fill_1 FILLER_53_1395 ();
 sg13g2_fill_2 FILLER_53_1414 ();
 sg13g2_fill_2 FILLER_53_1431 ();
 sg13g2_fill_1 FILLER_53_1459 ();
 sg13g2_decap_4 FILLER_53_1502 ();
 sg13g2_decap_8 FILLER_53_1510 ();
 sg13g2_decap_8 FILLER_53_1517 ();
 sg13g2_fill_1 FILLER_53_1524 ();
 sg13g2_fill_1 FILLER_53_1554 ();
 sg13g2_fill_1 FILLER_53_1568 ();
 sg13g2_fill_1 FILLER_53_1617 ();
 sg13g2_fill_2 FILLER_53_1635 ();
 sg13g2_decap_8 FILLER_53_1650 ();
 sg13g2_decap_4 FILLER_53_1657 ();
 sg13g2_fill_1 FILLER_53_1661 ();
 sg13g2_fill_2 FILLER_53_1680 ();
 sg13g2_decap_8 FILLER_53_1694 ();
 sg13g2_fill_2 FILLER_53_1710 ();
 sg13g2_fill_1 FILLER_53_1712 ();
 sg13g2_decap_8 FILLER_53_1744 ();
 sg13g2_fill_1 FILLER_53_1761 ();
 sg13g2_decap_4 FILLER_53_1779 ();
 sg13g2_fill_1 FILLER_53_1783 ();
 sg13g2_fill_2 FILLER_53_1789 ();
 sg13g2_fill_2 FILLER_53_1797 ();
 sg13g2_fill_1 FILLER_53_1807 ();
 sg13g2_fill_2 FILLER_53_1812 ();
 sg13g2_fill_1 FILLER_53_1826 ();
 sg13g2_fill_1 FILLER_53_1847 ();
 sg13g2_fill_1 FILLER_53_1853 ();
 sg13g2_decap_4 FILLER_53_1860 ();
 sg13g2_fill_2 FILLER_53_1864 ();
 sg13g2_fill_2 FILLER_53_1883 ();
 sg13g2_fill_1 FILLER_53_1885 ();
 sg13g2_fill_1 FILLER_53_1891 ();
 sg13g2_fill_1 FILLER_53_1897 ();
 sg13g2_fill_1 FILLER_53_1903 ();
 sg13g2_fill_1 FILLER_53_1910 ();
 sg13g2_fill_1 FILLER_53_1944 ();
 sg13g2_fill_1 FILLER_53_1950 ();
 sg13g2_fill_1 FILLER_53_1956 ();
 sg13g2_fill_1 FILLER_53_1962 ();
 sg13g2_fill_1 FILLER_53_1968 ();
 sg13g2_decap_8 FILLER_53_1974 ();
 sg13g2_decap_8 FILLER_53_1981 ();
 sg13g2_decap_8 FILLER_53_1988 ();
 sg13g2_decap_4 FILLER_53_2009 ();
 sg13g2_fill_2 FILLER_53_2043 ();
 sg13g2_fill_2 FILLER_53_2050 ();
 sg13g2_decap_4 FILLER_53_2082 ();
 sg13g2_fill_1 FILLER_53_2112 ();
 sg13g2_decap_8 FILLER_53_2117 ();
 sg13g2_decap_4 FILLER_53_2124 ();
 sg13g2_fill_1 FILLER_53_2128 ();
 sg13g2_decap_8 FILLER_53_2142 ();
 sg13g2_fill_1 FILLER_53_2149 ();
 sg13g2_fill_2 FILLER_53_2160 ();
 sg13g2_decap_4 FILLER_53_2166 ();
 sg13g2_fill_1 FILLER_53_2170 ();
 sg13g2_decap_8 FILLER_53_2175 ();
 sg13g2_decap_8 FILLER_53_2182 ();
 sg13g2_decap_8 FILLER_53_2189 ();
 sg13g2_fill_1 FILLER_53_2196 ();
 sg13g2_decap_8 FILLER_53_2223 ();
 sg13g2_decap_4 FILLER_53_2230 ();
 sg13g2_fill_2 FILLER_53_2254 ();
 sg13g2_fill_2 FILLER_53_2307 ();
 sg13g2_decap_4 FILLER_53_2314 ();
 sg13g2_fill_1 FILLER_53_2318 ();
 sg13g2_decap_4 FILLER_53_2323 ();
 sg13g2_fill_2 FILLER_53_2327 ();
 sg13g2_decap_8 FILLER_53_2333 ();
 sg13g2_decap_4 FILLER_53_2340 ();
 sg13g2_fill_1 FILLER_53_2344 ();
 sg13g2_fill_1 FILLER_53_2356 ();
 sg13g2_fill_2 FILLER_53_2360 ();
 sg13g2_fill_1 FILLER_53_2426 ();
 sg13g2_fill_2 FILLER_53_2473 ();
 sg13g2_fill_1 FILLER_53_2497 ();
 sg13g2_fill_2 FILLER_53_2528 ();
 sg13g2_fill_1 FILLER_53_2549 ();
 sg13g2_fill_2 FILLER_53_2554 ();
 sg13g2_fill_2 FILLER_53_2616 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_2 ();
 sg13g2_decap_4 FILLER_54_29 ();
 sg13g2_fill_1 FILLER_54_33 ();
 sg13g2_fill_1 FILLER_54_97 ();
 sg13g2_fill_1 FILLER_54_103 ();
 sg13g2_decap_8 FILLER_54_108 ();
 sg13g2_decap_8 FILLER_54_115 ();
 sg13g2_decap_8 FILLER_54_122 ();
 sg13g2_decap_8 FILLER_54_129 ();
 sg13g2_decap_8 FILLER_54_136 ();
 sg13g2_fill_1 FILLER_54_143 ();
 sg13g2_fill_1 FILLER_54_152 ();
 sg13g2_fill_1 FILLER_54_158 ();
 sg13g2_fill_1 FILLER_54_163 ();
 sg13g2_decap_8 FILLER_54_169 ();
 sg13g2_decap_8 FILLER_54_176 ();
 sg13g2_fill_2 FILLER_54_198 ();
 sg13g2_fill_1 FILLER_54_200 ();
 sg13g2_fill_2 FILLER_54_210 ();
 sg13g2_fill_1 FILLER_54_212 ();
 sg13g2_decap_8 FILLER_54_323 ();
 sg13g2_decap_8 FILLER_54_330 ();
 sg13g2_fill_1 FILLER_54_360 ();
 sg13g2_decap_8 FILLER_54_391 ();
 sg13g2_decap_8 FILLER_54_398 ();
 sg13g2_fill_1 FILLER_54_405 ();
 sg13g2_fill_1 FILLER_54_410 ();
 sg13g2_fill_2 FILLER_54_420 ();
 sg13g2_fill_2 FILLER_54_428 ();
 sg13g2_fill_1 FILLER_54_476 ();
 sg13g2_fill_2 FILLER_54_486 ();
 sg13g2_fill_1 FILLER_54_488 ();
 sg13g2_fill_1 FILLER_54_497 ();
 sg13g2_fill_2 FILLER_54_532 ();
 sg13g2_fill_2 FILLER_54_542 ();
 sg13g2_fill_1 FILLER_54_544 ();
 sg13g2_fill_1 FILLER_54_550 ();
 sg13g2_fill_2 FILLER_54_592 ();
 sg13g2_fill_2 FILLER_54_637 ();
 sg13g2_fill_1 FILLER_54_639 ();
 sg13g2_fill_2 FILLER_54_644 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_decap_8 FILLER_54_659 ();
 sg13g2_decap_8 FILLER_54_666 ();
 sg13g2_decap_8 FILLER_54_673 ();
 sg13g2_decap_4 FILLER_54_680 ();
 sg13g2_fill_2 FILLER_54_701 ();
 sg13g2_fill_1 FILLER_54_743 ();
 sg13g2_fill_1 FILLER_54_753 ();
 sg13g2_fill_2 FILLER_54_767 ();
 sg13g2_fill_1 FILLER_54_795 ();
 sg13g2_fill_1 FILLER_54_819 ();
 sg13g2_fill_1 FILLER_54_827 ();
 sg13g2_decap_4 FILLER_54_854 ();
 sg13g2_fill_1 FILLER_54_907 ();
 sg13g2_fill_2 FILLER_54_913 ();
 sg13g2_fill_1 FILLER_54_941 ();
 sg13g2_fill_1 FILLER_54_948 ();
 sg13g2_fill_2 FILLER_54_952 ();
 sg13g2_decap_8 FILLER_54_966 ();
 sg13g2_decap_8 FILLER_54_973 ();
 sg13g2_fill_2 FILLER_54_980 ();
 sg13g2_fill_1 FILLER_54_982 ();
 sg13g2_decap_8 FILLER_54_997 ();
 sg13g2_decap_8 FILLER_54_1004 ();
 sg13g2_decap_8 FILLER_54_1011 ();
 sg13g2_decap_4 FILLER_54_1018 ();
 sg13g2_fill_1 FILLER_54_1022 ();
 sg13g2_fill_2 FILLER_54_1049 ();
 sg13g2_fill_2 FILLER_54_1102 ();
 sg13g2_decap_4 FILLER_54_1108 ();
 sg13g2_fill_2 FILLER_54_1153 ();
 sg13g2_fill_1 FILLER_54_1155 ();
 sg13g2_fill_1 FILLER_54_1182 ();
 sg13g2_fill_1 FILLER_54_1209 ();
 sg13g2_fill_1 FILLER_54_1214 ();
 sg13g2_decap_8 FILLER_54_1230 ();
 sg13g2_fill_2 FILLER_54_1237 ();
 sg13g2_decap_4 FILLER_54_1277 ();
 sg13g2_fill_1 FILLER_54_1281 ();
 sg13g2_decap_8 FILLER_54_1305 ();
 sg13g2_decap_8 FILLER_54_1312 ();
 sg13g2_decap_4 FILLER_54_1319 ();
 sg13g2_fill_1 FILLER_54_1323 ();
 sg13g2_decap_8 FILLER_54_1334 ();
 sg13g2_fill_2 FILLER_54_1341 ();
 sg13g2_fill_1 FILLER_54_1352 ();
 sg13g2_decap_8 FILLER_54_1358 ();
 sg13g2_fill_1 FILLER_54_1365 ();
 sg13g2_decap_4 FILLER_54_1371 ();
 sg13g2_fill_2 FILLER_54_1375 ();
 sg13g2_decap_4 FILLER_54_1386 ();
 sg13g2_fill_1 FILLER_54_1414 ();
 sg13g2_fill_2 FILLER_54_1439 ();
 sg13g2_decap_8 FILLER_54_1450 ();
 sg13g2_fill_2 FILLER_54_1457 ();
 sg13g2_decap_4 FILLER_54_1472 ();
 sg13g2_fill_1 FILLER_54_1476 ();
 sg13g2_fill_1 FILLER_54_1480 ();
 sg13g2_decap_8 FILLER_54_1485 ();
 sg13g2_fill_2 FILLER_54_1492 ();
 sg13g2_decap_8 FILLER_54_1499 ();
 sg13g2_decap_8 FILLER_54_1506 ();
 sg13g2_fill_1 FILLER_54_1513 ();
 sg13g2_decap_8 FILLER_54_1518 ();
 sg13g2_fill_2 FILLER_54_1525 ();
 sg13g2_fill_1 FILLER_54_1527 ();
 sg13g2_fill_2 FILLER_54_1532 ();
 sg13g2_fill_1 FILLER_54_1538 ();
 sg13g2_fill_1 FILLER_54_1564 ();
 sg13g2_fill_1 FILLER_54_1579 ();
 sg13g2_fill_1 FILLER_54_1636 ();
 sg13g2_decap_8 FILLER_54_1650 ();
 sg13g2_decap_4 FILLER_54_1657 ();
 sg13g2_decap_8 FILLER_54_1676 ();
 sg13g2_decap_8 FILLER_54_1683 ();
 sg13g2_decap_4 FILLER_54_1690 ();
 sg13g2_fill_2 FILLER_54_1694 ();
 sg13g2_decap_8 FILLER_54_1716 ();
 sg13g2_decap_4 FILLER_54_1723 ();
 sg13g2_fill_2 FILLER_54_1727 ();
 sg13g2_fill_2 FILLER_54_1740 ();
 sg13g2_fill_1 FILLER_54_1742 ();
 sg13g2_decap_8 FILLER_54_1749 ();
 sg13g2_decap_4 FILLER_54_1756 ();
 sg13g2_decap_8 FILLER_54_1798 ();
 sg13g2_decap_4 FILLER_54_1805 ();
 sg13g2_fill_2 FILLER_54_1816 ();
 sg13g2_fill_1 FILLER_54_1851 ();
 sg13g2_fill_2 FILLER_54_1863 ();
 sg13g2_fill_2 FILLER_54_1870 ();
 sg13g2_fill_1 FILLER_54_1877 ();
 sg13g2_fill_1 FILLER_54_1899 ();
 sg13g2_fill_1 FILLER_54_1904 ();
 sg13g2_fill_1 FILLER_54_1910 ();
 sg13g2_fill_1 FILLER_54_1932 ();
 sg13g2_fill_1 FILLER_54_1938 ();
 sg13g2_fill_1 FILLER_54_1947 ();
 sg13g2_fill_1 FILLER_54_1957 ();
 sg13g2_fill_1 FILLER_54_1971 ();
 sg13g2_fill_1 FILLER_54_1983 ();
 sg13g2_fill_2 FILLER_54_1994 ();
 sg13g2_fill_1 FILLER_54_2004 ();
 sg13g2_decap_8 FILLER_54_2008 ();
 sg13g2_fill_2 FILLER_54_2015 ();
 sg13g2_decap_8 FILLER_54_2025 ();
 sg13g2_decap_8 FILLER_54_2032 ();
 sg13g2_decap_4 FILLER_54_2039 ();
 sg13g2_fill_1 FILLER_54_2043 ();
 sg13g2_decap_4 FILLER_54_2054 ();
 sg13g2_fill_1 FILLER_54_2058 ();
 sg13g2_decap_8 FILLER_54_2079 ();
 sg13g2_fill_2 FILLER_54_2086 ();
 sg13g2_fill_2 FILLER_54_2147 ();
 sg13g2_fill_1 FILLER_54_2149 ();
 sg13g2_fill_1 FILLER_54_2181 ();
 sg13g2_decap_8 FILLER_54_2186 ();
 sg13g2_decap_8 FILLER_54_2193 ();
 sg13g2_fill_2 FILLER_54_2200 ();
 sg13g2_fill_1 FILLER_54_2202 ();
 sg13g2_fill_2 FILLER_54_2243 ();
 sg13g2_fill_1 FILLER_54_2245 ();
 sg13g2_decap_8 FILLER_54_2283 ();
 sg13g2_decap_4 FILLER_54_2290 ();
 sg13g2_fill_2 FILLER_54_2294 ();
 sg13g2_fill_1 FILLER_54_2308 ();
 sg13g2_fill_2 FILLER_54_2343 ();
 sg13g2_fill_1 FILLER_54_2348 ();
 sg13g2_fill_1 FILLER_54_2353 ();
 sg13g2_fill_2 FILLER_54_2369 ();
 sg13g2_fill_1 FILLER_54_2384 ();
 sg13g2_fill_2 FILLER_54_2447 ();
 sg13g2_fill_1 FILLER_54_2455 ();
 sg13g2_fill_1 FILLER_54_2482 ();
 sg13g2_fill_2 FILLER_54_2487 ();
 sg13g2_fill_1 FILLER_54_2496 ();
 sg13g2_fill_1 FILLER_54_2523 ();
 sg13g2_fill_2 FILLER_54_2565 ();
 sg13g2_fill_2 FILLER_54_2646 ();
 sg13g2_fill_2 FILLER_54_2659 ();
 sg13g2_fill_1 FILLER_54_2664 ();
 sg13g2_fill_2 FILLER_54_2668 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_4 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_11 ();
 sg13g2_fill_2 FILLER_55_52 ();
 sg13g2_decap_8 FILLER_55_59 ();
 sg13g2_decap_8 FILLER_55_66 ();
 sg13g2_decap_4 FILLER_55_73 ();
 sg13g2_fill_1 FILLER_55_77 ();
 sg13g2_fill_1 FILLER_55_99 ();
 sg13g2_decap_4 FILLER_55_126 ();
 sg13g2_fill_2 FILLER_55_130 ();
 sg13g2_fill_1 FILLER_55_145 ();
 sg13g2_fill_1 FILLER_55_151 ();
 sg13g2_fill_1 FILLER_55_162 ();
 sg13g2_fill_2 FILLER_55_189 ();
 sg13g2_decap_8 FILLER_55_249 ();
 sg13g2_fill_1 FILLER_55_256 ();
 sg13g2_decap_4 FILLER_55_261 ();
 sg13g2_fill_1 FILLER_55_265 ();
 sg13g2_decap_8 FILLER_55_274 ();
 sg13g2_decap_4 FILLER_55_281 ();
 sg13g2_fill_2 FILLER_55_289 ();
 sg13g2_fill_1 FILLER_55_299 ();
 sg13g2_fill_1 FILLER_55_304 ();
 sg13g2_fill_1 FILLER_55_331 ();
 sg13g2_fill_1 FILLER_55_377 ();
 sg13g2_decap_8 FILLER_55_382 ();
 sg13g2_fill_1 FILLER_55_389 ();
 sg13g2_fill_1 FILLER_55_395 ();
 sg13g2_decap_8 FILLER_55_408 ();
 sg13g2_fill_1 FILLER_55_457 ();
 sg13g2_fill_1 FILLER_55_501 ();
 sg13g2_fill_1 FILLER_55_512 ();
 sg13g2_fill_1 FILLER_55_521 ();
 sg13g2_fill_2 FILLER_55_541 ();
 sg13g2_fill_1 FILLER_55_557 ();
 sg13g2_fill_1 FILLER_55_638 ();
 sg13g2_fill_1 FILLER_55_674 ();
 sg13g2_decap_8 FILLER_55_679 ();
 sg13g2_decap_8 FILLER_55_686 ();
 sg13g2_decap_4 FILLER_55_693 ();
 sg13g2_fill_1 FILLER_55_697 ();
 sg13g2_fill_1 FILLER_55_744 ();
 sg13g2_fill_1 FILLER_55_749 ();
 sg13g2_fill_1 FILLER_55_762 ();
 sg13g2_fill_1 FILLER_55_771 ();
 sg13g2_fill_2 FILLER_55_787 ();
 sg13g2_fill_1 FILLER_55_795 ();
 sg13g2_fill_1 FILLER_55_829 ();
 sg13g2_decap_8 FILLER_55_849 ();
 sg13g2_decap_4 FILLER_55_856 ();
 sg13g2_fill_1 FILLER_55_860 ();
 sg13g2_fill_1 FILLER_55_865 ();
 sg13g2_fill_1 FILLER_55_870 ();
 sg13g2_fill_2 FILLER_55_949 ();
 sg13g2_fill_1 FILLER_55_956 ();
 sg13g2_fill_2 FILLER_55_960 ();
 sg13g2_fill_1 FILLER_55_962 ();
 sg13g2_decap_4 FILLER_55_971 ();
 sg13g2_fill_2 FILLER_55_979 ();
 sg13g2_fill_1 FILLER_55_981 ();
 sg13g2_decap_4 FILLER_55_1008 ();
 sg13g2_decap_8 FILLER_55_1017 ();
 sg13g2_fill_1 FILLER_55_1083 ();
 sg13g2_fill_2 FILLER_55_1088 ();
 sg13g2_fill_1 FILLER_55_1100 ();
 sg13g2_decap_8 FILLER_55_1127 ();
 sg13g2_decap_8 FILLER_55_1134 ();
 sg13g2_fill_2 FILLER_55_1141 ();
 sg13g2_fill_1 FILLER_55_1182 ();
 sg13g2_fill_2 FILLER_55_1187 ();
 sg13g2_fill_2 FILLER_55_1193 ();
 sg13g2_fill_2 FILLER_55_1205 ();
 sg13g2_fill_1 FILLER_55_1207 ();
 sg13g2_decap_8 FILLER_55_1212 ();
 sg13g2_decap_4 FILLER_55_1219 ();
 sg13g2_fill_2 FILLER_55_1223 ();
 sg13g2_fill_2 FILLER_55_1230 ();
 sg13g2_fill_1 FILLER_55_1232 ();
 sg13g2_fill_2 FILLER_55_1238 ();
 sg13g2_decap_4 FILLER_55_1275 ();
 sg13g2_decap_8 FILLER_55_1297 ();
 sg13g2_decap_8 FILLER_55_1304 ();
 sg13g2_decap_4 FILLER_55_1311 ();
 sg13g2_decap_4 FILLER_55_1319 ();
 sg13g2_fill_2 FILLER_55_1323 ();
 sg13g2_decap_4 FILLER_55_1334 ();
 sg13g2_fill_2 FILLER_55_1338 ();
 sg13g2_decap_4 FILLER_55_1354 ();
 sg13g2_fill_2 FILLER_55_1429 ();
 sg13g2_fill_2 FILLER_55_1440 ();
 sg13g2_fill_1 FILLER_55_1442 ();
 sg13g2_decap_8 FILLER_55_1451 ();
 sg13g2_decap_8 FILLER_55_1458 ();
 sg13g2_fill_2 FILLER_55_1465 ();
 sg13g2_decap_4 FILLER_55_1507 ();
 sg13g2_decap_4 FILLER_55_1519 ();
 sg13g2_fill_1 FILLER_55_1574 ();
 sg13g2_fill_2 FILLER_55_1596 ();
 sg13g2_fill_1 FILLER_55_1618 ();
 sg13g2_fill_2 FILLER_55_1630 ();
 sg13g2_decap_8 FILLER_55_1639 ();
 sg13g2_decap_4 FILLER_55_1646 ();
 sg13g2_decap_8 FILLER_55_1678 ();
 sg13g2_decap_8 FILLER_55_1685 ();
 sg13g2_decap_4 FILLER_55_1696 ();
 sg13g2_fill_1 FILLER_55_1700 ();
 sg13g2_decap_8 FILLER_55_1704 ();
 sg13g2_fill_2 FILLER_55_1716 ();
 sg13g2_fill_1 FILLER_55_1718 ();
 sg13g2_decap_4 FILLER_55_1723 ();
 sg13g2_fill_2 FILLER_55_1754 ();
 sg13g2_fill_1 FILLER_55_1756 ();
 sg13g2_fill_1 FILLER_55_1773 ();
 sg13g2_fill_1 FILLER_55_1779 ();
 sg13g2_fill_1 FILLER_55_1791 ();
 sg13g2_decap_8 FILLER_55_1797 ();
 sg13g2_fill_2 FILLER_55_1804 ();
 sg13g2_fill_1 FILLER_55_1818 ();
 sg13g2_fill_2 FILLER_55_1829 ();
 sg13g2_fill_2 FILLER_55_1841 ();
 sg13g2_fill_1 FILLER_55_1848 ();
 sg13g2_fill_2 FILLER_55_1863 ();
 sg13g2_fill_1 FILLER_55_1873 ();
 sg13g2_fill_1 FILLER_55_1889 ();
 sg13g2_fill_1 FILLER_55_1898 ();
 sg13g2_fill_1 FILLER_55_1933 ();
 sg13g2_fill_1 FILLER_55_1944 ();
 sg13g2_fill_1 FILLER_55_1950 ();
 sg13g2_decap_8 FILLER_55_1956 ();
 sg13g2_fill_2 FILLER_55_1963 ();
 sg13g2_fill_1 FILLER_55_1977 ();
 sg13g2_fill_2 FILLER_55_1996 ();
 sg13g2_fill_1 FILLER_55_1998 ();
 sg13g2_fill_1 FILLER_55_2004 ();
 sg13g2_decap_4 FILLER_55_2021 ();
 sg13g2_fill_1 FILLER_55_2025 ();
 sg13g2_decap_8 FILLER_55_2068 ();
 sg13g2_decap_4 FILLER_55_2075 ();
 sg13g2_fill_1 FILLER_55_2079 ();
 sg13g2_fill_2 FILLER_55_2112 ();
 sg13g2_fill_2 FILLER_55_2166 ();
 sg13g2_fill_2 FILLER_55_2189 ();
 sg13g2_decap_4 FILLER_55_2238 ();
 sg13g2_fill_1 FILLER_55_2242 ();
 sg13g2_fill_2 FILLER_55_2264 ();
 sg13g2_fill_1 FILLER_55_2266 ();
 sg13g2_fill_1 FILLER_55_2339 ();
 sg13g2_fill_2 FILLER_55_2348 ();
 sg13g2_fill_1 FILLER_55_2359 ();
 sg13g2_fill_1 FILLER_55_2367 ();
 sg13g2_fill_1 FILLER_55_2389 ();
 sg13g2_fill_1 FILLER_55_2400 ();
 sg13g2_fill_2 FILLER_55_2409 ();
 sg13g2_fill_1 FILLER_55_2415 ();
 sg13g2_fill_1 FILLER_55_2422 ();
 sg13g2_fill_1 FILLER_55_2427 ();
 sg13g2_fill_1 FILLER_55_2437 ();
 sg13g2_fill_2 FILLER_55_2451 ();
 sg13g2_fill_2 FILLER_55_2479 ();
 sg13g2_fill_2 FILLER_55_2539 ();
 sg13g2_fill_2 FILLER_55_2569 ();
 sg13g2_fill_2 FILLER_55_2584 ();
 sg13g2_fill_1 FILLER_55_2590 ();
 sg13g2_fill_1 FILLER_55_2601 ();
 sg13g2_fill_1 FILLER_55_2612 ();
 sg13g2_fill_1 FILLER_55_2617 ();
 sg13g2_fill_1 FILLER_55_2628 ();
 sg13g2_fill_1 FILLER_55_2655 ();
 sg13g2_fill_1 FILLER_55_2663 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_4 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_11 ();
 sg13g2_fill_2 FILLER_56_29 ();
 sg13g2_fill_1 FILLER_56_31 ();
 sg13g2_decap_4 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_57 ();
 sg13g2_decap_4 FILLER_56_64 ();
 sg13g2_fill_1 FILLER_56_68 ();
 sg13g2_fill_2 FILLER_56_77 ();
 sg13g2_fill_1 FILLER_56_84 ();
 sg13g2_fill_2 FILLER_56_115 ();
 sg13g2_fill_2 FILLER_56_120 ();
 sg13g2_fill_1 FILLER_56_148 ();
 sg13g2_fill_1 FILLER_56_153 ();
 sg13g2_fill_2 FILLER_56_164 ();
 sg13g2_fill_1 FILLER_56_171 ();
 sg13g2_fill_2 FILLER_56_176 ();
 sg13g2_fill_2 FILLER_56_251 ();
 sg13g2_decap_8 FILLER_56_288 ();
 sg13g2_fill_1 FILLER_56_295 ();
 sg13g2_decap_4 FILLER_56_301 ();
 sg13g2_fill_2 FILLER_56_305 ();
 sg13g2_decap_8 FILLER_56_311 ();
 sg13g2_decap_8 FILLER_56_322 ();
 sg13g2_decap_8 FILLER_56_329 ();
 sg13g2_decap_4 FILLER_56_336 ();
 sg13g2_fill_1 FILLER_56_340 ();
 sg13g2_fill_2 FILLER_56_345 ();
 sg13g2_fill_2 FILLER_56_351 ();
 sg13g2_decap_8 FILLER_56_357 ();
 sg13g2_decap_8 FILLER_56_364 ();
 sg13g2_fill_1 FILLER_56_371 ();
 sg13g2_decap_4 FILLER_56_376 ();
 sg13g2_fill_1 FILLER_56_426 ();
 sg13g2_fill_2 FILLER_56_459 ();
 sg13g2_fill_2 FILLER_56_523 ();
 sg13g2_fill_2 FILLER_56_531 ();
 sg13g2_fill_1 FILLER_56_533 ();
 sg13g2_fill_2 FILLER_56_572 ();
 sg13g2_fill_2 FILLER_56_664 ();
 sg13g2_fill_2 FILLER_56_697 ();
 sg13g2_fill_1 FILLER_56_716 ();
 sg13g2_fill_1 FILLER_56_739 ();
 sg13g2_fill_1 FILLER_56_748 ();
 sg13g2_fill_2 FILLER_56_757 ();
 sg13g2_fill_2 FILLER_56_764 ();
 sg13g2_fill_1 FILLER_56_798 ();
 sg13g2_fill_2 FILLER_56_807 ();
 sg13g2_decap_8 FILLER_56_851 ();
 sg13g2_fill_2 FILLER_56_858 ();
 sg13g2_fill_1 FILLER_56_860 ();
 sg13g2_fill_1 FILLER_56_883 ();
 sg13g2_fill_1 FILLER_56_890 ();
 sg13g2_fill_2 FILLER_56_901 ();
 sg13g2_fill_2 FILLER_56_907 ();
 sg13g2_fill_2 FILLER_56_914 ();
 sg13g2_fill_2 FILLER_56_928 ();
 sg13g2_fill_1 FILLER_56_930 ();
 sg13g2_fill_1 FILLER_56_967 ();
 sg13g2_fill_2 FILLER_56_1016 ();
 sg13g2_decap_8 FILLER_56_1022 ();
 sg13g2_decap_8 FILLER_56_1029 ();
 sg13g2_fill_2 FILLER_56_1036 ();
 sg13g2_fill_2 FILLER_56_1062 ();
 sg13g2_decap_4 FILLER_56_1081 ();
 sg13g2_fill_2 FILLER_56_1085 ();
 sg13g2_fill_2 FILLER_56_1133 ();
 sg13g2_fill_1 FILLER_56_1135 ();
 sg13g2_decap_8 FILLER_56_1140 ();
 sg13g2_decap_8 FILLER_56_1147 ();
 sg13g2_decap_4 FILLER_56_1154 ();
 sg13g2_fill_1 FILLER_56_1168 ();
 sg13g2_decap_8 FILLER_56_1173 ();
 sg13g2_fill_2 FILLER_56_1194 ();
 sg13g2_fill_2 FILLER_56_1248 ();
 sg13g2_fill_2 FILLER_56_1258 ();
 sg13g2_fill_2 FILLER_56_1265 ();
 sg13g2_fill_1 FILLER_56_1273 ();
 sg13g2_fill_2 FILLER_56_1279 ();
 sg13g2_fill_1 FILLER_56_1286 ();
 sg13g2_fill_1 FILLER_56_1292 ();
 sg13g2_decap_4 FILLER_56_1297 ();
 sg13g2_fill_2 FILLER_56_1301 ();
 sg13g2_decap_4 FILLER_56_1307 ();
 sg13g2_fill_1 FILLER_56_1311 ();
 sg13g2_decap_4 FILLER_56_1332 ();
 sg13g2_fill_1 FILLER_56_1336 ();
 sg13g2_decap_8 FILLER_56_1355 ();
 sg13g2_decap_8 FILLER_56_1362 ();
 sg13g2_fill_2 FILLER_56_1369 ();
 sg13g2_decap_4 FILLER_56_1397 ();
 sg13g2_fill_1 FILLER_56_1401 ();
 sg13g2_fill_2 FILLER_56_1443 ();
 sg13g2_decap_8 FILLER_56_1460 ();
 sg13g2_fill_2 FILLER_56_1480 ();
 sg13g2_fill_2 FILLER_56_1508 ();
 sg13g2_decap_8 FILLER_56_1515 ();
 sg13g2_decap_8 FILLER_56_1522 ();
 sg13g2_decap_8 FILLER_56_1529 ();
 sg13g2_decap_4 FILLER_56_1536 ();
 sg13g2_fill_1 FILLER_56_1540 ();
 sg13g2_fill_1 FILLER_56_1547 ();
 sg13g2_fill_1 FILLER_56_1561 ();
 sg13g2_fill_1 FILLER_56_1572 ();
 sg13g2_fill_2 FILLER_56_1590 ();
 sg13g2_fill_1 FILLER_56_1604 ();
 sg13g2_fill_1 FILLER_56_1610 ();
 sg13g2_decap_8 FILLER_56_1631 ();
 sg13g2_decap_4 FILLER_56_1638 ();
 sg13g2_fill_1 FILLER_56_1642 ();
 sg13g2_fill_2 FILLER_56_1655 ();
 sg13g2_fill_1 FILLER_56_1657 ();
 sg13g2_fill_1 FILLER_56_1683 ();
 sg13g2_fill_2 FILLER_56_1708 ();
 sg13g2_fill_2 FILLER_56_1715 ();
 sg13g2_fill_1 FILLER_56_1757 ();
 sg13g2_fill_1 FILLER_56_1792 ();
 sg13g2_decap_4 FILLER_56_1801 ();
 sg13g2_fill_2 FILLER_56_1810 ();
 sg13g2_fill_1 FILLER_56_1812 ();
 sg13g2_decap_8 FILLER_56_1821 ();
 sg13g2_decap_8 FILLER_56_1828 ();
 sg13g2_fill_2 FILLER_56_1835 ();
 sg13g2_fill_2 FILLER_56_1851 ();
 sg13g2_fill_1 FILLER_56_1857 ();
 sg13g2_decap_4 FILLER_56_1863 ();
 sg13g2_fill_2 FILLER_56_1867 ();
 sg13g2_decap_4 FILLER_56_1883 ();
 sg13g2_decap_4 FILLER_56_1901 ();
 sg13g2_decap_4 FILLER_56_1910 ();
 sg13g2_decap_8 FILLER_56_1919 ();
 sg13g2_decap_4 FILLER_56_1926 ();
 sg13g2_decap_4 FILLER_56_1935 ();
 sg13g2_fill_1 FILLER_56_1939 ();
 sg13g2_fill_1 FILLER_56_1950 ();
 sg13g2_fill_2 FILLER_56_1955 ();
 sg13g2_fill_1 FILLER_56_1966 ();
 sg13g2_fill_1 FILLER_56_1977 ();
 sg13g2_fill_1 FILLER_56_1984 ();
 sg13g2_fill_2 FILLER_56_2015 ();
 sg13g2_fill_1 FILLER_56_2017 ();
 sg13g2_fill_2 FILLER_56_2044 ();
 sg13g2_fill_1 FILLER_56_2046 ();
 sg13g2_decap_4 FILLER_56_2150 ();
 sg13g2_fill_1 FILLER_56_2154 ();
 sg13g2_fill_2 FILLER_56_2233 ();
 sg13g2_fill_1 FILLER_56_2278 ();
 sg13g2_fill_2 FILLER_56_2311 ();
 sg13g2_fill_2 FILLER_56_2326 ();
 sg13g2_fill_2 FILLER_56_2416 ();
 sg13g2_fill_1 FILLER_56_2434 ();
 sg13g2_fill_1 FILLER_56_2470 ();
 sg13g2_fill_2 FILLER_56_2594 ();
 sg13g2_fill_1 FILLER_56_2669 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_4 FILLER_57_34 ();
 sg13g2_fill_1 FILLER_57_38 ();
 sg13g2_fill_2 FILLER_57_120 ();
 sg13g2_decap_4 FILLER_57_152 ();
 sg13g2_decap_8 FILLER_57_166 ();
 sg13g2_fill_1 FILLER_57_173 ();
 sg13g2_decap_4 FILLER_57_210 ();
 sg13g2_fill_1 FILLER_57_214 ();
 sg13g2_fill_2 FILLER_57_223 ();
 sg13g2_fill_1 FILLER_57_225 ();
 sg13g2_fill_2 FILLER_57_230 ();
 sg13g2_fill_2 FILLER_57_260 ();
 sg13g2_fill_2 FILLER_57_271 ();
 sg13g2_fill_1 FILLER_57_277 ();
 sg13g2_fill_1 FILLER_57_291 ();
 sg13g2_decap_8 FILLER_57_323 ();
 sg13g2_decap_4 FILLER_57_330 ();
 sg13g2_fill_2 FILLER_57_360 ();
 sg13g2_fill_1 FILLER_57_362 ();
 sg13g2_fill_1 FILLER_57_405 ();
 sg13g2_fill_1 FILLER_57_412 ();
 sg13g2_fill_1 FILLER_57_432 ();
 sg13g2_fill_2 FILLER_57_492 ();
 sg13g2_fill_1 FILLER_57_494 ();
 sg13g2_fill_1 FILLER_57_514 ();
 sg13g2_decap_8 FILLER_57_545 ();
 sg13g2_fill_1 FILLER_57_552 ();
 sg13g2_fill_2 FILLER_57_564 ();
 sg13g2_fill_2 FILLER_57_571 ();
 sg13g2_fill_2 FILLER_57_600 ();
 sg13g2_fill_1 FILLER_57_628 ();
 sg13g2_fill_2 FILLER_57_640 ();
 sg13g2_fill_1 FILLER_57_646 ();
 sg13g2_fill_1 FILLER_57_651 ();
 sg13g2_fill_2 FILLER_57_662 ();
 sg13g2_fill_2 FILLER_57_669 ();
 sg13g2_fill_2 FILLER_57_697 ();
 sg13g2_fill_1 FILLER_57_703 ();
 sg13g2_fill_1 FILLER_57_717 ();
 sg13g2_fill_2 FILLER_57_753 ();
 sg13g2_fill_1 FILLER_57_788 ();
 sg13g2_decap_8 FILLER_57_855 ();
 sg13g2_decap_4 FILLER_57_862 ();
 sg13g2_fill_1 FILLER_57_866 ();
 sg13g2_decap_8 FILLER_57_875 ();
 sg13g2_decap_8 FILLER_57_882 ();
 sg13g2_decap_4 FILLER_57_889 ();
 sg13g2_fill_1 FILLER_57_893 ();
 sg13g2_decap_8 FILLER_57_908 ();
 sg13g2_fill_1 FILLER_57_915 ();
 sg13g2_decap_8 FILLER_57_920 ();
 sg13g2_fill_2 FILLER_57_927 ();
 sg13g2_decap_4 FILLER_57_933 ();
 sg13g2_fill_1 FILLER_57_975 ();
 sg13g2_fill_1 FILLER_57_986 ();
 sg13g2_fill_1 FILLER_57_1003 ();
 sg13g2_fill_1 FILLER_57_1010 ();
 sg13g2_fill_1 FILLER_57_1037 ();
 sg13g2_decap_4 FILLER_57_1054 ();
 sg13g2_fill_2 FILLER_57_1088 ();
 sg13g2_fill_1 FILLER_57_1090 ();
 sg13g2_fill_2 FILLER_57_1101 ();
 sg13g2_fill_1 FILLER_57_1103 ();
 sg13g2_fill_2 FILLER_57_1120 ();
 sg13g2_fill_1 FILLER_57_1122 ();
 sg13g2_decap_8 FILLER_57_1149 ();
 sg13g2_decap_8 FILLER_57_1166 ();
 sg13g2_decap_4 FILLER_57_1183 ();
 sg13g2_decap_8 FILLER_57_1213 ();
 sg13g2_fill_1 FILLER_57_1220 ();
 sg13g2_fill_2 FILLER_57_1248 ();
 sg13g2_decap_4 FILLER_57_1271 ();
 sg13g2_decap_8 FILLER_57_1293 ();
 sg13g2_decap_8 FILLER_57_1300 ();
 sg13g2_decap_8 FILLER_57_1307 ();
 sg13g2_fill_1 FILLER_57_1314 ();
 sg13g2_fill_2 FILLER_57_1319 ();
 sg13g2_fill_1 FILLER_57_1366 ();
 sg13g2_decap_8 FILLER_57_1372 ();
 sg13g2_fill_2 FILLER_57_1379 ();
 sg13g2_decap_8 FILLER_57_1391 ();
 sg13g2_decap_8 FILLER_57_1398 ();
 sg13g2_fill_1 FILLER_57_1405 ();
 sg13g2_fill_1 FILLER_57_1445 ();
 sg13g2_fill_2 FILLER_57_1470 ();
 sg13g2_fill_2 FILLER_57_1481 ();
 sg13g2_fill_2 FILLER_57_1487 ();
 sg13g2_fill_2 FILLER_57_1493 ();
 sg13g2_fill_1 FILLER_57_1495 ();
 sg13g2_decap_8 FILLER_57_1514 ();
 sg13g2_decap_8 FILLER_57_1521 ();
 sg13g2_fill_1 FILLER_57_1532 ();
 sg13g2_decap_4 FILLER_57_1537 ();
 sg13g2_fill_1 FILLER_57_1546 ();
 sg13g2_fill_1 FILLER_57_1559 ();
 sg13g2_fill_2 FILLER_57_1603 ();
 sg13g2_fill_1 FILLER_57_1605 ();
 sg13g2_decap_4 FILLER_57_1621 ();
 sg13g2_fill_2 FILLER_57_1638 ();
 sg13g2_decap_4 FILLER_57_1645 ();
 sg13g2_fill_1 FILLER_57_1649 ();
 sg13g2_decap_4 FILLER_57_1663 ();
 sg13g2_fill_2 FILLER_57_1703 ();
 sg13g2_fill_1 FILLER_57_1705 ();
 sg13g2_decap_4 FILLER_57_1746 ();
 sg13g2_fill_2 FILLER_57_1755 ();
 sg13g2_fill_2 FILLER_57_1775 ();
 sg13g2_fill_2 FILLER_57_1787 ();
 sg13g2_fill_1 FILLER_57_1789 ();
 sg13g2_decap_8 FILLER_57_1795 ();
 sg13g2_fill_1 FILLER_57_1802 ();
 sg13g2_fill_2 FILLER_57_1813 ();
 sg13g2_decap_8 FILLER_57_1820 ();
 sg13g2_decap_4 FILLER_57_1827 ();
 sg13g2_fill_2 FILLER_57_1835 ();
 sg13g2_fill_1 FILLER_57_1837 ();
 sg13g2_decap_4 FILLER_57_1842 ();
 sg13g2_fill_1 FILLER_57_1846 ();
 sg13g2_fill_2 FILLER_57_1851 ();
 sg13g2_decap_8 FILLER_57_1861 ();
 sg13g2_decap_4 FILLER_57_1868 ();
 sg13g2_fill_1 FILLER_57_1872 ();
 sg13g2_decap_8 FILLER_57_1878 ();
 sg13g2_decap_8 FILLER_57_1885 ();
 sg13g2_decap_8 FILLER_57_1892 ();
 sg13g2_decap_8 FILLER_57_1899 ();
 sg13g2_decap_8 FILLER_57_1917 ();
 sg13g2_decap_4 FILLER_57_1924 ();
 sg13g2_fill_1 FILLER_57_1939 ();
 sg13g2_fill_1 FILLER_57_1945 ();
 sg13g2_fill_2 FILLER_57_1966 ();
 sg13g2_fill_1 FILLER_57_1968 ();
 sg13g2_fill_1 FILLER_57_1978 ();
 sg13g2_fill_1 FILLER_57_1983 ();
 sg13g2_decap_4 FILLER_57_2059 ();
 sg13g2_fill_2 FILLER_57_2063 ();
 sg13g2_decap_4 FILLER_57_2068 ();
 sg13g2_fill_2 FILLER_57_2072 ();
 sg13g2_fill_2 FILLER_57_2078 ();
 sg13g2_fill_1 FILLER_57_2080 ();
 sg13g2_decap_8 FILLER_57_2091 ();
 sg13g2_decap_4 FILLER_57_2098 ();
 sg13g2_fill_1 FILLER_57_2102 ();
 sg13g2_fill_2 FILLER_57_2107 ();
 sg13g2_fill_1 FILLER_57_2133 ();
 sg13g2_decap_4 FILLER_57_2138 ();
 sg13g2_fill_2 FILLER_57_2152 ();
 sg13g2_decap_4 FILLER_57_2168 ();
 sg13g2_fill_2 FILLER_57_2172 ();
 sg13g2_fill_1 FILLER_57_2184 ();
 sg13g2_fill_1 FILLER_57_2195 ();
 sg13g2_fill_1 FILLER_57_2200 ();
 sg13g2_fill_1 FILLER_57_2205 ();
 sg13g2_fill_1 FILLER_57_2216 ();
 sg13g2_fill_2 FILLER_57_2269 ();
 sg13g2_decap_4 FILLER_57_2279 ();
 sg13g2_fill_2 FILLER_57_2283 ();
 sg13g2_fill_2 FILLER_57_2289 ();
 sg13g2_fill_1 FILLER_57_2301 ();
 sg13g2_fill_1 FILLER_57_2316 ();
 sg13g2_fill_2 FILLER_57_2365 ();
 sg13g2_fill_1 FILLER_57_2381 ();
 sg13g2_fill_2 FILLER_57_2408 ();
 sg13g2_fill_1 FILLER_57_2414 ();
 sg13g2_fill_2 FILLER_57_2445 ();
 sg13g2_fill_2 FILLER_57_2499 ();
 sg13g2_fill_2 FILLER_57_2552 ();
 sg13g2_fill_2 FILLER_57_2565 ();
 sg13g2_fill_1 FILLER_57_2599 ();
 sg13g2_fill_1 FILLER_57_2604 ();
 sg13g2_fill_2 FILLER_57_2668 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_4 FILLER_58_7 ();
 sg13g2_fill_2 FILLER_58_11 ();
 sg13g2_fill_1 FILLER_58_47 ();
 sg13g2_fill_2 FILLER_58_66 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_fill_1 FILLER_58_84 ();
 sg13g2_fill_1 FILLER_58_94 ();
 sg13g2_fill_1 FILLER_58_105 ();
 sg13g2_fill_1 FILLER_58_128 ();
 sg13g2_fill_1 FILLER_58_133 ();
 sg13g2_decap_4 FILLER_58_138 ();
 sg13g2_decap_4 FILLER_58_176 ();
 sg13g2_fill_2 FILLER_58_189 ();
 sg13g2_fill_1 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_209 ();
 sg13g2_decap_8 FILLER_58_216 ();
 sg13g2_decap_8 FILLER_58_223 ();
 sg13g2_decap_4 FILLER_58_230 ();
 sg13g2_fill_2 FILLER_58_234 ();
 sg13g2_decap_4 FILLER_58_239 ();
 sg13g2_fill_2 FILLER_58_302 ();
 sg13g2_fill_1 FILLER_58_304 ();
 sg13g2_fill_2 FILLER_58_309 ();
 sg13g2_fill_1 FILLER_58_319 ();
 sg13g2_fill_2 FILLER_58_325 ();
 sg13g2_fill_1 FILLER_58_327 ();
 sg13g2_fill_2 FILLER_58_338 ();
 sg13g2_fill_2 FILLER_58_344 ();
 sg13g2_fill_2 FILLER_58_377 ();
 sg13g2_fill_1 FILLER_58_398 ();
 sg13g2_fill_1 FILLER_58_433 ();
 sg13g2_fill_2 FILLER_58_440 ();
 sg13g2_fill_2 FILLER_58_445 ();
 sg13g2_fill_2 FILLER_58_453 ();
 sg13g2_fill_1 FILLER_58_455 ();
 sg13g2_fill_2 FILLER_58_464 ();
 sg13g2_fill_2 FILLER_58_471 ();
 sg13g2_fill_1 FILLER_58_503 ();
 sg13g2_fill_2 FILLER_58_524 ();
 sg13g2_fill_1 FILLER_58_536 ();
 sg13g2_fill_1 FILLER_58_580 ();
 sg13g2_fill_1 FILLER_58_622 ();
 sg13g2_fill_1 FILLER_58_669 ();
 sg13g2_fill_1 FILLER_58_674 ();
 sg13g2_decap_8 FILLER_58_699 ();
 sg13g2_decap_8 FILLER_58_706 ();
 sg13g2_fill_2 FILLER_58_713 ();
 sg13g2_fill_2 FILLER_58_793 ();
 sg13g2_fill_1 FILLER_58_824 ();
 sg13g2_fill_1 FILLER_58_830 ();
 sg13g2_fill_2 FILLER_58_836 ();
 sg13g2_fill_2 FILLER_58_864 ();
 sg13g2_fill_2 FILLER_58_870 ();
 sg13g2_fill_2 FILLER_58_882 ();
 sg13g2_fill_1 FILLER_58_884 ();
 sg13g2_fill_2 FILLER_58_916 ();
 sg13g2_fill_2 FILLER_58_951 ();
 sg13g2_fill_2 FILLER_58_958 ();
 sg13g2_fill_1 FILLER_58_960 ();
 sg13g2_decap_8 FILLER_58_1029 ();
 sg13g2_fill_1 FILLER_58_1036 ();
 sg13g2_fill_1 FILLER_58_1047 ();
 sg13g2_fill_2 FILLER_58_1090 ();
 sg13g2_fill_2 FILLER_58_1118 ();
 sg13g2_fill_1 FILLER_58_1120 ();
 sg13g2_fill_2 FILLER_58_1126 ();
 sg13g2_fill_1 FILLER_58_1128 ();
 sg13g2_fill_2 FILLER_58_1133 ();
 sg13g2_fill_2 FILLER_58_1161 ();
 sg13g2_fill_2 FILLER_58_1231 ();
 sg13g2_fill_1 FILLER_58_1233 ();
 sg13g2_decap_4 FILLER_58_1241 ();
 sg13g2_fill_1 FILLER_58_1245 ();
 sg13g2_decap_4 FILLER_58_1264 ();
 sg13g2_fill_2 FILLER_58_1268 ();
 sg13g2_fill_2 FILLER_58_1276 ();
 sg13g2_fill_1 FILLER_58_1283 ();
 sg13g2_decap_8 FILLER_58_1293 ();
 sg13g2_decap_8 FILLER_58_1300 ();
 sg13g2_decap_8 FILLER_58_1307 ();
 sg13g2_decap_8 FILLER_58_1352 ();
 sg13g2_fill_2 FILLER_58_1359 ();
 sg13g2_fill_1 FILLER_58_1361 ();
 sg13g2_fill_2 FILLER_58_1369 ();
 sg13g2_fill_1 FILLER_58_1376 ();
 sg13g2_fill_2 FILLER_58_1409 ();
 sg13g2_decap_4 FILLER_58_1415 ();
 sg13g2_fill_1 FILLER_58_1419 ();
 sg13g2_fill_1 FILLER_58_1428 ();
 sg13g2_fill_2 FILLER_58_1433 ();
 sg13g2_fill_1 FILLER_58_1435 ();
 sg13g2_decap_8 FILLER_58_1485 ();
 sg13g2_decap_8 FILLER_58_1492 ();
 sg13g2_decap_8 FILLER_58_1499 ();
 sg13g2_fill_2 FILLER_58_1506 ();
 sg13g2_fill_1 FILLER_58_1508 ();
 sg13g2_decap_8 FILLER_58_1519 ();
 sg13g2_fill_2 FILLER_58_1526 ();
 sg13g2_fill_1 FILLER_58_1528 ();
 sg13g2_fill_2 FILLER_58_1535 ();
 sg13g2_fill_1 FILLER_58_1547 ();
 sg13g2_fill_1 FILLER_58_1552 ();
 sg13g2_fill_2 FILLER_58_1569 ();
 sg13g2_fill_2 FILLER_58_1583 ();
 sg13g2_decap_8 FILLER_58_1589 ();
 sg13g2_fill_1 FILLER_58_1596 ();
 sg13g2_fill_1 FILLER_58_1602 ();
 sg13g2_decap_8 FILLER_58_1613 ();
 sg13g2_fill_2 FILLER_58_1624 ();
 sg13g2_decap_8 FILLER_58_1631 ();
 sg13g2_fill_1 FILLER_58_1638 ();
 sg13g2_decap_8 FILLER_58_1644 ();
 sg13g2_decap_4 FILLER_58_1651 ();
 sg13g2_fill_1 FILLER_58_1655 ();
 sg13g2_decap_4 FILLER_58_1669 ();
 sg13g2_decap_4 FILLER_58_1677 ();
 sg13g2_fill_2 FILLER_58_1681 ();
 sg13g2_fill_1 FILLER_58_1699 ();
 sg13g2_fill_2 FILLER_58_1726 ();
 sg13g2_fill_2 FILLER_58_1737 ();
 sg13g2_decap_8 FILLER_58_1755 ();
 sg13g2_fill_1 FILLER_58_1762 ();
 sg13g2_decap_8 FILLER_58_1785 ();
 sg13g2_decap_4 FILLER_58_1792 ();
 sg13g2_fill_1 FILLER_58_1796 ();
 sg13g2_decap_4 FILLER_58_1801 ();
 sg13g2_fill_1 FILLER_58_1805 ();
 sg13g2_decap_4 FILLER_58_1811 ();
 sg13g2_fill_1 FILLER_58_1815 ();
 sg13g2_fill_2 FILLER_58_1821 ();
 sg13g2_decap_8 FILLER_58_1827 ();
 sg13g2_fill_1 FILLER_58_1834 ();
 sg13g2_decap_4 FILLER_58_1839 ();
 sg13g2_fill_1 FILLER_58_1843 ();
 sg13g2_fill_1 FILLER_58_1853 ();
 sg13g2_decap_8 FILLER_58_1866 ();
 sg13g2_decap_8 FILLER_58_1873 ();
 sg13g2_decap_8 FILLER_58_1880 ();
 sg13g2_decap_8 FILLER_58_1887 ();
 sg13g2_decap_8 FILLER_58_1894 ();
 sg13g2_decap_8 FILLER_58_1905 ();
 sg13g2_fill_1 FILLER_58_1912 ();
 sg13g2_fill_1 FILLER_58_1939 ();
 sg13g2_fill_1 FILLER_58_1946 ();
 sg13g2_fill_1 FILLER_58_1951 ();
 sg13g2_fill_1 FILLER_58_1962 ();
 sg13g2_fill_1 FILLER_58_1970 ();
 sg13g2_fill_1 FILLER_58_1978 ();
 sg13g2_fill_1 FILLER_58_1984 ();
 sg13g2_fill_1 FILLER_58_1997 ();
 sg13g2_decap_4 FILLER_58_2003 ();
 sg13g2_fill_2 FILLER_58_2013 ();
 sg13g2_decap_8 FILLER_58_2032 ();
 sg13g2_fill_1 FILLER_58_2039 ();
 sg13g2_decap_8 FILLER_58_2044 ();
 sg13g2_decap_4 FILLER_58_2054 ();
 sg13g2_fill_2 FILLER_58_2058 ();
 sg13g2_fill_1 FILLER_58_2064 ();
 sg13g2_decap_8 FILLER_58_2069 ();
 sg13g2_decap_8 FILLER_58_2076 ();
 sg13g2_decap_8 FILLER_58_2114 ();
 sg13g2_decap_8 FILLER_58_2121 ();
 sg13g2_fill_2 FILLER_58_2128 ();
 sg13g2_decap_8 FILLER_58_2166 ();
 sg13g2_decap_8 FILLER_58_2173 ();
 sg13g2_decap_4 FILLER_58_2180 ();
 sg13g2_fill_1 FILLER_58_2184 ();
 sg13g2_decap_8 FILLER_58_2194 ();
 sg13g2_fill_2 FILLER_58_2201 ();
 sg13g2_fill_1 FILLER_58_2203 ();
 sg13g2_fill_2 FILLER_58_2243 ();
 sg13g2_fill_1 FILLER_58_2255 ();
 sg13g2_fill_1 FILLER_58_2260 ();
 sg13g2_decap_4 FILLER_58_2265 ();
 sg13g2_fill_1 FILLER_58_2269 ();
 sg13g2_fill_1 FILLER_58_2294 ();
 sg13g2_fill_2 FILLER_58_2344 ();
 sg13g2_fill_2 FILLER_58_2368 ();
 sg13g2_fill_1 FILLER_58_2404 ();
 sg13g2_fill_1 FILLER_58_2411 ();
 sg13g2_fill_1 FILLER_58_2438 ();
 sg13g2_fill_1 FILLER_58_2471 ();
 sg13g2_fill_1 FILLER_58_2490 ();
 sg13g2_fill_2 FILLER_58_2495 ();
 sg13g2_fill_2 FILLER_58_2526 ();
 sg13g2_fill_2 FILLER_58_2543 ();
 sg13g2_fill_2 FILLER_58_2555 ();
 sg13g2_fill_2 FILLER_58_2571 ();
 sg13g2_fill_2 FILLER_58_2642 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_4 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_11 ();
 sg13g2_fill_2 FILLER_59_26 ();
 sg13g2_fill_1 FILLER_59_28 ();
 sg13g2_fill_1 FILLER_59_44 ();
 sg13g2_decap_8 FILLER_59_76 ();
 sg13g2_decap_8 FILLER_59_83 ();
 sg13g2_decap_8 FILLER_59_90 ();
 sg13g2_decap_8 FILLER_59_97 ();
 sg13g2_decap_4 FILLER_59_104 ();
 sg13g2_decap_4 FILLER_59_112 ();
 sg13g2_fill_1 FILLER_59_116 ();
 sg13g2_decap_8 FILLER_59_125 ();
 sg13g2_decap_8 FILLER_59_132 ();
 sg13g2_decap_8 FILLER_59_139 ();
 sg13g2_decap_4 FILLER_59_146 ();
 sg13g2_fill_2 FILLER_59_150 ();
 sg13g2_decap_8 FILLER_59_162 ();
 sg13g2_decap_8 FILLER_59_169 ();
 sg13g2_decap_8 FILLER_59_176 ();
 sg13g2_decap_8 FILLER_59_183 ();
 sg13g2_fill_2 FILLER_59_194 ();
 sg13g2_fill_1 FILLER_59_209 ();
 sg13g2_decap_8 FILLER_59_219 ();
 sg13g2_fill_1 FILLER_59_226 ();
 sg13g2_decap_8 FILLER_59_329 ();
 sg13g2_fill_2 FILLER_59_336 ();
 sg13g2_fill_1 FILLER_59_338 ();
 sg13g2_fill_1 FILLER_59_348 ();
 sg13g2_fill_1 FILLER_59_359 ();
 sg13g2_fill_1 FILLER_59_365 ();
 sg13g2_fill_1 FILLER_59_392 ();
 sg13g2_fill_2 FILLER_59_401 ();
 sg13g2_fill_2 FILLER_59_418 ();
 sg13g2_fill_1 FILLER_59_473 ();
 sg13g2_fill_2 FILLER_59_483 ();
 sg13g2_decap_4 FILLER_59_514 ();
 sg13g2_decap_4 FILLER_59_525 ();
 sg13g2_fill_1 FILLER_59_529 ();
 sg13g2_decap_8 FILLER_59_533 ();
 sg13g2_decap_8 FILLER_59_540 ();
 sg13g2_fill_2 FILLER_59_547 ();
 sg13g2_decap_4 FILLER_59_554 ();
 sg13g2_fill_1 FILLER_59_558 ();
 sg13g2_fill_1 FILLER_59_639 ();
 sg13g2_decap_4 FILLER_59_654 ();
 sg13g2_fill_1 FILLER_59_658 ();
 sg13g2_fill_2 FILLER_59_663 ();
 sg13g2_decap_8 FILLER_59_670 ();
 sg13g2_decap_8 FILLER_59_677 ();
 sg13g2_fill_1 FILLER_59_684 ();
 sg13g2_fill_1 FILLER_59_697 ();
 sg13g2_decap_8 FILLER_59_703 ();
 sg13g2_fill_2 FILLER_59_715 ();
 sg13g2_fill_1 FILLER_59_721 ();
 sg13g2_fill_1 FILLER_59_761 ();
 sg13g2_fill_2 FILLER_59_780 ();
 sg13g2_fill_2 FILLER_59_808 ();
 sg13g2_fill_2 FILLER_59_825 ();
 sg13g2_fill_1 FILLER_59_851 ();
 sg13g2_decap_4 FILLER_59_857 ();
 sg13g2_fill_1 FILLER_59_909 ();
 sg13g2_fill_1 FILLER_59_914 ();
 sg13g2_fill_1 FILLER_59_941 ();
 sg13g2_fill_1 FILLER_59_948 ();
 sg13g2_decap_8 FILLER_59_965 ();
 sg13g2_fill_2 FILLER_59_976 ();
 sg13g2_decap_4 FILLER_59_1004 ();
 sg13g2_decap_8 FILLER_59_1012 ();
 sg13g2_fill_2 FILLER_59_1019 ();
 sg13g2_decap_8 FILLER_59_1057 ();
 sg13g2_decap_4 FILLER_59_1094 ();
 sg13g2_fill_1 FILLER_59_1098 ();
 sg13g2_fill_2 FILLER_59_1103 ();
 sg13g2_decap_8 FILLER_59_1118 ();
 sg13g2_fill_2 FILLER_59_1125 ();
 sg13g2_decap_8 FILLER_59_1224 ();
 sg13g2_fill_2 FILLER_59_1231 ();
 sg13g2_fill_1 FILLER_59_1233 ();
 sg13g2_fill_2 FILLER_59_1243 ();
 sg13g2_decap_8 FILLER_59_1249 ();
 sg13g2_decap_4 FILLER_59_1266 ();
 sg13g2_fill_2 FILLER_59_1270 ();
 sg13g2_fill_1 FILLER_59_1287 ();
 sg13g2_fill_2 FILLER_59_1311 ();
 sg13g2_fill_1 FILLER_59_1318 ();
 sg13g2_decap_8 FILLER_59_1361 ();
 sg13g2_fill_2 FILLER_59_1368 ();
 sg13g2_fill_1 FILLER_59_1370 ();
 sg13g2_decap_8 FILLER_59_1393 ();
 sg13g2_decap_8 FILLER_59_1400 ();
 sg13g2_decap_8 FILLER_59_1407 ();
 sg13g2_decap_8 FILLER_59_1414 ();
 sg13g2_fill_2 FILLER_59_1421 ();
 sg13g2_fill_1 FILLER_59_1423 ();
 sg13g2_decap_8 FILLER_59_1462 ();
 sg13g2_decap_8 FILLER_59_1469 ();
 sg13g2_decap_4 FILLER_59_1476 ();
 sg13g2_fill_1 FILLER_59_1480 ();
 sg13g2_decap_8 FILLER_59_1489 ();
 sg13g2_decap_8 FILLER_59_1496 ();
 sg13g2_fill_1 FILLER_59_1503 ();
 sg13g2_fill_2 FILLER_59_1507 ();
 sg13g2_fill_1 FILLER_59_1528 ();
 sg13g2_fill_1 FILLER_59_1545 ();
 sg13g2_fill_1 FILLER_59_1551 ();
 sg13g2_fill_1 FILLER_59_1581 ();
 sg13g2_decap_8 FILLER_59_1598 ();
 sg13g2_decap_8 FILLER_59_1605 ();
 sg13g2_decap_8 FILLER_59_1612 ();
 sg13g2_fill_2 FILLER_59_1627 ();
 sg13g2_fill_1 FILLER_59_1629 ();
 sg13g2_fill_1 FILLER_59_1638 ();
 sg13g2_fill_1 FILLER_59_1643 ();
 sg13g2_fill_1 FILLER_59_1649 ();
 sg13g2_decap_8 FILLER_59_1659 ();
 sg13g2_decap_8 FILLER_59_1666 ();
 sg13g2_decap_4 FILLER_59_1673 ();
 sg13g2_fill_2 FILLER_59_1677 ();
 sg13g2_fill_1 FILLER_59_1709 ();
 sg13g2_decap_4 FILLER_59_1719 ();
 sg13g2_decap_4 FILLER_59_1729 ();
 sg13g2_decap_4 FILLER_59_1736 ();
 sg13g2_fill_2 FILLER_59_1740 ();
 sg13g2_fill_1 FILLER_59_1747 ();
 sg13g2_decap_4 FILLER_59_1753 ();
 sg13g2_decap_8 FILLER_59_1761 ();
 sg13g2_decap_8 FILLER_59_1768 ();
 sg13g2_decap_8 FILLER_59_1775 ();
 sg13g2_decap_4 FILLER_59_1782 ();
 sg13g2_fill_1 FILLER_59_1786 ();
 sg13g2_fill_1 FILLER_59_1807 ();
 sg13g2_fill_2 FILLER_59_1875 ();
 sg13g2_fill_1 FILLER_59_1877 ();
 sg13g2_fill_2 FILLER_59_1892 ();
 sg13g2_fill_2 FILLER_59_1900 ();
 sg13g2_fill_1 FILLER_59_1902 ();
 sg13g2_fill_1 FILLER_59_1908 ();
 sg13g2_fill_2 FILLER_59_1915 ();
 sg13g2_fill_1 FILLER_59_1917 ();
 sg13g2_fill_1 FILLER_59_1932 ();
 sg13g2_fill_2 FILLER_59_1943 ();
 sg13g2_fill_2 FILLER_59_2019 ();
 sg13g2_fill_1 FILLER_59_2050 ();
 sg13g2_fill_1 FILLER_59_2054 ();
 sg13g2_fill_2 FILLER_59_2061 ();
 sg13g2_fill_1 FILLER_59_2063 ();
 sg13g2_decap_8 FILLER_59_2078 ();
 sg13g2_decap_4 FILLER_59_2085 ();
 sg13g2_fill_2 FILLER_59_2089 ();
 sg13g2_fill_2 FILLER_59_2095 ();
 sg13g2_fill_1 FILLER_59_2097 ();
 sg13g2_decap_8 FILLER_59_2121 ();
 sg13g2_fill_2 FILLER_59_2128 ();
 sg13g2_decap_8 FILLER_59_2134 ();
 sg13g2_fill_1 FILLER_59_2141 ();
 sg13g2_decap_4 FILLER_59_2152 ();
 sg13g2_fill_1 FILLER_59_2156 ();
 sg13g2_fill_2 FILLER_59_2167 ();
 sg13g2_fill_2 FILLER_59_2179 ();
 sg13g2_fill_1 FILLER_59_2181 ();
 sg13g2_fill_2 FILLER_59_2192 ();
 sg13g2_fill_1 FILLER_59_2194 ();
 sg13g2_fill_2 FILLER_59_2216 ();
 sg13g2_fill_2 FILLER_59_2244 ();
 sg13g2_fill_2 FILLER_59_2299 ();
 sg13g2_fill_2 FILLER_59_2306 ();
 sg13g2_fill_1 FILLER_59_2324 ();
 sg13g2_fill_2 FILLER_59_2352 ();
 sg13g2_fill_1 FILLER_59_2359 ();
 sg13g2_fill_2 FILLER_59_2395 ();
 sg13g2_fill_1 FILLER_59_2403 ();
 sg13g2_fill_1 FILLER_59_2409 ();
 sg13g2_fill_2 FILLER_59_2417 ();
 sg13g2_fill_2 FILLER_59_2427 ();
 sg13g2_fill_1 FILLER_59_2429 ();
 sg13g2_fill_2 FILLER_59_2436 ();
 sg13g2_fill_1 FILLER_59_2438 ();
 sg13g2_fill_1 FILLER_59_2443 ();
 sg13g2_decap_4 FILLER_59_2448 ();
 sg13g2_fill_2 FILLER_59_2452 ();
 sg13g2_fill_1 FILLER_59_2458 ();
 sg13g2_fill_1 FILLER_59_2471 ();
 sg13g2_fill_1 FILLER_59_2501 ();
 sg13g2_fill_2 FILLER_59_2554 ();
 sg13g2_fill_1 FILLER_59_2585 ();
 sg13g2_fill_2 FILLER_59_2628 ();
 sg13g2_fill_1 FILLER_59_2640 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_34 ();
 sg13g2_fill_1 FILLER_60_41 ();
 sg13g2_fill_1 FILLER_60_46 ();
 sg13g2_fill_2 FILLER_60_83 ();
 sg13g2_decap_8 FILLER_60_95 ();
 sg13g2_decap_4 FILLER_60_102 ();
 sg13g2_fill_1 FILLER_60_106 ();
 sg13g2_fill_1 FILLER_60_126 ();
 sg13g2_fill_2 FILLER_60_157 ();
 sg13g2_fill_2 FILLER_60_204 ();
 sg13g2_fill_2 FILLER_60_232 ();
 sg13g2_fill_1 FILLER_60_234 ();
 sg13g2_fill_2 FILLER_60_239 ();
 sg13g2_fill_1 FILLER_60_241 ();
 sg13g2_fill_2 FILLER_60_246 ();
 sg13g2_fill_2 FILLER_60_279 ();
 sg13g2_fill_1 FILLER_60_281 ();
 sg13g2_fill_2 FILLER_60_286 ();
 sg13g2_fill_2 FILLER_60_293 ();
 sg13g2_fill_1 FILLER_60_295 ();
 sg13g2_decap_8 FILLER_60_331 ();
 sg13g2_decap_8 FILLER_60_338 ();
 sg13g2_fill_2 FILLER_60_345 ();
 sg13g2_fill_1 FILLER_60_347 ();
 sg13g2_fill_1 FILLER_60_358 ();
 sg13g2_fill_1 FILLER_60_364 ();
 sg13g2_fill_2 FILLER_60_431 ();
 sg13g2_fill_1 FILLER_60_468 ();
 sg13g2_fill_2 FILLER_60_493 ();
 sg13g2_fill_1 FILLER_60_495 ();
 sg13g2_decap_8 FILLER_60_500 ();
 sg13g2_decap_4 FILLER_60_507 ();
 sg13g2_fill_2 FILLER_60_524 ();
 sg13g2_fill_1 FILLER_60_526 ();
 sg13g2_fill_2 FILLER_60_535 ();
 sg13g2_fill_2 FILLER_60_542 ();
 sg13g2_fill_2 FILLER_60_549 ();
 sg13g2_decap_4 FILLER_60_635 ();
 sg13g2_fill_2 FILLER_60_639 ();
 sg13g2_decap_4 FILLER_60_653 ();
 sg13g2_fill_2 FILLER_60_657 ();
 sg13g2_decap_8 FILLER_60_663 ();
 sg13g2_decap_8 FILLER_60_670 ();
 sg13g2_fill_2 FILLER_60_677 ();
 sg13g2_fill_1 FILLER_60_679 ();
 sg13g2_decap_8 FILLER_60_692 ();
 sg13g2_fill_1 FILLER_60_704 ();
 sg13g2_fill_1 FILLER_60_709 ();
 sg13g2_fill_1 FILLER_60_755 ();
 sg13g2_fill_2 FILLER_60_782 ();
 sg13g2_fill_2 FILLER_60_821 ();
 sg13g2_fill_2 FILLER_60_829 ();
 sg13g2_fill_1 FILLER_60_839 ();
 sg13g2_decap_4 FILLER_60_856 ();
 sg13g2_fill_2 FILLER_60_860 ();
 sg13g2_fill_1 FILLER_60_906 ();
 sg13g2_fill_2 FILLER_60_939 ();
 sg13g2_fill_1 FILLER_60_941 ();
 sg13g2_decap_4 FILLER_60_968 ();
 sg13g2_fill_1 FILLER_60_972 ();
 sg13g2_decap_4 FILLER_60_983 ();
 sg13g2_fill_1 FILLER_60_987 ();
 sg13g2_fill_2 FILLER_60_1007 ();
 sg13g2_decap_8 FILLER_60_1049 ();
 sg13g2_fill_2 FILLER_60_1056 ();
 sg13g2_fill_1 FILLER_60_1058 ();
 sg13g2_decap_4 FILLER_60_1069 ();
 sg13g2_decap_8 FILLER_60_1077 ();
 sg13g2_decap_8 FILLER_60_1084 ();
 sg13g2_decap_8 FILLER_60_1091 ();
 sg13g2_decap_4 FILLER_60_1098 ();
 sg13g2_fill_1 FILLER_60_1102 ();
 sg13g2_decap_4 FILLER_60_1129 ();
 sg13g2_fill_2 FILLER_60_1133 ();
 sg13g2_decap_4 FILLER_60_1139 ();
 sg13g2_decap_8 FILLER_60_1147 ();
 sg13g2_fill_2 FILLER_60_1154 ();
 sg13g2_fill_1 FILLER_60_1156 ();
 sg13g2_fill_1 FILLER_60_1167 ();
 sg13g2_fill_1 FILLER_60_1172 ();
 sg13g2_fill_1 FILLER_60_1183 ();
 sg13g2_fill_2 FILLER_60_1262 ();
 sg13g2_fill_1 FILLER_60_1264 ();
 sg13g2_fill_1 FILLER_60_1270 ();
 sg13g2_fill_2 FILLER_60_1276 ();
 sg13g2_fill_1 FILLER_60_1283 ();
 sg13g2_fill_2 FILLER_60_1292 ();
 sg13g2_decap_8 FILLER_60_1311 ();
 sg13g2_fill_1 FILLER_60_1318 ();
 sg13g2_fill_2 FILLER_60_1344 ();
 sg13g2_fill_1 FILLER_60_1361 ();
 sg13g2_decap_8 FILLER_60_1369 ();
 sg13g2_decap_4 FILLER_60_1376 ();
 sg13g2_fill_2 FILLER_60_1389 ();
 sg13g2_fill_1 FILLER_60_1391 ();
 sg13g2_fill_1 FILLER_60_1400 ();
 sg13g2_fill_2 FILLER_60_1417 ();
 sg13g2_fill_1 FILLER_60_1424 ();
 sg13g2_fill_1 FILLER_60_1446 ();
 sg13g2_decap_4 FILLER_60_1463 ();
 sg13g2_fill_2 FILLER_60_1467 ();
 sg13g2_decap_4 FILLER_60_1473 ();
 sg13g2_decap_8 FILLER_60_1481 ();
 sg13g2_decap_8 FILLER_60_1488 ();
 sg13g2_decap_4 FILLER_60_1495 ();
 sg13g2_fill_1 FILLER_60_1576 ();
 sg13g2_decap_8 FILLER_60_1582 ();
 sg13g2_decap_8 FILLER_60_1589 ();
 sg13g2_decap_8 FILLER_60_1596 ();
 sg13g2_decap_8 FILLER_60_1608 ();
 sg13g2_decap_8 FILLER_60_1615 ();
 sg13g2_fill_2 FILLER_60_1630 ();
 sg13g2_fill_1 FILLER_60_1632 ();
 sg13g2_fill_1 FILLER_60_1638 ();
 sg13g2_fill_1 FILLER_60_1659 ();
 sg13g2_decap_8 FILLER_60_1664 ();
 sg13g2_decap_8 FILLER_60_1671 ();
 sg13g2_decap_8 FILLER_60_1678 ();
 sg13g2_decap_8 FILLER_60_1685 ();
 sg13g2_fill_1 FILLER_60_1692 ();
 sg13g2_decap_8 FILLER_60_1701 ();
 sg13g2_fill_1 FILLER_60_1708 ();
 sg13g2_fill_2 FILLER_60_1720 ();
 sg13g2_fill_1 FILLER_60_1722 ();
 sg13g2_fill_1 FILLER_60_1729 ();
 sg13g2_decap_8 FILLER_60_1775 ();
 sg13g2_decap_4 FILLER_60_1782 ();
 sg13g2_fill_2 FILLER_60_1786 ();
 sg13g2_decap_4 FILLER_60_1801 ();
 sg13g2_decap_4 FILLER_60_1834 ();
 sg13g2_fill_1 FILLER_60_1848 ();
 sg13g2_decap_4 FILLER_60_1861 ();
 sg13g2_fill_2 FILLER_60_1870 ();
 sg13g2_fill_1 FILLER_60_1872 ();
 sg13g2_fill_2 FILLER_60_1877 ();
 sg13g2_fill_1 FILLER_60_1879 ();
 sg13g2_fill_1 FILLER_60_1895 ();
 sg13g2_decap_8 FILLER_60_1906 ();
 sg13g2_fill_2 FILLER_60_1913 ();
 sg13g2_fill_2 FILLER_60_1928 ();
 sg13g2_fill_1 FILLER_60_1957 ();
 sg13g2_fill_2 FILLER_60_1995 ();
 sg13g2_fill_2 FILLER_60_2012 ();
 sg13g2_fill_1 FILLER_60_2014 ();
 sg13g2_fill_2 FILLER_60_2020 ();
 sg13g2_fill_1 FILLER_60_2022 ();
 sg13g2_fill_1 FILLER_60_2050 ();
 sg13g2_fill_1 FILLER_60_2068 ();
 sg13g2_fill_1 FILLER_60_2095 ();
 sg13g2_decap_4 FILLER_60_2122 ();
 sg13g2_fill_1 FILLER_60_2126 ();
 sg13g2_fill_2 FILLER_60_2174 ();
 sg13g2_decap_8 FILLER_60_2242 ();
 sg13g2_decap_4 FILLER_60_2249 ();
 sg13g2_fill_2 FILLER_60_2279 ();
 sg13g2_fill_1 FILLER_60_2286 ();
 sg13g2_fill_1 FILLER_60_2299 ();
 sg13g2_fill_2 FILLER_60_2310 ();
 sg13g2_fill_2 FILLER_60_2323 ();
 sg13g2_fill_1 FILLER_60_2351 ();
 sg13g2_fill_1 FILLER_60_2361 ();
 sg13g2_fill_1 FILLER_60_2376 ();
 sg13g2_fill_1 FILLER_60_2407 ();
 sg13g2_fill_2 FILLER_60_2413 ();
 sg13g2_decap_4 FILLER_60_2420 ();
 sg13g2_fill_1 FILLER_60_2424 ();
 sg13g2_decap_4 FILLER_60_2433 ();
 sg13g2_fill_1 FILLER_60_2437 ();
 sg13g2_fill_1 FILLER_60_2450 ();
 sg13g2_fill_1 FILLER_60_2471 ();
 sg13g2_fill_1 FILLER_60_2477 ();
 sg13g2_fill_1 FILLER_60_2504 ();
 sg13g2_fill_1 FILLER_60_2514 ();
 sg13g2_fill_2 FILLER_60_2524 ();
 sg13g2_fill_2 FILLER_60_2538 ();
 sg13g2_fill_1 FILLER_60_2584 ();
 sg13g2_fill_2 FILLER_60_2607 ();
 sg13g2_fill_1 FILLER_60_2615 ();
 sg13g2_fill_1 FILLER_60_2626 ();
 sg13g2_fill_1 FILLER_60_2631 ();
 sg13g2_fill_1 FILLER_60_2658 ();
 sg13g2_fill_1 FILLER_60_2669 ();
 sg13g2_decap_4 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_fill_2 FILLER_61_56 ();
 sg13g2_fill_1 FILLER_61_58 ();
 sg13g2_fill_2 FILLER_61_67 ();
 sg13g2_fill_1 FILLER_61_69 ();
 sg13g2_fill_1 FILLER_61_74 ();
 sg13g2_fill_1 FILLER_61_80 ();
 sg13g2_fill_1 FILLER_61_91 ();
 sg13g2_fill_1 FILLER_61_97 ();
 sg13g2_fill_1 FILLER_61_163 ();
 sg13g2_fill_1 FILLER_61_218 ();
 sg13g2_fill_2 FILLER_61_253 ();
 sg13g2_fill_1 FILLER_61_255 ();
 sg13g2_fill_2 FILLER_61_261 ();
 sg13g2_decap_4 FILLER_61_276 ();
 sg13g2_fill_1 FILLER_61_289 ();
 sg13g2_fill_2 FILLER_61_294 ();
 sg13g2_fill_1 FILLER_61_296 ();
 sg13g2_fill_2 FILLER_61_311 ();
 sg13g2_fill_1 FILLER_61_313 ();
 sg13g2_decap_8 FILLER_61_318 ();
 sg13g2_fill_1 FILLER_61_325 ();
 sg13g2_decap_8 FILLER_61_336 ();
 sg13g2_decap_8 FILLER_61_343 ();
 sg13g2_decap_4 FILLER_61_350 ();
 sg13g2_fill_1 FILLER_61_354 ();
 sg13g2_fill_2 FILLER_61_360 ();
 sg13g2_fill_1 FILLER_61_375 ();
 sg13g2_fill_1 FILLER_61_417 ();
 sg13g2_fill_1 FILLER_61_434 ();
 sg13g2_fill_1 FILLER_61_444 ();
 sg13g2_fill_2 FILLER_61_450 ();
 sg13g2_fill_1 FILLER_61_469 ();
 sg13g2_fill_2 FILLER_61_477 ();
 sg13g2_fill_1 FILLER_61_494 ();
 sg13g2_decap_8 FILLER_61_499 ();
 sg13g2_decap_4 FILLER_61_510 ();
 sg13g2_fill_1 FILLER_61_514 ();
 sg13g2_decap_4 FILLER_61_524 ();
 sg13g2_fill_2 FILLER_61_528 ();
 sg13g2_fill_2 FILLER_61_559 ();
 sg13g2_fill_2 FILLER_61_657 ();
 sg13g2_fill_2 FILLER_61_690 ();
 sg13g2_fill_1 FILLER_61_696 ();
 sg13g2_fill_1 FILLER_61_728 ();
 sg13g2_fill_2 FILLER_61_734 ();
 sg13g2_fill_2 FILLER_61_750 ();
 sg13g2_fill_2 FILLER_61_770 ();
 sg13g2_fill_2 FILLER_61_792 ();
 sg13g2_fill_2 FILLER_61_802 ();
 sg13g2_fill_1 FILLER_61_813 ();
 sg13g2_decap_8 FILLER_61_847 ();
 sg13g2_decap_8 FILLER_61_854 ();
 sg13g2_decap_8 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_61_868 ();
 sg13g2_fill_2 FILLER_61_875 ();
 sg13g2_fill_1 FILLER_61_885 ();
 sg13g2_decap_8 FILLER_61_894 ();
 sg13g2_decap_8 FILLER_61_901 ();
 sg13g2_fill_1 FILLER_61_937 ();
 sg13g2_fill_1 FILLER_61_942 ();
 sg13g2_fill_1 FILLER_61_953 ();
 sg13g2_fill_1 FILLER_61_980 ();
 sg13g2_fill_1 FILLER_61_1011 ();
 sg13g2_fill_2 FILLER_61_1022 ();
 sg13g2_decap_8 FILLER_61_1118 ();
 sg13g2_decap_8 FILLER_61_1125 ();
 sg13g2_fill_2 FILLER_61_1132 ();
 sg13g2_fill_2 FILLER_61_1183 ();
 sg13g2_fill_2 FILLER_61_1199 ();
 sg13g2_fill_1 FILLER_61_1201 ();
 sg13g2_fill_2 FILLER_61_1244 ();
 sg13g2_fill_2 FILLER_61_1259 ();
 sg13g2_fill_2 FILLER_61_1268 ();
 sg13g2_fill_1 FILLER_61_1270 ();
 sg13g2_fill_1 FILLER_61_1297 ();
 sg13g2_decap_8 FILLER_61_1303 ();
 sg13g2_fill_1 FILLER_61_1310 ();
 sg13g2_decap_8 FILLER_61_1319 ();
 sg13g2_fill_2 FILLER_61_1326 ();
 sg13g2_fill_1 FILLER_61_1328 ();
 sg13g2_decap_8 FILLER_61_1351 ();
 sg13g2_decap_4 FILLER_61_1358 ();
 sg13g2_fill_1 FILLER_61_1362 ();
 sg13g2_fill_2 FILLER_61_1387 ();
 sg13g2_fill_1 FILLER_61_1409 ();
 sg13g2_fill_1 FILLER_61_1418 ();
 sg13g2_fill_2 FILLER_61_1435 ();
 sg13g2_fill_1 FILLER_61_1437 ();
 sg13g2_decap_4 FILLER_61_1459 ();
 sg13g2_fill_2 FILLER_61_1463 ();
 sg13g2_decap_4 FILLER_61_1496 ();
 sg13g2_fill_1 FILLER_61_1500 ();
 sg13g2_fill_2 FILLER_61_1536 ();
 sg13g2_fill_1 FILLER_61_1578 ();
 sg13g2_decap_8 FILLER_61_1602 ();
 sg13g2_decap_8 FILLER_61_1609 ();
 sg13g2_fill_2 FILLER_61_1625 ();
 sg13g2_fill_1 FILLER_61_1636 ();
 sg13g2_fill_1 FILLER_61_1646 ();
 sg13g2_decap_8 FILLER_61_1661 ();
 sg13g2_decap_8 FILLER_61_1668 ();
 sg13g2_decap_8 FILLER_61_1675 ();
 sg13g2_decap_8 FILLER_61_1682 ();
 sg13g2_fill_2 FILLER_61_1689 ();
 sg13g2_fill_1 FILLER_61_1691 ();
 sg13g2_fill_1 FILLER_61_1701 ();
 sg13g2_fill_1 FILLER_61_1706 ();
 sg13g2_fill_1 FILLER_61_1727 ();
 sg13g2_fill_1 FILLER_61_1735 ();
 sg13g2_fill_1 FILLER_61_1748 ();
 sg13g2_fill_2 FILLER_61_1762 ();
 sg13g2_decap_8 FILLER_61_1769 ();
 sg13g2_decap_8 FILLER_61_1776 ();
 sg13g2_decap_4 FILLER_61_1783 ();
 sg13g2_fill_1 FILLER_61_1787 ();
 sg13g2_decap_8 FILLER_61_1793 ();
 sg13g2_fill_2 FILLER_61_1800 ();
 sg13g2_fill_1 FILLER_61_1802 ();
 sg13g2_decap_4 FILLER_61_1841 ();
 sg13g2_fill_2 FILLER_61_1845 ();
 sg13g2_fill_2 FILLER_61_1852 ();
 sg13g2_fill_2 FILLER_61_1867 ();
 sg13g2_fill_1 FILLER_61_1869 ();
 sg13g2_fill_2 FILLER_61_1874 ();
 sg13g2_fill_1 FILLER_61_1876 ();
 sg13g2_fill_2 FILLER_61_1889 ();
 sg13g2_fill_1 FILLER_61_1891 ();
 sg13g2_fill_1 FILLER_61_1905 ();
 sg13g2_decap_4 FILLER_61_1911 ();
 sg13g2_fill_2 FILLER_61_1915 ();
 sg13g2_decap_4 FILLER_61_1922 ();
 sg13g2_fill_1 FILLER_61_1926 ();
 sg13g2_fill_1 FILLER_61_2000 ();
 sg13g2_decap_8 FILLER_61_2025 ();
 sg13g2_fill_2 FILLER_61_2032 ();
 sg13g2_fill_1 FILLER_61_2056 ();
 sg13g2_fill_2 FILLER_61_2083 ();
 sg13g2_fill_2 FILLER_61_2095 ();
 sg13g2_fill_1 FILLER_61_2097 ();
 sg13g2_decap_8 FILLER_61_2106 ();
 sg13g2_decap_4 FILLER_61_2113 ();
 sg13g2_fill_2 FILLER_61_2157 ();
 sg13g2_fill_2 FILLER_61_2185 ();
 sg13g2_fill_2 FILLER_61_2226 ();
 sg13g2_decap_8 FILLER_61_2232 ();
 sg13g2_decap_8 FILLER_61_2239 ();
 sg13g2_fill_1 FILLER_61_2246 ();
 sg13g2_fill_2 FILLER_61_2283 ();
 sg13g2_fill_1 FILLER_61_2322 ();
 sg13g2_fill_1 FILLER_61_2328 ();
 sg13g2_fill_2 FILLER_61_2389 ();
 sg13g2_fill_2 FILLER_61_2408 ();
 sg13g2_decap_4 FILLER_61_2420 ();
 sg13g2_fill_2 FILLER_61_2424 ();
 sg13g2_fill_2 FILLER_61_2431 ();
 sg13g2_fill_1 FILLER_61_2433 ();
 sg13g2_fill_1 FILLER_61_2438 ();
 sg13g2_fill_2 FILLER_61_2443 ();
 sg13g2_decap_4 FILLER_61_2451 ();
 sg13g2_fill_1 FILLER_61_2455 ();
 sg13g2_fill_2 FILLER_61_2520 ();
 sg13g2_fill_2 FILLER_61_2609 ();
 sg13g2_fill_1 FILLER_61_2647 ();
 sg13g2_decap_4 FILLER_61_2655 ();
 sg13g2_fill_1 FILLER_61_2665 ();
 sg13g2_fill_1 FILLER_61_2669 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_7 ();
 sg13g2_fill_1 FILLER_62_9 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_4 FILLER_62_31 ();
 sg13g2_fill_2 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_41 ();
 sg13g2_decap_8 FILLER_62_48 ();
 sg13g2_decap_4 FILLER_62_55 ();
 sg13g2_fill_1 FILLER_62_59 ();
 sg13g2_fill_2 FILLER_62_90 ();
 sg13g2_fill_1 FILLER_62_92 ();
 sg13g2_fill_2 FILLER_62_124 ();
 sg13g2_fill_1 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_163 ();
 sg13g2_fill_2 FILLER_62_185 ();
 sg13g2_fill_2 FILLER_62_259 ();
 sg13g2_decap_4 FILLER_62_273 ();
 sg13g2_fill_1 FILLER_62_277 ();
 sg13g2_fill_2 FILLER_62_287 ();
 sg13g2_decap_8 FILLER_62_294 ();
 sg13g2_fill_1 FILLER_62_301 ();
 sg13g2_decap_8 FILLER_62_310 ();
 sg13g2_decap_8 FILLER_62_320 ();
 sg13g2_decap_4 FILLER_62_327 ();
 sg13g2_fill_1 FILLER_62_331 ();
 sg13g2_fill_1 FILLER_62_372 ();
 sg13g2_fill_2 FILLER_62_378 ();
 sg13g2_fill_1 FILLER_62_475 ();
 sg13g2_fill_1 FILLER_62_494 ();
 sg13g2_fill_2 FILLER_62_499 ();
 sg13g2_fill_1 FILLER_62_505 ();
 sg13g2_fill_2 FILLER_62_511 ();
 sg13g2_fill_2 FILLER_62_523 ();
 sg13g2_fill_2 FILLER_62_529 ();
 sg13g2_fill_1 FILLER_62_531 ();
 sg13g2_fill_2 FILLER_62_571 ();
 sg13g2_fill_1 FILLER_62_573 ();
 sg13g2_fill_1 FILLER_62_585 ();
 sg13g2_fill_2 FILLER_62_591 ();
 sg13g2_fill_2 FILLER_62_597 ();
 sg13g2_decap_4 FILLER_62_618 ();
 sg13g2_fill_1 FILLER_62_622 ();
 sg13g2_fill_1 FILLER_62_628 ();
 sg13g2_fill_1 FILLER_62_633 ();
 sg13g2_fill_1 FILLER_62_666 ();
 sg13g2_fill_1 FILLER_62_677 ();
 sg13g2_decap_8 FILLER_62_682 ();
 sg13g2_decap_8 FILLER_62_689 ();
 sg13g2_decap_4 FILLER_62_696 ();
 sg13g2_fill_1 FILLER_62_726 ();
 sg13g2_fill_1 FILLER_62_812 ();
 sg13g2_fill_1 FILLER_62_854 ();
 sg13g2_fill_2 FILLER_62_881 ();
 sg13g2_decap_8 FILLER_62_893 ();
 sg13g2_fill_1 FILLER_62_904 ();
 sg13g2_fill_2 FILLER_62_931 ();
 sg13g2_fill_1 FILLER_62_933 ();
 sg13g2_fill_2 FILLER_62_968 ();
 sg13g2_fill_2 FILLER_62_977 ();
 sg13g2_fill_1 FILLER_62_979 ();
 sg13g2_fill_2 FILLER_62_1016 ();
 sg13g2_fill_2 FILLER_62_1022 ();
 sg13g2_fill_1 FILLER_62_1024 ();
 sg13g2_fill_2 FILLER_62_1035 ();
 sg13g2_fill_1 FILLER_62_1037 ();
 sg13g2_fill_2 FILLER_62_1044 ();
 sg13g2_fill_2 FILLER_62_1072 ();
 sg13g2_fill_1 FILLER_62_1074 ();
 sg13g2_decap_4 FILLER_62_1079 ();
 sg13g2_fill_1 FILLER_62_1083 ();
 sg13g2_fill_1 FILLER_62_1104 ();
 sg13g2_decap_4 FILLER_62_1113 ();
 sg13g2_decap_4 FILLER_62_1148 ();
 sg13g2_fill_2 FILLER_62_1152 ();
 sg13g2_fill_2 FILLER_62_1158 ();
 sg13g2_fill_2 FILLER_62_1186 ();
 sg13g2_fill_1 FILLER_62_1188 ();
 sg13g2_fill_1 FILLER_62_1267 ();
 sg13g2_fill_2 FILLER_62_1278 ();
 sg13g2_fill_1 FILLER_62_1285 ();
 sg13g2_fill_1 FILLER_62_1293 ();
 sg13g2_fill_2 FILLER_62_1304 ();
 sg13g2_fill_1 FILLER_62_1306 ();
 sg13g2_decap_4 FILLER_62_1316 ();
 sg13g2_fill_2 FILLER_62_1327 ();
 sg13g2_fill_1 FILLER_62_1329 ();
 sg13g2_decap_4 FILLER_62_1349 ();
 sg13g2_decap_4 FILLER_62_1358 ();
 sg13g2_fill_1 FILLER_62_1362 ();
 sg13g2_fill_1 FILLER_62_1370 ();
 sg13g2_fill_2 FILLER_62_1387 ();
 sg13g2_fill_2 FILLER_62_1394 ();
 sg13g2_decap_4 FILLER_62_1411 ();
 sg13g2_fill_1 FILLER_62_1415 ();
 sg13g2_fill_2 FILLER_62_1439 ();
 sg13g2_fill_2 FILLER_62_1457 ();
 sg13g2_fill_1 FILLER_62_1459 ();
 sg13g2_fill_2 FILLER_62_1491 ();
 sg13g2_decap_8 FILLER_62_1503 ();
 sg13g2_decap_4 FILLER_62_1510 ();
 sg13g2_fill_1 FILLER_62_1514 ();
 sg13g2_fill_1 FILLER_62_1534 ();
 sg13g2_fill_2 FILLER_62_1613 ();
 sg13g2_decap_4 FILLER_62_1645 ();
 sg13g2_fill_1 FILLER_62_1649 ();
 sg13g2_fill_2 FILLER_62_1673 ();
 sg13g2_decap_8 FILLER_62_1679 ();
 sg13g2_fill_1 FILLER_62_1686 ();
 sg13g2_fill_2 FILLER_62_1695 ();
 sg13g2_fill_1 FILLER_62_1697 ();
 sg13g2_fill_2 FILLER_62_1702 ();
 sg13g2_fill_1 FILLER_62_1717 ();
 sg13g2_fill_1 FILLER_62_1722 ();
 sg13g2_fill_1 FILLER_62_1729 ();
 sg13g2_fill_1 FILLER_62_1739 ();
 sg13g2_fill_2 FILLER_62_1748 ();
 sg13g2_fill_1 FILLER_62_1750 ();
 sg13g2_fill_1 FILLER_62_1760 ();
 sg13g2_fill_2 FILLER_62_1764 ();
 sg13g2_decap_8 FILLER_62_1797 ();
 sg13g2_decap_8 FILLER_62_1804 ();
 sg13g2_decap_4 FILLER_62_1811 ();
 sg13g2_fill_1 FILLER_62_1815 ();
 sg13g2_decap_4 FILLER_62_1830 ();
 sg13g2_fill_1 FILLER_62_1834 ();
 sg13g2_fill_1 FILLER_62_1845 ();
 sg13g2_fill_1 FILLER_62_1870 ();
 sg13g2_fill_2 FILLER_62_1875 ();
 sg13g2_fill_2 FILLER_62_1885 ();
 sg13g2_decap_8 FILLER_62_1902 ();
 sg13g2_decap_8 FILLER_62_1909 ();
 sg13g2_decap_8 FILLER_62_1916 ();
 sg13g2_fill_1 FILLER_62_1936 ();
 sg13g2_fill_1 FILLER_62_1981 ();
 sg13g2_decap_8 FILLER_62_2022 ();
 sg13g2_fill_2 FILLER_62_2038 ();
 sg13g2_fill_2 FILLER_62_2108 ();
 sg13g2_fill_1 FILLER_62_2110 ();
 sg13g2_fill_2 FILLER_62_2121 ();
 sg13g2_fill_2 FILLER_62_2127 ();
 sg13g2_fill_2 FILLER_62_2159 ();
 sg13g2_fill_2 FILLER_62_2166 ();
 sg13g2_fill_1 FILLER_62_2168 ();
 sg13g2_decap_4 FILLER_62_2234 ();
 sg13g2_fill_1 FILLER_62_2238 ();
 sg13g2_decap_8 FILLER_62_2243 ();
 sg13g2_decap_4 FILLER_62_2250 ();
 sg13g2_fill_1 FILLER_62_2262 ();
 sg13g2_fill_2 FILLER_62_2277 ();
 sg13g2_fill_1 FILLER_62_2299 ();
 sg13g2_fill_1 FILLER_62_2312 ();
 sg13g2_fill_1 FILLER_62_2358 ();
 sg13g2_fill_2 FILLER_62_2362 ();
 sg13g2_fill_2 FILLER_62_2394 ();
 sg13g2_fill_2 FILLER_62_2422 ();
 sg13g2_fill_2 FILLER_62_2450 ();
 sg13g2_fill_1 FILLER_62_2521 ();
 sg13g2_fill_1 FILLER_62_2573 ();
 sg13g2_fill_1 FILLER_62_2612 ();
 sg13g2_fill_1 FILLER_62_2641 ();
 sg13g2_fill_2 FILLER_62_2668 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_4 FILLER_63_7 ();
 sg13g2_fill_2 FILLER_63_11 ();
 sg13g2_decap_4 FILLER_63_17 ();
 sg13g2_fill_2 FILLER_63_21 ();
 sg13g2_fill_2 FILLER_63_59 ();
 sg13g2_fill_1 FILLER_63_104 ();
 sg13g2_fill_1 FILLER_63_111 ();
 sg13g2_decap_8 FILLER_63_143 ();
 sg13g2_fill_2 FILLER_63_196 ();
 sg13g2_fill_1 FILLER_63_222 ();
 sg13g2_fill_1 FILLER_63_229 ();
 sg13g2_fill_1 FILLER_63_237 ();
 sg13g2_fill_1 FILLER_63_275 ();
 sg13g2_fill_2 FILLER_63_280 ();
 sg13g2_fill_2 FILLER_63_287 ();
 sg13g2_fill_1 FILLER_63_289 ();
 sg13g2_decap_8 FILLER_63_324 ();
 sg13g2_decap_4 FILLER_63_331 ();
 sg13g2_fill_2 FILLER_63_335 ();
 sg13g2_fill_2 FILLER_63_341 ();
 sg13g2_fill_1 FILLER_63_343 ();
 sg13g2_fill_2 FILLER_63_354 ();
 sg13g2_fill_1 FILLER_63_356 ();
 sg13g2_decap_8 FILLER_63_366 ();
 sg13g2_decap_4 FILLER_63_373 ();
 sg13g2_fill_1 FILLER_63_377 ();
 sg13g2_fill_1 FILLER_63_389 ();
 sg13g2_fill_1 FILLER_63_396 ();
 sg13g2_fill_1 FILLER_63_445 ();
 sg13g2_fill_2 FILLER_63_485 ();
 sg13g2_fill_2 FILLER_63_513 ();
 sg13g2_fill_1 FILLER_63_529 ();
 sg13g2_fill_2 FILLER_63_539 ();
 sg13g2_fill_2 FILLER_63_546 ();
 sg13g2_fill_2 FILLER_63_557 ();
 sg13g2_fill_1 FILLER_63_559 ();
 sg13g2_decap_4 FILLER_63_600 ();
 sg13g2_decap_8 FILLER_63_608 ();
 sg13g2_decap_4 FILLER_63_615 ();
 sg13g2_fill_2 FILLER_63_619 ();
 sg13g2_decap_4 FILLER_63_626 ();
 sg13g2_fill_1 FILLER_63_649 ();
 sg13g2_decap_8 FILLER_63_690 ();
 sg13g2_decap_8 FILLER_63_697 ();
 sg13g2_fill_2 FILLER_63_780 ();
 sg13g2_fill_2 FILLER_63_790 ();
 sg13g2_fill_2 FILLER_63_854 ();
 sg13g2_fill_1 FILLER_63_898 ();
 sg13g2_fill_1 FILLER_63_907 ();
 sg13g2_fill_1 FILLER_63_934 ();
 sg13g2_fill_1 FILLER_63_940 ();
 sg13g2_fill_1 FILLER_63_945 ();
 sg13g2_decap_8 FILLER_63_977 ();
 sg13g2_decap_8 FILLER_63_984 ();
 sg13g2_decap_8 FILLER_63_991 ();
 sg13g2_fill_1 FILLER_63_998 ();
 sg13g2_fill_2 FILLER_63_1003 ();
 sg13g2_fill_1 FILLER_63_1005 ();
 sg13g2_decap_4 FILLER_63_1021 ();
 sg13g2_fill_2 FILLER_63_1025 ();
 sg13g2_fill_2 FILLER_63_1035 ();
 sg13g2_decap_4 FILLER_63_1047 ();
 sg13g2_fill_1 FILLER_63_1051 ();
 sg13g2_decap_8 FILLER_63_1056 ();
 sg13g2_fill_2 FILLER_63_1063 ();
 sg13g2_decap_4 FILLER_63_1068 ();
 sg13g2_decap_8 FILLER_63_1076 ();
 sg13g2_decap_4 FILLER_63_1083 ();
 sg13g2_fill_2 FILLER_63_1087 ();
 sg13g2_decap_8 FILLER_63_1093 ();
 sg13g2_decap_4 FILLER_63_1100 ();
 sg13g2_fill_2 FILLER_63_1104 ();
 sg13g2_decap_4 FILLER_63_1160 ();
 sg13g2_fill_2 FILLER_63_1164 ();
 sg13g2_fill_1 FILLER_63_1202 ();
 sg13g2_fill_2 FILLER_63_1228 ();
 sg13g2_fill_1 FILLER_63_1240 ();
 sg13g2_fill_2 FILLER_63_1263 ();
 sg13g2_fill_1 FILLER_63_1265 ();
 sg13g2_fill_2 FILLER_63_1300 ();
 sg13g2_fill_1 FILLER_63_1307 ();
 sg13g2_decap_4 FILLER_63_1313 ();
 sg13g2_decap_8 FILLER_63_1325 ();
 sg13g2_decap_4 FILLER_63_1332 ();
 sg13g2_fill_2 FILLER_63_1340 ();
 sg13g2_fill_2 FILLER_63_1347 ();
 sg13g2_fill_1 FILLER_63_1349 ();
 sg13g2_fill_2 FILLER_63_1363 ();
 sg13g2_fill_2 FILLER_63_1373 ();
 sg13g2_fill_1 FILLER_63_1375 ();
 sg13g2_fill_1 FILLER_63_1381 ();
 sg13g2_fill_1 FILLER_63_1392 ();
 sg13g2_fill_1 FILLER_63_1398 ();
 sg13g2_fill_2 FILLER_63_1414 ();
 sg13g2_fill_2 FILLER_63_1435 ();
 sg13g2_fill_1 FILLER_63_1437 ();
 sg13g2_decap_8 FILLER_63_1453 ();
 sg13g2_fill_1 FILLER_63_1460 ();
 sg13g2_fill_2 FILLER_63_1470 ();
 sg13g2_fill_1 FILLER_63_1472 ();
 sg13g2_decap_8 FILLER_63_1503 ();
 sg13g2_decap_8 FILLER_63_1510 ();
 sg13g2_fill_2 FILLER_63_1517 ();
 sg13g2_fill_1 FILLER_63_1519 ();
 sg13g2_fill_1 FILLER_63_1529 ();
 sg13g2_fill_2 FILLER_63_1541 ();
 sg13g2_fill_2 FILLER_63_1551 ();
 sg13g2_decap_8 FILLER_63_1573 ();
 sg13g2_decap_8 FILLER_63_1580 ();
 sg13g2_decap_4 FILLER_63_1599 ();
 sg13g2_fill_2 FILLER_63_1603 ();
 sg13g2_decap_4 FILLER_63_1617 ();
 sg13g2_fill_1 FILLER_63_1642 ();
 sg13g2_fill_1 FILLER_63_1653 ();
 sg13g2_fill_2 FILLER_63_1663 ();
 sg13g2_fill_1 FILLER_63_1674 ();
 sg13g2_decap_4 FILLER_63_1680 ();
 sg13g2_fill_2 FILLER_63_1684 ();
 sg13g2_fill_1 FILLER_63_1690 ();
 sg13g2_fill_1 FILLER_63_1703 ();
 sg13g2_fill_1 FILLER_63_1708 ();
 sg13g2_fill_1 FILLER_63_1713 ();
 sg13g2_fill_1 FILLER_63_1719 ();
 sg13g2_fill_1 FILLER_63_1724 ();
 sg13g2_fill_1 FILLER_63_1729 ();
 sg13g2_fill_1 FILLER_63_1745 ();
 sg13g2_fill_1 FILLER_63_1750 ();
 sg13g2_fill_2 FILLER_63_1762 ();
 sg13g2_fill_2 FILLER_63_1783 ();
 sg13g2_decap_4 FILLER_63_1794 ();
 sg13g2_decap_8 FILLER_63_1802 ();
 sg13g2_decap_4 FILLER_63_1809 ();
 sg13g2_fill_1 FILLER_63_1817 ();
 sg13g2_decap_8 FILLER_63_1823 ();
 sg13g2_decap_8 FILLER_63_1830 ();
 sg13g2_decap_4 FILLER_63_1841 ();
 sg13g2_decap_8 FILLER_63_1856 ();
 sg13g2_fill_1 FILLER_63_1880 ();
 sg13g2_decap_8 FILLER_63_1898 ();
 sg13g2_decap_8 FILLER_63_1905 ();
 sg13g2_decap_4 FILLER_63_1912 ();
 sg13g2_fill_2 FILLER_63_1916 ();
 sg13g2_fill_1 FILLER_63_1956 ();
 sg13g2_fill_1 FILLER_63_1963 ();
 sg13g2_fill_1 FILLER_63_1970 ();
 sg13g2_fill_1 FILLER_63_1975 ();
 sg13g2_fill_1 FILLER_63_1981 ();
 sg13g2_fill_2 FILLER_63_1987 ();
 sg13g2_fill_2 FILLER_63_2019 ();
 sg13g2_fill_1 FILLER_63_2041 ();
 sg13g2_fill_1 FILLER_63_2046 ();
 sg13g2_fill_1 FILLER_63_2068 ();
 sg13g2_fill_2 FILLER_63_2090 ();
 sg13g2_fill_1 FILLER_63_2092 ();
 sg13g2_decap_4 FILLER_63_2176 ();
 sg13g2_fill_2 FILLER_63_2180 ();
 sg13g2_decap_4 FILLER_63_2190 ();
 sg13g2_fill_2 FILLER_63_2194 ();
 sg13g2_fill_1 FILLER_63_2206 ();
 sg13g2_decap_4 FILLER_63_2256 ();
 sg13g2_fill_2 FILLER_63_2260 ();
 sg13g2_fill_1 FILLER_63_2270 ();
 sg13g2_fill_1 FILLER_63_2296 ();
 sg13g2_fill_1 FILLER_63_2324 ();
 sg13g2_fill_2 FILLER_63_2330 ();
 sg13g2_fill_2 FILLER_63_2344 ();
 sg13g2_fill_2 FILLER_63_2494 ();
 sg13g2_fill_1 FILLER_63_2533 ();
 sg13g2_fill_2 FILLER_63_2549 ();
 sg13g2_fill_1 FILLER_63_2558 ();
 sg13g2_fill_1 FILLER_63_2636 ();
 sg13g2_fill_2 FILLER_63_2667 ();
 sg13g2_fill_1 FILLER_63_2669 ();
 sg13g2_decap_4 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_4 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_fill_2 FILLER_64_109 ();
 sg13g2_fill_2 FILLER_64_121 ();
 sg13g2_fill_1 FILLER_64_123 ();
 sg13g2_fill_1 FILLER_64_133 ();
 sg13g2_fill_2 FILLER_64_148 ();
 sg13g2_fill_1 FILLER_64_150 ();
 sg13g2_fill_2 FILLER_64_160 ();
 sg13g2_fill_1 FILLER_64_172 ();
 sg13g2_fill_2 FILLER_64_177 ();
 sg13g2_fill_2 FILLER_64_253 ();
 sg13g2_fill_1 FILLER_64_312 ();
 sg13g2_decap_8 FILLER_64_317 ();
 sg13g2_fill_2 FILLER_64_324 ();
 sg13g2_fill_2 FILLER_64_356 ();
 sg13g2_fill_2 FILLER_64_449 ();
 sg13g2_fill_2 FILLER_64_463 ();
 sg13g2_fill_1 FILLER_64_476 ();
 sg13g2_decap_8 FILLER_64_482 ();
 sg13g2_fill_2 FILLER_64_489 ();
 sg13g2_decap_4 FILLER_64_495 ();
 sg13g2_decap_4 FILLER_64_523 ();
 sg13g2_fill_2 FILLER_64_527 ();
 sg13g2_fill_1 FILLER_64_538 ();
 sg13g2_decap_8 FILLER_64_543 ();
 sg13g2_decap_4 FILLER_64_550 ();
 sg13g2_fill_2 FILLER_64_554 ();
 sg13g2_fill_1 FILLER_64_582 ();
 sg13g2_fill_2 FILLER_64_602 ();
 sg13g2_decap_8 FILLER_64_609 ();
 sg13g2_decap_4 FILLER_64_639 ();
 sg13g2_decap_8 FILLER_64_647 ();
 sg13g2_fill_2 FILLER_64_654 ();
 sg13g2_fill_1 FILLER_64_656 ();
 sg13g2_decap_8 FILLER_64_682 ();
 sg13g2_decap_8 FILLER_64_689 ();
 sg13g2_fill_1 FILLER_64_700 ();
 sg13g2_fill_1 FILLER_64_706 ();
 sg13g2_fill_1 FILLER_64_721 ();
 sg13g2_fill_2 FILLER_64_738 ();
 sg13g2_fill_1 FILLER_64_749 ();
 sg13g2_fill_1 FILLER_64_769 ();
 sg13g2_fill_2 FILLER_64_806 ();
 sg13g2_fill_1 FILLER_64_858 ();
 sg13g2_fill_2 FILLER_64_881 ();
 sg13g2_fill_1 FILLER_64_883 ();
 sg13g2_decap_8 FILLER_64_953 ();
 sg13g2_fill_2 FILLER_64_965 ();
 sg13g2_fill_1 FILLER_64_974 ();
 sg13g2_decap_4 FILLER_64_990 ();
 sg13g2_fill_1 FILLER_64_994 ();
 sg13g2_fill_2 FILLER_64_1030 ();
 sg13g2_decap_4 FILLER_64_1037 ();
 sg13g2_decap_8 FILLER_64_1050 ();
 sg13g2_fill_1 FILLER_64_1057 ();
 sg13g2_decap_8 FILLER_64_1108 ();
 sg13g2_decap_4 FILLER_64_1115 ();
 sg13g2_fill_2 FILLER_64_1119 ();
 sg13g2_fill_1 FILLER_64_1155 ();
 sg13g2_fill_1 FILLER_64_1164 ();
 sg13g2_fill_2 FILLER_64_1168 ();
 sg13g2_fill_1 FILLER_64_1174 ();
 sg13g2_fill_2 FILLER_64_1185 ();
 sg13g2_fill_2 FILLER_64_1213 ();
 sg13g2_decap_8 FILLER_64_1236 ();
 sg13g2_decap_8 FILLER_64_1243 ();
 sg13g2_decap_4 FILLER_64_1250 ();
 sg13g2_fill_1 FILLER_64_1261 ();
 sg13g2_fill_1 FILLER_64_1266 ();
 sg13g2_fill_2 FILLER_64_1284 ();
 sg13g2_fill_1 FILLER_64_1291 ();
 sg13g2_fill_1 FILLER_64_1296 ();
 sg13g2_fill_1 FILLER_64_1302 ();
 sg13g2_decap_8 FILLER_64_1316 ();
 sg13g2_decap_4 FILLER_64_1323 ();
 sg13g2_fill_1 FILLER_64_1332 ();
 sg13g2_fill_2 FILLER_64_1338 ();
 sg13g2_decap_4 FILLER_64_1351 ();
 sg13g2_fill_1 FILLER_64_1381 ();
 sg13g2_fill_2 FILLER_64_1399 ();
 sg13g2_fill_1 FILLER_64_1401 ();
 sg13g2_decap_8 FILLER_64_1407 ();
 sg13g2_decap_4 FILLER_64_1414 ();
 sg13g2_fill_1 FILLER_64_1428 ();
 sg13g2_decap_4 FILLER_64_1445 ();
 sg13g2_decap_8 FILLER_64_1458 ();
 sg13g2_decap_8 FILLER_64_1465 ();
 sg13g2_decap_8 FILLER_64_1472 ();
 sg13g2_decap_4 FILLER_64_1479 ();
 sg13g2_fill_1 FILLER_64_1483 ();
 sg13g2_decap_8 FILLER_64_1488 ();
 sg13g2_decap_8 FILLER_64_1495 ();
 sg13g2_fill_2 FILLER_64_1502 ();
 sg13g2_fill_1 FILLER_64_1504 ();
 sg13g2_decap_4 FILLER_64_1509 ();
 sg13g2_fill_1 FILLER_64_1534 ();
 sg13g2_fill_2 FILLER_64_1538 ();
 sg13g2_fill_2 FILLER_64_1561 ();
 sg13g2_fill_1 FILLER_64_1605 ();
 sg13g2_fill_1 FILLER_64_1628 ();
 sg13g2_fill_2 FILLER_64_1656 ();
 sg13g2_fill_1 FILLER_64_1658 ();
 sg13g2_decap_8 FILLER_64_1673 ();
 sg13g2_fill_1 FILLER_64_1680 ();
 sg13g2_fill_2 FILLER_64_1685 ();
 sg13g2_fill_1 FILLER_64_1687 ();
 sg13g2_fill_1 FILLER_64_1721 ();
 sg13g2_fill_1 FILLER_64_1727 ();
 sg13g2_fill_1 FILLER_64_1733 ();
 sg13g2_fill_2 FILLER_64_1764 ();
 sg13g2_decap_8 FILLER_64_1769 ();
 sg13g2_decap_8 FILLER_64_1776 ();
 sg13g2_fill_2 FILLER_64_1783 ();
 sg13g2_fill_1 FILLER_64_1785 ();
 sg13g2_decap_8 FILLER_64_1816 ();
 sg13g2_decap_8 FILLER_64_1823 ();
 sg13g2_decap_8 FILLER_64_1830 ();
 sg13g2_decap_8 FILLER_64_1837 ();
 sg13g2_fill_2 FILLER_64_1844 ();
 sg13g2_fill_1 FILLER_64_1846 ();
 sg13g2_decap_8 FILLER_64_1858 ();
 sg13g2_fill_1 FILLER_64_1865 ();
 sg13g2_decap_8 FILLER_64_1910 ();
 sg13g2_fill_1 FILLER_64_1927 ();
 sg13g2_fill_1 FILLER_64_1932 ();
 sg13g2_fill_1 FILLER_64_1948 ();
 sg13g2_decap_8 FILLER_64_1954 ();
 sg13g2_fill_2 FILLER_64_1969 ();
 sg13g2_fill_1 FILLER_64_1989 ();
 sg13g2_fill_1 FILLER_64_2019 ();
 sg13g2_fill_2 FILLER_64_2024 ();
 sg13g2_fill_1 FILLER_64_2042 ();
 sg13g2_fill_2 FILLER_64_2049 ();
 sg13g2_fill_2 FILLER_64_2080 ();
 sg13g2_fill_1 FILLER_64_2175 ();
 sg13g2_fill_2 FILLER_64_2202 ();
 sg13g2_fill_2 FILLER_64_2230 ();
 sg13g2_fill_1 FILLER_64_2232 ();
 sg13g2_decap_4 FILLER_64_2259 ();
 sg13g2_fill_1 FILLER_64_2263 ();
 sg13g2_fill_1 FILLER_64_2304 ();
 sg13g2_decap_4 FILLER_64_2361 ();
 sg13g2_fill_1 FILLER_64_2365 ();
 sg13g2_fill_1 FILLER_64_2435 ();
 sg13g2_decap_4 FILLER_64_2445 ();
 sg13g2_decap_8 FILLER_64_2454 ();
 sg13g2_fill_1 FILLER_64_2466 ();
 sg13g2_fill_2 FILLER_64_2479 ();
 sg13g2_decap_4 FILLER_64_2487 ();
 sg13g2_fill_1 FILLER_64_2491 ();
 sg13g2_decap_4 FILLER_64_2509 ();
 sg13g2_fill_2 FILLER_64_2519 ();
 sg13g2_fill_1 FILLER_64_2554 ();
 sg13g2_decap_8 FILLER_64_2565 ();
 sg13g2_fill_2 FILLER_64_2585 ();
 sg13g2_fill_2 FILLER_64_2591 ();
 sg13g2_fill_2 FILLER_64_2606 ();
 sg13g2_fill_1 FILLER_64_2614 ();
 sg13g2_fill_2 FILLER_64_2625 ();
 sg13g2_decap_8 FILLER_64_2657 ();
 sg13g2_decap_4 FILLER_64_2664 ();
 sg13g2_fill_2 FILLER_64_2668 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_28 ();
 sg13g2_fill_1 FILLER_65_30 ();
 sg13g2_decap_4 FILLER_65_35 ();
 sg13g2_fill_1 FILLER_65_39 ();
 sg13g2_decap_4 FILLER_65_50 ();
 sg13g2_fill_1 FILLER_65_54 ();
 sg13g2_fill_2 FILLER_65_65 ();
 sg13g2_fill_1 FILLER_65_67 ();
 sg13g2_decap_4 FILLER_65_72 ();
 sg13g2_decap_8 FILLER_65_85 ();
 sg13g2_decap_8 FILLER_65_92 ();
 sg13g2_fill_1 FILLER_65_99 ();
 sg13g2_decap_8 FILLER_65_115 ();
 sg13g2_decap_8 FILLER_65_122 ();
 sg13g2_fill_2 FILLER_65_129 ();
 sg13g2_fill_1 FILLER_65_131 ();
 sg13g2_fill_1 FILLER_65_136 ();
 sg13g2_fill_1 FILLER_65_163 ();
 sg13g2_fill_1 FILLER_65_185 ();
 sg13g2_fill_2 FILLER_65_210 ();
 sg13g2_fill_1 FILLER_65_212 ();
 sg13g2_decap_4 FILLER_65_217 ();
 sg13g2_decap_4 FILLER_65_225 ();
 sg13g2_fill_1 FILLER_65_260 ();
 sg13g2_fill_1 FILLER_65_265 ();
 sg13g2_fill_1 FILLER_65_288 ();
 sg13g2_fill_1 FILLER_65_293 ();
 sg13g2_fill_1 FILLER_65_303 ();
 sg13g2_fill_1 FILLER_65_330 ();
 sg13g2_fill_1 FILLER_65_345 ();
 sg13g2_fill_2 FILLER_65_356 ();
 sg13g2_fill_1 FILLER_65_398 ();
 sg13g2_fill_2 FILLER_65_402 ();
 sg13g2_fill_2 FILLER_65_416 ();
 sg13g2_fill_1 FILLER_65_449 ();
 sg13g2_fill_2 FILLER_65_476 ();
 sg13g2_fill_2 FILLER_65_484 ();
 sg13g2_decap_4 FILLER_65_492 ();
 sg13g2_fill_2 FILLER_65_496 ();
 sg13g2_fill_1 FILLER_65_513 ();
 sg13g2_decap_4 FILLER_65_549 ();
 sg13g2_fill_2 FILLER_65_553 ();
 sg13g2_decap_4 FILLER_65_630 ();
 sg13g2_fill_2 FILLER_65_638 ();
 sg13g2_fill_1 FILLER_65_655 ();
 sg13g2_fill_1 FILLER_65_661 ();
 sg13g2_decap_8 FILLER_65_672 ();
 sg13g2_decap_8 FILLER_65_679 ();
 sg13g2_decap_4 FILLER_65_686 ();
 sg13g2_fill_1 FILLER_65_690 ();
 sg13g2_fill_1 FILLER_65_717 ();
 sg13g2_fill_1 FILLER_65_756 ();
 sg13g2_fill_2 FILLER_65_769 ();
 sg13g2_fill_1 FILLER_65_779 ();
 sg13g2_fill_1 FILLER_65_803 ();
 sg13g2_fill_2 FILLER_65_813 ();
 sg13g2_fill_1 FILLER_65_815 ();
 sg13g2_fill_1 FILLER_65_835 ();
 sg13g2_fill_2 FILLER_65_843 ();
 sg13g2_decap_8 FILLER_65_849 ();
 sg13g2_decap_8 FILLER_65_856 ();
 sg13g2_fill_1 FILLER_65_863 ();
 sg13g2_fill_2 FILLER_65_896 ();
 sg13g2_fill_2 FILLER_65_938 ();
 sg13g2_fill_1 FILLER_65_949 ();
 sg13g2_fill_1 FILLER_65_963 ();
 sg13g2_fill_1 FILLER_65_974 ();
 sg13g2_fill_2 FILLER_65_1021 ();
 sg13g2_fill_1 FILLER_65_1023 ();
 sg13g2_fill_1 FILLER_65_1032 ();
 sg13g2_fill_2 FILLER_65_1059 ();
 sg13g2_fill_2 FILLER_65_1064 ();
 sg13g2_fill_2 FILLER_65_1092 ();
 sg13g2_fill_1 FILLER_65_1120 ();
 sg13g2_decap_4 FILLER_65_1125 ();
 sg13g2_fill_2 FILLER_65_1129 ();
 sg13g2_decap_8 FILLER_65_1139 ();
 sg13g2_decap_8 FILLER_65_1146 ();
 sg13g2_fill_2 FILLER_65_1153 ();
 sg13g2_decap_4 FILLER_65_1175 ();
 sg13g2_decap_8 FILLER_65_1183 ();
 sg13g2_fill_2 FILLER_65_1190 ();
 sg13g2_fill_1 FILLER_65_1192 ();
 sg13g2_decap_8 FILLER_65_1197 ();
 sg13g2_decap_8 FILLER_65_1235 ();
 sg13g2_decap_4 FILLER_65_1242 ();
 sg13g2_fill_2 FILLER_65_1261 ();
 sg13g2_fill_2 FILLER_65_1296 ();
 sg13g2_decap_4 FILLER_65_1313 ();
 sg13g2_fill_1 FILLER_65_1317 ();
 sg13g2_decap_4 FILLER_65_1368 ();
 sg13g2_fill_1 FILLER_65_1386 ();
 sg13g2_fill_1 FILLER_65_1402 ();
 sg13g2_fill_1 FILLER_65_1408 ();
 sg13g2_decap_8 FILLER_65_1416 ();
 sg13g2_fill_2 FILLER_65_1423 ();
 sg13g2_fill_1 FILLER_65_1429 ();
 sg13g2_decap_4 FILLER_65_1451 ();
 sg13g2_fill_2 FILLER_65_1455 ();
 sg13g2_decap_4 FILLER_65_1467 ();
 sg13g2_decap_8 FILLER_65_1484 ();
 sg13g2_decap_8 FILLER_65_1491 ();
 sg13g2_fill_2 FILLER_65_1498 ();
 sg13g2_fill_1 FILLER_65_1500 ();
 sg13g2_fill_1 FILLER_65_1505 ();
 sg13g2_fill_1 FILLER_65_1595 ();
 sg13g2_fill_1 FILLER_65_1620 ();
 sg13g2_decap_4 FILLER_65_1624 ();
 sg13g2_fill_1 FILLER_65_1641 ();
 sg13g2_fill_2 FILLER_65_1649 ();
 sg13g2_fill_1 FILLER_65_1651 ();
 sg13g2_fill_2 FILLER_65_1657 ();
 sg13g2_fill_1 FILLER_65_1659 ();
 sg13g2_decap_8 FILLER_65_1675 ();
 sg13g2_fill_2 FILLER_65_1691 ();
 sg13g2_fill_1 FILLER_65_1738 ();
 sg13g2_fill_1 FILLER_65_1775 ();
 sg13g2_fill_2 FILLER_65_1781 ();
 sg13g2_fill_1 FILLER_65_1805 ();
 sg13g2_decap_8 FILLER_65_1810 ();
 sg13g2_decap_8 FILLER_65_1826 ();
 sg13g2_decap_4 FILLER_65_1833 ();
 sg13g2_fill_2 FILLER_65_1842 ();
 sg13g2_fill_1 FILLER_65_1844 ();
 sg13g2_decap_4 FILLER_65_1849 ();
 sg13g2_decap_8 FILLER_65_1857 ();
 sg13g2_decap_4 FILLER_65_1864 ();
 sg13g2_fill_1 FILLER_65_1868 ();
 sg13g2_decap_8 FILLER_65_1886 ();
 sg13g2_fill_1 FILLER_65_1893 ();
 sg13g2_fill_2 FILLER_65_1913 ();
 sg13g2_fill_1 FILLER_65_1915 ();
 sg13g2_fill_2 FILLER_65_1962 ();
 sg13g2_fill_1 FILLER_65_1964 ();
 sg13g2_fill_1 FILLER_65_1970 ();
 sg13g2_fill_1 FILLER_65_1975 ();
 sg13g2_fill_1 FILLER_65_1982 ();
 sg13g2_fill_1 FILLER_65_1989 ();
 sg13g2_fill_1 FILLER_65_2000 ();
 sg13g2_fill_2 FILLER_65_2006 ();
 sg13g2_fill_1 FILLER_65_2014 ();
 sg13g2_fill_2 FILLER_65_2019 ();
 sg13g2_fill_1 FILLER_65_2021 ();
 sg13g2_decap_4 FILLER_65_2026 ();
 sg13g2_fill_2 FILLER_65_2030 ();
 sg13g2_fill_1 FILLER_65_2038 ();
 sg13g2_fill_2 FILLER_65_2094 ();
 sg13g2_fill_1 FILLER_65_2096 ();
 sg13g2_fill_2 FILLER_65_2133 ();
 sg13g2_decap_4 FILLER_65_2161 ();
 sg13g2_fill_2 FILLER_65_2165 ();
 sg13g2_decap_8 FILLER_65_2193 ();
 sg13g2_decap_4 FILLER_65_2200 ();
 sg13g2_fill_2 FILLER_65_2204 ();
 sg13g2_fill_2 FILLER_65_2216 ();
 sg13g2_fill_1 FILLER_65_2218 ();
 sg13g2_fill_1 FILLER_65_2255 ();
 sg13g2_fill_2 FILLER_65_2300 ();
 sg13g2_fill_1 FILLER_65_2308 ();
 sg13g2_fill_2 FILLER_65_2320 ();
 sg13g2_fill_2 FILLER_65_2332 ();
 sg13g2_decap_4 FILLER_65_2364 ();
 sg13g2_fill_2 FILLER_65_2368 ();
 sg13g2_fill_1 FILLER_65_2376 ();
 sg13g2_decap_8 FILLER_65_2415 ();
 sg13g2_decap_8 FILLER_65_2422 ();
 sg13g2_decap_4 FILLER_65_2433 ();
 sg13g2_fill_2 FILLER_65_2437 ();
 sg13g2_fill_1 FILLER_65_2444 ();
 sg13g2_fill_2 FILLER_65_2449 ();
 sg13g2_fill_1 FILLER_65_2456 ();
 sg13g2_fill_2 FILLER_65_2462 ();
 sg13g2_fill_1 FILLER_65_2464 ();
 sg13g2_fill_2 FILLER_65_2469 ();
 sg13g2_fill_1 FILLER_65_2471 ();
 sg13g2_decap_8 FILLER_65_2502 ();
 sg13g2_decap_8 FILLER_65_2509 ();
 sg13g2_fill_2 FILLER_65_2516 ();
 sg13g2_decap_8 FILLER_65_2521 ();
 sg13g2_decap_8 FILLER_65_2567 ();
 sg13g2_decap_8 FILLER_65_2574 ();
 sg13g2_decap_4 FILLER_65_2581 ();
 sg13g2_fill_1 FILLER_65_2585 ();
 sg13g2_fill_2 FILLER_65_2646 ();
 sg13g2_fill_1 FILLER_65_2648 ();
 sg13g2_decap_8 FILLER_65_2653 ();
 sg13g2_decap_8 FILLER_65_2660 ();
 sg13g2_fill_2 FILLER_65_2667 ();
 sg13g2_fill_1 FILLER_65_2669 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_7 ();
 sg13g2_fill_2 FILLER_66_15 ();
 sg13g2_decap_4 FILLER_66_53 ();
 sg13g2_fill_2 FILLER_66_57 ();
 sg13g2_fill_2 FILLER_66_103 ();
 sg13g2_fill_2 FILLER_66_131 ();
 sg13g2_fill_1 FILLER_66_133 ();
 sg13g2_fill_1 FILLER_66_138 ();
 sg13g2_fill_2 FILLER_66_165 ();
 sg13g2_fill_1 FILLER_66_167 ();
 sg13g2_fill_1 FILLER_66_198 ();
 sg13g2_decap_8 FILLER_66_230 ();
 sg13g2_decap_4 FILLER_66_237 ();
 sg13g2_fill_2 FILLER_66_241 ();
 sg13g2_fill_2 FILLER_66_246 ();
 sg13g2_fill_1 FILLER_66_278 ();
 sg13g2_decap_4 FILLER_66_327 ();
 sg13g2_fill_1 FILLER_66_331 ();
 sg13g2_fill_1 FILLER_66_340 ();
 sg13g2_fill_2 FILLER_66_367 ();
 sg13g2_fill_1 FILLER_66_369 ();
 sg13g2_decap_4 FILLER_66_376 ();
 sg13g2_decap_8 FILLER_66_384 ();
 sg13g2_decap_4 FILLER_66_391 ();
 sg13g2_fill_1 FILLER_66_395 ();
 sg13g2_decap_8 FILLER_66_407 ();
 sg13g2_decap_4 FILLER_66_427 ();
 sg13g2_fill_2 FILLER_66_431 ();
 sg13g2_decap_4 FILLER_66_437 ();
 sg13g2_fill_2 FILLER_66_441 ();
 sg13g2_fill_1 FILLER_66_507 ();
 sg13g2_fill_2 FILLER_66_527 ();
 sg13g2_fill_1 FILLER_66_529 ();
 sg13g2_decap_8 FILLER_66_539 ();
 sg13g2_decap_8 FILLER_66_546 ();
 sg13g2_decap_8 FILLER_66_553 ();
 sg13g2_fill_1 FILLER_66_560 ();
 sg13g2_decap_4 FILLER_66_566 ();
 sg13g2_fill_1 FILLER_66_570 ();
 sg13g2_fill_2 FILLER_66_586 ();
 sg13g2_fill_1 FILLER_66_588 ();
 sg13g2_fill_1 FILLER_66_607 ();
 sg13g2_fill_1 FILLER_66_612 ();
 sg13g2_fill_1 FILLER_66_643 ();
 sg13g2_fill_1 FILLER_66_654 ();
 sg13g2_decap_4 FILLER_66_681 ();
 sg13g2_fill_1 FILLER_66_685 ();
 sg13g2_fill_1 FILLER_66_692 ();
 sg13g2_fill_1 FILLER_66_778 ();
 sg13g2_decap_8 FILLER_66_805 ();
 sg13g2_decap_8 FILLER_66_850 ();
 sg13g2_decap_8 FILLER_66_857 ();
 sg13g2_fill_2 FILLER_66_864 ();
 sg13g2_fill_1 FILLER_66_866 ();
 sg13g2_decap_8 FILLER_66_877 ();
 sg13g2_fill_2 FILLER_66_884 ();
 sg13g2_fill_1 FILLER_66_896 ();
 sg13g2_fill_2 FILLER_66_907 ();
 sg13g2_fill_2 FILLER_66_929 ();
 sg13g2_decap_4 FILLER_66_957 ();
 sg13g2_fill_1 FILLER_66_961 ();
 sg13g2_fill_2 FILLER_66_966 ();
 sg13g2_fill_2 FILLER_66_994 ();
 sg13g2_fill_2 FILLER_66_1030 ();
 sg13g2_fill_2 FILLER_66_1044 ();
 sg13g2_fill_1 FILLER_66_1046 ();
 sg13g2_decap_4 FILLER_66_1053 ();
 sg13g2_fill_1 FILLER_66_1057 ();
 sg13g2_fill_2 FILLER_66_1064 ();
 sg13g2_fill_2 FILLER_66_1093 ();
 sg13g2_decap_8 FILLER_66_1121 ();
 sg13g2_decap_4 FILLER_66_1128 ();
 sg13g2_fill_2 FILLER_66_1132 ();
 sg13g2_decap_4 FILLER_66_1168 ();
 sg13g2_fill_2 FILLER_66_1172 ();
 sg13g2_fill_2 FILLER_66_1218 ();
 sg13g2_fill_1 FILLER_66_1220 ();
 sg13g2_fill_2 FILLER_66_1268 ();
 sg13g2_fill_1 FILLER_66_1270 ();
 sg13g2_fill_1 FILLER_66_1276 ();
 sg13g2_fill_1 FILLER_66_1285 ();
 sg13g2_fill_2 FILLER_66_1292 ();
 sg13g2_decap_4 FILLER_66_1299 ();
 sg13g2_decap_4 FILLER_66_1311 ();
 sg13g2_fill_2 FILLER_66_1320 ();
 sg13g2_fill_1 FILLER_66_1322 ();
 sg13g2_decap_8 FILLER_66_1338 ();
 sg13g2_decap_4 FILLER_66_1345 ();
 sg13g2_fill_1 FILLER_66_1349 ();
 sg13g2_fill_2 FILLER_66_1358 ();
 sg13g2_fill_1 FILLER_66_1409 ();
 sg13g2_fill_2 FILLER_66_1415 ();
 sg13g2_fill_1 FILLER_66_1440 ();
 sg13g2_fill_1 FILLER_66_1449 ();
 sg13g2_fill_1 FILLER_66_1460 ();
 sg13g2_decap_4 FILLER_66_1487 ();
 sg13g2_fill_2 FILLER_66_1491 ();
 sg13g2_fill_2 FILLER_66_1530 ();
 sg13g2_fill_2 FILLER_66_1538 ();
 sg13g2_fill_1 FILLER_66_1558 ();
 sg13g2_fill_2 FILLER_66_1582 ();
 sg13g2_decap_8 FILLER_66_1603 ();
 sg13g2_fill_1 FILLER_66_1610 ();
 sg13g2_fill_2 FILLER_66_1615 ();
 sg13g2_fill_1 FILLER_66_1630 ();
 sg13g2_fill_2 FILLER_66_1635 ();
 sg13g2_fill_1 FILLER_66_1642 ();
 sg13g2_fill_1 FILLER_66_1649 ();
 sg13g2_decap_4 FILLER_66_1680 ();
 sg13g2_fill_1 FILLER_66_1684 ();
 sg13g2_fill_2 FILLER_66_1690 ();
 sg13g2_decap_8 FILLER_66_1696 ();
 sg13g2_fill_1 FILLER_66_1719 ();
 sg13g2_decap_4 FILLER_66_1728 ();
 sg13g2_fill_2 FILLER_66_1732 ();
 sg13g2_decap_4 FILLER_66_1768 ();
 sg13g2_fill_1 FILLER_66_1772 ();
 sg13g2_decap_4 FILLER_66_1818 ();
 sg13g2_fill_2 FILLER_66_1822 ();
 sg13g2_decap_8 FILLER_66_1828 ();
 sg13g2_decap_8 FILLER_66_1835 ();
 sg13g2_fill_2 FILLER_66_1842 ();
 sg13g2_fill_1 FILLER_66_1844 ();
 sg13g2_decap_8 FILLER_66_1859 ();
 sg13g2_fill_2 FILLER_66_1866 ();
 sg13g2_fill_1 FILLER_66_1883 ();
 sg13g2_decap_4 FILLER_66_1888 ();
 sg13g2_fill_2 FILLER_66_1892 ();
 sg13g2_decap_8 FILLER_66_1900 ();
 sg13g2_decap_8 FILLER_66_1907 ();
 sg13g2_decap_4 FILLER_66_1914 ();
 sg13g2_fill_2 FILLER_66_1929 ();
 sg13g2_fill_1 FILLER_66_1931 ();
 sg13g2_decap_4 FILLER_66_1937 ();
 sg13g2_fill_1 FILLER_66_1941 ();
 sg13g2_fill_1 FILLER_66_1960 ();
 sg13g2_decap_4 FILLER_66_1973 ();
 sg13g2_decap_4 FILLER_66_1989 ();
 sg13g2_fill_1 FILLER_66_1993 ();
 sg13g2_fill_2 FILLER_66_2037 ();
 sg13g2_decap_4 FILLER_66_2092 ();
 sg13g2_fill_1 FILLER_66_2099 ();
 sg13g2_decap_8 FILLER_66_2160 ();
 sg13g2_decap_8 FILLER_66_2167 ();
 sg13g2_decap_8 FILLER_66_2178 ();
 sg13g2_fill_1 FILLER_66_2185 ();
 sg13g2_decap_8 FILLER_66_2206 ();
 sg13g2_fill_1 FILLER_66_2239 ();
 sg13g2_decap_4 FILLER_66_2248 ();
 sg13g2_fill_2 FILLER_66_2290 ();
 sg13g2_fill_2 FILLER_66_2370 ();
 sg13g2_fill_1 FILLER_66_2372 ();
 sg13g2_decap_8 FILLER_66_2413 ();
 sg13g2_decap_8 FILLER_66_2420 ();
 sg13g2_decap_8 FILLER_66_2427 ();
 sg13g2_decap_8 FILLER_66_2434 ();
 sg13g2_fill_1 FILLER_66_2441 ();
 sg13g2_fill_1 FILLER_66_2494 ();
 sg13g2_fill_1 FILLER_66_2499 ();
 sg13g2_decap_4 FILLER_66_2514 ();
 sg13g2_fill_2 FILLER_66_2526 ();
 sg13g2_decap_8 FILLER_66_2567 ();
 sg13g2_fill_2 FILLER_66_2574 ();
 sg13g2_fill_1 FILLER_66_2576 ();
 sg13g2_decap_4 FILLER_66_2612 ();
 sg13g2_fill_2 FILLER_66_2640 ();
 sg13g2_fill_2 FILLER_66_2668 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_fill_2 FILLER_67_35 ();
 sg13g2_fill_1 FILLER_67_68 ();
 sg13g2_fill_1 FILLER_67_111 ();
 sg13g2_fill_2 FILLER_67_116 ();
 sg13g2_fill_1 FILLER_67_118 ();
 sg13g2_decap_8 FILLER_67_155 ();
 sg13g2_fill_2 FILLER_67_162 ();
 sg13g2_fill_1 FILLER_67_189 ();
 sg13g2_fill_1 FILLER_67_223 ();
 sg13g2_fill_1 FILLER_67_229 ();
 sg13g2_fill_1 FILLER_67_244 ();
 sg13g2_fill_2 FILLER_67_257 ();
 sg13g2_fill_1 FILLER_67_269 ();
 sg13g2_fill_2 FILLER_67_275 ();
 sg13g2_fill_1 FILLER_67_277 ();
 sg13g2_fill_1 FILLER_67_290 ();
 sg13g2_decap_8 FILLER_67_295 ();
 sg13g2_decap_8 FILLER_67_302 ();
 sg13g2_fill_2 FILLER_67_313 ();
 sg13g2_decap_8 FILLER_67_327 ();
 sg13g2_decap_8 FILLER_67_334 ();
 sg13g2_fill_2 FILLER_67_341 ();
 sg13g2_decap_4 FILLER_67_369 ();
 sg13g2_fill_2 FILLER_67_373 ();
 sg13g2_fill_2 FILLER_67_390 ();
 sg13g2_decap_4 FILLER_67_396 ();
 sg13g2_decap_8 FILLER_67_404 ();
 sg13g2_fill_2 FILLER_67_411 ();
 sg13g2_fill_1 FILLER_67_413 ();
 sg13g2_fill_1 FILLER_67_418 ();
 sg13g2_decap_4 FILLER_67_424 ();
 sg13g2_fill_1 FILLER_67_428 ();
 sg13g2_fill_2 FILLER_67_442 ();
 sg13g2_fill_2 FILLER_67_449 ();
 sg13g2_fill_1 FILLER_67_451 ();
 sg13g2_fill_2 FILLER_67_458 ();
 sg13g2_decap_4 FILLER_67_474 ();
 sg13g2_fill_1 FILLER_67_478 ();
 sg13g2_fill_2 FILLER_67_484 ();
 sg13g2_fill_1 FILLER_67_486 ();
 sg13g2_decap_8 FILLER_67_490 ();
 sg13g2_decap_4 FILLER_67_497 ();
 sg13g2_fill_2 FILLER_67_516 ();
 sg13g2_fill_1 FILLER_67_518 ();
 sg13g2_fill_2 FILLER_67_524 ();
 sg13g2_fill_1 FILLER_67_526 ();
 sg13g2_decap_8 FILLER_67_553 ();
 sg13g2_fill_1 FILLER_67_560 ();
 sg13g2_decap_8 FILLER_67_565 ();
 sg13g2_fill_1 FILLER_67_572 ();
 sg13g2_decap_8 FILLER_67_590 ();
 sg13g2_fill_1 FILLER_67_597 ();
 sg13g2_decap_4 FILLER_67_602 ();
 sg13g2_decap_8 FILLER_67_611 ();
 sg13g2_decap_8 FILLER_67_618 ();
 sg13g2_decap_4 FILLER_67_625 ();
 sg13g2_fill_2 FILLER_67_736 ();
 sg13g2_fill_2 FILLER_67_760 ();
 sg13g2_fill_1 FILLER_67_778 ();
 sg13g2_fill_1 FILLER_67_783 ();
 sg13g2_fill_1 FILLER_67_789 ();
 sg13g2_fill_1 FILLER_67_821 ();
 sg13g2_fill_1 FILLER_67_827 ();
 sg13g2_fill_2 FILLER_67_833 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_fill_2 FILLER_67_888 ();
 sg13g2_fill_2 FILLER_67_922 ();
 sg13g2_fill_1 FILLER_67_939 ();
 sg13g2_fill_1 FILLER_67_944 ();
 sg13g2_fill_1 FILLER_67_971 ();
 sg13g2_decap_8 FILLER_67_998 ();
 sg13g2_fill_2 FILLER_67_1005 ();
 sg13g2_fill_1 FILLER_67_1024 ();
 sg13g2_fill_2 FILLER_67_1051 ();
 sg13g2_decap_4 FILLER_67_1131 ();
 sg13g2_decap_4 FILLER_67_1161 ();
 sg13g2_fill_1 FILLER_67_1165 ();
 sg13g2_fill_2 FILLER_67_1250 ();
 sg13g2_fill_1 FILLER_67_1252 ();
 sg13g2_fill_1 FILLER_67_1269 ();
 sg13g2_fill_2 FILLER_67_1320 ();
 sg13g2_fill_1 FILLER_67_1322 ();
 sg13g2_fill_2 FILLER_67_1334 ();
 sg13g2_fill_1 FILLER_67_1336 ();
 sg13g2_fill_2 FILLER_67_1343 ();
 sg13g2_fill_1 FILLER_67_1345 ();
 sg13g2_decap_4 FILLER_67_1361 ();
 sg13g2_fill_1 FILLER_67_1365 ();
 sg13g2_fill_1 FILLER_67_1374 ();
 sg13g2_fill_2 FILLER_67_1390 ();
 sg13g2_fill_1 FILLER_67_1392 ();
 sg13g2_fill_2 FILLER_67_1405 ();
 sg13g2_fill_1 FILLER_67_1411 ();
 sg13g2_fill_1 FILLER_67_1417 ();
 sg13g2_fill_2 FILLER_67_1430 ();
 sg13g2_fill_1 FILLER_67_1432 ();
 sg13g2_fill_2 FILLER_67_1454 ();
 sg13g2_fill_1 FILLER_67_1461 ();
 sg13g2_fill_2 FILLER_67_1480 ();
 sg13g2_decap_8 FILLER_67_1487 ();
 sg13g2_decap_4 FILLER_67_1494 ();
 sg13g2_fill_2 FILLER_67_1530 ();
 sg13g2_fill_1 FILLER_67_1552 ();
 sg13g2_fill_1 FILLER_67_1559 ();
 sg13g2_fill_2 FILLER_67_1578 ();
 sg13g2_fill_1 FILLER_67_1580 ();
 sg13g2_fill_2 FILLER_67_1587 ();
 sg13g2_fill_1 FILLER_67_1589 ();
 sg13g2_fill_2 FILLER_67_1595 ();
 sg13g2_fill_1 FILLER_67_1597 ();
 sg13g2_fill_2 FILLER_67_1617 ();
 sg13g2_fill_1 FILLER_67_1619 ();
 sg13g2_decap_4 FILLER_67_1625 ();
 sg13g2_fill_1 FILLER_67_1633 ();
 sg13g2_fill_2 FILLER_67_1639 ();
 sg13g2_fill_1 FILLER_67_1641 ();
 sg13g2_fill_1 FILLER_67_1647 ();
 sg13g2_fill_1 FILLER_67_1654 ();
 sg13g2_fill_2 FILLER_67_1660 ();
 sg13g2_fill_1 FILLER_67_1667 ();
 sg13g2_fill_2 FILLER_67_1673 ();
 sg13g2_fill_1 FILLER_67_1697 ();
 sg13g2_decap_4 FILLER_67_1702 ();
 sg13g2_fill_2 FILLER_67_1710 ();
 sg13g2_fill_1 FILLER_67_1712 ();
 sg13g2_fill_1 FILLER_67_1732 ();
 sg13g2_decap_8 FILLER_67_1738 ();
 sg13g2_fill_2 FILLER_67_1745 ();
 sg13g2_decap_4 FILLER_67_1755 ();
 sg13g2_fill_2 FILLER_67_1764 ();
 sg13g2_fill_1 FILLER_67_1766 ();
 sg13g2_fill_1 FILLER_67_1785 ();
 sg13g2_fill_1 FILLER_67_1795 ();
 sg13g2_fill_1 FILLER_67_1800 ();
 sg13g2_fill_2 FILLER_67_1805 ();
 sg13g2_decap_8 FILLER_67_1811 ();
 sg13g2_decap_4 FILLER_67_1822 ();
 sg13g2_fill_1 FILLER_67_1826 ();
 sg13g2_decap_4 FILLER_67_1831 ();
 sg13g2_fill_2 FILLER_67_1835 ();
 sg13g2_fill_1 FILLER_67_1841 ();
 sg13g2_decap_4 FILLER_67_1846 ();
 sg13g2_fill_1 FILLER_67_1850 ();
 sg13g2_fill_1 FILLER_67_1864 ();
 sg13g2_fill_1 FILLER_67_1871 ();
 sg13g2_fill_2 FILLER_67_1877 ();
 sg13g2_fill_1 FILLER_67_1879 ();
 sg13g2_fill_2 FILLER_67_1890 ();
 sg13g2_decap_4 FILLER_67_1897 ();
 sg13g2_decap_8 FILLER_67_1910 ();
 sg13g2_fill_2 FILLER_67_1917 ();
 sg13g2_fill_1 FILLER_67_1919 ();
 sg13g2_fill_1 FILLER_67_1925 ();
 sg13g2_fill_2 FILLER_67_1931 ();
 sg13g2_fill_1 FILLER_67_1937 ();
 sg13g2_fill_2 FILLER_67_1951 ();
 sg13g2_fill_2 FILLER_67_1978 ();
 sg13g2_fill_1 FILLER_67_1986 ();
 sg13g2_fill_1 FILLER_67_1993 ();
 sg13g2_decap_4 FILLER_67_2024 ();
 sg13g2_fill_1 FILLER_67_2028 ();
 sg13g2_decap_8 FILLER_67_2130 ();
 sg13g2_decap_4 FILLER_67_2137 ();
 sg13g2_decap_8 FILLER_67_2149 ();
 sg13g2_fill_2 FILLER_67_2156 ();
 sg13g2_fill_1 FILLER_67_2158 ();
 sg13g2_fill_2 FILLER_67_2169 ();
 sg13g2_decap_4 FILLER_67_2197 ();
 sg13g2_fill_2 FILLER_67_2241 ();
 sg13g2_fill_1 FILLER_67_2243 ();
 sg13g2_fill_1 FILLER_67_2294 ();
 sg13g2_fill_1 FILLER_67_2318 ();
 sg13g2_fill_2 FILLER_67_2323 ();
 sg13g2_decap_4 FILLER_67_2360 ();
 sg13g2_fill_2 FILLER_67_2364 ();
 sg13g2_fill_1 FILLER_67_2378 ();
 sg13g2_fill_2 FILLER_67_2410 ();
 sg13g2_fill_1 FILLER_67_2412 ();
 sg13g2_fill_1 FILLER_67_2448 ();
 sg13g2_fill_1 FILLER_67_2487 ();
 sg13g2_fill_1 FILLER_67_2532 ();
 sg13g2_fill_1 FILLER_67_2543 ();
 sg13g2_fill_1 FILLER_67_2555 ();
 sg13g2_fill_2 FILLER_67_2586 ();
 sg13g2_fill_2 FILLER_67_2592 ();
 sg13g2_fill_1 FILLER_67_2594 ();
 sg13g2_decap_4 FILLER_67_2605 ();
 sg13g2_fill_2 FILLER_67_2622 ();
 sg13g2_decap_8 FILLER_67_2643 ();
 sg13g2_decap_8 FILLER_67_2650 ();
 sg13g2_decap_8 FILLER_67_2657 ();
 sg13g2_decap_4 FILLER_67_2664 ();
 sg13g2_fill_2 FILLER_67_2668 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_fill_2 FILLER_68_14 ();
 sg13g2_fill_2 FILLER_68_20 ();
 sg13g2_fill_1 FILLER_68_22 ();
 sg13g2_decap_8 FILLER_68_27 ();
 sg13g2_fill_2 FILLER_68_34 ();
 sg13g2_fill_2 FILLER_68_71 ();
 sg13g2_fill_1 FILLER_68_73 ();
 sg13g2_fill_1 FILLER_68_115 ();
 sg13g2_decap_8 FILLER_68_130 ();
 sg13g2_decap_4 FILLER_68_137 ();
 sg13g2_fill_2 FILLER_68_141 ();
 sg13g2_decap_8 FILLER_68_159 ();
 sg13g2_decap_8 FILLER_68_166 ();
 sg13g2_decap_8 FILLER_68_173 ();
 sg13g2_decap_4 FILLER_68_180 ();
 sg13g2_fill_1 FILLER_68_189 ();
 sg13g2_fill_2 FILLER_68_204 ();
 sg13g2_fill_1 FILLER_68_226 ();
 sg13g2_fill_1 FILLER_68_232 ();
 sg13g2_fill_2 FILLER_68_238 ();
 sg13g2_fill_2 FILLER_68_245 ();
 sg13g2_fill_1 FILLER_68_247 ();
 sg13g2_fill_1 FILLER_68_253 ();
 sg13g2_fill_2 FILLER_68_260 ();
 sg13g2_fill_2 FILLER_68_278 ();
 sg13g2_fill_1 FILLER_68_280 ();
 sg13g2_fill_1 FILLER_68_292 ();
 sg13g2_fill_2 FILLER_68_298 ();
 sg13g2_fill_2 FILLER_68_305 ();
 sg13g2_fill_2 FILLER_68_312 ();
 sg13g2_decap_8 FILLER_68_318 ();
 sg13g2_decap_8 FILLER_68_325 ();
 sg13g2_decap_8 FILLER_68_332 ();
 sg13g2_decap_8 FILLER_68_339 ();
 sg13g2_decap_8 FILLER_68_354 ();
 sg13g2_decap_8 FILLER_68_361 ();
 sg13g2_fill_2 FILLER_68_372 ();
 sg13g2_fill_1 FILLER_68_379 ();
 sg13g2_fill_1 FILLER_68_390 ();
 sg13g2_fill_2 FILLER_68_456 ();
 sg13g2_fill_1 FILLER_68_463 ();
 sg13g2_fill_1 FILLER_68_493 ();
 sg13g2_fill_2 FILLER_68_530 ();
 sg13g2_fill_1 FILLER_68_536 ();
 sg13g2_decap_8 FILLER_68_541 ();
 sg13g2_decap_8 FILLER_68_548 ();
 sg13g2_decap_4 FILLER_68_555 ();
 sg13g2_fill_1 FILLER_68_590 ();
 sg13g2_decap_4 FILLER_68_600 ();
 sg13g2_fill_1 FILLER_68_604 ();
 sg13g2_decap_8 FILLER_68_623 ();
 sg13g2_fill_1 FILLER_68_644 ();
 sg13g2_fill_2 FILLER_68_685 ();
 sg13g2_fill_1 FILLER_68_687 ();
 sg13g2_fill_1 FILLER_68_700 ();
 sg13g2_fill_2 FILLER_68_706 ();
 sg13g2_decap_4 FILLER_68_721 ();
 sg13g2_fill_2 FILLER_68_725 ();
 sg13g2_decap_4 FILLER_68_750 ();
 sg13g2_fill_1 FILLER_68_754 ();
 sg13g2_fill_2 FILLER_68_761 ();
 sg13g2_fill_2 FILLER_68_799 ();
 sg13g2_fill_2 FILLER_68_833 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_fill_1 FILLER_68_866 ();
 sg13g2_fill_1 FILLER_68_899 ();
 sg13g2_fill_1 FILLER_68_905 ();
 sg13g2_fill_2 FILLER_68_932 ();
 sg13g2_decap_4 FILLER_68_944 ();
 sg13g2_fill_2 FILLER_68_968 ();
 sg13g2_fill_1 FILLER_68_970 ();
 sg13g2_decap_8 FILLER_68_985 ();
 sg13g2_decap_8 FILLER_68_992 ();
 sg13g2_fill_1 FILLER_68_999 ();
 sg13g2_fill_1 FILLER_68_1010 ();
 sg13g2_decap_8 FILLER_68_1017 ();
 sg13g2_decap_8 FILLER_68_1024 ();
 sg13g2_decap_8 FILLER_68_1031 ();
 sg13g2_decap_8 FILLER_68_1038 ();
 sg13g2_fill_1 FILLER_68_1045 ();
 sg13g2_fill_2 FILLER_68_1058 ();
 sg13g2_fill_1 FILLER_68_1060 ();
 sg13g2_decap_8 FILLER_68_1075 ();
 sg13g2_fill_2 FILLER_68_1082 ();
 sg13g2_fill_1 FILLER_68_1084 ();
 sg13g2_decap_8 FILLER_68_1095 ();
 sg13g2_fill_1 FILLER_68_1102 ();
 sg13g2_decap_4 FILLER_68_1107 ();
 sg13g2_fill_2 FILLER_68_1111 ();
 sg13g2_decap_8 FILLER_68_1117 ();
 sg13g2_decap_4 FILLER_68_1124 ();
 sg13g2_fill_2 FILLER_68_1128 ();
 sg13g2_decap_4 FILLER_68_1135 ();
 sg13g2_fill_2 FILLER_68_1159 ();
 sg13g2_fill_2 FILLER_68_1178 ();
 sg13g2_fill_2 FILLER_68_1206 ();
 sg13g2_fill_2 FILLER_68_1220 ();
 sg13g2_fill_1 FILLER_68_1222 ();
 sg13g2_fill_2 FILLER_68_1231 ();
 sg13g2_fill_1 FILLER_68_1305 ();
 sg13g2_fill_1 FILLER_68_1321 ();
 sg13g2_fill_1 FILLER_68_1327 ();
 sg13g2_fill_1 FILLER_68_1338 ();
 sg13g2_fill_2 FILLER_68_1344 ();
 sg13g2_fill_2 FILLER_68_1351 ();
 sg13g2_fill_1 FILLER_68_1365 ();
 sg13g2_fill_2 FILLER_68_1393 ();
 sg13g2_fill_1 FILLER_68_1395 ();
 sg13g2_fill_1 FILLER_68_1401 ();
 sg13g2_fill_2 FILLER_68_1428 ();
 sg13g2_fill_1 FILLER_68_1430 ();
 sg13g2_decap_8 FILLER_68_1452 ();
 sg13g2_fill_1 FILLER_68_1459 ();
 sg13g2_fill_2 FILLER_68_1504 ();
 sg13g2_fill_1 FILLER_68_1506 ();
 sg13g2_fill_2 FILLER_68_1511 ();
 sg13g2_fill_1 FILLER_68_1529 ();
 sg13g2_fill_1 FILLER_68_1544 ();
 sg13g2_decap_4 FILLER_68_1595 ();
 sg13g2_fill_1 FILLER_68_1607 ();
 sg13g2_decap_8 FILLER_68_1649 ();
 sg13g2_decap_8 FILLER_68_1656 ();
 sg13g2_decap_4 FILLER_68_1663 ();
 sg13g2_decap_8 FILLER_68_1672 ();
 sg13g2_decap_8 FILLER_68_1679 ();
 sg13g2_decap_4 FILLER_68_1695 ();
 sg13g2_decap_8 FILLER_68_1704 ();
 sg13g2_fill_1 FILLER_68_1711 ();
 sg13g2_fill_1 FILLER_68_1722 ();
 sg13g2_fill_1 FILLER_68_1729 ();
 sg13g2_fill_1 FILLER_68_1734 ();
 sg13g2_fill_1 FILLER_68_1739 ();
 sg13g2_decap_8 FILLER_68_1752 ();
 sg13g2_decap_8 FILLER_68_1759 ();
 sg13g2_decap_4 FILLER_68_1766 ();
 sg13g2_fill_1 FILLER_68_1770 ();
 sg13g2_fill_2 FILLER_68_1778 ();
 sg13g2_fill_1 FILLER_68_1794 ();
 sg13g2_decap_8 FILLER_68_1802 ();
 sg13g2_decap_8 FILLER_68_1809 ();
 sg13g2_decap_8 FILLER_68_1816 ();
 sg13g2_fill_2 FILLER_68_1823 ();
 sg13g2_fill_1 FILLER_68_1825 ();
 sg13g2_fill_2 FILLER_68_1834 ();
 sg13g2_fill_2 FILLER_68_1871 ();
 sg13g2_fill_1 FILLER_68_1873 ();
 sg13g2_decap_4 FILLER_68_1890 ();
 sg13g2_decap_4 FILLER_68_1899 ();
 sg13g2_fill_2 FILLER_68_1903 ();
 sg13g2_decap_8 FILLER_68_1910 ();
 sg13g2_fill_2 FILLER_68_1917 ();
 sg13g2_fill_1 FILLER_68_1923 ();
 sg13g2_fill_2 FILLER_68_1943 ();
 sg13g2_fill_1 FILLER_68_1945 ();
 sg13g2_fill_1 FILLER_68_1966 ();
 sg13g2_fill_2 FILLER_68_2015 ();
 sg13g2_fill_1 FILLER_68_2021 ();
 sg13g2_decap_4 FILLER_68_2026 ();
 sg13g2_fill_1 FILLER_68_2056 ();
 sg13g2_decap_8 FILLER_68_2073 ();
 sg13g2_fill_2 FILLER_68_2080 ();
 sg13g2_fill_1 FILLER_68_2082 ();
 sg13g2_decap_8 FILLER_68_2119 ();
 sg13g2_decap_4 FILLER_68_2126 ();
 sg13g2_fill_2 FILLER_68_2130 ();
 sg13g2_decap_8 FILLER_68_2153 ();
 sg13g2_decap_8 FILLER_68_2160 ();
 sg13g2_decap_4 FILLER_68_2167 ();
 sg13g2_fill_2 FILLER_68_2171 ();
 sg13g2_decap_8 FILLER_68_2235 ();
 sg13g2_decap_8 FILLER_68_2242 ();
 sg13g2_decap_8 FILLER_68_2249 ();
 sg13g2_decap_4 FILLER_68_2260 ();
 sg13g2_fill_1 FILLER_68_2264 ();
 sg13g2_decap_4 FILLER_68_2304 ();
 sg13g2_fill_2 FILLER_68_2308 ();
 sg13g2_decap_8 FILLER_68_2318 ();
 sg13g2_decap_4 FILLER_68_2325 ();
 sg13g2_fill_2 FILLER_68_2329 ();
 sg13g2_fill_2 FILLER_68_2369 ();
 sg13g2_fill_1 FILLER_68_2371 ();
 sg13g2_fill_1 FILLER_68_2414 ();
 sg13g2_fill_2 FILLER_68_2452 ();
 sg13g2_fill_1 FILLER_68_2459 ();
 sg13g2_fill_1 FILLER_68_2548 ();
 sg13g2_fill_1 FILLER_68_2557 ();
 sg13g2_fill_1 FILLER_68_2581 ();
 sg13g2_fill_2 FILLER_68_2587 ();
 sg13g2_fill_1 FILLER_68_2622 ();
 sg13g2_fill_2 FILLER_68_2637 ();
 sg13g2_fill_1 FILLER_68_2639 ();
 sg13g2_decap_4 FILLER_68_2666 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_4 FILLER_69_7 ();
 sg13g2_fill_2 FILLER_69_15 ();
 sg13g2_fill_2 FILLER_69_51 ();
 sg13g2_fill_1 FILLER_69_53 ();
 sg13g2_fill_1 FILLER_69_74 ();
 sg13g2_fill_1 FILLER_69_80 ();
 sg13g2_decap_4 FILLER_69_116 ();
 sg13g2_fill_2 FILLER_69_124 ();
 sg13g2_fill_1 FILLER_69_126 ();
 sg13g2_fill_2 FILLER_69_133 ();
 sg13g2_fill_1 FILLER_69_149 ();
 sg13g2_decap_8 FILLER_69_176 ();
 sg13g2_decap_8 FILLER_69_188 ();
 sg13g2_decap_4 FILLER_69_195 ();
 sg13g2_decap_8 FILLER_69_203 ();
 sg13g2_fill_1 FILLER_69_210 ();
 sg13g2_fill_1 FILLER_69_269 ();
 sg13g2_fill_1 FILLER_69_278 ();
 sg13g2_fill_1 FILLER_69_287 ();
 sg13g2_fill_2 FILLER_69_295 ();
 sg13g2_fill_2 FILLER_69_303 ();
 sg13g2_fill_2 FILLER_69_310 ();
 sg13g2_decap_8 FILLER_69_333 ();
 sg13g2_fill_2 FILLER_69_340 ();
 sg13g2_fill_1 FILLER_69_383 ();
 sg13g2_fill_1 FILLER_69_403 ();
 sg13g2_fill_2 FILLER_69_418 ();
 sg13g2_fill_1 FILLER_69_425 ();
 sg13g2_fill_2 FILLER_69_455 ();
 sg13g2_fill_2 FILLER_69_493 ();
 sg13g2_fill_1 FILLER_69_495 ();
 sg13g2_fill_1 FILLER_69_509 ();
 sg13g2_decap_8 FILLER_69_546 ();
 sg13g2_decap_4 FILLER_69_553 ();
 sg13g2_fill_2 FILLER_69_592 ();
 sg13g2_fill_1 FILLER_69_594 ();
 sg13g2_fill_2 FILLER_69_625 ();
 sg13g2_decap_4 FILLER_69_631 ();
 sg13g2_decap_8 FILLER_69_639 ();
 sg13g2_decap_8 FILLER_69_646 ();
 sg13g2_decap_8 FILLER_69_653 ();
 sg13g2_decap_8 FILLER_69_660 ();
 sg13g2_decap_8 FILLER_69_667 ();
 sg13g2_decap_8 FILLER_69_674 ();
 sg13g2_decap_8 FILLER_69_681 ();
 sg13g2_fill_2 FILLER_69_688 ();
 sg13g2_fill_1 FILLER_69_690 ();
 sg13g2_decap_4 FILLER_69_734 ();
 sg13g2_fill_1 FILLER_69_744 ();
 sg13g2_decap_4 FILLER_69_755 ();
 sg13g2_fill_1 FILLER_69_759 ();
 sg13g2_fill_1 FILLER_69_766 ();
 sg13g2_fill_1 FILLER_69_777 ();
 sg13g2_fill_1 FILLER_69_782 ();
 sg13g2_fill_1 FILLER_69_787 ();
 sg13g2_fill_1 FILLER_69_792 ();
 sg13g2_fill_1 FILLER_69_797 ();
 sg13g2_fill_2 FILLER_69_803 ();
 sg13g2_fill_1 FILLER_69_832 ();
 sg13g2_decap_8 FILLER_69_851 ();
 sg13g2_decap_4 FILLER_69_858 ();
 sg13g2_fill_2 FILLER_69_862 ();
 sg13g2_fill_1 FILLER_69_878 ();
 sg13g2_decap_8 FILLER_69_946 ();
 sg13g2_decap_8 FILLER_69_953 ();
 sg13g2_decap_8 FILLER_69_960 ();
 sg13g2_decap_4 FILLER_69_967 ();
 sg13g2_decap_8 FILLER_69_988 ();
 sg13g2_fill_1 FILLER_69_1005 ();
 sg13g2_decap_4 FILLER_69_1016 ();
 sg13g2_decap_8 FILLER_69_1056 ();
 sg13g2_decap_8 FILLER_69_1063 ();
 sg13g2_fill_2 FILLER_69_1070 ();
 sg13g2_decap_8 FILLER_69_1078 ();
 sg13g2_decap_8 FILLER_69_1085 ();
 sg13g2_decap_8 FILLER_69_1092 ();
 sg13g2_decap_8 FILLER_69_1099 ();
 sg13g2_decap_8 FILLER_69_1106 ();
 sg13g2_fill_1 FILLER_69_1113 ();
 sg13g2_decap_8 FILLER_69_1124 ();
 sg13g2_decap_8 FILLER_69_1131 ();
 sg13g2_fill_2 FILLER_69_1193 ();
 sg13g2_fill_2 FILLER_69_1247 ();
 sg13g2_fill_1 FILLER_69_1283 ();
 sg13g2_fill_1 FILLER_69_1288 ();
 sg13g2_fill_1 FILLER_69_1294 ();
 sg13g2_decap_4 FILLER_69_1305 ();
 sg13g2_decap_8 FILLER_69_1317 ();
 sg13g2_fill_1 FILLER_69_1329 ();
 sg13g2_fill_2 FILLER_69_1337 ();
 sg13g2_decap_4 FILLER_69_1354 ();
 sg13g2_decap_4 FILLER_69_1392 ();
 sg13g2_fill_2 FILLER_69_1396 ();
 sg13g2_decap_4 FILLER_69_1424 ();
 sg13g2_decap_8 FILLER_69_1433 ();
 sg13g2_decap_8 FILLER_69_1440 ();
 sg13g2_decap_8 FILLER_69_1447 ();
 sg13g2_fill_1 FILLER_69_1494 ();
 sg13g2_fill_1 FILLER_69_1526 ();
 sg13g2_fill_2 FILLER_69_1591 ();
 sg13g2_decap_8 FILLER_69_1634 ();
 sg13g2_decap_8 FILLER_69_1641 ();
 sg13g2_fill_2 FILLER_69_1648 ();
 sg13g2_decap_8 FILLER_69_1668 ();
 sg13g2_decap_8 FILLER_69_1675 ();
 sg13g2_decap_4 FILLER_69_1682 ();
 sg13g2_decap_8 FILLER_69_1690 ();
 sg13g2_fill_1 FILLER_69_1709 ();
 sg13g2_fill_2 FILLER_69_1719 ();
 sg13g2_fill_1 FILLER_69_1721 ();
 sg13g2_fill_1 FILLER_69_1727 ();
 sg13g2_decap_4 FILLER_69_1750 ();
 sg13g2_fill_1 FILLER_69_1754 ();
 sg13g2_fill_2 FILLER_69_1759 ();
 sg13g2_fill_1 FILLER_69_1765 ();
 sg13g2_fill_1 FILLER_69_1772 ();
 sg13g2_fill_2 FILLER_69_1800 ();
 sg13g2_fill_1 FILLER_69_1802 ();
 sg13g2_decap_8 FILLER_69_1807 ();
 sg13g2_decap_4 FILLER_69_1814 ();
 sg13g2_fill_1 FILLER_69_1818 ();
 sg13g2_fill_1 FILLER_69_1824 ();
 sg13g2_fill_2 FILLER_69_1830 ();
 sg13g2_fill_1 FILLER_69_1844 ();
 sg13g2_fill_1 FILLER_69_1864 ();
 sg13g2_fill_2 FILLER_69_1869 ();
 sg13g2_fill_2 FILLER_69_1874 ();
 sg13g2_fill_1 FILLER_69_1927 ();
 sg13g2_fill_1 FILLER_69_1933 ();
 sg13g2_fill_1 FILLER_69_1940 ();
 sg13g2_fill_1 FILLER_69_1956 ();
 sg13g2_fill_2 FILLER_69_1967 ();
 sg13g2_fill_1 FILLER_69_2000 ();
 sg13g2_fill_2 FILLER_69_2055 ();
 sg13g2_fill_2 FILLER_69_2071 ();
 sg13g2_fill_1 FILLER_69_2129 ();
 sg13g2_decap_8 FILLER_69_2155 ();
 sg13g2_fill_2 FILLER_69_2162 ();
 sg13g2_fill_2 FILLER_69_2174 ();
 sg13g2_fill_1 FILLER_69_2204 ();
 sg13g2_decap_4 FILLER_69_2259 ();
 sg13g2_decap_8 FILLER_69_2272 ();
 sg13g2_decap_4 FILLER_69_2279 ();
 sg13g2_fill_2 FILLER_69_2283 ();
 sg13g2_decap_4 FILLER_69_2288 ();
 sg13g2_fill_1 FILLER_69_2309 ();
 sg13g2_decap_4 FILLER_69_2323 ();
 sg13g2_fill_1 FILLER_69_2327 ();
 sg13g2_decap_8 FILLER_69_2333 ();
 sg13g2_decap_8 FILLER_69_2340 ();
 sg13g2_fill_2 FILLER_69_2357 ();
 sg13g2_decap_4 FILLER_69_2369 ();
 sg13g2_fill_2 FILLER_69_2373 ();
 sg13g2_fill_2 FILLER_69_2380 ();
 sg13g2_fill_2 FILLER_69_2390 ();
 sg13g2_fill_1 FILLER_69_2396 ();
 sg13g2_fill_1 FILLER_69_2401 ();
 sg13g2_fill_1 FILLER_69_2428 ();
 sg13g2_fill_1 FILLER_69_2433 ();
 sg13g2_fill_1 FILLER_69_2438 ();
 sg13g2_fill_2 FILLER_69_2449 ();
 sg13g2_fill_2 FILLER_69_2493 ();
 sg13g2_fill_2 FILLER_69_2505 ();
 sg13g2_fill_2 FILLER_69_2538 ();
 sg13g2_decap_8 FILLER_69_2580 ();
 sg13g2_fill_1 FILLER_69_2587 ();
 sg13g2_fill_2 FILLER_69_2621 ();
 sg13g2_fill_1 FILLER_69_2623 ();
 sg13g2_decap_8 FILLER_69_2660 ();
 sg13g2_fill_2 FILLER_69_2667 ();
 sg13g2_fill_1 FILLER_69_2669 ();
 sg13g2_decap_4 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_4 ();
 sg13g2_decap_4 FILLER_70_31 ();
 sg13g2_fill_1 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_51 ();
 sg13g2_fill_2 FILLER_70_58 ();
 sg13g2_fill_1 FILLER_70_60 ();
 sg13g2_fill_2 FILLER_70_84 ();
 sg13g2_fill_1 FILLER_70_86 ();
 sg13g2_decap_8 FILLER_70_108 ();
 sg13g2_decap_8 FILLER_70_115 ();
 sg13g2_decap_8 FILLER_70_122 ();
 sg13g2_decap_8 FILLER_70_129 ();
 sg13g2_decap_8 FILLER_70_136 ();
 sg13g2_decap_8 FILLER_70_185 ();
 sg13g2_decap_8 FILLER_70_192 ();
 sg13g2_fill_1 FILLER_70_203 ();
 sg13g2_fill_1 FILLER_70_208 ();
 sg13g2_fill_1 FILLER_70_213 ();
 sg13g2_fill_1 FILLER_70_233 ();
 sg13g2_fill_2 FILLER_70_269 ();
 sg13g2_fill_1 FILLER_70_271 ();
 sg13g2_fill_2 FILLER_70_310 ();
 sg13g2_decap_8 FILLER_70_333 ();
 sg13g2_decap_8 FILLER_70_340 ();
 sg13g2_decap_8 FILLER_70_347 ();
 sg13g2_fill_1 FILLER_70_354 ();
 sg13g2_fill_1 FILLER_70_407 ();
 sg13g2_fill_2 FILLER_70_412 ();
 sg13g2_fill_1 FILLER_70_440 ();
 sg13g2_fill_2 FILLER_70_467 ();
 sg13g2_fill_1 FILLER_70_469 ();
 sg13g2_fill_1 FILLER_70_480 ();
 sg13g2_fill_2 FILLER_70_512 ();
 sg13g2_fill_1 FILLER_70_514 ();
 sg13g2_fill_1 FILLER_70_524 ();
 sg13g2_decap_8 FILLER_70_556 ();
 sg13g2_fill_1 FILLER_70_563 ();
 sg13g2_fill_1 FILLER_70_592 ();
 sg13g2_fill_1 FILLER_70_598 ();
 sg13g2_fill_2 FILLER_70_614 ();
 sg13g2_decap_8 FILLER_70_622 ();
 sg13g2_fill_1 FILLER_70_629 ();
 sg13g2_fill_1 FILLER_70_653 ();
 sg13g2_fill_2 FILLER_70_673 ();
 sg13g2_fill_1 FILLER_70_675 ();
 sg13g2_decap_8 FILLER_70_686 ();
 sg13g2_decap_4 FILLER_70_693 ();
 sg13g2_fill_2 FILLER_70_697 ();
 sg13g2_fill_1 FILLER_70_725 ();
 sg13g2_fill_2 FILLER_70_742 ();
 sg13g2_decap_4 FILLER_70_770 ();
 sg13g2_decap_8 FILLER_70_779 ();
 sg13g2_decap_4 FILLER_70_786 ();
 sg13g2_fill_1 FILLER_70_795 ();
 sg13g2_fill_2 FILLER_70_801 ();
 sg13g2_decap_8 FILLER_70_807 ();
 sg13g2_decap_8 FILLER_70_819 ();
 sg13g2_decap_8 FILLER_70_826 ();
 sg13g2_decap_8 FILLER_70_833 ();
 sg13g2_decap_8 FILLER_70_840 ();
 sg13g2_decap_8 FILLER_70_847 ();
 sg13g2_decap_8 FILLER_70_854 ();
 sg13g2_fill_2 FILLER_70_861 ();
 sg13g2_fill_1 FILLER_70_863 ();
 sg13g2_decap_4 FILLER_70_894 ();
 sg13g2_decap_4 FILLER_70_901 ();
 sg13g2_fill_2 FILLER_70_921 ();
 sg13g2_fill_1 FILLER_70_923 ();
 sg13g2_decap_8 FILLER_70_935 ();
 sg13g2_decap_8 FILLER_70_942 ();
 sg13g2_decap_4 FILLER_70_949 ();
 sg13g2_fill_1 FILLER_70_963 ();
 sg13g2_fill_1 FILLER_70_970 ();
 sg13g2_fill_2 FILLER_70_981 ();
 sg13g2_fill_2 FILLER_70_987 ();
 sg13g2_fill_2 FILLER_70_995 ();
 sg13g2_fill_1 FILLER_70_997 ();
 sg13g2_fill_2 FILLER_70_1054 ();
 sg13g2_fill_1 FILLER_70_1056 ();
 sg13g2_fill_2 FILLER_70_1067 ();
 sg13g2_fill_2 FILLER_70_1075 ();
 sg13g2_fill_1 FILLER_70_1107 ();
 sg13g2_fill_2 FILLER_70_1118 ();
 sg13g2_fill_1 FILLER_70_1149 ();
 sg13g2_fill_2 FILLER_70_1155 ();
 sg13g2_fill_2 FILLER_70_1171 ();
 sg13g2_decap_4 FILLER_70_1183 ();
 sg13g2_fill_1 FILLER_70_1187 ();
 sg13g2_fill_2 FILLER_70_1236 ();
 sg13g2_decap_8 FILLER_70_1253 ();
 sg13g2_decap_8 FILLER_70_1260 ();
 sg13g2_decap_8 FILLER_70_1267 ();
 sg13g2_decap_8 FILLER_70_1274 ();
 sg13g2_decap_8 FILLER_70_1281 ();
 sg13g2_decap_4 FILLER_70_1288 ();
 sg13g2_decap_4 FILLER_70_1319 ();
 sg13g2_fill_1 FILLER_70_1323 ();
 sg13g2_fill_2 FILLER_70_1331 ();
 sg13g2_decap_4 FILLER_70_1340 ();
 sg13g2_decap_4 FILLER_70_1349 ();
 sg13g2_fill_2 FILLER_70_1376 ();
 sg13g2_fill_1 FILLER_70_1378 ();
 sg13g2_fill_2 FILLER_70_1392 ();
 sg13g2_fill_1 FILLER_70_1394 ();
 sg13g2_decap_8 FILLER_70_1403 ();
 sg13g2_decap_4 FILLER_70_1410 ();
 sg13g2_fill_1 FILLER_70_1414 ();
 sg13g2_fill_2 FILLER_70_1428 ();
 sg13g2_fill_1 FILLER_70_1430 ();
 sg13g2_decap_8 FILLER_70_1435 ();
 sg13g2_decap_4 FILLER_70_1442 ();
 sg13g2_fill_1 FILLER_70_1446 ();
 sg13g2_decap_4 FILLER_70_1461 ();
 sg13g2_fill_1 FILLER_70_1465 ();
 sg13g2_fill_2 FILLER_70_1471 ();
 sg13g2_fill_1 FILLER_70_1473 ();
 sg13g2_decap_8 FILLER_70_1478 ();
 sg13g2_decap_8 FILLER_70_1485 ();
 sg13g2_decap_8 FILLER_70_1492 ();
 sg13g2_decap_4 FILLER_70_1499 ();
 sg13g2_fill_1 FILLER_70_1541 ();
 sg13g2_fill_2 FILLER_70_1582 ();
 sg13g2_fill_1 FILLER_70_1584 ();
 sg13g2_fill_2 FILLER_70_1593 ();
 sg13g2_fill_1 FILLER_70_1595 ();
 sg13g2_decap_4 FILLER_70_1636 ();
 sg13g2_fill_2 FILLER_70_1658 ();
 sg13g2_fill_1 FILLER_70_1660 ();
 sg13g2_fill_2 FILLER_70_1666 ();
 sg13g2_fill_1 FILLER_70_1668 ();
 sg13g2_decap_8 FILLER_70_1674 ();
 sg13g2_decap_4 FILLER_70_1681 ();
 sg13g2_fill_1 FILLER_70_1685 ();
 sg13g2_decap_8 FILLER_70_1690 ();
 sg13g2_decap_4 FILLER_70_1697 ();
 sg13g2_fill_2 FILLER_70_1701 ();
 sg13g2_decap_4 FILLER_70_1707 ();
 sg13g2_decap_8 FILLER_70_1730 ();
 sg13g2_decap_4 FILLER_70_1742 ();
 sg13g2_fill_2 FILLER_70_1746 ();
 sg13g2_fill_1 FILLER_70_1769 ();
 sg13g2_fill_2 FILLER_70_1787 ();
 sg13g2_fill_1 FILLER_70_1795 ();
 sg13g2_fill_2 FILLER_70_1804 ();
 sg13g2_decap_8 FILLER_70_1811 ();
 sg13g2_decap_8 FILLER_70_1818 ();
 sg13g2_fill_2 FILLER_70_1825 ();
 sg13g2_fill_1 FILLER_70_1850 ();
 sg13g2_fill_2 FILLER_70_1871 ();
 sg13g2_decap_8 FILLER_70_1877 ();
 sg13g2_fill_1 FILLER_70_1884 ();
 sg13g2_decap_4 FILLER_70_1889 ();
 sg13g2_fill_1 FILLER_70_1906 ();
 sg13g2_fill_2 FILLER_70_1912 ();
 sg13g2_decap_8 FILLER_70_1917 ();
 sg13g2_decap_8 FILLER_70_1924 ();
 sg13g2_fill_1 FILLER_70_1931 ();
 sg13g2_fill_2 FILLER_70_1952 ();
 sg13g2_fill_2 FILLER_70_1959 ();
 sg13g2_fill_1 FILLER_70_1961 ();
 sg13g2_fill_2 FILLER_70_1967 ();
 sg13g2_fill_1 FILLER_70_1969 ();
 sg13g2_fill_1 FILLER_70_1978 ();
 sg13g2_fill_2 FILLER_70_2006 ();
 sg13g2_fill_1 FILLER_70_2008 ();
 sg13g2_fill_1 FILLER_70_2014 ();
 sg13g2_fill_2 FILLER_70_2051 ();
 sg13g2_decap_4 FILLER_70_2155 ();
 sg13g2_fill_2 FILLER_70_2159 ();
 sg13g2_fill_1 FILLER_70_2171 ();
 sg13g2_fill_1 FILLER_70_2217 ();
 sg13g2_decap_8 FILLER_70_2252 ();
 sg13g2_fill_1 FILLER_70_2259 ();
 sg13g2_fill_1 FILLER_70_2270 ();
 sg13g2_fill_1 FILLER_70_2284 ();
 sg13g2_fill_1 FILLER_70_2354 ();
 sg13g2_decap_8 FILLER_70_2387 ();
 sg13g2_decap_8 FILLER_70_2394 ();
 sg13g2_decap_8 FILLER_70_2401 ();
 sg13g2_decap_4 FILLER_70_2433 ();
 sg13g2_decap_8 FILLER_70_2467 ();
 sg13g2_fill_1 FILLER_70_2474 ();
 sg13g2_fill_1 FILLER_70_2486 ();
 sg13g2_fill_1 FILLER_70_2499 ();
 sg13g2_fill_1 FILLER_70_2526 ();
 sg13g2_fill_2 FILLER_70_2532 ();
 sg13g2_fill_2 FILLER_70_2548 ();
 sg13g2_fill_1 FILLER_70_2565 ();
 sg13g2_fill_2 FILLER_70_2592 ();
 sg13g2_fill_2 FILLER_70_2604 ();
 sg13g2_fill_1 FILLER_70_2606 ();
 sg13g2_decap_8 FILLER_70_2659 ();
 sg13g2_decap_4 FILLER_70_2666 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_42 ();
 sg13g2_fill_2 FILLER_71_69 ();
 sg13g2_decap_8 FILLER_71_110 ();
 sg13g2_decap_4 FILLER_71_117 ();
 sg13g2_fill_1 FILLER_71_121 ();
 sg13g2_fill_2 FILLER_71_179 ();
 sg13g2_fill_1 FILLER_71_216 ();
 sg13g2_fill_2 FILLER_71_221 ();
 sg13g2_fill_1 FILLER_71_228 ();
 sg13g2_fill_1 FILLER_71_235 ();
 sg13g2_fill_1 FILLER_71_240 ();
 sg13g2_decap_4 FILLER_71_272 ();
 sg13g2_fill_1 FILLER_71_276 ();
 sg13g2_fill_1 FILLER_71_282 ();
 sg13g2_decap_8 FILLER_71_327 ();
 sg13g2_decap_8 FILLER_71_334 ();
 sg13g2_decap_8 FILLER_71_341 ();
 sg13g2_fill_1 FILLER_71_348 ();
 sg13g2_fill_2 FILLER_71_359 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_fill_2 FILLER_71_415 ();
 sg13g2_fill_1 FILLER_71_417 ();
 sg13g2_fill_1 FILLER_71_422 ();
 sg13g2_decap_8 FILLER_71_428 ();
 sg13g2_fill_1 FILLER_71_435 ();
 sg13g2_decap_8 FILLER_71_440 ();
 sg13g2_fill_1 FILLER_71_447 ();
 sg13g2_decap_8 FILLER_71_452 ();
 sg13g2_decap_4 FILLER_71_459 ();
 sg13g2_decap_8 FILLER_71_468 ();
 sg13g2_decap_4 FILLER_71_475 ();
 sg13g2_fill_1 FILLER_71_479 ();
 sg13g2_decap_8 FILLER_71_490 ();
 sg13g2_decap_4 FILLER_71_497 ();
 sg13g2_fill_2 FILLER_71_505 ();
 sg13g2_fill_2 FILLER_71_511 ();
 sg13g2_fill_1 FILLER_71_513 ();
 sg13g2_decap_4 FILLER_71_524 ();
 sg13g2_fill_1 FILLER_71_528 ();
 sg13g2_fill_1 FILLER_71_544 ();
 sg13g2_decap_8 FILLER_71_550 ();
 sg13g2_decap_8 FILLER_71_557 ();
 sg13g2_fill_2 FILLER_71_564 ();
 sg13g2_decap_8 FILLER_71_570 ();
 sg13g2_fill_1 FILLER_71_577 ();
 sg13g2_fill_2 FILLER_71_582 ();
 sg13g2_fill_1 FILLER_71_584 ();
 sg13g2_fill_1 FILLER_71_594 ();
 sg13g2_fill_2 FILLER_71_621 ();
 sg13g2_fill_2 FILLER_71_689 ();
 sg13g2_fill_1 FILLER_71_691 ();
 sg13g2_fill_1 FILLER_71_753 ();
 sg13g2_fill_2 FILLER_71_758 ();
 sg13g2_fill_1 FILLER_71_760 ();
 sg13g2_fill_2 FILLER_71_780 ();
 sg13g2_fill_1 FILLER_71_786 ();
 sg13g2_decap_8 FILLER_71_792 ();
 sg13g2_fill_2 FILLER_71_799 ();
 sg13g2_decap_4 FILLER_71_805 ();
 sg13g2_decap_8 FILLER_71_813 ();
 sg13g2_decap_8 FILLER_71_820 ();
 sg13g2_fill_2 FILLER_71_827 ();
 sg13g2_decap_8 FILLER_71_834 ();
 sg13g2_decap_8 FILLER_71_841 ();
 sg13g2_decap_8 FILLER_71_848 ();
 sg13g2_decap_8 FILLER_71_855 ();
 sg13g2_decap_8 FILLER_71_862 ();
 sg13g2_decap_8 FILLER_71_873 ();
 sg13g2_decap_8 FILLER_71_880 ();
 sg13g2_fill_2 FILLER_71_895 ();
 sg13g2_fill_1 FILLER_71_897 ();
 sg13g2_fill_1 FILLER_71_904 ();
 sg13g2_fill_2 FILLER_71_911 ();
 sg13g2_fill_1 FILLER_71_913 ();
 sg13g2_fill_1 FILLER_71_948 ();
 sg13g2_fill_1 FILLER_71_1023 ();
 sg13g2_decap_8 FILLER_71_1052 ();
 sg13g2_fill_2 FILLER_71_1059 ();
 sg13g2_decap_8 FILLER_71_1148 ();
 sg13g2_decap_8 FILLER_71_1155 ();
 sg13g2_fill_2 FILLER_71_1166 ();
 sg13g2_fill_1 FILLER_71_1168 ();
 sg13g2_decap_4 FILLER_71_1250 ();
 sg13g2_fill_2 FILLER_71_1254 ();
 sg13g2_decap_8 FILLER_71_1266 ();
 sg13g2_decap_4 FILLER_71_1273 ();
 sg13g2_fill_1 FILLER_71_1277 ();
 sg13g2_decap_8 FILLER_71_1286 ();
 sg13g2_decap_8 FILLER_71_1293 ();
 sg13g2_fill_2 FILLER_71_1300 ();
 sg13g2_decap_8 FILLER_71_1307 ();
 sg13g2_decap_8 FILLER_71_1314 ();
 sg13g2_decap_8 FILLER_71_1321 ();
 sg13g2_decap_8 FILLER_71_1346 ();
 sg13g2_decap_4 FILLER_71_1353 ();
 sg13g2_fill_1 FILLER_71_1357 ();
 sg13g2_decap_8 FILLER_71_1363 ();
 sg13g2_decap_8 FILLER_71_1374 ();
 sg13g2_decap_4 FILLER_71_1381 ();
 sg13g2_fill_1 FILLER_71_1385 ();
 sg13g2_decap_8 FILLER_71_1389 ();
 sg13g2_decap_8 FILLER_71_1396 ();
 sg13g2_decap_4 FILLER_71_1403 ();
 sg13g2_fill_1 FILLER_71_1417 ();
 sg13g2_fill_1 FILLER_71_1444 ();
 sg13g2_fill_1 FILLER_71_1449 ();
 sg13g2_fill_1 FILLER_71_1460 ();
 sg13g2_decap_8 FILLER_71_1491 ();
 sg13g2_decap_4 FILLER_71_1498 ();
 sg13g2_fill_2 FILLER_71_1502 ();
 sg13g2_fill_2 FILLER_71_1523 ();
 sg13g2_fill_1 FILLER_71_1540 ();
 sg13g2_fill_2 FILLER_71_1550 ();
 sg13g2_fill_1 FILLER_71_1562 ();
 sg13g2_decap_4 FILLER_71_1607 ();
 sg13g2_fill_2 FILLER_71_1611 ();
 sg13g2_fill_2 FILLER_71_1623 ();
 sg13g2_decap_8 FILLER_71_1630 ();
 sg13g2_decap_8 FILLER_71_1637 ();
 sg13g2_decap_4 FILLER_71_1644 ();
 sg13g2_fill_1 FILLER_71_1648 ();
 sg13g2_fill_2 FILLER_71_1664 ();
 sg13g2_fill_1 FILLER_71_1666 ();
 sg13g2_decap_8 FILLER_71_1675 ();
 sg13g2_decap_8 FILLER_71_1682 ();
 sg13g2_decap_8 FILLER_71_1689 ();
 sg13g2_fill_2 FILLER_71_1696 ();
 sg13g2_fill_2 FILLER_71_1707 ();
 sg13g2_fill_1 FILLER_71_1709 ();
 sg13g2_fill_1 FILLER_71_1720 ();
 sg13g2_fill_1 FILLER_71_1746 ();
 sg13g2_fill_1 FILLER_71_1752 ();
 sg13g2_fill_1 FILLER_71_1763 ();
 sg13g2_fill_2 FILLER_71_1768 ();
 sg13g2_decap_8 FILLER_71_1813 ();
 sg13g2_fill_1 FILLER_71_1825 ();
 sg13g2_fill_1 FILLER_71_1831 ();
 sg13g2_fill_1 FILLER_71_1837 ();
 sg13g2_fill_1 FILLER_71_1843 ();
 sg13g2_fill_1 FILLER_71_1848 ();
 sg13g2_fill_1 FILLER_71_1854 ();
 sg13g2_fill_1 FILLER_71_1860 ();
 sg13g2_fill_1 FILLER_71_1865 ();
 sg13g2_fill_1 FILLER_71_1883 ();
 sg13g2_fill_1 FILLER_71_1890 ();
 sg13g2_decap_4 FILLER_71_1896 ();
 sg13g2_decap_8 FILLER_71_1909 ();
 sg13g2_decap_8 FILLER_71_1916 ();
 sg13g2_decap_8 FILLER_71_1923 ();
 sg13g2_fill_1 FILLER_71_1930 ();
 sg13g2_fill_2 FILLER_71_1952 ();
 sg13g2_fill_2 FILLER_71_1972 ();
 sg13g2_fill_1 FILLER_71_1974 ();
 sg13g2_fill_1 FILLER_71_1996 ();
 sg13g2_fill_2 FILLER_71_2001 ();
 sg13g2_fill_2 FILLER_71_2007 ();
 sg13g2_decap_4 FILLER_71_2019 ();
 sg13g2_fill_1 FILLER_71_2048 ();
 sg13g2_fill_2 FILLER_71_2075 ();
 sg13g2_fill_1 FILLER_71_2077 ();
 sg13g2_fill_2 FILLER_71_2134 ();
 sg13g2_fill_1 FILLER_71_2162 ();
 sg13g2_fill_1 FILLER_71_2167 ();
 sg13g2_decap_8 FILLER_71_2194 ();
 sg13g2_fill_1 FILLER_71_2220 ();
 sg13g2_decap_8 FILLER_71_2247 ();
 sg13g2_fill_2 FILLER_71_2254 ();
 sg13g2_decap_8 FILLER_71_2296 ();
 sg13g2_decap_4 FILLER_71_2303 ();
 sg13g2_fill_1 FILLER_71_2307 ();
 sg13g2_fill_1 FILLER_71_2324 ();
 sg13g2_fill_1 FILLER_71_2334 ();
 sg13g2_fill_1 FILLER_71_2339 ();
 sg13g2_fill_2 FILLER_71_2345 ();
 sg13g2_fill_1 FILLER_71_2347 ();
 sg13g2_fill_2 FILLER_71_2359 ();
 sg13g2_fill_1 FILLER_71_2361 ();
 sg13g2_fill_1 FILLER_71_2388 ();
 sg13g2_decap_8 FILLER_71_2398 ();
 sg13g2_fill_1 FILLER_71_2405 ();
 sg13g2_decap_8 FILLER_71_2410 ();
 sg13g2_decap_8 FILLER_71_2417 ();
 sg13g2_decap_8 FILLER_71_2424 ();
 sg13g2_fill_1 FILLER_71_2431 ();
 sg13g2_decap_8 FILLER_71_2436 ();
 sg13g2_decap_8 FILLER_71_2443 ();
 sg13g2_fill_2 FILLER_71_2450 ();
 sg13g2_fill_1 FILLER_71_2452 ();
 sg13g2_decap_4 FILLER_71_2458 ();
 sg13g2_fill_1 FILLER_71_2462 ();
 sg13g2_fill_2 FILLER_71_2482 ();
 sg13g2_fill_1 FILLER_71_2484 ();
 sg13g2_fill_2 FILLER_71_2513 ();
 sg13g2_fill_2 FILLER_71_2520 ();
 sg13g2_fill_1 FILLER_71_2522 ();
 sg13g2_fill_1 FILLER_71_2549 ();
 sg13g2_fill_1 FILLER_71_2560 ();
 sg13g2_fill_1 FILLER_71_2587 ();
 sg13g2_fill_1 FILLER_71_2592 ();
 sg13g2_fill_2 FILLER_71_2623 ();
 sg13g2_fill_1 FILLER_71_2625 ();
 sg13g2_decap_4 FILLER_71_2636 ();
 sg13g2_fill_1 FILLER_71_2640 ();
 sg13g2_decap_8 FILLER_71_2649 ();
 sg13g2_decap_8 FILLER_71_2656 ();
 sg13g2_decap_8 FILLER_71_2663 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_4 FILLER_72_7 ();
 sg13g2_fill_1 FILLER_72_11 ();
 sg13g2_decap_8 FILLER_72_16 ();
 sg13g2_decap_8 FILLER_72_23 ();
 sg13g2_decap_8 FILLER_72_30 ();
 sg13g2_decap_4 FILLER_72_37 ();
 sg13g2_fill_2 FILLER_72_71 ();
 sg13g2_fill_1 FILLER_72_73 ();
 sg13g2_fill_2 FILLER_72_79 ();
 sg13g2_fill_1 FILLER_72_81 ();
 sg13g2_fill_1 FILLER_72_103 ();
 sg13g2_fill_2 FILLER_72_109 ();
 sg13g2_fill_1 FILLER_72_111 ();
 sg13g2_decap_8 FILLER_72_137 ();
 sg13g2_fill_2 FILLER_72_144 ();
 sg13g2_fill_1 FILLER_72_146 ();
 sg13g2_fill_1 FILLER_72_213 ();
 sg13g2_decap_4 FILLER_72_221 ();
 sg13g2_decap_4 FILLER_72_238 ();
 sg13g2_fill_1 FILLER_72_242 ();
 sg13g2_fill_1 FILLER_72_249 ();
 sg13g2_fill_2 FILLER_72_265 ();
 sg13g2_fill_2 FILLER_72_280 ();
 sg13g2_decap_4 FILLER_72_288 ();
 sg13g2_fill_2 FILLER_72_298 ();
 sg13g2_decap_4 FILLER_72_306 ();
 sg13g2_decap_8 FILLER_72_315 ();
 sg13g2_decap_4 FILLER_72_322 ();
 sg13g2_fill_1 FILLER_72_362 ();
 sg13g2_fill_2 FILLER_72_410 ();
 sg13g2_decap_8 FILLER_72_421 ();
 sg13g2_fill_2 FILLER_72_428 ();
 sg13g2_fill_1 FILLER_72_430 ();
 sg13g2_fill_1 FILLER_72_470 ();
 sg13g2_decap_4 FILLER_72_514 ();
 sg13g2_decap_8 FILLER_72_522 ();
 sg13g2_fill_2 FILLER_72_529 ();
 sg13g2_fill_1 FILLER_72_531 ();
 sg13g2_decap_8 FILLER_72_541 ();
 sg13g2_decap_8 FILLER_72_548 ();
 sg13g2_decap_8 FILLER_72_555 ();
 sg13g2_fill_2 FILLER_72_562 ();
 sg13g2_fill_1 FILLER_72_568 ();
 sg13g2_fill_1 FILLER_72_574 ();
 sg13g2_fill_1 FILLER_72_580 ();
 sg13g2_fill_2 FILLER_72_592 ();
 sg13g2_fill_1 FILLER_72_637 ();
 sg13g2_decap_4 FILLER_72_664 ();
 sg13g2_fill_1 FILLER_72_668 ();
 sg13g2_fill_2 FILLER_72_678 ();
 sg13g2_fill_1 FILLER_72_680 ();
 sg13g2_decap_8 FILLER_72_687 ();
 sg13g2_fill_2 FILLER_72_694 ();
 sg13g2_fill_2 FILLER_72_704 ();
 sg13g2_fill_1 FILLER_72_706 ();
 sg13g2_decap_4 FILLER_72_711 ();
 sg13g2_fill_2 FILLER_72_715 ();
 sg13g2_fill_1 FILLER_72_725 ();
 sg13g2_fill_2 FILLER_72_730 ();
 sg13g2_fill_2 FILLER_72_736 ();
 sg13g2_fill_2 FILLER_72_744 ();
 sg13g2_decap_8 FILLER_72_750 ();
 sg13g2_fill_1 FILLER_72_851 ();
 sg13g2_decap_4 FILLER_72_903 ();
 sg13g2_fill_1 FILLER_72_907 ();
 sg13g2_fill_1 FILLER_72_938 ();
 sg13g2_fill_1 FILLER_72_975 ();
 sg13g2_fill_1 FILLER_72_982 ();
 sg13g2_fill_2 FILLER_72_1009 ();
 sg13g2_fill_1 FILLER_72_1011 ();
 sg13g2_decap_8 FILLER_72_1017 ();
 sg13g2_fill_2 FILLER_72_1024 ();
 sg13g2_fill_1 FILLER_72_1026 ();
 sg13g2_decap_8 FILLER_72_1051 ();
 sg13g2_decap_4 FILLER_72_1058 ();
 sg13g2_fill_1 FILLER_72_1062 ();
 sg13g2_fill_1 FILLER_72_1108 ();
 sg13g2_decap_8 FILLER_72_1139 ();
 sg13g2_fill_2 FILLER_72_1146 ();
 sg13g2_decap_8 FILLER_72_1184 ();
 sg13g2_fill_2 FILLER_72_1191 ();
 sg13g2_fill_1 FILLER_72_1193 ();
 sg13g2_fill_2 FILLER_72_1228 ();
 sg13g2_decap_8 FILLER_72_1240 ();
 sg13g2_fill_2 FILLER_72_1247 ();
 sg13g2_fill_1 FILLER_72_1249 ();
 sg13g2_fill_2 FILLER_72_1286 ();
 sg13g2_decap_8 FILLER_72_1317 ();
 sg13g2_decap_8 FILLER_72_1324 ();
 sg13g2_decap_4 FILLER_72_1357 ();
 sg13g2_fill_2 FILLER_72_1361 ();
 sg13g2_decap_8 FILLER_72_1389 ();
 sg13g2_decap_8 FILLER_72_1396 ();
 sg13g2_fill_1 FILLER_72_1403 ();
 sg13g2_fill_1 FILLER_72_1447 ();
 sg13g2_decap_8 FILLER_72_1486 ();
 sg13g2_fill_2 FILLER_72_1493 ();
 sg13g2_fill_1 FILLER_72_1495 ();
 sg13g2_fill_1 FILLER_72_1533 ();
 sg13g2_fill_2 FILLER_72_1542 ();
 sg13g2_fill_1 FILLER_72_1552 ();
 sg13g2_fill_2 FILLER_72_1562 ();
 sg13g2_fill_2 FILLER_72_1588 ();
 sg13g2_fill_1 FILLER_72_1590 ();
 sg13g2_fill_1 FILLER_72_1617 ();
 sg13g2_decap_4 FILLER_72_1622 ();
 sg13g2_fill_2 FILLER_72_1630 ();
 sg13g2_fill_2 FILLER_72_1640 ();
 sg13g2_fill_1 FILLER_72_1642 ();
 sg13g2_decap_4 FILLER_72_1656 ();
 sg13g2_fill_2 FILLER_72_1660 ();
 sg13g2_fill_2 FILLER_72_1667 ();
 sg13g2_decap_8 FILLER_72_1673 ();
 sg13g2_decap_8 FILLER_72_1680 ();
 sg13g2_fill_1 FILLER_72_1687 ();
 sg13g2_fill_2 FILLER_72_1692 ();
 sg13g2_fill_1 FILLER_72_1698 ();
 sg13g2_fill_1 FILLER_72_1704 ();
 sg13g2_decap_4 FILLER_72_1710 ();
 sg13g2_fill_2 FILLER_72_1722 ();
 sg13g2_fill_2 FILLER_72_1730 ();
 sg13g2_fill_1 FILLER_72_1732 ();
 sg13g2_fill_1 FILLER_72_1763 ();
 sg13g2_fill_2 FILLER_72_1775 ();
 sg13g2_fill_2 FILLER_72_1791 ();
 sg13g2_fill_2 FILLER_72_1828 ();
 sg13g2_fill_1 FILLER_72_1836 ();
 sg13g2_fill_2 FILLER_72_1841 ();
 sg13g2_fill_1 FILLER_72_1849 ();
 sg13g2_fill_1 FILLER_72_1858 ();
 sg13g2_fill_1 FILLER_72_1863 ();
 sg13g2_fill_1 FILLER_72_1873 ();
 sg13g2_fill_1 FILLER_72_1878 ();
 sg13g2_fill_1 FILLER_72_1884 ();
 sg13g2_fill_1 FILLER_72_1895 ();
 sg13g2_fill_1 FILLER_72_1901 ();
 sg13g2_fill_2 FILLER_72_1907 ();
 sg13g2_fill_2 FILLER_72_1914 ();
 sg13g2_fill_2 FILLER_72_1921 ();
 sg13g2_fill_2 FILLER_72_1938 ();
 sg13g2_fill_1 FILLER_72_1940 ();
 sg13g2_fill_1 FILLER_72_1952 ();
 sg13g2_fill_1 FILLER_72_1988 ();
 sg13g2_decap_8 FILLER_72_1994 ();
 sg13g2_decap_8 FILLER_72_2001 ();
 sg13g2_fill_2 FILLER_72_2016 ();
 sg13g2_fill_1 FILLER_72_2044 ();
 sg13g2_fill_1 FILLER_72_2055 ();
 sg13g2_fill_1 FILLER_72_2082 ();
 sg13g2_fill_1 FILLER_72_2087 ();
 sg13g2_fill_2 FILLER_72_2105 ();
 sg13g2_fill_2 FILLER_72_2166 ();
 sg13g2_fill_1 FILLER_72_2220 ();
 sg13g2_fill_1 FILLER_72_2231 ();
 sg13g2_fill_2 FILLER_72_2309 ();
 sg13g2_fill_2 FILLER_72_2319 ();
 sg13g2_fill_1 FILLER_72_2358 ();
 sg13g2_fill_1 FILLER_72_2382 ();
 sg13g2_fill_1 FILLER_72_2388 ();
 sg13g2_fill_2 FILLER_72_2415 ();
 sg13g2_fill_1 FILLER_72_2423 ();
 sg13g2_fill_1 FILLER_72_2450 ();
 sg13g2_fill_1 FILLER_72_2477 ();
 sg13g2_fill_1 FILLER_72_2509 ();
 sg13g2_fill_2 FILLER_72_2515 ();
 sg13g2_fill_1 FILLER_72_2562 ();
 sg13g2_decap_8 FILLER_72_2607 ();
 sg13g2_decap_8 FILLER_72_2614 ();
 sg13g2_decap_8 FILLER_72_2621 ();
 sg13g2_decap_8 FILLER_72_2628 ();
 sg13g2_decap_8 FILLER_72_2635 ();
 sg13g2_decap_8 FILLER_72_2642 ();
 sg13g2_decap_8 FILLER_72_2649 ();
 sg13g2_decap_8 FILLER_72_2656 ();
 sg13g2_decap_8 FILLER_72_2663 ();
 sg13g2_decap_4 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_30 ();
 sg13g2_fill_1 FILLER_73_36 ();
 sg13g2_fill_2 FILLER_73_47 ();
 sg13g2_fill_1 FILLER_73_49 ();
 sg13g2_fill_2 FILLER_73_59 ();
 sg13g2_fill_1 FILLER_73_61 ();
 sg13g2_fill_1 FILLER_73_76 ();
 sg13g2_fill_1 FILLER_73_81 ();
 sg13g2_fill_1 FILLER_73_103 ();
 sg13g2_decap_8 FILLER_73_109 ();
 sg13g2_fill_1 FILLER_73_125 ();
 sg13g2_decap_4 FILLER_73_134 ();
 sg13g2_fill_2 FILLER_73_138 ();
 sg13g2_decap_4 FILLER_73_144 ();
 sg13g2_fill_2 FILLER_73_148 ();
 sg13g2_decap_8 FILLER_73_155 ();
 sg13g2_fill_1 FILLER_73_162 ();
 sg13g2_decap_4 FILLER_73_168 ();
 sg13g2_fill_2 FILLER_73_172 ();
 sg13g2_fill_2 FILLER_73_189 ();
 sg13g2_fill_2 FILLER_73_216 ();
 sg13g2_decap_8 FILLER_73_226 ();
 sg13g2_decap_8 FILLER_73_233 ();
 sg13g2_fill_2 FILLER_73_240 ();
 sg13g2_fill_1 FILLER_73_242 ();
 sg13g2_decap_4 FILLER_73_251 ();
 sg13g2_decap_8 FILLER_73_260 ();
 sg13g2_decap_8 FILLER_73_267 ();
 sg13g2_decap_4 FILLER_73_300 ();
 sg13g2_decap_4 FILLER_73_309 ();
 sg13g2_fill_1 FILLER_73_323 ();
 sg13g2_fill_1 FILLER_73_420 ();
 sg13g2_fill_1 FILLER_73_430 ();
 sg13g2_fill_1 FILLER_73_441 ();
 sg13g2_fill_1 FILLER_73_473 ();
 sg13g2_fill_2 FILLER_73_504 ();
 sg13g2_fill_2 FILLER_73_515 ();
 sg13g2_fill_1 FILLER_73_517 ();
 sg13g2_fill_2 FILLER_73_522 ();
 sg13g2_fill_2 FILLER_73_529 ();
 sg13g2_fill_2 FILLER_73_536 ();
 sg13g2_fill_2 FILLER_73_542 ();
 sg13g2_fill_2 FILLER_73_549 ();
 sg13g2_fill_1 FILLER_73_558 ();
 sg13g2_decap_4 FILLER_73_585 ();
 sg13g2_fill_2 FILLER_73_615 ();
 sg13g2_fill_1 FILLER_73_617 ();
 sg13g2_fill_2 FILLER_73_623 ();
 sg13g2_decap_8 FILLER_73_681 ();
 sg13g2_fill_1 FILLER_73_688 ();
 sg13g2_decap_8 FILLER_73_693 ();
 sg13g2_decap_8 FILLER_73_705 ();
 sg13g2_fill_1 FILLER_73_712 ();
 sg13g2_decap_8 FILLER_73_718 ();
 sg13g2_fill_2 FILLER_73_725 ();
 sg13g2_fill_1 FILLER_73_732 ();
 sg13g2_decap_8 FILLER_73_750 ();
 sg13g2_fill_2 FILLER_73_822 ();
 sg13g2_fill_2 FILLER_73_850 ();
 sg13g2_fill_1 FILLER_73_852 ();
 sg13g2_fill_1 FILLER_73_883 ();
 sg13g2_decap_4 FILLER_73_924 ();
 sg13g2_fill_1 FILLER_73_928 ();
 sg13g2_fill_1 FILLER_73_943 ();
 sg13g2_decap_8 FILLER_73_952 ();
 sg13g2_decap_8 FILLER_73_959 ();
 sg13g2_fill_1 FILLER_73_966 ();
 sg13g2_decap_8 FILLER_73_1000 ();
 sg13g2_decap_4 FILLER_73_1007 ();
 sg13g2_fill_2 FILLER_73_1011 ();
 sg13g2_decap_8 FILLER_73_1029 ();
 sg13g2_fill_1 FILLER_73_1036 ();
 sg13g2_decap_4 FILLER_73_1045 ();
 sg13g2_fill_2 FILLER_73_1049 ();
 sg13g2_fill_2 FILLER_73_1061 ();
 sg13g2_fill_1 FILLER_73_1063 ();
 sg13g2_fill_2 FILLER_73_1090 ();
 sg13g2_fill_2 FILLER_73_1119 ();
 sg13g2_decap_8 FILLER_73_1125 ();
 sg13g2_decap_4 FILLER_73_1132 ();
 sg13g2_fill_1 FILLER_73_1136 ();
 sg13g2_decap_4 FILLER_73_1184 ();
 sg13g2_decap_8 FILLER_73_1215 ();
 sg13g2_fill_2 FILLER_73_1222 ();
 sg13g2_fill_1 FILLER_73_1224 ();
 sg13g2_decap_4 FILLER_73_1255 ();
 sg13g2_fill_2 FILLER_73_1324 ();
 sg13g2_decap_8 FILLER_73_1356 ();
 sg13g2_fill_2 FILLER_73_1363 ();
 sg13g2_fill_2 FILLER_73_1411 ();
 sg13g2_fill_2 FILLER_73_1479 ();
 sg13g2_decap_8 FILLER_73_1486 ();
 sg13g2_fill_2 FILLER_73_1493 ();
 sg13g2_fill_1 FILLER_73_1495 ();
 sg13g2_fill_1 FILLER_73_1500 ();
 sg13g2_fill_1 FILLER_73_1508 ();
 sg13g2_fill_2 FILLER_73_1540 ();
 sg13g2_fill_2 FILLER_73_1566 ();
 sg13g2_decap_4 FILLER_73_1576 ();
 sg13g2_fill_1 FILLER_73_1580 ();
 sg13g2_fill_2 FILLER_73_1587 ();
 sg13g2_fill_1 FILLER_73_1589 ();
 sg13g2_fill_1 FILLER_73_1603 ();
 sg13g2_decap_8 FILLER_73_1608 ();
 sg13g2_fill_1 FILLER_73_1615 ();
 sg13g2_fill_1 FILLER_73_1638 ();
 sg13g2_decap_4 FILLER_73_1643 ();
 sg13g2_fill_2 FILLER_73_1647 ();
 sg13g2_decap_8 FILLER_73_1653 ();
 sg13g2_decap_4 FILLER_73_1660 ();
 sg13g2_fill_1 FILLER_73_1664 ();
 sg13g2_decap_4 FILLER_73_1678 ();
 sg13g2_fill_2 FILLER_73_1682 ();
 sg13g2_decap_4 FILLER_73_1692 ();
 sg13g2_decap_8 FILLER_73_1701 ();
 sg13g2_decap_4 FILLER_73_1708 ();
 sg13g2_fill_2 FILLER_73_1724 ();
 sg13g2_fill_2 FILLER_73_1756 ();
 sg13g2_decap_8 FILLER_73_1780 ();
 sg13g2_decap_8 FILLER_73_1787 ();
 sg13g2_fill_2 FILLER_73_1794 ();
 sg13g2_fill_1 FILLER_73_1796 ();
 sg13g2_decap_8 FILLER_73_1805 ();
 sg13g2_decap_8 FILLER_73_1812 ();
 sg13g2_decap_4 FILLER_73_1819 ();
 sg13g2_fill_2 FILLER_73_1823 ();
 sg13g2_fill_2 FILLER_73_1829 ();
 sg13g2_fill_1 FILLER_73_1842 ();
 sg13g2_decap_8 FILLER_73_1853 ();
 sg13g2_fill_2 FILLER_73_1860 ();
 sg13g2_decap_4 FILLER_73_1886 ();
 sg13g2_fill_2 FILLER_73_1911 ();
 sg13g2_decap_4 FILLER_73_1919 ();
 sg13g2_fill_2 FILLER_73_1923 ();
 sg13g2_fill_2 FILLER_73_1930 ();
 sg13g2_fill_1 FILLER_73_1947 ();
 sg13g2_fill_2 FILLER_73_1963 ();
 sg13g2_fill_2 FILLER_73_1979 ();
 sg13g2_fill_2 FILLER_73_1986 ();
 sg13g2_decap_4 FILLER_73_1993 ();
 sg13g2_fill_1 FILLER_73_1997 ();
 sg13g2_decap_8 FILLER_73_2034 ();
 sg13g2_decap_8 FILLER_73_2041 ();
 sg13g2_decap_4 FILLER_73_2048 ();
 sg13g2_fill_2 FILLER_73_2152 ();
 sg13g2_fill_2 FILLER_73_2158 ();
 sg13g2_decap_4 FILLER_73_2170 ();
 sg13g2_fill_2 FILLER_73_2178 ();
 sg13g2_decap_4 FILLER_73_2184 ();
 sg13g2_fill_1 FILLER_73_2188 ();
 sg13g2_fill_2 FILLER_73_2204 ();
 sg13g2_fill_1 FILLER_73_2206 ();
 sg13g2_decap_4 FILLER_73_2212 ();
 sg13g2_fill_2 FILLER_73_2216 ();
 sg13g2_fill_1 FILLER_73_2235 ();
 sg13g2_fill_1 FILLER_73_2262 ();
 sg13g2_fill_2 FILLER_73_2368 ();
 sg13g2_fill_1 FILLER_73_2370 ();
 sg13g2_fill_2 FILLER_73_2382 ();
 sg13g2_fill_1 FILLER_73_2384 ();
 sg13g2_fill_2 FILLER_73_2482 ();
 sg13g2_fill_2 FILLER_73_2488 ();
 sg13g2_fill_1 FILLER_73_2490 ();
 sg13g2_decap_8 FILLER_73_2549 ();
 sg13g2_decap_8 FILLER_73_2556 ();
 sg13g2_decap_8 FILLER_73_2563 ();
 sg13g2_decap_4 FILLER_73_2570 ();
 sg13g2_fill_1 FILLER_73_2574 ();
 sg13g2_decap_8 FILLER_73_2609 ();
 sg13g2_decap_8 FILLER_73_2616 ();
 sg13g2_decap_8 FILLER_73_2623 ();
 sg13g2_decap_8 FILLER_73_2630 ();
 sg13g2_decap_8 FILLER_73_2637 ();
 sg13g2_decap_8 FILLER_73_2644 ();
 sg13g2_decap_8 FILLER_73_2651 ();
 sg13g2_decap_8 FILLER_73_2658 ();
 sg13g2_decap_4 FILLER_73_2665 ();
 sg13g2_fill_1 FILLER_73_2669 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_fill_2 FILLER_74_14 ();
 sg13g2_fill_2 FILLER_74_26 ();
 sg13g2_fill_2 FILLER_74_54 ();
 sg13g2_decap_4 FILLER_74_61 ();
 sg13g2_decap_4 FILLER_74_75 ();
 sg13g2_fill_1 FILLER_74_84 ();
 sg13g2_fill_1 FILLER_74_106 ();
 sg13g2_fill_2 FILLER_74_112 ();
 sg13g2_fill_1 FILLER_74_114 ();
 sg13g2_decap_8 FILLER_74_156 ();
 sg13g2_decap_8 FILLER_74_163 ();
 sg13g2_decap_8 FILLER_74_170 ();
 sg13g2_fill_2 FILLER_74_177 ();
 sg13g2_fill_1 FILLER_74_179 ();
 sg13g2_fill_2 FILLER_74_193 ();
 sg13g2_fill_2 FILLER_74_239 ();
 sg13g2_fill_2 FILLER_74_267 ();
 sg13g2_decap_4 FILLER_74_278 ();
 sg13g2_decap_8 FILLER_74_316 ();
 sg13g2_decap_8 FILLER_74_323 ();
 sg13g2_decap_4 FILLER_74_330 ();
 sg13g2_fill_2 FILLER_74_365 ();
 sg13g2_fill_1 FILLER_74_415 ();
 sg13g2_fill_1 FILLER_74_424 ();
 sg13g2_fill_1 FILLER_74_434 ();
 sg13g2_decap_4 FILLER_74_444 ();
 sg13g2_fill_1 FILLER_74_448 ();
 sg13g2_fill_2 FILLER_74_453 ();
 sg13g2_decap_8 FILLER_74_464 ();
 sg13g2_decap_4 FILLER_74_471 ();
 sg13g2_fill_1 FILLER_74_475 ();
 sg13g2_fill_1 FILLER_74_480 ();
 sg13g2_fill_1 FILLER_74_499 ();
 sg13g2_fill_2 FILLER_74_510 ();
 sg13g2_fill_1 FILLER_74_527 ();
 sg13g2_decap_4 FILLER_74_594 ();
 sg13g2_fill_2 FILLER_74_608 ();
 sg13g2_fill_2 FILLER_74_640 ();
 sg13g2_fill_1 FILLER_74_652 ();
 sg13g2_fill_2 FILLER_74_666 ();
 sg13g2_fill_1 FILLER_74_668 ();
 sg13g2_decap_8 FILLER_74_708 ();
 sg13g2_fill_2 FILLER_74_715 ();
 sg13g2_fill_1 FILLER_74_717 ();
 sg13g2_fill_2 FILLER_74_751 ();
 sg13g2_fill_2 FILLER_74_779 ();
 sg13g2_fill_1 FILLER_74_785 ();
 sg13g2_fill_1 FILLER_74_799 ();
 sg13g2_fill_2 FILLER_74_804 ();
 sg13g2_fill_1 FILLER_74_806 ();
 sg13g2_fill_1 FILLER_74_816 ();
 sg13g2_fill_1 FILLER_74_839 ();
 sg13g2_decap_8 FILLER_74_853 ();
 sg13g2_fill_1 FILLER_74_860 ();
 sg13g2_fill_1 FILLER_74_875 ();
 sg13g2_fill_2 FILLER_74_918 ();
 sg13g2_fill_1 FILLER_74_920 ();
 sg13g2_decap_4 FILLER_74_953 ();
 sg13g2_fill_1 FILLER_74_957 ();
 sg13g2_decap_8 FILLER_74_977 ();
 sg13g2_decap_8 FILLER_74_984 ();
 sg13g2_fill_2 FILLER_74_991 ();
 sg13g2_fill_1 FILLER_74_993 ();
 sg13g2_fill_2 FILLER_74_998 ();
 sg13g2_fill_2 FILLER_74_1004 ();
 sg13g2_fill_2 FILLER_74_1032 ();
 sg13g2_fill_1 FILLER_74_1034 ();
 sg13g2_fill_2 FILLER_74_1083 ();
 sg13g2_fill_2 FILLER_74_1111 ();
 sg13g2_fill_1 FILLER_74_1113 ();
 sg13g2_decap_4 FILLER_74_1124 ();
 sg13g2_decap_8 FILLER_74_1132 ();
 sg13g2_decap_8 FILLER_74_1139 ();
 sg13g2_fill_1 FILLER_74_1146 ();
 sg13g2_fill_2 FILLER_74_1177 ();
 sg13g2_fill_1 FILLER_74_1179 ();
 sg13g2_decap_8 FILLER_74_1210 ();
 sg13g2_decap_8 FILLER_74_1217 ();
 sg13g2_decap_8 FILLER_74_1224 ();
 sg13g2_fill_2 FILLER_74_1231 ();
 sg13g2_fill_1 FILLER_74_1233 ();
 sg13g2_decap_4 FILLER_74_1238 ();
 sg13g2_decap_8 FILLER_74_1310 ();
 sg13g2_decap_8 FILLER_74_1317 ();
 sg13g2_decap_4 FILLER_74_1372 ();
 sg13g2_decap_8 FILLER_74_1402 ();
 sg13g2_decap_8 FILLER_74_1409 ();
 sg13g2_decap_4 FILLER_74_1416 ();
 sg13g2_decap_8 FILLER_74_1430 ();
 sg13g2_fill_1 FILLER_74_1437 ();
 sg13g2_decap_8 FILLER_74_1442 ();
 sg13g2_fill_2 FILLER_74_1449 ();
 sg13g2_fill_2 FILLER_74_1455 ();
 sg13g2_decap_4 FILLER_74_1461 ();
 sg13g2_fill_2 FILLER_74_1465 ();
 sg13g2_decap_8 FILLER_74_1571 ();
 sg13g2_decap_4 FILLER_74_1578 ();
 sg13g2_fill_1 FILLER_74_1582 ();
 sg13g2_decap_8 FILLER_74_1606 ();
 sg13g2_decap_8 FILLER_74_1613 ();
 sg13g2_fill_2 FILLER_74_1620 ();
 sg13g2_decap_4 FILLER_74_1631 ();
 sg13g2_fill_2 FILLER_74_1648 ();
 sg13g2_decap_8 FILLER_74_1654 ();
 sg13g2_decap_8 FILLER_74_1661 ();
 sg13g2_decap_8 FILLER_74_1668 ();
 sg13g2_fill_2 FILLER_74_1675 ();
 sg13g2_fill_1 FILLER_74_1677 ();
 sg13g2_fill_2 FILLER_74_1692 ();
 sg13g2_fill_1 FILLER_74_1707 ();
 sg13g2_fill_2 FILLER_74_1744 ();
 sg13g2_fill_1 FILLER_74_1764 ();
 sg13g2_fill_2 FILLER_74_1774 ();
 sg13g2_decap_4 FILLER_74_1787 ();
 sg13g2_fill_1 FILLER_74_1791 ();
 sg13g2_decap_8 FILLER_74_1801 ();
 sg13g2_decap_8 FILLER_74_1808 ();
 sg13g2_decap_8 FILLER_74_1815 ();
 sg13g2_decap_8 FILLER_74_1822 ();
 sg13g2_fill_1 FILLER_74_1829 ();
 sg13g2_decap_4 FILLER_74_1858 ();
 sg13g2_fill_2 FILLER_74_1889 ();
 sg13g2_fill_1 FILLER_74_1896 ();
 sg13g2_decap_4 FILLER_74_1901 ();
 sg13g2_fill_2 FILLER_74_1905 ();
 sg13g2_fill_2 FILLER_74_1913 ();
 sg13g2_fill_1 FILLER_74_1915 ();
 sg13g2_fill_2 FILLER_74_1920 ();
 sg13g2_fill_1 FILLER_74_1922 ();
 sg13g2_decap_4 FILLER_74_1927 ();
 sg13g2_fill_2 FILLER_74_1931 ();
 sg13g2_fill_1 FILLER_74_1938 ();
 sg13g2_fill_2 FILLER_74_1943 ();
 sg13g2_fill_2 FILLER_74_1950 ();
 sg13g2_fill_2 FILLER_74_1957 ();
 sg13g2_fill_2 FILLER_74_1963 ();
 sg13g2_fill_1 FILLER_74_1965 ();
 sg13g2_fill_1 FILLER_74_1970 ();
 sg13g2_fill_2 FILLER_74_1976 ();
 sg13g2_fill_2 FILLER_74_1983 ();
 sg13g2_fill_2 FILLER_74_1989 ();
 sg13g2_decap_4 FILLER_74_1996 ();
 sg13g2_fill_2 FILLER_74_2000 ();
 sg13g2_decap_8 FILLER_74_2042 ();
 sg13g2_decap_8 FILLER_74_2049 ();
 sg13g2_fill_2 FILLER_74_2056 ();
 sg13g2_fill_1 FILLER_74_2058 ();
 sg13g2_decap_8 FILLER_74_2076 ();
 sg13g2_decap_8 FILLER_74_2083 ();
 sg13g2_decap_8 FILLER_74_2090 ();
 sg13g2_fill_1 FILLER_74_2097 ();
 sg13g2_decap_4 FILLER_74_2102 ();
 sg13g2_fill_1 FILLER_74_2106 ();
 sg13g2_decap_8 FILLER_74_2110 ();
 sg13g2_decap_4 FILLER_74_2117 ();
 sg13g2_decap_8 FILLER_74_2135 ();
 sg13g2_decap_8 FILLER_74_2142 ();
 sg13g2_decap_8 FILLER_74_2149 ();
 sg13g2_decap_8 FILLER_74_2156 ();
 sg13g2_decap_8 FILLER_74_2184 ();
 sg13g2_decap_8 FILLER_74_2191 ();
 sg13g2_fill_2 FILLER_74_2198 ();
 sg13g2_decap_8 FILLER_74_2204 ();
 sg13g2_decap_8 FILLER_74_2211 ();
 sg13g2_decap_8 FILLER_74_2218 ();
 sg13g2_decap_4 FILLER_74_2225 ();
 sg13g2_fill_2 FILLER_74_2239 ();
 sg13g2_fill_2 FILLER_74_2267 ();
 sg13g2_fill_2 FILLER_74_2295 ();
 sg13g2_decap_4 FILLER_74_2356 ();
 sg13g2_fill_1 FILLER_74_2402 ();
 sg13g2_decap_4 FILLER_74_2407 ();
 sg13g2_fill_2 FILLER_74_2437 ();
 sg13g2_fill_2 FILLER_74_2448 ();
 sg13g2_decap_8 FILLER_74_2468 ();
 sg13g2_decap_4 FILLER_74_2485 ();
 sg13g2_fill_1 FILLER_74_2489 ();
 sg13g2_decap_8 FILLER_74_2504 ();
 sg13g2_fill_1 FILLER_74_2511 ();
 sg13g2_fill_2 FILLER_74_2537 ();
 sg13g2_decap_8 FILLER_74_2565 ();
 sg13g2_decap_8 FILLER_74_2572 ();
 sg13g2_decap_8 FILLER_74_2579 ();
 sg13g2_decap_8 FILLER_74_2586 ();
 sg13g2_decap_8 FILLER_74_2593 ();
 sg13g2_decap_8 FILLER_74_2600 ();
 sg13g2_decap_8 FILLER_74_2607 ();
 sg13g2_decap_8 FILLER_74_2614 ();
 sg13g2_decap_8 FILLER_74_2621 ();
 sg13g2_decap_8 FILLER_74_2628 ();
 sg13g2_decap_8 FILLER_74_2635 ();
 sg13g2_decap_8 FILLER_74_2642 ();
 sg13g2_decap_8 FILLER_74_2649 ();
 sg13g2_decap_8 FILLER_74_2656 ();
 sg13g2_decap_8 FILLER_74_2663 ();
 sg13g2_decap_4 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_4 ();
 sg13g2_fill_1 FILLER_75_31 ();
 sg13g2_fill_1 FILLER_75_37 ();
 sg13g2_fill_1 FILLER_75_42 ();
 sg13g2_fill_2 FILLER_75_53 ();
 sg13g2_decap_4 FILLER_75_65 ();
 sg13g2_fill_1 FILLER_75_69 ();
 sg13g2_decap_4 FILLER_75_80 ();
 sg13g2_decap_8 FILLER_75_110 ();
 sg13g2_decap_4 FILLER_75_158 ();
 sg13g2_fill_2 FILLER_75_229 ();
 sg13g2_fill_1 FILLER_75_244 ();
 sg13g2_decap_8 FILLER_75_253 ();
 sg13g2_decap_4 FILLER_75_260 ();
 sg13g2_fill_2 FILLER_75_264 ();
 sg13g2_fill_2 FILLER_75_299 ();
 sg13g2_decap_4 FILLER_75_314 ();
 sg13g2_fill_2 FILLER_75_318 ();
 sg13g2_decap_8 FILLER_75_324 ();
 sg13g2_fill_2 FILLER_75_331 ();
 sg13g2_fill_2 FILLER_75_343 ();
 sg13g2_fill_1 FILLER_75_345 ();
 sg13g2_decap_4 FILLER_75_426 ();
 sg13g2_fill_2 FILLER_75_430 ();
 sg13g2_fill_1 FILLER_75_443 ();
 sg13g2_fill_1 FILLER_75_479 ();
 sg13g2_fill_2 FILLER_75_485 ();
 sg13g2_fill_1 FILLER_75_487 ();
 sg13g2_fill_2 FILLER_75_492 ();
 sg13g2_fill_2 FILLER_75_506 ();
 sg13g2_fill_2 FILLER_75_537 ();
 sg13g2_fill_1 FILLER_75_539 ();
 sg13g2_fill_2 FILLER_75_561 ();
 sg13g2_decap_4 FILLER_75_572 ();
 sg13g2_fill_2 FILLER_75_581 ();
 sg13g2_fill_2 FILLER_75_587 ();
 sg13g2_fill_1 FILLER_75_589 ();
 sg13g2_fill_2 FILLER_75_594 ();
 sg13g2_fill_1 FILLER_75_601 ();
 sg13g2_fill_1 FILLER_75_607 ();
 sg13g2_fill_2 FILLER_75_629 ();
 sg13g2_fill_1 FILLER_75_636 ();
 sg13g2_fill_2 FILLER_75_641 ();
 sg13g2_fill_2 FILLER_75_647 ();
 sg13g2_fill_2 FILLER_75_653 ();
 sg13g2_decap_8 FILLER_75_661 ();
 sg13g2_fill_2 FILLER_75_668 ();
 sg13g2_fill_2 FILLER_75_675 ();
 sg13g2_decap_4 FILLER_75_712 ();
 sg13g2_decap_8 FILLER_75_754 ();
 sg13g2_fill_1 FILLER_75_761 ();
 sg13g2_decap_8 FILLER_75_794 ();
 sg13g2_decap_8 FILLER_75_801 ();
 sg13g2_decap_4 FILLER_75_808 ();
 sg13g2_decap_8 FILLER_75_838 ();
 sg13g2_decap_8 FILLER_75_845 ();
 sg13g2_decap_8 FILLER_75_852 ();
 sg13g2_decap_4 FILLER_75_859 ();
 sg13g2_fill_1 FILLER_75_863 ();
 sg13g2_decap_8 FILLER_75_883 ();
 sg13g2_fill_1 FILLER_75_890 ();
 sg13g2_fill_2 FILLER_75_895 ();
 sg13g2_fill_1 FILLER_75_904 ();
 sg13g2_fill_2 FILLER_75_922 ();
 sg13g2_fill_1 FILLER_75_924 ();
 sg13g2_fill_2 FILLER_75_955 ();
 sg13g2_fill_1 FILLER_75_957 ();
 sg13g2_fill_2 FILLER_75_995 ();
 sg13g2_decap_8 FILLER_75_1027 ();
 sg13g2_decap_4 FILLER_75_1050 ();
 sg13g2_fill_1 FILLER_75_1088 ();
 sg13g2_fill_2 FILLER_75_1104 ();
 sg13g2_fill_1 FILLER_75_1106 ();
 sg13g2_decap_4 FILLER_75_1148 ();
 sg13g2_fill_2 FILLER_75_1152 ();
 sg13g2_decap_8 FILLER_75_1158 ();
 sg13g2_fill_2 FILLER_75_1165 ();
 sg13g2_fill_1 FILLER_75_1167 ();
 sg13g2_fill_2 FILLER_75_1182 ();
 sg13g2_fill_1 FILLER_75_1220 ();
 sg13g2_fill_1 FILLER_75_1264 ();
 sg13g2_fill_1 FILLER_75_1286 ();
 sg13g2_decap_8 FILLER_75_1313 ();
 sg13g2_decap_8 FILLER_75_1320 ();
 sg13g2_decap_4 FILLER_75_1327 ();
 sg13g2_decap_8 FILLER_75_1341 ();
 sg13g2_fill_2 FILLER_75_1348 ();
 sg13g2_fill_1 FILLER_75_1350 ();
 sg13g2_decap_4 FILLER_75_1395 ();
 sg13g2_fill_1 FILLER_75_1399 ();
 sg13g2_decap_8 FILLER_75_1456 ();
 sg13g2_decap_4 FILLER_75_1463 ();
 sg13g2_decap_8 FILLER_75_1477 ();
 sg13g2_decap_4 FILLER_75_1484 ();
 sg13g2_decap_8 FILLER_75_1492 ();
 sg13g2_fill_2 FILLER_75_1499 ();
 sg13g2_fill_1 FILLER_75_1501 ();
 sg13g2_fill_2 FILLER_75_1506 ();
 sg13g2_decap_4 FILLER_75_1554 ();
 sg13g2_fill_1 FILLER_75_1558 ();
 sg13g2_fill_2 FILLER_75_1562 ();
 sg13g2_fill_1 FILLER_75_1564 ();
 sg13g2_decap_8 FILLER_75_1579 ();
 sg13g2_decap_4 FILLER_75_1586 ();
 sg13g2_decap_4 FILLER_75_1599 ();
 sg13g2_fill_2 FILLER_75_1603 ();
 sg13g2_fill_1 FILLER_75_1620 ();
 sg13g2_fill_1 FILLER_75_1626 ();
 sg13g2_fill_2 FILLER_75_1645 ();
 sg13g2_decap_4 FILLER_75_1656 ();
 sg13g2_decap_8 FILLER_75_1666 ();
 sg13g2_fill_1 FILLER_75_1688 ();
 sg13g2_decap_4 FILLER_75_1703 ();
 sg13g2_fill_2 FILLER_75_1707 ();
 sg13g2_fill_1 FILLER_75_1721 ();
 sg13g2_decap_4 FILLER_75_1731 ();
 sg13g2_fill_2 FILLER_75_1781 ();
 sg13g2_fill_1 FILLER_75_1787 ();
 sg13g2_decap_8 FILLER_75_1818 ();
 sg13g2_decap_8 FILLER_75_1825 ();
 sg13g2_fill_1 FILLER_75_1832 ();
 sg13g2_fill_2 FILLER_75_1848 ();
 sg13g2_fill_2 FILLER_75_1874 ();
 sg13g2_fill_1 FILLER_75_1903 ();
 sg13g2_fill_2 FILLER_75_1909 ();
 sg13g2_fill_2 FILLER_75_1926 ();
 sg13g2_fill_1 FILLER_75_1937 ();
 sg13g2_decap_8 FILLER_75_1955 ();
 sg13g2_decap_8 FILLER_75_1962 ();
 sg13g2_decap_8 FILLER_75_1969 ();
 sg13g2_decap_8 FILLER_75_1976 ();
 sg13g2_decap_8 FILLER_75_1983 ();
 sg13g2_decap_8 FILLER_75_1990 ();
 sg13g2_decap_8 FILLER_75_1997 ();
 sg13g2_decap_8 FILLER_75_2008 ();
 sg13g2_fill_1 FILLER_75_2015 ();
 sg13g2_decap_8 FILLER_75_2020 ();
 sg13g2_decap_8 FILLER_75_2027 ();
 sg13g2_decap_8 FILLER_75_2034 ();
 sg13g2_decap_8 FILLER_75_2041 ();
 sg13g2_fill_1 FILLER_75_2062 ();
 sg13g2_decap_8 FILLER_75_2104 ();
 sg13g2_decap_8 FILLER_75_2111 ();
 sg13g2_fill_1 FILLER_75_2118 ();
 sg13g2_decap_8 FILLER_75_2180 ();
 sg13g2_fill_2 FILLER_75_2187 ();
 sg13g2_fill_1 FILLER_75_2189 ();
 sg13g2_fill_2 FILLER_75_2200 ();
 sg13g2_decap_8 FILLER_75_2223 ();
 sg13g2_decap_8 FILLER_75_2230 ();
 sg13g2_fill_2 FILLER_75_2237 ();
 sg13g2_fill_2 FILLER_75_2253 ();
 sg13g2_fill_2 FILLER_75_2265 ();
 sg13g2_fill_1 FILLER_75_2329 ();
 sg13g2_decap_8 FILLER_75_2334 ();
 sg13g2_fill_2 FILLER_75_2341 ();
 sg13g2_fill_1 FILLER_75_2347 ();
 sg13g2_fill_2 FILLER_75_2353 ();
 sg13g2_fill_1 FILLER_75_2381 ();
 sg13g2_fill_2 FILLER_75_2430 ();
 sg13g2_decap_4 FILLER_75_2445 ();
 sg13g2_fill_1 FILLER_75_2449 ();
 sg13g2_fill_2 FILLER_75_2455 ();
 sg13g2_fill_2 FILLER_75_2461 ();
 sg13g2_decap_8 FILLER_75_2467 ();
 sg13g2_decap_8 FILLER_75_2478 ();
 sg13g2_decap_8 FILLER_75_2485 ();
 sg13g2_decap_4 FILLER_75_2492 ();
 sg13g2_fill_2 FILLER_75_2496 ();
 sg13g2_fill_1 FILLER_75_2533 ();
 sg13g2_fill_2 FILLER_75_2538 ();
 sg13g2_fill_1 FILLER_75_2540 ();
 sg13g2_decap_8 FILLER_75_2549 ();
 sg13g2_decap_8 FILLER_75_2556 ();
 sg13g2_decap_8 FILLER_75_2563 ();
 sg13g2_decap_8 FILLER_75_2570 ();
 sg13g2_decap_8 FILLER_75_2577 ();
 sg13g2_decap_8 FILLER_75_2584 ();
 sg13g2_decap_8 FILLER_75_2591 ();
 sg13g2_decap_8 FILLER_75_2598 ();
 sg13g2_decap_8 FILLER_75_2605 ();
 sg13g2_decap_8 FILLER_75_2612 ();
 sg13g2_decap_8 FILLER_75_2619 ();
 sg13g2_decap_8 FILLER_75_2626 ();
 sg13g2_decap_8 FILLER_75_2633 ();
 sg13g2_decap_8 FILLER_75_2640 ();
 sg13g2_decap_8 FILLER_75_2647 ();
 sg13g2_decap_8 FILLER_75_2654 ();
 sg13g2_decap_8 FILLER_75_2661 ();
 sg13g2_fill_2 FILLER_75_2668 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_4 FILLER_76_7 ();
 sg13g2_decap_4 FILLER_76_15 ();
 sg13g2_decap_4 FILLER_76_49 ();
 sg13g2_fill_1 FILLER_76_53 ();
 sg13g2_fill_1 FILLER_76_89 ();
 sg13g2_fill_2 FILLER_76_95 ();
 sg13g2_fill_2 FILLER_76_102 ();
 sg13g2_fill_1 FILLER_76_109 ();
 sg13g2_fill_2 FILLER_76_115 ();
 sg13g2_fill_1 FILLER_76_117 ();
 sg13g2_fill_1 FILLER_76_165 ();
 sg13g2_fill_1 FILLER_76_192 ();
 sg13g2_decap_4 FILLER_76_277 ();
 sg13g2_fill_1 FILLER_76_281 ();
 sg13g2_decap_8 FILLER_76_339 ();
 sg13g2_decap_4 FILLER_76_346 ();
 sg13g2_fill_1 FILLER_76_380 ();
 sg13g2_fill_2 FILLER_76_393 ();
 sg13g2_fill_2 FILLER_76_422 ();
 sg13g2_decap_4 FILLER_76_429 ();
 sg13g2_fill_2 FILLER_76_433 ();
 sg13g2_fill_2 FILLER_76_439 ();
 sg13g2_fill_1 FILLER_76_450 ();
 sg13g2_fill_2 FILLER_76_456 ();
 sg13g2_decap_8 FILLER_76_462 ();
 sg13g2_fill_1 FILLER_76_469 ();
 sg13g2_fill_1 FILLER_76_475 ();
 sg13g2_fill_2 FILLER_76_486 ();
 sg13g2_fill_1 FILLER_76_516 ();
 sg13g2_fill_1 FILLER_76_522 ();
 sg13g2_fill_1 FILLER_76_557 ();
 sg13g2_fill_2 FILLER_76_563 ();
 sg13g2_fill_1 FILLER_76_565 ();
 sg13g2_decap_4 FILLER_76_570 ();
 sg13g2_fill_2 FILLER_76_574 ();
 sg13g2_fill_1 FILLER_76_580 ();
 sg13g2_decap_4 FILLER_76_586 ();
 sg13g2_fill_2 FILLER_76_590 ();
 sg13g2_decap_4 FILLER_76_597 ();
 sg13g2_fill_2 FILLER_76_601 ();
 sg13g2_fill_2 FILLER_76_608 ();
 sg13g2_fill_1 FILLER_76_610 ();
 sg13g2_fill_1 FILLER_76_615 ();
 sg13g2_fill_1 FILLER_76_620 ();
 sg13g2_decap_4 FILLER_76_626 ();
 sg13g2_fill_1 FILLER_76_630 ();
 sg13g2_fill_1 FILLER_76_687 ();
 sg13g2_fill_2 FILLER_76_698 ();
 sg13g2_decap_8 FILLER_76_706 ();
 sg13g2_decap_4 FILLER_76_713 ();
 sg13g2_fill_1 FILLER_76_717 ();
 sg13g2_fill_2 FILLER_76_792 ();
 sg13g2_fill_1 FILLER_76_794 ();
 sg13g2_fill_1 FILLER_76_804 ();
 sg13g2_decap_4 FILLER_76_809 ();
 sg13g2_fill_1 FILLER_76_817 ();
 sg13g2_fill_1 FILLER_76_823 ();
 sg13g2_fill_1 FILLER_76_829 ();
 sg13g2_fill_2 FILLER_76_856 ();
 sg13g2_fill_2 FILLER_76_862 ();
 sg13g2_fill_2 FILLER_76_914 ();
 sg13g2_fill_1 FILLER_76_916 ();
 sg13g2_fill_2 FILLER_76_932 ();
 sg13g2_fill_1 FILLER_76_989 ();
 sg13g2_decap_8 FILLER_76_994 ();
 sg13g2_fill_2 FILLER_76_1001 ();
 sg13g2_fill_1 FILLER_76_1003 ();
 sg13g2_decap_8 FILLER_76_1020 ();
 sg13g2_decap_4 FILLER_76_1027 ();
 sg13g2_fill_1 FILLER_76_1031 ();
 sg13g2_fill_2 FILLER_76_1081 ();
 sg13g2_fill_1 FILLER_76_1083 ();
 sg13g2_decap_8 FILLER_76_1156 ();
 sg13g2_decap_8 FILLER_76_1163 ();
 sg13g2_fill_2 FILLER_76_1170 ();
 sg13g2_decap_4 FILLER_76_1220 ();
 sg13g2_fill_2 FILLER_76_1224 ();
 sg13g2_decap_8 FILLER_76_1229 ();
 sg13g2_fill_2 FILLER_76_1236 ();
 sg13g2_decap_4 FILLER_76_1241 ();
 sg13g2_fill_2 FILLER_76_1245 ();
 sg13g2_decap_4 FILLER_76_1283 ();
 sg13g2_fill_2 FILLER_76_1304 ();
 sg13g2_fill_1 FILLER_76_1306 ();
 sg13g2_decap_8 FILLER_76_1343 ();
 sg13g2_decap_8 FILLER_76_1350 ();
 sg13g2_fill_1 FILLER_76_1357 ();
 sg13g2_decap_8 FILLER_76_1368 ();
 sg13g2_fill_1 FILLER_76_1392 ();
 sg13g2_decap_8 FILLER_76_1429 ();
 sg13g2_fill_2 FILLER_76_1436 ();
 sg13g2_fill_1 FILLER_76_1438 ();
 sg13g2_decap_4 FILLER_76_1449 ();
 sg13g2_fill_2 FILLER_76_1493 ();
 sg13g2_fill_2 FILLER_76_1569 ();
 sg13g2_fill_1 FILLER_76_1571 ();
 sg13g2_fill_2 FILLER_76_1577 ();
 sg13g2_fill_1 FILLER_76_1579 ();
 sg13g2_fill_1 FILLER_76_1604 ();
 sg13g2_fill_1 FILLER_76_1618 ();
 sg13g2_fill_1 FILLER_76_1624 ();
 sg13g2_fill_2 FILLER_76_1650 ();
 sg13g2_decap_4 FILLER_76_1662 ();
 sg13g2_fill_2 FILLER_76_1706 ();
 sg13g2_fill_1 FILLER_76_1753 ();
 sg13g2_fill_1 FILLER_76_1759 ();
 sg13g2_fill_1 FILLER_76_1782 ();
 sg13g2_fill_1 FILLER_76_1788 ();
 sg13g2_fill_2 FILLER_76_1799 ();
 sg13g2_fill_1 FILLER_76_1801 ();
 sg13g2_decap_8 FILLER_76_1812 ();
 sg13g2_decap_8 FILLER_76_1819 ();
 sg13g2_decap_8 FILLER_76_1826 ();
 sg13g2_decap_4 FILLER_76_1833 ();
 sg13g2_fill_1 FILLER_76_1837 ();
 sg13g2_fill_1 FILLER_76_1871 ();
 sg13g2_fill_2 FILLER_76_1880 ();
 sg13g2_fill_2 FILLER_76_1887 ();
 sg13g2_fill_2 FILLER_76_1894 ();
 sg13g2_fill_2 FILLER_76_1902 ();
 sg13g2_fill_1 FILLER_76_1920 ();
 sg13g2_decap_8 FILLER_76_1956 ();
 sg13g2_decap_8 FILLER_76_1967 ();
 sg13g2_decap_8 FILLER_76_1974 ();
 sg13g2_decap_4 FILLER_76_1981 ();
 sg13g2_fill_2 FILLER_76_1985 ();
 sg13g2_decap_8 FILLER_76_2023 ();
 sg13g2_fill_1 FILLER_76_2030 ();
 sg13g2_fill_1 FILLER_76_2041 ();
 sg13g2_fill_1 FILLER_76_2068 ();
 sg13g2_fill_1 FILLER_76_2079 ();
 sg13g2_fill_1 FILLER_76_2106 ();
 sg13g2_decap_8 FILLER_76_2133 ();
 sg13g2_fill_1 FILLER_76_2140 ();
 sg13g2_fill_2 FILLER_76_2151 ();
 sg13g2_decap_4 FILLER_76_2179 ();
 sg13g2_decap_4 FILLER_76_2193 ();
 sg13g2_fill_2 FILLER_76_2223 ();
 sg13g2_fill_1 FILLER_76_2225 ();
 sg13g2_fill_2 FILLER_76_2262 ();
 sg13g2_fill_2 FILLER_76_2303 ();
 sg13g2_fill_2 FILLER_76_2319 ();
 sg13g2_fill_1 FILLER_76_2347 ();
 sg13g2_fill_1 FILLER_76_2354 ();
 sg13g2_fill_2 FILLER_76_2360 ();
 sg13g2_fill_1 FILLER_76_2362 ();
 sg13g2_fill_1 FILLER_76_2380 ();
 sg13g2_decap_8 FILLER_76_2388 ();
 sg13g2_fill_2 FILLER_76_2445 ();
 sg13g2_fill_1 FILLER_76_2447 ();
 sg13g2_decap_4 FILLER_76_2483 ();
 sg13g2_fill_2 FILLER_76_2492 ();
 sg13g2_fill_1 FILLER_76_2494 ();
 sg13g2_decap_8 FILLER_76_2499 ();
 sg13g2_fill_2 FILLER_76_2506 ();
 sg13g2_decap_4 FILLER_76_2512 ();
 sg13g2_decap_4 FILLER_76_2525 ();
 sg13g2_fill_1 FILLER_76_2529 ();
 sg13g2_decap_8 FILLER_76_2556 ();
 sg13g2_decap_8 FILLER_76_2563 ();
 sg13g2_decap_8 FILLER_76_2570 ();
 sg13g2_decap_8 FILLER_76_2577 ();
 sg13g2_decap_8 FILLER_76_2584 ();
 sg13g2_decap_8 FILLER_76_2591 ();
 sg13g2_decap_8 FILLER_76_2598 ();
 sg13g2_decap_8 FILLER_76_2605 ();
 sg13g2_decap_8 FILLER_76_2612 ();
 sg13g2_decap_8 FILLER_76_2619 ();
 sg13g2_decap_8 FILLER_76_2626 ();
 sg13g2_decap_8 FILLER_76_2633 ();
 sg13g2_decap_8 FILLER_76_2640 ();
 sg13g2_decap_8 FILLER_76_2647 ();
 sg13g2_decap_8 FILLER_76_2654 ();
 sg13g2_decap_8 FILLER_76_2661 ();
 sg13g2_fill_2 FILLER_76_2668 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_4 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_29 ();
 sg13g2_fill_1 FILLER_77_36 ();
 sg13g2_fill_1 FILLER_77_47 ();
 sg13g2_fill_2 FILLER_77_58 ();
 sg13g2_fill_2 FILLER_77_87 ();
 sg13g2_fill_1 FILLER_77_99 ();
 sg13g2_fill_1 FILLER_77_110 ();
 sg13g2_fill_1 FILLER_77_116 ();
 sg13g2_fill_2 FILLER_77_121 ();
 sg13g2_fill_2 FILLER_77_126 ();
 sg13g2_fill_2 FILLER_77_159 ();
 sg13g2_fill_1 FILLER_77_248 ();
 sg13g2_fill_2 FILLER_77_284 ();
 sg13g2_fill_1 FILLER_77_286 ();
 sg13g2_fill_1 FILLER_77_308 ();
 sg13g2_fill_2 FILLER_77_314 ();
 sg13g2_decap_4 FILLER_77_337 ();
 sg13g2_fill_1 FILLER_77_341 ();
 sg13g2_decap_4 FILLER_77_346 ();
 sg13g2_fill_1 FILLER_77_350 ();
 sg13g2_fill_2 FILLER_77_381 ();
 sg13g2_fill_1 FILLER_77_386 ();
 sg13g2_fill_2 FILLER_77_395 ();
 sg13g2_fill_1 FILLER_77_424 ();
 sg13g2_fill_1 FILLER_77_504 ();
 sg13g2_decap_8 FILLER_77_550 ();
 sg13g2_decap_4 FILLER_77_593 ();
 sg13g2_fill_1 FILLER_77_597 ();
 sg13g2_fill_2 FILLER_77_613 ();
 sg13g2_fill_1 FILLER_77_620 ();
 sg13g2_fill_1 FILLER_77_720 ();
 sg13g2_fill_2 FILLER_77_726 ();
 sg13g2_fill_2 FILLER_77_738 ();
 sg13g2_fill_2 FILLER_77_748 ();
 sg13g2_fill_1 FILLER_77_750 ();
 sg13g2_fill_2 FILLER_77_777 ();
 sg13g2_fill_2 FILLER_77_789 ();
 sg13g2_fill_2 FILLER_77_795 ();
 sg13g2_fill_1 FILLER_77_797 ();
 sg13g2_fill_1 FILLER_77_853 ();
 sg13g2_fill_2 FILLER_77_880 ();
 sg13g2_fill_1 FILLER_77_882 ();
 sg13g2_decap_8 FILLER_77_912 ();
 sg13g2_decap_4 FILLER_77_919 ();
 sg13g2_fill_1 FILLER_77_949 ();
 sg13g2_decap_4 FILLER_77_1055 ();
 sg13g2_fill_1 FILLER_77_1059 ();
 sg13g2_fill_2 FILLER_77_1112 ();
 sg13g2_fill_1 FILLER_77_1114 ();
 sg13g2_decap_4 FILLER_77_1155 ();
 sg13g2_fill_2 FILLER_77_1206 ();
 sg13g2_fill_1 FILLER_77_1208 ();
 sg13g2_fill_1 FILLER_77_1219 ();
 sg13g2_fill_2 FILLER_77_1224 ();
 sg13g2_fill_2 FILLER_77_1236 ();
 sg13g2_decap_4 FILLER_77_1248 ();
 sg13g2_fill_1 FILLER_77_1252 ();
 sg13g2_fill_1 FILLER_77_1257 ();
 sg13g2_decap_8 FILLER_77_1262 ();
 sg13g2_decap_8 FILLER_77_1269 ();
 sg13g2_fill_1 FILLER_77_1276 ();
 sg13g2_decap_8 FILLER_77_1313 ();
 sg13g2_fill_1 FILLER_77_1334 ();
 sg13g2_decap_4 FILLER_77_1371 ();
 sg13g2_fill_1 FILLER_77_1375 ();
 sg13g2_decap_4 FILLER_77_1402 ();
 sg13g2_fill_2 FILLER_77_1406 ();
 sg13g2_fill_1 FILLER_77_1412 ();
 sg13g2_decap_8 FILLER_77_1423 ();
 sg13g2_fill_2 FILLER_77_1490 ();
 sg13g2_fill_1 FILLER_77_1492 ();
 sg13g2_fill_1 FILLER_77_1549 ();
 sg13g2_fill_2 FILLER_77_1556 ();
 sg13g2_fill_1 FILLER_77_1581 ();
 sg13g2_fill_1 FILLER_77_1588 ();
 sg13g2_fill_2 FILLER_77_1594 ();
 sg13g2_fill_2 FILLER_77_1601 ();
 sg13g2_fill_1 FILLER_77_1644 ();
 sg13g2_decap_4 FILLER_77_1666 ();
 sg13g2_fill_2 FILLER_77_1670 ();
 sg13g2_fill_1 FILLER_77_1680 ();
 sg13g2_fill_2 FILLER_77_1686 ();
 sg13g2_fill_1 FILLER_77_1688 ();
 sg13g2_fill_2 FILLER_77_1753 ();
 sg13g2_fill_1 FILLER_77_1765 ();
 sg13g2_decap_8 FILLER_77_1823 ();
 sg13g2_decap_4 FILLER_77_1830 ();
 sg13g2_decap_4 FILLER_77_1838 ();
 sg13g2_fill_2 FILLER_77_1842 ();
 sg13g2_fill_1 FILLER_77_1875 ();
 sg13g2_fill_1 FILLER_77_1914 ();
 sg13g2_decap_8 FILLER_77_1964 ();
 sg13g2_decap_8 FILLER_77_1971 ();
 sg13g2_fill_1 FILLER_77_1978 ();
 sg13g2_fill_1 FILLER_77_2025 ();
 sg13g2_fill_1 FILLER_77_2030 ();
 sg13g2_fill_1 FILLER_77_2078 ();
 sg13g2_fill_1 FILLER_77_2100 ();
 sg13g2_fill_1 FILLER_77_2111 ();
 sg13g2_fill_1 FILLER_77_2122 ();
 sg13g2_fill_2 FILLER_77_2149 ();
 sg13g2_fill_2 FILLER_77_2155 ();
 sg13g2_fill_2 FILLER_77_2183 ();
 sg13g2_fill_1 FILLER_77_2231 ();
 sg13g2_fill_2 FILLER_77_2253 ();
 sg13g2_fill_1 FILLER_77_2314 ();
 sg13g2_fill_2 FILLER_77_2325 ();
 sg13g2_fill_2 FILLER_77_2358 ();
 sg13g2_fill_1 FILLER_77_2377 ();
 sg13g2_fill_1 FILLER_77_2384 ();
 sg13g2_fill_2 FILLER_77_2435 ();
 sg13g2_decap_8 FILLER_77_2463 ();
 sg13g2_fill_2 FILLER_77_2479 ();
 sg13g2_fill_1 FILLER_77_2481 ();
 sg13g2_decap_8 FILLER_77_2543 ();
 sg13g2_decap_8 FILLER_77_2550 ();
 sg13g2_decap_8 FILLER_77_2557 ();
 sg13g2_decap_8 FILLER_77_2564 ();
 sg13g2_decap_8 FILLER_77_2571 ();
 sg13g2_decap_8 FILLER_77_2578 ();
 sg13g2_decap_8 FILLER_77_2585 ();
 sg13g2_decap_8 FILLER_77_2592 ();
 sg13g2_decap_8 FILLER_77_2599 ();
 sg13g2_decap_8 FILLER_77_2606 ();
 sg13g2_decap_8 FILLER_77_2613 ();
 sg13g2_decap_8 FILLER_77_2620 ();
 sg13g2_decap_8 FILLER_77_2627 ();
 sg13g2_decap_8 FILLER_77_2634 ();
 sg13g2_decap_8 FILLER_77_2641 ();
 sg13g2_decap_8 FILLER_77_2648 ();
 sg13g2_decap_8 FILLER_77_2655 ();
 sg13g2_decap_8 FILLER_77_2662 ();
 sg13g2_fill_1 FILLER_77_2669 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_4 FILLER_78_42 ();
 sg13g2_fill_2 FILLER_78_77 ();
 sg13g2_fill_1 FILLER_78_89 ();
 sg13g2_fill_2 FILLER_78_132 ();
 sg13g2_fill_2 FILLER_78_146 ();
 sg13g2_fill_1 FILLER_78_194 ();
 sg13g2_fill_2 FILLER_78_244 ();
 sg13g2_fill_2 FILLER_78_272 ();
 sg13g2_fill_1 FILLER_78_300 ();
 sg13g2_fill_1 FILLER_78_311 ();
 sg13g2_fill_2 FILLER_78_317 ();
 sg13g2_decap_8 FILLER_78_340 ();
 sg13g2_decap_8 FILLER_78_347 ();
 sg13g2_decap_8 FILLER_78_354 ();
 sg13g2_fill_1 FILLER_78_361 ();
 sg13g2_fill_2 FILLER_78_434 ();
 sg13g2_fill_1 FILLER_78_436 ();
 sg13g2_fill_1 FILLER_78_513 ();
 sg13g2_fill_1 FILLER_78_527 ();
 sg13g2_fill_2 FILLER_78_554 ();
 sg13g2_fill_2 FILLER_78_591 ();
 sg13g2_fill_1 FILLER_78_632 ();
 sg13g2_fill_1 FILLER_78_642 ();
 sg13g2_fill_1 FILLER_78_653 ();
 sg13g2_fill_2 FILLER_78_664 ();
 sg13g2_fill_2 FILLER_78_671 ();
 sg13g2_decap_4 FILLER_78_709 ();
 sg13g2_fill_1 FILLER_78_713 ();
 sg13g2_fill_1 FILLER_78_745 ();
 sg13g2_fill_1 FILLER_78_751 ();
 sg13g2_fill_1 FILLER_78_778 ();
 sg13g2_decap_8 FILLER_78_846 ();
 sg13g2_fill_1 FILLER_78_853 ();
 sg13g2_fill_2 FILLER_78_884 ();
 sg13g2_fill_2 FILLER_78_912 ();
 sg13g2_fill_1 FILLER_78_914 ();
 sg13g2_fill_2 FILLER_78_925 ();
 sg13g2_fill_2 FILLER_78_953 ();
 sg13g2_fill_1 FILLER_78_955 ();
 sg13g2_decap_4 FILLER_78_995 ();
 sg13g2_decap_4 FILLER_78_1029 ();
 sg13g2_fill_1 FILLER_78_1115 ();
 sg13g2_decap_4 FILLER_78_1120 ();
 sg13g2_fill_2 FILLER_78_1124 ();
 sg13g2_decap_4 FILLER_78_1152 ();
 sg13g2_fill_2 FILLER_78_1156 ();
 sg13g2_fill_1 FILLER_78_1184 ();
 sg13g2_decap_4 FILLER_78_1223 ();
 sg13g2_fill_1 FILLER_78_1227 ();
 sg13g2_fill_1 FILLER_78_1254 ();
 sg13g2_decap_4 FILLER_78_1314 ();
 sg13g2_fill_2 FILLER_78_1384 ();
 sg13g2_decap_4 FILLER_78_1458 ();
 sg13g2_fill_1 FILLER_78_1462 ();
 sg13g2_fill_1 FILLER_78_1506 ();
 sg13g2_fill_1 FILLER_78_1533 ();
 sg13g2_fill_1 FILLER_78_1543 ();
 sg13g2_decap_4 FILLER_78_1560 ();
 sg13g2_fill_1 FILLER_78_1564 ();
 sg13g2_fill_1 FILLER_78_1613 ();
 sg13g2_decap_4 FILLER_78_1650 ();
 sg13g2_decap_8 FILLER_78_1659 ();
 sg13g2_decap_8 FILLER_78_1666 ();
 sg13g2_fill_1 FILLER_78_1673 ();
 sg13g2_fill_1 FILLER_78_1683 ();
 sg13g2_fill_1 FILLER_78_1732 ();
 sg13g2_fill_1 FILLER_78_1741 ();
 sg13g2_fill_2 FILLER_78_1758 ();
 sg13g2_fill_1 FILLER_78_1760 ();
 sg13g2_fill_1 FILLER_78_1777 ();
 sg13g2_fill_2 FILLER_78_1782 ();
 sg13g2_fill_1 FILLER_78_1789 ();
 sg13g2_fill_2 FILLER_78_1794 ();
 sg13g2_fill_1 FILLER_78_1796 ();
 sg13g2_fill_1 FILLER_78_1801 ();
 sg13g2_fill_2 FILLER_78_1805 ();
 sg13g2_decap_8 FILLER_78_1837 ();
 sg13g2_decap_8 FILLER_78_1844 ();
 sg13g2_fill_2 FILLER_78_1851 ();
 sg13g2_fill_1 FILLER_78_1853 ();
 sg13g2_fill_1 FILLER_78_1868 ();
 sg13g2_fill_1 FILLER_78_1878 ();
 sg13g2_fill_1 FILLER_78_1883 ();
 sg13g2_fill_2 FILLER_78_1912 ();
 sg13g2_fill_1 FILLER_78_1926 ();
 sg13g2_fill_1 FILLER_78_1956 ();
 sg13g2_decap_8 FILLER_78_1961 ();
 sg13g2_decap_8 FILLER_78_1968 ();
 sg13g2_fill_1 FILLER_78_1975 ();
 sg13g2_decap_4 FILLER_78_2038 ();
 sg13g2_fill_1 FILLER_78_2068 ();
 sg13g2_fill_1 FILLER_78_2108 ();
 sg13g2_fill_1 FILLER_78_2139 ();
 sg13g2_fill_1 FILLER_78_2144 ();
 sg13g2_fill_1 FILLER_78_2155 ();
 sg13g2_fill_1 FILLER_78_2176 ();
 sg13g2_fill_1 FILLER_78_2190 ();
 sg13g2_fill_1 FILLER_78_2221 ();
 sg13g2_decap_8 FILLER_78_2252 ();
 sg13g2_fill_2 FILLER_78_2259 ();
 sg13g2_fill_1 FILLER_78_2265 ();
 sg13g2_decap_4 FILLER_78_2270 ();
 sg13g2_fill_1 FILLER_78_2313 ();
 sg13g2_fill_1 FILLER_78_2340 ();
 sg13g2_fill_2 FILLER_78_2371 ();
 sg13g2_fill_2 FILLER_78_2482 ();
 sg13g2_fill_2 FILLER_78_2489 ();
 sg13g2_fill_1 FILLER_78_2491 ();
 sg13g2_decap_8 FILLER_78_2535 ();
 sg13g2_decap_8 FILLER_78_2542 ();
 sg13g2_decap_8 FILLER_78_2549 ();
 sg13g2_decap_8 FILLER_78_2556 ();
 sg13g2_decap_8 FILLER_78_2563 ();
 sg13g2_decap_8 FILLER_78_2570 ();
 sg13g2_decap_8 FILLER_78_2577 ();
 sg13g2_decap_8 FILLER_78_2584 ();
 sg13g2_decap_8 FILLER_78_2591 ();
 sg13g2_decap_8 FILLER_78_2598 ();
 sg13g2_decap_8 FILLER_78_2605 ();
 sg13g2_decap_8 FILLER_78_2612 ();
 sg13g2_decap_8 FILLER_78_2619 ();
 sg13g2_decap_8 FILLER_78_2626 ();
 sg13g2_decap_8 FILLER_78_2633 ();
 sg13g2_decap_8 FILLER_78_2640 ();
 sg13g2_decap_8 FILLER_78_2647 ();
 sg13g2_decap_8 FILLER_78_2654 ();
 sg13g2_decap_8 FILLER_78_2661 ();
 sg13g2_fill_2 FILLER_78_2668 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_fill_2 FILLER_79_42 ();
 sg13g2_fill_1 FILLER_79_44 ();
 sg13g2_fill_2 FILLER_79_80 ();
 sg13g2_fill_2 FILLER_79_138 ();
 sg13g2_fill_1 FILLER_79_147 ();
 sg13g2_fill_1 FILLER_79_231 ();
 sg13g2_fill_1 FILLER_79_241 ();
 sg13g2_fill_1 FILLER_79_271 ();
 sg13g2_fill_1 FILLER_79_286 ();
 sg13g2_fill_1 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_335 ();
 sg13g2_decap_8 FILLER_79_342 ();
 sg13g2_decap_4 FILLER_79_349 ();
 sg13g2_fill_1 FILLER_79_353 ();
 sg13g2_decap_8 FILLER_79_358 ();
 sg13g2_fill_2 FILLER_79_365 ();
 sg13g2_fill_2 FILLER_79_374 ();
 sg13g2_fill_1 FILLER_79_386 ();
 sg13g2_decap_8 FILLER_79_448 ();
 sg13g2_fill_1 FILLER_79_459 ();
 sg13g2_fill_1 FILLER_79_465 ();
 sg13g2_fill_1 FILLER_79_492 ();
 sg13g2_fill_1 FILLER_79_497 ();
 sg13g2_fill_2 FILLER_79_529 ();
 sg13g2_fill_2 FILLER_79_539 ();
 sg13g2_decap_8 FILLER_79_545 ();
 sg13g2_decap_8 FILLER_79_552 ();
 sg13g2_fill_2 FILLER_79_559 ();
 sg13g2_fill_1 FILLER_79_565 ();
 sg13g2_decap_4 FILLER_79_571 ();
 sg13g2_fill_2 FILLER_79_575 ();
 sg13g2_fill_1 FILLER_79_618 ();
 sg13g2_fill_2 FILLER_79_679 ();
 sg13g2_fill_2 FILLER_79_711 ();
 sg13g2_fill_1 FILLER_79_713 ();
 sg13g2_decap_8 FILLER_79_718 ();
 sg13g2_fill_1 FILLER_79_725 ();
 sg13g2_fill_1 FILLER_79_730 ();
 sg13g2_fill_1 FILLER_79_795 ();
 sg13g2_decap_4 FILLER_79_805 ();
 sg13g2_fill_1 FILLER_79_814 ();
 sg13g2_fill_1 FILLER_79_820 ();
 sg13g2_decap_8 FILLER_79_826 ();
 sg13g2_decap_8 FILLER_79_845 ();
 sg13g2_decap_4 FILLER_79_874 ();
 sg13g2_fill_1 FILLER_79_878 ();
 sg13g2_decap_4 FILLER_79_915 ();
 sg13g2_fill_1 FILLER_79_919 ();
 sg13g2_fill_2 FILLER_79_956 ();
 sg13g2_fill_1 FILLER_79_958 ();
 sg13g2_fill_1 FILLER_79_969 ();
 sg13g2_fill_1 FILLER_79_977 ();
 sg13g2_decap_8 FILLER_79_991 ();
 sg13g2_decap_8 FILLER_79_998 ();
 sg13g2_fill_2 FILLER_79_1009 ();
 sg13g2_fill_1 FILLER_79_1011 ();
 sg13g2_decap_4 FILLER_79_1022 ();
 sg13g2_fill_2 FILLER_79_1026 ();
 sg13g2_fill_2 FILLER_79_1032 ();
 sg13g2_fill_2 FILLER_79_1044 ();
 sg13g2_fill_1 FILLER_79_1046 ();
 sg13g2_fill_2 FILLER_79_1051 ();
 sg13g2_fill_1 FILLER_79_1053 ();
 sg13g2_decap_8 FILLER_79_1061 ();
 sg13g2_decap_8 FILLER_79_1068 ();
 sg13g2_fill_1 FILLER_79_1114 ();
 sg13g2_decap_8 FILLER_79_1125 ();
 sg13g2_fill_2 FILLER_79_1132 ();
 sg13g2_decap_8 FILLER_79_1138 ();
 sg13g2_decap_8 FILLER_79_1145 ();
 sg13g2_decap_4 FILLER_79_1152 ();
 sg13g2_fill_2 FILLER_79_1182 ();
 sg13g2_fill_1 FILLER_79_1184 ();
 sg13g2_fill_2 FILLER_79_1219 ();
 sg13g2_fill_1 FILLER_79_1221 ();
 sg13g2_fill_2 FILLER_79_1248 ();
 sg13g2_fill_1 FILLER_79_1250 ();
 sg13g2_fill_1 FILLER_79_1306 ();
 sg13g2_fill_1 FILLER_79_1317 ();
 sg13g2_decap_4 FILLER_79_1348 ();
 sg13g2_fill_2 FILLER_79_1352 ();
 sg13g2_fill_2 FILLER_79_1385 ();
 sg13g2_decap_8 FILLER_79_1413 ();
 sg13g2_decap_8 FILLER_79_1420 ();
 sg13g2_fill_2 FILLER_79_1427 ();
 sg13g2_decap_8 FILLER_79_1459 ();
 sg13g2_fill_1 FILLER_79_1466 ();
 sg13g2_fill_1 FILLER_79_1505 ();
 sg13g2_decap_8 FILLER_79_1540 ();
 sg13g2_fill_2 FILLER_79_1547 ();
 sg13g2_decap_8 FILLER_79_1556 ();
 sg13g2_decap_4 FILLER_79_1563 ();
 sg13g2_fill_2 FILLER_79_1567 ();
 sg13g2_fill_2 FILLER_79_1606 ();
 sg13g2_fill_1 FILLER_79_1608 ();
 sg13g2_decap_8 FILLER_79_1624 ();
 sg13g2_decap_4 FILLER_79_1641 ();
 sg13g2_decap_4 FILLER_79_1650 ();
 sg13g2_fill_2 FILLER_79_1654 ();
 sg13g2_fill_2 FILLER_79_1682 ();
 sg13g2_fill_1 FILLER_79_1684 ();
 sg13g2_decap_4 FILLER_79_1690 ();
 sg13g2_fill_2 FILLER_79_1694 ();
 sg13g2_fill_2 FILLER_79_1735 ();
 sg13g2_fill_2 FILLER_79_1742 ();
 sg13g2_fill_2 FILLER_79_1748 ();
 sg13g2_fill_1 FILLER_79_1750 ();
 sg13g2_decap_4 FILLER_79_1762 ();
 sg13g2_fill_1 FILLER_79_1766 ();
 sg13g2_decap_8 FILLER_79_1838 ();
 sg13g2_decap_8 FILLER_79_1845 ();
 sg13g2_decap_8 FILLER_79_1852 ();
 sg13g2_decap_4 FILLER_79_1859 ();
 sg13g2_fill_1 FILLER_79_1863 ();
 sg13g2_fill_2 FILLER_79_1885 ();
 sg13g2_fill_1 FILLER_79_1887 ();
 sg13g2_fill_1 FILLER_79_1896 ();
 sg13g2_fill_1 FILLER_79_1901 ();
 sg13g2_fill_1 FILLER_79_1907 ();
 sg13g2_fill_1 FILLER_79_1914 ();
 sg13g2_fill_2 FILLER_79_1920 ();
 sg13g2_fill_1 FILLER_79_1927 ();
 sg13g2_fill_2 FILLER_79_1933 ();
 sg13g2_fill_1 FILLER_79_1935 ();
 sg13g2_fill_2 FILLER_79_1948 ();
 sg13g2_decap_8 FILLER_79_1976 ();
 sg13g2_fill_1 FILLER_79_1983 ();
 sg13g2_decap_8 FILLER_79_2014 ();
 sg13g2_decap_8 FILLER_79_2025 ();
 sg13g2_fill_2 FILLER_79_2032 ();
 sg13g2_decap_4 FILLER_79_2044 ();
 sg13g2_fill_2 FILLER_79_2048 ();
 sg13g2_fill_2 FILLER_79_2054 ();
 sg13g2_fill_2 FILLER_79_2066 ();
 sg13g2_fill_2 FILLER_79_2078 ();
 sg13g2_fill_1 FILLER_79_2080 ();
 sg13g2_fill_2 FILLER_79_2107 ();
 sg13g2_fill_1 FILLER_79_2109 ();
 sg13g2_decap_8 FILLER_79_2175 ();
 sg13g2_fill_1 FILLER_79_2182 ();
 sg13g2_fill_2 FILLER_79_2209 ();
 sg13g2_fill_2 FILLER_79_2215 ();
 sg13g2_fill_1 FILLER_79_2217 ();
 sg13g2_fill_1 FILLER_79_2251 ();
 sg13g2_fill_2 FILLER_79_2278 ();
 sg13g2_fill_1 FILLER_79_2310 ();
 sg13g2_fill_1 FILLER_79_2389 ();
 sg13g2_fill_1 FILLER_79_2416 ();
 sg13g2_fill_1 FILLER_79_2443 ();
 sg13g2_fill_2 FILLER_79_2448 ();
 sg13g2_decap_8 FILLER_79_2454 ();
 sg13g2_fill_1 FILLER_79_2461 ();
 sg13g2_decap_8 FILLER_79_2522 ();
 sg13g2_decap_8 FILLER_79_2529 ();
 sg13g2_decap_8 FILLER_79_2536 ();
 sg13g2_decap_8 FILLER_79_2543 ();
 sg13g2_decap_8 FILLER_79_2550 ();
 sg13g2_decap_8 FILLER_79_2557 ();
 sg13g2_decap_8 FILLER_79_2564 ();
 sg13g2_decap_8 FILLER_79_2571 ();
 sg13g2_decap_8 FILLER_79_2578 ();
 sg13g2_decap_8 FILLER_79_2585 ();
 sg13g2_decap_8 FILLER_79_2592 ();
 sg13g2_decap_8 FILLER_79_2599 ();
 sg13g2_decap_8 FILLER_79_2606 ();
 sg13g2_decap_8 FILLER_79_2613 ();
 sg13g2_decap_8 FILLER_79_2620 ();
 sg13g2_decap_8 FILLER_79_2627 ();
 sg13g2_decap_8 FILLER_79_2634 ();
 sg13g2_decap_8 FILLER_79_2641 ();
 sg13g2_decap_8 FILLER_79_2648 ();
 sg13g2_decap_8 FILLER_79_2655 ();
 sg13g2_decap_8 FILLER_79_2662 ();
 sg13g2_fill_1 FILLER_79_2669 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_60 ();
 sg13g2_decap_8 FILLER_80_67 ();
 sg13g2_decap_8 FILLER_80_74 ();
 sg13g2_fill_1 FILLER_80_81 ();
 sg13g2_fill_1 FILLER_80_98 ();
 sg13g2_fill_1 FILLER_80_134 ();
 sg13g2_fill_2 FILLER_80_170 ();
 sg13g2_fill_1 FILLER_80_199 ();
 sg13g2_fill_2 FILLER_80_215 ();
 sg13g2_fill_1 FILLER_80_264 ();
 sg13g2_fill_1 FILLER_80_276 ();
 sg13g2_fill_2 FILLER_80_281 ();
 sg13g2_decap_8 FILLER_80_307 ();
 sg13g2_decap_4 FILLER_80_314 ();
 sg13g2_decap_8 FILLER_80_342 ();
 sg13g2_decap_4 FILLER_80_349 ();
 sg13g2_fill_1 FILLER_80_353 ();
 sg13g2_decap_8 FILLER_80_366 ();
 sg13g2_decap_4 FILLER_80_373 ();
 sg13g2_fill_2 FILLER_80_381 ();
 sg13g2_fill_1 FILLER_80_383 ();
 sg13g2_fill_2 FILLER_80_390 ();
 sg13g2_decap_4 FILLER_80_395 ();
 sg13g2_fill_1 FILLER_80_399 ();
 sg13g2_decap_8 FILLER_80_408 ();
 sg13g2_fill_1 FILLER_80_415 ();
 sg13g2_decap_4 FILLER_80_425 ();
 sg13g2_decap_8 FILLER_80_437 ();
 sg13g2_decap_4 FILLER_80_444 ();
 sg13g2_fill_1 FILLER_80_448 ();
 sg13g2_decap_4 FILLER_80_454 ();
 sg13g2_fill_2 FILLER_80_458 ();
 sg13g2_decap_8 FILLER_80_464 ();
 sg13g2_fill_1 FILLER_80_471 ();
 sg13g2_decap_8 FILLER_80_476 ();
 sg13g2_decap_8 FILLER_80_483 ();
 sg13g2_decap_8 FILLER_80_490 ();
 sg13g2_decap_8 FILLER_80_497 ();
 sg13g2_fill_2 FILLER_80_504 ();
 sg13g2_fill_1 FILLER_80_506 ();
 sg13g2_decap_8 FILLER_80_511 ();
 sg13g2_decap_8 FILLER_80_528 ();
 sg13g2_decap_8 FILLER_80_535 ();
 sg13g2_decap_8 FILLER_80_542 ();
 sg13g2_decap_8 FILLER_80_549 ();
 sg13g2_decap_8 FILLER_80_556 ();
 sg13g2_decap_8 FILLER_80_563 ();
 sg13g2_decap_8 FILLER_80_570 ();
 sg13g2_decap_8 FILLER_80_577 ();
 sg13g2_decap_8 FILLER_80_584 ();
 sg13g2_decap_8 FILLER_80_591 ();
 sg13g2_decap_8 FILLER_80_606 ();
 sg13g2_decap_8 FILLER_80_613 ();
 sg13g2_decap_8 FILLER_80_624 ();
 sg13g2_fill_2 FILLER_80_631 ();
 sg13g2_fill_2 FILLER_80_637 ();
 sg13g2_decap_4 FILLER_80_644 ();
 sg13g2_decap_8 FILLER_80_652 ();
 sg13g2_decap_8 FILLER_80_667 ();
 sg13g2_decap_8 FILLER_80_674 ();
 sg13g2_decap_8 FILLER_80_681 ();
 sg13g2_fill_2 FILLER_80_688 ();
 sg13g2_decap_8 FILLER_80_694 ();
 sg13g2_decap_8 FILLER_80_701 ();
 sg13g2_decap_8 FILLER_80_708 ();
 sg13g2_decap_8 FILLER_80_715 ();
 sg13g2_decap_8 FILLER_80_722 ();
 sg13g2_decap_8 FILLER_80_729 ();
 sg13g2_fill_2 FILLER_80_736 ();
 sg13g2_fill_1 FILLER_80_738 ();
 sg13g2_decap_8 FILLER_80_743 ();
 sg13g2_decap_8 FILLER_80_750 ();
 sg13g2_decap_8 FILLER_80_757 ();
 sg13g2_fill_1 FILLER_80_764 ();
 sg13g2_fill_1 FILLER_80_787 ();
 sg13g2_decap_8 FILLER_80_818 ();
 sg13g2_decap_8 FILLER_80_825 ();
 sg13g2_decap_8 FILLER_80_832 ();
 sg13g2_decap_8 FILLER_80_839 ();
 sg13g2_decap_8 FILLER_80_846 ();
 sg13g2_decap_8 FILLER_80_853 ();
 sg13g2_decap_8 FILLER_80_860 ();
 sg13g2_decap_8 FILLER_80_867 ();
 sg13g2_decap_8 FILLER_80_874 ();
 sg13g2_fill_2 FILLER_80_881 ();
 sg13g2_fill_2 FILLER_80_887 ();
 sg13g2_fill_1 FILLER_80_889 ();
 sg13g2_fill_1 FILLER_80_894 ();
 sg13g2_decap_4 FILLER_80_899 ();
 sg13g2_decap_8 FILLER_80_913 ();
 sg13g2_decap_8 FILLER_80_920 ();
 sg13g2_fill_1 FILLER_80_927 ();
 sg13g2_fill_2 FILLER_80_936 ();
 sg13g2_fill_1 FILLER_80_938 ();
 sg13g2_decap_8 FILLER_80_943 ();
 sg13g2_decap_8 FILLER_80_950 ();
 sg13g2_decap_4 FILLER_80_957 ();
 sg13g2_fill_2 FILLER_80_973 ();
 sg13g2_fill_1 FILLER_80_988 ();
 sg13g2_decap_8 FILLER_80_1015 ();
 sg13g2_decap_8 FILLER_80_1022 ();
 sg13g2_fill_2 FILLER_80_1029 ();
 sg13g2_decap_8 FILLER_80_1061 ();
 sg13g2_decap_8 FILLER_80_1068 ();
 sg13g2_decap_4 FILLER_80_1075 ();
 sg13g2_fill_1 FILLER_80_1079 ();
 sg13g2_fill_2 FILLER_80_1084 ();
 sg13g2_fill_1 FILLER_80_1086 ();
 sg13g2_decap_8 FILLER_80_1091 ();
 sg13g2_fill_2 FILLER_80_1098 ();
 sg13g2_fill_1 FILLER_80_1100 ();
 sg13g2_fill_2 FILLER_80_1105 ();
 sg13g2_fill_1 FILLER_80_1107 ();
 sg13g2_decap_8 FILLER_80_1138 ();
 sg13g2_decap_8 FILLER_80_1145 ();
 sg13g2_decap_8 FILLER_80_1152 ();
 sg13g2_fill_2 FILLER_80_1159 ();
 sg13g2_fill_1 FILLER_80_1161 ();
 sg13g2_decap_8 FILLER_80_1166 ();
 sg13g2_decap_8 FILLER_80_1173 ();
 sg13g2_decap_8 FILLER_80_1180 ();
 sg13g2_decap_4 FILLER_80_1187 ();
 sg13g2_fill_1 FILLER_80_1191 ();
 sg13g2_decap_4 FILLER_80_1196 ();
 sg13g2_fill_2 FILLER_80_1200 ();
 sg13g2_decap_8 FILLER_80_1206 ();
 sg13g2_decap_8 FILLER_80_1213 ();
 sg13g2_decap_8 FILLER_80_1220 ();
 sg13g2_decap_4 FILLER_80_1227 ();
 sg13g2_decap_4 FILLER_80_1239 ();
 sg13g2_fill_2 FILLER_80_1243 ();
 sg13g2_fill_1 FILLER_80_1274 ();
 sg13g2_fill_1 FILLER_80_1282 ();
 sg13g2_fill_1 FILLER_80_1297 ();
 sg13g2_decap_8 FILLER_80_1302 ();
 sg13g2_decap_8 FILLER_80_1309 ();
 sg13g2_decap_8 FILLER_80_1316 ();
 sg13g2_fill_2 FILLER_80_1323 ();
 sg13g2_fill_1 FILLER_80_1325 ();
 sg13g2_decap_8 FILLER_80_1330 ();
 sg13g2_decap_8 FILLER_80_1337 ();
 sg13g2_decap_8 FILLER_80_1344 ();
 sg13g2_decap_8 FILLER_80_1351 ();
 sg13g2_fill_1 FILLER_80_1358 ();
 sg13g2_fill_1 FILLER_80_1363 ();
 sg13g2_decap_8 FILLER_80_1368 ();
 sg13g2_decap_8 FILLER_80_1375 ();
 sg13g2_fill_1 FILLER_80_1382 ();
 sg13g2_decap_8 FILLER_80_1397 ();
 sg13g2_fill_1 FILLER_80_1404 ();
 sg13g2_decap_8 FILLER_80_1409 ();
 sg13g2_decap_8 FILLER_80_1416 ();
 sg13g2_decap_8 FILLER_80_1423 ();
 sg13g2_fill_1 FILLER_80_1430 ();
 sg13g2_fill_2 FILLER_80_1452 ();
 sg13g2_fill_1 FILLER_80_1480 ();
 sg13g2_fill_1 FILLER_80_1510 ();
 sg13g2_fill_1 FILLER_80_1515 ();
 sg13g2_decap_8 FILLER_80_1544 ();
 sg13g2_decap_8 FILLER_80_1551 ();
 sg13g2_decap_8 FILLER_80_1558 ();
 sg13g2_decap_8 FILLER_80_1565 ();
 sg13g2_decap_4 FILLER_80_1572 ();
 sg13g2_fill_2 FILLER_80_1576 ();
 sg13g2_decap_8 FILLER_80_1591 ();
 sg13g2_decap_4 FILLER_80_1598 ();
 sg13g2_fill_2 FILLER_80_1602 ();
 sg13g2_decap_8 FILLER_80_1608 ();
 sg13g2_decap_8 FILLER_80_1615 ();
 sg13g2_decap_8 FILLER_80_1622 ();
 sg13g2_decap_8 FILLER_80_1629 ();
 sg13g2_decap_8 FILLER_80_1636 ();
 sg13g2_decap_8 FILLER_80_1643 ();
 sg13g2_decap_8 FILLER_80_1650 ();
 sg13g2_decap_4 FILLER_80_1657 ();
 sg13g2_fill_1 FILLER_80_1661 ();
 sg13g2_decap_8 FILLER_80_1666 ();
 sg13g2_decap_8 FILLER_80_1673 ();
 sg13g2_decap_8 FILLER_80_1680 ();
 sg13g2_decap_8 FILLER_80_1687 ();
 sg13g2_decap_8 FILLER_80_1694 ();
 sg13g2_decap_8 FILLER_80_1701 ();
 sg13g2_fill_2 FILLER_80_1708 ();
 sg13g2_fill_1 FILLER_80_1710 ();
 sg13g2_decap_8 FILLER_80_1716 ();
 sg13g2_fill_1 FILLER_80_1723 ();
 sg13g2_decap_4 FILLER_80_1733 ();
 sg13g2_decap_8 FILLER_80_1741 ();
 sg13g2_decap_8 FILLER_80_1748 ();
 sg13g2_decap_8 FILLER_80_1755 ();
 sg13g2_decap_8 FILLER_80_1762 ();
 sg13g2_decap_8 FILLER_80_1769 ();
 sg13g2_fill_2 FILLER_80_1780 ();
 sg13g2_decap_8 FILLER_80_1790 ();
 sg13g2_decap_8 FILLER_80_1797 ();
 sg13g2_fill_2 FILLER_80_1804 ();
 sg13g2_fill_2 FILLER_80_1812 ();
 sg13g2_decap_8 FILLER_80_1822 ();
 sg13g2_decap_8 FILLER_80_1829 ();
 sg13g2_decap_8 FILLER_80_1836 ();
 sg13g2_decap_8 FILLER_80_1843 ();
 sg13g2_decap_8 FILLER_80_1850 ();
 sg13g2_decap_8 FILLER_80_1857 ();
 sg13g2_decap_8 FILLER_80_1864 ();
 sg13g2_decap_4 FILLER_80_1871 ();
 sg13g2_fill_1 FILLER_80_1875 ();
 sg13g2_decap_8 FILLER_80_1880 ();
 sg13g2_fill_2 FILLER_80_1887 ();
 sg13g2_decap_8 FILLER_80_1899 ();
 sg13g2_fill_2 FILLER_80_1906 ();
 sg13g2_fill_1 FILLER_80_1908 ();
 sg13g2_decap_8 FILLER_80_1913 ();
 sg13g2_decap_8 FILLER_80_1920 ();
 sg13g2_decap_8 FILLER_80_1927 ();
 sg13g2_decap_8 FILLER_80_1934 ();
 sg13g2_decap_8 FILLER_80_1941 ();
 sg13g2_decap_8 FILLER_80_1948 ();
 sg13g2_decap_8 FILLER_80_1955 ();
 sg13g2_decap_8 FILLER_80_1962 ();
 sg13g2_decap_8 FILLER_80_1969 ();
 sg13g2_decap_8 FILLER_80_1976 ();
 sg13g2_decap_8 FILLER_80_1983 ();
 sg13g2_fill_2 FILLER_80_1994 ();
 sg13g2_decap_8 FILLER_80_2000 ();
 sg13g2_decap_8 FILLER_80_2007 ();
 sg13g2_decap_8 FILLER_80_2040 ();
 sg13g2_decap_8 FILLER_80_2047 ();
 sg13g2_decap_8 FILLER_80_2054 ();
 sg13g2_decap_8 FILLER_80_2061 ();
 sg13g2_fill_2 FILLER_80_2068 ();
 sg13g2_fill_1 FILLER_80_2070 ();
 sg13g2_decap_8 FILLER_80_2097 ();
 sg13g2_decap_4 FILLER_80_2104 ();
 sg13g2_decap_8 FILLER_80_2136 ();
 sg13g2_decap_8 FILLER_80_2143 ();
 sg13g2_decap_4 FILLER_80_2150 ();
 sg13g2_fill_2 FILLER_80_2154 ();
 sg13g2_fill_2 FILLER_80_2160 ();
 sg13g2_fill_1 FILLER_80_2162 ();
 sg13g2_decap_8 FILLER_80_2167 ();
 sg13g2_decap_8 FILLER_80_2174 ();
 sg13g2_decap_8 FILLER_80_2181 ();
 sg13g2_fill_2 FILLER_80_2188 ();
 sg13g2_decap_4 FILLER_80_2194 ();
 sg13g2_fill_2 FILLER_80_2198 ();
 sg13g2_decap_8 FILLER_80_2204 ();
 sg13g2_decap_8 FILLER_80_2211 ();
 sg13g2_fill_2 FILLER_80_2218 ();
 sg13g2_fill_1 FILLER_80_2220 ();
 sg13g2_decap_8 FILLER_80_2255 ();
 sg13g2_decap_8 FILLER_80_2262 ();
 sg13g2_decap_8 FILLER_80_2269 ();
 sg13g2_decap_8 FILLER_80_2276 ();
 sg13g2_decap_4 FILLER_80_2283 ();
 sg13g2_fill_1 FILLER_80_2287 ();
 sg13g2_fill_2 FILLER_80_2298 ();
 sg13g2_decap_8 FILLER_80_2312 ();
 sg13g2_decap_8 FILLER_80_2327 ();
 sg13g2_decap_8 FILLER_80_2334 ();
 sg13g2_fill_2 FILLER_80_2341 ();
 sg13g2_fill_1 FILLER_80_2343 ();
 sg13g2_decap_8 FILLER_80_2352 ();
 sg13g2_decap_8 FILLER_80_2359 ();
 sg13g2_fill_2 FILLER_80_2366 ();
 sg13g2_fill_1 FILLER_80_2368 ();
 sg13g2_decap_8 FILLER_80_2373 ();
 sg13g2_decap_4 FILLER_80_2380 ();
 sg13g2_decap_8 FILLER_80_2388 ();
 sg13g2_fill_1 FILLER_80_2395 ();
 sg13g2_decap_8 FILLER_80_2410 ();
 sg13g2_fill_2 FILLER_80_2428 ();
 sg13g2_decap_8 FILLER_80_2451 ();
 sg13g2_decap_8 FILLER_80_2458 ();
 sg13g2_decap_8 FILLER_80_2465 ();
 sg13g2_decap_8 FILLER_80_2476 ();
 sg13g2_decap_8 FILLER_80_2487 ();
 sg13g2_fill_1 FILLER_80_2494 ();
 sg13g2_fill_2 FILLER_80_2499 ();
 sg13g2_fill_1 FILLER_80_2501 ();
 sg13g2_decap_8 FILLER_80_2506 ();
 sg13g2_decap_8 FILLER_80_2513 ();
 sg13g2_decap_8 FILLER_80_2520 ();
 sg13g2_decap_8 FILLER_80_2527 ();
 sg13g2_decap_8 FILLER_80_2534 ();
 sg13g2_decap_8 FILLER_80_2541 ();
 sg13g2_decap_8 FILLER_80_2548 ();
 sg13g2_decap_8 FILLER_80_2555 ();
 sg13g2_decap_8 FILLER_80_2562 ();
 sg13g2_decap_8 FILLER_80_2569 ();
 sg13g2_decap_8 FILLER_80_2576 ();
 sg13g2_decap_8 FILLER_80_2583 ();
 sg13g2_decap_8 FILLER_80_2590 ();
 sg13g2_decap_8 FILLER_80_2597 ();
 sg13g2_decap_8 FILLER_80_2604 ();
 sg13g2_decap_8 FILLER_80_2611 ();
 sg13g2_decap_8 FILLER_80_2618 ();
 sg13g2_decap_8 FILLER_80_2625 ();
 sg13g2_decap_8 FILLER_80_2632 ();
 sg13g2_decap_8 FILLER_80_2639 ();
 sg13g2_decap_8 FILLER_80_2646 ();
 sg13g2_decap_8 FILLER_80_2653 ();
 sg13g2_decap_8 FILLER_80_2660 ();
 sg13g2_fill_2 FILLER_80_2667 ();
 sg13g2_fill_1 FILLER_80_2669 ();
endmodule
