module tt_um_rejunity_sn76489 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire clknet_0_clk;
 wire net86;
 wire \chan[0].attenuation.control[0] ;
 wire \chan[0].attenuation.control[1] ;
 wire \chan[0].attenuation.control[2] ;
 wire \chan[0].attenuation.control[3] ;
 wire \chan[0].attenuation.in ;
 wire \chan[1].attenuation.control[0] ;
 wire \chan[1].attenuation.control[1] ;
 wire \chan[1].attenuation.control[2] ;
 wire \chan[1].attenuation.control[3] ;
 wire \chan[1].attenuation.in ;
 wire \chan[2].attenuation.control[0] ;
 wire \chan[2].attenuation.control[1] ;
 wire \chan[2].attenuation.control[2] ;
 wire \chan[2].attenuation.control[3] ;
 wire \chan[2].attenuation.in ;
 wire \chan[3].attenuation.control[0] ;
 wire \chan[3].attenuation.control[1] ;
 wire \chan[3].attenuation.control[2] ;
 wire \chan[3].attenuation.control[3] ;
 wire \chan[3].attenuation.in ;
 wire \clk_counter[0] ;
 wire \clk_counter[1] ;
 wire \clk_counter[2] ;
 wire \clk_counter[3] ;
 wire \clk_counter[4] ;
 wire \clk_counter[5] ;
 wire \clk_counter[6] ;
 wire \control_noise[0][0] ;
 wire \control_noise[0][1] ;
 wire \control_noise[0][2] ;
 wire \control_tone_freq[0][0] ;
 wire \control_tone_freq[0][1] ;
 wire \control_tone_freq[0][2] ;
 wire \control_tone_freq[0][3] ;
 wire \control_tone_freq[0][4] ;
 wire \control_tone_freq[0][5] ;
 wire \control_tone_freq[0][6] ;
 wire \control_tone_freq[0][7] ;
 wire \control_tone_freq[0][8] ;
 wire \control_tone_freq[0][9] ;
 wire \control_tone_freq[1][0] ;
 wire \control_tone_freq[1][1] ;
 wire \control_tone_freq[1][2] ;
 wire \control_tone_freq[1][3] ;
 wire \control_tone_freq[1][4] ;
 wire \control_tone_freq[1][5] ;
 wire \control_tone_freq[1][6] ;
 wire \control_tone_freq[1][7] ;
 wire \control_tone_freq[1][8] ;
 wire \control_tone_freq[1][9] ;
 wire \control_tone_freq[2][0] ;
 wire \control_tone_freq[2][1] ;
 wire \control_tone_freq[2][2] ;
 wire \control_tone_freq[2][3] ;
 wire \control_tone_freq[2][4] ;
 wire \control_tone_freq[2][5] ;
 wire \control_tone_freq[2][6] ;
 wire \control_tone_freq[2][7] ;
 wire \control_tone_freq[2][8] ;
 wire \control_tone_freq[2][9] ;
 wire \genblk4[0].pwm.accumulator[0] ;
 wire \genblk4[0].pwm.accumulator[10] ;
 wire \genblk4[0].pwm.accumulator[1] ;
 wire \genblk4[0].pwm.accumulator[2] ;
 wire \genblk4[0].pwm.accumulator[3] ;
 wire \genblk4[0].pwm.accumulator[4] ;
 wire \genblk4[0].pwm.accumulator[5] ;
 wire \genblk4[0].pwm.accumulator[6] ;
 wire \genblk4[0].pwm.accumulator[7] ;
 wire \genblk4[0].pwm.accumulator[8] ;
 wire \genblk4[0].pwm.accumulator[9] ;
 wire \genblk4[1].pwm.accumulator[0] ;
 wire \genblk4[1].pwm.accumulator[10] ;
 wire \genblk4[1].pwm.accumulator[1] ;
 wire \genblk4[1].pwm.accumulator[2] ;
 wire \genblk4[1].pwm.accumulator[3] ;
 wire \genblk4[1].pwm.accumulator[4] ;
 wire \genblk4[1].pwm.accumulator[5] ;
 wire \genblk4[1].pwm.accumulator[6] ;
 wire \genblk4[1].pwm.accumulator[7] ;
 wire \genblk4[1].pwm.accumulator[8] ;
 wire \genblk4[1].pwm.accumulator[9] ;
 wire \genblk4[2].pwm.accumulator[0] ;
 wire \genblk4[2].pwm.accumulator[10] ;
 wire \genblk4[2].pwm.accumulator[1] ;
 wire \genblk4[2].pwm.accumulator[2] ;
 wire \genblk4[2].pwm.accumulator[3] ;
 wire \genblk4[2].pwm.accumulator[4] ;
 wire \genblk4[2].pwm.accumulator[5] ;
 wire \genblk4[2].pwm.accumulator[6] ;
 wire \genblk4[2].pwm.accumulator[7] ;
 wire \genblk4[2].pwm.accumulator[8] ;
 wire \genblk4[2].pwm.accumulator[9] ;
 wire \genblk4[3].pwm.accumulator[0] ;
 wire \genblk4[3].pwm.accumulator[10] ;
 wire \genblk4[3].pwm.accumulator[1] ;
 wire \genblk4[3].pwm.accumulator[2] ;
 wire \genblk4[3].pwm.accumulator[3] ;
 wire \genblk4[3].pwm.accumulator[4] ;
 wire \genblk4[3].pwm.accumulator[5] ;
 wire \genblk4[3].pwm.accumulator[6] ;
 wire \genblk4[3].pwm.accumulator[7] ;
 wire \genblk4[3].pwm.accumulator[8] ;
 wire \genblk4[3].pwm.accumulator[9] ;
 wire \latch_control_reg[0] ;
 wire \latch_control_reg[1] ;
 wire \latch_control_reg[2] ;
 wire \noise[0].gen.counter[0] ;
 wire \noise[0].gen.counter[1] ;
 wire \noise[0].gen.counter[2] ;
 wire \noise[0].gen.counter[3] ;
 wire \noise[0].gen.counter[4] ;
 wire \noise[0].gen.counter[5] ;
 wire \noise[0].gen.counter[6] ;
 wire \noise[0].gen.lfsr[10] ;
 wire \noise[0].gen.lfsr[11] ;
 wire \noise[0].gen.lfsr[12] ;
 wire \noise[0].gen.lfsr[13] ;
 wire \noise[0].gen.lfsr[14] ;
 wire \noise[0].gen.lfsr[1] ;
 wire \noise[0].gen.lfsr[2] ;
 wire \noise[0].gen.lfsr[3] ;
 wire \noise[0].gen.lfsr[4] ;
 wire \noise[0].gen.lfsr[5] ;
 wire \noise[0].gen.lfsr[6] ;
 wire \noise[0].gen.lfsr[7] ;
 wire \noise[0].gen.lfsr[8] ;
 wire \noise[0].gen.lfsr[9] ;
 wire \noise[0].gen.restart_noise ;
 wire \noise[0].gen.signal_edge.previous_signal_state_0 ;
 wire \pwm.accumulator[0] ;
 wire \pwm.accumulator[10] ;
 wire \pwm.accumulator[11] ;
 wire \pwm.accumulator[12] ;
 wire \pwm.accumulator[1] ;
 wire \pwm.accumulator[2] ;
 wire \pwm.accumulator[3] ;
 wire \pwm.accumulator[4] ;
 wire \pwm.accumulator[5] ;
 wire \pwm.accumulator[6] ;
 wire \pwm.accumulator[7] ;
 wire \pwm.accumulator[8] ;
 wire \pwm.accumulator[9] ;
 wire \tone[0].gen.counter[0] ;
 wire \tone[0].gen.counter[1] ;
 wire \tone[0].gen.counter[2] ;
 wire \tone[0].gen.counter[3] ;
 wire \tone[0].gen.counter[4] ;
 wire \tone[0].gen.counter[5] ;
 wire \tone[0].gen.counter[6] ;
 wire \tone[0].gen.counter[7] ;
 wire \tone[0].gen.counter[8] ;
 wire \tone[0].gen.counter[9] ;
 wire \tone[1].gen.counter[0] ;
 wire \tone[1].gen.counter[1] ;
 wire \tone[1].gen.counter[2] ;
 wire \tone[1].gen.counter[3] ;
 wire \tone[1].gen.counter[4] ;
 wire \tone[1].gen.counter[5] ;
 wire \tone[1].gen.counter[6] ;
 wire \tone[1].gen.counter[7] ;
 wire \tone[1].gen.counter[8] ;
 wire \tone[1].gen.counter[9] ;
 wire \tone[2].gen.counter[0] ;
 wire \tone[2].gen.counter[1] ;
 wire \tone[2].gen.counter[2] ;
 wire \tone[2].gen.counter[3] ;
 wire \tone[2].gen.counter[4] ;
 wire \tone[2].gen.counter[5] ;
 wire \tone[2].gen.counter[6] ;
 wire \tone[2].gen.counter[7] ;
 wire \tone[2].gen.counter[8] ;
 wire \tone[2].gen.counter[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_inv_1 _1509_ (.Y(_0811_),
    .A(_0004_));
 sg13g2_buf_1 _1510_ (.A(\chan[2].attenuation.in ),
    .X(_0812_));
 sg13g2_mux4_1 _1511_ (.S0(\control_noise[0][0] ),
    .A0(_0811_),
    .A1(\noise[0].gen.counter[5] ),
    .A2(\noise[0].gen.counter[6] ),
    .A3(net75),
    .S1(\control_noise[0][1] ),
    .X(_0813_));
 sg13g2_nor2b_1 _1512_ (.A(\noise[0].gen.signal_edge.previous_signal_state_0 ),
    .B_N(_0813_),
    .Y(_0814_));
 sg13g2_buf_2 _1513_ (.A(_0814_),
    .X(_0815_));
 sg13g2_buf_1 _1514_ (.A(_0815_),
    .X(_0816_));
 sg13g2_nand2_1 _1515_ (.Y(_0817_),
    .A(\noise[0].gen.lfsr[1] ),
    .B(net29));
 sg13g2_buf_1 _1516_ (.A(\chan[3].attenuation.in ),
    .X(_0818_));
 sg13g2_nand2b_1 _1517_ (.Y(_0819_),
    .B(_0813_),
    .A_N(\noise[0].gen.signal_edge.previous_signal_state_0 ));
 sg13g2_buf_1 _1518_ (.A(_0819_),
    .X(_0820_));
 sg13g2_buf_1 _1519_ (.A(_0820_),
    .X(_0821_));
 sg13g2_nand2_1 _1520_ (.Y(_0822_),
    .A(net74),
    .B(net28));
 sg13g2_buf_1 _1521_ (.A(rst_n),
    .X(_0823_));
 sg13g2_nand2b_1 _1522_ (.Y(_0824_),
    .B(_0823_),
    .A_N(\noise[0].gen.restart_noise ));
 sg13g2_buf_1 _1523_ (.A(_0824_),
    .X(_0825_));
 sg13g2_buf_1 _1524_ (.A(_0825_),
    .X(_0826_));
 sg13g2_a21oi_1 _1525_ (.A1(_0817_),
    .A2(_0822_),
    .Y(_0117_),
    .B1(net38));
 sg13g2_nand2_1 _1526_ (.Y(_0827_),
    .A(\noise[0].gen.lfsr[11] ),
    .B(net29));
 sg13g2_nand2_1 _1527_ (.Y(_0828_),
    .A(\noise[0].gen.lfsr[10] ),
    .B(net28));
 sg13g2_a21oi_1 _1528_ (.A1(_0827_),
    .A2(_0828_),
    .Y(_0118_),
    .B1(net38));
 sg13g2_nand2_1 _1529_ (.Y(_0829_),
    .A(\noise[0].gen.lfsr[12] ),
    .B(_0816_));
 sg13g2_nand2_1 _1530_ (.Y(_0830_),
    .A(\noise[0].gen.lfsr[11] ),
    .B(net28));
 sg13g2_a21oi_1 _1531_ (.A1(_0829_),
    .A2(_0830_),
    .Y(_0119_),
    .B1(net38));
 sg13g2_nand2_1 _1532_ (.Y(_0831_),
    .A(\noise[0].gen.lfsr[13] ),
    .B(_0816_));
 sg13g2_nand2_1 _1533_ (.Y(_0832_),
    .A(\noise[0].gen.lfsr[12] ),
    .B(_0821_));
 sg13g2_a21oi_1 _1534_ (.A1(_0831_),
    .A2(_0832_),
    .Y(_0120_),
    .B1(_0826_));
 sg13g2_nand2_1 _1535_ (.Y(_0833_),
    .A(\noise[0].gen.lfsr[14] ),
    .B(net29));
 sg13g2_nand2_1 _1536_ (.Y(_0834_),
    .A(\noise[0].gen.lfsr[13] ),
    .B(_0821_));
 sg13g2_a21oi_1 _1537_ (.A1(_0833_),
    .A2(_0834_),
    .Y(_0121_),
    .B1(_0826_));
 sg13g2_inv_1 _1538_ (.Y(_0835_),
    .A(_0818_));
 sg13g2_nand2_1 _1539_ (.Y(_0836_),
    .A(\noise[0].gen.lfsr[1] ),
    .B(\control_noise[0][2] ));
 sg13g2_xnor2_1 _1540_ (.Y(_0837_),
    .A(_0835_),
    .B(_0836_));
 sg13g2_nand2_1 _1541_ (.Y(_0838_),
    .A(_0815_),
    .B(_0837_));
 sg13g2_o21ai_1 _1542_ (.B1(_0838_),
    .Y(_0839_),
    .A1(\noise[0].gen.lfsr[14] ),
    .A2(_0815_));
 sg13g2_nand2b_1 _1543_ (.Y(_0122_),
    .B(_0839_),
    .A_N(_0825_));
 sg13g2_nand2_1 _1544_ (.Y(_0840_),
    .A(\noise[0].gen.lfsr[2] ),
    .B(net29));
 sg13g2_nand2_1 _1545_ (.Y(_0841_),
    .A(\noise[0].gen.lfsr[1] ),
    .B(net28));
 sg13g2_a21oi_1 _1546_ (.A1(_0840_),
    .A2(_0841_),
    .Y(_0123_),
    .B1(net38));
 sg13g2_nand2_1 _1547_ (.Y(_0842_),
    .A(\noise[0].gen.lfsr[3] ),
    .B(net29));
 sg13g2_nand2_1 _1548_ (.Y(_0843_),
    .A(\noise[0].gen.lfsr[2] ),
    .B(net28));
 sg13g2_a21oi_1 _1549_ (.A1(_0842_),
    .A2(_0843_),
    .Y(_0124_),
    .B1(net38));
 sg13g2_nand2_1 _1550_ (.Y(_0844_),
    .A(\noise[0].gen.lfsr[4] ),
    .B(net29));
 sg13g2_nand2_1 _1551_ (.Y(_0845_),
    .A(\noise[0].gen.lfsr[3] ),
    .B(net28));
 sg13g2_a21oi_1 _1552_ (.A1(_0844_),
    .A2(_0845_),
    .Y(_0125_),
    .B1(net38));
 sg13g2_nand2_1 _1553_ (.Y(_0846_),
    .A(\noise[0].gen.lfsr[5] ),
    .B(net29));
 sg13g2_nand2_1 _1554_ (.Y(_0847_),
    .A(\noise[0].gen.lfsr[4] ),
    .B(net28));
 sg13g2_a21oi_1 _1555_ (.A1(_0846_),
    .A2(_0847_),
    .Y(_0126_),
    .B1(net38));
 sg13g2_nand2_1 _1556_ (.Y(_0848_),
    .A(\noise[0].gen.lfsr[6] ),
    .B(net29));
 sg13g2_nand2_1 _1557_ (.Y(_0849_),
    .A(\noise[0].gen.lfsr[5] ),
    .B(net28));
 sg13g2_a21oi_1 _1558_ (.A1(_0848_),
    .A2(_0849_),
    .Y(_0127_),
    .B1(net38));
 sg13g2_nand2_1 _1559_ (.Y(_0850_),
    .A(\noise[0].gen.lfsr[7] ),
    .B(_0815_));
 sg13g2_nand2_1 _1560_ (.Y(_0851_),
    .A(\noise[0].gen.lfsr[6] ),
    .B(_0820_));
 sg13g2_a21oi_1 _1561_ (.A1(_0850_),
    .A2(_0851_),
    .Y(_0128_),
    .B1(_0825_));
 sg13g2_nand2_1 _1562_ (.Y(_0852_),
    .A(\noise[0].gen.lfsr[8] ),
    .B(_0815_));
 sg13g2_nand2_1 _1563_ (.Y(_0853_),
    .A(\noise[0].gen.lfsr[7] ),
    .B(_0820_));
 sg13g2_a21oi_1 _1564_ (.A1(_0852_),
    .A2(_0853_),
    .Y(_0129_),
    .B1(_0825_));
 sg13g2_nand2_1 _1565_ (.Y(_0854_),
    .A(\noise[0].gen.lfsr[9] ),
    .B(_0815_));
 sg13g2_nand2_1 _1566_ (.Y(_0855_),
    .A(\noise[0].gen.lfsr[8] ),
    .B(_0820_));
 sg13g2_a21oi_1 _1567_ (.A1(_0854_),
    .A2(_0855_),
    .Y(_0130_),
    .B1(_0825_));
 sg13g2_nand2_1 _1568_ (.Y(_0856_),
    .A(\noise[0].gen.lfsr[10] ),
    .B(_0815_));
 sg13g2_nand2_1 _1569_ (.Y(_0857_),
    .A(\noise[0].gen.lfsr[9] ),
    .B(_0820_));
 sg13g2_a21oi_1 _1570_ (.A1(_0856_),
    .A2(_0857_),
    .Y(_0131_),
    .B1(_0825_));
 sg13g2_inv_1 _1571_ (.Y(_0858_),
    .A(_0823_));
 sg13g2_buf_1 _1572_ (.A(net73),
    .X(_0859_));
 sg13g2_buf_1 _1573_ (.A(net59),
    .X(_0860_));
 sg13g2_buf_2 _1574_ (.A(ui_in[5]),
    .X(_0861_));
 sg13g2_buf_2 _1575_ (.A(ui_in[4]),
    .X(_0862_));
 sg13g2_buf_2 _1576_ (.A(uio_in[0]),
    .X(_0863_));
 sg13g2_nand2b_1 _1577_ (.Y(_0864_),
    .B(net5),
    .A_N(_0863_));
 sg13g2_buf_2 _1578_ (.A(_0864_),
    .X(_0865_));
 sg13g2_nor2_1 _1579_ (.A(_0862_),
    .B(_0865_),
    .Y(_0866_));
 sg13g2_nand3_1 _1580_ (.B(net4),
    .C(_0866_),
    .A(_0861_),
    .Y(_0867_));
 sg13g2_buf_1 _1581_ (.A(_0867_),
    .X(_0868_));
 sg13g2_nor2_1 _1582_ (.A(net37),
    .B(_0868_),
    .Y(_0146_));
 sg13g2_buf_1 _1583_ (.A(_0823_),
    .X(_0869_));
 sg13g2_and2_1 _1584_ (.A(_0869_),
    .B(_0005_),
    .X(_0007_));
 sg13g2_xnor2_1 _1585_ (.Y(_0870_),
    .A(\clk_counter[1] ),
    .B(\clk_counter[0] ));
 sg13g2_nor2_1 _1586_ (.A(net37),
    .B(_0870_),
    .Y(_0008_));
 sg13g2_nand2_1 _1587_ (.Y(_0871_),
    .A(\clk_counter[1] ),
    .B(\clk_counter[0] ));
 sg13g2_xor2_1 _1588_ (.B(_0871_),
    .A(\clk_counter[2] ),
    .X(_0872_));
 sg13g2_nor2_1 _1589_ (.A(net37),
    .B(_0872_),
    .Y(_0009_));
 sg13g2_inv_1 _1590_ (.Y(_0873_),
    .A(\clk_counter[3] ));
 sg13g2_nand3_1 _1591_ (.B(\clk_counter[0] ),
    .C(\clk_counter[2] ),
    .A(\clk_counter[1] ),
    .Y(_0874_));
 sg13g2_xnor2_1 _1592_ (.Y(_0875_),
    .A(_0873_),
    .B(_0874_));
 sg13g2_nor2_1 _1593_ (.A(net37),
    .B(_0875_),
    .Y(_0010_));
 sg13g2_nor2_1 _1594_ (.A(_0873_),
    .B(_0874_),
    .Y(_0876_));
 sg13g2_xnor2_1 _1595_ (.Y(_0877_),
    .A(\clk_counter[4] ),
    .B(_0876_));
 sg13g2_nor2_1 _1596_ (.A(net37),
    .B(_0877_),
    .Y(_0011_));
 sg13g2_nand2_1 _1597_ (.Y(_0878_),
    .A(\clk_counter[4] ),
    .B(_0876_));
 sg13g2_xor2_1 _1598_ (.B(_0878_),
    .A(\clk_counter[5] ),
    .X(_0879_));
 sg13g2_nor2_1 _1599_ (.A(_0860_),
    .B(_0879_),
    .Y(_0012_));
 sg13g2_nand3_1 _1600_ (.B(\clk_counter[4] ),
    .C(_0876_),
    .A(\clk_counter[5] ),
    .Y(_0880_));
 sg13g2_xor2_1 _1601_ (.B(_0880_),
    .A(\clk_counter[6] ),
    .X(_0881_));
 sg13g2_nor2_1 _1602_ (.A(_0860_),
    .B(_0881_),
    .Y(_0013_));
 sg13g2_buf_1 _1603_ (.A(_0823_),
    .X(_0882_));
 sg13g2_buf_1 _1604_ (.A(_0863_),
    .X(_0883_));
 sg13g2_nor2b_2 _1605_ (.A(net5),
    .B_N(\latch_control_reg[0] ),
    .Y(_0884_));
 sg13g2_buf_1 _1606_ (.A(\latch_control_reg[1] ),
    .X(_0885_));
 sg13g2_nor2_1 _1607_ (.A(_0885_),
    .B(\latch_control_reg[2] ),
    .Y(_0886_));
 sg13g2_and2_1 _1608_ (.A(net5),
    .B(_0862_),
    .X(_0887_));
 sg13g2_buf_1 _1609_ (.A(_0887_),
    .X(_0888_));
 sg13g2_nor2_1 _1610_ (.A(_0861_),
    .B(net4),
    .Y(_0889_));
 sg13g2_a22oi_1 _1611_ (.Y(_0890_),
    .B1(_0888_),
    .B2(_0889_),
    .A2(_0886_),
    .A1(_0884_));
 sg13g2_buf_1 _1612_ (.A(_0890_),
    .X(_0891_));
 sg13g2_buf_1 _1613_ (.A(\chan[0].attenuation.control[0] ),
    .X(_0892_));
 sg13g2_o21ai_1 _1614_ (.B1(_0892_),
    .Y(_0893_),
    .A1(net70),
    .A2(_0891_));
 sg13g2_buf_1 _1615_ (.A(net1),
    .X(_0894_));
 sg13g2_nor2_1 _1616_ (.A(net70),
    .B(_0891_),
    .Y(_0895_));
 sg13g2_nand2_1 _1617_ (.Y(_0896_),
    .A(net79),
    .B(_0895_));
 sg13g2_nand3_1 _1618_ (.B(_0893_),
    .C(_0896_),
    .A(net71),
    .Y(_0014_));
 sg13g2_buf_8 _1619_ (.A(\chan[0].attenuation.control[1] ),
    .X(_0897_));
 sg13g2_o21ai_1 _1620_ (.B1(_0897_),
    .Y(_0898_),
    .A1(net70),
    .A2(_0891_));
 sg13g2_buf_1 _1621_ (.A(net2),
    .X(_0899_));
 sg13g2_nand2_1 _1622_ (.Y(_0900_),
    .A(net78),
    .B(_0895_));
 sg13g2_nand3_1 _1623_ (.B(_0898_),
    .C(_0900_),
    .A(net71),
    .Y(_0015_));
 sg13g2_buf_8 _1624_ (.A(\chan[0].attenuation.control[2] ),
    .X(_0901_));
 sg13g2_buf_8 _1625_ (.A(_0901_),
    .X(_0902_));
 sg13g2_o21ai_1 _1626_ (.B1(_0902_),
    .Y(_0903_),
    .A1(_0883_),
    .A2(_0891_));
 sg13g2_buf_1 _1627_ (.A(net3),
    .X(_0904_));
 sg13g2_nand2_1 _1628_ (.Y(_0905_),
    .A(net77),
    .B(_0895_));
 sg13g2_nand3_1 _1629_ (.B(_0903_),
    .C(_0905_),
    .A(_0882_),
    .Y(_0016_));
 sg13g2_buf_8 _1630_ (.A(\chan[0].attenuation.control[3] ),
    .X(_0906_));
 sg13g2_buf_1 _1631_ (.A(_0906_),
    .X(_0907_));
 sg13g2_o21ai_1 _1632_ (.B1(_0907_),
    .Y(_0908_),
    .A1(_0883_),
    .A2(_0891_));
 sg13g2_buf_1 _1633_ (.A(ui_in[3]),
    .X(_0909_));
 sg13g2_nand2_1 _1634_ (.Y(_0910_),
    .A(net76),
    .B(_0895_));
 sg13g2_nand3_1 _1635_ (.B(_0908_),
    .C(_0910_),
    .A(_0882_),
    .Y(_0017_));
 sg13g2_nand3b_1 _1636_ (.B(_0884_),
    .C(_0885_),
    .Y(_0911_),
    .A_N(\latch_control_reg[2] ));
 sg13g2_inv_1 _1637_ (.Y(_0912_),
    .A(net4));
 sg13g2_nand3_1 _1638_ (.B(_0912_),
    .C(_0888_),
    .A(_0861_),
    .Y(_0913_));
 sg13g2_a21oi_2 _1639_ (.B1(_0863_),
    .Y(_0914_),
    .A2(_0913_),
    .A1(_0911_));
 sg13g2_buf_2 _1640_ (.A(\chan[1].attenuation.control[0] ),
    .X(_0915_));
 sg13g2_buf_1 _1641_ (.A(_0915_),
    .X(_0916_));
 sg13g2_nand2b_1 _1642_ (.Y(_0917_),
    .B(_0916_),
    .A_N(_0914_));
 sg13g2_nand2_1 _1643_ (.Y(_0918_),
    .A(net79),
    .B(_0914_));
 sg13g2_nand3_1 _1644_ (.B(_0917_),
    .C(_0918_),
    .A(net71),
    .Y(_0018_));
 sg13g2_buf_2 _1645_ (.A(\chan[1].attenuation.control[1] ),
    .X(_0919_));
 sg13g2_buf_1 _1646_ (.A(_0919_),
    .X(_0920_));
 sg13g2_nand2b_1 _1647_ (.Y(_0921_),
    .B(_0920_),
    .A_N(_0914_));
 sg13g2_nand2_1 _1648_ (.Y(_0922_),
    .A(net78),
    .B(_0914_));
 sg13g2_nand3_1 _1649_ (.B(_0921_),
    .C(_0922_),
    .A(net71),
    .Y(_0019_));
 sg13g2_buf_1 _1650_ (.A(\chan[1].attenuation.control[2] ),
    .X(_0923_));
 sg13g2_buf_1 _1651_ (.A(_0923_),
    .X(_0924_));
 sg13g2_nand2b_1 _1652_ (.Y(_0925_),
    .B(_0924_),
    .A_N(_0914_));
 sg13g2_nand2_1 _1653_ (.Y(_0926_),
    .A(net77),
    .B(_0914_));
 sg13g2_nand3_1 _1654_ (.B(_0925_),
    .C(_0926_),
    .A(net71),
    .Y(_0020_));
 sg13g2_buf_1 _1655_ (.A(\chan[1].attenuation.control[3] ),
    .X(_0927_));
 sg13g2_nand2b_1 _1656_ (.Y(_0928_),
    .B(net67),
    .A_N(_0914_));
 sg13g2_nand2_1 _1657_ (.Y(_0929_),
    .A(net76),
    .B(_0914_));
 sg13g2_nand3_1 _1658_ (.B(_0928_),
    .C(_0929_),
    .A(net71),
    .Y(_0021_));
 sg13g2_nor2_1 _1659_ (.A(_0861_),
    .B(_0912_),
    .Y(_0930_));
 sg13g2_nor2_1 _1660_ (.A(_0885_),
    .B(_0003_),
    .Y(_0931_));
 sg13g2_a22oi_1 _1661_ (.Y(_0932_),
    .B1(_0931_),
    .B2(_0884_),
    .A2(_0930_),
    .A1(_0888_));
 sg13g2_buf_1 _1662_ (.A(_0932_),
    .X(_0933_));
 sg13g2_buf_8 _1663_ (.A(\chan[2].attenuation.control[0] ),
    .X(_0934_));
 sg13g2_buf_1 _1664_ (.A(_0934_),
    .X(_0935_));
 sg13g2_o21ai_1 _1665_ (.B1(_0935_),
    .Y(_0936_),
    .A1(net70),
    .A2(_0933_));
 sg13g2_nor2_1 _1666_ (.A(net70),
    .B(_0933_),
    .Y(_0937_));
 sg13g2_nand2_1 _1667_ (.Y(_0938_),
    .A(_0894_),
    .B(_0937_));
 sg13g2_nand3_1 _1668_ (.B(_0936_),
    .C(_0938_),
    .A(net71),
    .Y(_0022_));
 sg13g2_buf_1 _1669_ (.A(_0823_),
    .X(_0939_));
 sg13g2_buf_1 _1670_ (.A(\chan[2].attenuation.control[1] ),
    .X(_0940_));
 sg13g2_buf_1 _1671_ (.A(_0940_),
    .X(_0941_));
 sg13g2_o21ai_1 _1672_ (.B1(_0941_),
    .Y(_0942_),
    .A1(net70),
    .A2(_0933_));
 sg13g2_nand2_1 _1673_ (.Y(_0943_),
    .A(net78),
    .B(_0937_));
 sg13g2_nand3_1 _1674_ (.B(_0942_),
    .C(_0943_),
    .A(net66),
    .Y(_0023_));
 sg13g2_buf_1 _1675_ (.A(\chan[2].attenuation.control[2] ),
    .X(_0944_));
 sg13g2_buf_1 _1676_ (.A(net65),
    .X(_0945_));
 sg13g2_o21ai_1 _1677_ (.B1(_0945_),
    .Y(_0946_),
    .A1(net70),
    .A2(_0933_));
 sg13g2_nand2_1 _1678_ (.Y(_0947_),
    .A(_0904_),
    .B(_0937_));
 sg13g2_nand3_1 _1679_ (.B(_0946_),
    .C(_0947_),
    .A(net66),
    .Y(_0024_));
 sg13g2_buf_2 _1680_ (.A(\chan[2].attenuation.control[3] ),
    .X(_0948_));
 sg13g2_buf_8 _1681_ (.A(_0948_),
    .X(_0949_));
 sg13g2_o21ai_1 _1682_ (.B1(_0949_),
    .Y(_0950_),
    .A1(net70),
    .A2(_0933_));
 sg13g2_nand2_1 _1683_ (.Y(_0951_),
    .A(net76),
    .B(_0937_));
 sg13g2_nand3_1 _1684_ (.B(_0950_),
    .C(_0951_),
    .A(net66),
    .Y(_0025_));
 sg13g2_nand3_1 _1685_ (.B(net4),
    .C(_0888_),
    .A(_0861_),
    .Y(_0952_));
 sg13g2_nand3b_1 _1686_ (.B(_0884_),
    .C(_0885_),
    .Y(_0953_),
    .A_N(_0003_));
 sg13g2_a21oi_2 _1687_ (.B1(_0863_),
    .Y(_0954_),
    .A2(_0953_),
    .A1(_0952_));
 sg13g2_buf_1 _1688_ (.A(\chan[3].attenuation.control[0] ),
    .X(_0955_));
 sg13g2_nand2b_1 _1689_ (.Y(_0956_),
    .B(_0955_),
    .A_N(_0954_));
 sg13g2_nand2_1 _1690_ (.Y(_0957_),
    .A(net79),
    .B(_0954_));
 sg13g2_nand3_1 _1691_ (.B(_0956_),
    .C(_0957_),
    .A(net66),
    .Y(_0026_));
 sg13g2_buf_2 _1692_ (.A(\chan[3].attenuation.control[1] ),
    .X(_0958_));
 sg13g2_buf_1 _1693_ (.A(_0958_),
    .X(_0959_));
 sg13g2_nand2b_1 _1694_ (.Y(_0960_),
    .B(_0959_),
    .A_N(_0954_));
 sg13g2_nand2_1 _1695_ (.Y(_0961_),
    .A(net78),
    .B(_0954_));
 sg13g2_nand3_1 _1696_ (.B(_0960_),
    .C(_0961_),
    .A(net66),
    .Y(_0027_));
 sg13g2_buf_2 _1697_ (.A(\chan[3].attenuation.control[2] ),
    .X(_0962_));
 sg13g2_buf_1 _1698_ (.A(_0962_),
    .X(_0963_));
 sg13g2_nand2b_1 _1699_ (.Y(_0964_),
    .B(_0963_),
    .A_N(_0954_));
 sg13g2_nand2_1 _1700_ (.Y(_0965_),
    .A(net77),
    .B(_0954_));
 sg13g2_nand3_1 _1701_ (.B(_0964_),
    .C(_0965_),
    .A(net66),
    .Y(_0028_));
 sg13g2_buf_2 _1702_ (.A(\chan[3].attenuation.control[3] ),
    .X(_0966_));
 sg13g2_buf_1 _1703_ (.A(_0966_),
    .X(_0967_));
 sg13g2_nand2b_1 _1704_ (.Y(_0968_),
    .B(_0967_),
    .A_N(_0954_));
 sg13g2_nand2_1 _1705_ (.Y(_0969_),
    .A(net76),
    .B(_0954_));
 sg13g2_nand3_1 _1706_ (.B(_0968_),
    .C(_0969_),
    .A(net66),
    .Y(_0029_));
 sg13g2_mux2_1 _1707_ (.A0(net79),
    .A1(\control_noise[0][0] ),
    .S(_0868_),
    .X(_0970_));
 sg13g2_and2_1 _1708_ (.A(net72),
    .B(_0970_),
    .X(_0030_));
 sg13g2_mux2_1 _1709_ (.A0(net78),
    .A1(\control_noise[0][1] ),
    .S(_0868_),
    .X(_0971_));
 sg13g2_and2_1 _1710_ (.A(net72),
    .B(_0971_),
    .X(_0031_));
 sg13g2_nor2_1 _1711_ (.A(net77),
    .B(_0868_),
    .Y(_0972_));
 sg13g2_nor2b_1 _1712_ (.A(\control_noise[0][2] ),
    .B_N(_0868_),
    .Y(_0973_));
 sg13g2_o21ai_1 _1713_ (.B1(net71),
    .Y(_0032_),
    .A1(_0972_),
    .A2(_0973_));
 sg13g2_and2_1 _1714_ (.A(_0866_),
    .B(_0889_),
    .X(_0974_));
 sg13g2_buf_2 _1715_ (.A(_0974_),
    .X(_0975_));
 sg13g2_nand2b_1 _1716_ (.Y(_0976_),
    .B(\control_tone_freq[0][0] ),
    .A_N(_0975_));
 sg13g2_nand2_1 _1717_ (.Y(_0977_),
    .A(net79),
    .B(_0975_));
 sg13g2_nand3_1 _1718_ (.B(_0976_),
    .C(_0977_),
    .A(net66),
    .Y(_0033_));
 sg13g2_nand2_1 _1719_ (.Y(_0978_),
    .A(net78),
    .B(_0975_));
 sg13g2_nand2b_1 _1720_ (.Y(_0979_),
    .B(\control_tone_freq[0][1] ),
    .A_N(_0975_));
 sg13g2_buf_1 _1721_ (.A(net73),
    .X(_0980_));
 sg13g2_a21oi_1 _1722_ (.A1(_0978_),
    .A2(_0979_),
    .Y(_0034_),
    .B1(net46));
 sg13g2_nand2_1 _1723_ (.Y(_0981_),
    .A(net77),
    .B(_0975_));
 sg13g2_nand2b_1 _1724_ (.Y(_0982_),
    .B(\control_tone_freq[0][2] ),
    .A_N(_0975_));
 sg13g2_a21oi_1 _1725_ (.A1(_0981_),
    .A2(_0982_),
    .Y(_0035_),
    .B1(net46));
 sg13g2_nand2_1 _1726_ (.Y(_0983_),
    .A(net76),
    .B(_0975_));
 sg13g2_nand2b_1 _1727_ (.Y(_0984_),
    .B(\control_tone_freq[0][3] ),
    .A_N(_0975_));
 sg13g2_buf_1 _1728_ (.A(net73),
    .X(_0985_));
 sg13g2_a21oi_1 _1729_ (.A1(_0983_),
    .A2(_0984_),
    .Y(_0036_),
    .B1(net45));
 sg13g2_nor3_2 _1730_ (.A(net5),
    .B(_0863_),
    .C(\latch_control_reg[0] ),
    .Y(_0986_));
 sg13g2_and2_1 _1731_ (.A(_0886_),
    .B(_0986_),
    .X(_0987_));
 sg13g2_buf_1 _1732_ (.A(_0987_),
    .X(_0988_));
 sg13g2_nand2_1 _1733_ (.Y(_0989_),
    .A(net79),
    .B(net35));
 sg13g2_nand2b_1 _1734_ (.Y(_0990_),
    .B(\control_tone_freq[0][4] ),
    .A_N(net35));
 sg13g2_a21oi_1 _1735_ (.A1(_0989_),
    .A2(_0990_),
    .Y(_0037_),
    .B1(net45));
 sg13g2_nand2_1 _1736_ (.Y(_0991_),
    .A(_0899_),
    .B(net35));
 sg13g2_nand2b_1 _1737_ (.Y(_0992_),
    .B(\control_tone_freq[0][5] ),
    .A_N(net35));
 sg13g2_a21oi_1 _1738_ (.A1(_0991_),
    .A2(_0992_),
    .Y(_0038_),
    .B1(net45));
 sg13g2_nand2_1 _1739_ (.Y(_0993_),
    .A(net77),
    .B(net35));
 sg13g2_nand2b_1 _1740_ (.Y(_0994_),
    .B(\control_tone_freq[0][6] ),
    .A_N(net35));
 sg13g2_a21oi_1 _1741_ (.A1(_0993_),
    .A2(_0994_),
    .Y(_0039_),
    .B1(net45));
 sg13g2_nand2_1 _1742_ (.Y(_0995_),
    .A(net76),
    .B(net35));
 sg13g2_nand2b_1 _1743_ (.Y(_0996_),
    .B(\control_tone_freq[0][7] ),
    .A_N(net35));
 sg13g2_a21oi_1 _1744_ (.A1(_0995_),
    .A2(_0996_),
    .Y(_0040_),
    .B1(net45));
 sg13g2_nand2_1 _1745_ (.Y(_0997_),
    .A(_0862_),
    .B(_0988_));
 sg13g2_nand2b_1 _1746_ (.Y(_0998_),
    .B(\control_tone_freq[0][8] ),
    .A_N(_0987_));
 sg13g2_a21oi_1 _1747_ (.A1(_0997_),
    .A2(_0998_),
    .Y(_0041_),
    .B1(_0985_));
 sg13g2_nand2_1 _1748_ (.Y(_0999_),
    .A(_0861_),
    .B(_0988_));
 sg13g2_nand2b_1 _1749_ (.Y(_1000_),
    .B(\control_tone_freq[0][9] ),
    .A_N(_0987_));
 sg13g2_a21oi_1 _1750_ (.A1(_0999_),
    .A2(_1000_),
    .Y(_0042_),
    .B1(_0985_));
 sg13g2_inv_1 _1751_ (.Y(_1001_),
    .A(_0861_));
 sg13g2_nor4_2 _1752_ (.A(_1001_),
    .B(_0862_),
    .C(net4),
    .Y(_1002_),
    .D(_0865_));
 sg13g2_nand2b_1 _1753_ (.Y(_1003_),
    .B(\control_tone_freq[1][0] ),
    .A_N(_1002_));
 sg13g2_nand2_1 _1754_ (.Y(_1004_),
    .A(net79),
    .B(_1002_));
 sg13g2_nand3_1 _1755_ (.B(_1003_),
    .C(_1004_),
    .A(_0939_),
    .Y(_0043_));
 sg13g2_nand2_1 _1756_ (.Y(_1005_),
    .A(net78),
    .B(_1002_));
 sg13g2_nand2b_1 _1757_ (.Y(_1006_),
    .B(\control_tone_freq[1][1] ),
    .A_N(_1002_));
 sg13g2_a21oi_1 _1758_ (.A1(_1005_),
    .A2(_1006_),
    .Y(_0044_),
    .B1(net45));
 sg13g2_nand2_1 _1759_ (.Y(_1007_),
    .A(net77),
    .B(_1002_));
 sg13g2_nand2b_1 _1760_ (.Y(_1008_),
    .B(\control_tone_freq[1][2] ),
    .A_N(_1002_));
 sg13g2_a21oi_1 _1761_ (.A1(_1007_),
    .A2(_1008_),
    .Y(_0045_),
    .B1(net45));
 sg13g2_nand2_1 _1762_ (.Y(_1009_),
    .A(net76),
    .B(_1002_));
 sg13g2_nand2b_1 _1763_ (.Y(_1010_),
    .B(\control_tone_freq[1][3] ),
    .A_N(_1002_));
 sg13g2_a21oi_1 _1764_ (.A1(_1009_),
    .A2(_1010_),
    .Y(_0046_),
    .B1(net45));
 sg13g2_nor2b_1 _1765_ (.A(\latch_control_reg[2] ),
    .B_N(_0986_),
    .Y(_1011_));
 sg13g2_nand2_2 _1766_ (.Y(_1012_),
    .A(_0885_),
    .B(_1011_));
 sg13g2_mux2_1 _1767_ (.A0(net79),
    .A1(\control_tone_freq[1][4] ),
    .S(_1012_),
    .X(_1013_));
 sg13g2_and2_1 _1768_ (.A(net72),
    .B(_1013_),
    .X(_0047_));
 sg13g2_mux2_1 _1769_ (.A0(net78),
    .A1(\control_tone_freq[1][5] ),
    .S(_1012_),
    .X(_1014_));
 sg13g2_and2_1 _1770_ (.A(net72),
    .B(_1014_),
    .X(_0048_));
 sg13g2_mux2_1 _1771_ (.A0(net77),
    .A1(\control_tone_freq[1][6] ),
    .S(_1012_),
    .X(_1015_));
 sg13g2_and2_1 _1772_ (.A(net72),
    .B(_1015_),
    .X(_0049_));
 sg13g2_mux2_1 _1773_ (.A0(net76),
    .A1(\control_tone_freq[1][7] ),
    .S(_1012_),
    .X(_1016_));
 sg13g2_and2_1 _1774_ (.A(net72),
    .B(_1016_),
    .X(_0050_));
 sg13g2_mux2_1 _1775_ (.A0(_0862_),
    .A1(\control_tone_freq[1][8] ),
    .S(_1012_),
    .X(_1017_));
 sg13g2_and2_1 _1776_ (.A(net72),
    .B(_1017_),
    .X(_0051_));
 sg13g2_nand2_1 _1777_ (.Y(_1018_),
    .A(\control_tone_freq[1][9] ),
    .B(_1012_));
 sg13g2_o21ai_1 _1778_ (.B1(_1018_),
    .Y(_1019_),
    .A1(_1001_),
    .A2(_1012_));
 sg13g2_and2_1 _1779_ (.A(net72),
    .B(_1019_),
    .X(_0052_));
 sg13g2_and2_1 _1780_ (.A(_0866_),
    .B(_0930_),
    .X(_1020_));
 sg13g2_buf_2 _1781_ (.A(_1020_),
    .X(_1021_));
 sg13g2_nand2b_1 _1782_ (.Y(_1022_),
    .B(\control_tone_freq[2][0] ),
    .A_N(_1021_));
 sg13g2_nand2_1 _1783_ (.Y(_1023_),
    .A(_0894_),
    .B(_1021_));
 sg13g2_nand3_1 _1784_ (.B(_1022_),
    .C(_1023_),
    .A(_0939_),
    .Y(_0053_));
 sg13g2_nand2_1 _1785_ (.Y(_1024_),
    .A(_0899_),
    .B(_1021_));
 sg13g2_nand2b_1 _1786_ (.Y(_1025_),
    .B(\control_tone_freq[2][1] ),
    .A_N(_1021_));
 sg13g2_buf_1 _1787_ (.A(_0858_),
    .X(_1026_));
 sg13g2_a21oi_1 _1788_ (.A1(_1024_),
    .A2(_1025_),
    .Y(_0054_),
    .B1(net44));
 sg13g2_nand2_1 _1789_ (.Y(_1027_),
    .A(_0904_),
    .B(_1021_));
 sg13g2_nand2b_1 _1790_ (.Y(_1028_),
    .B(\control_tone_freq[2][2] ),
    .A_N(_1021_));
 sg13g2_a21oi_1 _1791_ (.A1(_1027_),
    .A2(_1028_),
    .Y(_0055_),
    .B1(net44));
 sg13g2_nand2_1 _1792_ (.Y(_1029_),
    .A(_0909_),
    .B(_1021_));
 sg13g2_nand2b_1 _1793_ (.Y(_1030_),
    .B(\control_tone_freq[2][3] ),
    .A_N(_1021_));
 sg13g2_a21oi_1 _1794_ (.A1(_1029_),
    .A2(_1030_),
    .Y(_0056_),
    .B1(net44));
 sg13g2_nand2_2 _1795_ (.Y(_1031_),
    .A(_0931_),
    .B(_0986_));
 sg13g2_mux2_1 _1796_ (.A0(net1),
    .A1(\control_tone_freq[2][4] ),
    .S(_1031_),
    .X(_1032_));
 sg13g2_and2_1 _1797_ (.A(_0869_),
    .B(_1032_),
    .X(_0057_));
 sg13g2_buf_1 _1798_ (.A(_0823_),
    .X(_1033_));
 sg13g2_mux2_1 _1799_ (.A0(net2),
    .A1(\control_tone_freq[2][5] ),
    .S(_1031_),
    .X(_1034_));
 sg13g2_and2_1 _1800_ (.A(net63),
    .B(_1034_),
    .X(_0058_));
 sg13g2_mux2_1 _1801_ (.A0(net3),
    .A1(\control_tone_freq[2][6] ),
    .S(_1031_),
    .X(_1035_));
 sg13g2_and2_1 _1802_ (.A(net63),
    .B(_1035_),
    .X(_0059_));
 sg13g2_mux2_1 _1803_ (.A0(_0909_),
    .A1(\control_tone_freq[2][7] ),
    .S(_1031_),
    .X(_1036_));
 sg13g2_and2_1 _1804_ (.A(net63),
    .B(_1036_),
    .X(_0060_));
 sg13g2_mux2_1 _1805_ (.A0(_0862_),
    .A1(\control_tone_freq[2][8] ),
    .S(_1031_),
    .X(_1037_));
 sg13g2_and2_1 _1806_ (.A(_1033_),
    .B(_1037_),
    .X(_0061_));
 sg13g2_nand2_1 _1807_ (.Y(_1038_),
    .A(\control_tone_freq[2][9] ),
    .B(_1031_));
 sg13g2_o21ai_1 _1808_ (.B1(_1038_),
    .Y(_1039_),
    .A1(_1001_),
    .A2(_1031_));
 sg13g2_and2_1 _1809_ (.A(_1033_),
    .B(_1039_),
    .X(_0062_));
 sg13g2_buf_1 _1810_ (.A(\chan[0].attenuation.in ),
    .X(_1040_));
 sg13g2_nand2_1 _1811_ (.Y(_1041_),
    .A(_0897_),
    .B(_0907_));
 sg13g2_nand3b_1 _1812_ (.B(_1041_),
    .C(_0892_),
    .Y(_1042_),
    .A_N(_0902_));
 sg13g2_nor2b_1 _1813_ (.A(\chan[0].attenuation.control[0] ),
    .B_N(_0906_),
    .Y(_1043_));
 sg13g2_a21oi_1 _1814_ (.A1(net58),
    .A2(net68),
    .Y(_1044_),
    .B1(_1043_));
 sg13g2_and3_1 _1815_ (.X(_1045_),
    .A(net62),
    .B(_1042_),
    .C(_1044_));
 sg13g2_xnor2_1 _1816_ (.Y(_1046_),
    .A(\genblk4[0].pwm.accumulator[0] ),
    .B(_1045_));
 sg13g2_nor2_1 _1817_ (.A(net37),
    .B(_1046_),
    .Y(_0063_));
 sg13g2_xor2_1 _1818_ (.B(_0906_),
    .A(net58),
    .X(_1047_));
 sg13g2_nor3_1 _1819_ (.A(net69),
    .B(net68),
    .C(_1047_),
    .Y(_1048_));
 sg13g2_nand2b_1 _1820_ (.Y(_1049_),
    .B(net68),
    .A_N(net58));
 sg13g2_a21oi_1 _1821_ (.A1(net69),
    .A2(net58),
    .Y(_1050_),
    .B1(net57));
 sg13g2_a21oi_1 _1822_ (.A1(net57),
    .A2(_1049_),
    .Y(_1051_),
    .B1(_1050_));
 sg13g2_o21ai_1 _1823_ (.B1(net62),
    .Y(_1052_),
    .A1(_1048_),
    .A2(_1051_));
 sg13g2_buf_1 _1824_ (.A(_1052_),
    .X(_1053_));
 sg13g2_inv_2 _1825_ (.Y(_1054_),
    .A(net62));
 sg13g2_mux2_1 _1826_ (.A0(\chan[0].attenuation.control[1] ),
    .A1(_0901_),
    .S(_0906_),
    .X(_1055_));
 sg13g2_nand2b_1 _1827_ (.Y(_1056_),
    .B(_0901_),
    .A_N(\chan[0].attenuation.control[1] ));
 sg13g2_mux2_1 _1828_ (.A0(_1055_),
    .A1(_1056_),
    .S(\chan[0].attenuation.control[0] ),
    .X(_1057_));
 sg13g2_inv_1 _1829_ (.Y(_1058_),
    .A(\genblk4[0].pwm.accumulator[1] ));
 sg13g2_o21ai_1 _1830_ (.B1(_1058_),
    .Y(_1059_),
    .A1(_1054_),
    .A2(_1057_));
 sg13g2_and4_1 _1831_ (.A(net62),
    .B(\genblk4[0].pwm.accumulator[0] ),
    .C(_1042_),
    .D(_1044_),
    .X(_1060_));
 sg13g2_nor2_1 _1832_ (.A(_0901_),
    .B(net68),
    .Y(_1061_));
 sg13g2_and3_1 _1833_ (.X(_1062_),
    .A(\chan[0].attenuation.control[0] ),
    .B(_0901_),
    .C(\chan[0].attenuation.control[1] ));
 sg13g2_inv_1 _1834_ (.Y(_1063_),
    .A(_0906_));
 sg13g2_o21ai_1 _1835_ (.B1(_1063_),
    .Y(_1064_),
    .A1(_1061_),
    .A2(_1062_));
 sg13g2_or2_1 _1836_ (.X(_1065_),
    .B(_0906_),
    .A(\chan[0].attenuation.control[1] ));
 sg13g2_a21o_1 _1837_ (.A2(_1065_),
    .A1(_1049_),
    .B1(net69),
    .X(_1066_));
 sg13g2_a21oi_2 _1838_ (.B1(_1054_),
    .Y(_1067_),
    .A2(_1066_),
    .A1(_1064_));
 sg13g2_nor3_1 _1839_ (.A(_1054_),
    .B(_1058_),
    .C(_1057_),
    .Y(_1068_));
 sg13g2_a221oi_1 _1840_ (.B2(\genblk4[0].pwm.accumulator[2] ),
    .C1(_1068_),
    .B1(_1067_),
    .A1(_1059_),
    .Y(_1069_),
    .A2(_1060_));
 sg13g2_nor2_1 _1841_ (.A(\genblk4[0].pwm.accumulator[2] ),
    .B(_1067_),
    .Y(_1070_));
 sg13g2_nand2_1 _1842_ (.Y(_1071_),
    .A(net58),
    .B(net68));
 sg13g2_nand2b_1 _1843_ (.Y(_1072_),
    .B(_1043_),
    .A_N(_1071_));
 sg13g2_a21o_1 _1844_ (.A2(_1072_),
    .A1(_1064_),
    .B1(_1054_),
    .X(_1073_));
 sg13g2_buf_2 _1845_ (.A(_1073_),
    .X(_1074_));
 sg13g2_o21ai_1 _1846_ (.B1(_1074_),
    .Y(_1075_),
    .A1(_1069_),
    .A2(_1070_));
 sg13g2_nor3_1 _1847_ (.A(_1074_),
    .B(_1069_),
    .C(_1070_),
    .Y(_1076_));
 sg13g2_a21oi_2 _1848_ (.B1(_1076_),
    .Y(_1077_),
    .A2(_1075_),
    .A1(\genblk4[0].pwm.accumulator[3] ));
 sg13g2_nor2_1 _1849_ (.A(net69),
    .B(_1065_),
    .Y(_1078_));
 sg13g2_xor2_1 _1850_ (.B(net68),
    .A(_0901_),
    .X(_1079_));
 sg13g2_and3_1 _1851_ (.X(_1080_),
    .A(net69),
    .B(net57),
    .C(_1079_));
 sg13g2_o21ai_1 _1852_ (.B1(net62),
    .Y(_1081_),
    .A1(_1078_),
    .A2(_1080_));
 sg13g2_buf_1 _1853_ (.A(_1081_),
    .X(_1082_));
 sg13g2_nor2_1 _1854_ (.A(_1077_),
    .B(_1082_),
    .Y(_1083_));
 sg13g2_inv_1 _1855_ (.Y(_1084_),
    .A(\genblk4[0].pwm.accumulator[4] ));
 sg13g2_a21oi_1 _1856_ (.A1(_1077_),
    .A2(_1082_),
    .Y(_1085_),
    .B1(_1084_));
 sg13g2_or2_1 _1857_ (.X(_1086_),
    .B(_1085_),
    .A(_1083_));
 sg13g2_xor2_1 _1858_ (.B(_1056_),
    .A(net69),
    .X(_1087_));
 sg13g2_nor3_1 _1859_ (.A(net58),
    .B(net68),
    .C(net57),
    .Y(_1088_));
 sg13g2_a21oi_1 _1860_ (.A1(net57),
    .A2(_1087_),
    .Y(_1089_),
    .B1(_1088_));
 sg13g2_nor2_2 _1861_ (.A(_1054_),
    .B(_1089_),
    .Y(_1090_));
 sg13g2_a21o_1 _1862_ (.A2(_1090_),
    .A1(_1086_),
    .B1(\genblk4[0].pwm.accumulator[5] ),
    .X(_1091_));
 sg13g2_o21ai_1 _1863_ (.B1(_1091_),
    .Y(_1092_),
    .A1(_1086_),
    .A2(_1090_));
 sg13g2_nand2_1 _1864_ (.Y(_1093_),
    .A(_1053_),
    .B(_1092_));
 sg13g2_inv_1 _1865_ (.Y(_1094_),
    .A(\genblk4[0].pwm.accumulator[6] ));
 sg13g2_o21ai_1 _1866_ (.B1(_1094_),
    .Y(_1095_),
    .A1(_1053_),
    .A2(_1092_));
 sg13g2_nand2_1 _1867_ (.Y(_1096_),
    .A(_1093_),
    .B(_1095_));
 sg13g2_xnor2_1 _1868_ (.Y(_1097_),
    .A(net69),
    .B(_1071_));
 sg13g2_nand2_1 _1869_ (.Y(_1098_),
    .A(net57),
    .B(_1061_));
 sg13g2_o21ai_1 _1870_ (.B1(_1098_),
    .Y(_1099_),
    .A1(net57),
    .A2(_1097_));
 sg13g2_nand2_2 _1871_ (.Y(_1100_),
    .A(net62),
    .B(_1099_));
 sg13g2_nand2_1 _1872_ (.Y(_1101_),
    .A(_1096_),
    .B(_1100_));
 sg13g2_nor2_1 _1873_ (.A(_1096_),
    .B(_1100_),
    .Y(_1102_));
 sg13g2_a21oi_2 _1874_ (.B1(_1102_),
    .Y(_1103_),
    .A2(_1101_),
    .A1(\genblk4[0].pwm.accumulator[7] ));
 sg13g2_nand2b_1 _1875_ (.Y(_1104_),
    .B(net58),
    .A_N(net69));
 sg13g2_nand2b_1 _1876_ (.Y(_1105_),
    .B(net62),
    .A_N(net57));
 sg13g2_a21oi_2 _1877_ (.B1(_1105_),
    .Y(_1106_),
    .A2(_1104_),
    .A1(net68));
 sg13g2_inv_1 _1878_ (.Y(_1107_),
    .A(_1106_));
 sg13g2_nor2_1 _1879_ (.A(_1103_),
    .B(_1107_),
    .Y(_1108_));
 sg13g2_nand2_1 _1880_ (.Y(_1109_),
    .A(_1103_),
    .B(_1107_));
 sg13g2_o21ai_1 _1881_ (.B1(_1109_),
    .Y(_1110_),
    .A1(\genblk4[0].pwm.accumulator[8] ),
    .A2(_1108_));
 sg13g2_nor2_2 _1882_ (.A(net58),
    .B(_1105_),
    .Y(_1111_));
 sg13g2_nor2_1 _1883_ (.A(\genblk4[0].pwm.accumulator[9] ),
    .B(_1111_),
    .Y(_1112_));
 sg13g2_nand2_1 _1884_ (.Y(_1113_),
    .A(\genblk4[0].pwm.accumulator[9] ),
    .B(_1111_));
 sg13g2_o21ai_1 _1885_ (.B1(_1113_),
    .Y(_1114_),
    .A1(_1110_),
    .A2(_1112_));
 sg13g2_and2_1 _1886_ (.A(net63),
    .B(_1114_),
    .X(_0064_));
 sg13g2_nor2_2 _1887_ (.A(_1054_),
    .B(_1057_),
    .Y(_1115_));
 sg13g2_xnor2_1 _1888_ (.Y(_1116_),
    .A(_1115_),
    .B(_1060_));
 sg13g2_xnor2_1 _1889_ (.Y(_1117_),
    .A(_1058_),
    .B(_1116_));
 sg13g2_nor2_1 _1890_ (.A(net37),
    .B(_1117_),
    .Y(_0065_));
 sg13g2_nand2_1 _1891_ (.Y(_1118_),
    .A(\genblk4[0].pwm.accumulator[1] ),
    .B(_1115_));
 sg13g2_nand2_1 _1892_ (.Y(_1119_),
    .A(_1059_),
    .B(_1060_));
 sg13g2_xnor2_1 _1893_ (.Y(_1120_),
    .A(\genblk4[0].pwm.accumulator[2] ),
    .B(_1067_));
 sg13g2_and3_1 _1894_ (.X(_1121_),
    .A(_1118_),
    .B(_1119_),
    .C(_1120_));
 sg13g2_a21oi_1 _1895_ (.A1(_1118_),
    .A2(_1119_),
    .Y(_1122_),
    .B1(_1120_));
 sg13g2_nor3_1 _1896_ (.A(net59),
    .B(_1121_),
    .C(_1122_),
    .Y(_0066_));
 sg13g2_nor2_1 _1897_ (.A(_1069_),
    .B(_1070_),
    .Y(_1123_));
 sg13g2_xnor2_1 _1898_ (.Y(_1124_),
    .A(\genblk4[0].pwm.accumulator[3] ),
    .B(_1074_));
 sg13g2_xnor2_1 _1899_ (.Y(_1125_),
    .A(_1123_),
    .B(_1124_));
 sg13g2_nor2_1 _1900_ (.A(net37),
    .B(_1125_),
    .Y(_0067_));
 sg13g2_buf_1 _1901_ (.A(net59),
    .X(_1126_));
 sg13g2_xnor2_1 _1902_ (.Y(_1127_),
    .A(_1084_),
    .B(_1082_));
 sg13g2_xnor2_1 _1903_ (.Y(_1128_),
    .A(_1077_),
    .B(_1127_));
 sg13g2_nor2_1 _1904_ (.A(_1126_),
    .B(_1128_),
    .Y(_0068_));
 sg13g2_xnor2_1 _1905_ (.Y(_1129_),
    .A(\genblk4[0].pwm.accumulator[5] ),
    .B(_1090_));
 sg13g2_xnor2_1 _1906_ (.Y(_1130_),
    .A(_1086_),
    .B(_1129_));
 sg13g2_and2_1 _1907_ (.A(net63),
    .B(_1130_),
    .X(_0069_));
 sg13g2_xnor2_1 _1908_ (.Y(_1131_),
    .A(_1094_),
    .B(_1053_));
 sg13g2_xnor2_1 _1909_ (.Y(_1132_),
    .A(_1092_),
    .B(_1131_));
 sg13g2_nor2_1 _1910_ (.A(net36),
    .B(_1132_),
    .Y(_0070_));
 sg13g2_xor2_1 _1911_ (.B(_1100_),
    .A(\genblk4[0].pwm.accumulator[7] ),
    .X(_1133_));
 sg13g2_xnor2_1 _1912_ (.Y(_1134_),
    .A(_1096_),
    .B(_1133_));
 sg13g2_nor2_1 _1913_ (.A(net36),
    .B(_1134_),
    .Y(_0071_));
 sg13g2_xnor2_1 _1914_ (.Y(_1135_),
    .A(\genblk4[0].pwm.accumulator[8] ),
    .B(_1106_));
 sg13g2_xnor2_1 _1915_ (.Y(_1136_),
    .A(_1103_),
    .B(_1135_));
 sg13g2_nor2_1 _1916_ (.A(_1126_),
    .B(_1136_),
    .Y(_0072_));
 sg13g2_xnor2_1 _1917_ (.Y(_1137_),
    .A(\genblk4[0].pwm.accumulator[9] ),
    .B(_1111_));
 sg13g2_xnor2_1 _1918_ (.Y(_1138_),
    .A(_1110_),
    .B(_1137_));
 sg13g2_nor2_1 _1919_ (.A(net36),
    .B(_1138_),
    .Y(_0073_));
 sg13g2_nor2b_1 _1920_ (.A(net67),
    .B_N(net56),
    .Y(_1139_));
 sg13g2_o21ai_1 _1921_ (.B1(net55),
    .Y(_1140_),
    .A1(net54),
    .A2(_1139_));
 sg13g2_inv_1 _1922_ (.Y(_1141_),
    .A(net56));
 sg13g2_inv_1 _1923_ (.Y(_1142_),
    .A(\chan[1].attenuation.in ));
 sg13g2_a21oi_1 _1924_ (.A1(_1141_),
    .A2(net67),
    .Y(_1143_),
    .B1(_1142_));
 sg13g2_nor2_1 _1925_ (.A(_0919_),
    .B(_0923_),
    .Y(_1144_));
 sg13g2_nand2_1 _1926_ (.Y(_1145_),
    .A(net56),
    .B(_1144_));
 sg13g2_and3_1 _1927_ (.X(_1146_),
    .A(_1140_),
    .B(_1143_),
    .C(_1145_));
 sg13g2_xnor2_1 _1928_ (.Y(_1147_),
    .A(\genblk4[1].pwm.accumulator[0] ),
    .B(_1146_));
 sg13g2_nor2_1 _1929_ (.A(net36),
    .B(_1147_),
    .Y(_0074_));
 sg13g2_buf_1 _1930_ (.A(\chan[1].attenuation.in ),
    .X(_1148_));
 sg13g2_inv_2 _1931_ (.Y(_1149_),
    .A(_0927_));
 sg13g2_nand2_1 _1932_ (.Y(_1150_),
    .A(net61),
    .B(_1149_));
 sg13g2_nor2_2 _1933_ (.A(net54),
    .B(_1150_),
    .Y(_1151_));
 sg13g2_or2_1 _1934_ (.X(_1152_),
    .B(_0923_),
    .A(_0915_));
 sg13g2_nand3_1 _1935_ (.B(net56),
    .C(net54),
    .A(net55),
    .Y(_1153_));
 sg13g2_a21oi_1 _1936_ (.A1(_1152_),
    .A2(_1153_),
    .Y(_1154_),
    .B1(net67));
 sg13g2_nand2b_1 _1937_ (.Y(_1155_),
    .B(net67),
    .A_N(net54));
 sg13g2_or2_1 _1938_ (.X(_1156_),
    .B(\chan[1].attenuation.control[3] ),
    .A(_0915_));
 sg13g2_a21oi_1 _1939_ (.A1(_1155_),
    .A2(_1156_),
    .Y(_1157_),
    .B1(net55));
 sg13g2_o21ai_1 _1940_ (.B1(net61),
    .Y(_1158_),
    .A1(_1154_),
    .A2(_1157_));
 sg13g2_buf_2 _1941_ (.A(_1158_),
    .X(_1159_));
 sg13g2_xor2_1 _1942_ (.B(net67),
    .A(net54),
    .X(_1160_));
 sg13g2_nor3_1 _1943_ (.A(net55),
    .B(net56),
    .C(_1160_),
    .Y(_1161_));
 sg13g2_nand3b_1 _1944_ (.B(_0923_),
    .C(_0915_),
    .Y(_1162_),
    .A_N(\chan[1].attenuation.control[3] ));
 sg13g2_nand3b_1 _1945_ (.B(net67),
    .C(_0919_),
    .Y(_1163_),
    .A_N(net54));
 sg13g2_nand2_1 _1946_ (.Y(_1164_),
    .A(_1162_),
    .B(_1163_));
 sg13g2_o21ai_1 _1947_ (.B1(net61),
    .Y(_1165_),
    .A1(_1161_),
    .A2(_1164_));
 sg13g2_buf_2 _1948_ (.A(_1165_),
    .X(_1166_));
 sg13g2_xor2_1 _1949_ (.B(\chan[1].attenuation.control[3] ),
    .A(_0915_),
    .X(_1167_));
 sg13g2_and2_1 _1950_ (.A(_0919_),
    .B(_0923_),
    .X(_1168_));
 sg13g2_a22oi_1 _1951_ (.Y(_1169_),
    .B1(_1167_),
    .B2(_1168_),
    .A2(_1144_),
    .A1(_1149_));
 sg13g2_nand2b_1 _1952_ (.Y(_1170_),
    .B(net61),
    .A_N(_1169_));
 sg13g2_buf_2 _1953_ (.A(_1170_),
    .X(_1171_));
 sg13g2_nand2_1 _1954_ (.Y(_1172_),
    .A(_0915_),
    .B(_0923_));
 sg13g2_a21o_1 _1955_ (.A2(_1172_),
    .A1(_1149_),
    .B1(_0919_),
    .X(_1173_));
 sg13g2_nand3_1 _1956_ (.B(_1152_),
    .C(_1162_),
    .A(net55),
    .Y(_1174_));
 sg13g2_nand3_1 _1957_ (.B(_1173_),
    .C(_1174_),
    .A(net61),
    .Y(_1175_));
 sg13g2_nand2b_1 _1958_ (.Y(_1176_),
    .B(net61),
    .A_N(_0919_));
 sg13g2_a21o_1 _1959_ (.A2(_1156_),
    .A1(_1172_),
    .B1(_1176_),
    .X(_1177_));
 sg13g2_or3_1 _1960_ (.A(_1142_),
    .B(_1149_),
    .C(_1152_),
    .X(_1178_));
 sg13g2_nand2_2 _1961_ (.Y(_1179_),
    .A(_1177_),
    .B(_1178_));
 sg13g2_and4_1 _1962_ (.A(\genblk4[1].pwm.accumulator[0] ),
    .B(_1140_),
    .C(_1143_),
    .D(_1145_),
    .X(_1180_));
 sg13g2_nand2_1 _1963_ (.Y(_1181_),
    .A(_1179_),
    .B(_1180_));
 sg13g2_o21ai_1 _1964_ (.B1(\genblk4[1].pwm.accumulator[1] ),
    .Y(_1182_),
    .A1(_1179_),
    .A2(_1180_));
 sg13g2_nand3_1 _1965_ (.B(_1181_),
    .C(_1182_),
    .A(_1175_),
    .Y(_1183_));
 sg13g2_a21oi_1 _1966_ (.A1(_1181_),
    .A2(_1182_),
    .Y(_1184_),
    .B1(_1175_));
 sg13g2_a21oi_1 _1967_ (.A1(\genblk4[1].pwm.accumulator[2] ),
    .A2(_1183_),
    .Y(_1185_),
    .B1(_1184_));
 sg13g2_or2_1 _1968_ (.X(_1186_),
    .B(_1185_),
    .A(_1171_));
 sg13g2_inv_1 _1969_ (.Y(_1187_),
    .A(\genblk4[1].pwm.accumulator[3] ));
 sg13g2_a21o_1 _1970_ (.A2(_1185_),
    .A1(_1171_),
    .B1(_1187_),
    .X(_1188_));
 sg13g2_nand3_1 _1971_ (.B(net54),
    .C(net67),
    .A(net56),
    .Y(_1189_));
 sg13g2_a21oi_1 _1972_ (.A1(_1156_),
    .A2(_1189_),
    .Y(_1190_),
    .B1(net55));
 sg13g2_nor2_1 _1973_ (.A(_1141_),
    .B(_1163_),
    .Y(_1191_));
 sg13g2_o21ai_1 _1974_ (.B1(net61),
    .Y(_1192_),
    .A1(_1190_),
    .A2(_1191_));
 sg13g2_buf_2 _1975_ (.A(_1192_),
    .X(_1193_));
 sg13g2_a21oi_1 _1976_ (.A1(_1186_),
    .A2(_1188_),
    .Y(_1194_),
    .B1(_1193_));
 sg13g2_nand3_1 _1977_ (.B(_1188_),
    .C(_1193_),
    .A(_1186_),
    .Y(_1195_));
 sg13g2_o21ai_1 _1978_ (.B1(_1195_),
    .Y(_1196_),
    .A1(\genblk4[1].pwm.accumulator[4] ),
    .A2(_1194_));
 sg13g2_nand2b_1 _1979_ (.Y(_1197_),
    .B(net55),
    .A_N(_0916_));
 sg13g2_nand3b_1 _1980_ (.B(net56),
    .C(_0924_),
    .Y(_1198_),
    .A_N(_0920_));
 sg13g2_a21oi_1 _1981_ (.A1(_1197_),
    .A2(_1198_),
    .Y(_1199_),
    .B1(_1149_));
 sg13g2_nand2_1 _1982_ (.Y(_1200_),
    .A(net56),
    .B(_0927_));
 sg13g2_and2_1 _1983_ (.A(_1144_),
    .B(_1200_),
    .X(_1201_));
 sg13g2_o21ai_1 _1984_ (.B1(_1148_),
    .Y(_1202_),
    .A1(_1199_),
    .A2(_1201_));
 sg13g2_buf_2 _1985_ (.A(_1202_),
    .X(_1203_));
 sg13g2_nand2_1 _1986_ (.Y(_1204_),
    .A(_1196_),
    .B(_1203_));
 sg13g2_nor2_1 _1987_ (.A(_1196_),
    .B(_1203_),
    .Y(_1205_));
 sg13g2_a21oi_2 _1988_ (.B1(_1205_),
    .Y(_1206_),
    .A2(_1204_),
    .A1(\genblk4[1].pwm.accumulator[5] ));
 sg13g2_nand2_1 _1989_ (.Y(_1207_),
    .A(_1166_),
    .B(_1206_));
 sg13g2_nor2_1 _1990_ (.A(_1166_),
    .B(_1206_),
    .Y(_1208_));
 sg13g2_a21oi_2 _1991_ (.B1(_1208_),
    .Y(_1209_),
    .A2(_1207_),
    .A1(\genblk4[1].pwm.accumulator[6] ));
 sg13g2_nand2_1 _1992_ (.Y(_1210_),
    .A(_1159_),
    .B(_1209_));
 sg13g2_nor2_1 _1993_ (.A(_1159_),
    .B(_1209_),
    .Y(_1211_));
 sg13g2_a21oi_1 _1994_ (.A1(\genblk4[1].pwm.accumulator[7] ),
    .A2(_1210_),
    .Y(_1212_),
    .B1(_1211_));
 sg13g2_nand2_1 _1995_ (.Y(_1213_),
    .A(_1141_),
    .B(net54));
 sg13g2_a21oi_2 _1996_ (.B1(_1150_),
    .Y(_1214_),
    .A2(_1213_),
    .A1(net55));
 sg13g2_nor2_1 _1997_ (.A(\genblk4[1].pwm.accumulator[8] ),
    .B(_1214_),
    .Y(_1215_));
 sg13g2_nand2_1 _1998_ (.Y(_1216_),
    .A(\genblk4[1].pwm.accumulator[8] ),
    .B(_1214_));
 sg13g2_o21ai_1 _1999_ (.B1(_1216_),
    .Y(_1217_),
    .A1(_1212_),
    .A2(_1215_));
 sg13g2_o21ai_1 _2000_ (.B1(_1217_),
    .Y(_1218_),
    .A1(\genblk4[1].pwm.accumulator[9] ),
    .A2(_1151_));
 sg13g2_nand2_1 _2001_ (.Y(_1219_),
    .A(\genblk4[1].pwm.accumulator[9] ),
    .B(_1151_));
 sg13g2_a21oi_1 _2002_ (.A1(_1218_),
    .A2(_1219_),
    .Y(_0075_),
    .B1(net44));
 sg13g2_xnor2_1 _2003_ (.Y(_1220_),
    .A(_1179_),
    .B(_1180_));
 sg13g2_xor2_1 _2004_ (.B(_1220_),
    .A(\genblk4[1].pwm.accumulator[1] ),
    .X(_1221_));
 sg13g2_nor2_1 _2005_ (.A(net36),
    .B(_1221_),
    .Y(_0076_));
 sg13g2_and3_1 _2006_ (.X(_1222_),
    .A(net61),
    .B(_1173_),
    .C(_1174_));
 sg13g2_buf_2 _2007_ (.A(_1222_),
    .X(_1223_));
 sg13g2_xnor2_1 _2008_ (.Y(_1224_),
    .A(\genblk4[1].pwm.accumulator[2] ),
    .B(_1223_));
 sg13g2_and3_1 _2009_ (.X(_1225_),
    .A(_1181_),
    .B(_1182_),
    .C(_1224_));
 sg13g2_a21oi_1 _2010_ (.A1(_1181_),
    .A2(_1182_),
    .Y(_1226_),
    .B1(_1224_));
 sg13g2_nor3_1 _2011_ (.A(net59),
    .B(_1225_),
    .C(_1226_),
    .Y(_0077_));
 sg13g2_xnor2_1 _2012_ (.Y(_1227_),
    .A(_1187_),
    .B(_1171_));
 sg13g2_xnor2_1 _2013_ (.Y(_1228_),
    .A(_1185_),
    .B(_1227_));
 sg13g2_nor2_1 _2014_ (.A(net36),
    .B(_1228_),
    .Y(_0078_));
 sg13g2_nand2_1 _2015_ (.Y(_1229_),
    .A(_1186_),
    .B(_1188_));
 sg13g2_xnor2_1 _2016_ (.Y(_1230_),
    .A(\genblk4[1].pwm.accumulator[4] ),
    .B(_1193_));
 sg13g2_xnor2_1 _2017_ (.Y(_1231_),
    .A(_1229_),
    .B(_1230_));
 sg13g2_nor2_1 _2018_ (.A(net36),
    .B(_1231_),
    .Y(_0079_));
 sg13g2_xor2_1 _2019_ (.B(_1203_),
    .A(\genblk4[1].pwm.accumulator[5] ),
    .X(_1232_));
 sg13g2_xnor2_1 _2020_ (.Y(_1233_),
    .A(_1196_),
    .B(_1232_));
 sg13g2_nor2_1 _2021_ (.A(net36),
    .B(_1233_),
    .Y(_0080_));
 sg13g2_buf_1 _2022_ (.A(net73),
    .X(_1234_));
 sg13g2_xor2_1 _2023_ (.B(_1166_),
    .A(\genblk4[1].pwm.accumulator[6] ),
    .X(_1235_));
 sg13g2_xnor2_1 _2024_ (.Y(_1236_),
    .A(_1206_),
    .B(_1235_));
 sg13g2_nor2_1 _2025_ (.A(net43),
    .B(_1236_),
    .Y(_0081_));
 sg13g2_xor2_1 _2026_ (.B(_1159_),
    .A(\genblk4[1].pwm.accumulator[7] ),
    .X(_1237_));
 sg13g2_xnor2_1 _2027_ (.Y(_1238_),
    .A(_1209_),
    .B(_1237_));
 sg13g2_nor2_1 _2028_ (.A(net43),
    .B(_1238_),
    .Y(_0082_));
 sg13g2_xnor2_1 _2029_ (.Y(_1239_),
    .A(\genblk4[1].pwm.accumulator[8] ),
    .B(_1214_));
 sg13g2_xnor2_1 _2030_ (.Y(_1240_),
    .A(_1212_),
    .B(_1239_));
 sg13g2_nor2_1 _2031_ (.A(net43),
    .B(_1240_),
    .Y(_0083_));
 sg13g2_xor2_1 _2032_ (.B(_1151_),
    .A(\genblk4[1].pwm.accumulator[9] ),
    .X(_1241_));
 sg13g2_xnor2_1 _2033_ (.Y(_1242_),
    .A(_1217_),
    .B(_1241_));
 sg13g2_nor2_1 _2034_ (.A(_1234_),
    .B(_1242_),
    .Y(_0084_));
 sg13g2_inv_2 _2035_ (.Y(_1243_),
    .A(_0948_));
 sg13g2_nand3b_1 _2036_ (.B(_1243_),
    .C(_0935_),
    .Y(_1244_),
    .A_N(net51));
 sg13g2_inv_2 _2037_ (.Y(_1245_),
    .A(net75));
 sg13g2_a21oi_1 _2038_ (.A1(_0941_),
    .A2(net51),
    .Y(_1246_),
    .B1(_1245_));
 sg13g2_o21ai_1 _2039_ (.B1(net53),
    .Y(_1247_),
    .A1(net52),
    .A2(_0945_));
 sg13g2_nand2_1 _2040_ (.Y(_1248_),
    .A(_0949_),
    .B(_1247_));
 sg13g2_and3_1 _2041_ (.X(_1249_),
    .A(_1244_),
    .B(_1246_),
    .C(_1248_));
 sg13g2_buf_1 _2042_ (.A(_1249_),
    .X(_1250_));
 sg13g2_xnor2_1 _2043_ (.Y(_1251_),
    .A(\genblk4[2].pwm.accumulator[0] ),
    .B(_1250_));
 sg13g2_nor2_1 _2044_ (.A(_1234_),
    .B(_1251_),
    .Y(_0085_));
 sg13g2_nand2_1 _2045_ (.Y(_1252_),
    .A(net75),
    .B(_1243_));
 sg13g2_nor2_2 _2046_ (.A(net51),
    .B(_1252_),
    .Y(_1253_));
 sg13g2_nor2_1 _2047_ (.A(\genblk4[2].pwm.accumulator[9] ),
    .B(_1253_),
    .Y(_1254_));
 sg13g2_nand2b_1 _2048_ (.Y(_1255_),
    .B(net65),
    .A_N(net53));
 sg13g2_a21oi_2 _2049_ (.B1(_1252_),
    .Y(_1256_),
    .A2(_1255_),
    .A1(net52));
 sg13g2_inv_1 _2050_ (.Y(_1257_),
    .A(\genblk4[2].pwm.accumulator[8] ));
 sg13g2_mux2_1 _2051_ (.A0(net53),
    .A1(net51),
    .S(net50),
    .X(_1258_));
 sg13g2_nor2_1 _2052_ (.A(net52),
    .B(_1258_),
    .Y(_1259_));
 sg13g2_or2_1 _2053_ (.X(_1260_),
    .B(net65),
    .A(_0934_));
 sg13g2_nand3_1 _2054_ (.B(net53),
    .C(net51),
    .A(net52),
    .Y(_1261_));
 sg13g2_a21oi_1 _2055_ (.A1(_1260_),
    .A2(_1261_),
    .Y(_1262_),
    .B1(net50));
 sg13g2_o21ai_1 _2056_ (.B1(net75),
    .Y(_1263_),
    .A1(_1259_),
    .A2(_1262_));
 sg13g2_buf_2 _2057_ (.A(_1263_),
    .X(_1264_));
 sg13g2_inv_1 _2058_ (.Y(_1265_),
    .A(_0940_));
 sg13g2_mux2_1 _2059_ (.A0(net51),
    .A1(_1255_),
    .S(_1265_),
    .X(_1266_));
 sg13g2_nor3_1 _2060_ (.A(net52),
    .B(net53),
    .C(net51),
    .Y(_1267_));
 sg13g2_a21o_1 _2061_ (.A2(net65),
    .A1(_0934_),
    .B1(net50),
    .X(_1268_));
 sg13g2_o21ai_1 _2062_ (.B1(net75),
    .Y(_1269_),
    .A1(_1267_),
    .A2(_1268_));
 sg13g2_a21o_1 _2063_ (.A2(_1266_),
    .A1(net50),
    .B1(_1269_),
    .X(_1270_));
 sg13g2_buf_2 _2064_ (.A(_1270_),
    .X(_1271_));
 sg13g2_nor2b_1 _2065_ (.A(net52),
    .B_N(net65),
    .Y(_1272_));
 sg13g2_nor3_1 _2066_ (.A(net53),
    .B(_1243_),
    .C(_1272_),
    .Y(_1273_));
 sg13g2_or2_1 _2067_ (.X(_1274_),
    .B(net50),
    .A(net65));
 sg13g2_nand3_1 _2068_ (.B(net65),
    .C(net50),
    .A(net53),
    .Y(_1275_));
 sg13g2_a21oi_1 _2069_ (.A1(_1274_),
    .A2(_1275_),
    .Y(_1276_),
    .B1(net52));
 sg13g2_o21ai_1 _2070_ (.B1(net75),
    .Y(_1277_),
    .A1(_1273_),
    .A2(_1276_));
 sg13g2_buf_2 _2071_ (.A(_1277_),
    .X(_1278_));
 sg13g2_inv_1 _2072_ (.Y(_1279_),
    .A(\genblk4[2].pwm.accumulator[4] ));
 sg13g2_nand2b_1 _2073_ (.Y(_1280_),
    .B(_1265_),
    .A_N(_1268_));
 sg13g2_nand3b_1 _2074_ (.B(_0944_),
    .C(_0934_),
    .Y(_1281_),
    .A_N(_0948_));
 sg13g2_a21o_1 _2075_ (.A2(_1281_),
    .A1(_1260_),
    .B1(_1265_),
    .X(_1282_));
 sg13g2_a21o_1 _2076_ (.A2(_1282_),
    .A1(_1280_),
    .B1(_1245_),
    .X(_1283_));
 sg13g2_buf_2 _2077_ (.A(_1283_),
    .X(_1284_));
 sg13g2_nor2_1 _2078_ (.A(_0934_),
    .B(_0948_),
    .Y(_1285_));
 sg13g2_and2_1 _2079_ (.A(_0934_),
    .B(net65),
    .X(_1286_));
 sg13g2_nor2b_1 _2080_ (.A(_0940_),
    .B_N(net75),
    .Y(_1287_));
 sg13g2_o21ai_1 _2081_ (.B1(_1287_),
    .Y(_1288_),
    .A1(_1285_),
    .A2(_1286_));
 sg13g2_or3_1 _2082_ (.A(_1245_),
    .B(_1243_),
    .C(_1260_),
    .X(_1289_));
 sg13g2_nand2_2 _2083_ (.Y(_1290_),
    .A(_1288_),
    .B(_1289_));
 sg13g2_and4_1 _2084_ (.A(\genblk4[2].pwm.accumulator[0] ),
    .B(_1244_),
    .C(_1246_),
    .D(_1248_),
    .X(_1291_));
 sg13g2_nand2_1 _2085_ (.Y(_1292_),
    .A(_1290_),
    .B(_1291_));
 sg13g2_o21ai_1 _2086_ (.B1(\genblk4[2].pwm.accumulator[1] ),
    .Y(_1293_),
    .A1(_1290_),
    .A2(_1291_));
 sg13g2_nand3_1 _2087_ (.B(_1292_),
    .C(_1293_),
    .A(_1284_),
    .Y(_1294_));
 sg13g2_a21oi_1 _2088_ (.A1(_1292_),
    .A2(_1293_),
    .Y(_1295_),
    .B1(_1284_));
 sg13g2_a21oi_2 _2089_ (.B1(_1295_),
    .Y(_1296_),
    .A2(_1294_),
    .A1(\genblk4[2].pwm.accumulator[2] ));
 sg13g2_and3_1 _2090_ (.X(_1297_),
    .A(_0940_),
    .B(_0934_),
    .C(\chan[2].attenuation.control[2] ));
 sg13g2_and2_1 _2091_ (.A(_0940_),
    .B(_0948_),
    .X(_1298_));
 sg13g2_nor2b_1 _2092_ (.A(_0934_),
    .B_N(\chan[2].attenuation.control[2] ),
    .Y(_1299_));
 sg13g2_nor3_1 _2093_ (.A(_0940_),
    .B(_0944_),
    .C(_0948_),
    .Y(_1300_));
 sg13g2_a221oi_1 _2094_ (.B2(_1299_),
    .C1(_1300_),
    .B1(_1298_),
    .A1(_1243_),
    .Y(_1301_),
    .A2(_1297_));
 sg13g2_or2_1 _2095_ (.X(_1302_),
    .B(_1301_),
    .A(_1245_));
 sg13g2_buf_8 _2096_ (.A(_1302_),
    .X(_1303_));
 sg13g2_nor2_1 _2097_ (.A(_1296_),
    .B(_1303_),
    .Y(_1304_));
 sg13g2_inv_1 _2098_ (.Y(_1305_),
    .A(\genblk4[2].pwm.accumulator[3] ));
 sg13g2_a21oi_1 _2099_ (.A1(_1296_),
    .A2(_1303_),
    .Y(_1306_),
    .B1(_1305_));
 sg13g2_xor2_1 _2100_ (.B(net51),
    .A(net52),
    .X(_1307_));
 sg13g2_and2_1 _2101_ (.A(net53),
    .B(net50),
    .X(_1308_));
 sg13g2_a22oi_1 _2102_ (.Y(_1309_),
    .B1(_1307_),
    .B2(_1308_),
    .A2(_1285_),
    .A1(_1265_));
 sg13g2_nor2_2 _2103_ (.A(_1245_),
    .B(_1309_),
    .Y(_1310_));
 sg13g2_o21ai_1 _2104_ (.B1(_1310_),
    .Y(_1311_),
    .A1(_1304_),
    .A2(_1306_));
 sg13g2_nor3_1 _2105_ (.A(_1310_),
    .B(_1304_),
    .C(_1306_),
    .Y(_1312_));
 sg13g2_a21o_1 _2106_ (.A2(_1311_),
    .A1(_1279_),
    .B1(_1312_),
    .X(_1313_));
 sg13g2_or2_1 _2107_ (.X(_1314_),
    .B(_1313_),
    .A(_1278_));
 sg13g2_inv_1 _2108_ (.Y(_1315_),
    .A(\genblk4[2].pwm.accumulator[5] ));
 sg13g2_a21o_1 _2109_ (.A2(_1313_),
    .A1(_1278_),
    .B1(_1315_),
    .X(_1316_));
 sg13g2_nand3_1 _2110_ (.B(_1314_),
    .C(_1316_),
    .A(_1271_),
    .Y(_1317_));
 sg13g2_a21oi_1 _2111_ (.A1(_1314_),
    .A2(_1316_),
    .Y(_1318_),
    .B1(_1271_));
 sg13g2_a21oi_2 _2112_ (.B1(_1318_),
    .Y(_1319_),
    .A2(_1317_),
    .A1(\genblk4[2].pwm.accumulator[6] ));
 sg13g2_nand2_1 _2113_ (.Y(_1320_),
    .A(_1264_),
    .B(_1319_));
 sg13g2_nor2_1 _2114_ (.A(_1264_),
    .B(_1319_),
    .Y(_1321_));
 sg13g2_a21oi_2 _2115_ (.B1(_1321_),
    .Y(_1322_),
    .A2(_1320_),
    .A1(\genblk4[2].pwm.accumulator[7] ));
 sg13g2_nand2_1 _2116_ (.Y(_1323_),
    .A(_1257_),
    .B(_1322_));
 sg13g2_nor2_1 _2117_ (.A(_1257_),
    .B(_1322_),
    .Y(_1324_));
 sg13g2_a21oi_1 _2118_ (.A1(_1256_),
    .A2(_1323_),
    .Y(_1325_),
    .B1(_1324_));
 sg13g2_nand2_1 _2119_ (.Y(_1326_),
    .A(\genblk4[2].pwm.accumulator[9] ),
    .B(_1253_));
 sg13g2_o21ai_1 _2120_ (.B1(_1326_),
    .Y(_1327_),
    .A1(_1254_),
    .A2(_1325_));
 sg13g2_and2_1 _2121_ (.A(net63),
    .B(_1327_),
    .X(_0086_));
 sg13g2_xnor2_1 _2122_ (.Y(_1328_),
    .A(_1290_),
    .B(_1291_));
 sg13g2_xor2_1 _2123_ (.B(_1328_),
    .A(\genblk4[2].pwm.accumulator[1] ),
    .X(_1329_));
 sg13g2_nor2_1 _2124_ (.A(net43),
    .B(_1329_),
    .Y(_0087_));
 sg13g2_nand2_1 _2125_ (.Y(_1330_),
    .A(_1292_),
    .B(_1293_));
 sg13g2_xnor2_1 _2126_ (.Y(_1331_),
    .A(\genblk4[2].pwm.accumulator[2] ),
    .B(_1284_));
 sg13g2_xnor2_1 _2127_ (.Y(_1332_),
    .A(_1330_),
    .B(_1331_));
 sg13g2_nor2_1 _2128_ (.A(net43),
    .B(_1332_),
    .Y(_0088_));
 sg13g2_xnor2_1 _2129_ (.Y(_1333_),
    .A(_1305_),
    .B(_1303_));
 sg13g2_xnor2_1 _2130_ (.Y(_1334_),
    .A(_1296_),
    .B(_1333_));
 sg13g2_nor2_1 _2131_ (.A(net43),
    .B(_1334_),
    .Y(_0089_));
 sg13g2_nor2_1 _2132_ (.A(_1304_),
    .B(_1306_),
    .Y(_1335_));
 sg13g2_xnor2_1 _2133_ (.Y(_1336_),
    .A(\genblk4[2].pwm.accumulator[4] ),
    .B(_1310_));
 sg13g2_xnor2_1 _2134_ (.Y(_1337_),
    .A(_1335_),
    .B(_1336_));
 sg13g2_nor2_1 _2135_ (.A(net43),
    .B(_1337_),
    .Y(_0090_));
 sg13g2_xnor2_1 _2136_ (.Y(_1338_),
    .A(_1315_),
    .B(_1278_));
 sg13g2_xnor2_1 _2137_ (.Y(_1339_),
    .A(_1313_),
    .B(_1338_));
 sg13g2_nor2_1 _2138_ (.A(net43),
    .B(_1339_),
    .Y(_0091_));
 sg13g2_buf_1 _2139_ (.A(net73),
    .X(_1340_));
 sg13g2_nand2_1 _2140_ (.Y(_0180_),
    .A(_1314_),
    .B(_1316_));
 sg13g2_xnor2_1 _2141_ (.Y(_0181_),
    .A(\genblk4[2].pwm.accumulator[6] ),
    .B(_1271_));
 sg13g2_xnor2_1 _2142_ (.Y(_0182_),
    .A(_0180_),
    .B(_0181_));
 sg13g2_nor2_1 _2143_ (.A(_1340_),
    .B(_0182_),
    .Y(_0092_));
 sg13g2_xor2_1 _2144_ (.B(_1264_),
    .A(\genblk4[2].pwm.accumulator[7] ),
    .X(_0183_));
 sg13g2_xnor2_1 _2145_ (.Y(_0184_),
    .A(_1319_),
    .B(_0183_));
 sg13g2_nor2_1 _2146_ (.A(_1340_),
    .B(_0184_),
    .Y(_0093_));
 sg13g2_xnor2_1 _2147_ (.Y(_0185_),
    .A(\genblk4[2].pwm.accumulator[8] ),
    .B(_1256_));
 sg13g2_xnor2_1 _2148_ (.Y(_0186_),
    .A(_1322_),
    .B(_0185_));
 sg13g2_nor2_1 _2149_ (.A(net42),
    .B(_0186_),
    .Y(_0094_));
 sg13g2_nor2b_1 _2150_ (.A(_1254_),
    .B_N(_1326_),
    .Y(_0187_));
 sg13g2_xnor2_1 _2151_ (.Y(_0188_),
    .A(_1325_),
    .B(_0187_));
 sg13g2_and2_1 _2152_ (.A(net63),
    .B(_0188_),
    .X(_0095_));
 sg13g2_nor2_1 _2153_ (.A(_0962_),
    .B(_0966_),
    .Y(_0189_));
 sg13g2_a221oi_1 _2154_ (.B2(net64),
    .C1(_0835_),
    .B1(_0189_),
    .A1(_0958_),
    .Y(_0190_),
    .A2(_0963_));
 sg13g2_or2_1 _2155_ (.X(_0191_),
    .B(_0962_),
    .A(_0958_));
 sg13g2_inv_1 _2156_ (.Y(_0192_),
    .A(_0966_));
 sg13g2_a21o_1 _2157_ (.A2(_0191_),
    .A1(net64),
    .B1(_0192_),
    .X(_0193_));
 sg13g2_and2_1 _2158_ (.A(_0190_),
    .B(_0193_),
    .X(_0194_));
 sg13g2_buf_1 _2159_ (.A(_0194_),
    .X(_0195_));
 sg13g2_xnor2_1 _2160_ (.Y(_0196_),
    .A(\genblk4[3].pwm.accumulator[0] ),
    .B(net27));
 sg13g2_nor2_1 _2161_ (.A(net42),
    .B(_0196_),
    .Y(_0096_));
 sg13g2_nand2_1 _2162_ (.Y(_0197_),
    .A(net74),
    .B(_0192_));
 sg13g2_nor2_2 _2163_ (.A(net48),
    .B(_0197_),
    .Y(_0198_));
 sg13g2_nor2_1 _2164_ (.A(\genblk4[3].pwm.accumulator[9] ),
    .B(_0198_),
    .Y(_0199_));
 sg13g2_nand2b_2 _2165_ (.Y(_0200_),
    .B(_0962_),
    .A_N(\chan[3].attenuation.control[0] ));
 sg13g2_a21o_1 _2166_ (.A2(_0200_),
    .A1(net49),
    .B1(_0197_),
    .X(_0201_));
 sg13g2_or2_1 _2167_ (.X(_0202_),
    .B(_0966_),
    .A(\chan[3].attenuation.control[0] ));
 sg13g2_nand2b_1 _2168_ (.Y(_0203_),
    .B(net47),
    .A_N(net48));
 sg13g2_a21oi_1 _2169_ (.A1(_0202_),
    .A2(_0203_),
    .Y(_0204_),
    .B1(net49));
 sg13g2_or2_1 _2170_ (.X(_0205_),
    .B(_0962_),
    .A(\chan[3].attenuation.control[0] ));
 sg13g2_nand3_1 _2171_ (.B(net64),
    .C(_0962_),
    .A(_0958_),
    .Y(_0206_));
 sg13g2_a21oi_1 _2172_ (.A1(_0205_),
    .A2(_0206_),
    .Y(_0207_),
    .B1(net47));
 sg13g2_o21ai_1 _2173_ (.B1(net74),
    .Y(_0208_),
    .A1(_0204_),
    .A2(_0207_));
 sg13g2_buf_2 _2174_ (.A(_0208_),
    .X(_0209_));
 sg13g2_mux2_1 _2175_ (.A0(_0200_),
    .A1(net48),
    .S(net49),
    .X(_0210_));
 sg13g2_nor3_1 _2176_ (.A(net49),
    .B(net64),
    .C(net48),
    .Y(_0211_));
 sg13g2_a21o_1 _2177_ (.A2(net48),
    .A1(net64),
    .B1(net47),
    .X(_0212_));
 sg13g2_o21ai_1 _2178_ (.B1(net74),
    .Y(_0213_),
    .A1(_0211_),
    .A2(_0212_));
 sg13g2_a21oi_2 _2179_ (.B1(_0213_),
    .Y(_0214_),
    .A2(_0210_),
    .A1(net47));
 sg13g2_inv_1 _2180_ (.Y(_0215_),
    .A(_0214_));
 sg13g2_nor2b_1 _2181_ (.A(net49),
    .B_N(net48),
    .Y(_0216_));
 sg13g2_nor3_1 _2182_ (.A(net64),
    .B(_0192_),
    .C(_0216_),
    .Y(_0217_));
 sg13g2_or2_1 _2183_ (.X(_0218_),
    .B(net47),
    .A(net48));
 sg13g2_nand3_1 _2184_ (.B(net48),
    .C(net47),
    .A(net64),
    .Y(_0219_));
 sg13g2_a21oi_1 _2185_ (.A1(_0218_),
    .A2(_0219_),
    .Y(_0220_),
    .B1(net49));
 sg13g2_o21ai_1 _2186_ (.B1(net74),
    .Y(_0221_),
    .A1(_0217_),
    .A2(_0220_));
 sg13g2_xor2_1 _2187_ (.B(_0962_),
    .A(_0958_),
    .X(_0222_));
 sg13g2_and3_1 _2188_ (.X(_0223_),
    .A(net64),
    .B(net47),
    .C(_0222_));
 sg13g2_nor2_1 _2189_ (.A(_0958_),
    .B(_0202_),
    .Y(_0224_));
 sg13g2_o21ai_1 _2190_ (.B1(net74),
    .Y(_0225_),
    .A1(_0223_),
    .A2(_0224_));
 sg13g2_buf_2 _2191_ (.A(_0225_),
    .X(_0226_));
 sg13g2_nand2_1 _2192_ (.Y(_0227_),
    .A(_0955_),
    .B(_0962_));
 sg13g2_o21ai_1 _2193_ (.B1(_0205_),
    .Y(_0228_),
    .A1(_0967_),
    .A2(_0227_));
 sg13g2_nor2_1 _2194_ (.A(net49),
    .B(_0212_),
    .Y(_0229_));
 sg13g2_a21oi_1 _2195_ (.A1(_0959_),
    .A2(_0228_),
    .Y(_0230_),
    .B1(_0229_));
 sg13g2_nand2b_1 _2196_ (.Y(_0231_),
    .B(net74),
    .A_N(_0230_));
 sg13g2_buf_2 _2197_ (.A(_0231_),
    .X(_0232_));
 sg13g2_or2_1 _2198_ (.X(_0233_),
    .B(_0205_),
    .A(_0192_));
 sg13g2_a21o_1 _2199_ (.A2(_0227_),
    .A1(_0202_),
    .B1(_0958_),
    .X(_0234_));
 sg13g2_a21oi_2 _2200_ (.B1(_0835_),
    .Y(_0235_),
    .A2(_0234_),
    .A1(_0233_));
 sg13g2_and3_1 _2201_ (.X(_0236_),
    .A(\genblk4[3].pwm.accumulator[0] ),
    .B(_0190_),
    .C(_0193_));
 sg13g2_nand2_1 _2202_ (.Y(_0237_),
    .A(_0235_),
    .B(_0236_));
 sg13g2_o21ai_1 _2203_ (.B1(\genblk4[3].pwm.accumulator[1] ),
    .Y(_0238_),
    .A1(_0235_),
    .A2(_0236_));
 sg13g2_nand3_1 _2204_ (.B(_0237_),
    .C(_0238_),
    .A(_0232_),
    .Y(_0239_));
 sg13g2_a21oi_1 _2205_ (.A1(_0237_),
    .A2(_0238_),
    .Y(_0240_),
    .B1(_0232_));
 sg13g2_a21oi_1 _2206_ (.A1(\genblk4[3].pwm.accumulator[2] ),
    .A2(_0239_),
    .Y(_0241_),
    .B1(_0240_));
 sg13g2_nand2_1 _2207_ (.Y(_0242_),
    .A(_0958_),
    .B(_0966_));
 sg13g2_or2_1 _2208_ (.X(_0243_),
    .B(_0242_),
    .A(_0200_));
 sg13g2_a21o_1 _2209_ (.A2(_0206_),
    .A1(_0191_),
    .B1(net47),
    .X(_0244_));
 sg13g2_a21o_1 _2210_ (.A2(_0244_),
    .A1(_0243_),
    .B1(_0835_),
    .X(_0245_));
 sg13g2_buf_2 _2211_ (.A(_0245_),
    .X(_0246_));
 sg13g2_or2_1 _2212_ (.X(_0247_),
    .B(_0246_),
    .A(_0241_));
 sg13g2_inv_1 _2213_ (.Y(_0248_),
    .A(\genblk4[3].pwm.accumulator[3] ));
 sg13g2_a21o_1 _2214_ (.A2(_0246_),
    .A1(_0241_),
    .B1(_0248_),
    .X(_0249_));
 sg13g2_nand3_1 _2215_ (.B(_0247_),
    .C(_0249_),
    .A(_0226_),
    .Y(_0250_));
 sg13g2_a21oi_1 _2216_ (.A1(_0247_),
    .A2(_0249_),
    .Y(_0251_),
    .B1(_0226_));
 sg13g2_a21oi_1 _2217_ (.A1(\genblk4[3].pwm.accumulator[4] ),
    .A2(_0250_),
    .Y(_0252_),
    .B1(_0251_));
 sg13g2_or2_1 _2218_ (.X(_0253_),
    .B(_0252_),
    .A(_0221_));
 sg13g2_buf_1 _2219_ (.A(_0253_),
    .X(_0254_));
 sg13g2_inv_1 _2220_ (.Y(_0255_),
    .A(\genblk4[3].pwm.accumulator[5] ));
 sg13g2_a21o_1 _2221_ (.A2(_0252_),
    .A1(_0221_),
    .B1(_0255_),
    .X(_0256_));
 sg13g2_nand3_1 _2222_ (.B(_0254_),
    .C(_0256_),
    .A(_0215_),
    .Y(_0257_));
 sg13g2_a21oi_1 _2223_ (.A1(_0254_),
    .A2(_0256_),
    .Y(_0258_),
    .B1(_0215_));
 sg13g2_a21oi_2 _2224_ (.B1(_0258_),
    .Y(_0259_),
    .A2(_0257_),
    .A1(\genblk4[3].pwm.accumulator[6] ));
 sg13g2_nand2_1 _2225_ (.Y(_0260_),
    .A(_0209_),
    .B(_0259_));
 sg13g2_nor2_1 _2226_ (.A(_0209_),
    .B(_0259_),
    .Y(_0261_));
 sg13g2_a21oi_2 _2227_ (.B1(_0261_),
    .Y(_0262_),
    .A2(_0260_),
    .A1(\genblk4[3].pwm.accumulator[7] ));
 sg13g2_nor2_1 _2228_ (.A(_0201_),
    .B(_0262_),
    .Y(_0263_));
 sg13g2_nand2_1 _2229_ (.Y(_0264_),
    .A(_0201_),
    .B(_0262_));
 sg13g2_o21ai_1 _2230_ (.B1(_0264_),
    .Y(_0265_),
    .A1(\genblk4[3].pwm.accumulator[8] ),
    .A2(_0263_));
 sg13g2_nand2_1 _2231_ (.Y(_0266_),
    .A(\genblk4[3].pwm.accumulator[9] ),
    .B(_0198_));
 sg13g2_o21ai_1 _2232_ (.B1(_0266_),
    .Y(_0267_),
    .A1(_0199_),
    .A2(_0265_));
 sg13g2_and2_1 _2233_ (.A(net63),
    .B(_0267_),
    .X(_0097_));
 sg13g2_xnor2_1 _2234_ (.Y(_0268_),
    .A(_0235_),
    .B(_0236_));
 sg13g2_xor2_1 _2235_ (.B(_0268_),
    .A(\genblk4[3].pwm.accumulator[1] ),
    .X(_0269_));
 sg13g2_nor2_1 _2236_ (.A(net42),
    .B(_0269_),
    .Y(_0098_));
 sg13g2_xor2_1 _2237_ (.B(_0232_),
    .A(\genblk4[3].pwm.accumulator[2] ),
    .X(_0270_));
 sg13g2_and3_1 _2238_ (.X(_0271_),
    .A(_0237_),
    .B(_0238_),
    .C(_0270_));
 sg13g2_a21oi_1 _2239_ (.A1(_0237_),
    .A2(_0238_),
    .Y(_0272_),
    .B1(_0270_));
 sg13g2_nor3_1 _2240_ (.A(net59),
    .B(_0271_),
    .C(_0272_),
    .Y(_0099_));
 sg13g2_xnor2_1 _2241_ (.Y(_0273_),
    .A(_0248_),
    .B(_0246_));
 sg13g2_xnor2_1 _2242_ (.Y(_0274_),
    .A(_0241_),
    .B(_0273_));
 sg13g2_nor2_1 _2243_ (.A(net42),
    .B(_0274_),
    .Y(_0100_));
 sg13g2_nand2_1 _2244_ (.Y(_0275_),
    .A(_0247_),
    .B(_0249_));
 sg13g2_xnor2_1 _2245_ (.Y(_0276_),
    .A(\genblk4[3].pwm.accumulator[4] ),
    .B(_0226_));
 sg13g2_xnor2_1 _2246_ (.Y(_0277_),
    .A(_0275_),
    .B(_0276_));
 sg13g2_nor2_1 _2247_ (.A(net42),
    .B(_0277_),
    .Y(_0101_));
 sg13g2_xnor2_1 _2248_ (.Y(_0278_),
    .A(_0255_),
    .B(_0221_));
 sg13g2_xnor2_1 _2249_ (.Y(_0279_),
    .A(_0252_),
    .B(_0278_));
 sg13g2_nor2_1 _2250_ (.A(net42),
    .B(_0279_),
    .Y(_0102_));
 sg13g2_xnor2_1 _2251_ (.Y(_0280_),
    .A(\genblk4[3].pwm.accumulator[6] ),
    .B(_0214_));
 sg13g2_and3_1 _2252_ (.X(_0281_),
    .A(_0254_),
    .B(_0256_),
    .C(_0280_));
 sg13g2_a21oi_1 _2253_ (.A1(_0254_),
    .A2(_0256_),
    .Y(_0282_),
    .B1(_0280_));
 sg13g2_nor3_1 _2254_ (.A(net59),
    .B(_0281_),
    .C(_0282_),
    .Y(_0103_));
 sg13g2_xor2_1 _2255_ (.B(_0209_),
    .A(\genblk4[3].pwm.accumulator[7] ),
    .X(_0283_));
 sg13g2_xnor2_1 _2256_ (.Y(_0284_),
    .A(_0259_),
    .B(_0283_));
 sg13g2_nor2_1 _2257_ (.A(net42),
    .B(_0284_),
    .Y(_0104_));
 sg13g2_a21oi_2 _2258_ (.B1(_0197_),
    .Y(_0285_),
    .A2(_0200_),
    .A1(net49));
 sg13g2_xnor2_1 _2259_ (.Y(_0286_),
    .A(\genblk4[3].pwm.accumulator[8] ),
    .B(_0285_));
 sg13g2_xnor2_1 _2260_ (.Y(_0287_),
    .A(_0262_),
    .B(_0286_));
 sg13g2_nor2_1 _2261_ (.A(net42),
    .B(_0287_),
    .Y(_0105_));
 sg13g2_buf_1 _2262_ (.A(_0823_),
    .X(_0288_));
 sg13g2_nor2b_1 _2263_ (.A(_0199_),
    .B_N(_0266_),
    .Y(_0289_));
 sg13g2_xnor2_1 _2264_ (.Y(_0290_),
    .A(_0265_),
    .B(_0289_));
 sg13g2_and2_1 _2265_ (.A(net60),
    .B(_0290_),
    .X(_0106_));
 sg13g2_mux2_1 _2266_ (.A0(_0862_),
    .A1(\latch_control_reg[0] ),
    .S(_0865_),
    .X(_0291_));
 sg13g2_and2_1 _2267_ (.A(net60),
    .B(_0291_),
    .X(_0107_));
 sg13g2_buf_1 _2268_ (.A(net73),
    .X(_0292_));
 sg13g2_nor2_1 _2269_ (.A(_1001_),
    .B(_0865_),
    .Y(_0293_));
 sg13g2_a21oi_1 _2270_ (.A1(_0885_),
    .A2(_0865_),
    .Y(_0294_),
    .B1(_0293_));
 sg13g2_nor2_1 _2271_ (.A(net41),
    .B(_0294_),
    .Y(_0108_));
 sg13g2_nor2_1 _2272_ (.A(_0912_),
    .B(_0865_),
    .Y(_0295_));
 sg13g2_a21oi_1 _2273_ (.A1(\latch_control_reg[2] ),
    .A2(_0865_),
    .Y(_0296_),
    .B1(_0295_));
 sg13g2_nor2_1 _2274_ (.A(net41),
    .B(_0296_),
    .Y(_0109_));
 sg13g2_nor3_1 _2275_ (.A(\clk_counter[5] ),
    .B(\clk_counter[4] ),
    .C(\clk_counter[6] ),
    .Y(_0297_));
 sg13g2_nor4_1 _2276_ (.A(\clk_counter[1] ),
    .B(\clk_counter[0] ),
    .C(\clk_counter[3] ),
    .D(\clk_counter[2] ),
    .Y(_0298_));
 sg13g2_o21ai_1 _2277_ (.B1(_0298_),
    .Y(_0299_),
    .A1(net6),
    .A2(_0297_));
 sg13g2_nor2_1 _2278_ (.A(net6),
    .B(_0298_),
    .Y(_0300_));
 sg13g2_a21oi_2 _2279_ (.B1(_0300_),
    .Y(_0301_),
    .A2(_0299_),
    .A1(net7));
 sg13g2_buf_1 _2280_ (.A(_0301_),
    .X(_0302_));
 sg13g2_buf_1 _2281_ (.A(net34),
    .X(_0303_));
 sg13g2_nand2_1 _2282_ (.Y(_0304_),
    .A(_0006_),
    .B(net26));
 sg13g2_a21o_1 _2283_ (.A2(_0299_),
    .A1(net7),
    .B1(_0300_),
    .X(_0305_));
 sg13g2_buf_1 _2284_ (.A(_0305_),
    .X(_0306_));
 sg13g2_buf_1 _2285_ (.A(net33),
    .X(_0307_));
 sg13g2_nand2_1 _2286_ (.Y(_0308_),
    .A(\noise[0].gen.counter[0] ),
    .B(net25));
 sg13g2_a21oi_1 _2287_ (.A1(_0304_),
    .A2(_0308_),
    .Y(_0110_),
    .B1(net44));
 sg13g2_nand2_1 _2288_ (.Y(_0309_),
    .A(\noise[0].gen.counter[0] ),
    .B(net34));
 sg13g2_xor2_1 _2289_ (.B(_0309_),
    .A(\noise[0].gen.counter[1] ),
    .X(_0310_));
 sg13g2_nor2_1 _2290_ (.A(_0292_),
    .B(_0310_),
    .Y(_0111_));
 sg13g2_inv_1 _2291_ (.Y(_0311_),
    .A(\noise[0].gen.counter[2] ));
 sg13g2_nand3_1 _2292_ (.B(\noise[0].gen.counter[0] ),
    .C(_0301_),
    .A(\noise[0].gen.counter[1] ),
    .Y(_0312_));
 sg13g2_xnor2_1 _2293_ (.Y(_0313_),
    .A(_0311_),
    .B(_0312_));
 sg13g2_nor2_1 _2294_ (.A(net41),
    .B(_0313_),
    .Y(_0112_));
 sg13g2_nor2_2 _2295_ (.A(_0311_),
    .B(_0312_),
    .Y(_0314_));
 sg13g2_xnor2_1 _2296_ (.Y(_0315_),
    .A(\noise[0].gen.counter[3] ),
    .B(_0314_));
 sg13g2_nor2_1 _2297_ (.A(net41),
    .B(_0315_),
    .Y(_0113_));
 sg13g2_nand2_1 _2298_ (.Y(_0316_),
    .A(\noise[0].gen.counter[3] ),
    .B(_0314_));
 sg13g2_xor2_1 _2299_ (.B(_0316_),
    .A(\noise[0].gen.counter[4] ),
    .X(_0317_));
 sg13g2_nor2_1 _2300_ (.A(net41),
    .B(_0317_),
    .Y(_0114_));
 sg13g2_nand3_1 _2301_ (.B(\noise[0].gen.counter[4] ),
    .C(_0314_),
    .A(\noise[0].gen.counter[3] ),
    .Y(_0318_));
 sg13g2_xor2_1 _2302_ (.B(_0318_),
    .A(\noise[0].gen.counter[5] ),
    .X(_0319_));
 sg13g2_nor2_1 _2303_ (.A(net41),
    .B(_0319_),
    .Y(_0115_));
 sg13g2_nand4_1 _2304_ (.B(\noise[0].gen.counter[3] ),
    .C(\noise[0].gen.counter[4] ),
    .A(\noise[0].gen.counter[5] ),
    .Y(_0320_),
    .D(_0314_));
 sg13g2_xor2_1 _2305_ (.B(_0320_),
    .A(\noise[0].gen.counter[6] ),
    .X(_0321_));
 sg13g2_nor2_1 _2306_ (.A(net41),
    .B(_0321_),
    .Y(_0116_));
 sg13g2_and2_1 _2307_ (.A(_0288_),
    .B(_0813_),
    .X(_0132_));
 sg13g2_nand3_1 _2308_ (.B(_1042_),
    .C(_1044_),
    .A(net62),
    .Y(_0322_));
 sg13g2_buf_1 _2309_ (.A(_0322_),
    .X(_0323_));
 sg13g2_xnor2_1 _2310_ (.Y(_0324_),
    .A(_1146_),
    .B(_1250_));
 sg13g2_xnor2_1 _2311_ (.Y(_0325_),
    .A(_0323_),
    .B(_0324_));
 sg13g2_xnor2_1 _2312_ (.Y(_0326_),
    .A(net27),
    .B(_0325_));
 sg13g2_xnor2_1 _2313_ (.Y(_0327_),
    .A(\pwm.accumulator[0] ),
    .B(_0326_));
 sg13g2_nor2_1 _2314_ (.A(net41),
    .B(_0327_),
    .Y(_0133_));
 sg13g2_nand2_1 _2315_ (.Y(_0328_),
    .A(_1159_),
    .B(_1264_));
 sg13g2_o21ai_1 _2316_ (.B1(_1100_),
    .Y(_0329_),
    .A1(_1159_),
    .A2(_1264_));
 sg13g2_xnor2_1 _2317_ (.Y(_0330_),
    .A(_1214_),
    .B(_1256_));
 sg13g2_xnor2_1 _2318_ (.Y(_0331_),
    .A(_1106_),
    .B(_0330_));
 sg13g2_a21oi_1 _2319_ (.A1(_0328_),
    .A2(_0329_),
    .Y(_0332_),
    .B1(_0331_));
 sg13g2_nand3_1 _2320_ (.B(_0329_),
    .C(_0331_),
    .A(_0328_),
    .Y(_0333_));
 sg13g2_o21ai_1 _2321_ (.B1(_0333_),
    .Y(_0334_),
    .A1(_0201_),
    .A2(_0332_));
 sg13g2_buf_1 _2322_ (.A(_0334_),
    .X(_0335_));
 sg13g2_a21o_1 _2323_ (.A2(_1256_),
    .A1(_1214_),
    .B1(_1106_),
    .X(_0336_));
 sg13g2_o21ai_1 _2324_ (.B1(_0336_),
    .Y(_0337_),
    .A1(_1214_),
    .A2(_1256_));
 sg13g2_buf_1 _2325_ (.A(_0337_),
    .X(_0338_));
 sg13g2_xnor2_1 _2326_ (.Y(_0339_),
    .A(_1151_),
    .B(_1253_));
 sg13g2_xor2_1 _2327_ (.B(_0339_),
    .A(_1111_),
    .X(_0340_));
 sg13g2_xor2_1 _2328_ (.B(_0340_),
    .A(_0198_),
    .X(_0341_));
 sg13g2_xnor2_1 _2329_ (.Y(_0342_),
    .A(_0338_),
    .B(_0341_));
 sg13g2_xnor2_1 _2330_ (.Y(_0343_),
    .A(_0335_),
    .B(_0342_));
 sg13g2_nand2b_1 _2331_ (.Y(_0344_),
    .B(_0343_),
    .A_N(\pwm.accumulator[9] ));
 sg13g2_or2_1 _2332_ (.X(_0345_),
    .B(_0343_),
    .A(\pwm.accumulator[9] ));
 sg13g2_nand2_1 _2333_ (.Y(_0346_),
    .A(_0328_),
    .B(_0329_));
 sg13g2_xnor2_1 _2334_ (.Y(_0347_),
    .A(_0285_),
    .B(_0331_));
 sg13g2_xnor2_1 _2335_ (.Y(_0348_),
    .A(_0346_),
    .B(_0347_));
 sg13g2_nand2_1 _2336_ (.Y(_0349_),
    .A(_1166_),
    .B(_1271_));
 sg13g2_o21ai_1 _2337_ (.B1(_1053_),
    .Y(_0350_),
    .A1(_1166_),
    .A2(_1271_));
 sg13g2_nand2_1 _2338_ (.Y(_0351_),
    .A(_0349_),
    .B(_0350_));
 sg13g2_xnor2_1 _2339_ (.Y(_0352_),
    .A(_1159_),
    .B(_1264_));
 sg13g2_xnor2_1 _2340_ (.Y(_0353_),
    .A(_1100_),
    .B(_0352_));
 sg13g2_nand2_1 _2341_ (.Y(_0354_),
    .A(_0351_),
    .B(_0353_));
 sg13g2_o21ai_1 _2342_ (.B1(_0209_),
    .Y(_0355_),
    .A1(_0351_),
    .A2(_0353_));
 sg13g2_nand2_1 _2343_ (.Y(_0356_),
    .A(_0354_),
    .B(_0355_));
 sg13g2_nand2_1 _2344_ (.Y(_0357_),
    .A(_0348_),
    .B(_0356_));
 sg13g2_xnor2_1 _2345_ (.Y(_0358_),
    .A(_0209_),
    .B(_0351_));
 sg13g2_xnor2_1 _2346_ (.Y(_0359_),
    .A(_0353_),
    .B(_0358_));
 sg13g2_nand2_1 _2347_ (.Y(_0360_),
    .A(_1203_),
    .B(_1278_));
 sg13g2_nor2_1 _2348_ (.A(_1203_),
    .B(_1278_),
    .Y(_0361_));
 sg13g2_a21o_1 _2349_ (.A2(_0360_),
    .A1(_1090_),
    .B1(_0361_),
    .X(_0362_));
 sg13g2_xor2_1 _2350_ (.B(_1166_),
    .A(_1053_),
    .X(_0363_));
 sg13g2_xnor2_1 _2351_ (.Y(_0364_),
    .A(_1271_),
    .B(_0363_));
 sg13g2_a21oi_1 _2352_ (.A1(_0214_),
    .A2(_0362_),
    .Y(_0365_),
    .B1(_0364_));
 sg13g2_nor2_1 _2353_ (.A(_0214_),
    .B(_0362_),
    .Y(_0366_));
 sg13g2_nor2_1 _2354_ (.A(_0365_),
    .B(_0366_),
    .Y(_0367_));
 sg13g2_nor2b_1 _2355_ (.A(_0359_),
    .B_N(_0367_),
    .Y(_0368_));
 sg13g2_a21o_1 _2356_ (.A2(_1066_),
    .A1(_1064_),
    .B1(_1054_),
    .X(_0369_));
 sg13g2_a21oi_2 _2357_ (.B1(_1245_),
    .Y(_0370_),
    .A2(_1282_),
    .A1(_1280_));
 sg13g2_xnor2_1 _2358_ (.Y(_0371_),
    .A(_1223_),
    .B(_0370_));
 sg13g2_xnor2_1 _2359_ (.Y(_0372_),
    .A(_0369_),
    .B(_0371_));
 sg13g2_a22oi_1 _2360_ (.Y(_0373_),
    .B1(_1288_),
    .B2(_1289_),
    .A2(_1178_),
    .A1(_1177_));
 sg13g2_nand4_1 _2361_ (.B(_1178_),
    .C(_1288_),
    .A(_1177_),
    .Y(_0374_),
    .D(_1289_));
 sg13g2_o21ai_1 _2362_ (.B1(_0374_),
    .Y(_0375_),
    .A1(_1115_),
    .A2(_0373_));
 sg13g2_or2_1 _2363_ (.X(_0376_),
    .B(_0375_),
    .A(_0232_));
 sg13g2_and2_1 _2364_ (.A(_0232_),
    .B(_0375_),
    .X(_0377_));
 sg13g2_a21oi_2 _2365_ (.B1(_0377_),
    .Y(_0378_),
    .A2(_0376_),
    .A1(_0372_));
 sg13g2_nand3_1 _2366_ (.B(_1143_),
    .C(_1145_),
    .A(_1140_),
    .Y(_0379_));
 sg13g2_buf_2 _2367_ (.A(_0379_),
    .X(_0380_));
 sg13g2_nand3_1 _2368_ (.B(_1246_),
    .C(_1248_),
    .A(_1244_),
    .Y(_0381_));
 sg13g2_and2_1 _2369_ (.A(_0381_),
    .B(net27),
    .X(_0382_));
 sg13g2_nand3_1 _2370_ (.B(_0380_),
    .C(_0382_),
    .A(_1045_),
    .Y(_0383_));
 sg13g2_nand3_1 _2371_ (.B(_1146_),
    .C(_0382_),
    .A(_0323_),
    .Y(_0384_));
 sg13g2_xor2_1 _2372_ (.B(_1179_),
    .A(_1115_),
    .X(_0385_));
 sg13g2_xor2_1 _2373_ (.B(_0235_),
    .A(_1290_),
    .X(_0386_));
 sg13g2_xnor2_1 _2374_ (.Y(_0387_),
    .A(_0385_),
    .B(_0386_));
 sg13g2_a21oi_2 _2375_ (.B1(_0387_),
    .Y(_0388_),
    .A2(_0384_),
    .A1(_0383_));
 sg13g2_and4_1 _2376_ (.A(_0323_),
    .B(_0380_),
    .C(_1250_),
    .D(net27),
    .X(_0389_));
 sg13g2_nor2_1 _2377_ (.A(_0323_),
    .B(_0380_),
    .Y(_0390_));
 sg13g2_and3_1 _2378_ (.X(_0391_),
    .A(_1250_),
    .B(net27),
    .C(_0390_));
 sg13g2_mux2_1 _2379_ (.A0(_0389_),
    .A1(_0391_),
    .S(_0387_),
    .X(_0392_));
 sg13g2_xnor2_1 _2380_ (.Y(_0393_),
    .A(_0232_),
    .B(_0375_));
 sg13g2_xor2_1 _2381_ (.B(_0393_),
    .A(_0372_),
    .X(_0394_));
 sg13g2_nor4_1 _2382_ (.A(_0378_),
    .B(_0388_),
    .C(_0392_),
    .D(_0394_),
    .Y(_0395_));
 sg13g2_xnor2_1 _2383_ (.Y(_0396_),
    .A(_1171_),
    .B(_1303_));
 sg13g2_xnor2_1 _2384_ (.Y(_0397_),
    .A(_1074_),
    .B(_0396_));
 sg13g2_nand2_1 _2385_ (.Y(_0398_),
    .A(_1175_),
    .B(_1284_));
 sg13g2_nor2_1 _2386_ (.A(_0369_),
    .B(_0246_),
    .Y(_0399_));
 sg13g2_nand2_1 _2387_ (.Y(_0400_),
    .A(_0243_),
    .B(_0244_));
 sg13g2_a22oi_1 _2388_ (.Y(_0401_),
    .B1(_0400_),
    .B2(net74),
    .A2(_0370_),
    .A1(_1223_));
 sg13g2_o21ai_1 _2389_ (.B1(_1067_),
    .Y(_0402_),
    .A1(_1223_),
    .A2(_0370_));
 sg13g2_nor3_1 _2390_ (.A(_1175_),
    .B(_1284_),
    .C(_0246_),
    .Y(_0403_));
 sg13g2_a221oi_1 _2391_ (.B2(_0402_),
    .C1(_0403_),
    .B1(_0401_),
    .A1(_0398_),
    .Y(_0404_),
    .A2(_0399_));
 sg13g2_xnor2_1 _2392_ (.Y(_0405_),
    .A(_0397_),
    .B(_0404_));
 sg13g2_nor4_1 _2393_ (.A(_0405_),
    .B(_0388_),
    .C(_0392_),
    .D(_0394_),
    .Y(_0406_));
 sg13g2_xnor2_1 _2394_ (.Y(_0407_),
    .A(_1290_),
    .B(_0385_));
 sg13g2_nor2_1 _2395_ (.A(_0380_),
    .B(_0381_),
    .Y(_0408_));
 sg13g2_a21oi_1 _2396_ (.A1(_0380_),
    .A2(_0381_),
    .Y(_0409_),
    .B1(_0323_));
 sg13g2_o21ai_1 _2397_ (.B1(_0235_),
    .Y(_0410_),
    .A1(_0408_),
    .A2(_0409_));
 sg13g2_nor3_1 _2398_ (.A(_0235_),
    .B(_0408_),
    .C(_0409_),
    .Y(_0411_));
 sg13g2_a21oi_2 _2399_ (.B1(_0411_),
    .Y(_0412_),
    .A2(_0410_),
    .A1(_0407_));
 sg13g2_nor4_1 _2400_ (.A(_0378_),
    .B(_0388_),
    .C(_0392_),
    .D(_0412_),
    .Y(_0413_));
 sg13g2_nor4_1 _2401_ (.A(_0405_),
    .B(_0388_),
    .C(_0392_),
    .D(_0412_),
    .Y(_0414_));
 sg13g2_nor4_2 _2402_ (.A(_0395_),
    .B(_0406_),
    .C(_0413_),
    .Y(_0415_),
    .D(_0414_));
 sg13g2_nor2_1 _2403_ (.A(_0378_),
    .B(_0405_),
    .Y(_0416_));
 sg13g2_nor3_1 _2404_ (.A(_0378_),
    .B(_0394_),
    .C(_0412_),
    .Y(_0417_));
 sg13g2_nor3_1 _2405_ (.A(_0405_),
    .B(_0394_),
    .C(_0412_),
    .Y(_0418_));
 sg13g2_nor3_1 _2406_ (.A(_0416_),
    .B(_0417_),
    .C(_0418_),
    .Y(_0419_));
 sg13g2_xor2_1 _2407_ (.B(_1278_),
    .A(_1203_),
    .X(_0420_));
 sg13g2_xnor2_1 _2408_ (.Y(_0421_),
    .A(_1090_),
    .B(_0420_));
 sg13g2_inv_1 _2409_ (.Y(_0422_),
    .A(_0221_));
 sg13g2_nand2b_1 _2410_ (.Y(_0423_),
    .B(net75),
    .A_N(_1309_));
 sg13g2_nor2_1 _2411_ (.A(_1193_),
    .B(_0423_),
    .Y(_0424_));
 sg13g2_a21oi_1 _2412_ (.A1(_1193_),
    .A2(_0423_),
    .Y(_0425_),
    .B1(_1082_));
 sg13g2_nor3_1 _2413_ (.A(_0422_),
    .B(_0424_),
    .C(_0425_),
    .Y(_0426_));
 sg13g2_o21ai_1 _2414_ (.B1(_0422_),
    .Y(_0427_),
    .A1(_0424_),
    .A2(_0425_));
 sg13g2_nor2b_1 _2415_ (.A(_0426_),
    .B_N(_0427_),
    .Y(_0428_));
 sg13g2_xor2_1 _2416_ (.B(_0428_),
    .A(_0421_),
    .X(_0429_));
 sg13g2_a21oi_2 _2417_ (.B1(_0426_),
    .Y(_0430_),
    .A2(_0427_),
    .A1(_0421_));
 sg13g2_nor2_1 _2418_ (.A(_1271_),
    .B(_0214_),
    .Y(_0431_));
 sg13g2_and2_1 _2419_ (.A(_1271_),
    .B(_0214_),
    .X(_0432_));
 sg13g2_o21ai_1 _2420_ (.B1(_0363_),
    .Y(_0433_),
    .A1(_0431_),
    .A2(_0432_));
 sg13g2_a21oi_1 _2421_ (.A1(net50),
    .A2(_1266_),
    .Y(_0434_),
    .B1(_1269_));
 sg13g2_or2_1 _2422_ (.X(_0435_),
    .B(_0214_),
    .A(_0434_));
 sg13g2_nand2_1 _2423_ (.Y(_0436_),
    .A(_0434_),
    .B(_0214_));
 sg13g2_a21o_1 _2424_ (.A2(_0436_),
    .A1(_0435_),
    .B1(_0363_),
    .X(_0437_));
 sg13g2_a21o_1 _2425_ (.A2(_0437_),
    .A1(_0433_),
    .B1(_0362_),
    .X(_0438_));
 sg13g2_nand3_1 _2426_ (.B(_0433_),
    .C(_0437_),
    .A(_0362_),
    .Y(_0439_));
 sg13g2_nand3_1 _2427_ (.B(_0438_),
    .C(_0439_),
    .A(_0430_),
    .Y(_0440_));
 sg13g2_or2_1 _2428_ (.X(_0441_),
    .B(_0397_),
    .A(_0246_));
 sg13g2_nand2_1 _2429_ (.Y(_0442_),
    .A(_1223_),
    .B(_0370_));
 sg13g2_and2_1 _2430_ (.A(_0442_),
    .B(_0402_),
    .X(_0443_));
 sg13g2_a21o_1 _2431_ (.A2(_0397_),
    .A1(_0246_),
    .B1(_0443_),
    .X(_0444_));
 sg13g2_xnor2_1 _2432_ (.Y(_0445_),
    .A(_1082_),
    .B(_1193_));
 sg13g2_xnor2_1 _2433_ (.Y(_0446_),
    .A(_1310_),
    .B(_0445_));
 sg13g2_a21o_1 _2434_ (.A2(_1303_),
    .A1(_1171_),
    .B1(_1074_),
    .X(_0447_));
 sg13g2_or4_1 _2435_ (.A(_1245_),
    .B(_1142_),
    .C(_1169_),
    .D(_1301_),
    .X(_0448_));
 sg13g2_and2_1 _2436_ (.A(_0226_),
    .B(_0448_),
    .X(_0449_));
 sg13g2_nor2_1 _2437_ (.A(_1074_),
    .B(_0226_),
    .Y(_0450_));
 sg13g2_nand2_1 _2438_ (.Y(_0451_),
    .A(_1171_),
    .B(_1303_));
 sg13g2_nor2_1 _2439_ (.A(_0226_),
    .B(_0448_),
    .Y(_0452_));
 sg13g2_a221oi_1 _2440_ (.B2(_0451_),
    .C1(_0452_),
    .B1(_0450_),
    .A1(_0447_),
    .Y(_0453_),
    .A2(_0449_));
 sg13g2_xnor2_1 _2441_ (.Y(_0454_),
    .A(_0446_),
    .B(_0453_));
 sg13g2_a21o_1 _2442_ (.A2(_0444_),
    .A1(_0441_),
    .B1(_0454_),
    .X(_0455_));
 sg13g2_buf_1 _2443_ (.A(_0455_),
    .X(_0456_));
 sg13g2_nand3_1 _2444_ (.B(_0440_),
    .C(net22),
    .A(_0429_),
    .Y(_0457_));
 sg13g2_and2_1 _2445_ (.A(_0448_),
    .B(_0447_),
    .X(_0458_));
 sg13g2_nand2b_1 _2446_ (.Y(_0459_),
    .B(_0446_),
    .A_N(_0226_));
 sg13g2_nor2b_1 _2447_ (.A(_0446_),
    .B_N(_0226_),
    .Y(_0460_));
 sg13g2_a21o_1 _2448_ (.A2(_0459_),
    .A1(_0458_),
    .B1(_0460_),
    .X(_0461_));
 sg13g2_nand3_1 _2449_ (.B(_0440_),
    .C(net22),
    .A(_0461_),
    .Y(_0462_));
 sg13g2_a22oi_1 _2450_ (.Y(_0463_),
    .B1(_0457_),
    .B2(_0462_),
    .A2(_0419_),
    .A1(_0415_));
 sg13g2_a21oi_2 _2451_ (.B1(_0460_),
    .Y(_0464_),
    .A2(_0459_),
    .A1(_0458_));
 sg13g2_nand3_1 _2452_ (.B(_0441_),
    .C(_0444_),
    .A(_0454_),
    .Y(_0465_));
 sg13g2_buf_2 _2453_ (.A(_0465_),
    .X(_0466_));
 sg13g2_nor2_1 _2454_ (.A(_0464_),
    .B(_0466_),
    .Y(_0467_));
 sg13g2_and2_1 _2455_ (.A(_0438_),
    .B(_0439_),
    .X(_0468_));
 sg13g2_xnor2_1 _2456_ (.Y(_0469_),
    .A(_0421_),
    .B(_0428_));
 sg13g2_a221oi_1 _2457_ (.B2(_0464_),
    .C1(_0469_),
    .B1(_0466_),
    .A1(_0430_),
    .Y(_0470_),
    .A2(_0468_));
 sg13g2_a21o_1 _2458_ (.A2(_0467_),
    .A1(_0440_),
    .B1(_0470_),
    .X(_0471_));
 sg13g2_nor2_1 _2459_ (.A(_0463_),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_nand2b_1 _2460_ (.Y(_0473_),
    .B(_0359_),
    .A_N(_0367_));
 sg13g2_or2_1 _2461_ (.X(_0474_),
    .B(_0468_),
    .A(_0430_));
 sg13g2_and3_1 _2462_ (.X(_0475_),
    .A(_0357_),
    .B(_0473_),
    .C(_0474_));
 sg13g2_nor2_1 _2463_ (.A(_0348_),
    .B(_0356_),
    .Y(_0476_));
 sg13g2_a221oi_1 _2464_ (.B2(_0475_),
    .C1(_0476_),
    .B1(_0472_),
    .A1(_0357_),
    .Y(_0477_),
    .A2(_0368_));
 sg13g2_buf_2 _2465_ (.A(_0477_),
    .X(_0478_));
 sg13g2_mux2_1 _2466_ (.A0(_0344_),
    .A1(_0345_),
    .S(_0478_),
    .X(_0479_));
 sg13g2_buf_2 _2467_ (.A(_0479_),
    .X(_0480_));
 sg13g2_xnor2_1 _2468_ (.Y(_0481_),
    .A(_0348_),
    .B(_0356_));
 sg13g2_or2_1 _2469_ (.X(_0482_),
    .B(_0481_),
    .A(_0368_));
 sg13g2_and3_1 _2470_ (.X(_0483_),
    .A(_0473_),
    .B(_0474_),
    .C(_0481_));
 sg13g2_inv_1 _2471_ (.Y(_0484_),
    .A(_0483_));
 sg13g2_mux2_1 _2472_ (.A0(_0482_),
    .A1(_0484_),
    .S(_0472_),
    .X(_0485_));
 sg13g2_or2_1 _2473_ (.X(_0486_),
    .B(_0474_),
    .A(_0368_));
 sg13g2_a21oi_1 _2474_ (.A1(_0473_),
    .A2(_0486_),
    .Y(_0487_),
    .B1(_0481_));
 sg13g2_a21oi_1 _2475_ (.A1(_0368_),
    .A2(_0481_),
    .Y(_0488_),
    .B1(_0487_));
 sg13g2_nand2_1 _2476_ (.Y(net17),
    .A(_0485_),
    .B(_0488_));
 sg13g2_nand2_1 _2477_ (.Y(_0489_),
    .A(_0474_),
    .B(_0472_));
 sg13g2_xnor2_1 _2478_ (.Y(_0490_),
    .A(_0359_),
    .B(_0367_));
 sg13g2_xnor2_1 _2479_ (.Y(net16),
    .A(_0489_),
    .B(_0490_));
 sg13g2_and3_1 _2480_ (.X(_0491_),
    .A(_0480_),
    .B(net17),
    .C(net16));
 sg13g2_and3_1 _2481_ (.X(_0492_),
    .A(\pwm.accumulator[8] ),
    .B(_0480_),
    .C(net16));
 sg13g2_inv_1 _2482_ (.Y(_0493_),
    .A(_0466_));
 sg13g2_xnor2_1 _2483_ (.Y(_0494_),
    .A(_0430_),
    .B(_0468_));
 sg13g2_or3_1 _2484_ (.A(_0429_),
    .B(_0493_),
    .C(net21),
    .X(_0495_));
 sg13g2_nand3b_1 _2485_ (.B(_0464_),
    .C(_0466_),
    .Y(_0496_),
    .A_N(net21));
 sg13g2_nand2_1 _2486_ (.Y(_0497_),
    .A(_0415_),
    .B(_0419_));
 sg13g2_a21oi_1 _2487_ (.A1(_0495_),
    .A2(_0496_),
    .Y(_0498_),
    .B1(_0497_));
 sg13g2_or3_1 _2488_ (.A(_0429_),
    .B(net22),
    .C(net21),
    .X(_0499_));
 sg13g2_or3_1 _2489_ (.A(_0461_),
    .B(net22),
    .C(net21),
    .X(_0500_));
 sg13g2_nand3b_1 _2490_ (.B(_0464_),
    .C(_0469_),
    .Y(_0501_),
    .A_N(net21));
 sg13g2_nand3_1 _2491_ (.B(_0493_),
    .C(net21),
    .A(_0429_),
    .Y(_0502_));
 sg13g2_nand4_1 _2492_ (.B(_0500_),
    .C(_0501_),
    .A(_0499_),
    .Y(_0503_),
    .D(_0502_));
 sg13g2_and4_1 _2493_ (.A(_0429_),
    .B(_0497_),
    .C(net22),
    .D(_0494_),
    .X(_0504_));
 sg13g2_a21o_1 _2494_ (.A2(_0384_),
    .A1(_0383_),
    .B1(_0387_),
    .X(_0505_));
 sg13g2_nand4_1 _2495_ (.B(_0380_),
    .C(_1250_),
    .A(_0323_),
    .Y(_0506_),
    .D(net27));
 sg13g2_nand3_1 _2496_ (.B(net27),
    .C(_0390_),
    .A(_1250_),
    .Y(_0507_));
 sg13g2_mux2_1 _2497_ (.A0(_0506_),
    .A1(_0507_),
    .S(_0387_),
    .X(_0508_));
 sg13g2_xnor2_1 _2498_ (.Y(_0509_),
    .A(_0372_),
    .B(_0393_));
 sg13g2_nand3_1 _2499_ (.B(_0508_),
    .C(_0509_),
    .A(_0505_),
    .Y(_0510_));
 sg13g2_a21oi_1 _2500_ (.A1(_0505_),
    .A2(_0508_),
    .Y(_0511_),
    .B1(_0509_));
 sg13g2_a221oi_1 _2501_ (.B2(_0412_),
    .C1(_0511_),
    .B1(_0510_),
    .A1(_0378_),
    .Y(_0512_),
    .A2(_0405_));
 sg13g2_nor2_1 _2502_ (.A(_0416_),
    .B(_0512_),
    .Y(_0513_));
 sg13g2_nand3_1 _2503_ (.B(net22),
    .C(net21),
    .A(_0461_),
    .Y(_0514_));
 sg13g2_nor2_1 _2504_ (.A(_0464_),
    .B(_0469_),
    .Y(_0515_));
 sg13g2_o21ai_1 _2505_ (.B1(net21),
    .Y(_0516_),
    .A1(_0467_),
    .A2(_0515_));
 sg13g2_o21ai_1 _2506_ (.B1(_0516_),
    .Y(_0517_),
    .A1(_0513_),
    .A2(_0514_));
 sg13g2_nor4_2 _2507_ (.A(_0498_),
    .B(_0503_),
    .C(_0504_),
    .Y(net15),
    .D(_0517_));
 sg13g2_a21oi_1 _2508_ (.A1(_0510_),
    .A2(_0412_),
    .Y(_0518_),
    .B1(_0511_));
 sg13g2_xor2_1 _2509_ (.B(_0405_),
    .A(_0378_),
    .X(_0519_));
 sg13g2_xnor2_1 _2510_ (.Y(_0520_),
    .A(_0518_),
    .B(_0519_));
 sg13g2_nor2_1 _2511_ (.A(_0408_),
    .B(_0409_),
    .Y(_0521_));
 sg13g2_xor2_1 _2512_ (.B(_0521_),
    .A(_0387_),
    .X(_0522_));
 sg13g2_and3_1 _2513_ (.X(_0523_),
    .A(\pwm.accumulator[0] ),
    .B(_0326_),
    .C(_0522_));
 sg13g2_nor3_1 _2514_ (.A(\pwm.accumulator[1] ),
    .B(\pwm.accumulator[2] ),
    .C(_0523_),
    .Y(_0524_));
 sg13g2_nor2_1 _2515_ (.A(_0388_),
    .B(_0392_),
    .Y(_0525_));
 sg13g2_xnor2_1 _2516_ (.Y(_0526_),
    .A(_0509_),
    .B(_0412_));
 sg13g2_nor2b_1 _2517_ (.A(_0525_),
    .B_N(_0526_),
    .Y(_0527_));
 sg13g2_nand2_1 _2518_ (.Y(_0528_),
    .A(\pwm.accumulator[0] ),
    .B(net27));
 sg13g2_nor2_1 _2519_ (.A(\pwm.accumulator[0] ),
    .B(_0195_),
    .Y(_0529_));
 sg13g2_a21oi_1 _2520_ (.A1(_0325_),
    .A2(_0528_),
    .Y(_0530_),
    .B1(_0529_));
 sg13g2_or2_1 _2521_ (.X(_0531_),
    .B(_0530_),
    .A(_0522_));
 sg13g2_a21o_1 _2522_ (.A2(_0530_),
    .A1(_0522_),
    .B1(\pwm.accumulator[1] ),
    .X(_0532_));
 sg13g2_a21oi_1 _2523_ (.A1(_0531_),
    .A2(_0532_),
    .Y(_0533_),
    .B1(_0526_));
 sg13g2_a21oi_1 _2524_ (.A1(_0531_),
    .A2(_0526_),
    .Y(_0534_),
    .B1(\pwm.accumulator[2] ));
 sg13g2_nor4_2 _2525_ (.A(_0524_),
    .B(_0527_),
    .C(_0533_),
    .Y(_0535_),
    .D(_0534_));
 sg13g2_a21oi_1 _2526_ (.A1(_0520_),
    .A2(_0535_),
    .Y(_0536_),
    .B1(\pwm.accumulator[3] ));
 sg13g2_nor2_1 _2527_ (.A(_0520_),
    .B(_0535_),
    .Y(_0537_));
 sg13g2_nand2_1 _2528_ (.Y(_0538_),
    .A(_0466_),
    .B(net22));
 sg13g2_o21ai_1 _2529_ (.B1(_0538_),
    .Y(_0539_),
    .A1(_0416_),
    .A2(_0512_));
 sg13g2_nand4_1 _2530_ (.B(_0415_),
    .C(_0419_),
    .A(_0466_),
    .Y(_0540_),
    .D(net22));
 sg13g2_nand3_1 _2531_ (.B(_0539_),
    .C(_0540_),
    .A(\pwm.accumulator[4] ),
    .Y(_0541_));
 sg13g2_o21ai_1 _2532_ (.B1(_0541_),
    .Y(_0542_),
    .A1(_0536_),
    .A2(_0537_));
 sg13g2_nand2_1 _2533_ (.Y(_0543_),
    .A(_0539_),
    .B(_0540_));
 sg13g2_nand2b_1 _2534_ (.Y(_0544_),
    .B(_0543_),
    .A_N(\pwm.accumulator[4] ));
 sg13g2_o21ai_1 _2535_ (.B1(_0456_),
    .Y(_0545_),
    .A1(_0416_),
    .A2(_0512_));
 sg13g2_xnor2_1 _2536_ (.Y(_0546_),
    .A(_0464_),
    .B(_0429_));
 sg13g2_a21oi_2 _2537_ (.B1(_0546_),
    .Y(_0547_),
    .A2(_0545_),
    .A1(_0466_));
 sg13g2_and3_1 _2538_ (.X(_0548_),
    .A(_0466_),
    .B(_0545_),
    .C(_0546_));
 sg13g2_inv_1 _2539_ (.Y(_0549_),
    .A(\pwm.accumulator[5] ));
 sg13g2_o21ai_1 _2540_ (.B1(_0549_),
    .Y(_0550_),
    .A1(_0547_),
    .A2(_0548_));
 sg13g2_nand4_1 _2541_ (.B(_0542_),
    .C(_0544_),
    .A(net15),
    .Y(_0551_),
    .D(_0550_));
 sg13g2_nor3_2 _2542_ (.A(_0549_),
    .B(_0547_),
    .C(_0548_),
    .Y(_0552_));
 sg13g2_o21ai_1 _2543_ (.B1(net15),
    .Y(_0553_),
    .A1(\pwm.accumulator[6] ),
    .A2(_0552_));
 sg13g2_nand2_1 _2544_ (.Y(_0554_),
    .A(\pwm.accumulator[6] ),
    .B(_0552_));
 sg13g2_nand4_1 _2545_ (.B(_0542_),
    .C(_0544_),
    .A(\pwm.accumulator[6] ),
    .Y(_0555_),
    .D(_0550_));
 sg13g2_nand4_1 _2546_ (.B(_0553_),
    .C(_0554_),
    .A(_0551_),
    .Y(_0556_),
    .D(_0555_));
 sg13g2_buf_2 _2547_ (.A(_0556_),
    .X(_0557_));
 sg13g2_o21ai_1 _2548_ (.B1(_0557_),
    .Y(_0558_),
    .A1(_0491_),
    .A2(_0492_));
 sg13g2_buf_1 _2549_ (.A(\pwm.accumulator[7] ),
    .X(_0559_));
 sg13g2_and3_1 _2550_ (.X(_0560_),
    .A(_0559_),
    .B(_0480_),
    .C(net17));
 sg13g2_and3_1 _2551_ (.X(_0561_),
    .A(_0559_),
    .B(\pwm.accumulator[8] ),
    .C(_0480_));
 sg13g2_o21ai_1 _2552_ (.B1(_0557_),
    .Y(_0562_),
    .A1(_0560_),
    .A2(_0561_));
 sg13g2_inv_1 _2553_ (.Y(_0563_),
    .A(\pwm.accumulator[8] ));
 sg13g2_a21oi_1 _2554_ (.A1(_0485_),
    .A2(_0488_),
    .Y(_0564_),
    .B1(_0563_));
 sg13g2_and4_1 _2555_ (.A(_0559_),
    .B(\pwm.accumulator[8] ),
    .C(_0480_),
    .D(net16),
    .X(_0565_));
 sg13g2_a221oi_1 _2556_ (.B2(_0559_),
    .C1(_0565_),
    .B1(_0491_),
    .A1(_0480_),
    .Y(_0566_),
    .A2(_0564_));
 sg13g2_xnor2_1 _2557_ (.Y(net18),
    .A(_0478_),
    .B(_0343_));
 sg13g2_nand2_1 _2558_ (.Y(_0567_),
    .A(\pwm.accumulator[9] ),
    .B(net18));
 sg13g2_nand4_1 _2559_ (.B(_0562_),
    .C(_0566_),
    .A(_0558_),
    .Y(_0568_),
    .D(_0567_));
 sg13g2_nor2_1 _2560_ (.A(_1151_),
    .B(_1253_),
    .Y(_0569_));
 sg13g2_a21oi_1 _2561_ (.A1(_1151_),
    .A2(_1253_),
    .Y(_0570_),
    .B1(_1111_));
 sg13g2_nor2_2 _2562_ (.A(_0569_),
    .B(_0570_),
    .Y(_0571_));
 sg13g2_nand2_1 _2563_ (.Y(_0572_),
    .A(_0338_),
    .B(_0340_));
 sg13g2_nor2_1 _2564_ (.A(_0335_),
    .B(_0572_),
    .Y(_0573_));
 sg13g2_nor2_1 _2565_ (.A(_0338_),
    .B(_0340_),
    .Y(_0574_));
 sg13g2_o21ai_1 _2566_ (.B1(_0572_),
    .Y(_0575_),
    .A1(_0335_),
    .A2(_0574_));
 sg13g2_or2_1 _2567_ (.X(_0576_),
    .B(_0573_),
    .A(_0198_));
 sg13g2_a21o_1 _2568_ (.A2(_0575_),
    .A1(_0478_),
    .B1(_0576_),
    .X(_0577_));
 sg13g2_inv_1 _2569_ (.Y(_0578_),
    .A(_0338_));
 sg13g2_nand2_1 _2570_ (.Y(_0579_),
    .A(_0335_),
    .B(_0578_));
 sg13g2_nor2_1 _2571_ (.A(_0340_),
    .B(_0579_),
    .Y(_0580_));
 sg13g2_nor2b_1 _2572_ (.A(_0580_),
    .B_N(_0198_),
    .Y(_0581_));
 sg13g2_o21ai_1 _2573_ (.B1(_0581_),
    .Y(_0582_),
    .A1(_0478_),
    .A2(_0575_));
 sg13g2_nor2b_1 _2574_ (.A(_0478_),
    .B_N(_0580_),
    .Y(_0583_));
 sg13g2_a221oi_1 _2575_ (.B2(_0582_),
    .C1(_0583_),
    .B1(_0577_),
    .A1(_0478_),
    .Y(_0584_),
    .A2(_0573_));
 sg13g2_xor2_1 _2576_ (.B(_0584_),
    .A(_0571_),
    .X(net19));
 sg13g2_and2_1 _2577_ (.A(\pwm.accumulator[10] ),
    .B(net19),
    .X(_0585_));
 sg13g2_inv_1 _2578_ (.Y(_0586_),
    .A(\pwm.accumulator[10] ));
 sg13g2_nand2b_1 _2579_ (.Y(_0587_),
    .B(_0586_),
    .A_N(net19));
 sg13g2_nand2b_1 _2580_ (.Y(_0588_),
    .B(_0587_),
    .A_N(_0585_));
 sg13g2_xnor2_1 _2581_ (.Y(_0589_),
    .A(_0568_),
    .B(_0588_));
 sg13g2_and2_1 _2582_ (.A(net60),
    .B(_0589_),
    .X(_0134_));
 sg13g2_a21oi_1 _2583_ (.A1(_0568_),
    .A2(_0587_),
    .Y(_0590_),
    .B1(_0585_));
 sg13g2_nand2b_1 _2584_ (.Y(_0591_),
    .B(_0338_),
    .A_N(_0335_));
 sg13g2_inv_1 _2585_ (.Y(_0592_),
    .A(_0579_));
 sg13g2_a21oi_1 _2586_ (.A1(_0198_),
    .A2(_0591_),
    .Y(_0593_),
    .B1(_0592_));
 sg13g2_nor2_1 _2587_ (.A(_0478_),
    .B(_0340_),
    .Y(_0594_));
 sg13g2_nor2_1 _2588_ (.A(_0571_),
    .B(_0594_),
    .Y(_0595_));
 sg13g2_nand2b_1 _2589_ (.Y(_0596_),
    .B(_0579_),
    .A_N(_0571_));
 sg13g2_a22oi_1 _2590_ (.Y(_0597_),
    .B1(_0596_),
    .B2(_0198_),
    .A2(_0591_),
    .A1(_0571_));
 sg13g2_a21oi_1 _2591_ (.A1(_0478_),
    .A2(_0340_),
    .Y(_0598_),
    .B1(_0597_));
 sg13g2_a21oi_1 _2592_ (.A1(_0571_),
    .A2(_0594_),
    .Y(_0599_),
    .B1(_0598_));
 sg13g2_o21ai_1 _2593_ (.B1(_0599_),
    .Y(net20),
    .A1(_0593_),
    .A2(_0595_));
 sg13g2_nand2_1 _2594_ (.Y(_0600_),
    .A(\pwm.accumulator[11] ),
    .B(net20));
 sg13g2_or2_1 _2595_ (.X(_0601_),
    .B(net20),
    .A(\pwm.accumulator[11] ));
 sg13g2_and2_1 _2596_ (.A(_0600_),
    .B(_0601_),
    .X(_0602_));
 sg13g2_xnor2_1 _2597_ (.Y(_0603_),
    .A(_0590_),
    .B(_0602_));
 sg13g2_and2_1 _2598_ (.A(net60),
    .B(_0603_),
    .X(_0135_));
 sg13g2_and3_1 _2599_ (.X(_0604_),
    .A(_0558_),
    .B(_0562_),
    .C(_0566_));
 sg13g2_nor2b_1 _2600_ (.A(net19),
    .B_N(_0567_),
    .Y(_0605_));
 sg13g2_a21oi_1 _2601_ (.A1(_0604_),
    .A2(_0605_),
    .Y(_0606_),
    .B1(_0586_));
 sg13g2_and2_1 _2602_ (.A(_0568_),
    .B(net19),
    .X(_0607_));
 sg13g2_o21ai_1 _2603_ (.B1(_0601_),
    .Y(_0608_),
    .A1(_0606_),
    .A2(_0607_));
 sg13g2_a21oi_1 _2604_ (.A1(_0600_),
    .A2(_0608_),
    .Y(_0136_),
    .B1(net44));
 sg13g2_xor2_1 _2605_ (.B(_0530_),
    .A(\pwm.accumulator[1] ),
    .X(_0609_));
 sg13g2_xnor2_1 _2606_ (.Y(_0610_),
    .A(_0522_),
    .B(_0609_));
 sg13g2_nor2_1 _2607_ (.A(_0292_),
    .B(_0610_),
    .Y(_0137_));
 sg13g2_buf_1 _2608_ (.A(net73),
    .X(_0611_));
 sg13g2_nand2_1 _2609_ (.Y(_0612_),
    .A(_0531_),
    .B(_0532_));
 sg13g2_xnor2_1 _2610_ (.Y(_0613_),
    .A(\pwm.accumulator[2] ),
    .B(_0526_));
 sg13g2_xnor2_1 _2611_ (.Y(_0614_),
    .A(_0612_),
    .B(_0613_));
 sg13g2_nor2_1 _2612_ (.A(_0611_),
    .B(_0614_),
    .Y(_0138_));
 sg13g2_xnor2_1 _2613_ (.Y(_0615_),
    .A(_0520_),
    .B(_0535_));
 sg13g2_xnor2_1 _2614_ (.Y(_0616_),
    .A(\pwm.accumulator[3] ),
    .B(_0615_));
 sg13g2_and2_1 _2615_ (.A(net60),
    .B(_0616_),
    .X(_0139_));
 sg13g2_nor2_1 _2616_ (.A(_0536_),
    .B(_0537_),
    .Y(_0617_));
 sg13g2_and2_1 _2617_ (.A(_0541_),
    .B(_0544_),
    .X(_0618_));
 sg13g2_xnor2_1 _2618_ (.Y(_0619_),
    .A(_0617_),
    .B(_0618_));
 sg13g2_nor2_1 _2619_ (.A(net40),
    .B(_0619_),
    .Y(_0140_));
 sg13g2_and2_1 _2620_ (.A(_0542_),
    .B(_0544_),
    .X(_0620_));
 sg13g2_nand2b_1 _2621_ (.Y(_0621_),
    .B(_0550_),
    .A_N(_0552_));
 sg13g2_xnor2_1 _2622_ (.Y(_0622_),
    .A(_0620_),
    .B(_0621_));
 sg13g2_and2_1 _2623_ (.A(net60),
    .B(_0622_),
    .X(_0141_));
 sg13g2_a21oi_1 _2624_ (.A1(_0620_),
    .A2(_0550_),
    .Y(_0623_),
    .B1(_0552_));
 sg13g2_xnor2_1 _2625_ (.Y(_0624_),
    .A(\pwm.accumulator[6] ),
    .B(net15));
 sg13g2_xnor2_1 _2626_ (.Y(_0625_),
    .A(_0623_),
    .B(_0624_));
 sg13g2_nor2_1 _2627_ (.A(net40),
    .B(_0625_),
    .Y(_0142_));
 sg13g2_xor2_1 _2628_ (.B(net16),
    .A(_0559_),
    .X(_0626_));
 sg13g2_xnor2_1 _2629_ (.Y(_0627_),
    .A(_0557_),
    .B(_0626_));
 sg13g2_nor2_1 _2630_ (.A(net40),
    .B(_0627_),
    .Y(_0143_));
 sg13g2_nand2_1 _2631_ (.Y(_0628_),
    .A(_0557_),
    .B(net16));
 sg13g2_o21ai_1 _2632_ (.B1(_0559_),
    .Y(_0629_),
    .A1(_0557_),
    .A2(net16));
 sg13g2_nand2_1 _2633_ (.Y(_0630_),
    .A(_0628_),
    .B(_0629_));
 sg13g2_xnor2_1 _2634_ (.Y(_0631_),
    .A(_0563_),
    .B(net17));
 sg13g2_xnor2_1 _2635_ (.Y(_0632_),
    .A(_0630_),
    .B(_0631_));
 sg13g2_nor2_1 _2636_ (.A(net40),
    .B(_0632_),
    .Y(_0144_));
 sg13g2_nand3_1 _2637_ (.B(_0485_),
    .C(_0488_),
    .A(_0563_),
    .Y(_0633_));
 sg13g2_a21oi_1 _2638_ (.A1(_0633_),
    .A2(_0630_),
    .Y(_0634_),
    .B1(_0564_));
 sg13g2_nand2_1 _2639_ (.Y(_0635_),
    .A(_0480_),
    .B(_0567_));
 sg13g2_xnor2_1 _2640_ (.Y(_0636_),
    .A(_0634_),
    .B(_0635_));
 sg13g2_nor2_1 _2641_ (.A(net40),
    .B(_0636_),
    .Y(_0145_));
 sg13g2_nor2_1 _2642_ (.A(\tone[0].gen.counter[1] ),
    .B(\tone[0].gen.counter[0] ),
    .Y(_0637_));
 sg13g2_nor4_1 _2643_ (.A(\tone[0].gen.counter[3] ),
    .B(\tone[0].gen.counter[6] ),
    .C(\tone[0].gen.counter[9] ),
    .D(\tone[0].gen.counter[8] ),
    .Y(_0638_));
 sg13g2_nor4_1 _2644_ (.A(\tone[0].gen.counter[2] ),
    .B(\tone[0].gen.counter[5] ),
    .C(\tone[0].gen.counter[4] ),
    .D(\tone[0].gen.counter[7] ),
    .Y(_0639_));
 sg13g2_and3_1 _2645_ (.X(_0640_),
    .A(_0637_),
    .B(_0638_),
    .C(_0639_));
 sg13g2_buf_1 _2646_ (.A(_0640_),
    .X(_0641_));
 sg13g2_buf_1 _2647_ (.A(_0641_),
    .X(_0642_));
 sg13g2_a21oi_1 _2648_ (.A1(\control_tone_freq[0][0] ),
    .A2(net32),
    .Y(_0643_),
    .B1(\tone[0].gen.counter[0] ));
 sg13g2_nand2_1 _2649_ (.Y(_0644_),
    .A(net26),
    .B(_0643_));
 sg13g2_nand2_1 _2650_ (.Y(_0645_),
    .A(\tone[0].gen.counter[0] ),
    .B(net25));
 sg13g2_a21oi_1 _2651_ (.A1(_0644_),
    .A2(_0645_),
    .Y(_0147_),
    .B1(net44));
 sg13g2_buf_1 _2652_ (.A(net34),
    .X(_0646_));
 sg13g2_xor2_1 _2653_ (.B(\control_tone_freq[0][1] ),
    .A(\control_tone_freq[0][0] ),
    .X(_0647_));
 sg13g2_a21oi_1 _2654_ (.A1(net32),
    .A2(_0647_),
    .Y(_0648_),
    .B1(\tone[0].gen.counter[1] ));
 sg13g2_nand3b_1 _2655_ (.B(net24),
    .C(_0648_),
    .Y(_0649_),
    .A_N(\tone[0].gen.counter[0] ));
 sg13g2_o21ai_1 _2656_ (.B1(\tone[0].gen.counter[1] ),
    .Y(_0650_),
    .A1(\tone[0].gen.counter[0] ),
    .A2(net25));
 sg13g2_a21oi_1 _2657_ (.A1(_0649_),
    .A2(_0650_),
    .Y(_0148_),
    .B1(net44));
 sg13g2_o21ai_1 _2658_ (.B1(_0641_),
    .Y(_0651_),
    .A1(\control_tone_freq[0][0] ),
    .A2(\control_tone_freq[0][1] ));
 sg13g2_a21oi_1 _2659_ (.A1(\control_tone_freq[0][2] ),
    .A2(_0641_),
    .Y(_0652_),
    .B1(\tone[0].gen.counter[2] ));
 sg13g2_nand3_1 _2660_ (.B(_0651_),
    .C(_0652_),
    .A(_0637_),
    .Y(_0653_));
 sg13g2_nand2_1 _2661_ (.Y(_0654_),
    .A(_0637_),
    .B(_0651_));
 sg13g2_nand3_1 _2662_ (.B(net32),
    .C(_0654_),
    .A(\control_tone_freq[0][2] ),
    .Y(_0655_));
 sg13g2_buf_1 _2663_ (.A(net33),
    .X(_0656_));
 sg13g2_a21o_1 _2664_ (.A2(_0655_),
    .A1(_0653_),
    .B1(net23),
    .X(_0657_));
 sg13g2_o21ai_1 _2665_ (.B1(\tone[0].gen.counter[2] ),
    .Y(_0658_),
    .A1(net25),
    .A2(_0654_));
 sg13g2_a21oi_1 _2666_ (.A1(_0657_),
    .A2(_0658_),
    .Y(_0149_),
    .B1(_1026_));
 sg13g2_and2_1 _2667_ (.A(\control_tone_freq[0][3] ),
    .B(_0641_),
    .X(_0659_));
 sg13g2_nor3_2 _2668_ (.A(\tone[0].gen.counter[3] ),
    .B(_0653_),
    .C(_0659_),
    .Y(_0660_));
 sg13g2_and2_1 _2669_ (.A(_0653_),
    .B(_0659_),
    .X(_0661_));
 sg13g2_o21ai_1 _2670_ (.B1(net24),
    .Y(_0662_),
    .A1(_0660_),
    .A2(_0661_));
 sg13g2_o21ai_1 _2671_ (.B1(\tone[0].gen.counter[3] ),
    .Y(_0663_),
    .A1(net25),
    .A2(_0653_));
 sg13g2_a21oi_1 _2672_ (.A1(_0662_),
    .A2(_0663_),
    .Y(_0150_),
    .B1(_1026_));
 sg13g2_a21oi_1 _2673_ (.A1(\control_tone_freq[0][4] ),
    .A2(_0641_),
    .Y(_0664_),
    .B1(\tone[0].gen.counter[4] ));
 sg13g2_and2_1 _2674_ (.A(_0660_),
    .B(_0664_),
    .X(_0665_));
 sg13g2_nand3b_1 _2675_ (.B(net32),
    .C(\control_tone_freq[0][4] ),
    .Y(_0666_),
    .A_N(_0660_));
 sg13g2_nand2b_1 _2676_ (.Y(_0667_),
    .B(_0666_),
    .A_N(_0665_));
 sg13g2_nand2_1 _2677_ (.Y(_0668_),
    .A(net24),
    .B(_0660_));
 sg13g2_a22oi_1 _2678_ (.Y(_0669_),
    .B1(_0668_),
    .B2(\tone[0].gen.counter[4] ),
    .A2(_0667_),
    .A1(net26));
 sg13g2_nor2_1 _2679_ (.A(net40),
    .B(_0669_),
    .Y(_0151_));
 sg13g2_nand2_1 _2680_ (.Y(_0670_),
    .A(\control_tone_freq[0][5] ),
    .B(_0642_));
 sg13g2_nand3b_1 _2681_ (.B(_0665_),
    .C(_0670_),
    .Y(_0671_),
    .A_N(\tone[0].gen.counter[5] ));
 sg13g2_o21ai_1 _2682_ (.B1(_0671_),
    .Y(_0672_),
    .A1(_0665_),
    .A2(_0670_));
 sg13g2_nand2_1 _2683_ (.Y(_0673_),
    .A(net34),
    .B(_0665_));
 sg13g2_a22oi_1 _2684_ (.Y(_0674_),
    .B1(_0673_),
    .B2(\tone[0].gen.counter[5] ),
    .A2(_0672_),
    .A1(net26));
 sg13g2_nor2_1 _2685_ (.A(net40),
    .B(_0674_),
    .Y(_0152_));
 sg13g2_a21oi_1 _2686_ (.A1(\control_tone_freq[0][6] ),
    .A2(net32),
    .Y(_0675_),
    .B1(\tone[0].gen.counter[6] ));
 sg13g2_nand2b_2 _2687_ (.Y(_0676_),
    .B(_0675_),
    .A_N(_0671_));
 sg13g2_nand3_1 _2688_ (.B(net32),
    .C(_0671_),
    .A(\control_tone_freq[0][6] ),
    .Y(_0677_));
 sg13g2_a21o_1 _2689_ (.A2(_0677_),
    .A1(_0676_),
    .B1(net23),
    .X(_0678_));
 sg13g2_o21ai_1 _2690_ (.B1(\tone[0].gen.counter[6] ),
    .Y(_0679_),
    .A1(net25),
    .A2(_0671_));
 sg13g2_buf_1 _2691_ (.A(net73),
    .X(_0680_));
 sg13g2_a21oi_1 _2692_ (.A1(_0678_),
    .A2(_0679_),
    .Y(_0153_),
    .B1(net39));
 sg13g2_and2_1 _2693_ (.A(\control_tone_freq[0][7] ),
    .B(_0642_),
    .X(_0681_));
 sg13g2_nor3_2 _2694_ (.A(\tone[0].gen.counter[7] ),
    .B(_0676_),
    .C(_0681_),
    .Y(_0682_));
 sg13g2_a21oi_1 _2695_ (.A1(_0676_),
    .A2(_0681_),
    .Y(_0683_),
    .B1(_0682_));
 sg13g2_o21ai_1 _2696_ (.B1(\tone[0].gen.counter[7] ),
    .Y(_0684_),
    .A1(net33),
    .A2(_0676_));
 sg13g2_o21ai_1 _2697_ (.B1(_0684_),
    .Y(_0685_),
    .A1(net33),
    .A2(_0683_));
 sg13g2_and2_1 _2698_ (.A(net60),
    .B(_0685_),
    .X(_0154_));
 sg13g2_and2_1 _2699_ (.A(\control_tone_freq[0][8] ),
    .B(net32),
    .X(_0686_));
 sg13g2_nor2_1 _2700_ (.A(\tone[0].gen.counter[8] ),
    .B(_0686_),
    .Y(_0687_));
 sg13g2_mux2_1 _2701_ (.A0(_0686_),
    .A1(_0687_),
    .S(_0682_),
    .X(_0688_));
 sg13g2_nand2_1 _2702_ (.Y(_0689_),
    .A(net34),
    .B(_0682_));
 sg13g2_a22oi_1 _2703_ (.Y(_0690_),
    .B1(_0689_),
    .B2(\tone[0].gen.counter[8] ),
    .A2(_0688_),
    .A1(_0303_));
 sg13g2_nor2_1 _2704_ (.A(_0611_),
    .B(_0690_),
    .Y(_0155_));
 sg13g2_nor3_1 _2705_ (.A(\tone[0].gen.counter[8] ),
    .B(_0686_),
    .C(_0689_),
    .Y(_0691_));
 sg13g2_and2_1 _2706_ (.A(_0301_),
    .B(net32),
    .X(_0692_));
 sg13g2_a21oi_1 _2707_ (.A1(\control_tone_freq[0][9] ),
    .A2(_0692_),
    .Y(_0693_),
    .B1(\tone[0].gen.counter[9] ));
 sg13g2_xor2_1 _2708_ (.B(_0693_),
    .A(_0691_),
    .X(_0694_));
 sg13g2_nor2_1 _2709_ (.A(net40),
    .B(_0694_),
    .Y(_0156_));
 sg13g2_nand2_1 _2710_ (.Y(_0695_),
    .A(_0000_),
    .B(_0692_));
 sg13g2_nand2b_1 _2711_ (.Y(_0696_),
    .B(_1040_),
    .A_N(_0692_));
 sg13g2_a21oi_1 _2712_ (.A1(_0695_),
    .A2(_0696_),
    .Y(_0157_),
    .B1(net39));
 sg13g2_nor2_1 _2713_ (.A(\tone[1].gen.counter[1] ),
    .B(\tone[1].gen.counter[0] ),
    .Y(_0697_));
 sg13g2_nor4_1 _2714_ (.A(\tone[1].gen.counter[3] ),
    .B(\tone[1].gen.counter[6] ),
    .C(\tone[1].gen.counter[9] ),
    .D(\tone[1].gen.counter[8] ),
    .Y(_0698_));
 sg13g2_nor4_1 _2715_ (.A(\tone[1].gen.counter[2] ),
    .B(\tone[1].gen.counter[5] ),
    .C(\tone[1].gen.counter[4] ),
    .D(\tone[1].gen.counter[7] ),
    .Y(_0699_));
 sg13g2_and3_1 _2716_ (.X(_0700_),
    .A(_0697_),
    .B(_0698_),
    .C(_0699_));
 sg13g2_buf_1 _2717_ (.A(_0700_),
    .X(_0701_));
 sg13g2_buf_1 _2718_ (.A(_0701_),
    .X(_0702_));
 sg13g2_a21oi_1 _2719_ (.A1(\control_tone_freq[1][0] ),
    .A2(net31),
    .Y(_0703_),
    .B1(\tone[1].gen.counter[0] ));
 sg13g2_nand2_1 _2720_ (.Y(_0704_),
    .A(net26),
    .B(_0703_));
 sg13g2_nand2_1 _2721_ (.Y(_0705_),
    .A(\tone[1].gen.counter[0] ),
    .B(net25));
 sg13g2_a21oi_1 _2722_ (.A1(_0704_),
    .A2(_0705_),
    .Y(_0158_),
    .B1(net39));
 sg13g2_xor2_1 _2723_ (.B(\control_tone_freq[1][1] ),
    .A(\control_tone_freq[1][0] ),
    .X(_0706_));
 sg13g2_a21oi_1 _2724_ (.A1(net31),
    .A2(_0706_),
    .Y(_0707_),
    .B1(\tone[1].gen.counter[1] ));
 sg13g2_nand3b_1 _2725_ (.B(net24),
    .C(_0707_),
    .Y(_0708_),
    .A_N(\tone[1].gen.counter[0] ));
 sg13g2_o21ai_1 _2726_ (.B1(\tone[1].gen.counter[1] ),
    .Y(_0709_),
    .A1(\tone[1].gen.counter[0] ),
    .A2(net25));
 sg13g2_a21oi_1 _2727_ (.A1(_0708_),
    .A2(_0709_),
    .Y(_0159_),
    .B1(net39));
 sg13g2_o21ai_1 _2728_ (.B1(_0701_),
    .Y(_0710_),
    .A1(\control_tone_freq[1][0] ),
    .A2(\control_tone_freq[1][1] ));
 sg13g2_a21oi_1 _2729_ (.A1(\control_tone_freq[1][2] ),
    .A2(_0701_),
    .Y(_0711_),
    .B1(\tone[1].gen.counter[2] ));
 sg13g2_nand3_1 _2730_ (.B(_0710_),
    .C(_0711_),
    .A(_0697_),
    .Y(_0712_));
 sg13g2_nand2_1 _2731_ (.Y(_0713_),
    .A(_0697_),
    .B(_0710_));
 sg13g2_nand3_1 _2732_ (.B(net31),
    .C(_0713_),
    .A(\control_tone_freq[1][2] ),
    .Y(_0714_));
 sg13g2_a21o_1 _2733_ (.A2(_0714_),
    .A1(_0712_),
    .B1(net23),
    .X(_0715_));
 sg13g2_o21ai_1 _2734_ (.B1(\tone[1].gen.counter[2] ),
    .Y(_0716_),
    .A1(net23),
    .A2(_0713_));
 sg13g2_a21oi_1 _2735_ (.A1(_0715_),
    .A2(_0716_),
    .Y(_0160_),
    .B1(net39));
 sg13g2_and2_1 _2736_ (.A(\control_tone_freq[1][3] ),
    .B(_0701_),
    .X(_0717_));
 sg13g2_nor3_2 _2737_ (.A(\tone[1].gen.counter[3] ),
    .B(_0712_),
    .C(_0717_),
    .Y(_0718_));
 sg13g2_and2_1 _2738_ (.A(_0712_),
    .B(_0717_),
    .X(_0719_));
 sg13g2_o21ai_1 _2739_ (.B1(net24),
    .Y(_0720_),
    .A1(_0718_),
    .A2(_0719_));
 sg13g2_o21ai_1 _2740_ (.B1(\tone[1].gen.counter[3] ),
    .Y(_0721_),
    .A1(net23),
    .A2(_0712_));
 sg13g2_a21oi_1 _2741_ (.A1(_0720_),
    .A2(_0721_),
    .Y(_0161_),
    .B1(net39));
 sg13g2_a21oi_1 _2742_ (.A1(\control_tone_freq[1][4] ),
    .A2(_0701_),
    .Y(_0722_),
    .B1(\tone[1].gen.counter[4] ));
 sg13g2_and2_1 _2743_ (.A(_0718_),
    .B(_0722_),
    .X(_0723_));
 sg13g2_nand3b_1 _2744_ (.B(net31),
    .C(\control_tone_freq[1][4] ),
    .Y(_0724_),
    .A_N(_0718_));
 sg13g2_nand2b_1 _2745_ (.Y(_0725_),
    .B(_0724_),
    .A_N(_0723_));
 sg13g2_nand2_1 _2746_ (.Y(_0726_),
    .A(net34),
    .B(_0718_));
 sg13g2_a22oi_1 _2747_ (.Y(_0727_),
    .B1(_0726_),
    .B2(\tone[1].gen.counter[4] ),
    .A2(_0725_),
    .A1(net26));
 sg13g2_nor2_1 _2748_ (.A(net46),
    .B(_0727_),
    .Y(_0162_));
 sg13g2_nand2_1 _2749_ (.Y(_0728_),
    .A(\control_tone_freq[1][5] ),
    .B(net31));
 sg13g2_nand3b_1 _2750_ (.B(_0723_),
    .C(_0728_),
    .Y(_0729_),
    .A_N(\tone[1].gen.counter[5] ));
 sg13g2_o21ai_1 _2751_ (.B1(_0729_),
    .Y(_0730_),
    .A1(_0723_),
    .A2(_0728_));
 sg13g2_nand2_1 _2752_ (.Y(_0731_),
    .A(net34),
    .B(_0723_));
 sg13g2_a22oi_1 _2753_ (.Y(_0732_),
    .B1(_0731_),
    .B2(\tone[1].gen.counter[5] ),
    .A2(_0730_),
    .A1(net26));
 sg13g2_nor2_1 _2754_ (.A(net46),
    .B(_0732_),
    .Y(_0163_));
 sg13g2_a21oi_1 _2755_ (.A1(\control_tone_freq[1][6] ),
    .A2(_0702_),
    .Y(_0733_),
    .B1(\tone[1].gen.counter[6] ));
 sg13g2_nand2b_2 _2756_ (.Y(_0734_),
    .B(_0733_),
    .A_N(_0729_));
 sg13g2_nand3_1 _2757_ (.B(_0702_),
    .C(_0729_),
    .A(\control_tone_freq[1][6] ),
    .Y(_0735_));
 sg13g2_a21o_1 _2758_ (.A2(_0735_),
    .A1(_0734_),
    .B1(net23),
    .X(_0736_));
 sg13g2_o21ai_1 _2759_ (.B1(\tone[1].gen.counter[6] ),
    .Y(_0737_),
    .A1(net23),
    .A2(_0729_));
 sg13g2_a21oi_1 _2760_ (.A1(_0736_),
    .A2(_0737_),
    .Y(_0164_),
    .B1(net39));
 sg13g2_and2_1 _2761_ (.A(\control_tone_freq[1][7] ),
    .B(net31),
    .X(_0738_));
 sg13g2_nor3_2 _2762_ (.A(\tone[1].gen.counter[7] ),
    .B(_0734_),
    .C(_0738_),
    .Y(_0739_));
 sg13g2_a21oi_1 _2763_ (.A1(_0734_),
    .A2(_0738_),
    .Y(_0740_),
    .B1(_0739_));
 sg13g2_o21ai_1 _2764_ (.B1(\tone[1].gen.counter[7] ),
    .Y(_0741_),
    .A1(net33),
    .A2(_0734_));
 sg13g2_o21ai_1 _2765_ (.B1(_0741_),
    .Y(_0742_),
    .A1(net33),
    .A2(_0740_));
 sg13g2_and2_1 _2766_ (.A(net60),
    .B(_0742_),
    .X(_0165_));
 sg13g2_and2_1 _2767_ (.A(\control_tone_freq[1][8] ),
    .B(net31),
    .X(_0743_));
 sg13g2_nor2_1 _2768_ (.A(\tone[1].gen.counter[8] ),
    .B(_0743_),
    .Y(_0744_));
 sg13g2_mux2_1 _2769_ (.A0(_0743_),
    .A1(_0744_),
    .S(_0739_),
    .X(_0745_));
 sg13g2_nand2_1 _2770_ (.Y(_0746_),
    .A(net34),
    .B(_0739_));
 sg13g2_a22oi_1 _2771_ (.Y(_0747_),
    .B1(_0746_),
    .B2(\tone[1].gen.counter[8] ),
    .A2(_0745_),
    .A1(net26));
 sg13g2_nor2_1 _2772_ (.A(net46),
    .B(_0747_),
    .Y(_0166_));
 sg13g2_nor3_1 _2773_ (.A(\tone[1].gen.counter[8] ),
    .B(_0743_),
    .C(_0746_),
    .Y(_0748_));
 sg13g2_and2_1 _2774_ (.A(_0301_),
    .B(net31),
    .X(_0749_));
 sg13g2_a21oi_1 _2775_ (.A1(\control_tone_freq[1][9] ),
    .A2(_0749_),
    .Y(_0750_),
    .B1(\tone[1].gen.counter[9] ));
 sg13g2_xor2_1 _2776_ (.B(_0750_),
    .A(_0748_),
    .X(_0751_));
 sg13g2_nor2_1 _2777_ (.A(net46),
    .B(_0751_),
    .Y(_0167_));
 sg13g2_nand2_1 _2778_ (.Y(_0752_),
    .A(_0001_),
    .B(_0749_));
 sg13g2_nand2b_1 _2779_ (.Y(_0753_),
    .B(_1148_),
    .A_N(_0749_));
 sg13g2_a21oi_1 _2780_ (.A1(_0752_),
    .A2(_0753_),
    .Y(_0168_),
    .B1(net39));
 sg13g2_nor2_1 _2781_ (.A(\tone[2].gen.counter[1] ),
    .B(\tone[2].gen.counter[0] ),
    .Y(_0754_));
 sg13g2_nor4_1 _2782_ (.A(\tone[2].gen.counter[3] ),
    .B(\tone[2].gen.counter[6] ),
    .C(\tone[2].gen.counter[9] ),
    .D(\tone[2].gen.counter[8] ),
    .Y(_0755_));
 sg13g2_nor4_1 _2783_ (.A(\tone[2].gen.counter[2] ),
    .B(\tone[2].gen.counter[5] ),
    .C(\tone[2].gen.counter[4] ),
    .D(\tone[2].gen.counter[7] ),
    .Y(_0756_));
 sg13g2_and3_1 _2784_ (.X(_0757_),
    .A(_0754_),
    .B(_0755_),
    .C(_0756_));
 sg13g2_buf_1 _2785_ (.A(_0757_),
    .X(_0758_));
 sg13g2_buf_1 _2786_ (.A(_0758_),
    .X(_0759_));
 sg13g2_a21oi_1 _2787_ (.A1(\control_tone_freq[2][0] ),
    .A2(net30),
    .Y(_0760_),
    .B1(\tone[2].gen.counter[0] ));
 sg13g2_nand2_1 _2788_ (.Y(_0761_),
    .A(_0303_),
    .B(_0760_));
 sg13g2_nand2_1 _2789_ (.Y(_0762_),
    .A(\tone[2].gen.counter[0] ),
    .B(_0307_));
 sg13g2_a21oi_1 _2790_ (.A1(_0761_),
    .A2(_0762_),
    .Y(_0169_),
    .B1(_0680_));
 sg13g2_xor2_1 _2791_ (.B(\control_tone_freq[2][1] ),
    .A(\control_tone_freq[2][0] ),
    .X(_0763_));
 sg13g2_a21oi_1 _2792_ (.A1(net30),
    .A2(_0763_),
    .Y(_0764_),
    .B1(\tone[2].gen.counter[1] ));
 sg13g2_nand3b_1 _2793_ (.B(net24),
    .C(_0764_),
    .Y(_0765_),
    .A_N(\tone[2].gen.counter[0] ));
 sg13g2_o21ai_1 _2794_ (.B1(\tone[2].gen.counter[1] ),
    .Y(_0766_),
    .A1(\tone[2].gen.counter[0] ),
    .A2(_0307_));
 sg13g2_a21oi_1 _2795_ (.A1(_0765_),
    .A2(_0766_),
    .Y(_0170_),
    .B1(_0680_));
 sg13g2_o21ai_1 _2796_ (.B1(_0758_),
    .Y(_0767_),
    .A1(\control_tone_freq[2][0] ),
    .A2(\control_tone_freq[2][1] ));
 sg13g2_a21oi_1 _2797_ (.A1(\control_tone_freq[2][2] ),
    .A2(_0758_),
    .Y(_0768_),
    .B1(\tone[2].gen.counter[2] ));
 sg13g2_nand3_1 _2798_ (.B(_0767_),
    .C(_0768_),
    .A(_0754_),
    .Y(_0769_));
 sg13g2_nand2_1 _2799_ (.Y(_0770_),
    .A(_0754_),
    .B(_0767_));
 sg13g2_nand3_1 _2800_ (.B(net30),
    .C(_0770_),
    .A(\control_tone_freq[2][2] ),
    .Y(_0771_));
 sg13g2_a21o_1 _2801_ (.A2(_0771_),
    .A1(_0769_),
    .B1(net33),
    .X(_0772_));
 sg13g2_o21ai_1 _2802_ (.B1(\tone[2].gen.counter[2] ),
    .Y(_0773_),
    .A1(net23),
    .A2(_0770_));
 sg13g2_a21oi_1 _2803_ (.A1(_0772_),
    .A2(_0773_),
    .Y(_0171_),
    .B1(net59));
 sg13g2_and2_1 _2804_ (.A(\control_tone_freq[2][3] ),
    .B(_0758_),
    .X(_0774_));
 sg13g2_nor3_2 _2805_ (.A(\tone[2].gen.counter[3] ),
    .B(_0769_),
    .C(_0774_),
    .Y(_0775_));
 sg13g2_and2_1 _2806_ (.A(_0769_),
    .B(_0774_),
    .X(_0776_));
 sg13g2_o21ai_1 _2807_ (.B1(net24),
    .Y(_0777_),
    .A1(_0775_),
    .A2(_0776_));
 sg13g2_o21ai_1 _2808_ (.B1(\tone[2].gen.counter[3] ),
    .Y(_0778_),
    .A1(_0656_),
    .A2(_0769_));
 sg13g2_a21oi_1 _2809_ (.A1(_0777_),
    .A2(_0778_),
    .Y(_0172_),
    .B1(net59));
 sg13g2_a21oi_1 _2810_ (.A1(\control_tone_freq[2][4] ),
    .A2(_0758_),
    .Y(_0779_),
    .B1(\tone[2].gen.counter[4] ));
 sg13g2_and2_1 _2811_ (.A(_0775_),
    .B(_0779_),
    .X(_0780_));
 sg13g2_nand3b_1 _2812_ (.B(net30),
    .C(\control_tone_freq[2][4] ),
    .Y(_0781_),
    .A_N(_0775_));
 sg13g2_nand2b_1 _2813_ (.Y(_0782_),
    .B(_0781_),
    .A_N(_0780_));
 sg13g2_nand2_1 _2814_ (.Y(_0783_),
    .A(_0302_),
    .B(_0775_));
 sg13g2_a22oi_1 _2815_ (.Y(_0784_),
    .B1(_0783_),
    .B2(\tone[2].gen.counter[4] ),
    .A2(_0782_),
    .A1(net24));
 sg13g2_nor2_1 _2816_ (.A(net46),
    .B(_0784_),
    .Y(_0173_));
 sg13g2_nand2_1 _2817_ (.Y(_0785_),
    .A(\control_tone_freq[2][5] ),
    .B(net30));
 sg13g2_nand3b_1 _2818_ (.B(_0780_),
    .C(_0785_),
    .Y(_0786_),
    .A_N(\tone[2].gen.counter[5] ));
 sg13g2_o21ai_1 _2819_ (.B1(_0786_),
    .Y(_0787_),
    .A1(_0780_),
    .A2(_0785_));
 sg13g2_nand2_1 _2820_ (.Y(_0788_),
    .A(_0302_),
    .B(_0780_));
 sg13g2_a22oi_1 _2821_ (.Y(_0789_),
    .B1(_0788_),
    .B2(\tone[2].gen.counter[5] ),
    .A2(_0787_),
    .A1(_0646_));
 sg13g2_nor2_1 _2822_ (.A(net46),
    .B(_0789_),
    .Y(_0174_));
 sg13g2_a21oi_1 _2823_ (.A1(\control_tone_freq[2][6] ),
    .A2(net30),
    .Y(_0790_),
    .B1(\tone[2].gen.counter[6] ));
 sg13g2_nand2b_2 _2824_ (.Y(_0791_),
    .B(_0790_),
    .A_N(_0786_));
 sg13g2_nand3_1 _2825_ (.B(net30),
    .C(_0786_),
    .A(\control_tone_freq[2][6] ),
    .Y(_0792_));
 sg13g2_a21o_1 _2826_ (.A2(_0792_),
    .A1(_0791_),
    .B1(net33),
    .X(_0793_));
 sg13g2_o21ai_1 _2827_ (.B1(\tone[2].gen.counter[6] ),
    .Y(_0794_),
    .A1(_0656_),
    .A2(_0786_));
 sg13g2_a21oi_1 _2828_ (.A1(_0793_),
    .A2(_0794_),
    .Y(_0175_),
    .B1(_0859_));
 sg13g2_and2_1 _2829_ (.A(\control_tone_freq[2][7] ),
    .B(_0759_),
    .X(_0795_));
 sg13g2_nor3_2 _2830_ (.A(\tone[2].gen.counter[7] ),
    .B(_0791_),
    .C(_0795_),
    .Y(_0796_));
 sg13g2_a21oi_1 _2831_ (.A1(_0791_),
    .A2(_0795_),
    .Y(_0797_),
    .B1(_0796_));
 sg13g2_o21ai_1 _2832_ (.B1(\tone[2].gen.counter[7] ),
    .Y(_0798_),
    .A1(_0306_),
    .A2(_0791_));
 sg13g2_o21ai_1 _2833_ (.B1(_0798_),
    .Y(_0799_),
    .A1(_0306_),
    .A2(_0797_));
 sg13g2_and2_1 _2834_ (.A(_0288_),
    .B(_0799_),
    .X(_0176_));
 sg13g2_and2_1 _2835_ (.A(\control_tone_freq[2][8] ),
    .B(_0759_),
    .X(_0800_));
 sg13g2_nor2_1 _2836_ (.A(\tone[2].gen.counter[8] ),
    .B(_0800_),
    .Y(_0801_));
 sg13g2_mux2_1 _2837_ (.A0(_0800_),
    .A1(_0801_),
    .S(_0796_),
    .X(_0802_));
 sg13g2_nand2_1 _2838_ (.Y(_0803_),
    .A(_0301_),
    .B(_0796_));
 sg13g2_a22oi_1 _2839_ (.Y(_0804_),
    .B1(_0803_),
    .B2(\tone[2].gen.counter[8] ),
    .A2(_0802_),
    .A1(_0646_));
 sg13g2_nor2_1 _2840_ (.A(_0980_),
    .B(_0804_),
    .Y(_0177_));
 sg13g2_nor3_1 _2841_ (.A(\tone[2].gen.counter[8] ),
    .B(_0800_),
    .C(_0803_),
    .Y(_0805_));
 sg13g2_and2_1 _2842_ (.A(_0301_),
    .B(net30),
    .X(_0806_));
 sg13g2_a21oi_1 _2843_ (.A1(\control_tone_freq[2][9] ),
    .A2(_0806_),
    .Y(_0807_),
    .B1(\tone[2].gen.counter[9] ));
 sg13g2_xor2_1 _2844_ (.B(_0807_),
    .A(_0805_),
    .X(_0808_));
 sg13g2_nor2_1 _2845_ (.A(_0980_),
    .B(_0808_),
    .Y(_0178_));
 sg13g2_nand2_1 _2846_ (.Y(_0809_),
    .A(_0002_),
    .B(_0806_));
 sg13g2_nand2b_1 _2847_ (.Y(_0810_),
    .B(_0812_),
    .A_N(_0806_));
 sg13g2_a21oi_1 _2848_ (.A1(_0809_),
    .A2(_0810_),
    .Y(_0179_),
    .B1(_0859_));
 sg13g2_inv_1 _2849_ (.Y(net13),
    .A(_0543_));
 sg13g2_nor2_1 _2850_ (.A(_0547_),
    .B(_0548_),
    .Y(net14));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _2856__86 (.L_HI(net86));
 sg13g2_buf_1 _2853_ (.A(net80),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2854_ (.A(net81),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2855_ (.A(net82),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2856_ (.A(net86),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2857_ (.A(net87),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2858_ (.A(net88),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2859_ (.A(net89),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2860_ (.A(net90),
    .X(uio_oe[7]));
 sg13g2_buf_1 _2861_ (.A(net83),
    .X(uio_out[0]));
 sg13g2_buf_1 _2862_ (.A(net84),
    .X(uio_out[1]));
 sg13g2_buf_1 _2863_ (.A(net85),
    .X(uio_out[2]));
 sg13g2_buf_1 _2864_ (.A(\genblk4[0].pwm.accumulator[10] ),
    .X(net8));
 sg13g2_buf_1 _2865_ (.A(\genblk4[1].pwm.accumulator[10] ),
    .X(net9));
 sg13g2_buf_1 _2866_ (.A(\genblk4[2].pwm.accumulator[10] ),
    .X(net10));
 sg13g2_buf_1 _2867_ (.A(\genblk4[3].pwm.accumulator[10] ),
    .X(net11));
 sg13g2_buf_1 _2868_ (.A(\pwm.accumulator[12] ),
    .X(net12));
 sg13g2_dfrbp_1 \clk_counter[0]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net91),
    .D(_0007_),
    .Q_N(_0005_),
    .Q(\clk_counter[0] ));
 sg13g2_dfrbp_1 \clk_counter[1]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net92),
    .D(_0008_),
    .Q_N(_1506_),
    .Q(\clk_counter[1] ));
 sg13g2_dfrbp_1 \clk_counter[2]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net93),
    .D(_0009_),
    .Q_N(_1505_),
    .Q(\clk_counter[2] ));
 sg13g2_dfrbp_1 \clk_counter[3]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net94),
    .D(_0010_),
    .Q_N(_1504_),
    .Q(\clk_counter[3] ));
 sg13g2_dfrbp_1 \clk_counter[4]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net95),
    .D(_0011_),
    .Q_N(_1503_),
    .Q(\clk_counter[4] ));
 sg13g2_dfrbp_1 \clk_counter[5]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net96),
    .D(_0012_),
    .Q_N(_1502_),
    .Q(\clk_counter[5] ));
 sg13g2_dfrbp_1 \clk_counter[6]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net97),
    .D(_0013_),
    .Q_N(_1501_),
    .Q(\clk_counter[6] ));
 sg13g2_dfrbp_1 \control_attn[0][0]$_SDFFE_PN1P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net98),
    .D(_0014_),
    .Q_N(_1500_),
    .Q(\chan[0].attenuation.control[0] ));
 sg13g2_dfrbp_1 \control_attn[0][1]$_SDFFE_PN1P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net99),
    .D(_0015_),
    .Q_N(_1499_),
    .Q(\chan[0].attenuation.control[1] ));
 sg13g2_dfrbp_1 \control_attn[0][2]$_SDFFE_PN1P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net100),
    .D(_0016_),
    .Q_N(_1498_),
    .Q(\chan[0].attenuation.control[2] ));
 sg13g2_dfrbp_1 \control_attn[0][3]$_SDFFE_PN1P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net101),
    .D(_0017_),
    .Q_N(_1497_),
    .Q(\chan[0].attenuation.control[3] ));
 sg13g2_dfrbp_1 \control_attn[1][0]$_SDFFE_PN1P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net102),
    .D(_0018_),
    .Q_N(_1496_),
    .Q(\chan[1].attenuation.control[0] ));
 sg13g2_dfrbp_1 \control_attn[1][1]$_SDFFE_PN1P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net103),
    .D(_0019_),
    .Q_N(_1495_),
    .Q(\chan[1].attenuation.control[1] ));
 sg13g2_dfrbp_1 \control_attn[1][2]$_SDFFE_PN1P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net104),
    .D(_0020_),
    .Q_N(_1494_),
    .Q(\chan[1].attenuation.control[2] ));
 sg13g2_dfrbp_1 \control_attn[1][3]$_SDFFE_PN1P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net105),
    .D(_0021_),
    .Q_N(_1493_),
    .Q(\chan[1].attenuation.control[3] ));
 sg13g2_dfrbp_1 \control_attn[2][0]$_SDFFE_PN1P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net106),
    .D(_0022_),
    .Q_N(_1492_),
    .Q(\chan[2].attenuation.control[0] ));
 sg13g2_dfrbp_1 \control_attn[2][1]$_SDFFE_PN1P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net107),
    .D(_0023_),
    .Q_N(_1491_),
    .Q(\chan[2].attenuation.control[1] ));
 sg13g2_dfrbp_1 \control_attn[2][2]$_SDFFE_PN1P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net108),
    .D(_0024_),
    .Q_N(_1490_),
    .Q(\chan[2].attenuation.control[2] ));
 sg13g2_dfrbp_1 \control_attn[2][3]$_SDFFE_PN1P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net109),
    .D(_0025_),
    .Q_N(_1489_),
    .Q(\chan[2].attenuation.control[3] ));
 sg13g2_dfrbp_1 \control_attn[3][0]$_SDFFE_PN1P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net110),
    .D(_0026_),
    .Q_N(_1488_),
    .Q(\chan[3].attenuation.control[0] ));
 sg13g2_dfrbp_1 \control_attn[3][1]$_SDFFE_PN1P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net111),
    .D(_0027_),
    .Q_N(_1487_),
    .Q(\chan[3].attenuation.control[1] ));
 sg13g2_dfrbp_1 \control_attn[3][2]$_SDFFE_PN1P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net112),
    .D(_0028_),
    .Q_N(_1486_),
    .Q(\chan[3].attenuation.control[2] ));
 sg13g2_dfrbp_1 \control_attn[3][3]$_SDFFE_PN1P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net113),
    .D(_0029_),
    .Q_N(_1485_),
    .Q(\chan[3].attenuation.control[3] ));
 sg13g2_dfrbp_1 \control_noise[0][0]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net114),
    .D(_0030_),
    .Q_N(_1484_),
    .Q(\control_noise[0][0] ));
 sg13g2_dfrbp_1 \control_noise[0][1]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net115),
    .D(_0031_),
    .Q_N(_1483_),
    .Q(\control_noise[0][1] ));
 sg13g2_dfrbp_1 \control_noise[0][2]$_SDFFE_PN1P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net116),
    .D(_0032_),
    .Q_N(_1482_),
    .Q(\control_noise[0][2] ));
 sg13g2_dfrbp_1 \control_tone_freq[0][0]$_SDFFE_PN1P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net117),
    .D(_0033_),
    .Q_N(_1481_),
    .Q(\control_tone_freq[0][0] ));
 sg13g2_dfrbp_1 \control_tone_freq[0][1]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net118),
    .D(_0034_),
    .Q_N(_1480_),
    .Q(\control_tone_freq[0][1] ));
 sg13g2_dfrbp_1 \control_tone_freq[0][2]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net119),
    .D(_0035_),
    .Q_N(_1479_),
    .Q(\control_tone_freq[0][2] ));
 sg13g2_dfrbp_1 \control_tone_freq[0][3]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net120),
    .D(_0036_),
    .Q_N(_1478_),
    .Q(\control_tone_freq[0][3] ));
 sg13g2_dfrbp_1 \control_tone_freq[0][4]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net121),
    .D(_0037_),
    .Q_N(_1477_),
    .Q(\control_tone_freq[0][4] ));
 sg13g2_dfrbp_1 \control_tone_freq[0][5]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net122),
    .D(_0038_),
    .Q_N(_1476_),
    .Q(\control_tone_freq[0][5] ));
 sg13g2_dfrbp_1 \control_tone_freq[0][6]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net123),
    .D(_0039_),
    .Q_N(_1475_),
    .Q(\control_tone_freq[0][6] ));
 sg13g2_dfrbp_1 \control_tone_freq[0][7]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net124),
    .D(_0040_),
    .Q_N(_1474_),
    .Q(\control_tone_freq[0][7] ));
 sg13g2_dfrbp_1 \control_tone_freq[0][8]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net125),
    .D(_0041_),
    .Q_N(_1473_),
    .Q(\control_tone_freq[0][8] ));
 sg13g2_dfrbp_1 \control_tone_freq[0][9]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net126),
    .D(_0042_),
    .Q_N(_1472_),
    .Q(\control_tone_freq[0][9] ));
 sg13g2_dfrbp_1 \control_tone_freq[1][0]$_SDFFE_PN1P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net127),
    .D(_0043_),
    .Q_N(_1471_),
    .Q(\control_tone_freq[1][0] ));
 sg13g2_dfrbp_1 \control_tone_freq[1][1]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net128),
    .D(_0044_),
    .Q_N(_1470_),
    .Q(\control_tone_freq[1][1] ));
 sg13g2_dfrbp_1 \control_tone_freq[1][2]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net129),
    .D(_0045_),
    .Q_N(_1469_),
    .Q(\control_tone_freq[1][2] ));
 sg13g2_dfrbp_1 \control_tone_freq[1][3]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net130),
    .D(_0046_),
    .Q_N(_1468_),
    .Q(\control_tone_freq[1][3] ));
 sg13g2_dfrbp_1 \control_tone_freq[1][4]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net131),
    .D(_0047_),
    .Q_N(_1467_),
    .Q(\control_tone_freq[1][4] ));
 sg13g2_dfrbp_1 \control_tone_freq[1][5]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net132),
    .D(_0048_),
    .Q_N(_1466_),
    .Q(\control_tone_freq[1][5] ));
 sg13g2_dfrbp_1 \control_tone_freq[1][6]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net133),
    .D(_0049_),
    .Q_N(_1465_),
    .Q(\control_tone_freq[1][6] ));
 sg13g2_dfrbp_1 \control_tone_freq[1][7]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net134),
    .D(_0050_),
    .Q_N(_1464_),
    .Q(\control_tone_freq[1][7] ));
 sg13g2_dfrbp_1 \control_tone_freq[1][8]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net135),
    .D(_0051_),
    .Q_N(_1463_),
    .Q(\control_tone_freq[1][8] ));
 sg13g2_dfrbp_1 \control_tone_freq[1][9]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net136),
    .D(_0052_),
    .Q_N(_1462_),
    .Q(\control_tone_freq[1][9] ));
 sg13g2_dfrbp_1 \control_tone_freq[2][0]$_SDFFE_PN1P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net137),
    .D(_0053_),
    .Q_N(_1461_),
    .Q(\control_tone_freq[2][0] ));
 sg13g2_dfrbp_1 \control_tone_freq[2][1]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net138),
    .D(_0054_),
    .Q_N(_1460_),
    .Q(\control_tone_freq[2][1] ));
 sg13g2_dfrbp_1 \control_tone_freq[2][2]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net139),
    .D(_0055_),
    .Q_N(_1459_),
    .Q(\control_tone_freq[2][2] ));
 sg13g2_dfrbp_1 \control_tone_freq[2][3]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net140),
    .D(_0056_),
    .Q_N(_1458_),
    .Q(\control_tone_freq[2][3] ));
 sg13g2_dfrbp_1 \control_tone_freq[2][4]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net141),
    .D(_0057_),
    .Q_N(_1457_),
    .Q(\control_tone_freq[2][4] ));
 sg13g2_dfrbp_1 \control_tone_freq[2][5]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net142),
    .D(_0058_),
    .Q_N(_1456_),
    .Q(\control_tone_freq[2][5] ));
 sg13g2_dfrbp_1 \control_tone_freq[2][6]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net143),
    .D(_0059_),
    .Q_N(_1455_),
    .Q(\control_tone_freq[2][6] ));
 sg13g2_dfrbp_1 \control_tone_freq[2][7]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net144),
    .D(_0060_),
    .Q_N(_1454_),
    .Q(\control_tone_freq[2][7] ));
 sg13g2_dfrbp_1 \control_tone_freq[2][8]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net145),
    .D(_0061_),
    .Q_N(_1453_),
    .Q(\control_tone_freq[2][8] ));
 sg13g2_dfrbp_1 \control_tone_freq[2][9]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net146),
    .D(_0062_),
    .Q_N(_1452_),
    .Q(\control_tone_freq[2][9] ));
 sg13g2_dfrbp_1 \genblk4[0].pwm.accumulator[0]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net147),
    .D(_0063_),
    .Q_N(_1451_),
    .Q(\genblk4[0].pwm.accumulator[0] ));
 sg13g2_dfrbp_1 \genblk4[0].pwm.accumulator[10]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net148),
    .D(_0064_),
    .Q_N(_1450_),
    .Q(\genblk4[0].pwm.accumulator[10] ));
 sg13g2_dfrbp_1 \genblk4[0].pwm.accumulator[1]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net149),
    .D(_0065_),
    .Q_N(_1449_),
    .Q(\genblk4[0].pwm.accumulator[1] ));
 sg13g2_dfrbp_1 \genblk4[0].pwm.accumulator[2]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net150),
    .D(_0066_),
    .Q_N(_1448_),
    .Q(\genblk4[0].pwm.accumulator[2] ));
 sg13g2_dfrbp_1 \genblk4[0].pwm.accumulator[3]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net151),
    .D(_0067_),
    .Q_N(_1447_),
    .Q(\genblk4[0].pwm.accumulator[3] ));
 sg13g2_dfrbp_1 \genblk4[0].pwm.accumulator[4]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net152),
    .D(_0068_),
    .Q_N(_1446_),
    .Q(\genblk4[0].pwm.accumulator[4] ));
 sg13g2_dfrbp_1 \genblk4[0].pwm.accumulator[5]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net153),
    .D(_0069_),
    .Q_N(_1445_),
    .Q(\genblk4[0].pwm.accumulator[5] ));
 sg13g2_dfrbp_1 \genblk4[0].pwm.accumulator[6]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net154),
    .D(_0070_),
    .Q_N(_1444_),
    .Q(\genblk4[0].pwm.accumulator[6] ));
 sg13g2_dfrbp_1 \genblk4[0].pwm.accumulator[7]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net155),
    .D(_0071_),
    .Q_N(_1443_),
    .Q(\genblk4[0].pwm.accumulator[7] ));
 sg13g2_dfrbp_1 \genblk4[0].pwm.accumulator[8]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net156),
    .D(_0072_),
    .Q_N(_1442_),
    .Q(\genblk4[0].pwm.accumulator[8] ));
 sg13g2_dfrbp_1 \genblk4[0].pwm.accumulator[9]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net157),
    .D(_0073_),
    .Q_N(_1441_),
    .Q(\genblk4[0].pwm.accumulator[9] ));
 sg13g2_dfrbp_1 \genblk4[1].pwm.accumulator[0]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net158),
    .D(_0074_),
    .Q_N(_1440_),
    .Q(\genblk4[1].pwm.accumulator[0] ));
 sg13g2_dfrbp_1 \genblk4[1].pwm.accumulator[10]$_SDFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net159),
    .D(_0075_),
    .Q_N(_1439_),
    .Q(\genblk4[1].pwm.accumulator[10] ));
 sg13g2_dfrbp_1 \genblk4[1].pwm.accumulator[1]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net160),
    .D(_0076_),
    .Q_N(_1438_),
    .Q(\genblk4[1].pwm.accumulator[1] ));
 sg13g2_dfrbp_1 \genblk4[1].pwm.accumulator[2]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net161),
    .D(_0077_),
    .Q_N(_1437_),
    .Q(\genblk4[1].pwm.accumulator[2] ));
 sg13g2_dfrbp_1 \genblk4[1].pwm.accumulator[3]$_SDFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net162),
    .D(_0078_),
    .Q_N(_1436_),
    .Q(\genblk4[1].pwm.accumulator[3] ));
 sg13g2_dfrbp_1 \genblk4[1].pwm.accumulator[4]$_SDFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net163),
    .D(_0079_),
    .Q_N(_1435_),
    .Q(\genblk4[1].pwm.accumulator[4] ));
 sg13g2_dfrbp_1 \genblk4[1].pwm.accumulator[5]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net164),
    .D(_0080_),
    .Q_N(_1434_),
    .Q(\genblk4[1].pwm.accumulator[5] ));
 sg13g2_dfrbp_1 \genblk4[1].pwm.accumulator[6]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net165),
    .D(_0081_),
    .Q_N(_1433_),
    .Q(\genblk4[1].pwm.accumulator[6] ));
 sg13g2_dfrbp_1 \genblk4[1].pwm.accumulator[7]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net166),
    .D(_0082_),
    .Q_N(_1432_),
    .Q(\genblk4[1].pwm.accumulator[7] ));
 sg13g2_dfrbp_1 \genblk4[1].pwm.accumulator[8]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net167),
    .D(_0083_),
    .Q_N(_1431_),
    .Q(\genblk4[1].pwm.accumulator[8] ));
 sg13g2_dfrbp_1 \genblk4[1].pwm.accumulator[9]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net168),
    .D(_0084_),
    .Q_N(_1430_),
    .Q(\genblk4[1].pwm.accumulator[9] ));
 sg13g2_dfrbp_1 \genblk4[2].pwm.accumulator[0]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net169),
    .D(_0085_),
    .Q_N(_1429_),
    .Q(\genblk4[2].pwm.accumulator[0] ));
 sg13g2_dfrbp_1 \genblk4[2].pwm.accumulator[10]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net170),
    .D(_0086_),
    .Q_N(_1428_),
    .Q(\genblk4[2].pwm.accumulator[10] ));
 sg13g2_dfrbp_1 \genblk4[2].pwm.accumulator[1]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net171),
    .D(_0087_),
    .Q_N(_1427_),
    .Q(\genblk4[2].pwm.accumulator[1] ));
 sg13g2_dfrbp_1 \genblk4[2].pwm.accumulator[2]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net172),
    .D(_0088_),
    .Q_N(_1426_),
    .Q(\genblk4[2].pwm.accumulator[2] ));
 sg13g2_dfrbp_1 \genblk4[2].pwm.accumulator[3]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net173),
    .D(_0089_),
    .Q_N(_1425_),
    .Q(\genblk4[2].pwm.accumulator[3] ));
 sg13g2_dfrbp_1 \genblk4[2].pwm.accumulator[4]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net174),
    .D(_0090_),
    .Q_N(_1424_),
    .Q(\genblk4[2].pwm.accumulator[4] ));
 sg13g2_dfrbp_1 \genblk4[2].pwm.accumulator[5]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net175),
    .D(_0091_),
    .Q_N(_1423_),
    .Q(\genblk4[2].pwm.accumulator[5] ));
 sg13g2_dfrbp_1 \genblk4[2].pwm.accumulator[6]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net176),
    .D(_0092_),
    .Q_N(_1422_),
    .Q(\genblk4[2].pwm.accumulator[6] ));
 sg13g2_dfrbp_1 \genblk4[2].pwm.accumulator[7]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net177),
    .D(_0093_),
    .Q_N(_1421_),
    .Q(\genblk4[2].pwm.accumulator[7] ));
 sg13g2_dfrbp_1 \genblk4[2].pwm.accumulator[8]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net178),
    .D(_0094_),
    .Q_N(_1420_),
    .Q(\genblk4[2].pwm.accumulator[8] ));
 sg13g2_dfrbp_1 \genblk4[2].pwm.accumulator[9]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net179),
    .D(_0095_),
    .Q_N(_1419_),
    .Q(\genblk4[2].pwm.accumulator[9] ));
 sg13g2_dfrbp_1 \genblk4[3].pwm.accumulator[0]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net180),
    .D(_0096_),
    .Q_N(_1418_),
    .Q(\genblk4[3].pwm.accumulator[0] ));
 sg13g2_dfrbp_1 \genblk4[3].pwm.accumulator[10]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net181),
    .D(_0097_),
    .Q_N(_1417_),
    .Q(\genblk4[3].pwm.accumulator[10] ));
 sg13g2_dfrbp_1 \genblk4[3].pwm.accumulator[1]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net182),
    .D(_0098_),
    .Q_N(_1416_),
    .Q(\genblk4[3].pwm.accumulator[1] ));
 sg13g2_dfrbp_1 \genblk4[3].pwm.accumulator[2]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net183),
    .D(_0099_),
    .Q_N(_1415_),
    .Q(\genblk4[3].pwm.accumulator[2] ));
 sg13g2_dfrbp_1 \genblk4[3].pwm.accumulator[3]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net184),
    .D(_0100_),
    .Q_N(_1414_),
    .Q(\genblk4[3].pwm.accumulator[3] ));
 sg13g2_dfrbp_1 \genblk4[3].pwm.accumulator[4]$_SDFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net185),
    .D(_0101_),
    .Q_N(_1413_),
    .Q(\genblk4[3].pwm.accumulator[4] ));
 sg13g2_dfrbp_1 \genblk4[3].pwm.accumulator[5]$_SDFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net186),
    .D(_0102_),
    .Q_N(_1412_),
    .Q(\genblk4[3].pwm.accumulator[5] ));
 sg13g2_dfrbp_1 \genblk4[3].pwm.accumulator[6]$_SDFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net187),
    .D(_0103_),
    .Q_N(_1411_),
    .Q(\genblk4[3].pwm.accumulator[6] ));
 sg13g2_dfrbp_1 \genblk4[3].pwm.accumulator[7]$_SDFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net188),
    .D(_0104_),
    .Q_N(_1410_),
    .Q(\genblk4[3].pwm.accumulator[7] ));
 sg13g2_dfrbp_1 \genblk4[3].pwm.accumulator[8]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net189),
    .D(_0105_),
    .Q_N(_1409_),
    .Q(\genblk4[3].pwm.accumulator[8] ));
 sg13g2_dfrbp_1 \genblk4[3].pwm.accumulator[9]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net190),
    .D(_0106_),
    .Q_N(_1408_),
    .Q(\genblk4[3].pwm.accumulator[9] ));
 sg13g2_dfrbp_1 \latch_control_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net191),
    .D(_0107_),
    .Q_N(_1407_),
    .Q(\latch_control_reg[0] ));
 sg13g2_dfrbp_1 \latch_control_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net192),
    .D(_0108_),
    .Q_N(_1406_),
    .Q(\latch_control_reg[1] ));
 sg13g2_dfrbp_1 \latch_control_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net193),
    .D(_0109_),
    .Q_N(_0003_),
    .Q(\latch_control_reg[2] ));
 sg13g2_dfrbp_1 \noise[0].gen.counter[0]$_SDFFE_PN0N_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net194),
    .D(_0110_),
    .Q_N(_0006_),
    .Q(\noise[0].gen.counter[0] ));
 sg13g2_dfrbp_1 \noise[0].gen.counter[1]$_SDFFE_PN0N_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net195),
    .D(_0111_),
    .Q_N(_1405_),
    .Q(\noise[0].gen.counter[1] ));
 sg13g2_dfrbp_1 \noise[0].gen.counter[2]$_SDFFE_PN0N_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net196),
    .D(_0112_),
    .Q_N(_1404_),
    .Q(\noise[0].gen.counter[2] ));
 sg13g2_dfrbp_1 \noise[0].gen.counter[3]$_SDFFE_PN0N_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net197),
    .D(_0113_),
    .Q_N(_1403_),
    .Q(\noise[0].gen.counter[3] ));
 sg13g2_dfrbp_1 \noise[0].gen.counter[4]$_SDFFE_PN0N_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net198),
    .D(_0114_),
    .Q_N(_0004_),
    .Q(\noise[0].gen.counter[4] ));
 sg13g2_dfrbp_1 \noise[0].gen.counter[5]$_SDFFE_PN0N_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net199),
    .D(_0115_),
    .Q_N(_1402_),
    .Q(\noise[0].gen.counter[5] ));
 sg13g2_dfrbp_1 \noise[0].gen.counter[6]$_SDFFE_PN0N_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net200),
    .D(_0116_),
    .Q_N(_1401_),
    .Q(\noise[0].gen.counter[6] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[0]$_SDFFE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net201),
    .D(_0117_),
    .Q_N(_1400_),
    .Q(\chan[3].attenuation.in ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[10]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net202),
    .D(_0118_),
    .Q_N(_1399_),
    .Q(\noise[0].gen.lfsr[10] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[11]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net203),
    .D(_0119_),
    .Q_N(_1398_),
    .Q(\noise[0].gen.lfsr[11] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[12]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net204),
    .D(_0120_),
    .Q_N(_1397_),
    .Q(\noise[0].gen.lfsr[12] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[13]$_SDFFE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net205),
    .D(_0121_),
    .Q_N(_1396_),
    .Q(\noise[0].gen.lfsr[13] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[14]$_SDFFE_PP1P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net206),
    .D(_0122_),
    .Q_N(_1395_),
    .Q(\noise[0].gen.lfsr[14] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[1]$_SDFFE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net207),
    .D(_0123_),
    .Q_N(_1394_),
    .Q(\noise[0].gen.lfsr[1] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[2]$_SDFFE_PP0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net208),
    .D(_0124_),
    .Q_N(_1393_),
    .Q(\noise[0].gen.lfsr[2] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[3]$_SDFFE_PP0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net209),
    .D(_0125_),
    .Q_N(_1392_),
    .Q(\noise[0].gen.lfsr[3] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[4]$_SDFFE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net210),
    .D(_0126_),
    .Q_N(_1391_),
    .Q(\noise[0].gen.lfsr[4] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[5]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net211),
    .D(_0127_),
    .Q_N(_1390_),
    .Q(\noise[0].gen.lfsr[5] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[6]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net212),
    .D(_0128_),
    .Q_N(_1389_),
    .Q(\noise[0].gen.lfsr[6] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[7]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net213),
    .D(_0129_),
    .Q_N(_1388_),
    .Q(\noise[0].gen.lfsr[7] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[8]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net214),
    .D(_0130_),
    .Q_N(_1387_),
    .Q(\noise[0].gen.lfsr[8] ));
 sg13g2_dfrbp_1 \noise[0].gen.lfsr[9]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net215),
    .D(_0131_),
    .Q_N(_1386_),
    .Q(\noise[0].gen.lfsr[9] ));
 sg13g2_dfrbp_1 \noise[0].gen.signal_edge.previous_signal_state_0$_SDFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net216),
    .D(_0132_),
    .Q_N(_1385_),
    .Q(\noise[0].gen.signal_edge.previous_signal_state_0 ));
 sg13g2_dfrbp_1 \pwm.accumulator[0]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net217),
    .D(_0133_),
    .Q_N(_1384_),
    .Q(\pwm.accumulator[0] ));
 sg13g2_dfrbp_1 \pwm.accumulator[10]$_SDFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net218),
    .D(_0134_),
    .Q_N(_1383_),
    .Q(\pwm.accumulator[10] ));
 sg13g2_dfrbp_1 \pwm.accumulator[11]$_SDFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net219),
    .D(_0135_),
    .Q_N(_1382_),
    .Q(\pwm.accumulator[11] ));
 sg13g2_dfrbp_1 \pwm.accumulator[12]$_SDFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net220),
    .D(_0136_),
    .Q_N(_1381_),
    .Q(\pwm.accumulator[12] ));
 sg13g2_dfrbp_1 \pwm.accumulator[1]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net221),
    .D(_0137_),
    .Q_N(_1380_),
    .Q(\pwm.accumulator[1] ));
 sg13g2_dfrbp_1 \pwm.accumulator[2]$_SDFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net222),
    .D(_0138_),
    .Q_N(_1379_),
    .Q(\pwm.accumulator[2] ));
 sg13g2_dfrbp_1 \pwm.accumulator[3]$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net223),
    .D(_0139_),
    .Q_N(_1378_),
    .Q(\pwm.accumulator[3] ));
 sg13g2_dfrbp_1 \pwm.accumulator[4]$_SDFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net224),
    .D(_0140_),
    .Q_N(_1377_),
    .Q(\pwm.accumulator[4] ));
 sg13g2_dfrbp_1 \pwm.accumulator[5]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net225),
    .D(_0141_),
    .Q_N(_1376_),
    .Q(\pwm.accumulator[5] ));
 sg13g2_dfrbp_1 \pwm.accumulator[6]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net226),
    .D(_0142_),
    .Q_N(_1375_),
    .Q(\pwm.accumulator[6] ));
 sg13g2_dfrbp_1 \pwm.accumulator[7]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net227),
    .D(_0143_),
    .Q_N(_1374_),
    .Q(\pwm.accumulator[7] ));
 sg13g2_dfrbp_1 \pwm.accumulator[8]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net228),
    .D(_0144_),
    .Q_N(_1373_),
    .Q(\pwm.accumulator[8] ));
 sg13g2_dfrbp_1 \pwm.accumulator[9]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net229),
    .D(_0145_),
    .Q_N(_1372_),
    .Q(\pwm.accumulator[9] ));
 sg13g2_dfrbp_1 \restart_noise$_SDFF_PP0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net230),
    .D(_0146_),
    .Q_N(_1371_),
    .Q(\noise[0].gen.restart_noise ));
 sg13g2_dfrbp_1 \tone[0].gen.counter[0]$_SDFFE_PN0N_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net231),
    .D(_0147_),
    .Q_N(_1370_),
    .Q(\tone[0].gen.counter[0] ));
 sg13g2_dfrbp_1 \tone[0].gen.counter[1]$_SDFFE_PN0N_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net232),
    .D(_0148_),
    .Q_N(_1369_),
    .Q(\tone[0].gen.counter[1] ));
 sg13g2_dfrbp_1 \tone[0].gen.counter[2]$_SDFFE_PN0N_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net233),
    .D(_0149_),
    .Q_N(_1368_),
    .Q(\tone[0].gen.counter[2] ));
 sg13g2_dfrbp_1 \tone[0].gen.counter[3]$_SDFFE_PN0N_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net234),
    .D(_0150_),
    .Q_N(_1367_),
    .Q(\tone[0].gen.counter[3] ));
 sg13g2_dfrbp_1 \tone[0].gen.counter[4]$_SDFFE_PN0N_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net235),
    .D(_0151_),
    .Q_N(_1366_),
    .Q(\tone[0].gen.counter[4] ));
 sg13g2_dfrbp_1 \tone[0].gen.counter[5]$_SDFFE_PN0N_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net236),
    .D(_0152_),
    .Q_N(_1365_),
    .Q(\tone[0].gen.counter[5] ));
 sg13g2_dfrbp_1 \tone[0].gen.counter[6]$_SDFFE_PN0N_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net237),
    .D(_0153_),
    .Q_N(_1364_),
    .Q(\tone[0].gen.counter[6] ));
 sg13g2_dfrbp_1 \tone[0].gen.counter[7]$_SDFFE_PN0N_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net238),
    .D(_0154_),
    .Q_N(_1363_),
    .Q(\tone[0].gen.counter[7] ));
 sg13g2_dfrbp_1 \tone[0].gen.counter[8]$_SDFFE_PN0N_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net239),
    .D(_0155_),
    .Q_N(_1362_),
    .Q(\tone[0].gen.counter[8] ));
 sg13g2_dfrbp_1 \tone[0].gen.counter[9]$_SDFFE_PN0N_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net240),
    .D(_0156_),
    .Q_N(_1361_),
    .Q(\tone[0].gen.counter[9] ));
 sg13g2_dfrbp_1 \tone[0].gen.state$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net241),
    .D(_0157_),
    .Q_N(_0000_),
    .Q(\chan[0].attenuation.in ));
 sg13g2_dfrbp_1 \tone[1].gen.counter[0]$_SDFFE_PN0N_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net242),
    .D(_0158_),
    .Q_N(_1360_),
    .Q(\tone[1].gen.counter[0] ));
 sg13g2_dfrbp_1 \tone[1].gen.counter[1]$_SDFFE_PN0N_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net243),
    .D(_0159_),
    .Q_N(_1359_),
    .Q(\tone[1].gen.counter[1] ));
 sg13g2_dfrbp_1 \tone[1].gen.counter[2]$_SDFFE_PN0N_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net244),
    .D(_0160_),
    .Q_N(_1358_),
    .Q(\tone[1].gen.counter[2] ));
 sg13g2_dfrbp_1 \tone[1].gen.counter[3]$_SDFFE_PN0N_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net245),
    .D(_0161_),
    .Q_N(_1357_),
    .Q(\tone[1].gen.counter[3] ));
 sg13g2_dfrbp_1 \tone[1].gen.counter[4]$_SDFFE_PN0N_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net246),
    .D(_0162_),
    .Q_N(_1356_),
    .Q(\tone[1].gen.counter[4] ));
 sg13g2_dfrbp_1 \tone[1].gen.counter[5]$_SDFFE_PN0N_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net247),
    .D(_0163_),
    .Q_N(_1355_),
    .Q(\tone[1].gen.counter[5] ));
 sg13g2_dfrbp_1 \tone[1].gen.counter[6]$_SDFFE_PN0N_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net248),
    .D(_0164_),
    .Q_N(_1354_),
    .Q(\tone[1].gen.counter[6] ));
 sg13g2_dfrbp_1 \tone[1].gen.counter[7]$_SDFFE_PN0N_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net249),
    .D(_0165_),
    .Q_N(_1353_),
    .Q(\tone[1].gen.counter[7] ));
 sg13g2_dfrbp_1 \tone[1].gen.counter[8]$_SDFFE_PN0N_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net250),
    .D(_0166_),
    .Q_N(_1352_),
    .Q(\tone[1].gen.counter[8] ));
 sg13g2_dfrbp_1 \tone[1].gen.counter[9]$_SDFFE_PN0N_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net251),
    .D(_0167_),
    .Q_N(_1351_),
    .Q(\tone[1].gen.counter[9] ));
 sg13g2_dfrbp_1 \tone[1].gen.state$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net252),
    .D(_0168_),
    .Q_N(_0001_),
    .Q(\chan[1].attenuation.in ));
 sg13g2_dfrbp_1 \tone[2].gen.counter[0]$_SDFFE_PN0N_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net253),
    .D(_0169_),
    .Q_N(_1350_),
    .Q(\tone[2].gen.counter[0] ));
 sg13g2_dfrbp_1 \tone[2].gen.counter[1]$_SDFFE_PN0N_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net254),
    .D(_0170_),
    .Q_N(_1349_),
    .Q(\tone[2].gen.counter[1] ));
 sg13g2_dfrbp_1 \tone[2].gen.counter[2]$_SDFFE_PN0N_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net255),
    .D(_0171_),
    .Q_N(_1348_),
    .Q(\tone[2].gen.counter[2] ));
 sg13g2_dfrbp_1 \tone[2].gen.counter[3]$_SDFFE_PN0N_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net256),
    .D(_0172_),
    .Q_N(_1347_),
    .Q(\tone[2].gen.counter[3] ));
 sg13g2_dfrbp_1 \tone[2].gen.counter[4]$_SDFFE_PN0N_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net257),
    .D(_0173_),
    .Q_N(_1346_),
    .Q(\tone[2].gen.counter[4] ));
 sg13g2_dfrbp_1 \tone[2].gen.counter[5]$_SDFFE_PN0N_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net258),
    .D(_0174_),
    .Q_N(_1345_),
    .Q(\tone[2].gen.counter[5] ));
 sg13g2_dfrbp_1 \tone[2].gen.counter[6]$_SDFFE_PN0N_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net259),
    .D(_0175_),
    .Q_N(_1344_),
    .Q(\tone[2].gen.counter[6] ));
 sg13g2_dfrbp_1 \tone[2].gen.counter[7]$_SDFFE_PN0N_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net260),
    .D(_0176_),
    .Q_N(_1343_),
    .Q(\tone[2].gen.counter[7] ));
 sg13g2_dfrbp_1 \tone[2].gen.counter[8]$_SDFFE_PN0N_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net261),
    .D(_0177_),
    .Q_N(_1342_),
    .Q(\tone[2].gen.counter[8] ));
 sg13g2_dfrbp_1 \tone[2].gen.counter[9]$_SDFFE_PN0N_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net262),
    .D(_0178_),
    .Q_N(_1341_),
    .Q(\tone[2].gen.counter[9] ));
 sg13g2_dfrbp_1 \tone[2].gen.state$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net263),
    .D(_0179_),
    .Q_N(_0002_),
    .Q(\chan[2].attenuation.in ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[6]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[7]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[1]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[2]),
    .X(net7));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[3]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[4]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[5]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[6]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[7]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[0]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[1]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[2]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[3]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[4]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[5]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[6]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout21 (.A(_0494_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0456_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0656_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0646_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0307_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0303_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0195_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0821_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0816_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0759_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0702_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0642_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0306_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0302_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0988_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1126_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0860_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0826_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0680_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0611_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0292_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1340_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1234_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1026_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0985_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0980_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0967_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0963_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0959_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0949_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0945_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0941_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0935_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0924_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0920_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0916_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0907_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0902_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0859_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0288_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1148_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1040_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1033_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0955_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0944_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0939_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0927_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0897_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0892_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0883_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0882_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0869_),
    .X(net72));
 sg13g2_buf_1 fanout73 (.A(_0858_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0818_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0812_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0909_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0904_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0899_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0894_),
    .X(net79));
 sg13g2_tielo _2853__80 (.L_LO(net80));
 sg13g2_tielo _2854__81 (.L_LO(net81));
 sg13g2_tielo _2855__82 (.L_LO(net82));
 sg13g2_tielo _2861__83 (.L_LO(net83));
 sg13g2_tielo _2862__84 (.L_LO(net84));
 sg13g2_tielo _2863__85 (.L_LO(net85));
 sg13g2_tiehi _2857__87 (.L_HI(net87));
 sg13g2_tiehi _2858__88 (.L_HI(net88));
 sg13g2_tiehi _2859__89 (.L_HI(net89));
 sg13g2_tiehi _2860__90 (.L_HI(net90));
 sg13g2_tiehi \clk_counter[0]$_SDFF_PN0__91  (.L_HI(net91));
 sg13g2_tiehi \clk_counter[1]$_SDFF_PN0__92  (.L_HI(net92));
 sg13g2_tiehi \clk_counter[2]$_SDFF_PN0__93  (.L_HI(net93));
 sg13g2_tiehi \clk_counter[3]$_SDFF_PN0__94  (.L_HI(net94));
 sg13g2_tiehi \clk_counter[4]$_SDFF_PN0__95  (.L_HI(net95));
 sg13g2_tiehi \clk_counter[5]$_SDFF_PN0__96  (.L_HI(net96));
 sg13g2_tiehi \clk_counter[6]$_SDFF_PN0__97  (.L_HI(net97));
 sg13g2_tiehi \control_attn[0][0]$_SDFFE_PN1P__98  (.L_HI(net98));
 sg13g2_tiehi \control_attn[0][1]$_SDFFE_PN1P__99  (.L_HI(net99));
 sg13g2_tiehi \control_attn[0][2]$_SDFFE_PN1P__100  (.L_HI(net100));
 sg13g2_tiehi \control_attn[0][3]$_SDFFE_PN1P__101  (.L_HI(net101));
 sg13g2_tiehi \control_attn[1][0]$_SDFFE_PN1P__102  (.L_HI(net102));
 sg13g2_tiehi \control_attn[1][1]$_SDFFE_PN1P__103  (.L_HI(net103));
 sg13g2_tiehi \control_attn[1][2]$_SDFFE_PN1P__104  (.L_HI(net104));
 sg13g2_tiehi \control_attn[1][3]$_SDFFE_PN1P__105  (.L_HI(net105));
 sg13g2_tiehi \control_attn[2][0]$_SDFFE_PN1P__106  (.L_HI(net106));
 sg13g2_tiehi \control_attn[2][1]$_SDFFE_PN1P__107  (.L_HI(net107));
 sg13g2_tiehi \control_attn[2][2]$_SDFFE_PN1P__108  (.L_HI(net108));
 sg13g2_tiehi \control_attn[2][3]$_SDFFE_PN1P__109  (.L_HI(net109));
 sg13g2_tiehi \control_attn[3][0]$_SDFFE_PN1P__110  (.L_HI(net110));
 sg13g2_tiehi \control_attn[3][1]$_SDFFE_PN1P__111  (.L_HI(net111));
 sg13g2_tiehi \control_attn[3][2]$_SDFFE_PN1P__112  (.L_HI(net112));
 sg13g2_tiehi \control_attn[3][3]$_SDFFE_PN1P__113  (.L_HI(net113));
 sg13g2_tiehi \control_noise[0][0]$_SDFFE_PN0P__114  (.L_HI(net114));
 sg13g2_tiehi \control_noise[0][1]$_SDFFE_PN0P__115  (.L_HI(net115));
 sg13g2_tiehi \control_noise[0][2]$_SDFFE_PN1P__116  (.L_HI(net116));
 sg13g2_tiehi \control_tone_freq[0][0]$_SDFFE_PN1P__117  (.L_HI(net117));
 sg13g2_tiehi \control_tone_freq[0][1]$_SDFFE_PN0P__118  (.L_HI(net118));
 sg13g2_tiehi \control_tone_freq[0][2]$_SDFFE_PN0P__119  (.L_HI(net119));
 sg13g2_tiehi \control_tone_freq[0][3]$_SDFFE_PN0P__120  (.L_HI(net120));
 sg13g2_tiehi \control_tone_freq[0][4]$_SDFFE_PN0P__121  (.L_HI(net121));
 sg13g2_tiehi \control_tone_freq[0][5]$_SDFFE_PN0P__122  (.L_HI(net122));
 sg13g2_tiehi \control_tone_freq[0][6]$_SDFFE_PN0P__123  (.L_HI(net123));
 sg13g2_tiehi \control_tone_freq[0][7]$_SDFFE_PN0P__124  (.L_HI(net124));
 sg13g2_tiehi \control_tone_freq[0][8]$_SDFFE_PN0P__125  (.L_HI(net125));
 sg13g2_tiehi \control_tone_freq[0][9]$_SDFFE_PN0P__126  (.L_HI(net126));
 sg13g2_tiehi \control_tone_freq[1][0]$_SDFFE_PN1P__127  (.L_HI(net127));
 sg13g2_tiehi \control_tone_freq[1][1]$_SDFFE_PN0P__128  (.L_HI(net128));
 sg13g2_tiehi \control_tone_freq[1][2]$_SDFFE_PN0P__129  (.L_HI(net129));
 sg13g2_tiehi \control_tone_freq[1][3]$_SDFFE_PN0P__130  (.L_HI(net130));
 sg13g2_tiehi \control_tone_freq[1][4]$_SDFFE_PN0P__131  (.L_HI(net131));
 sg13g2_tiehi \control_tone_freq[1][5]$_SDFFE_PN0P__132  (.L_HI(net132));
 sg13g2_tiehi \control_tone_freq[1][6]$_SDFFE_PN0P__133  (.L_HI(net133));
 sg13g2_tiehi \control_tone_freq[1][7]$_SDFFE_PN0P__134  (.L_HI(net134));
 sg13g2_tiehi \control_tone_freq[1][8]$_SDFFE_PN0P__135  (.L_HI(net135));
 sg13g2_tiehi \control_tone_freq[1][9]$_SDFFE_PN0P__136  (.L_HI(net136));
 sg13g2_tiehi \control_tone_freq[2][0]$_SDFFE_PN1P__137  (.L_HI(net137));
 sg13g2_tiehi \control_tone_freq[2][1]$_SDFFE_PN0P__138  (.L_HI(net138));
 sg13g2_tiehi \control_tone_freq[2][2]$_SDFFE_PN0P__139  (.L_HI(net139));
 sg13g2_tiehi \control_tone_freq[2][3]$_SDFFE_PN0P__140  (.L_HI(net140));
 sg13g2_tiehi \control_tone_freq[2][4]$_SDFFE_PN0P__141  (.L_HI(net141));
 sg13g2_tiehi \control_tone_freq[2][5]$_SDFFE_PN0P__142  (.L_HI(net142));
 sg13g2_tiehi \control_tone_freq[2][6]$_SDFFE_PN0P__143  (.L_HI(net143));
 sg13g2_tiehi \control_tone_freq[2][7]$_SDFFE_PN0P__144  (.L_HI(net144));
 sg13g2_tiehi \control_tone_freq[2][8]$_SDFFE_PN0P__145  (.L_HI(net145));
 sg13g2_tiehi \control_tone_freq[2][9]$_SDFFE_PN0P__146  (.L_HI(net146));
 sg13g2_tiehi \genblk4[0].pwm.accumulator[0]$_SDFF_PN0__147  (.L_HI(net147));
 sg13g2_tiehi \genblk4[0].pwm.accumulator[10]$_SDFF_PN0__148  (.L_HI(net148));
 sg13g2_tiehi \genblk4[0].pwm.accumulator[1]$_SDFF_PN0__149  (.L_HI(net149));
 sg13g2_tiehi \genblk4[0].pwm.accumulator[2]$_SDFF_PN0__150  (.L_HI(net150));
 sg13g2_tiehi \genblk4[0].pwm.accumulator[3]$_SDFF_PN0__151  (.L_HI(net151));
 sg13g2_tiehi \genblk4[0].pwm.accumulator[4]$_SDFF_PN0__152  (.L_HI(net152));
 sg13g2_tiehi \genblk4[0].pwm.accumulator[5]$_SDFF_PN0__153  (.L_HI(net153));
 sg13g2_tiehi \genblk4[0].pwm.accumulator[6]$_SDFF_PN0__154  (.L_HI(net154));
 sg13g2_tiehi \genblk4[0].pwm.accumulator[7]$_SDFF_PN0__155  (.L_HI(net155));
 sg13g2_tiehi \genblk4[0].pwm.accumulator[8]$_SDFF_PN0__156  (.L_HI(net156));
 sg13g2_tiehi \genblk4[0].pwm.accumulator[9]$_SDFF_PN0__157  (.L_HI(net157));
 sg13g2_tiehi \genblk4[1].pwm.accumulator[0]$_SDFF_PN0__158  (.L_HI(net158));
 sg13g2_tiehi \genblk4[1].pwm.accumulator[10]$_SDFF_PN0__159  (.L_HI(net159));
 sg13g2_tiehi \genblk4[1].pwm.accumulator[1]$_SDFF_PN0__160  (.L_HI(net160));
 sg13g2_tiehi \genblk4[1].pwm.accumulator[2]$_SDFF_PN0__161  (.L_HI(net161));
 sg13g2_tiehi \genblk4[1].pwm.accumulator[3]$_SDFF_PN0__162  (.L_HI(net162));
 sg13g2_tiehi \genblk4[1].pwm.accumulator[4]$_SDFF_PN0__163  (.L_HI(net163));
 sg13g2_tiehi \genblk4[1].pwm.accumulator[5]$_SDFF_PN0__164  (.L_HI(net164));
 sg13g2_tiehi \genblk4[1].pwm.accumulator[6]$_SDFF_PN0__165  (.L_HI(net165));
 sg13g2_tiehi \genblk4[1].pwm.accumulator[7]$_SDFF_PN0__166  (.L_HI(net166));
 sg13g2_tiehi \genblk4[1].pwm.accumulator[8]$_SDFF_PN0__167  (.L_HI(net167));
 sg13g2_tiehi \genblk4[1].pwm.accumulator[9]$_SDFF_PN0__168  (.L_HI(net168));
 sg13g2_tiehi \genblk4[2].pwm.accumulator[0]$_SDFF_PN0__169  (.L_HI(net169));
 sg13g2_tiehi \genblk4[2].pwm.accumulator[10]$_SDFF_PN0__170  (.L_HI(net170));
 sg13g2_tiehi \genblk4[2].pwm.accumulator[1]$_SDFF_PN0__171  (.L_HI(net171));
 sg13g2_tiehi \genblk4[2].pwm.accumulator[2]$_SDFF_PN0__172  (.L_HI(net172));
 sg13g2_tiehi \genblk4[2].pwm.accumulator[3]$_SDFF_PN0__173  (.L_HI(net173));
 sg13g2_tiehi \genblk4[2].pwm.accumulator[4]$_SDFF_PN0__174  (.L_HI(net174));
 sg13g2_tiehi \genblk4[2].pwm.accumulator[5]$_SDFF_PN0__175  (.L_HI(net175));
 sg13g2_tiehi \genblk4[2].pwm.accumulator[6]$_SDFF_PN0__176  (.L_HI(net176));
 sg13g2_tiehi \genblk4[2].pwm.accumulator[7]$_SDFF_PN0__177  (.L_HI(net177));
 sg13g2_tiehi \genblk4[2].pwm.accumulator[8]$_SDFF_PN0__178  (.L_HI(net178));
 sg13g2_tiehi \genblk4[2].pwm.accumulator[9]$_SDFF_PN0__179  (.L_HI(net179));
 sg13g2_tiehi \genblk4[3].pwm.accumulator[0]$_SDFF_PN0__180  (.L_HI(net180));
 sg13g2_tiehi \genblk4[3].pwm.accumulator[10]$_SDFF_PN0__181  (.L_HI(net181));
 sg13g2_tiehi \genblk4[3].pwm.accumulator[1]$_SDFF_PN0__182  (.L_HI(net182));
 sg13g2_tiehi \genblk4[3].pwm.accumulator[2]$_SDFF_PN0__183  (.L_HI(net183));
 sg13g2_tiehi \genblk4[3].pwm.accumulator[3]$_SDFF_PN0__184  (.L_HI(net184));
 sg13g2_tiehi \genblk4[3].pwm.accumulator[4]$_SDFF_PN0__185  (.L_HI(net185));
 sg13g2_tiehi \genblk4[3].pwm.accumulator[5]$_SDFF_PN0__186  (.L_HI(net186));
 sg13g2_tiehi \genblk4[3].pwm.accumulator[6]$_SDFF_PN0__187  (.L_HI(net187));
 sg13g2_tiehi \genblk4[3].pwm.accumulator[7]$_SDFF_PN0__188  (.L_HI(net188));
 sg13g2_tiehi \genblk4[3].pwm.accumulator[8]$_SDFF_PN0__189  (.L_HI(net189));
 sg13g2_tiehi \genblk4[3].pwm.accumulator[9]$_SDFF_PN0__190  (.L_HI(net190));
 sg13g2_tiehi \latch_control_reg[0]$_SDFFE_PN0P__191  (.L_HI(net191));
 sg13g2_tiehi \latch_control_reg[1]$_SDFFE_PN0P__192  (.L_HI(net192));
 sg13g2_tiehi \latch_control_reg[2]$_SDFFE_PN0P__193  (.L_HI(net193));
 sg13g2_tiehi \noise[0].gen.counter[0]$_SDFFE_PN0N__194  (.L_HI(net194));
 sg13g2_tiehi \noise[0].gen.counter[1]$_SDFFE_PN0N__195  (.L_HI(net195));
 sg13g2_tiehi \noise[0].gen.counter[2]$_SDFFE_PN0N__196  (.L_HI(net196));
 sg13g2_tiehi \noise[0].gen.counter[3]$_SDFFE_PN0N__197  (.L_HI(net197));
 sg13g2_tiehi \noise[0].gen.counter[4]$_SDFFE_PN0N__198  (.L_HI(net198));
 sg13g2_tiehi \noise[0].gen.counter[5]$_SDFFE_PN0N__199  (.L_HI(net199));
 sg13g2_tiehi \noise[0].gen.counter[6]$_SDFFE_PN0N__200  (.L_HI(net200));
 sg13g2_tiehi \noise[0].gen.lfsr[0]$_SDFFE_PP0P__201  (.L_HI(net201));
 sg13g2_tiehi \noise[0].gen.lfsr[10]$_SDFFE_PP0P__202  (.L_HI(net202));
 sg13g2_tiehi \noise[0].gen.lfsr[11]$_SDFFE_PP0P__203  (.L_HI(net203));
 sg13g2_tiehi \noise[0].gen.lfsr[12]$_SDFFE_PP0P__204  (.L_HI(net204));
 sg13g2_tiehi \noise[0].gen.lfsr[13]$_SDFFE_PP0P__205  (.L_HI(net205));
 sg13g2_tiehi \noise[0].gen.lfsr[14]$_SDFFE_PP1P__206  (.L_HI(net206));
 sg13g2_tiehi \noise[0].gen.lfsr[1]$_SDFFE_PP0P__207  (.L_HI(net207));
 sg13g2_tiehi \noise[0].gen.lfsr[2]$_SDFFE_PP0P__208  (.L_HI(net208));
 sg13g2_tiehi \noise[0].gen.lfsr[3]$_SDFFE_PP0P__209  (.L_HI(net209));
 sg13g2_tiehi \noise[0].gen.lfsr[4]$_SDFFE_PP0P__210  (.L_HI(net210));
 sg13g2_tiehi \noise[0].gen.lfsr[5]$_SDFFE_PP0P__211  (.L_HI(net211));
 sg13g2_tiehi \noise[0].gen.lfsr[6]$_SDFFE_PP0P__212  (.L_HI(net212));
 sg13g2_tiehi \noise[0].gen.lfsr[7]$_SDFFE_PP0P__213  (.L_HI(net213));
 sg13g2_tiehi \noise[0].gen.lfsr[8]$_SDFFE_PP0P__214  (.L_HI(net214));
 sg13g2_tiehi \noise[0].gen.lfsr[9]$_SDFFE_PP0P__215  (.L_HI(net215));
 sg13g2_tiehi \noise[0].gen.signal_edge.previous_signal_state_0$_SDFF_PN0__216  (.L_HI(net216));
 sg13g2_tiehi \pwm.accumulator[0]$_SDFF_PN0__217  (.L_HI(net217));
 sg13g2_tiehi \pwm.accumulator[10]$_SDFF_PN0__218  (.L_HI(net218));
 sg13g2_tiehi \pwm.accumulator[11]$_SDFF_PN0__219  (.L_HI(net219));
 sg13g2_tiehi \pwm.accumulator[12]$_SDFF_PN0__220  (.L_HI(net220));
 sg13g2_tiehi \pwm.accumulator[1]$_SDFF_PN0__221  (.L_HI(net221));
 sg13g2_tiehi \pwm.accumulator[2]$_SDFF_PN0__222  (.L_HI(net222));
 sg13g2_tiehi \pwm.accumulator[3]$_SDFF_PN0__223  (.L_HI(net223));
 sg13g2_tiehi \pwm.accumulator[4]$_SDFF_PN0__224  (.L_HI(net224));
 sg13g2_tiehi \pwm.accumulator[5]$_SDFF_PN0__225  (.L_HI(net225));
 sg13g2_tiehi \pwm.accumulator[6]$_SDFF_PN0__226  (.L_HI(net226));
 sg13g2_tiehi \pwm.accumulator[7]$_SDFF_PN0__227  (.L_HI(net227));
 sg13g2_tiehi \pwm.accumulator[8]$_SDFF_PN0__228  (.L_HI(net228));
 sg13g2_tiehi \pwm.accumulator[9]$_SDFF_PN0__229  (.L_HI(net229));
 sg13g2_tiehi \restart_noise$_SDFF_PP0__230  (.L_HI(net230));
 sg13g2_tiehi \tone[0].gen.counter[0]$_SDFFE_PN0N__231  (.L_HI(net231));
 sg13g2_tiehi \tone[0].gen.counter[1]$_SDFFE_PN0N__232  (.L_HI(net232));
 sg13g2_tiehi \tone[0].gen.counter[2]$_SDFFE_PN0N__233  (.L_HI(net233));
 sg13g2_tiehi \tone[0].gen.counter[3]$_SDFFE_PN0N__234  (.L_HI(net234));
 sg13g2_tiehi \tone[0].gen.counter[4]$_SDFFE_PN0N__235  (.L_HI(net235));
 sg13g2_tiehi \tone[0].gen.counter[5]$_SDFFE_PN0N__236  (.L_HI(net236));
 sg13g2_tiehi \tone[0].gen.counter[6]$_SDFFE_PN0N__237  (.L_HI(net237));
 sg13g2_tiehi \tone[0].gen.counter[7]$_SDFFE_PN0N__238  (.L_HI(net238));
 sg13g2_tiehi \tone[0].gen.counter[8]$_SDFFE_PN0N__239  (.L_HI(net239));
 sg13g2_tiehi \tone[0].gen.counter[9]$_SDFFE_PN0N__240  (.L_HI(net240));
 sg13g2_tiehi \tone[0].gen.state$_SDFFE_PN0P__241  (.L_HI(net241));
 sg13g2_tiehi \tone[1].gen.counter[0]$_SDFFE_PN0N__242  (.L_HI(net242));
 sg13g2_tiehi \tone[1].gen.counter[1]$_SDFFE_PN0N__243  (.L_HI(net243));
 sg13g2_tiehi \tone[1].gen.counter[2]$_SDFFE_PN0N__244  (.L_HI(net244));
 sg13g2_tiehi \tone[1].gen.counter[3]$_SDFFE_PN0N__245  (.L_HI(net245));
 sg13g2_tiehi \tone[1].gen.counter[4]$_SDFFE_PN0N__246  (.L_HI(net246));
 sg13g2_tiehi \tone[1].gen.counter[5]$_SDFFE_PN0N__247  (.L_HI(net247));
 sg13g2_tiehi \tone[1].gen.counter[6]$_SDFFE_PN0N__248  (.L_HI(net248));
 sg13g2_tiehi \tone[1].gen.counter[7]$_SDFFE_PN0N__249  (.L_HI(net249));
 sg13g2_tiehi \tone[1].gen.counter[8]$_SDFFE_PN0N__250  (.L_HI(net250));
 sg13g2_tiehi \tone[1].gen.counter[9]$_SDFFE_PN0N__251  (.L_HI(net251));
 sg13g2_tiehi \tone[1].gen.state$_SDFFE_PN0P__252  (.L_HI(net252));
 sg13g2_tiehi \tone[2].gen.counter[0]$_SDFFE_PN0N__253  (.L_HI(net253));
 sg13g2_tiehi \tone[2].gen.counter[1]$_SDFFE_PN0N__254  (.L_HI(net254));
 sg13g2_tiehi \tone[2].gen.counter[2]$_SDFFE_PN0N__255  (.L_HI(net255));
 sg13g2_tiehi \tone[2].gen.counter[3]$_SDFFE_PN0N__256  (.L_HI(net256));
 sg13g2_tiehi \tone[2].gen.counter[4]$_SDFFE_PN0N__257  (.L_HI(net257));
 sg13g2_tiehi \tone[2].gen.counter[5]$_SDFFE_PN0N__258  (.L_HI(net258));
 sg13g2_tiehi \tone[2].gen.counter[6]$_SDFFE_PN0N__259  (.L_HI(net259));
 sg13g2_tiehi \tone[2].gen.counter[7]$_SDFFE_PN0N__260  (.L_HI(net260));
 sg13g2_tiehi \tone[2].gen.counter[8]$_SDFFE_PN0N__261  (.L_HI(net261));
 sg13g2_tiehi \tone[2].gen.counter[9]$_SDFFE_PN0N__262  (.L_HI(net262));
 sg13g2_tiehi \tone[2].gen.state$_SDFFE_PN0P__263  (.L_HI(net263));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_29__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_fill_2 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_256 ();
 sg13g2_decap_8 FILLER_1_263 ();
 sg13g2_decap_8 FILLER_1_270 ();
 sg13g2_decap_8 FILLER_1_277 ();
 sg13g2_decap_8 FILLER_1_284 ();
 sg13g2_decap_8 FILLER_1_291 ();
 sg13g2_decap_8 FILLER_1_298 ();
 sg13g2_decap_8 FILLER_1_305 ();
 sg13g2_decap_8 FILLER_1_312 ();
 sg13g2_decap_8 FILLER_1_319 ();
 sg13g2_fill_2 FILLER_1_326 ();
 sg13g2_fill_1 FILLER_1_328 ();
 sg13g2_decap_8 FILLER_1_337 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_decap_8 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_4 FILLER_2_210 ();
 sg13g2_fill_1 FILLER_2_214 ();
 sg13g2_decap_4 FILLER_2_246 ();
 sg13g2_fill_2 FILLER_2_254 ();
 sg13g2_decap_4 FILLER_2_261 ();
 sg13g2_fill_1 FILLER_2_299 ();
 sg13g2_fill_1 FILLER_2_309 ();
 sg13g2_decap_8 FILLER_2_344 ();
 sg13g2_decap_8 FILLER_2_351 ();
 sg13g2_decap_8 FILLER_2_358 ();
 sg13g2_decap_8 FILLER_2_365 ();
 sg13g2_decap_8 FILLER_2_372 ();
 sg13g2_decap_8 FILLER_2_379 ();
 sg13g2_decap_8 FILLER_2_386 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_decap_8 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_2_414 ();
 sg13g2_decap_8 FILLER_2_421 ();
 sg13g2_fill_2 FILLER_2_428 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_fill_1 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_103 ();
 sg13g2_decap_8 FILLER_3_110 ();
 sg13g2_decap_8 FILLER_3_117 ();
 sg13g2_fill_1 FILLER_3_124 ();
 sg13g2_decap_8 FILLER_3_129 ();
 sg13g2_decap_8 FILLER_3_136 ();
 sg13g2_decap_8 FILLER_3_143 ();
 sg13g2_decap_8 FILLER_3_150 ();
 sg13g2_decap_8 FILLER_3_157 ();
 sg13g2_decap_8 FILLER_3_164 ();
 sg13g2_decap_8 FILLER_3_171 ();
 sg13g2_decap_8 FILLER_3_178 ();
 sg13g2_decap_8 FILLER_3_185 ();
 sg13g2_decap_8 FILLER_3_192 ();
 sg13g2_decap_8 FILLER_3_199 ();
 sg13g2_decap_8 FILLER_3_206 ();
 sg13g2_decap_8 FILLER_3_213 ();
 sg13g2_decap_4 FILLER_3_228 ();
 sg13g2_fill_2 FILLER_3_232 ();
 sg13g2_decap_4 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_258 ();
 sg13g2_decap_4 FILLER_3_265 ();
 sg13g2_decap_8 FILLER_3_282 ();
 sg13g2_fill_1 FILLER_3_289 ();
 sg13g2_fill_1 FILLER_3_326 ();
 sg13g2_fill_2 FILLER_3_331 ();
 sg13g2_fill_1 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_360 ();
 sg13g2_decap_8 FILLER_3_367 ();
 sg13g2_decap_8 FILLER_3_374 ();
 sg13g2_decap_8 FILLER_3_381 ();
 sg13g2_decap_8 FILLER_3_388 ();
 sg13g2_decap_8 FILLER_3_395 ();
 sg13g2_decap_8 FILLER_3_402 ();
 sg13g2_decap_8 FILLER_3_409 ();
 sg13g2_decap_8 FILLER_3_416 ();
 sg13g2_decap_8 FILLER_3_423 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_fill_1 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_75 ();
 sg13g2_decap_8 FILLER_4_82 ();
 sg13g2_fill_2 FILLER_4_89 ();
 sg13g2_fill_1 FILLER_4_91 ();
 sg13g2_fill_2 FILLER_4_144 ();
 sg13g2_fill_1 FILLER_4_146 ();
 sg13g2_decap_8 FILLER_4_159 ();
 sg13g2_decap_8 FILLER_4_166 ();
 sg13g2_decap_4 FILLER_4_173 ();
 sg13g2_fill_2 FILLER_4_177 ();
 sg13g2_decap_8 FILLER_4_209 ();
 sg13g2_fill_1 FILLER_4_216 ();
 sg13g2_fill_2 FILLER_4_248 ();
 sg13g2_fill_1 FILLER_4_250 ();
 sg13g2_decap_8 FILLER_4_268 ();
 sg13g2_decap_8 FILLER_4_275 ();
 sg13g2_fill_1 FILLER_4_345 ();
 sg13g2_fill_2 FILLER_4_350 ();
 sg13g2_fill_1 FILLER_4_352 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_8 FILLER_4_416 ();
 sg13g2_decap_8 FILLER_4_423 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_4 FILLER_5_14 ();
 sg13g2_fill_1 FILLER_5_18 ();
 sg13g2_fill_2 FILLER_5_52 ();
 sg13g2_fill_1 FILLER_5_54 ();
 sg13g2_fill_1 FILLER_5_81 ();
 sg13g2_fill_1 FILLER_5_96 ();
 sg13g2_decap_4 FILLER_5_105 ();
 sg13g2_fill_1 FILLER_5_109 ();
 sg13g2_fill_1 FILLER_5_113 ();
 sg13g2_fill_2 FILLER_5_141 ();
 sg13g2_fill_2 FILLER_5_160 ();
 sg13g2_fill_2 FILLER_5_193 ();
 sg13g2_fill_1 FILLER_5_200 ();
 sg13g2_fill_2 FILLER_5_240 ();
 sg13g2_fill_1 FILLER_5_247 ();
 sg13g2_fill_1 FILLER_5_252 ();
 sg13g2_fill_1 FILLER_5_279 ();
 sg13g2_fill_2 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_8 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_5_412 ();
 sg13g2_decap_8 FILLER_5_419 ();
 sg13g2_decap_4 FILLER_5_426 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_fill_1 FILLER_6_28 ();
 sg13g2_decap_4 FILLER_6_41 ();
 sg13g2_fill_2 FILLER_6_87 ();
 sg13g2_fill_1 FILLER_6_89 ();
 sg13g2_fill_2 FILLER_6_94 ();
 sg13g2_fill_1 FILLER_6_139 ();
 sg13g2_fill_1 FILLER_6_185 ();
 sg13g2_fill_1 FILLER_6_193 ();
 sg13g2_fill_1 FILLER_6_198 ();
 sg13g2_fill_2 FILLER_6_203 ();
 sg13g2_fill_2 FILLER_6_209 ();
 sg13g2_fill_2 FILLER_6_215 ();
 sg13g2_fill_2 FILLER_6_221 ();
 sg13g2_fill_1 FILLER_6_223 ();
 sg13g2_fill_2 FILLER_6_228 ();
 sg13g2_fill_1 FILLER_6_230 ();
 sg13g2_fill_2 FILLER_6_236 ();
 sg13g2_fill_2 FILLER_6_268 ();
 sg13g2_fill_1 FILLER_6_270 ();
 sg13g2_fill_1 FILLER_6_314 ();
 sg13g2_fill_1 FILLER_6_319 ();
 sg13g2_fill_1 FILLER_6_324 ();
 sg13g2_fill_1 FILLER_6_330 ();
 sg13g2_fill_1 FILLER_6_335 ();
 sg13g2_fill_2 FILLER_6_345 ();
 sg13g2_fill_1 FILLER_6_347 ();
 sg13g2_fill_1 FILLER_6_353 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_decap_8 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_6_415 ();
 sg13g2_decap_8 FILLER_6_422 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_fill_2 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_27 ();
 sg13g2_decap_4 FILLER_7_34 ();
 sg13g2_fill_1 FILLER_7_38 ();
 sg13g2_decap_8 FILLER_7_64 ();
 sg13g2_fill_2 FILLER_7_83 ();
 sg13g2_fill_1 FILLER_7_85 ();
 sg13g2_fill_2 FILLER_7_96 ();
 sg13g2_decap_4 FILLER_7_113 ();
 sg13g2_fill_2 FILLER_7_122 ();
 sg13g2_fill_2 FILLER_7_128 ();
 sg13g2_fill_1 FILLER_7_157 ();
 sg13g2_decap_4 FILLER_7_163 ();
 sg13g2_fill_1 FILLER_7_178 ();
 sg13g2_fill_2 FILLER_7_184 ();
 sg13g2_fill_1 FILLER_7_241 ();
 sg13g2_fill_2 FILLER_7_260 ();
 sg13g2_fill_2 FILLER_7_266 ();
 sg13g2_fill_1 FILLER_7_272 ();
 sg13g2_fill_2 FILLER_7_277 ();
 sg13g2_fill_2 FILLER_7_288 ();
 sg13g2_fill_1 FILLER_7_290 ();
 sg13g2_fill_2 FILLER_7_304 ();
 sg13g2_fill_1 FILLER_7_340 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_7_409 ();
 sg13g2_decap_8 FILLER_7_416 ();
 sg13g2_decap_8 FILLER_7_423 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_fill_2 FILLER_8_14 ();
 sg13g2_fill_2 FILLER_8_42 ();
 sg13g2_fill_2 FILLER_8_69 ();
 sg13g2_fill_1 FILLER_8_71 ();
 sg13g2_decap_4 FILLER_8_102 ();
 sg13g2_fill_1 FILLER_8_134 ();
 sg13g2_fill_2 FILLER_8_157 ();
 sg13g2_fill_1 FILLER_8_170 ();
 sg13g2_fill_2 FILLER_8_196 ();
 sg13g2_fill_1 FILLER_8_207 ();
 sg13g2_fill_1 FILLER_8_218 ();
 sg13g2_fill_1 FILLER_8_224 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_fill_1 FILLER_8_339 ();
 sg13g2_fill_2 FILLER_8_345 ();
 sg13g2_fill_2 FILLER_8_352 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_decap_8 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_8_415 ();
 sg13g2_decap_8 FILLER_8_422 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_18 ();
 sg13g2_fill_1 FILLER_9_23 ();
 sg13g2_fill_1 FILLER_9_52 ();
 sg13g2_fill_1 FILLER_9_57 ();
 sg13g2_fill_1 FILLER_9_88 ();
 sg13g2_decap_4 FILLER_9_101 ();
 sg13g2_decap_4 FILLER_9_142 ();
 sg13g2_fill_1 FILLER_9_146 ();
 sg13g2_fill_2 FILLER_9_157 ();
 sg13g2_fill_1 FILLER_9_159 ();
 sg13g2_fill_1 FILLER_9_216 ();
 sg13g2_fill_1 FILLER_9_221 ();
 sg13g2_fill_1 FILLER_9_226 ();
 sg13g2_fill_2 FILLER_9_231 ();
 sg13g2_fill_2 FILLER_9_242 ();
 sg13g2_fill_2 FILLER_9_248 ();
 sg13g2_fill_2 FILLER_9_255 ();
 sg13g2_fill_1 FILLER_9_265 ();
 sg13g2_decap_4 FILLER_9_270 ();
 sg13g2_fill_1 FILLER_9_274 ();
 sg13g2_fill_1 FILLER_9_280 ();
 sg13g2_fill_1 FILLER_9_298 ();
 sg13g2_fill_1 FILLER_9_315 ();
 sg13g2_fill_1 FILLER_9_319 ();
 sg13g2_fill_1 FILLER_9_367 ();
 sg13g2_fill_1 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_58 ();
 sg13g2_fill_2 FILLER_10_64 ();
 sg13g2_fill_1 FILLER_10_66 ();
 sg13g2_fill_2 FILLER_10_71 ();
 sg13g2_fill_2 FILLER_10_165 ();
 sg13g2_fill_2 FILLER_10_197 ();
 sg13g2_fill_1 FILLER_10_331 ();
 sg13g2_fill_1 FILLER_10_347 ();
 sg13g2_fill_2 FILLER_10_362 ();
 sg13g2_fill_1 FILLER_10_378 ();
 sg13g2_fill_1 FILLER_10_410 ();
 sg13g2_decap_8 FILLER_10_415 ();
 sg13g2_decap_8 FILLER_10_422 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_fill_1 FILLER_11_32 ();
 sg13g2_fill_1 FILLER_11_59 ();
 sg13g2_fill_1 FILLER_11_141 ();
 sg13g2_fill_2 FILLER_11_210 ();
 sg13g2_decap_4 FILLER_11_225 ();
 sg13g2_fill_1 FILLER_11_229 ();
 sg13g2_fill_1 FILLER_11_234 ();
 sg13g2_decap_8 FILLER_11_240 ();
 sg13g2_decap_4 FILLER_11_247 ();
 sg13g2_fill_2 FILLER_11_251 ();
 sg13g2_fill_1 FILLER_11_261 ();
 sg13g2_fill_1 FILLER_11_267 ();
 sg13g2_fill_1 FILLER_11_273 ();
 sg13g2_fill_1 FILLER_11_282 ();
 sg13g2_fill_2 FILLER_11_326 ();
 sg13g2_fill_1 FILLER_11_332 ();
 sg13g2_fill_1 FILLER_11_348 ();
 sg13g2_fill_1 FILLER_11_375 ();
 sg13g2_fill_2 FILLER_11_386 ();
 sg13g2_fill_2 FILLER_11_416 ();
 sg13g2_fill_1 FILLER_11_418 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_34 ();
 sg13g2_decap_8 FILLER_12_60 ();
 sg13g2_fill_1 FILLER_12_67 ();
 sg13g2_fill_1 FILLER_12_82 ();
 sg13g2_fill_1 FILLER_12_96 ();
 sg13g2_fill_2 FILLER_12_102 ();
 sg13g2_fill_2 FILLER_12_189 ();
 sg13g2_fill_1 FILLER_12_203 ();
 sg13g2_decap_4 FILLER_12_240 ();
 sg13g2_fill_1 FILLER_12_251 ();
 sg13g2_decap_4 FILLER_12_282 ();
 sg13g2_fill_1 FILLER_12_286 ();
 sg13g2_fill_1 FILLER_12_357 ();
 sg13g2_fill_2 FILLER_12_363 ();
 sg13g2_fill_1 FILLER_12_391 ();
 sg13g2_fill_2 FILLER_12_402 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_8 ();
 sg13g2_fill_1 FILLER_13_40 ();
 sg13g2_fill_1 FILLER_13_45 ();
 sg13g2_decap_4 FILLER_13_59 ();
 sg13g2_fill_2 FILLER_13_89 ();
 sg13g2_fill_2 FILLER_13_112 ();
 sg13g2_fill_1 FILLER_13_134 ();
 sg13g2_fill_1 FILLER_13_143 ();
 sg13g2_fill_1 FILLER_13_150 ();
 sg13g2_fill_1 FILLER_13_158 ();
 sg13g2_fill_2 FILLER_13_165 ();
 sg13g2_fill_2 FILLER_13_172 ();
 sg13g2_decap_4 FILLER_13_182 ();
 sg13g2_fill_2 FILLER_13_214 ();
 sg13g2_fill_1 FILLER_13_224 ();
 sg13g2_fill_1 FILLER_13_237 ();
 sg13g2_decap_4 FILLER_13_242 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_260 ();
 sg13g2_fill_1 FILLER_13_269 ();
 sg13g2_fill_1 FILLER_13_296 ();
 sg13g2_fill_1 FILLER_13_301 ();
 sg13g2_decap_4 FILLER_13_308 ();
 sg13g2_fill_1 FILLER_13_312 ();
 sg13g2_decap_4 FILLER_13_317 ();
 sg13g2_fill_2 FILLER_13_321 ();
 sg13g2_fill_2 FILLER_13_332 ();
 sg13g2_fill_1 FILLER_13_334 ();
 sg13g2_fill_1 FILLER_13_402 ();
 sg13g2_fill_1 FILLER_13_416 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_fill_1 FILLER_14_34 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_fill_1 FILLER_14_45 ();
 sg13g2_fill_2 FILLER_14_54 ();
 sg13g2_fill_1 FILLER_14_64 ();
 sg13g2_fill_2 FILLER_14_69 ();
 sg13g2_fill_2 FILLER_14_119 ();
 sg13g2_fill_2 FILLER_14_130 ();
 sg13g2_decap_4 FILLER_14_138 ();
 sg13g2_fill_2 FILLER_14_142 ();
 sg13g2_fill_1 FILLER_14_162 ();
 sg13g2_fill_2 FILLER_14_216 ();
 sg13g2_fill_1 FILLER_14_252 ();
 sg13g2_fill_1 FILLER_14_261 ();
 sg13g2_fill_1 FILLER_14_269 ();
 sg13g2_fill_2 FILLER_14_278 ();
 sg13g2_fill_2 FILLER_14_284 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_fill_1 FILLER_14_343 ();
 sg13g2_decap_4 FILLER_14_371 ();
 sg13g2_fill_2 FILLER_14_375 ();
 sg13g2_fill_2 FILLER_14_382 ();
 sg13g2_fill_1 FILLER_14_423 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_62 ();
 sg13g2_fill_2 FILLER_15_94 ();
 sg13g2_fill_1 FILLER_15_96 ();
 sg13g2_fill_2 FILLER_15_105 ();
 sg13g2_fill_2 FILLER_15_112 ();
 sg13g2_fill_1 FILLER_15_114 ();
 sg13g2_decap_4 FILLER_15_123 ();
 sg13g2_fill_1 FILLER_15_127 ();
 sg13g2_fill_1 FILLER_15_141 ();
 sg13g2_fill_1 FILLER_15_150 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_195 ();
 sg13g2_fill_1 FILLER_15_205 ();
 sg13g2_fill_2 FILLER_15_222 ();
 sg13g2_decap_8 FILLER_15_236 ();
 sg13g2_decap_4 FILLER_15_243 ();
 sg13g2_fill_2 FILLER_15_247 ();
 sg13g2_fill_2 FILLER_15_259 ();
 sg13g2_fill_1 FILLER_15_261 ();
 sg13g2_fill_2 FILLER_15_267 ();
 sg13g2_fill_2 FILLER_15_320 ();
 sg13g2_fill_1 FILLER_15_332 ();
 sg13g2_fill_2 FILLER_15_343 ();
 sg13g2_fill_1 FILLER_15_345 ();
 sg13g2_fill_2 FILLER_15_354 ();
 sg13g2_fill_2 FILLER_15_382 ();
 sg13g2_fill_1 FILLER_15_384 ();
 sg13g2_fill_1 FILLER_15_419 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_fill_1 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_27 ();
 sg13g2_fill_2 FILLER_16_32 ();
 sg13g2_decap_4 FILLER_16_50 ();
 sg13g2_fill_1 FILLER_16_54 ();
 sg13g2_fill_1 FILLER_16_73 ();
 sg13g2_fill_2 FILLER_16_78 ();
 sg13g2_decap_8 FILLER_16_89 ();
 sg13g2_fill_2 FILLER_16_96 ();
 sg13g2_fill_1 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_124 ();
 sg13g2_fill_1 FILLER_16_126 ();
 sg13g2_fill_1 FILLER_16_131 ();
 sg13g2_decap_4 FILLER_16_140 ();
 sg13g2_fill_2 FILLER_16_144 ();
 sg13g2_fill_1 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_175 ();
 sg13g2_fill_2 FILLER_16_235 ();
 sg13g2_fill_1 FILLER_16_254 ();
 sg13g2_fill_2 FILLER_16_266 ();
 sg13g2_decap_4 FILLER_16_276 ();
 sg13g2_decap_8 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_298 ();
 sg13g2_fill_2 FILLER_16_303 ();
 sg13g2_fill_2 FILLER_16_314 ();
 sg13g2_fill_1 FILLER_16_353 ();
 sg13g2_fill_2 FILLER_16_358 ();
 sg13g2_fill_2 FILLER_16_386 ();
 sg13g2_fill_1 FILLER_16_388 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_4 ();
 sg13g2_decap_8 FILLER_17_13 ();
 sg13g2_fill_2 FILLER_17_20 ();
 sg13g2_decap_8 FILLER_17_26 ();
 sg13g2_fill_1 FILLER_17_33 ();
 sg13g2_decap_4 FILLER_17_51 ();
 sg13g2_fill_2 FILLER_17_68 ();
 sg13g2_fill_1 FILLER_17_74 ();
 sg13g2_fill_1 FILLER_17_82 ();
 sg13g2_fill_1 FILLER_17_91 ();
 sg13g2_fill_1 FILLER_17_100 ();
 sg13g2_fill_1 FILLER_17_106 ();
 sg13g2_fill_1 FILLER_17_111 ();
 sg13g2_fill_2 FILLER_17_120 ();
 sg13g2_decap_4 FILLER_17_151 ();
 sg13g2_fill_1 FILLER_17_155 ();
 sg13g2_decap_4 FILLER_17_184 ();
 sg13g2_fill_2 FILLER_17_188 ();
 sg13g2_fill_2 FILLER_17_213 ();
 sg13g2_fill_1 FILLER_17_215 ();
 sg13g2_fill_2 FILLER_17_227 ();
 sg13g2_fill_1 FILLER_17_229 ();
 sg13g2_fill_2 FILLER_17_234 ();
 sg13g2_decap_4 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_257 ();
 sg13g2_decap_4 FILLER_17_294 ();
 sg13g2_fill_2 FILLER_17_328 ();
 sg13g2_fill_1 FILLER_17_330 ();
 sg13g2_decap_4 FILLER_17_357 ();
 sg13g2_fill_1 FILLER_17_361 ();
 sg13g2_fill_1 FILLER_17_420 ();
 sg13g2_decap_4 FILLER_17_425 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_34 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_fill_1 FILLER_18_96 ();
 sg13g2_fill_2 FILLER_18_101 ();
 sg13g2_decap_4 FILLER_18_109 ();
 sg13g2_fill_1 FILLER_18_113 ();
 sg13g2_fill_1 FILLER_18_138 ();
 sg13g2_decap_8 FILLER_18_167 ();
 sg13g2_fill_2 FILLER_18_174 ();
 sg13g2_fill_1 FILLER_18_176 ();
 sg13g2_fill_2 FILLER_18_184 ();
 sg13g2_fill_1 FILLER_18_261 ();
 sg13g2_fill_2 FILLER_18_266 ();
 sg13g2_fill_1 FILLER_18_268 ();
 sg13g2_fill_1 FILLER_18_273 ();
 sg13g2_fill_2 FILLER_18_333 ();
 sg13g2_fill_1 FILLER_18_354 ();
 sg13g2_fill_2 FILLER_18_386 ();
 sg13g2_fill_1 FILLER_18_388 ();
 sg13g2_fill_1 FILLER_18_394 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_27 ();
 sg13g2_fill_1 FILLER_19_40 ();
 sg13g2_decap_8 FILLER_19_44 ();
 sg13g2_fill_2 FILLER_19_56 ();
 sg13g2_fill_1 FILLER_19_66 ();
 sg13g2_fill_2 FILLER_19_109 ();
 sg13g2_fill_1 FILLER_19_121 ();
 sg13g2_fill_2 FILLER_19_127 ();
 sg13g2_fill_2 FILLER_19_134 ();
 sg13g2_fill_2 FILLER_19_143 ();
 sg13g2_fill_1 FILLER_19_145 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_fill_2 FILLER_19_186 ();
 sg13g2_fill_2 FILLER_19_220 ();
 sg13g2_fill_2 FILLER_19_226 ();
 sg13g2_fill_1 FILLER_19_228 ();
 sg13g2_fill_2 FILLER_19_233 ();
 sg13g2_fill_1 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_240 ();
 sg13g2_fill_2 FILLER_19_267 ();
 sg13g2_fill_2 FILLER_19_273 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_fill_2 FILLER_19_332 ();
 sg13g2_fill_1 FILLER_19_334 ();
 sg13g2_fill_1 FILLER_19_340 ();
 sg13g2_fill_1 FILLER_19_395 ();
 sg13g2_fill_1 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_414 ();
 sg13g2_decap_8 FILLER_19_419 ();
 sg13g2_decap_4 FILLER_19_426 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_49 ();
 sg13g2_fill_1 FILLER_20_53 ();
 sg13g2_fill_2 FILLER_20_70 ();
 sg13g2_fill_1 FILLER_20_104 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_fill_1 FILLER_20_125 ();
 sg13g2_fill_2 FILLER_20_154 ();
 sg13g2_fill_1 FILLER_20_170 ();
 sg13g2_decap_4 FILLER_20_187 ();
 sg13g2_fill_1 FILLER_20_191 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_fill_1 FILLER_20_216 ();
 sg13g2_fill_1 FILLER_20_222 ();
 sg13g2_fill_1 FILLER_20_228 ();
 sg13g2_fill_1 FILLER_20_234 ();
 sg13g2_fill_1 FILLER_20_239 ();
 sg13g2_fill_2 FILLER_20_245 ();
 sg13g2_decap_4 FILLER_20_251 ();
 sg13g2_fill_1 FILLER_20_255 ();
 sg13g2_decap_4 FILLER_20_260 ();
 sg13g2_fill_1 FILLER_20_264 ();
 sg13g2_fill_1 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_316 ();
 sg13g2_fill_1 FILLER_20_321 ();
 sg13g2_fill_2 FILLER_20_327 ();
 sg13g2_fill_2 FILLER_20_333 ();
 sg13g2_fill_1 FILLER_20_335 ();
 sg13g2_fill_2 FILLER_20_341 ();
 sg13g2_fill_2 FILLER_20_351 ();
 sg13g2_fill_1 FILLER_20_358 ();
 sg13g2_fill_1 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_107 ();
 sg13g2_fill_2 FILLER_21_116 ();
 sg13g2_fill_2 FILLER_21_123 ();
 sg13g2_fill_1 FILLER_21_125 ();
 sg13g2_fill_2 FILLER_21_130 ();
 sg13g2_fill_1 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_138 ();
 sg13g2_fill_1 FILLER_21_143 ();
 sg13g2_decap_4 FILLER_21_159 ();
 sg13g2_fill_1 FILLER_21_167 ();
 sg13g2_decap_8 FILLER_21_173 ();
 sg13g2_decap_4 FILLER_21_180 ();
 sg13g2_fill_1 FILLER_21_210 ();
 sg13g2_fill_1 FILLER_21_216 ();
 sg13g2_fill_2 FILLER_21_235 ();
 sg13g2_decap_8 FILLER_21_254 ();
 sg13g2_decap_4 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_265 ();
 sg13g2_fill_2 FILLER_21_324 ();
 sg13g2_fill_2 FILLER_21_347 ();
 sg13g2_fill_1 FILLER_21_380 ();
 sg13g2_fill_1 FILLER_21_385 ();
 sg13g2_fill_1 FILLER_21_414 ();
 sg13g2_fill_2 FILLER_21_419 ();
 sg13g2_decap_4 FILLER_21_425 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_fill_2 FILLER_22_34 ();
 sg13g2_fill_1 FILLER_22_36 ();
 sg13g2_decap_4 FILLER_22_61 ();
 sg13g2_fill_2 FILLER_22_65 ();
 sg13g2_decap_4 FILLER_22_87 ();
 sg13g2_decap_4 FILLER_22_108 ();
 sg13g2_fill_2 FILLER_22_112 ();
 sg13g2_fill_2 FILLER_22_149 ();
 sg13g2_fill_2 FILLER_22_171 ();
 sg13g2_fill_1 FILLER_22_173 ();
 sg13g2_decap_8 FILLER_22_195 ();
 sg13g2_fill_2 FILLER_22_202 ();
 sg13g2_fill_1 FILLER_22_214 ();
 sg13g2_fill_1 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_225 ();
 sg13g2_fill_1 FILLER_22_257 ();
 sg13g2_fill_1 FILLER_22_262 ();
 sg13g2_fill_2 FILLER_22_275 ();
 sg13g2_fill_1 FILLER_22_281 ();
 sg13g2_fill_1 FILLER_22_341 ();
 sg13g2_fill_1 FILLER_22_345 ();
 sg13g2_fill_2 FILLER_22_384 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_fill_2 FILLER_23_36 ();
 sg13g2_fill_1 FILLER_23_38 ();
 sg13g2_fill_2 FILLER_23_53 ();
 sg13g2_fill_1 FILLER_23_64 ();
 sg13g2_fill_2 FILLER_23_81 ();
 sg13g2_decap_4 FILLER_23_88 ();
 sg13g2_fill_2 FILLER_23_103 ();
 sg13g2_fill_1 FILLER_23_121 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_fill_1 FILLER_23_135 ();
 sg13g2_fill_2 FILLER_23_144 ();
 sg13g2_decap_8 FILLER_23_151 ();
 sg13g2_fill_2 FILLER_23_158 ();
 sg13g2_fill_1 FILLER_23_194 ();
 sg13g2_fill_1 FILLER_23_208 ();
 sg13g2_fill_1 FILLER_23_247 ();
 sg13g2_fill_1 FILLER_23_321 ();
 sg13g2_fill_1 FILLER_23_326 ();
 sg13g2_fill_2 FILLER_23_337 ();
 sg13g2_fill_1 FILLER_23_339 ();
 sg13g2_fill_2 FILLER_23_366 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_34 ();
 sg13g2_fill_1 FILLER_24_41 ();
 sg13g2_decap_4 FILLER_24_58 ();
 sg13g2_fill_2 FILLER_24_62 ();
 sg13g2_fill_1 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_100 ();
 sg13g2_fill_2 FILLER_24_105 ();
 sg13g2_fill_1 FILLER_24_124 ();
 sg13g2_fill_2 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_fill_2 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_fill_1 FILLER_24_199 ();
 sg13g2_fill_1 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_fill_2 FILLER_24_226 ();
 sg13g2_fill_1 FILLER_24_258 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_fill_2 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_61 ();
 sg13g2_fill_1 FILLER_25_70 ();
 sg13g2_fill_1 FILLER_25_100 ();
 sg13g2_fill_2 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_fill_2 FILLER_25_112 ();
 sg13g2_fill_1 FILLER_25_124 ();
 sg13g2_decap_4 FILLER_25_155 ();
 sg13g2_fill_2 FILLER_25_189 ();
 sg13g2_fill_1 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_fill_1 FILLER_25_209 ();
 sg13g2_decap_8 FILLER_25_226 ();
 sg13g2_fill_2 FILLER_25_237 ();
 sg13g2_fill_2 FILLER_25_243 ();
 sg13g2_fill_1 FILLER_25_245 ();
 sg13g2_fill_1 FILLER_25_285 ();
 sg13g2_fill_2 FILLER_25_329 ();
 sg13g2_fill_1 FILLER_25_331 ();
 sg13g2_fill_2 FILLER_25_374 ();
 sg13g2_fill_2 FILLER_25_396 ();
 sg13g2_decap_8 FILLER_26_38 ();
 sg13g2_decap_4 FILLER_26_45 ();
 sg13g2_fill_2 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_62 ();
 sg13g2_fill_2 FILLER_26_75 ();
 sg13g2_fill_1 FILLER_26_111 ();
 sg13g2_decap_8 FILLER_26_117 ();
 sg13g2_fill_1 FILLER_26_124 ();
 sg13g2_fill_1 FILLER_26_129 ();
 sg13g2_fill_1 FILLER_26_137 ();
 sg13g2_fill_1 FILLER_26_153 ();
 sg13g2_fill_2 FILLER_26_203 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_226 ();
 sg13g2_fill_2 FILLER_26_265 ();
 sg13g2_fill_2 FILLER_26_281 ();
 sg13g2_fill_1 FILLER_26_283 ();
 sg13g2_fill_1 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_312 ();
 sg13g2_fill_2 FILLER_26_346 ();
 sg13g2_fill_2 FILLER_26_352 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_fill_2 FILLER_26_364 ();
 sg13g2_fill_2 FILLER_26_397 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_fill_1 FILLER_27_60 ();
 sg13g2_fill_2 FILLER_27_74 ();
 sg13g2_decap_4 FILLER_27_100 ();
 sg13g2_fill_1 FILLER_27_108 ();
 sg13g2_decap_8 FILLER_27_113 ();
 sg13g2_fill_1 FILLER_27_125 ();
 sg13g2_fill_2 FILLER_27_146 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_fill_2 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_207 ();
 sg13g2_fill_1 FILLER_27_212 ();
 sg13g2_fill_1 FILLER_27_220 ();
 sg13g2_fill_2 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_fill_2 FILLER_27_316 ();
 sg13g2_fill_1 FILLER_27_323 ();
 sg13g2_fill_1 FILLER_27_331 ();
 sg13g2_fill_1 FILLER_27_358 ();
 sg13g2_fill_1 FILLER_27_390 ();
 sg13g2_fill_1 FILLER_27_423 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_30 ();
 sg13g2_decap_4 FILLER_28_37 ();
 sg13g2_fill_1 FILLER_28_41 ();
 sg13g2_decap_4 FILLER_28_50 ();
 sg13g2_fill_1 FILLER_28_91 ();
 sg13g2_fill_2 FILLER_28_100 ();
 sg13g2_fill_1 FILLER_28_102 ();
 sg13g2_fill_1 FILLER_28_124 ();
 sg13g2_fill_1 FILLER_28_138 ();
 sg13g2_fill_2 FILLER_28_144 ();
 sg13g2_fill_1 FILLER_28_146 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_188 ();
 sg13g2_fill_2 FILLER_28_202 ();
 sg13g2_fill_1 FILLER_28_223 ();
 sg13g2_fill_1 FILLER_28_250 ();
 sg13g2_fill_2 FILLER_28_264 ();
 sg13g2_fill_1 FILLER_28_271 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_fill_2 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_311 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_fill_2 FILLER_28_319 ();
 sg13g2_fill_2 FILLER_28_340 ();
 sg13g2_decap_4 FILLER_28_350 ();
 sg13g2_fill_1 FILLER_28_359 ();
 sg13g2_fill_1 FILLER_28_365 ();
 sg13g2_fill_1 FILLER_28_370 ();
 sg13g2_fill_2 FILLER_28_393 ();
 sg13g2_fill_2 FILLER_29_64 ();
 sg13g2_fill_2 FILLER_29_70 ();
 sg13g2_fill_1 FILLER_29_86 ();
 sg13g2_fill_2 FILLER_29_103 ();
 sg13g2_fill_1 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_124 ();
 sg13g2_fill_2 FILLER_29_133 ();
 sg13g2_fill_2 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_160 ();
 sg13g2_fill_1 FILLER_29_204 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_fill_2 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_7 ();
 sg13g2_fill_2 FILLER_30_29 ();
 sg13g2_fill_1 FILLER_30_31 ();
 sg13g2_decap_4 FILLER_30_36 ();
 sg13g2_fill_1 FILLER_30_40 ();
 sg13g2_fill_2 FILLER_30_48 ();
 sg13g2_fill_1 FILLER_30_50 ();
 sg13g2_fill_2 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_65 ();
 sg13g2_decap_8 FILLER_30_104 ();
 sg13g2_fill_2 FILLER_30_111 ();
 sg13g2_decap_4 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_fill_1 FILLER_30_160 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_fill_1 FILLER_30_170 ();
 sg13g2_fill_2 FILLER_30_175 ();
 sg13g2_fill_2 FILLER_30_182 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_fill_2 FILLER_30_193 ();
 sg13g2_fill_1 FILLER_30_195 ();
 sg13g2_fill_2 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_202 ();
 sg13g2_decap_4 FILLER_30_233 ();
 sg13g2_fill_1 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_261 ();
 sg13g2_fill_1 FILLER_30_289 ();
 sg13g2_fill_1 FILLER_30_370 ();
 sg13g2_fill_2 FILLER_30_375 ();
 sg13g2_fill_1 FILLER_30_386 ();
 sg13g2_fill_1 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_12 ();
 sg13g2_fill_1 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_27 ();
 sg13g2_fill_1 FILLER_31_34 ();
 sg13g2_fill_1 FILLER_31_48 ();
 sg13g2_fill_1 FILLER_31_57 ();
 sg13g2_fill_1 FILLER_31_66 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_fill_2 FILLER_31_85 ();
 sg13g2_fill_2 FILLER_31_104 ();
 sg13g2_fill_1 FILLER_31_131 ();
 sg13g2_fill_1 FILLER_31_153 ();
 sg13g2_fill_2 FILLER_31_184 ();
 sg13g2_fill_2 FILLER_31_264 ();
 sg13g2_fill_1 FILLER_31_266 ();
 sg13g2_fill_1 FILLER_31_298 ();
 sg13g2_fill_1 FILLER_31_304 ();
 sg13g2_fill_1 FILLER_31_318 ();
 sg13g2_fill_1 FILLER_31_329 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_fill_2 FILLER_32_103 ();
 sg13g2_fill_1 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_114 ();
 sg13g2_fill_2 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_125 ();
 sg13g2_decap_4 FILLER_32_129 ();
 sg13g2_fill_1 FILLER_32_171 ();
 sg13g2_fill_1 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_227 ();
 sg13g2_fill_2 FILLER_32_234 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_decap_8 FILLER_32_254 ();
 sg13g2_decap_4 FILLER_32_261 ();
 sg13g2_fill_1 FILLER_32_265 ();
 sg13g2_fill_1 FILLER_32_270 ();
 sg13g2_fill_1 FILLER_32_275 ();
 sg13g2_fill_1 FILLER_32_280 ();
 sg13g2_fill_1 FILLER_32_285 ();
 sg13g2_fill_2 FILLER_32_291 ();
 sg13g2_fill_2 FILLER_32_348 ();
 sg13g2_fill_1 FILLER_32_350 ();
 sg13g2_fill_2 FILLER_32_390 ();
 sg13g2_fill_2 FILLER_32_397 ();
 sg13g2_fill_2 FILLER_33_30 ();
 sg13g2_decap_4 FILLER_33_36 ();
 sg13g2_fill_2 FILLER_33_44 ();
 sg13g2_fill_2 FILLER_33_83 ();
 sg13g2_fill_1 FILLER_33_111 ();
 sg13g2_fill_1 FILLER_33_125 ();
 sg13g2_fill_2 FILLER_33_138 ();
 sg13g2_fill_1 FILLER_33_140 ();
 sg13g2_fill_2 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_153 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_decap_8 FILLER_33_228 ();
 sg13g2_fill_2 FILLER_33_265 ();
 sg13g2_fill_1 FILLER_33_267 ();
 sg13g2_fill_1 FILLER_33_272 ();
 sg13g2_fill_2 FILLER_33_324 ();
 sg13g2_fill_2 FILLER_33_348 ();
 sg13g2_fill_2 FILLER_33_354 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_fill_2 FILLER_34_78 ();
 sg13g2_fill_1 FILLER_34_88 ();
 sg13g2_fill_1 FILLER_34_117 ();
 sg13g2_fill_2 FILLER_34_146 ();
 sg13g2_fill_1 FILLER_34_153 ();
 sg13g2_decap_4 FILLER_34_180 ();
 sg13g2_fill_2 FILLER_34_243 ();
 sg13g2_fill_2 FILLER_34_319 ();
 sg13g2_fill_2 FILLER_34_427 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_29 ();
 sg13g2_fill_1 FILLER_35_31 ();
 sg13g2_fill_2 FILLER_35_49 ();
 sg13g2_fill_2 FILLER_35_60 ();
 sg13g2_fill_2 FILLER_35_67 ();
 sg13g2_fill_1 FILLER_35_73 ();
 sg13g2_fill_1 FILLER_35_114 ();
 sg13g2_fill_1 FILLER_35_135 ();
 sg13g2_fill_1 FILLER_35_145 ();
 sg13g2_fill_1 FILLER_35_151 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_fill_1 FILLER_35_162 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_decap_8 FILLER_35_177 ();
 sg13g2_decap_4 FILLER_35_234 ();
 sg13g2_fill_1 FILLER_35_242 ();
 sg13g2_fill_1 FILLER_35_274 ();
 sg13g2_fill_2 FILLER_35_280 ();
 sg13g2_fill_2 FILLER_35_294 ();
 sg13g2_fill_1 FILLER_35_306 ();
 sg13g2_fill_1 FILLER_35_316 ();
 sg13g2_fill_2 FILLER_35_347 ();
 sg13g2_fill_1 FILLER_35_359 ();
 sg13g2_fill_1 FILLER_36_47 ();
 sg13g2_fill_1 FILLER_36_55 ();
 sg13g2_fill_1 FILLER_36_78 ();
 sg13g2_fill_1 FILLER_36_83 ();
 sg13g2_fill_1 FILLER_36_88 ();
 sg13g2_fill_1 FILLER_36_93 ();
 sg13g2_fill_1 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_104 ();
 sg13g2_fill_1 FILLER_36_117 ();
 sg13g2_fill_1 FILLER_36_141 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_fill_2 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_37_26 ();
 sg13g2_fill_1 FILLER_37_28 ();
 sg13g2_fill_1 FILLER_37_33 ();
 sg13g2_fill_2 FILLER_37_38 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_fill_2 FILLER_37_137 ();
 sg13g2_fill_2 FILLER_37_163 ();
 sg13g2_fill_1 FILLER_37_185 ();
 sg13g2_fill_1 FILLER_37_218 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_fill_2 FILLER_37_259 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_fill_2 FILLER_37_307 ();
 sg13g2_fill_1 FILLER_37_321 ();
 sg13g2_fill_1 FILLER_37_353 ();
 sg13g2_fill_2 FILLER_37_384 ();
 sg13g2_fill_1 FILLER_37_396 ();
 sg13g2_fill_2 FILLER_37_428 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_2 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_75 ();
 sg13g2_fill_2 FILLER_38_177 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_fill_1 FILLER_38_188 ();
 sg13g2_fill_1 FILLER_38_193 ();
 sg13g2_fill_1 FILLER_38_273 ();
 sg13g2_fill_1 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_305 ();
 sg13g2_fill_1 FILLER_38_310 ();
 sg13g2_fill_1 FILLER_38_348 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_fill_1 FILLER_38_429 ();
endmodule
