module tt_um_rtfb_collatz (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire clknet_0_clk;
 wire net344;
 wire \collatz.busy ;
 wire \collatz.comp ;
 wire \collatz.iter[0] ;
 wire \collatz.iter[100] ;
 wire \collatz.iter[101] ;
 wire \collatz.iter[102] ;
 wire \collatz.iter[103] ;
 wire \collatz.iter[104] ;
 wire \collatz.iter[105] ;
 wire \collatz.iter[106] ;
 wire \collatz.iter[107] ;
 wire \collatz.iter[108] ;
 wire \collatz.iter[109] ;
 wire \collatz.iter[10] ;
 wire \collatz.iter[110] ;
 wire \collatz.iter[111] ;
 wire \collatz.iter[112] ;
 wire \collatz.iter[113] ;
 wire \collatz.iter[114] ;
 wire \collatz.iter[115] ;
 wire \collatz.iter[116] ;
 wire \collatz.iter[117] ;
 wire \collatz.iter[118] ;
 wire \collatz.iter[119] ;
 wire \collatz.iter[11] ;
 wire \collatz.iter[120] ;
 wire \collatz.iter[121] ;
 wire \collatz.iter[122] ;
 wire \collatz.iter[123] ;
 wire \collatz.iter[124] ;
 wire \collatz.iter[125] ;
 wire \collatz.iter[126] ;
 wire \collatz.iter[127] ;
 wire \collatz.iter[128] ;
 wire \collatz.iter[129] ;
 wire \collatz.iter[12] ;
 wire \collatz.iter[130] ;
 wire \collatz.iter[131] ;
 wire \collatz.iter[132] ;
 wire \collatz.iter[133] ;
 wire \collatz.iter[134] ;
 wire \collatz.iter[135] ;
 wire \collatz.iter[136] ;
 wire \collatz.iter[137] ;
 wire \collatz.iter[138] ;
 wire \collatz.iter[139] ;
 wire \collatz.iter[13] ;
 wire \collatz.iter[140] ;
 wire \collatz.iter[141] ;
 wire \collatz.iter[142] ;
 wire \collatz.iter[143] ;
 wire \collatz.iter[14] ;
 wire \collatz.iter[15] ;
 wire \collatz.iter[16] ;
 wire \collatz.iter[17] ;
 wire \collatz.iter[18] ;
 wire \collatz.iter[19] ;
 wire \collatz.iter[1] ;
 wire \collatz.iter[20] ;
 wire \collatz.iter[21] ;
 wire \collatz.iter[22] ;
 wire \collatz.iter[23] ;
 wire \collatz.iter[24] ;
 wire \collatz.iter[25] ;
 wire \collatz.iter[26] ;
 wire \collatz.iter[27] ;
 wire \collatz.iter[28] ;
 wire \collatz.iter[29] ;
 wire \collatz.iter[2] ;
 wire \collatz.iter[30] ;
 wire \collatz.iter[31] ;
 wire \collatz.iter[32] ;
 wire \collatz.iter[33] ;
 wire \collatz.iter[34] ;
 wire \collatz.iter[35] ;
 wire \collatz.iter[36] ;
 wire \collatz.iter[37] ;
 wire \collatz.iter[38] ;
 wire \collatz.iter[39] ;
 wire \collatz.iter[3] ;
 wire \collatz.iter[40] ;
 wire \collatz.iter[41] ;
 wire \collatz.iter[42] ;
 wire \collatz.iter[43] ;
 wire \collatz.iter[44] ;
 wire \collatz.iter[45] ;
 wire \collatz.iter[46] ;
 wire \collatz.iter[47] ;
 wire \collatz.iter[48] ;
 wire \collatz.iter[49] ;
 wire \collatz.iter[4] ;
 wire \collatz.iter[50] ;
 wire \collatz.iter[51] ;
 wire \collatz.iter[52] ;
 wire \collatz.iter[53] ;
 wire \collatz.iter[54] ;
 wire \collatz.iter[55] ;
 wire \collatz.iter[56] ;
 wire \collatz.iter[57] ;
 wire \collatz.iter[58] ;
 wire \collatz.iter[59] ;
 wire \collatz.iter[5] ;
 wire \collatz.iter[60] ;
 wire \collatz.iter[61] ;
 wire \collatz.iter[62] ;
 wire \collatz.iter[63] ;
 wire \collatz.iter[64] ;
 wire \collatz.iter[65] ;
 wire \collatz.iter[66] ;
 wire \collatz.iter[67] ;
 wire \collatz.iter[68] ;
 wire \collatz.iter[69] ;
 wire \collatz.iter[6] ;
 wire \collatz.iter[70] ;
 wire \collatz.iter[71] ;
 wire \collatz.iter[72] ;
 wire \collatz.iter[73] ;
 wire \collatz.iter[74] ;
 wire \collatz.iter[75] ;
 wire \collatz.iter[76] ;
 wire \collatz.iter[77] ;
 wire \collatz.iter[78] ;
 wire \collatz.iter[79] ;
 wire \collatz.iter[7] ;
 wire \collatz.iter[80] ;
 wire \collatz.iter[81] ;
 wire \collatz.iter[82] ;
 wire \collatz.iter[83] ;
 wire \collatz.iter[84] ;
 wire \collatz.iter[85] ;
 wire \collatz.iter[86] ;
 wire \collatz.iter[87] ;
 wire \collatz.iter[88] ;
 wire \collatz.iter[89] ;
 wire \collatz.iter[8] ;
 wire \collatz.iter[90] ;
 wire \collatz.iter[91] ;
 wire \collatz.iter[92] ;
 wire \collatz.iter[93] ;
 wire \collatz.iter[94] ;
 wire \collatz.iter[95] ;
 wire \collatz.iter[96] ;
 wire \collatz.iter[97] ;
 wire \collatz.iter[98] ;
 wire \collatz.iter[99] ;
 wire \collatz.iter[9] ;
 wire \collatz.orbit_len[0] ;
 wire \collatz.orbit_len[10] ;
 wire \collatz.orbit_len[11] ;
 wire \collatz.orbit_len[12] ;
 wire \collatz.orbit_len[13] ;
 wire \collatz.orbit_len[14] ;
 wire \collatz.orbit_len[15] ;
 wire \collatz.orbit_len[1] ;
 wire \collatz.orbit_len[2] ;
 wire \collatz.orbit_len[3] ;
 wire \collatz.orbit_len[4] ;
 wire \collatz.orbit_len[5] ;
 wire \collatz.orbit_len[6] ;
 wire \collatz.orbit_len[7] ;
 wire \collatz.orbit_len[8] ;
 wire \collatz.orbit_len[9] ;
 wire \collatz.path_record_h16[0] ;
 wire \collatz.path_record_h16[10] ;
 wire \collatz.path_record_h16[11] ;
 wire \collatz.path_record_h16[12] ;
 wire \collatz.path_record_h16[13] ;
 wire \collatz.path_record_h16[14] ;
 wire \collatz.path_record_h16[15] ;
 wire \collatz.path_record_h16[1] ;
 wire \collatz.path_record_h16[2] ;
 wire \collatz.path_record_h16[3] ;
 wire \collatz.path_record_h16[4] ;
 wire \collatz.path_record_h16[5] ;
 wire \collatz.path_record_h16[6] ;
 wire \collatz.path_record_h16[7] ;
 wire \collatz.path_record_h16[8] ;
 wire \collatz.path_record_h16[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_1 _4386_ (.A(\collatz.comp ),
    .X(_3161_));
 sg13g2_inv_1 _4387_ (.Y(_3171_),
    .A(\collatz.orbit_len[5] ));
 sg13g2_inv_1 _4388_ (.Y(_3181_),
    .A(\collatz.orbit_len[3] ));
 sg13g2_buf_1 _4389_ (.A(\collatz.orbit_len[1] ),
    .X(_3191_));
 sg13g2_buf_1 _4390_ (.A(\collatz.orbit_len[0] ),
    .X(_3201_));
 sg13g2_buf_1 _4391_ (.A(\collatz.orbit_len[2] ),
    .X(_3211_));
 sg13g2_nand3_1 _4392_ (.B(_3201_),
    .C(_3211_),
    .A(_3191_),
    .Y(_3220_));
 sg13g2_nor2_1 _4393_ (.A(_3181_),
    .B(_3220_),
    .Y(_3231_));
 sg13g2_nand2_1 _4394_ (.Y(_3241_),
    .A(\collatz.orbit_len[4] ),
    .B(_3231_));
 sg13g2_nor2_1 _4395_ (.A(_3171_),
    .B(_3241_),
    .Y(_3251_));
 sg13g2_buf_1 _4396_ (.A(\collatz.orbit_len[7] ),
    .X(_3261_));
 sg13g2_buf_1 _4397_ (.A(\collatz.orbit_len[8] ),
    .X(_3271_));
 sg13g2_and3_1 _4398_ (.X(_3280_),
    .A(_3261_),
    .B(\collatz.orbit_len[9] ),
    .C(_3271_));
 sg13g2_buf_1 _4399_ (.A(_3280_),
    .X(_3290_));
 sg13g2_buf_1 _4400_ (.A(\collatz.orbit_len[6] ),
    .X(_3300_));
 sg13g2_buf_1 _4401_ (.A(\collatz.orbit_len[10] ),
    .X(_3310_));
 sg13g2_buf_1 _4402_ (.A(\collatz.orbit_len[14] ),
    .X(_3320_));
 sg13g2_nand4_1 _4403_ (.B(_3310_),
    .C(_3320_),
    .A(_3300_),
    .Y(_3330_),
    .D(\collatz.orbit_len[15] ));
 sg13g2_buf_1 _4404_ (.A(\collatz.orbit_len[11] ),
    .X(_3340_));
 sg13g2_buf_1 _4405_ (.A(\collatz.orbit_len[12] ),
    .X(_3349_));
 sg13g2_nand3_1 _4406_ (.B(\collatz.orbit_len[13] ),
    .C(_3349_),
    .A(_3340_),
    .Y(_3359_));
 sg13g2_nor2_1 _4407_ (.A(_3330_),
    .B(_3359_),
    .Y(_3369_));
 sg13g2_nand3_1 _4408_ (.B(_3290_),
    .C(_3369_),
    .A(_3251_),
    .Y(_3379_));
 sg13g2_buf_1 _4409_ (.A(\collatz.iter[116] ),
    .X(_3389_));
 sg13g2_buf_2 _4410_ (.A(\collatz.iter[118] ),
    .X(_3399_));
 sg13g2_nor2_1 _4411_ (.A(net322),
    .B(_3399_),
    .Y(_3409_));
 sg13g2_buf_2 _4412_ (.A(\collatz.iter[123] ),
    .X(_3419_));
 sg13g2_buf_2 _4413_ (.A(\collatz.iter[125] ),
    .X(_3429_));
 sg13g2_nor2_2 _4414_ (.A(_3419_),
    .B(_3429_),
    .Y(_3438_));
 sg13g2_buf_2 _4415_ (.A(\collatz.iter[103] ),
    .X(_3447_));
 sg13g2_buf_2 _4416_ (.A(\collatz.iter[105] ),
    .X(_3456_));
 sg13g2_nor2_2 _4417_ (.A(net321),
    .B(_3456_),
    .Y(_3464_));
 sg13g2_buf_1 _4418_ (.A(\collatz.iter[117] ),
    .X(_3473_));
 sg13g2_buf_1 _4419_ (.A(_3473_),
    .X(_3481_));
 sg13g2_buf_1 _4420_ (.A(\collatz.iter[119] ),
    .X(_3489_));
 sg13g2_buf_1 _4421_ (.A(_3489_),
    .X(_3500_));
 sg13g2_nor2_1 _4422_ (.A(_3481_),
    .B(net260),
    .Y(_3511_));
 sg13g2_nand4_1 _4423_ (.B(_3438_),
    .C(_3464_),
    .A(_3409_),
    .Y(_3522_),
    .D(_3511_));
 sg13g2_buf_2 _4424_ (.A(\collatz.iter[39] ),
    .X(_3533_));
 sg13g2_buf_2 _4425_ (.A(\collatz.iter[41] ),
    .X(_3544_));
 sg13g2_nor2_2 _4426_ (.A(_3533_),
    .B(_3544_),
    .Y(_3555_));
 sg13g2_buf_8 _4427_ (.A(\collatz.iter[107] ),
    .X(_3566_));
 sg13g2_buf_1 _4428_ (.A(\collatz.iter[109] ),
    .X(_3577_));
 sg13g2_nor2_2 _4429_ (.A(_3566_),
    .B(_3577_),
    .Y(_3588_));
 sg13g2_buf_2 _4430_ (.A(\collatz.iter[122] ),
    .X(_3599_));
 sg13g2_buf_2 _4431_ (.A(\collatz.iter[124] ),
    .X(_3610_));
 sg13g2_nor2_2 _4432_ (.A(_3599_),
    .B(_3610_),
    .Y(_3621_));
 sg13g2_buf_2 _4433_ (.A(\collatz.iter[57] ),
    .X(_3632_));
 sg13g2_buf_1 _4434_ (.A(\collatz.iter[59] ),
    .X(_3641_));
 sg13g2_nor2_2 _4435_ (.A(_3632_),
    .B(net320),
    .Y(_3650_));
 sg13g2_nand4_1 _4436_ (.B(_3588_),
    .C(_3621_),
    .A(_3555_),
    .Y(_3659_),
    .D(_3650_));
 sg13g2_buf_2 _4437_ (.A(\collatz.iter[10] ),
    .X(_3667_));
 sg13g2_buf_2 _4438_ (.A(\collatz.iter[12] ),
    .X(_3676_));
 sg13g2_nor2_1 _4439_ (.A(_3667_),
    .B(_3676_),
    .Y(_3684_));
 sg13g2_buf_1 _4440_ (.A(\collatz.iter[48] ),
    .X(_3690_));
 sg13g2_buf_1 _4441_ (.A(\collatz.iter[50] ),
    .X(_3691_));
 sg13g2_nor2_1 _4442_ (.A(net319),
    .B(net318),
    .Y(_3692_));
 sg13g2_buf_1 _4443_ (.A(\collatz.iter[72] ),
    .X(_3693_));
 sg13g2_buf_1 _4444_ (.A(\collatz.iter[74] ),
    .X(_3694_));
 sg13g2_nor2_1 _4445_ (.A(net317),
    .B(_3694_),
    .Y(_3695_));
 sg13g2_buf_8 _4446_ (.A(\collatz.iter[100] ),
    .X(_3696_));
 sg13g2_buf_8 _4447_ (.A(\collatz.iter[102] ),
    .X(_3697_));
 sg13g2_nor2_2 _4448_ (.A(_3696_),
    .B(_3697_),
    .Y(_3698_));
 sg13g2_nand4_1 _4449_ (.B(_3692_),
    .C(_3695_),
    .A(_3684_),
    .Y(_3699_),
    .D(_3698_));
 sg13g2_buf_1 _4450_ (.A(\collatz.iter[80] ),
    .X(_3700_));
 sg13g2_buf_1 _4451_ (.A(\collatz.iter[82] ),
    .X(_3701_));
 sg13g2_nor2_1 _4452_ (.A(net315),
    .B(_3701_),
    .Y(_3702_));
 sg13g2_buf_1 _4453_ (.A(\collatz.iter[44] ),
    .X(_3703_));
 sg13g2_buf_1 _4454_ (.A(net313),
    .X(_3704_));
 sg13g2_buf_1 _4455_ (.A(\collatz.iter[46] ),
    .X(_3705_));
 sg13g2_buf_1 _4456_ (.A(net312),
    .X(_3706_));
 sg13g2_nor2_1 _4457_ (.A(_3704_),
    .B(net258),
    .Y(_3707_));
 sg13g2_buf_1 _4458_ (.A(\collatz.iter[2] ),
    .X(_3708_));
 sg13g2_buf_1 _4459_ (.A(_3708_),
    .X(_3709_));
 sg13g2_buf_1 _4460_ (.A(\collatz.iter[4] ),
    .X(_3710_));
 sg13g2_buf_1 _4461_ (.A(_3710_),
    .X(_3711_));
 sg13g2_or2_1 _4462_ (.X(_3712_),
    .B(net256),
    .A(net257));
 sg13g2_buf_2 _4463_ (.A(\collatz.iter[5] ),
    .X(_3713_));
 sg13g2_buf_1 _4464_ (.A(\collatz.iter[7] ),
    .X(_3714_));
 sg13g2_or2_1 _4465_ (.X(_3715_),
    .B(_3714_),
    .A(_3713_));
 sg13g2_buf_1 _4466_ (.A(_3715_),
    .X(_3716_));
 sg13g2_nor2_1 _4467_ (.A(_3712_),
    .B(_3716_),
    .Y(_3717_));
 sg13g2_nand3_1 _4468_ (.B(_3707_),
    .C(_3717_),
    .A(_3702_),
    .Y(_3718_));
 sg13g2_or4_1 _4469_ (.A(_3522_),
    .B(_3659_),
    .C(_3699_),
    .D(_3718_),
    .X(_3719_));
 sg13g2_buf_1 _4470_ (.A(\collatz.iter[92] ),
    .X(_3720_));
 sg13g2_buf_8 _4471_ (.A(\collatz.iter[94] ),
    .X(_3721_));
 sg13g2_nor2_1 _4472_ (.A(net311),
    .B(net310),
    .Y(_3722_));
 sg13g2_buf_8 _4473_ (.A(\collatz.iter[128] ),
    .X(_3723_));
 sg13g2_buf_1 _4474_ (.A(\collatz.iter[130] ),
    .X(_3724_));
 sg13g2_nor2_2 _4475_ (.A(_3723_),
    .B(net309),
    .Y(_3725_));
 sg13g2_buf_1 _4476_ (.A(\collatz.iter[23] ),
    .X(_3726_));
 sg13g2_buf_1 _4477_ (.A(_3726_),
    .X(_3727_));
 sg13g2_buf_1 _4478_ (.A(\collatz.iter[53] ),
    .X(_3728_));
 sg13g2_buf_1 _4479_ (.A(net307),
    .X(_3729_));
 sg13g2_buf_1 _4480_ (.A(\collatz.iter[55] ),
    .X(_3730_));
 sg13g2_buf_1 _4481_ (.A(net306),
    .X(_3731_));
 sg13g2_buf_1 _4482_ (.A(\collatz.iter[63] ),
    .X(_3732_));
 sg13g2_buf_1 _4483_ (.A(_3732_),
    .X(_3733_));
 sg13g2_buf_1 _4484_ (.A(net252),
    .X(_3734_));
 sg13g2_nor4_1 _4485_ (.A(_3727_),
    .B(_3729_),
    .C(_3731_),
    .D(net116),
    .Y(_3735_));
 sg13g2_nand3_1 _4486_ (.B(_3725_),
    .C(_3735_),
    .A(_3722_),
    .Y(_3736_));
 sg13g2_buf_1 _4487_ (.A(\collatz.iter[40] ),
    .X(_3737_));
 sg13g2_buf_1 _4488_ (.A(\collatz.iter[42] ),
    .X(_3738_));
 sg13g2_nor2_1 _4489_ (.A(net305),
    .B(_3738_),
    .Y(_3739_));
 sg13g2_buf_1 _4490_ (.A(\collatz.iter[52] ),
    .X(_3740_));
 sg13g2_buf_1 _4491_ (.A(\collatz.iter[54] ),
    .X(_3741_));
 sg13g2_nor2_2 _4492_ (.A(net303),
    .B(net302),
    .Y(_3742_));
 sg13g2_buf_2 _4493_ (.A(\collatz.iter[104] ),
    .X(_3743_));
 sg13g2_buf_1 _4494_ (.A(\collatz.iter[106] ),
    .X(_3744_));
 sg13g2_nor2_1 _4495_ (.A(_3743_),
    .B(net301),
    .Y(_3745_));
 sg13g2_buf_2 _4496_ (.A(\collatz.iter[129] ),
    .X(_3746_));
 sg13g2_buf_2 _4497_ (.A(\collatz.iter[131] ),
    .X(_3747_));
 sg13g2_nor2_1 _4498_ (.A(_3746_),
    .B(_3747_),
    .Y(_3748_));
 sg13g2_buf_2 _4499_ (.A(_3748_),
    .X(_3749_));
 sg13g2_nand4_1 _4500_ (.B(_3742_),
    .C(_3745_),
    .A(_3739_),
    .Y(_3750_),
    .D(_3749_));
 sg13g2_buf_8 _4501_ (.A(\collatz.iter[9] ),
    .X(_3751_));
 sg13g2_buf_1 _4502_ (.A(_3751_),
    .X(_3752_));
 sg13g2_buf_8 _4503_ (.A(\collatz.iter[11] ),
    .X(_3753_));
 sg13g2_buf_2 _4504_ (.A(\collatz.iter[13] ),
    .X(_3754_));
 sg13g2_buf_8 _4505_ (.A(_3754_),
    .X(_3755_));
 sg13g2_nor3_1 _4506_ (.A(net251),
    .B(net300),
    .C(net250),
    .Y(_3756_));
 sg13g2_buf_2 _4507_ (.A(\collatz.iter[3] ),
    .X(_3757_));
 sg13g2_buf_1 _4508_ (.A(_3757_),
    .X(_3758_));
 sg13g2_buf_1 _4509_ (.A(\collatz.iter[22] ),
    .X(_3759_));
 sg13g2_buf_1 _4510_ (.A(_3759_),
    .X(_3760_));
 sg13g2_buf_1 _4511_ (.A(net248),
    .X(_3761_));
 sg13g2_buf_8 _4512_ (.A(\collatz.iter[29] ),
    .X(_3762_));
 sg13g2_buf_1 _4513_ (.A(_3762_),
    .X(_3763_));
 sg13g2_buf_8 _4514_ (.A(\collatz.iter[31] ),
    .X(_3764_));
 sg13g2_buf_1 _4515_ (.A(_3764_),
    .X(_3765_));
 sg13g2_nor4_1 _4516_ (.A(net249),
    .B(net115),
    .C(net247),
    .D(net246),
    .Y(_3766_));
 sg13g2_buf_1 _4517_ (.A(\collatz.iter[60] ),
    .X(_3767_));
 sg13g2_buf_1 _4518_ (.A(\collatz.iter[62] ),
    .X(_3768_));
 sg13g2_buf_1 _4519_ (.A(\collatz.iter[64] ),
    .X(_3769_));
 sg13g2_nor3_2 _4520_ (.A(net299),
    .B(_3768_),
    .C(net298),
    .Y(_3770_));
 sg13g2_buf_1 _4521_ (.A(\collatz.iter[132] ),
    .X(_3771_));
 sg13g2_buf_1 _4522_ (.A(\collatz.iter[134] ),
    .X(_3772_));
 sg13g2_or2_1 _4523_ (.X(_3773_),
    .B(_3772_),
    .A(net297));
 sg13g2_buf_1 _4524_ (.A(_3773_),
    .X(_3774_));
 sg13g2_buf_8 _4525_ (.A(\collatz.iter[95] ),
    .X(_3775_));
 sg13g2_buf_1 _4526_ (.A(\collatz.iter[97] ),
    .X(_3776_));
 sg13g2_nor2_1 _4527_ (.A(_3775_),
    .B(net296),
    .Y(_3777_));
 sg13g2_nor2b_1 _4528_ (.A(_3774_),
    .B_N(_3777_),
    .Y(_3778_));
 sg13g2_nand4_1 _4529_ (.B(_3766_),
    .C(_3770_),
    .A(_3756_),
    .Y(_3779_),
    .D(_3778_));
 sg13g2_nor4_1 _4530_ (.A(_3719_),
    .B(_3736_),
    .C(_3750_),
    .D(_3779_),
    .Y(_3780_));
 sg13g2_buf_1 _4531_ (.A(\collatz.iter[66] ),
    .X(_3781_));
 sg13g2_buf_1 _4532_ (.A(_3781_),
    .X(_3782_));
 sg13g2_buf_1 _4533_ (.A(_3782_),
    .X(_3783_));
 sg13g2_buf_1 _4534_ (.A(\collatz.iter[71] ),
    .X(_3784_));
 sg13g2_buf_1 _4535_ (.A(net295),
    .X(_3785_));
 sg13g2_buf_2 _4536_ (.A(\collatz.iter[90] ),
    .X(_3786_));
 sg13g2_buf_1 _4537_ (.A(_3786_),
    .X(_3787_));
 sg13g2_buf_8 _4538_ (.A(\collatz.iter[99] ),
    .X(_3788_));
 sg13g2_buf_1 _4539_ (.A(_3788_),
    .X(_3789_));
 sg13g2_nor4_1 _4540_ (.A(_3783_),
    .B(_3785_),
    .C(_3787_),
    .D(_3789_),
    .Y(_3790_));
 sg13g2_buf_8 _4541_ (.A(\collatz.iter[27] ),
    .X(_3791_));
 sg13g2_buf_1 _4542_ (.A(_3791_),
    .X(_3792_));
 sg13g2_buf_2 _4543_ (.A(\collatz.iter[30] ),
    .X(_3793_));
 sg13g2_buf_1 _4544_ (.A(_3793_),
    .X(_3794_));
 sg13g2_buf_8 _4545_ (.A(\collatz.iter[35] ),
    .X(_3795_));
 sg13g2_buf_1 _4546_ (.A(_3795_),
    .X(_3796_));
 sg13g2_buf_2 _4547_ (.A(\collatz.iter[67] ),
    .X(_3797_));
 sg13g2_buf_1 _4548_ (.A(_3797_),
    .X(_3798_));
 sg13g2_nor4_1 _4549_ (.A(_3792_),
    .B(_3794_),
    .C(net239),
    .D(_3798_),
    .Y(_3799_));
 sg13g2_nand2_1 _4550_ (.Y(_3800_),
    .A(_3790_),
    .B(_3799_));
 sg13g2_buf_8 _4551_ (.A(\collatz.iter[86] ),
    .X(_3801_));
 sg13g2_buf_8 _4552_ (.A(\collatz.iter[88] ),
    .X(_3802_));
 sg13g2_nor2_1 _4553_ (.A(_3801_),
    .B(_3802_),
    .Y(_3803_));
 sg13g2_buf_2 _4554_ (.A(\collatz.iter[112] ),
    .X(_3804_));
 sg13g2_buf_1 _4555_ (.A(\collatz.iter[114] ),
    .X(_3805_));
 sg13g2_nor2_1 _4556_ (.A(_3804_),
    .B(_3805_),
    .Y(_3806_));
 sg13g2_buf_2 _4557_ (.A(_3806_),
    .X(_3807_));
 sg13g2_buf_8 _4558_ (.A(\collatz.iter[6] ),
    .X(_3808_));
 sg13g2_buf_1 _4559_ (.A(_3808_),
    .X(_3809_));
 sg13g2_buf_2 _4560_ (.A(\collatz.iter[8] ),
    .X(_3810_));
 sg13g2_buf_8 _4561_ (.A(_3810_),
    .X(_3811_));
 sg13g2_or2_1 _4562_ (.X(_3812_),
    .B(net236),
    .A(net237));
 sg13g2_buf_8 _4563_ (.A(\collatz.iter[96] ),
    .X(_3813_));
 sg13g2_buf_1 _4564_ (.A(\collatz.iter[98] ),
    .X(_3814_));
 sg13g2_buf_1 _4565_ (.A(_3814_),
    .X(_3815_));
 sg13g2_or2_1 _4566_ (.X(_3816_),
    .B(net235),
    .A(_3813_));
 sg13g2_buf_1 _4567_ (.A(_3816_),
    .X(_3817_));
 sg13g2_nor2_1 _4568_ (.A(_3812_),
    .B(_3817_),
    .Y(_3818_));
 sg13g2_nand3_1 _4569_ (.B(_3807_),
    .C(_3818_),
    .A(_3803_),
    .Y(_3819_));
 sg13g2_buf_1 _4570_ (.A(\collatz.iter[56] ),
    .X(_3820_));
 sg13g2_buf_1 _4571_ (.A(\collatz.iter[58] ),
    .X(_3821_));
 sg13g2_nor2_1 _4572_ (.A(net294),
    .B(_3821_),
    .Y(_3822_));
 sg13g2_buf_1 _4573_ (.A(\collatz.iter[18] ),
    .X(_3823_));
 sg13g2_nor2_2 _4574_ (.A(\collatz.iter[16] ),
    .B(net292),
    .Y(_3824_));
 sg13g2_buf_1 _4575_ (.A(\collatz.iter[26] ),
    .X(_3825_));
 sg13g2_buf_8 _4576_ (.A(\collatz.iter[28] ),
    .X(_3826_));
 sg13g2_nor2_1 _4577_ (.A(net291),
    .B(_3826_),
    .Y(_3827_));
 sg13g2_nand3_1 _4578_ (.B(_3824_),
    .C(_3827_),
    .A(_3822_),
    .Y(_3828_));
 sg13g2_nor3_1 _4579_ (.A(_3800_),
    .B(_3819_),
    .C(_3828_),
    .Y(_3829_));
 sg13g2_buf_2 _4580_ (.A(\collatz.iter[140] ),
    .X(_3830_));
 sg13g2_inv_1 _4581_ (.Y(_3831_),
    .A(_3830_));
 sg13g2_buf_2 _4582_ (.A(\collatz.iter[142] ),
    .X(_3832_));
 sg13g2_inv_1 _4583_ (.Y(_3833_),
    .A(_3832_));
 sg13g2_buf_8 _4584_ (.A(\collatz.iter[79] ),
    .X(_3834_));
 sg13g2_nor2_1 _4585_ (.A(\collatz.iter[77] ),
    .B(_3834_),
    .Y(_3835_));
 sg13g2_buf_2 _4586_ (.A(\collatz.iter[15] ),
    .X(_3836_));
 sg13g2_buf_1 _4587_ (.A(_3836_),
    .X(_3837_));
 sg13g2_buf_1 _4588_ (.A(\collatz.iter[17] ),
    .X(_3838_));
 sg13g2_buf_1 _4589_ (.A(net290),
    .X(_3839_));
 sg13g2_buf_1 _4590_ (.A(\collatz.iter[36] ),
    .X(_3840_));
 sg13g2_buf_1 _4591_ (.A(net289),
    .X(_3841_));
 sg13g2_buf_8 _4592_ (.A(\collatz.iter[38] ),
    .X(_3842_));
 sg13g2_buf_1 _4593_ (.A(net288),
    .X(_3843_));
 sg13g2_nor4_1 _4594_ (.A(_3837_),
    .B(_3839_),
    .C(_3841_),
    .D(net231),
    .Y(_3844_));
 sg13g2_nand4_1 _4595_ (.B(_3833_),
    .C(_3835_),
    .A(_3831_),
    .Y(_3845_),
    .D(_3844_));
 sg13g2_buf_1 _4596_ (.A(\collatz.iter[68] ),
    .X(_3846_));
 sg13g2_buf_2 _4597_ (.A(\collatz.iter[70] ),
    .X(_3847_));
 sg13g2_nor2_2 _4598_ (.A(_3846_),
    .B(_3847_),
    .Y(_3848_));
 sg13g2_buf_1 _4599_ (.A(\collatz.iter[108] ),
    .X(_3849_));
 sg13g2_buf_1 _4600_ (.A(\collatz.iter[110] ),
    .X(_3850_));
 sg13g2_nor2_1 _4601_ (.A(net286),
    .B(_3850_),
    .Y(_3851_));
 sg13g2_buf_8 _4602_ (.A(\collatz.iter[83] ),
    .X(_3852_));
 sg13g2_buf_8 _4603_ (.A(\collatz.iter[85] ),
    .X(_3853_));
 sg13g2_nor2_2 _4604_ (.A(_3852_),
    .B(_3853_),
    .Y(_3854_));
 sg13g2_buf_1 _4605_ (.A(\collatz.iter[137] ),
    .X(_3855_));
 sg13g2_buf_1 _4606_ (.A(\collatz.iter[139] ),
    .X(_3856_));
 sg13g2_nor2_1 _4607_ (.A(_3855_),
    .B(_3856_),
    .Y(_3857_));
 sg13g2_nand4_1 _4608_ (.B(_3851_),
    .C(_3854_),
    .A(_3848_),
    .Y(_3858_),
    .D(_3857_));
 sg13g2_buf_1 _4609_ (.A(\collatz.iter[1] ),
    .X(_3859_));
 sg13g2_buf_1 _4610_ (.A(\collatz.iter[0] ),
    .X(_3860_));
 sg13g2_inv_2 _4611_ (.Y(_3861_),
    .A(net283));
 sg13g2_buf_1 _4612_ (.A(_3861_),
    .X(_3862_));
 sg13g2_buf_1 _4613_ (.A(_3862_),
    .X(_3863_));
 sg13g2_buf_1 _4614_ (.A(\collatz.iter[65] ),
    .X(_3864_));
 sg13g2_buf_1 _4615_ (.A(net282),
    .X(_3865_));
 sg13g2_buf_2 _4616_ (.A(\collatz.iter[69] ),
    .X(_3866_));
 sg13g2_buf_1 _4617_ (.A(_3866_),
    .X(_3867_));
 sg13g2_buf_1 _4618_ (.A(\collatz.iter[138] ),
    .X(_3868_));
 sg13g2_buf_1 _4619_ (.A(_3868_),
    .X(_3869_));
 sg13g2_buf_1 _4620_ (.A(\collatz.iter[141] ),
    .X(_3870_));
 sg13g2_nor4_1 _4621_ (.A(_3865_),
    .B(_3867_),
    .C(net228),
    .D(_3870_),
    .Y(_3871_));
 sg13g2_buf_1 _4622_ (.A(\collatz.iter[73] ),
    .X(_3872_));
 sg13g2_buf_2 _4623_ (.A(\collatz.iter[75] ),
    .X(_3873_));
 sg13g2_buf_8 _4624_ (.A(_3873_),
    .X(_3874_));
 sg13g2_nor2_1 _4625_ (.A(_3872_),
    .B(net227),
    .Y(_3875_));
 sg13g2_nand4_1 _4626_ (.B(net84),
    .C(_3871_),
    .A(net284),
    .Y(_3876_),
    .D(_3875_));
 sg13g2_buf_1 _4627_ (.A(\collatz.iter[133] ),
    .X(_3877_));
 sg13g2_buf_1 _4628_ (.A(\collatz.iter[135] ),
    .X(_3878_));
 sg13g2_nor2_1 _4629_ (.A(_3877_),
    .B(_3878_),
    .Y(_3879_));
 sg13g2_buf_1 _4630_ (.A(\collatz.iter[49] ),
    .X(_3880_));
 sg13g2_buf_2 _4631_ (.A(\collatz.iter[51] ),
    .X(_3881_));
 sg13g2_nor2_2 _4632_ (.A(_3880_),
    .B(_3881_),
    .Y(_3882_));
 sg13g2_buf_2 _4633_ (.A(\collatz.iter[32] ),
    .X(_3883_));
 sg13g2_buf_8 _4634_ (.A(_3883_),
    .X(_3884_));
 sg13g2_buf_2 _4635_ (.A(\collatz.iter[34] ),
    .X(_3885_));
 sg13g2_buf_1 _4636_ (.A(_3885_),
    .X(_3886_));
 sg13g2_nor2_1 _4637_ (.A(net226),
    .B(net225),
    .Y(_3887_));
 sg13g2_buf_2 _4638_ (.A(\collatz.iter[19] ),
    .X(_3888_));
 sg13g2_nor2_2 _4639_ (.A(_3888_),
    .B(\collatz.iter[21] ),
    .Y(_3889_));
 sg13g2_nand4_1 _4640_ (.B(_3882_),
    .C(_3887_),
    .A(_3879_),
    .Y(_3890_),
    .D(_3889_));
 sg13g2_nor4_1 _4641_ (.A(_3845_),
    .B(_3858_),
    .C(_3876_),
    .D(_3890_),
    .Y(_3891_));
 sg13g2_buf_2 _4642_ (.A(\collatz.iter[43] ),
    .X(_3892_));
 sg13g2_buf_2 _4643_ (.A(\collatz.iter[45] ),
    .X(_3893_));
 sg13g2_buf_2 _4644_ (.A(\collatz.iter[47] ),
    .X(_3894_));
 sg13g2_nor3_1 _4645_ (.A(_3892_),
    .B(_3893_),
    .C(_3894_),
    .Y(_3895_));
 sg13g2_buf_8 _4646_ (.A(\collatz.iter[89] ),
    .X(_3896_));
 sg13g2_buf_1 _4647_ (.A(\collatz.iter[91] ),
    .X(_3897_));
 sg13g2_buf_1 _4648_ (.A(_3897_),
    .X(_3898_));
 sg13g2_buf_8 _4649_ (.A(\collatz.iter[93] ),
    .X(_3899_));
 sg13g2_nor3_1 _4650_ (.A(_3896_),
    .B(net224),
    .C(_3899_),
    .Y(_3900_));
 sg13g2_buf_2 _4651_ (.A(\collatz.iter[111] ),
    .X(_3901_));
 sg13g2_buf_1 _4652_ (.A(_3901_),
    .X(_3902_));
 sg13g2_buf_1 _4653_ (.A(\collatz.iter[113] ),
    .X(_3903_));
 sg13g2_buf_1 _4654_ (.A(\collatz.iter[115] ),
    .X(_3904_));
 sg13g2_nor3_2 _4655_ (.A(net223),
    .B(_3903_),
    .C(net279),
    .Y(_3905_));
 sg13g2_buf_1 _4656_ (.A(\collatz.iter[14] ),
    .X(_3906_));
 sg13g2_buf_1 _4657_ (.A(net278),
    .X(_3907_));
 sg13g2_buf_1 _4658_ (.A(\collatz.iter[20] ),
    .X(_3908_));
 sg13g2_buf_1 _4659_ (.A(_3908_),
    .X(_3909_));
 sg13g2_buf_1 _4660_ (.A(net221),
    .X(_3910_));
 sg13g2_buf_1 _4661_ (.A(\collatz.iter[25] ),
    .X(_3911_));
 sg13g2_buf_1 _4662_ (.A(net277),
    .X(_3912_));
 sg13g2_nor3_1 _4663_ (.A(net222),
    .B(net112),
    .C(_3912_),
    .Y(_3913_));
 sg13g2_nand4_1 _4664_ (.B(_3900_),
    .C(_3905_),
    .A(_3895_),
    .Y(_3914_),
    .D(_3913_));
 sg13g2_buf_1 _4665_ (.A(\collatz.iter[81] ),
    .X(_3915_));
 sg13g2_buf_1 _4666_ (.A(_3915_),
    .X(_3916_));
 sg13g2_buf_1 _4667_ (.A(net219),
    .X(_3917_));
 sg13g2_buf_1 _4668_ (.A(\collatz.iter[84] ),
    .X(_3918_));
 sg13g2_buf_1 _4669_ (.A(net276),
    .X(_3919_));
 sg13g2_buf_8 _4670_ (.A(\collatz.iter[101] ),
    .X(_3920_));
 sg13g2_buf_1 _4671_ (.A(_3920_),
    .X(_3921_));
 sg13g2_buf_1 _4672_ (.A(\collatz.iter[143] ),
    .X(_3922_));
 sg13g2_nor4_1 _4673_ (.A(_3917_),
    .B(_3919_),
    .C(_3921_),
    .D(_3922_),
    .Y(_3923_));
 sg13g2_buf_2 _4674_ (.A(\collatz.iter[24] ),
    .X(_3924_));
 sg13g2_buf_1 _4675_ (.A(_3924_),
    .X(_3925_));
 sg13g2_buf_1 _4676_ (.A(_3925_),
    .X(_3926_));
 sg13g2_buf_1 _4677_ (.A(\collatz.iter[33] ),
    .X(_3927_));
 sg13g2_buf_1 _4678_ (.A(_3927_),
    .X(_3928_));
 sg13g2_buf_8 _4679_ (.A(\collatz.iter[37] ),
    .X(_3929_));
 sg13g2_buf_1 _4680_ (.A(_3929_),
    .X(_3930_));
 sg13g2_buf_1 _4681_ (.A(\collatz.iter[61] ),
    .X(_3931_));
 sg13g2_buf_1 _4682_ (.A(net275),
    .X(_3932_));
 sg13g2_nor4_1 _4683_ (.A(net110),
    .B(net215),
    .C(net214),
    .D(_3932_),
    .Y(_3933_));
 sg13g2_buf_8 _4684_ (.A(\collatz.iter[121] ),
    .X(_3934_));
 sg13g2_buf_1 _4685_ (.A(_3934_),
    .X(_3935_));
 sg13g2_buf_8 _4686_ (.A(\collatz.iter[120] ),
    .X(_3936_));
 sg13g2_buf_1 _4687_ (.A(_3936_),
    .X(_3937_));
 sg13g2_buf_1 _4688_ (.A(\collatz.iter[127] ),
    .X(_3938_));
 sg13g2_buf_1 _4689_ (.A(_3938_),
    .X(_3939_));
 sg13g2_buf_2 _4690_ (.A(\collatz.iter[126] ),
    .X(_3940_));
 sg13g2_buf_1 _4691_ (.A(_3940_),
    .X(_3941_));
 sg13g2_nor4_1 _4692_ (.A(net212),
    .B(net211),
    .C(net210),
    .D(net209),
    .Y(_3942_));
 sg13g2_buf_2 _4693_ (.A(\collatz.iter[76] ),
    .X(_3943_));
 sg13g2_buf_1 _4694_ (.A(_3943_),
    .X(_3944_));
 sg13g2_buf_2 _4695_ (.A(\collatz.iter[78] ),
    .X(_3945_));
 sg13g2_buf_1 _4696_ (.A(_3945_),
    .X(_3946_));
 sg13g2_buf_2 _4697_ (.A(\collatz.iter[87] ),
    .X(_3947_));
 sg13g2_buf_1 _4698_ (.A(_3947_),
    .X(_3948_));
 sg13g2_buf_1 _4699_ (.A(\collatz.iter[136] ),
    .X(_3949_));
 sg13g2_buf_1 _4700_ (.A(_3949_),
    .X(_3950_));
 sg13g2_nor4_1 _4701_ (.A(net208),
    .B(net207),
    .C(_3948_),
    .D(_3950_),
    .Y(_3951_));
 sg13g2_nand4_1 _4702_ (.B(_3933_),
    .C(_3942_),
    .A(_3923_),
    .Y(_3952_),
    .D(_3951_));
 sg13g2_nor2_1 _4703_ (.A(_3914_),
    .B(_3952_),
    .Y(_3953_));
 sg13g2_nand4_1 _4704_ (.B(_3829_),
    .C(_3891_),
    .A(_3780_),
    .Y(_3954_),
    .D(_3953_));
 sg13g2_nand3_1 _4705_ (.B(_3379_),
    .C(_3954_),
    .A(_3161_),
    .Y(_3955_));
 sg13g2_inv_1 _4706_ (.Y(\collatz.busy ),
    .A(_3955_));
 sg13g2_buf_1 _4707_ (.A(rst_n),
    .X(_3956_));
 sg13g2_inv_1 _4708_ (.Y(_3957_),
    .A(_3161_));
 sg13g2_buf_1 _4709_ (.A(_3957_),
    .X(_3958_));
 sg13g2_buf_1 _4710_ (.A(uio_in[6]),
    .X(_3959_));
 sg13g2_nand3_1 _4711_ (.B(net109),
    .C(_3959_),
    .A(_3956_),
    .Y(_3960_));
 sg13g2_buf_1 _4712_ (.A(_3960_),
    .X(_3961_));
 sg13g2_buf_1 _4713_ (.A(_3961_),
    .X(_3962_));
 sg13g2_inv_1 _4714_ (.Y(_3963_),
    .A(_3956_));
 sg13g2_buf_1 _4715_ (.A(_3963_),
    .X(_3964_));
 sg13g2_buf_1 _4716_ (.A(_3964_),
    .X(_3965_));
 sg13g2_a21oi_1 _4717_ (.A1(_3955_),
    .A2(net53),
    .Y(_0027_),
    .B1(net108));
 sg13g2_buf_1 _4718_ (.A(_3963_),
    .X(_3966_));
 sg13g2_buf_1 _4719_ (.A(net204),
    .X(_3967_));
 sg13g2_nor2_1 _4720_ (.A(_0016_),
    .B(_0017_),
    .Y(_3968_));
 sg13g2_buf_1 _4721_ (.A(net84),
    .X(_3969_));
 sg13g2_buf_1 _4722_ (.A(_3161_),
    .X(_3970_));
 sg13g2_buf_1 _4723_ (.A(_3970_),
    .X(_3971_));
 sg13g2_nand3_1 _4724_ (.B(net257),
    .C(net106),
    .A(_3969_),
    .Y(_3972_));
 sg13g2_buf_1 _4725_ (.A(ui_in[1]),
    .X(_3973_));
 sg13g2_buf_1 _4726_ (.A(_3973_),
    .X(_3974_));
 sg13g2_buf_1 _4727_ (.A(uio_in[7]),
    .X(_3975_));
 sg13g2_buf_1 _4728_ (.A(uio_in[4]),
    .X(_3976_));
 sg13g2_buf_1 _4729_ (.A(uio_in[3]),
    .X(_3977_));
 sg13g2_buf_2 _4730_ (.A(uio_in[0]),
    .X(_3978_));
 sg13g2_inv_1 _4731_ (.Y(_3979_),
    .A(_3978_));
 sg13g2_buf_1 _4732_ (.A(uio_in[1]),
    .X(_3980_));
 sg13g2_buf_1 _4733_ (.A(uio_in[2]),
    .X(_3981_));
 sg13g2_nor2_1 _4734_ (.A(net329),
    .B(_3981_),
    .Y(_3982_));
 sg13g2_nand2_1 _4735_ (.Y(_3983_),
    .A(_3979_),
    .B(_3982_));
 sg13g2_or3_1 _4736_ (.A(_3976_),
    .B(_3977_),
    .C(_3983_),
    .X(_3984_));
 sg13g2_buf_1 _4737_ (.A(_3984_),
    .X(_3985_));
 sg13g2_inv_1 _4738_ (.Y(_3986_),
    .A(net83));
 sg13g2_nand2_1 _4739_ (.Y(_3987_),
    .A(_3975_),
    .B(_3986_));
 sg13g2_buf_4 _4740_ (.X(_3988_),
    .A(_3987_));
 sg13g2_mux2_1 _4741_ (.A0(net274),
    .A1(_3859_),
    .S(_3988_),
    .X(_3989_));
 sg13g2_nand2_1 _4742_ (.Y(_3990_),
    .A(net109),
    .B(_3989_));
 sg13g2_a21oi_1 _4743_ (.A1(_3972_),
    .A2(_3990_),
    .Y(_3991_),
    .B1(_3968_));
 sg13g2_a21oi_1 _4744_ (.A1(net284),
    .A2(_3968_),
    .Y(_3992_),
    .B1(_3991_));
 sg13g2_nor2_1 _4745_ (.A(net107),
    .B(_3992_),
    .Y(_0018_));
 sg13g2_or2_1 _4746_ (.X(_3993_),
    .B(_3975_),
    .A(_3161_));
 sg13g2_buf_1 _4747_ (.A(_3993_),
    .X(_3994_));
 sg13g2_buf_2 _4748_ (.A(\collatz.path_record_h16[0] ),
    .X(_3995_));
 sg13g2_buf_1 _4749_ (.A(\collatz.path_record_h16[8] ),
    .X(_3996_));
 sg13g2_buf_2 _4750_ (.A(_3978_),
    .X(_3997_));
 sg13g2_buf_4 _4751_ (.X(_3998_),
    .A(uio_in[5]));
 sg13g2_mux4_1 _4752_ (.S0(net273),
    .A0(_3201_),
    .A1(_3271_),
    .A2(_3995_),
    .A3(_3996_),
    .S1(_3998_),
    .X(_3999_));
 sg13g2_buf_1 _4753_ (.A(_3981_),
    .X(_4000_));
 sg13g2_nor3_1 _4754_ (.A(net329),
    .B(_4000_),
    .C(net105),
    .Y(_4001_));
 sg13g2_buf_2 _4755_ (.A(_4001_),
    .X(_4002_));
 sg13g2_a22oi_1 _4756_ (.Y(_4003_),
    .B1(_3999_),
    .B2(_4002_),
    .A2(net105),
    .A1(net5));
 sg13g2_nor2_1 _4757_ (.A(net107),
    .B(_4003_),
    .Y(_0019_));
 sg13g2_mux4_1 _4758_ (.S0(net273),
    .A0(_3191_),
    .A1(\collatz.orbit_len[9] ),
    .A2(\collatz.path_record_h16[1] ),
    .A3(\collatz.path_record_h16[9] ),
    .S1(_3998_),
    .X(_4004_));
 sg13g2_a22oi_1 _4759_ (.Y(_4005_),
    .B1(_4002_),
    .B2(_4004_),
    .A2(net105),
    .A1(net6));
 sg13g2_nor2_1 _4760_ (.A(net107),
    .B(_4005_),
    .Y(_0020_));
 sg13g2_buf_2 _4761_ (.A(\collatz.path_record_h16[2] ),
    .X(_4006_));
 sg13g2_mux4_1 _4762_ (.S0(net273),
    .A0(_3211_),
    .A1(_3310_),
    .A2(_4006_),
    .A3(\collatz.path_record_h16[10] ),
    .S1(_3998_),
    .X(_4007_));
 sg13g2_a22oi_1 _4763_ (.Y(_4008_),
    .B1(_4002_),
    .B2(_4007_),
    .A2(net105),
    .A1(net7));
 sg13g2_nor2_1 _4764_ (.A(net107),
    .B(_4008_),
    .Y(_0021_));
 sg13g2_buf_2 _4765_ (.A(\collatz.path_record_h16[11] ),
    .X(_4009_));
 sg13g2_mux4_1 _4766_ (.S0(net273),
    .A0(\collatz.orbit_len[3] ),
    .A1(_3340_),
    .A2(\collatz.path_record_h16[3] ),
    .A3(_4009_),
    .S1(_3998_),
    .X(_4010_));
 sg13g2_a22oi_1 _4767_ (.Y(_4011_),
    .B1(_4002_),
    .B2(_4010_),
    .A2(_3994_),
    .A1(net8));
 sg13g2_nor2_1 _4768_ (.A(net107),
    .B(_4011_),
    .Y(_0022_));
 sg13g2_buf_2 _4769_ (.A(\collatz.path_record_h16[4] ),
    .X(_4012_));
 sg13g2_mux4_1 _4770_ (.S0(net273),
    .A0(\collatz.orbit_len[4] ),
    .A1(_3349_),
    .A2(_4012_),
    .A3(\collatz.path_record_h16[12] ),
    .S1(_3998_),
    .X(_4013_));
 sg13g2_a22oi_1 _4771_ (.Y(_4014_),
    .B1(_4002_),
    .B2(_4013_),
    .A2(net105),
    .A1(net9));
 sg13g2_nor2_1 _4772_ (.A(net107),
    .B(_4014_),
    .Y(_0023_));
 sg13g2_buf_1 _4773_ (.A(\collatz.path_record_h16[5] ),
    .X(_4015_));
 sg13g2_buf_1 _4774_ (.A(\collatz.path_record_h16[13] ),
    .X(_4016_));
 sg13g2_mux4_1 _4775_ (.S0(net273),
    .A0(\collatz.orbit_len[5] ),
    .A1(\collatz.orbit_len[13] ),
    .A2(_4015_),
    .A3(_4016_),
    .S1(_3998_),
    .X(_4017_));
 sg13g2_a22oi_1 _4776_ (.Y(_4018_),
    .B1(_4002_),
    .B2(_4017_),
    .A2(net105),
    .A1(net10));
 sg13g2_nor2_1 _4777_ (.A(net107),
    .B(_4018_),
    .Y(_0024_));
 sg13g2_buf_2 _4778_ (.A(\collatz.path_record_h16[6] ),
    .X(_4019_));
 sg13g2_buf_2 _4779_ (.A(\collatz.path_record_h16[14] ),
    .X(_4020_));
 sg13g2_mux4_1 _4780_ (.S0(_3997_),
    .A0(_3300_),
    .A1(_3320_),
    .A2(_4019_),
    .A3(_4020_),
    .S1(_3998_),
    .X(_4021_));
 sg13g2_a22oi_1 _4781_ (.Y(_4022_),
    .B1(_4002_),
    .B2(_4021_),
    .A2(net105),
    .A1(net11));
 sg13g2_nor2_1 _4782_ (.A(_3967_),
    .B(_4022_),
    .Y(_0025_));
 sg13g2_buf_1 _4783_ (.A(\collatz.path_record_h16[7] ),
    .X(_4023_));
 sg13g2_mux4_1 _4784_ (.S0(_3997_),
    .A0(_3261_),
    .A1(\collatz.orbit_len[15] ),
    .A2(_4023_),
    .A3(\collatz.path_record_h16[15] ),
    .S1(_3998_),
    .X(_4024_));
 sg13g2_a22oi_1 _4785_ (.Y(_4025_),
    .B1(_4002_),
    .B2(_4024_),
    .A2(net105),
    .A1(net12));
 sg13g2_nor2_1 _4786_ (.A(_3967_),
    .B(_4025_),
    .Y(_0026_));
 sg13g2_buf_1 _4787_ (.A(net203),
    .X(_4026_));
 sg13g2_buf_1 _4788_ (.A(net104),
    .X(_4027_));
 sg13g2_buf_1 _4789_ (.A(net1),
    .X(_4028_));
 sg13g2_buf_1 _4790_ (.A(net283),
    .X(_4029_));
 sg13g2_buf_1 _4791_ (.A(net202),
    .X(_4030_));
 sg13g2_buf_1 _4792_ (.A(net103),
    .X(_4031_));
 sg13g2_buf_1 _4793_ (.A(net81),
    .X(_4032_));
 sg13g2_buf_1 _4794_ (.A(_4032_),
    .X(_4033_));
 sg13g2_buf_1 _4795_ (.A(_4033_),
    .X(_4034_));
 sg13g2_mux2_1 _4796_ (.A0(net328),
    .A1(net42),
    .S(_3988_),
    .X(_4035_));
 sg13g2_inv_1 _4797_ (.Y(_4036_),
    .A(net284));
 sg13g2_buf_1 _4798_ (.A(net67),
    .X(_4037_));
 sg13g2_buf_1 _4799_ (.A(net51),
    .X(_4038_));
 sg13g2_buf_1 _4800_ (.A(net106),
    .X(_4039_));
 sg13g2_o21ai_1 _4801_ (.B1(net80),
    .Y(_4040_),
    .A1(_4036_),
    .A2(_4038_));
 sg13g2_o21ai_1 _4802_ (.B1(_4040_),
    .Y(_4041_),
    .A1(_4027_),
    .A2(_4035_));
 sg13g2_nor2_1 _4803_ (.A(net107),
    .B(_4041_),
    .Y(_0028_));
 sg13g2_buf_1 _4804_ (.A(_3956_),
    .X(_4042_));
 sg13g2_buf_1 _4805_ (.A(net270),
    .X(_4043_));
 sg13g2_buf_1 _4806_ (.A(net203),
    .X(_4044_));
 sg13g2_buf_1 _4807_ (.A(net102),
    .X(_4045_));
 sg13g2_buf_1 _4808_ (.A(_4033_),
    .X(_4046_));
 sg13g2_buf_1 _4809_ (.A(net67),
    .X(_4047_));
 sg13g2_buf_1 _4810_ (.A(_3696_),
    .X(_4048_));
 sg13g2_xnor2_1 _4811_ (.Y(_4049_),
    .A(net242),
    .B(_4048_));
 sg13g2_buf_1 _4812_ (.A(_3775_),
    .X(_4050_));
 sg13g2_nor2b_1 _4813_ (.A(_3814_),
    .B_N(_3788_),
    .Y(_4051_));
 sg13g2_buf_2 _4814_ (.A(_4051_),
    .X(_4052_));
 sg13g2_nor2b_1 _4815_ (.A(_3813_),
    .B_N(net296),
    .Y(_4053_));
 sg13g2_nand3_1 _4816_ (.B(_4052_),
    .C(_4053_),
    .A(net199),
    .Y(_4054_));
 sg13g2_nor2b_1 _4817_ (.A(_3788_),
    .B_N(_3814_),
    .Y(_4055_));
 sg13g2_buf_2 _4818_ (.A(_4055_),
    .X(_4056_));
 sg13g2_nand3_1 _4819_ (.B(_3777_),
    .C(_4056_),
    .A(_3813_),
    .Y(_4057_));
 sg13g2_nand2_1 _4820_ (.Y(_4058_),
    .A(_4054_),
    .B(_4057_));
 sg13g2_nor2_1 _4821_ (.A(_3897_),
    .B(_3899_),
    .Y(_4059_));
 sg13g2_nor2b_1 _4822_ (.A(_3775_),
    .B_N(_3721_),
    .Y(_4060_));
 sg13g2_nand3_1 _4823_ (.B(_4059_),
    .C(_4060_),
    .A(net311),
    .Y(_4061_));
 sg13g2_nor2b_1 _4824_ (.A(\collatz.iter[94] ),
    .B_N(_3775_),
    .Y(_4062_));
 sg13g2_buf_2 _4825_ (.A(_4062_),
    .X(_4063_));
 sg13g2_nor2b_1 _4826_ (.A(net311),
    .B_N(_3899_),
    .Y(_4064_));
 sg13g2_nand3_1 _4827_ (.B(_4063_),
    .C(_4064_),
    .A(_3898_),
    .Y(_4065_));
 sg13g2_nand2_1 _4828_ (.Y(_4066_),
    .A(_4061_),
    .B(_4065_));
 sg13g2_nor2b_1 _4829_ (.A(_3802_),
    .B_N(_3896_),
    .Y(_4067_));
 sg13g2_buf_2 _4830_ (.A(_4067_),
    .X(_4068_));
 sg13g2_nor2b_1 _4831_ (.A(_3786_),
    .B_N(_3897_),
    .Y(_4069_));
 sg13g2_nand3_1 _4832_ (.B(_4068_),
    .C(_4069_),
    .A(net206),
    .Y(_4070_));
 sg13g2_nor2_1 _4833_ (.A(_3947_),
    .B(_3897_),
    .Y(_4071_));
 sg13g2_nor2b_1 _4834_ (.A(_3896_),
    .B_N(_3802_),
    .Y(_4072_));
 sg13g2_buf_2 _4835_ (.A(_4072_),
    .X(_4073_));
 sg13g2_nand3_1 _4836_ (.B(_4071_),
    .C(_4073_),
    .A(_3786_),
    .Y(_4074_));
 sg13g2_nand2_1 _4837_ (.Y(_4075_),
    .A(_4070_),
    .B(_4074_));
 sg13g2_nor2b_1 _4838_ (.A(net276),
    .B_N(_3853_),
    .Y(_4076_));
 sg13g2_buf_2 _4839_ (.A(_4076_),
    .X(_4077_));
 sg13g2_nor2b_1 _4840_ (.A(_3801_),
    .B_N(_3947_),
    .Y(_4078_));
 sg13g2_nand3_1 _4841_ (.B(_4077_),
    .C(_4078_),
    .A(_3852_),
    .Y(_4079_));
 sg13g2_nor2b_1 _4842_ (.A(_3947_),
    .B_N(_3801_),
    .Y(_4080_));
 sg13g2_buf_2 _4843_ (.A(_4080_),
    .X(_4081_));
 sg13g2_nand3_1 _4844_ (.B(_3854_),
    .C(_4081_),
    .A(net276),
    .Y(_4082_));
 sg13g2_nand2_1 _4845_ (.Y(_4083_),
    .A(_4079_),
    .B(_4082_));
 sg13g2_and4_1 _4846_ (.A(_4058_),
    .B(_4066_),
    .C(_4075_),
    .D(_4083_),
    .X(_4084_));
 sg13g2_buf_1 _4847_ (.A(_4084_),
    .X(_4085_));
 sg13g2_inv_1 _4848_ (.Y(_4086_),
    .A(_3852_));
 sg13g2_nor2_1 _4849_ (.A(_3834_),
    .B(_3915_),
    .Y(_4087_));
 sg13g2_nand4_1 _4850_ (.B(_4086_),
    .C(net314),
    .A(net315),
    .Y(_4088_),
    .D(_4087_));
 sg13g2_buf_1 _4851_ (.A(_3852_),
    .X(_4089_));
 sg13g2_inv_1 _4852_ (.Y(_4090_),
    .A(net314));
 sg13g2_nor2b_1 _4853_ (.A(_3700_),
    .B_N(_3834_),
    .Y(_4091_));
 sg13g2_nand4_1 _4854_ (.B(net198),
    .C(_4090_),
    .A(net219),
    .Y(_4092_),
    .D(_4091_));
 sg13g2_nand2_1 _4855_ (.Y(_4093_),
    .A(_4088_),
    .B(_4092_));
 sg13g2_inv_1 _4856_ (.Y(_4094_),
    .A(_3834_));
 sg13g2_and2_1 _4857_ (.A(_3943_),
    .B(_3945_),
    .X(_4095_));
 sg13g2_buf_1 _4858_ (.A(_4095_),
    .X(_4096_));
 sg13g2_buf_1 _4859_ (.A(\collatz.iter[77] ),
    .X(_4097_));
 sg13g2_nor2_1 _4860_ (.A(_3873_),
    .B(net269),
    .Y(_4098_));
 sg13g2_nand3_1 _4861_ (.B(_4096_),
    .C(_4098_),
    .A(_4094_),
    .Y(_4099_));
 sg13g2_nor2_1 _4862_ (.A(_3943_),
    .B(_3945_),
    .Y(_4100_));
 sg13g2_nand4_1 _4863_ (.B(net269),
    .C(_3834_),
    .A(net227),
    .Y(_4101_),
    .D(_4100_));
 sg13g2_nand2_1 _4864_ (.Y(_4102_),
    .A(_4099_),
    .B(_4101_));
 sg13g2_nand2_1 _4865_ (.Y(_4103_),
    .A(_4093_),
    .B(_4102_));
 sg13g2_a21o_1 _4866_ (.A2(net317),
    .A1(net295),
    .B1(net227),
    .X(_4104_));
 sg13g2_a21o_1 _4867_ (.A2(_3874_),
    .A1(net317),
    .B1(net316),
    .X(_4105_));
 sg13g2_buf_1 _4868_ (.A(_3872_),
    .X(_4106_));
 sg13g2_a22oi_1 _4869_ (.Y(_4107_),
    .B1(_4105_),
    .B2(net197),
    .A2(_4104_),
    .A1(net316));
 sg13g2_inv_1 _4870_ (.Y(_4108_),
    .A(_4107_));
 sg13g2_and2_1 _4871_ (.A(_3872_),
    .B(_3873_),
    .X(_4109_));
 sg13g2_buf_1 _4872_ (.A(_4109_),
    .X(_4110_));
 sg13g2_nand3_1 _4873_ (.B(_3695_),
    .C(_4110_),
    .A(net244),
    .Y(_4111_));
 sg13g2_inv_1 _4874_ (.Y(_4112_),
    .A(net295));
 sg13g2_nand4_1 _4875_ (.B(net317),
    .C(net316),
    .A(_4112_),
    .Y(_4113_),
    .D(_3875_));
 sg13g2_nand2_1 _4876_ (.Y(_4114_),
    .A(_4111_),
    .B(_4113_));
 sg13g2_buf_1 _4877_ (.A(_3768_),
    .X(_4115_));
 sg13g2_buf_1 _4878_ (.A(net196),
    .X(_4116_));
 sg13g2_inv_1 _4879_ (.Y(_4117_),
    .A(net299));
 sg13g2_a21o_1 _4880_ (.A2(net294),
    .A1(net306),
    .B1(net320),
    .X(_4118_));
 sg13g2_a21o_1 _4881_ (.A2(net320),
    .A1(net294),
    .B1(net293),
    .X(_4119_));
 sg13g2_buf_2 _4882_ (.A(_3632_),
    .X(_4120_));
 sg13g2_a22oi_1 _4883_ (.Y(_4121_),
    .B1(_4119_),
    .B2(net195),
    .A2(_4118_),
    .A1(net293));
 sg13g2_inv_1 _4884_ (.Y(_4122_),
    .A(_3732_));
 sg13g2_o21ai_1 _4885_ (.B1(_4122_),
    .Y(_4123_),
    .A1(_4117_),
    .A2(_4121_));
 sg13g2_nand2_1 _4886_ (.Y(_4124_),
    .A(net275),
    .B(net252));
 sg13g2_nand2_1 _4887_ (.Y(_4125_),
    .A(net299),
    .B(net196));
 sg13g2_o21ai_1 _4888_ (.B1(_4125_),
    .Y(_4126_),
    .A1(_4124_),
    .A2(_4121_));
 sg13g2_buf_1 _4889_ (.A(net320),
    .X(_4127_));
 sg13g2_a21o_1 _4890_ (.A2(_3732_),
    .A1(net299),
    .B1(net196),
    .X(_4128_));
 sg13g2_and2_1 _4891_ (.A(net213),
    .B(_4128_),
    .X(_4129_));
 sg13g2_a221oi_1 _4892_ (.B2(net194),
    .C1(_4129_),
    .B1(_4126_),
    .A1(net101),
    .Y(_4130_),
    .A2(_4123_));
 sg13g2_nor2_1 _4893_ (.A(_3866_),
    .B(\collatz.iter[71] ),
    .Y(_4131_));
 sg13g2_nor2b_1 _4894_ (.A(_3797_),
    .B_N(\collatz.iter[68] ),
    .Y(_4132_));
 sg13g2_buf_1 _4895_ (.A(_4132_),
    .X(_4133_));
 sg13g2_nand3_1 _4896_ (.B(_4131_),
    .C(_4133_),
    .A(_3847_),
    .Y(_4134_));
 sg13g2_and2_1 _4897_ (.A(_3797_),
    .B(_3866_),
    .X(_4135_));
 sg13g2_buf_1 _4898_ (.A(_4135_),
    .X(_4136_));
 sg13g2_nand3_1 _4899_ (.B(_3848_),
    .C(_4136_),
    .A(net295),
    .Y(_4137_));
 sg13g2_nand2_1 _4900_ (.Y(_4138_),
    .A(_4134_),
    .B(_4137_));
 sg13g2_nor2_1 _4901_ (.A(net298),
    .B(_3781_),
    .Y(_4139_));
 sg13g2_nand4_1 _4902_ (.B(net282),
    .C(_3797_),
    .A(net252),
    .Y(_4140_),
    .D(_4139_));
 sg13g2_buf_1 _4903_ (.A(_4140_),
    .X(_4141_));
 sg13g2_inv_1 _4904_ (.Y(_4142_),
    .A(_3797_));
 sg13g2_nor2b_1 _4905_ (.A(_3864_),
    .B_N(\collatz.iter[64] ),
    .Y(_4143_));
 sg13g2_nand4_1 _4906_ (.B(_4142_),
    .C(_3782_),
    .A(_4122_),
    .Y(_4144_),
    .D(_4143_));
 sg13g2_buf_1 _4907_ (.A(_4144_),
    .X(_4145_));
 sg13g2_nand2_1 _4908_ (.Y(_4146_),
    .A(_4141_),
    .B(_4145_));
 sg13g2_nand2_1 _4909_ (.Y(_4147_),
    .A(_4138_),
    .B(_4146_));
 sg13g2_inv_2 _4910_ (.Y(_4148_),
    .A(net245));
 sg13g2_a21oi_1 _4911_ (.A1(net252),
    .A2(net298),
    .Y(_4149_),
    .B1(net238));
 sg13g2_nor2_1 _4912_ (.A(_4148_),
    .B(_4149_),
    .Y(_4150_));
 sg13g2_a21oi_1 _4913_ (.A1(net298),
    .A2(net238),
    .Y(_4151_),
    .B1(net245));
 sg13g2_nand2b_1 _4914_ (.Y(_4152_),
    .B(net282),
    .A_N(_4151_));
 sg13g2_nand2b_1 _4915_ (.Y(_4153_),
    .B(_4152_),
    .A_N(_4150_));
 sg13g2_inv_1 _4916_ (.Y(_4154_),
    .A(_3866_));
 sg13g2_buf_1 _4917_ (.A(_3847_),
    .X(_4155_));
 sg13g2_a21oi_1 _4918_ (.A1(net287),
    .A2(net295),
    .Y(_4156_),
    .B1(net192));
 sg13g2_a21oi_1 _4919_ (.A1(net238),
    .A2(net287),
    .Y(_4157_),
    .B1(net295));
 sg13g2_nand2b_1 _4920_ (.Y(_4158_),
    .B(net192),
    .A_N(_4157_));
 sg13g2_o21ai_1 _4921_ (.B1(_4158_),
    .Y(_4159_),
    .A1(net193),
    .A2(_4156_));
 sg13g2_a21oi_1 _4922_ (.A1(_4138_),
    .A2(_4153_),
    .Y(_4160_),
    .B1(_4159_));
 sg13g2_o21ai_1 _4923_ (.B1(_4160_),
    .Y(_4161_),
    .A1(_4130_),
    .A2(_4147_));
 sg13g2_and2_1 _4924_ (.A(_4114_),
    .B(_4161_),
    .X(_4162_));
 sg13g2_buf_1 _4925_ (.A(_4162_),
    .X(_4163_));
 sg13g2_o21ai_1 _4926_ (.B1(net302),
    .Y(_4164_),
    .A1(net307),
    .A2(net306));
 sg13g2_buf_1 _4927_ (.A(_3881_),
    .X(_4165_));
 sg13g2_nand3_1 _4928_ (.B(net303),
    .C(net302),
    .A(net191),
    .Y(_4166_));
 sg13g2_nand3_1 _4929_ (.B(net303),
    .C(net306),
    .A(net307),
    .Y(_4167_));
 sg13g2_nand3_1 _4930_ (.B(_4166_),
    .C(_4167_),
    .A(_4164_),
    .Y(_4168_));
 sg13g2_buf_1 _4931_ (.A(net303),
    .X(_4169_));
 sg13g2_buf_1 _4932_ (.A(net302),
    .X(_4170_));
 sg13g2_nand2_1 _4933_ (.Y(_4171_),
    .A(net190),
    .B(net189));
 sg13g2_nand3_1 _4934_ (.B(net254),
    .C(net253),
    .A(net191),
    .Y(_4172_));
 sg13g2_buf_1 _4935_ (.A(net318),
    .X(_4173_));
 sg13g2_a21o_1 _4936_ (.A2(net319),
    .A1(_3894_),
    .B1(_3881_),
    .X(_4174_));
 sg13g2_a21o_1 _4937_ (.A2(_3881_),
    .A1(net319),
    .B1(net318),
    .X(_4175_));
 sg13g2_buf_1 _4938_ (.A(_3880_),
    .X(_4176_));
 sg13g2_a22oi_1 _4939_ (.Y(_4177_),
    .B1(_4175_),
    .B2(_4176_),
    .A2(_4174_),
    .A1(net188));
 sg13g2_buf_1 _4940_ (.A(_4177_),
    .X(_4178_));
 sg13g2_a21oi_1 _4941_ (.A1(_4171_),
    .A2(_4172_),
    .Y(_4179_),
    .B1(_4178_));
 sg13g2_nor2_1 _4942_ (.A(_4168_),
    .B(_4179_),
    .Y(_4180_));
 sg13g2_a21o_1 _4943_ (.A2(_3737_),
    .A1(_3533_),
    .B1(_3892_),
    .X(_4181_));
 sg13g2_a21o_1 _4944_ (.A2(_3892_),
    .A1(_3737_),
    .B1(net304),
    .X(_4182_));
 sg13g2_a22oi_1 _4945_ (.Y(_4183_),
    .B1(_4182_),
    .B2(_3544_),
    .A2(_4181_),
    .A1(net304));
 sg13g2_buf_1 _4946_ (.A(_4183_),
    .X(_4184_));
 sg13g2_inv_1 _4947_ (.Y(_4185_),
    .A(_3892_));
 sg13g2_nand4_1 _4948_ (.B(_4185_),
    .C(net304),
    .A(net305),
    .Y(_4186_),
    .D(_3555_));
 sg13g2_nor2b_1 _4949_ (.A(_3738_),
    .B_N(_3892_),
    .Y(_4187_));
 sg13g2_nor2b_1 _4950_ (.A(net305),
    .B_N(_3544_),
    .Y(_4188_));
 sg13g2_nand3_1 _4951_ (.B(_4187_),
    .C(_4188_),
    .A(_3533_),
    .Y(_4189_));
 sg13g2_and2_1 _4952_ (.A(_4186_),
    .B(_4189_),
    .X(_4190_));
 sg13g2_inv_1 _4953_ (.Y(_4191_),
    .A(_3795_));
 sg13g2_inv_1 _4954_ (.Y(_4192_),
    .A(_3533_));
 sg13g2_nor2b_1 _4955_ (.A(_3929_),
    .B_N(net289),
    .Y(_4193_));
 sg13g2_buf_8 _4956_ (.A(_4193_),
    .X(_4194_));
 sg13g2_nand4_1 _4957_ (.B(_4192_),
    .C(net288),
    .A(_4191_),
    .Y(_4195_),
    .D(_4194_));
 sg13g2_inv_1 _4958_ (.Y(_4196_),
    .A(net288));
 sg13g2_nor2b_1 _4959_ (.A(net289),
    .B_N(_3929_),
    .Y(_4197_));
 sg13g2_nand4_1 _4960_ (.B(_3533_),
    .C(_4196_),
    .A(net239),
    .Y(_4198_),
    .D(_4197_));
 sg13g2_a21o_1 _4961_ (.A2(_3883_),
    .A1(_3764_),
    .B1(net239),
    .X(_4199_));
 sg13g2_a21o_1 _4962_ (.A2(net239),
    .A1(_3883_),
    .B1(_3885_),
    .X(_4200_));
 sg13g2_a22oi_1 _4963_ (.Y(_4201_),
    .B1(_4200_),
    .B2(net215),
    .A2(_4199_),
    .A1(net225));
 sg13g2_a21o_1 _4964_ (.A2(_4198_),
    .A1(_4195_),
    .B1(_4201_),
    .X(_4202_));
 sg13g2_a21o_1 _4965_ (.A2(net289),
    .A1(_3795_),
    .B1(_3533_),
    .X(_4203_));
 sg13g2_a21o_1 _4966_ (.A2(_3533_),
    .A1(net289),
    .B1(net288),
    .X(_4204_));
 sg13g2_a22oi_1 _4967_ (.Y(_4205_),
    .B1(_4204_),
    .B2(net214),
    .A2(_4203_),
    .A1(net288));
 sg13g2_buf_1 _4968_ (.A(_4205_),
    .X(_4206_));
 sg13g2_and2_1 _4969_ (.A(_4184_),
    .B(_4206_),
    .X(_4207_));
 sg13g2_nand3_1 _4970_ (.B(_3705_),
    .C(_3895_),
    .A(net313),
    .Y(_4208_));
 sg13g2_buf_1 _4971_ (.A(_3892_),
    .X(_4209_));
 sg13g2_nor2b_1 _4972_ (.A(net312),
    .B_N(_3894_),
    .Y(_4210_));
 sg13g2_nor2b_1 _4973_ (.A(net313),
    .B_N(_3893_),
    .Y(_4211_));
 sg13g2_nand3_1 _4974_ (.B(_4210_),
    .C(_4211_),
    .A(_4209_),
    .Y(_4212_));
 sg13g2_and2_1 _4975_ (.A(_4208_),
    .B(_4212_),
    .X(_4213_));
 sg13g2_a221oi_1 _4976_ (.B2(_4207_),
    .C1(_4213_),
    .B1(_4202_),
    .A1(_4184_),
    .Y(_4214_),
    .A2(_4190_));
 sg13g2_a22oi_1 _4977_ (.Y(_4215_),
    .B1(_4195_),
    .B2(_4198_),
    .A2(_4189_),
    .A1(_4186_));
 sg13g2_buf_8 _4978_ (.A(_4215_),
    .X(_4216_));
 sg13g2_nor2b_1 _4979_ (.A(_3885_),
    .B_N(_3795_),
    .Y(_0203_));
 sg13g2_buf_2 _4980_ (.A(_0203_),
    .X(_0204_));
 sg13g2_nor2b_1 _4981_ (.A(_3883_),
    .B_N(_3927_),
    .Y(_0205_));
 sg13g2_nand3_1 _4982_ (.B(_0204_),
    .C(_0205_),
    .A(_3764_),
    .Y(_0206_));
 sg13g2_nor2_1 _4983_ (.A(_3764_),
    .B(_3927_),
    .Y(_0207_));
 sg13g2_nand4_1 _4984_ (.B(_4191_),
    .C(_3885_),
    .A(net226),
    .Y(_0208_),
    .D(_0207_));
 sg13g2_a22oi_1 _4985_ (.Y(_0209_),
    .B1(_4208_),
    .B2(_4212_),
    .A2(_0208_),
    .A1(_0206_));
 sg13g2_buf_1 _4986_ (.A(_3894_),
    .X(_0210_));
 sg13g2_a21o_1 _4987_ (.A2(net313),
    .A1(net186),
    .B1(net185),
    .X(_0211_));
 sg13g2_a21o_1 _4988_ (.A2(_3894_),
    .A1(_3703_),
    .B1(net312),
    .X(_0212_));
 sg13g2_buf_1 _4989_ (.A(_3893_),
    .X(_0213_));
 sg13g2_a22oi_1 _4990_ (.Y(_0214_),
    .B1(_0212_),
    .B2(net184),
    .A2(_0211_),
    .A1(_3705_));
 sg13g2_inv_1 _4991_ (.Y(_0215_),
    .A(_0214_));
 sg13g2_a21o_1 _4992_ (.A2(_0209_),
    .A1(_4216_),
    .B1(_0215_),
    .X(_0216_));
 sg13g2_nor2b_1 _4993_ (.A(net318),
    .B_N(_3881_),
    .Y(_0217_));
 sg13g2_nor2b_1 _4994_ (.A(_3690_),
    .B_N(_3880_),
    .Y(_0218_));
 sg13g2_nand3_1 _4995_ (.B(_0217_),
    .C(_0218_),
    .A(net185),
    .Y(_0219_));
 sg13g2_buf_1 _4996_ (.A(net319),
    .X(_0220_));
 sg13g2_nor2b_1 _4997_ (.A(_3894_),
    .B_N(net318),
    .Y(_0221_));
 sg13g2_nand3_1 _4998_ (.B(_3882_),
    .C(_0221_),
    .A(net183),
    .Y(_0222_));
 sg13g2_inv_1 _4999_ (.Y(_0223_),
    .A(net253));
 sg13g2_nor2_1 _5000_ (.A(_3881_),
    .B(net307),
    .Y(_0224_));
 sg13g2_nand4_1 _5001_ (.B(_0223_),
    .C(net189),
    .A(net190),
    .Y(_0225_),
    .D(_0224_));
 sg13g2_nand4_1 _5002_ (.B(_3729_),
    .C(_3731_),
    .A(net191),
    .Y(_0226_),
    .D(_3742_));
 sg13g2_a22oi_1 _5003_ (.Y(_0227_),
    .B1(_0225_),
    .B2(_0226_),
    .A2(_0222_),
    .A1(_0219_));
 sg13g2_o21ai_1 _5004_ (.B1(_0227_),
    .Y(_0228_),
    .A1(_4214_),
    .A2(_0216_));
 sg13g2_nor4_1 _5005_ (.A(_4168_),
    .B(_0215_),
    .C(_4179_),
    .D(_4214_),
    .Y(_0229_));
 sg13g2_a21o_1 _5006_ (.A2(_3676_),
    .A1(net300),
    .B1(_3836_),
    .X(_0230_));
 sg13g2_a21o_1 _5007_ (.A2(_3836_),
    .A1(_3676_),
    .B1(\collatz.iter[14] ),
    .X(_0231_));
 sg13g2_a22oi_1 _5008_ (.Y(_0232_),
    .B1(_0231_),
    .B2(_3755_),
    .A2(_0230_),
    .A1(net278));
 sg13g2_nor2_1 _5009_ (.A(\collatz.iter[17] ),
    .B(_3888_),
    .Y(_0233_));
 sg13g2_a21o_1 _5010_ (.A2(_0232_),
    .A1(_0233_),
    .B1(_3824_),
    .X(_0234_));
 sg13g2_inv_1 _5011_ (.Y(_0235_),
    .A(_3836_));
 sg13g2_buf_1 _5012_ (.A(_3888_),
    .X(_0236_));
 sg13g2_buf_1 _5013_ (.A(net292),
    .X(_0237_));
 sg13g2_buf_1 _5014_ (.A(\collatz.iter[16] ),
    .X(_0238_));
 sg13g2_o21ai_1 _5015_ (.B1(net292),
    .Y(_0239_),
    .A1(net268),
    .A2(_3888_));
 sg13g2_nand2b_1 _5016_ (.Y(_0240_),
    .B(_0239_),
    .A_N(net290));
 sg13g2_o21ai_1 _5017_ (.B1(_0240_),
    .Y(_0241_),
    .A1(net182),
    .A2(net181));
 sg13g2_a221oi_1 _5018_ (.B2(_0235_),
    .C1(_0241_),
    .B1(_0234_),
    .A1(_3824_),
    .Y(_0242_),
    .A2(_0232_));
 sg13g2_nor2b_1 _5019_ (.A(_3924_),
    .B_N(net277),
    .Y(_0243_));
 sg13g2_nor2b_1 _5020_ (.A(_3825_),
    .B_N(_3791_),
    .Y(_0244_));
 sg13g2_nand3_1 _5021_ (.B(_0243_),
    .C(_0244_),
    .A(net308),
    .Y(_0245_));
 sg13g2_nor2_1 _5022_ (.A(net277),
    .B(_3791_),
    .Y(_0246_));
 sg13g2_nor2b_1 _5023_ (.A(net308),
    .B_N(\collatz.iter[26] ),
    .Y(_0247_));
 sg13g2_nand3_1 _5024_ (.B(_0246_),
    .C(_0247_),
    .A(_3924_),
    .Y(_0248_));
 sg13g2_buf_1 _5025_ (.A(\collatz.iter[21] ),
    .X(_0249_));
 sg13g2_nor2_1 _5026_ (.A(_3908_),
    .B(_3759_),
    .Y(_0250_));
 sg13g2_nand4_1 _5027_ (.B(net267),
    .C(net308),
    .A(_3888_),
    .Y(_0251_),
    .D(_0250_));
 sg13g2_inv_1 _5028_ (.Y(_0252_),
    .A(_3726_));
 sg13g2_nand4_1 _5029_ (.B(_0252_),
    .C(_3759_),
    .A(net221),
    .Y(_0253_),
    .D(_3889_));
 sg13g2_a22oi_1 _5030_ (.Y(_0254_),
    .B1(_0251_),
    .B2(_0253_),
    .A2(_0248_),
    .A1(_0245_));
 sg13g2_buf_1 _5031_ (.A(_0254_),
    .X(_0255_));
 sg13g2_inv_1 _5032_ (.Y(_0256_),
    .A(_3791_));
 sg13g2_nor2b_1 _5033_ (.A(_3764_),
    .B_N(_3793_),
    .Y(_0257_));
 sg13g2_nor2b_1 _5034_ (.A(_3762_),
    .B_N(_3826_),
    .Y(_0258_));
 sg13g2_buf_2 _5035_ (.A(_0258_),
    .X(_0259_));
 sg13g2_nand3_1 _5036_ (.B(_0257_),
    .C(_0259_),
    .A(_0256_),
    .Y(_0260_));
 sg13g2_buf_1 _5037_ (.A(_0260_),
    .X(_0261_));
 sg13g2_nor2b_1 _5038_ (.A(_3793_),
    .B_N(_3764_),
    .Y(_0262_));
 sg13g2_buf_2 _5039_ (.A(_0262_),
    .X(_0263_));
 sg13g2_nor2b_1 _5040_ (.A(_3826_),
    .B_N(_3762_),
    .Y(_0264_));
 sg13g2_buf_2 _5041_ (.A(_0264_),
    .X(_0265_));
 sg13g2_nand3_1 _5042_ (.B(_0263_),
    .C(_0265_),
    .A(_3791_),
    .Y(_0266_));
 sg13g2_buf_1 _5043_ (.A(_0266_),
    .X(_0267_));
 sg13g2_nand2_1 _5044_ (.Y(_0268_),
    .A(_0261_),
    .B(_0267_));
 sg13g2_and2_1 _5045_ (.A(_0255_),
    .B(_0268_),
    .X(_0269_));
 sg13g2_nand4_1 _5046_ (.B(net268),
    .C(net292),
    .A(_0235_),
    .Y(_0270_),
    .D(_0233_));
 sg13g2_nand4_1 _5047_ (.B(net290),
    .C(net182),
    .A(net234),
    .Y(_0271_),
    .D(_3824_));
 sg13g2_nor2b_1 _5048_ (.A(net278),
    .B_N(_3836_),
    .Y(_0272_));
 sg13g2_nor2b_1 _5049_ (.A(_3676_),
    .B_N(_3754_),
    .Y(_0273_));
 sg13g2_nand3_1 _5050_ (.B(_0272_),
    .C(_0273_),
    .A(net300),
    .Y(_0274_));
 sg13g2_inv_2 _5051_ (.Y(_0275_),
    .A(_3753_));
 sg13g2_buf_1 _5052_ (.A(_3676_),
    .X(_0276_));
 sg13g2_nor2_2 _5053_ (.A(_3754_),
    .B(_3836_),
    .Y(_0277_));
 sg13g2_nand4_1 _5054_ (.B(net180),
    .C(net278),
    .A(_0275_),
    .Y(_0278_),
    .D(_0277_));
 sg13g2_a22oi_1 _5055_ (.Y(_0279_),
    .B1(_0274_),
    .B2(_0278_),
    .A2(_0271_),
    .A1(_0270_));
 sg13g2_and3_1 _5056_ (.X(_0280_),
    .A(_0255_),
    .B(_0279_),
    .C(_0268_));
 sg13g2_inv_2 _5057_ (.Y(_0281_),
    .A(_3714_));
 sg13g2_nor2_1 _5058_ (.A(_3751_),
    .B(net300),
    .Y(_0282_));
 sg13g2_nand4_1 _5059_ (.B(_3810_),
    .C(_3667_),
    .A(_0281_),
    .Y(_0283_),
    .D(_0282_));
 sg13g2_buf_1 _5060_ (.A(_3714_),
    .X(_0284_));
 sg13g2_inv_1 _5061_ (.Y(_0285_),
    .A(_3810_));
 sg13g2_inv_1 _5062_ (.Y(_0286_),
    .A(_3667_));
 sg13g2_and2_1 _5063_ (.A(_3751_),
    .B(\collatz.iter[11] ),
    .X(_0287_));
 sg13g2_buf_1 _5064_ (.A(_0287_),
    .X(_0288_));
 sg13g2_nand4_1 _5065_ (.B(_0285_),
    .C(_0286_),
    .A(net179),
    .Y(_0289_),
    .D(_0288_));
 sg13g2_nor2_1 _5066_ (.A(_3757_),
    .B(_3713_),
    .Y(_0290_));
 sg13g2_nand4_1 _5067_ (.B(_0281_),
    .C(_3809_),
    .A(net256),
    .Y(_0291_),
    .D(_0290_));
 sg13g2_buf_1 _5068_ (.A(_3713_),
    .X(_0292_));
 sg13g2_nor2_1 _5069_ (.A(_3710_),
    .B(_3808_),
    .Y(_0293_));
 sg13g2_nand4_1 _5070_ (.B(net178),
    .C(net179),
    .A(net249),
    .Y(_0294_),
    .D(_0293_));
 sg13g2_a21o_1 _5071_ (.A2(_3757_),
    .A1(\collatz.iter[0] ),
    .B1(_3708_),
    .X(_0295_));
 sg13g2_or2_1 _5072_ (.X(_0296_),
    .B(_3757_),
    .A(net283));
 sg13g2_a22oi_1 _5073_ (.Y(_0297_),
    .B1(_0296_),
    .B2(net257),
    .A2(_0295_),
    .A1(net284));
 sg13g2_a221oi_1 _5074_ (.B2(_0294_),
    .C1(_0297_),
    .B1(_0291_),
    .A1(_0283_),
    .Y(_0298_),
    .A2(_0289_));
 sg13g2_a21o_1 _5075_ (.A2(_3710_),
    .A1(_3757_),
    .B1(net179),
    .X(_0299_));
 sg13g2_a21o_1 _5076_ (.A2(_3714_),
    .A1(_3710_),
    .B1(_3808_),
    .X(_0300_));
 sg13g2_a22oi_1 _5077_ (.Y(_0301_),
    .B1(_0300_),
    .B2(net178),
    .A2(_0299_),
    .A1(_3809_));
 sg13g2_a21o_1 _5078_ (.A2(_0289_),
    .A1(_0283_),
    .B1(_0301_),
    .X(_0302_));
 sg13g2_buf_1 _5079_ (.A(_3667_),
    .X(_0303_));
 sg13g2_o21ai_1 _5080_ (.B1(_0275_),
    .Y(_0304_),
    .A1(_0281_),
    .A2(_0285_));
 sg13g2_o21ai_1 _5081_ (.B1(_0286_),
    .Y(_0305_),
    .A1(_0285_),
    .A2(_0275_));
 sg13g2_a22oi_1 _5082_ (.Y(_0306_),
    .B1(_0305_),
    .B2(net251),
    .A2(_0304_),
    .A1(net177));
 sg13g2_nand3b_1 _5083_ (.B(_0302_),
    .C(_0306_),
    .Y(_0307_),
    .A_N(_0298_));
 sg13g2_buf_2 _5084_ (.A(_0307_),
    .X(_0308_));
 sg13g2_a21o_1 _5085_ (.A2(net221),
    .A1(net182),
    .B1(net308),
    .X(_0309_));
 sg13g2_a21o_1 _5086_ (.A2(net308),
    .A1(net221),
    .B1(net248),
    .X(_0310_));
 sg13g2_a22oi_1 _5087_ (.Y(_0311_),
    .B1(_0310_),
    .B2(net267),
    .A2(_0309_),
    .A1(net248));
 sg13g2_a221oi_1 _5088_ (.B2(_0267_),
    .C1(_0311_),
    .B1(_0261_),
    .A1(_0245_),
    .Y(_0312_),
    .A2(_0248_));
 sg13g2_buf_1 _5089_ (.A(net291),
    .X(_0313_));
 sg13g2_a21o_1 _5090_ (.A2(_3924_),
    .A1(net308),
    .B1(_3791_),
    .X(_0314_));
 sg13g2_a21o_1 _5091_ (.A2(_3791_),
    .A1(net216),
    .B1(_3825_),
    .X(_0315_));
 sg13g2_a22oi_1 _5092_ (.Y(_0316_),
    .B1(_0315_),
    .B2(_3911_),
    .A2(_0314_),
    .A1(net176));
 sg13g2_a21o_1 _5093_ (.A2(_0267_),
    .A1(_0261_),
    .B1(_0316_),
    .X(_0317_));
 sg13g2_buf_1 _5094_ (.A(_3826_),
    .X(_0318_));
 sg13g2_a21o_1 _5095_ (.A2(net175),
    .A1(net241),
    .B1(net246),
    .X(_0319_));
 sg13g2_a21o_1 _5096_ (.A2(net246),
    .A1(net175),
    .B1(_3793_),
    .X(_0320_));
 sg13g2_a22oi_1 _5097_ (.Y(_0321_),
    .B1(_0320_),
    .B2(net247),
    .A2(_0319_),
    .A1(net240));
 sg13g2_nand3b_1 _5098_ (.B(_0317_),
    .C(_0321_),
    .Y(_0322_),
    .A_N(_0312_));
 sg13g2_a221oi_1 _5099_ (.B2(_0308_),
    .C1(_0322_),
    .B1(_0280_),
    .A1(_0242_),
    .Y(_0323_),
    .A2(_0269_));
 sg13g2_buf_2 _5100_ (.A(_0323_),
    .X(_0324_));
 sg13g2_and2_1 _5101_ (.A(_4111_),
    .B(_4113_),
    .X(_0325_));
 sg13g2_or4_1 _5102_ (.A(net194),
    .B(net275),
    .C(net252),
    .D(_4125_),
    .X(_0326_));
 sg13g2_buf_1 _5103_ (.A(net299),
    .X(_0327_));
 sg13g2_nor2_1 _5104_ (.A(net174),
    .B(net196),
    .Y(_0328_));
 sg13g2_nand4_1 _5105_ (.B(net213),
    .C(net116),
    .A(_4127_),
    .Y(_0329_),
    .D(_0328_));
 sg13g2_nor2b_1 _5106_ (.A(net306),
    .B_N(\collatz.iter[56] ),
    .Y(_0330_));
 sg13g2_and2_1 _5107_ (.A(net293),
    .B(_0330_),
    .X(_0331_));
 sg13g2_nand3b_1 _5108_ (.B(net320),
    .C(_3632_),
    .Y(_0332_),
    .A_N(net294));
 sg13g2_nor2_1 _5109_ (.A(net293),
    .B(_0332_),
    .Y(_0333_));
 sg13g2_a22oi_1 _5110_ (.Y(_0334_),
    .B1(_0333_),
    .B2(net253),
    .A2(_0331_),
    .A1(_3650_));
 sg13g2_buf_1 _5111_ (.A(_0334_),
    .X(_0335_));
 sg13g2_a21o_1 _5112_ (.A2(_0329_),
    .A1(_0326_),
    .B1(_0335_),
    .X(_0336_));
 sg13g2_or3_1 _5113_ (.A(_0325_),
    .B(_4147_),
    .C(_0336_),
    .X(_0337_));
 sg13g2_a221oi_1 _5114_ (.B2(_0324_),
    .C1(_0337_),
    .B1(_0229_),
    .A1(_4180_),
    .Y(_0338_),
    .A2(_0228_));
 sg13g2_nor3_1 _5115_ (.A(_4108_),
    .B(_4163_),
    .C(_0338_),
    .Y(_0339_));
 sg13g2_inv_1 _5116_ (.Y(_0340_),
    .A(net207));
 sg13g2_a21oi_1 _5117_ (.A1(net227),
    .A2(_3943_),
    .Y(_0341_),
    .B1(_3834_));
 sg13g2_and2_1 _5118_ (.A(_3943_),
    .B(_3834_),
    .X(_0342_));
 sg13g2_o21ai_1 _5119_ (.B1(net269),
    .Y(_0343_),
    .A1(net207),
    .A2(_0342_));
 sg13g2_o21ai_1 _5120_ (.B1(_0343_),
    .Y(_0344_),
    .A1(_0340_),
    .A2(_0341_));
 sg13g2_buf_1 _5121_ (.A(_3834_),
    .X(_0345_));
 sg13g2_a21oi_1 _5122_ (.A1(net173),
    .A2(net315),
    .Y(_0346_),
    .B1(net198));
 sg13g2_buf_1 _5123_ (.A(net314),
    .X(_0347_));
 sg13g2_and2_1 _5124_ (.A(net315),
    .B(_3852_),
    .X(_0348_));
 sg13g2_o21ai_1 _5125_ (.B1(net219),
    .Y(_0349_),
    .A1(_0347_),
    .A2(_0348_));
 sg13g2_o21ai_1 _5126_ (.B1(_0349_),
    .Y(_0350_),
    .A1(_4090_),
    .A2(_0346_));
 sg13g2_a21oi_1 _5127_ (.A1(_4093_),
    .A2(_0344_),
    .Y(_0351_),
    .B1(_0350_));
 sg13g2_o21ai_1 _5128_ (.B1(_0351_),
    .Y(_0352_),
    .A1(_4103_),
    .A2(_0339_));
 sg13g2_a21o_1 _5129_ (.A2(net276),
    .A1(_3852_),
    .B1(_3947_),
    .X(_0353_));
 sg13g2_a21o_1 _5130_ (.A2(_3947_),
    .A1(net276),
    .B1(_3801_),
    .X(_0354_));
 sg13g2_buf_1 _5131_ (.A(_3853_),
    .X(_0355_));
 sg13g2_a22oi_1 _5132_ (.Y(_0356_),
    .B1(_0354_),
    .B2(net171),
    .A2(_0353_),
    .A1(_3801_));
 sg13g2_a21o_1 _5133_ (.A2(_4074_),
    .A1(_4070_),
    .B1(_0356_),
    .X(_0357_));
 sg13g2_a21o_1 _5134_ (.A2(net311),
    .A1(_3897_),
    .B1(_3775_),
    .X(_0358_));
 sg13g2_a21o_1 _5135_ (.A2(_3775_),
    .A1(net311),
    .B1(net310),
    .X(_0359_));
 sg13g2_a22oi_1 _5136_ (.Y(_0360_),
    .B1(_0359_),
    .B2(_3899_),
    .A2(_0358_),
    .A1(net310));
 sg13g2_a21oi_1 _5137_ (.A1(_3947_),
    .A2(_3802_),
    .Y(_0361_),
    .B1(net224));
 sg13g2_nand2b_1 _5138_ (.Y(_0362_),
    .B(_3786_),
    .A_N(_0361_));
 sg13g2_and2_1 _5139_ (.A(_3802_),
    .B(_3897_),
    .X(_0363_));
 sg13g2_buf_1 _5140_ (.A(_3896_),
    .X(_0364_));
 sg13g2_o21ai_1 _5141_ (.B1(_0364_),
    .Y(_0365_),
    .A1(_3786_),
    .A2(_0363_));
 sg13g2_and3_1 _5142_ (.X(_0366_),
    .A(_0360_),
    .B(_0362_),
    .C(_0365_));
 sg13g2_and3_1 _5143_ (.X(_0367_),
    .A(_0360_),
    .B(_4061_),
    .C(_4065_));
 sg13g2_a221oi_1 _5144_ (.B2(_0366_),
    .C1(_0367_),
    .B1(_0357_),
    .A1(_4054_),
    .Y(_0368_),
    .A2(_4057_));
 sg13g2_inv_1 _5145_ (.Y(_0369_),
    .A(net235));
 sg13g2_buf_1 _5146_ (.A(_3813_),
    .X(_0370_));
 sg13g2_a21oi_1 _5147_ (.A1(net199),
    .A2(_0370_),
    .Y(_0371_),
    .B1(net242));
 sg13g2_nor2_1 _5148_ (.A(_0369_),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_a21oi_1 _5149_ (.A1(_0370_),
    .A2(net242),
    .Y(_0373_),
    .B1(net235));
 sg13g2_buf_1 _5150_ (.A(net296),
    .X(_0374_));
 sg13g2_nand2b_1 _5151_ (.Y(_0375_),
    .B(_0374_),
    .A_N(_0373_));
 sg13g2_nor2b_1 _5152_ (.A(_0372_),
    .B_N(_0375_),
    .Y(_0376_));
 sg13g2_nand2b_1 _5153_ (.Y(_0377_),
    .B(_0376_),
    .A_N(_0368_));
 sg13g2_a21oi_1 _5154_ (.A1(_4085_),
    .A2(_0352_),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_xnor2_1 _5155_ (.Y(_0379_),
    .A(_4049_),
    .B(_0378_));
 sg13g2_nand2_1 _5156_ (.Y(_0380_),
    .A(net50),
    .B(_0379_));
 sg13g2_o21ai_1 _5157_ (.B1(_0380_),
    .Y(_0381_),
    .A1(net40),
    .A2(_3921_));
 sg13g2_buf_1 _5158_ (.A(ui_in[4]),
    .X(_0382_));
 sg13g2_inv_1 _5159_ (.Y(_0383_),
    .A(net329));
 sg13g2_nor3_2 _5160_ (.A(_3978_),
    .B(net329),
    .C(_3981_),
    .Y(_0384_));
 sg13g2_nand2b_1 _5161_ (.Y(_0385_),
    .B(_3977_),
    .A_N(_3976_));
 sg13g2_nand3b_1 _5162_ (.B(_0384_),
    .C(_3976_),
    .Y(_0386_),
    .A_N(_3977_));
 sg13g2_o21ai_1 _5163_ (.B1(_0386_),
    .Y(_0387_),
    .A1(_0384_),
    .A2(_0385_));
 sg13g2_and2_1 _5164_ (.A(_3975_),
    .B(_0387_),
    .X(_0388_));
 sg13g2_buf_1 _5165_ (.A(_0388_),
    .X(_0389_));
 sg13g2_and4_1 _5166_ (.A(_3979_),
    .B(_0383_),
    .C(net272),
    .D(net66),
    .X(_0390_));
 sg13g2_buf_1 _5167_ (.A(_0390_),
    .X(_0391_));
 sg13g2_buf_1 _5168_ (.A(_0391_),
    .X(_0392_));
 sg13g2_nand2_1 _5169_ (.Y(_0393_),
    .A(_3956_),
    .B(_3161_));
 sg13g2_nand2b_1 _5170_ (.Y(_0394_),
    .B(_3955_),
    .A_N(_0393_));
 sg13g2_buf_1 _5171_ (.A(_0394_),
    .X(_0395_));
 sg13g2_buf_1 _5172_ (.A(_0395_),
    .X(_0396_));
 sg13g2_inv_2 _5173_ (.Y(_0397_),
    .A(_3696_));
 sg13g2_nor2_1 _5174_ (.A(_0397_),
    .B(_0391_),
    .Y(_0398_));
 sg13g2_buf_1 _5175_ (.A(net203),
    .X(_0399_));
 sg13g2_buf_1 _5176_ (.A(_0399_),
    .X(_0400_));
 sg13g2_a221oi_1 _5177_ (.B2(_0398_),
    .C1(_0400_),
    .B1(net19),
    .A1(net327),
    .Y(_0401_),
    .A2(_0392_));
 sg13g2_a21oi_1 _5178_ (.A1(_4045_),
    .A2(_0381_),
    .Y(_0402_),
    .B1(_0401_));
 sg13g2_and2_1 _5179_ (.A(_4043_),
    .B(_0402_),
    .X(_0029_));
 sg13g2_buf_1 _5180_ (.A(_3964_),
    .X(_0403_));
 sg13g2_buf_1 _5181_ (.A(net109),
    .X(_0404_));
 sg13g2_buf_1 _5182_ (.A(net77),
    .X(_0405_));
 sg13g2_buf_1 _5183_ (.A(net52),
    .X(_0406_));
 sg13g2_nor2b_1 _5184_ (.A(_3920_),
    .B_N(_3696_),
    .Y(_0407_));
 sg13g2_nor2b_1 _5185_ (.A(_3696_),
    .B_N(_3920_),
    .Y(_0408_));
 sg13g2_nor2_1 _5186_ (.A(_0407_),
    .B(_0408_),
    .Y(_0409_));
 sg13g2_inv_1 _5187_ (.Y(_0410_),
    .A(net315));
 sg13g2_nand2_1 _5188_ (.Y(_0411_),
    .A(net314),
    .B(net276));
 sg13g2_or4_1 _5189_ (.A(net219),
    .B(_0410_),
    .C(_3852_),
    .D(_0411_),
    .X(_0412_));
 sg13g2_nor2_1 _5190_ (.A(net314),
    .B(_3918_),
    .Y(_0413_));
 sg13g2_nand4_1 _5191_ (.B(_0410_),
    .C(net198),
    .A(net219),
    .Y(_0414_),
    .D(_0413_));
 sg13g2_and2_1 _5192_ (.A(_3945_),
    .B(net315),
    .X(_0415_));
 sg13g2_buf_1 _5193_ (.A(_0415_),
    .X(_0416_));
 sg13g2_nand3_1 _5194_ (.B(_3835_),
    .C(_0416_),
    .A(net208),
    .Y(_0417_));
 sg13g2_buf_1 _5195_ (.A(net269),
    .X(_0418_));
 sg13g2_nand3_1 _5196_ (.B(_4100_),
    .C(_4091_),
    .A(net167),
    .Y(_0419_));
 sg13g2_a22oi_1 _5197_ (.Y(_0420_),
    .B1(_0417_),
    .B2(_0419_),
    .A2(_0414_),
    .A1(_0412_));
 sg13g2_nand3_1 _5198_ (.B(_4133_),
    .C(_4143_),
    .A(net245),
    .Y(_0421_));
 sg13g2_inv_1 _5199_ (.Y(_0422_),
    .A(net298));
 sg13g2_nor2_1 _5200_ (.A(_3781_),
    .B(net287),
    .Y(_0423_));
 sg13g2_nand4_1 _5201_ (.B(_0422_),
    .C(net238),
    .A(net282),
    .Y(_0424_),
    .D(_0423_));
 sg13g2_nand2_1 _5202_ (.Y(_0425_),
    .A(_0421_),
    .B(_0424_));
 sg13g2_buf_1 _5203_ (.A(net298),
    .X(_0426_));
 sg13g2_o21ai_1 _5204_ (.B1(net116),
    .Y(_0427_),
    .A1(_4116_),
    .A2(net166));
 sg13g2_a22oi_1 _5205_ (.Y(_0428_),
    .B1(net196),
    .B2(net166),
    .A2(net252),
    .A1(net174));
 sg13g2_nand2b_1 _5206_ (.Y(_0429_),
    .B(net213),
    .A_N(_0428_));
 sg13g2_nand2_1 _5207_ (.Y(_0430_),
    .A(_0427_),
    .B(_0429_));
 sg13g2_a22oi_1 _5208_ (.Y(_0431_),
    .B1(net248),
    .B2(net216),
    .A2(net255),
    .A1(net221));
 sg13g2_buf_1 _5209_ (.A(_0249_),
    .X(_0432_));
 sg13g2_nand2b_1 _5210_ (.Y(_0433_),
    .B(net165),
    .A_N(_0431_));
 sg13g2_and2_1 _5211_ (.A(net277),
    .B(_3791_),
    .X(_0434_));
 sg13g2_buf_1 _5212_ (.A(_0434_),
    .X(_0435_));
 sg13g2_o21ai_1 _5213_ (.B1(net255),
    .Y(_0436_),
    .A1(net248),
    .A2(_3925_));
 sg13g2_nor2b_1 _5214_ (.A(_0435_),
    .B_N(_0436_),
    .Y(_0437_));
 sg13g2_and2_1 _5215_ (.A(net291),
    .B(_3826_),
    .X(_0438_));
 sg13g2_buf_1 _5216_ (.A(_0438_),
    .X(_0439_));
 sg13g2_o21ai_1 _5217_ (.B1(net110),
    .Y(_0440_),
    .A1(_0435_),
    .A2(_0439_));
 sg13g2_a21o_1 _5218_ (.A2(_0437_),
    .A1(_0433_),
    .B1(_0440_),
    .X(_0441_));
 sg13g2_o21ai_1 _5219_ (.B1(net241),
    .Y(_0442_),
    .A1(net291),
    .A2(_3826_));
 sg13g2_inv_1 _5220_ (.Y(_0443_),
    .A(net165));
 sg13g2_o21ai_1 _5221_ (.B1(_0436_),
    .Y(_0444_),
    .A1(_0443_),
    .A2(_0431_));
 sg13g2_a22oi_1 _5222_ (.Y(_0445_),
    .B1(_0444_),
    .B2(_0435_),
    .A2(_0439_),
    .A1(_3912_));
 sg13g2_and3_1 _5223_ (.X(_0446_),
    .A(_0441_),
    .B(_0442_),
    .C(_0445_));
 sg13g2_buf_1 _5224_ (.A(_0446_),
    .X(_0447_));
 sg13g2_buf_1 _5225_ (.A(net268),
    .X(_0448_));
 sg13g2_nand4_1 _5226_ (.B(net181),
    .C(net221),
    .A(net164),
    .Y(_0449_),
    .D(_0233_));
 sg13g2_inv_1 _5227_ (.Y(_0450_),
    .A(net268));
 sg13g2_nor2_1 _5228_ (.A(net292),
    .B(_3908_),
    .Y(_0451_));
 sg13g2_nand4_1 _5229_ (.B(_0450_),
    .C(net182),
    .A(net233),
    .Y(_0452_),
    .D(_0451_));
 sg13g2_nand2_1 _5230_ (.Y(_0453_),
    .A(_0449_),
    .B(_0452_));
 sg13g2_inv_1 _5231_ (.Y(_0454_),
    .A(_0276_));
 sg13g2_a22oi_1 _5232_ (.Y(_0455_),
    .B1(_3667_),
    .B2(_3676_),
    .A2(net300),
    .A1(net236));
 sg13g2_nand2b_1 _5233_ (.Y(_0456_),
    .B(_3752_),
    .A_N(_0455_));
 sg13g2_nor2_1 _5234_ (.A(net278),
    .B(net268),
    .Y(_0457_));
 sg13g2_o21ai_1 _5235_ (.B1(net300),
    .Y(_0458_),
    .A1(_3667_),
    .A2(_3676_));
 sg13g2_and3_1 _5236_ (.X(_0459_),
    .A(_0454_),
    .B(_0457_),
    .C(_0458_));
 sg13g2_a22oi_1 _5237_ (.Y(_0460_),
    .B1(_0456_),
    .B2(_0459_),
    .A2(_0277_),
    .A1(_0454_));
 sg13g2_inv_1 _5238_ (.Y(_0461_),
    .A(_3754_));
 sg13g2_and2_1 _5239_ (.A(_0277_),
    .B(_0458_),
    .X(_0462_));
 sg13g2_a21oi_1 _5240_ (.A1(net222),
    .A2(net164),
    .Y(_0463_),
    .B1(net234));
 sg13g2_a221oi_1 _5241_ (.B2(_0462_),
    .C1(_0463_),
    .B1(_0456_),
    .A1(_0461_),
    .Y(_0464_),
    .A2(_0457_));
 sg13g2_nand3_1 _5242_ (.B(_0460_),
    .C(_0464_),
    .A(_0453_),
    .Y(_0465_));
 sg13g2_and2_1 _5243_ (.A(net283),
    .B(net249),
    .X(_0466_));
 sg13g2_and2_1 _5244_ (.A(_3708_),
    .B(_3710_),
    .X(_0467_));
 sg13g2_buf_2 _5245_ (.A(_0467_),
    .X(_0468_));
 sg13g2_o21ai_1 _5246_ (.B1(net284),
    .Y(_0469_),
    .A1(_0466_),
    .A2(_0468_));
 sg13g2_a22oi_1 _5247_ (.Y(_0470_),
    .B1(_0468_),
    .B2(net283),
    .A2(_3712_),
    .A1(net249));
 sg13g2_or2_1 _5248_ (.X(_0471_),
    .B(_3808_),
    .A(_3710_));
 sg13g2_o21ai_1 _5249_ (.B1(_3716_),
    .Y(_0472_),
    .A1(net236),
    .A2(_0471_));
 sg13g2_nand3_1 _5250_ (.B(_0470_),
    .C(_0472_),
    .A(_0469_),
    .Y(_0473_));
 sg13g2_buf_1 _5251_ (.A(_0473_),
    .X(_0474_));
 sg13g2_nand4_1 _5252_ (.B(net177),
    .C(net180),
    .A(net236),
    .Y(_0475_),
    .D(_0282_));
 sg13g2_nand3_1 _5253_ (.B(_3684_),
    .C(_0288_),
    .A(_0285_),
    .Y(_0476_));
 sg13g2_nand2_1 _5254_ (.Y(_0477_),
    .A(_3808_),
    .B(_3810_));
 sg13g2_or2_1 _5255_ (.X(_0478_),
    .B(net179),
    .A(_3711_));
 sg13g2_a21oi_1 _5256_ (.A1(_3812_),
    .A2(_0478_),
    .Y(_0479_),
    .B1(net178));
 sg13g2_a221oi_1 _5257_ (.B2(_0281_),
    .C1(_0479_),
    .B1(_0477_),
    .A1(_0475_),
    .Y(_0480_),
    .A2(_0476_));
 sg13g2_nand3_1 _5258_ (.B(net222),
    .C(_0277_),
    .A(net180),
    .Y(_0481_));
 sg13g2_nand3_1 _5259_ (.B(_0272_),
    .C(_0273_),
    .A(_0450_),
    .Y(_0482_));
 sg13g2_o21ai_1 _5260_ (.B1(_0482_),
    .Y(_0483_),
    .A1(_0450_),
    .A2(_0481_));
 sg13g2_nand4_1 _5261_ (.B(_0474_),
    .C(_0480_),
    .A(_0453_),
    .Y(_0484_),
    .D(_0483_));
 sg13g2_inv_1 _5262_ (.Y(_0485_),
    .A(_3927_));
 sg13g2_a22oi_1 _5263_ (.Y(_0486_),
    .B1(net225),
    .B2(net289),
    .A2(net239),
    .A1(net226));
 sg13g2_o21ai_1 _5264_ (.B1(net239),
    .Y(_0487_),
    .A1(net225),
    .A2(net232));
 sg13g2_o21ai_1 _5265_ (.B1(_0487_),
    .Y(_0488_),
    .A1(_0485_),
    .A2(_0486_));
 sg13g2_buf_1 _5266_ (.A(_0488_),
    .X(_0489_));
 sg13g2_nor2b_1 _5267_ (.A(net215),
    .B_N(_3883_),
    .Y(_0490_));
 sg13g2_nor2b_1 _5268_ (.A(_3795_),
    .B_N(_3885_),
    .Y(_0491_));
 sg13g2_nand3_1 _5269_ (.B(_0490_),
    .C(_0491_),
    .A(_3841_),
    .Y(_0492_));
 sg13g2_nand3b_1 _5270_ (.B(_0204_),
    .C(_0205_),
    .Y(_0493_),
    .A_N(net289));
 sg13g2_o21ai_1 _5271_ (.B1(net246),
    .Y(_0494_),
    .A1(_3794_),
    .A2(net226));
 sg13g2_and2_1 _5272_ (.A(_3793_),
    .B(_3883_),
    .X(_0495_));
 sg13g2_buf_2 _5273_ (.A(_0495_),
    .X(_0496_));
 sg13g2_and2_1 _5274_ (.A(net247),
    .B(_3764_),
    .X(_0497_));
 sg13g2_a22oi_1 _5275_ (.Y(_0498_),
    .B1(_0497_),
    .B2(net175),
    .A2(_0496_),
    .A1(_3763_));
 sg13g2_a22oi_1 _5276_ (.Y(_0499_),
    .B1(_0494_),
    .B2(_0498_),
    .A2(_0493_),
    .A1(_0492_));
 sg13g2_inv_1 _5277_ (.Y(_0500_),
    .A(_3888_));
 sg13g2_a22oi_1 _5278_ (.Y(_0501_),
    .B1(net181),
    .B2(net221),
    .A2(net182),
    .A1(net268));
 sg13g2_nand2b_1 _5279_ (.Y(_0502_),
    .B(net233),
    .A_N(_0501_));
 sg13g2_o21ai_1 _5280_ (.B1(_0502_),
    .Y(_0503_),
    .A1(_0500_),
    .A2(_0451_));
 sg13g2_nor3_1 _5281_ (.A(_0489_),
    .B(_0499_),
    .C(_0503_),
    .Y(_0504_));
 sg13g2_nand4_1 _5282_ (.B(_0465_),
    .C(_0484_),
    .A(_0447_),
    .Y(_0505_),
    .D(_0504_));
 sg13g2_nor2_1 _5283_ (.A(_0489_),
    .B(_0499_),
    .Y(_0506_));
 sg13g2_nand3b_1 _5284_ (.B(_0263_),
    .C(_0265_),
    .Y(_0507_),
    .A_N(net226));
 sg13g2_nand3b_1 _5285_ (.B(_0259_),
    .C(_0496_),
    .Y(_0508_),
    .A_N(net246));
 sg13g2_and2_1 _5286_ (.A(_0507_),
    .B(_0508_),
    .X(_0509_));
 sg13g2_a21o_1 _5287_ (.A2(_0493_),
    .A1(_0492_),
    .B1(_0509_),
    .X(_0510_));
 sg13g2_nand2_1 _5288_ (.Y(_0511_),
    .A(_0492_),
    .B(_0493_));
 sg13g2_nand2_1 _5289_ (.Y(_0512_),
    .A(_0494_),
    .B(_0498_));
 sg13g2_nor2_1 _5290_ (.A(net267),
    .B(net308),
    .Y(_0513_));
 sg13g2_nand4_1 _5291_ (.B(net248),
    .C(net216),
    .A(net112),
    .Y(_0514_),
    .D(_0513_));
 sg13g2_nand2_1 _5292_ (.Y(_0515_),
    .A(net267),
    .B(net308));
 sg13g2_or2_1 _5293_ (.X(_0516_),
    .B(_3759_),
    .A(_3908_));
 sg13g2_buf_1 _5294_ (.A(_0516_),
    .X(_0517_));
 sg13g2_or3_1 _5295_ (.A(net216),
    .B(_0515_),
    .C(_0517_),
    .X(_0518_));
 sg13g2_nand2_1 _5296_ (.Y(_0519_),
    .A(_0514_),
    .B(_0518_));
 sg13g2_nand3_1 _5297_ (.B(_0246_),
    .C(_0439_),
    .A(net216),
    .Y(_0520_));
 sg13g2_nand3_1 _5298_ (.B(_3827_),
    .C(_0243_),
    .A(net241),
    .Y(_0521_));
 sg13g2_nand2_1 _5299_ (.Y(_0522_),
    .A(_0520_),
    .B(_0521_));
 sg13g2_a221oi_1 _5300_ (.B2(_0522_),
    .C1(_0489_),
    .B1(_0519_),
    .A1(_0511_),
    .Y(_0523_),
    .A2(_0512_));
 sg13g2_a22oi_1 _5301_ (.Y(_0524_),
    .B1(_0447_),
    .B2(_0523_),
    .A2(_0510_),
    .A1(_0506_));
 sg13g2_nand2_2 _5302_ (.Y(_0525_),
    .A(_0505_),
    .B(_0524_));
 sg13g2_nor2_1 _5303_ (.A(\collatz.iter[58] ),
    .B(net299),
    .Y(_0526_));
 sg13g2_nand2b_1 _5304_ (.Y(_0527_),
    .B(_0526_),
    .A_N(_0332_));
 sg13g2_buf_1 _5305_ (.A(net293),
    .X(_0528_));
 sg13g2_nand4_1 _5306_ (.B(net163),
    .C(net174),
    .A(_3820_),
    .Y(_0529_),
    .D(_3650_));
 sg13g2_buf_1 _5307_ (.A(net294),
    .X(_0530_));
 sg13g2_nor2_1 _5308_ (.A(net307),
    .B(net306),
    .Y(_0531_));
 sg13g2_nand4_1 _5309_ (.B(_3741_),
    .C(net162),
    .A(net303),
    .Y(_0532_),
    .D(_0531_));
 sg13g2_inv_1 _5310_ (.Y(_0533_),
    .A(net294));
 sg13g2_nand4_1 _5311_ (.B(net306),
    .C(_0533_),
    .A(net254),
    .Y(_0534_),
    .D(_3742_));
 sg13g2_a22oi_1 _5312_ (.Y(_0535_),
    .B1(_0532_),
    .B2(_0534_),
    .A2(_0529_),
    .A1(_0527_));
 sg13g2_buf_1 _5313_ (.A(_0535_),
    .X(_0536_));
 sg13g2_nand2_1 _5314_ (.Y(_0537_),
    .A(_4187_),
    .B(_4188_));
 sg13g2_inv_1 _5315_ (.Y(_0538_),
    .A(net305));
 sg13g2_nand2_1 _5316_ (.Y(_0539_),
    .A(net304),
    .B(\collatz.iter[44] ));
 sg13g2_or4_1 _5317_ (.A(_3544_),
    .B(_0538_),
    .C(_3892_),
    .D(_0539_),
    .X(_0540_));
 sg13g2_o21ai_1 _5318_ (.B1(_0540_),
    .Y(_0541_),
    .A1(net259),
    .A2(_0537_));
 sg13g2_buf_2 _5319_ (.A(_0541_),
    .X(_0542_));
 sg13g2_nand4_1 _5320_ (.B(_3691_),
    .C(net303),
    .A(_3690_),
    .Y(_0543_),
    .D(_3882_));
 sg13g2_inv_1 _5321_ (.Y(_0544_),
    .A(\collatz.iter[52] ));
 sg13g2_nand3_1 _5322_ (.B(_0217_),
    .C(_0218_),
    .A(_0544_),
    .Y(_0545_));
 sg13g2_nor2_1 _5323_ (.A(_3893_),
    .B(_3894_),
    .Y(_0546_));
 sg13g2_nand4_1 _5324_ (.B(net312),
    .C(net319),
    .A(net313),
    .Y(_0547_),
    .D(_0546_));
 sg13g2_inv_1 _5325_ (.Y(_0548_),
    .A(net319));
 sg13g2_nand3_1 _5326_ (.B(_4210_),
    .C(_4211_),
    .A(_0548_),
    .Y(_0549_));
 sg13g2_a22oi_1 _5327_ (.Y(_0550_),
    .B1(_0547_),
    .B2(_0549_),
    .A2(_0545_),
    .A1(_0543_));
 sg13g2_buf_2 _5328_ (.A(_0550_),
    .X(_0551_));
 sg13g2_buf_1 _5329_ (.A(_3533_),
    .X(_0552_));
 sg13g2_nand3_1 _5330_ (.B(net305),
    .C(_4194_),
    .A(_3842_),
    .Y(_0553_));
 sg13g2_nor2_1 _5331_ (.A(net288),
    .B(net305),
    .Y(_0554_));
 sg13g2_nand3_1 _5332_ (.B(_4197_),
    .C(_0554_),
    .A(net161),
    .Y(_0555_));
 sg13g2_o21ai_1 _5333_ (.B1(_0555_),
    .Y(_0556_),
    .A1(net161),
    .A2(_0553_));
 sg13g2_buf_1 _5334_ (.A(_0556_),
    .X(_0557_));
 sg13g2_nand4_1 _5335_ (.B(_0542_),
    .C(_0551_),
    .A(_0536_),
    .Y(_0558_),
    .D(_0557_));
 sg13g2_nand2_1 _5336_ (.Y(_0559_),
    .A(_0543_),
    .B(_0545_));
 sg13g2_inv_1 _5337_ (.Y(_0560_),
    .A(net184));
 sg13g2_a22oi_1 _5338_ (.Y(_0561_),
    .B1(net312),
    .B2(_0220_),
    .A2(_0210_),
    .A1(net313));
 sg13g2_o21ai_1 _5339_ (.B1(_0210_),
    .Y(_0562_),
    .A1(net258),
    .A2(net183));
 sg13g2_o21ai_1 _5340_ (.B1(_0562_),
    .Y(_0563_),
    .A1(_0560_),
    .A2(_0561_));
 sg13g2_inv_1 _5341_ (.Y(_0564_),
    .A(net187));
 sg13g2_a22oi_1 _5342_ (.Y(_0565_),
    .B1(net188),
    .B2(_4169_),
    .A2(_4165_),
    .A1(net183));
 sg13g2_o21ai_1 _5343_ (.B1(net191),
    .Y(_0566_),
    .A1(net188),
    .A2(_4169_));
 sg13g2_o21ai_1 _5344_ (.B1(_0566_),
    .Y(_0567_),
    .A1(_0564_),
    .A2(_0565_));
 sg13g2_a21o_1 _5345_ (.A2(_0563_),
    .A1(_0559_),
    .B1(_0567_),
    .X(_0568_));
 sg13g2_inv_1 _5346_ (.Y(_0569_),
    .A(net214));
 sg13g2_buf_1 _5347_ (.A(net305),
    .X(_0570_));
 sg13g2_a22oi_1 _5348_ (.Y(_0571_),
    .B1(net288),
    .B2(net160),
    .A2(_0552_),
    .A1(net232));
 sg13g2_o21ai_1 _5349_ (.B1(net161),
    .Y(_0572_),
    .A1(net288),
    .A2(net160));
 sg13g2_o21ai_1 _5350_ (.B1(_0572_),
    .Y(_0573_),
    .A1(_0569_),
    .A2(_0571_));
 sg13g2_buf_1 _5351_ (.A(_3544_),
    .X(_0574_));
 sg13g2_inv_1 _5352_ (.Y(_0575_),
    .A(net159));
 sg13g2_a22oi_1 _5353_ (.Y(_0576_),
    .B1(net304),
    .B2(_3703_),
    .A2(net186),
    .A1(_0570_));
 sg13g2_buf_1 _5354_ (.A(net304),
    .X(_0577_));
 sg13g2_o21ai_1 _5355_ (.B1(net186),
    .Y(_0578_),
    .A1(net158),
    .A2(net259));
 sg13g2_o21ai_1 _5356_ (.B1(_0578_),
    .Y(_0579_),
    .A1(_0575_),
    .A2(_0576_));
 sg13g2_a21o_1 _5357_ (.A2(_0573_),
    .A1(_0542_),
    .B1(_0579_),
    .X(_0580_));
 sg13g2_and2_1 _5358_ (.A(_0536_),
    .B(_0551_),
    .X(_0581_));
 sg13g2_inv_1 _5359_ (.Y(_0582_),
    .A(net307));
 sg13g2_a22oi_1 _5360_ (.Y(_0583_),
    .B1(_3741_),
    .B2(net162),
    .A2(net253),
    .A1(net190));
 sg13g2_o21ai_1 _5361_ (.B1(net253),
    .Y(_0584_),
    .A1(net189),
    .A2(net162));
 sg13g2_o21ai_1 _5362_ (.B1(_0584_),
    .Y(_0585_),
    .A1(_0582_),
    .A2(_0583_));
 sg13g2_nand2_1 _5363_ (.Y(_0586_),
    .A(_0527_),
    .B(_0529_));
 sg13g2_o21ai_1 _5364_ (.B1(net320),
    .Y(_0587_),
    .A1(net163),
    .A2(_0327_));
 sg13g2_a22oi_1 _5365_ (.Y(_0588_),
    .B1(net163),
    .B2(net174),
    .A2(net320),
    .A1(net162));
 sg13g2_nand2b_1 _5366_ (.Y(_0589_),
    .B(net195),
    .A_N(_0588_));
 sg13g2_nand2_1 _5367_ (.Y(_0590_),
    .A(_0587_),
    .B(_0589_));
 sg13g2_a21o_1 _5368_ (.A2(_0586_),
    .A1(_0585_),
    .B1(_0590_),
    .X(_0591_));
 sg13g2_a221oi_1 _5369_ (.B2(_0581_),
    .C1(_0591_),
    .B1(_0580_),
    .A1(_0536_),
    .Y(_0592_),
    .A2(_0568_));
 sg13g2_o21ai_1 _5370_ (.B1(_0592_),
    .Y(_0593_),
    .A1(_0525_),
    .A2(_0558_));
 sg13g2_nor2_1 _5371_ (.A(net275),
    .B(net252),
    .Y(_0594_));
 sg13g2_nand4_1 _5372_ (.B(net101),
    .C(net166),
    .A(net174),
    .Y(_0595_),
    .D(_0594_));
 sg13g2_nand3_1 _5373_ (.B(net116),
    .C(_3770_),
    .A(net213),
    .Y(_0596_));
 sg13g2_a22oi_1 _5374_ (.Y(_0597_),
    .B1(_0595_),
    .B2(_0596_),
    .A2(_0424_),
    .A1(_0421_));
 sg13g2_inv_1 _5375_ (.Y(_0598_),
    .A(net282));
 sg13g2_a22oi_1 _5376_ (.Y(_0599_),
    .B1(net245),
    .B2(net287),
    .A2(_3797_),
    .A1(net298));
 sg13g2_o21ai_1 _5377_ (.B1(_3797_),
    .Y(_0600_),
    .A1(net245),
    .A2(net287));
 sg13g2_o21ai_1 _5378_ (.B1(_0600_),
    .Y(_0601_),
    .A1(_0598_),
    .A2(_0599_));
 sg13g2_buf_1 _5379_ (.A(_0601_),
    .X(_0602_));
 sg13g2_a221oi_1 _5380_ (.B2(_0597_),
    .C1(_0602_),
    .B1(_0593_),
    .A1(_0425_),
    .Y(_0603_),
    .A2(_0430_));
 sg13g2_buf_1 _5381_ (.A(net317),
    .X(_0604_));
 sg13g2_and2_1 _5382_ (.A(\collatz.iter[74] ),
    .B(_3943_),
    .X(_0605_));
 sg13g2_buf_2 _5383_ (.A(_0605_),
    .X(_0606_));
 sg13g2_nand3_1 _5384_ (.B(_3875_),
    .C(_0606_),
    .A(net157),
    .Y(_0607_));
 sg13g2_nand3b_1 _5385_ (.B(_3695_),
    .C(_4110_),
    .Y(_0608_),
    .A_N(net208));
 sg13g2_and2_1 _5386_ (.A(_0607_),
    .B(_0608_),
    .X(_0609_));
 sg13g2_nand4_1 _5387_ (.B(_3847_),
    .C(net317),
    .A(net287),
    .Y(_0610_),
    .D(_4131_));
 sg13g2_inv_1 _5388_ (.Y(_0611_),
    .A(net317));
 sg13g2_nand4_1 _5389_ (.B(_3784_),
    .C(_0611_),
    .A(_3866_),
    .Y(_0612_),
    .D(_3848_));
 sg13g2_nand2_1 _5390_ (.Y(_0613_),
    .A(_0610_),
    .B(_0612_));
 sg13g2_nand2b_1 _5391_ (.Y(_0614_),
    .B(_0613_),
    .A_N(_0609_));
 sg13g2_buf_1 _5392_ (.A(net197),
    .X(_0615_));
 sg13g2_nand3_1 _5393_ (.B(net157),
    .C(net227),
    .A(net98),
    .Y(_0616_));
 sg13g2_o21ai_1 _5394_ (.B1(net295),
    .Y(_0617_),
    .A1(net192),
    .A2(net317));
 sg13g2_nand2_1 _5395_ (.Y(_0618_),
    .A(_0616_),
    .B(_0617_));
 sg13g2_a22oi_1 _5396_ (.Y(_0619_),
    .B1(net192),
    .B2(net157),
    .A2(net295),
    .A1(net287));
 sg13g2_buf_1 _5397_ (.A(_3874_),
    .X(_0620_));
 sg13g2_nand3_1 _5398_ (.B(net98),
    .C(net97),
    .A(net229),
    .Y(_0621_));
 sg13g2_nor2_1 _5399_ (.A(_0619_),
    .B(_0621_),
    .Y(_0622_));
 sg13g2_a221oi_1 _5400_ (.B2(_4110_),
    .C1(_0622_),
    .B1(_0618_),
    .A1(net98),
    .Y(_0623_),
    .A2(_0606_));
 sg13g2_buf_1 _5401_ (.A(_3694_),
    .X(_0624_));
 sg13g2_o21ai_1 _5402_ (.B1(net97),
    .Y(_0625_),
    .A1(net156),
    .A2(net208));
 sg13g2_nor2_1 _5403_ (.A(net193),
    .B(_0619_),
    .Y(_0626_));
 sg13g2_buf_1 _5404_ (.A(net157),
    .X(_0627_));
 sg13g2_and2_1 _5405_ (.A(net96),
    .B(_0606_),
    .X(_0628_));
 sg13g2_o21ai_1 _5406_ (.B1(_0628_),
    .Y(_0629_),
    .A1(_0618_),
    .A2(_0626_));
 sg13g2_and3_1 _5407_ (.X(_0630_),
    .A(_0623_),
    .B(_0625_),
    .C(_0629_));
 sg13g2_o21ai_1 _5408_ (.B1(_0630_),
    .Y(_0631_),
    .A1(_0603_),
    .A2(_0614_));
 sg13g2_and2_1 _5409_ (.A(_0412_),
    .B(_0414_),
    .X(_0632_));
 sg13g2_buf_1 _5410_ (.A(_0632_),
    .X(_0633_));
 sg13g2_buf_1 _5411_ (.A(net315),
    .X(_0634_));
 sg13g2_o21ai_1 _5412_ (.B1(_0345_),
    .Y(_0635_),
    .A1(net207),
    .A2(_0634_));
 sg13g2_o21ai_1 _5413_ (.B1(net167),
    .Y(_0636_),
    .A1(_0342_),
    .A2(_0416_));
 sg13g2_and2_1 _5414_ (.A(_0635_),
    .B(_0636_),
    .X(_0637_));
 sg13g2_or2_1 _5415_ (.X(_0638_),
    .B(net276),
    .A(net314));
 sg13g2_buf_1 _5416_ (.A(_0638_),
    .X(_0639_));
 sg13g2_nand2b_1 _5417_ (.Y(_0640_),
    .B(_0411_),
    .A_N(_0348_));
 sg13g2_a22oi_1 _5418_ (.Y(_0641_),
    .B1(_0640_),
    .B2(net111),
    .A2(_0639_),
    .A1(_4089_));
 sg13g2_o21ai_1 _5419_ (.B1(_0641_),
    .Y(_0642_),
    .A1(_0633_),
    .A2(_0637_));
 sg13g2_a21oi_1 _5420_ (.A1(_0420_),
    .A2(_0631_),
    .Y(_0643_),
    .B1(_0642_));
 sg13g2_inv_1 _5421_ (.Y(_0644_),
    .A(_3813_));
 sg13g2_nand3_1 _5422_ (.B(_4063_),
    .C(_4064_),
    .A(_0644_),
    .Y(_0645_));
 sg13g2_inv_1 _5423_ (.Y(_0646_),
    .A(_3899_));
 sg13g2_nand4_1 _5424_ (.B(net311),
    .C(_3813_),
    .A(_0646_),
    .Y(_0647_),
    .D(_4060_));
 sg13g2_buf_1 _5425_ (.A(_0647_),
    .X(_0648_));
 sg13g2_inv_1 _5426_ (.Y(_0649_),
    .A(_3898_));
 sg13g2_and2_1 _5427_ (.A(_3786_),
    .B(_3720_),
    .X(_0650_));
 sg13g2_buf_1 _5428_ (.A(_0650_),
    .X(_0651_));
 sg13g2_nand3_1 _5429_ (.B(_4073_),
    .C(_0651_),
    .A(_0649_),
    .Y(_0652_));
 sg13g2_nand3b_1 _5430_ (.B(_4068_),
    .C(_4069_),
    .Y(_0653_),
    .A_N(net311));
 sg13g2_a22oi_1 _5431_ (.Y(_0654_),
    .B1(_0652_),
    .B2(_0653_),
    .A2(_0648_),
    .A1(_0645_));
 sg13g2_buf_1 _5432_ (.A(_0654_),
    .X(_0655_));
 sg13g2_nand3_1 _5433_ (.B(_4052_),
    .C(_4053_),
    .A(_0397_),
    .Y(_0656_));
 sg13g2_nor2b_1 _5434_ (.A(net296),
    .B_N(_3813_),
    .Y(_0657_));
 sg13g2_nand3_1 _5435_ (.B(_4056_),
    .C(_0657_),
    .A(net200),
    .Y(_0658_));
 sg13g2_buf_1 _5436_ (.A(_3802_),
    .X(_0659_));
 sg13g2_nor2b_1 _5437_ (.A(_3853_),
    .B_N(net276),
    .Y(_0660_));
 sg13g2_nand3_1 _5438_ (.B(_4081_),
    .C(_0660_),
    .A(net154),
    .Y(_0661_));
 sg13g2_nand3_1 _5439_ (.B(_3803_),
    .C(_4077_),
    .A(net206),
    .Y(_0662_));
 sg13g2_a22oi_1 _5440_ (.Y(_0663_),
    .B1(_0661_),
    .B2(_0662_),
    .A2(_0658_),
    .A1(_0656_));
 sg13g2_nand2_1 _5441_ (.Y(_0664_),
    .A(_0655_),
    .B(_0663_));
 sg13g2_nand2_1 _5442_ (.Y(_0665_),
    .A(_0656_),
    .B(_0658_));
 sg13g2_nand2_1 _5443_ (.Y(_0666_),
    .A(_0645_),
    .B(_0648_));
 sg13g2_nand2_1 _5444_ (.Y(_0667_),
    .A(_0652_),
    .B(_0653_));
 sg13g2_inv_1 _5445_ (.Y(_0668_),
    .A(_3853_));
 sg13g2_buf_1 _5446_ (.A(_3801_),
    .X(_0669_));
 sg13g2_a22oi_1 _5447_ (.Y(_0670_),
    .B1(net153),
    .B2(net154),
    .A2(net206),
    .A1(net218));
 sg13g2_o21ai_1 _5448_ (.B1(net206),
    .Y(_0671_),
    .A1(net153),
    .A2(net154));
 sg13g2_o21ai_1 _5449_ (.B1(_0671_),
    .Y(_0672_),
    .A1(_0668_),
    .A2(_0670_));
 sg13g2_buf_1 _5450_ (.A(net311),
    .X(_0673_));
 sg13g2_o21ai_1 _5451_ (.B1(net224),
    .Y(_0674_),
    .A1(net243),
    .A2(_0673_));
 sg13g2_o21ai_1 _5452_ (.B1(_0364_),
    .Y(_0675_),
    .A1(_0363_),
    .A2(_0651_));
 sg13g2_nand2_1 _5453_ (.Y(_0676_),
    .A(_0674_),
    .B(_0675_));
 sg13g2_a21o_1 _5454_ (.A2(_0672_),
    .A1(_0667_),
    .B1(_0676_),
    .X(_0677_));
 sg13g2_buf_1 _5455_ (.A(net310),
    .X(_0678_));
 sg13g2_a22oi_1 _5456_ (.Y(_0679_),
    .B1(net151),
    .B2(net169),
    .A2(_4050_),
    .A1(net152));
 sg13g2_o21ai_1 _5457_ (.B1(_4050_),
    .Y(_0680_),
    .A1(net151),
    .A2(net169));
 sg13g2_o21ai_1 _5458_ (.B1(_0680_),
    .Y(_0681_),
    .A1(_0646_),
    .A2(_0679_));
 sg13g2_buf_1 _5459_ (.A(_0681_),
    .X(_0682_));
 sg13g2_a21o_1 _5460_ (.A2(_0677_),
    .A1(_0666_),
    .B1(_0682_),
    .X(_0683_));
 sg13g2_inv_1 _5461_ (.Y(_0684_),
    .A(net296));
 sg13g2_a22oi_1 _5462_ (.Y(_0685_),
    .B1(net235),
    .B2(_3696_),
    .A2(_3788_),
    .A1(net169));
 sg13g2_o21ai_1 _5463_ (.B1(_3788_),
    .Y(_0686_),
    .A1(net235),
    .A2(_4048_));
 sg13g2_o21ai_1 _5464_ (.B1(_0686_),
    .Y(_0687_),
    .A1(_0684_),
    .A2(_0685_));
 sg13g2_buf_1 _5465_ (.A(_0687_),
    .X(_0688_));
 sg13g2_a21oi_1 _5466_ (.A1(_0665_),
    .A2(_0683_),
    .Y(_0689_),
    .B1(_0688_));
 sg13g2_o21ai_1 _5467_ (.B1(_0689_),
    .Y(_0690_),
    .A1(_0643_),
    .A2(_0664_));
 sg13g2_xor2_1 _5468_ (.B(_0690_),
    .A(_0409_),
    .X(_0691_));
 sg13g2_buf_1 _5469_ (.A(net67),
    .X(_0692_));
 sg13g2_buf_1 _5470_ (.A(_0692_),
    .X(_0693_));
 sg13g2_buf_1 _5471_ (.A(_3697_),
    .X(_0694_));
 sg13g2_nor2_1 _5472_ (.A(net38),
    .B(_0694_),
    .Y(_0695_));
 sg13g2_a21oi_1 _5473_ (.A1(net39),
    .A2(_0691_),
    .Y(_0696_),
    .B1(_0695_));
 sg13g2_nor2_1 _5474_ (.A(net65),
    .B(_0696_),
    .Y(_0697_));
 sg13g2_buf_1 _5475_ (.A(ui_in[5]),
    .X(_0698_));
 sg13g2_buf_1 _5476_ (.A(_0698_),
    .X(_0699_));
 sg13g2_buf_1 _5477_ (.A(_0395_),
    .X(_0700_));
 sg13g2_inv_2 _5478_ (.Y(_0701_),
    .A(_3920_));
 sg13g2_nor2_1 _5479_ (.A(_0701_),
    .B(net20),
    .Y(_0702_));
 sg13g2_buf_1 _5480_ (.A(net203),
    .X(_0703_));
 sg13g2_buf_1 _5481_ (.A(net95),
    .X(_0704_));
 sg13g2_a221oi_1 _5482_ (.B2(_0702_),
    .C1(net76),
    .B1(net18),
    .A1(net266),
    .Y(_0705_),
    .A2(net20));
 sg13g2_nor3_1 _5483_ (.A(_0403_),
    .B(_0697_),
    .C(_0705_),
    .Y(_0030_));
 sg13g2_buf_1 _5484_ (.A(_3971_),
    .X(_0706_));
 sg13g2_buf_1 _5485_ (.A(ui_in[6]),
    .X(_0707_));
 sg13g2_inv_1 _5486_ (.Y(_0708_),
    .A(_3697_));
 sg13g2_nor2_1 _5487_ (.A(_0708_),
    .B(_0391_),
    .Y(_0709_));
 sg13g2_a22oi_1 _5488_ (.Y(_0710_),
    .B1(net19),
    .B2(_0709_),
    .A2(net20),
    .A1(net325));
 sg13g2_xor2_1 _5489_ (.B(net150),
    .A(net217),
    .X(_0711_));
 sg13g2_nand3_1 _5490_ (.B(_4056_),
    .C(_0407_),
    .A(_0684_),
    .Y(_0712_));
 sg13g2_buf_1 _5491_ (.A(_0712_),
    .X(_0713_));
 sg13g2_nand3_1 _5492_ (.B(_4052_),
    .C(_0408_),
    .A(net296),
    .Y(_0714_));
 sg13g2_buf_1 _5493_ (.A(_0714_),
    .X(_0715_));
 sg13g2_nand2_1 _5494_ (.Y(_0716_),
    .A(_0713_),
    .B(_0715_));
 sg13g2_buf_1 _5495_ (.A(_3899_),
    .X(_0717_));
 sg13g2_nand3_1 _5496_ (.B(_4053_),
    .C(_4063_),
    .A(net149),
    .Y(_0718_));
 sg13g2_nand3_1 _5497_ (.B(_4060_),
    .C(_0657_),
    .A(_0646_),
    .Y(_0719_));
 sg13g2_nand2_1 _5498_ (.Y(_0720_),
    .A(_0718_),
    .B(_0719_));
 sg13g2_a21oi_1 _5499_ (.A1(net170),
    .A2(net243),
    .Y(_0721_),
    .B1(net149));
 sg13g2_nor2b_1 _5500_ (.A(_0721_),
    .B_N(net152),
    .Y(_0722_));
 sg13g2_and2_1 _5501_ (.A(_3786_),
    .B(_3899_),
    .X(_0723_));
 sg13g2_o21ai_1 _5502_ (.B1(net224),
    .Y(_0724_),
    .A1(net152),
    .A2(_0723_));
 sg13g2_nand2b_1 _5503_ (.Y(_0725_),
    .B(_0724_),
    .A_N(_0722_));
 sg13g2_a21oi_1 _5504_ (.A1(net149),
    .A2(net151),
    .Y(_0726_),
    .B1(net168));
 sg13g2_nand2b_1 _5505_ (.Y(_0727_),
    .B(net169),
    .A_N(_0726_));
 sg13g2_and2_1 _5506_ (.A(net310),
    .B(net296),
    .X(_0728_));
 sg13g2_o21ai_1 _5507_ (.B1(net199),
    .Y(_0729_),
    .A1(net169),
    .A2(_0728_));
 sg13g2_nand2_1 _5508_ (.Y(_0730_),
    .A(_0727_),
    .B(_0729_));
 sg13g2_a21o_1 _5509_ (.A2(_0725_),
    .A1(_0720_),
    .B1(_0730_),
    .X(_0731_));
 sg13g2_a21oi_1 _5510_ (.A1(_3776_),
    .A2(net235),
    .Y(_0732_),
    .B1(net217));
 sg13g2_and2_1 _5511_ (.A(_3815_),
    .B(_3920_),
    .X(_0733_));
 sg13g2_o21ai_1 _5512_ (.B1(net242),
    .Y(_0734_),
    .A1(net200),
    .A2(_0733_));
 sg13g2_o21ai_1 _5513_ (.B1(_0734_),
    .Y(_0735_),
    .A1(_0397_),
    .A2(_0732_));
 sg13g2_buf_1 _5514_ (.A(_0735_),
    .X(_0736_));
 sg13g2_a21o_1 _5515_ (.A2(_0731_),
    .A1(_0716_),
    .B1(_0736_),
    .X(_0737_));
 sg13g2_nand4_1 _5516_ (.B(net114),
    .C(net193),
    .A(_0598_),
    .Y(_0738_),
    .D(_4133_));
 sg13g2_nand3_1 _5517_ (.B(_4136_),
    .C(_0423_),
    .A(net230),
    .Y(_0739_));
 sg13g2_nor2b_1 _5518_ (.A(_3754_),
    .B_N(_3676_),
    .Y(_0740_));
 sg13g2_nand3_1 _5519_ (.B(_0282_),
    .C(_0740_),
    .A(net177),
    .Y(_0741_));
 sg13g2_nand3_1 _5520_ (.B(_3684_),
    .C(_0288_),
    .A(net250),
    .Y(_0742_));
 sg13g2_nand2_1 _5521_ (.Y(_0743_),
    .A(_0741_),
    .B(_0742_));
 sg13g2_a21oi_1 _5522_ (.A1(net178),
    .A2(net237),
    .Y(_0744_),
    .B1(net251));
 sg13g2_and2_1 _5523_ (.A(_3808_),
    .B(_3751_),
    .X(_0745_));
 sg13g2_o21ai_1 _5524_ (.B1(net179),
    .Y(_0746_),
    .A1(net236),
    .A2(_0745_));
 sg13g2_o21ai_1 _5525_ (.B1(_0746_),
    .Y(_0747_),
    .A1(_0285_),
    .A2(_0744_));
 sg13g2_a21o_1 _5526_ (.A2(_3713_),
    .A1(net257),
    .B1(net256),
    .X(_0748_));
 sg13g2_a21o_1 _5527_ (.A2(net257),
    .A1(net283),
    .B1(_3713_),
    .X(_0749_));
 sg13g2_a22oi_1 _5528_ (.Y(_0750_),
    .B1(_0749_),
    .B2(net256),
    .A2(_0748_),
    .A1(net249));
 sg13g2_and3_1 _5529_ (.X(_0751_),
    .A(_3860_),
    .B(_3757_),
    .C(_3713_));
 sg13g2_o21ai_1 _5530_ (.B1(net284),
    .Y(_0752_),
    .A1(_0468_),
    .A2(_0751_));
 sg13g2_nand2_1 _5531_ (.Y(_0753_),
    .A(_0750_),
    .B(_0752_));
 sg13g2_nor2_1 _5532_ (.A(_3808_),
    .B(_3810_),
    .Y(_0754_));
 sg13g2_nand4_1 _5533_ (.B(net179),
    .C(_3751_),
    .A(_0292_),
    .Y(_0755_),
    .D(_0754_));
 sg13g2_or3_1 _5534_ (.A(_3751_),
    .B(_3716_),
    .C(_0477_),
    .X(_0756_));
 sg13g2_a22oi_1 _5535_ (.Y(_0757_),
    .B1(_0755_),
    .B2(_0756_),
    .A2(_0742_),
    .A1(_0741_));
 sg13g2_a21oi_1 _5536_ (.A1(_3752_),
    .A2(net177),
    .Y(_0758_),
    .B1(net250));
 sg13g2_and2_1 _5537_ (.A(_3667_),
    .B(net250),
    .X(_0759_));
 sg13g2_o21ai_1 _5538_ (.B1(net300),
    .Y(_0760_),
    .A1(net180),
    .A2(_0759_));
 sg13g2_o21ai_1 _5539_ (.B1(_0760_),
    .Y(_0761_),
    .A1(_0454_),
    .A2(_0758_));
 sg13g2_a221oi_1 _5540_ (.B2(_0757_),
    .C1(_0761_),
    .B1(_0753_),
    .A1(_0743_),
    .Y(_0762_),
    .A2(_0747_));
 sg13g2_buf_2 _5541_ (.A(_0762_),
    .X(_0763_));
 sg13g2_nand3_1 _5542_ (.B(net233),
    .C(_0457_),
    .A(net234),
    .Y(_0764_));
 sg13g2_nor2b_1 _5543_ (.A(net290),
    .B_N(net278),
    .Y(_0765_));
 sg13g2_nand3_1 _5544_ (.B(_0277_),
    .C(_0765_),
    .A(net164),
    .Y(_0766_));
 sg13g2_o21ai_1 _5545_ (.B1(_0766_),
    .Y(_0767_),
    .A1(_0461_),
    .A2(_0764_));
 sg13g2_inv_1 _5546_ (.Y(_0768_),
    .A(_0767_));
 sg13g2_nand3_1 _5547_ (.B(net216),
    .C(_0513_),
    .A(_3760_),
    .Y(_0769_));
 sg13g2_inv_1 _5548_ (.Y(_0770_),
    .A(net277));
 sg13g2_or2_1 _5549_ (.X(_0771_),
    .B(_3924_),
    .A(_3759_));
 sg13g2_or3_1 _5550_ (.A(_0770_),
    .B(_0515_),
    .C(_0771_),
    .X(_0772_));
 sg13g2_o21ai_1 _5551_ (.B1(_0772_),
    .Y(_0773_),
    .A1(net277),
    .A2(_0769_));
 sg13g2_buf_1 _5552_ (.A(_0773_),
    .X(_0774_));
 sg13g2_or3_1 _5553_ (.A(net290),
    .B(_3888_),
    .C(net267),
    .X(_0775_));
 sg13g2_nand2_1 _5554_ (.Y(_0776_),
    .A(net181),
    .B(net112));
 sg13g2_nand4_1 _5555_ (.B(net182),
    .C(net267),
    .A(net233),
    .Y(_0777_),
    .D(_0451_));
 sg13g2_o21ai_1 _5556_ (.B1(_0777_),
    .Y(_0778_),
    .A1(_0775_),
    .A2(_0776_));
 sg13g2_nand2_1 _5557_ (.Y(_0779_),
    .A(_0774_),
    .B(_0778_));
 sg13g2_nand3_1 _5558_ (.B(_4194_),
    .C(_0491_),
    .A(_0485_),
    .Y(_0780_));
 sg13g2_nand3_1 _5559_ (.B(_4197_),
    .C(_0204_),
    .A(_3927_),
    .Y(_0781_));
 sg13g2_nand3b_1 _5560_ (.B(_0207_),
    .C(_0496_),
    .Y(_0782_),
    .A_N(_3762_));
 sg13g2_buf_1 _5561_ (.A(_0782_),
    .X(_0783_));
 sg13g2_nand3_1 _5562_ (.B(_0205_),
    .C(_0263_),
    .A(_3762_),
    .Y(_0784_));
 sg13g2_a22oi_1 _5563_ (.Y(_0785_),
    .B1(_0783_),
    .B2(_0784_),
    .A2(_0781_),
    .A1(_0780_));
 sg13g2_buf_1 _5564_ (.A(_0785_),
    .X(_0786_));
 sg13g2_nand4_1 _5565_ (.B(_3842_),
    .C(net305),
    .A(_0569_),
    .Y(_0787_),
    .D(_3555_));
 sg13g2_nand4_1 _5566_ (.B(_0552_),
    .C(net159),
    .A(_3930_),
    .Y(_0788_),
    .D(_0554_));
 sg13g2_nand3_1 _5567_ (.B(_0244_),
    .C(_0265_),
    .A(net277),
    .Y(_0789_));
 sg13g2_nand3_1 _5568_ (.B(_0246_),
    .C(_0259_),
    .A(net291),
    .Y(_0790_));
 sg13g2_a22oi_1 _5569_ (.Y(_0791_),
    .B1(_0789_),
    .B2(_0790_),
    .A2(_0788_),
    .A1(_0787_));
 sg13g2_nand2_1 _5570_ (.Y(_0792_),
    .A(_0786_),
    .B(_0791_));
 sg13g2_nor4_2 _5571_ (.A(_0763_),
    .B(_0768_),
    .C(_0779_),
    .Y(_0793_),
    .D(_0792_));
 sg13g2_a21o_1 _5572_ (.A2(net248),
    .A1(net165),
    .B1(net220),
    .X(_0794_));
 sg13g2_a21o_1 _5573_ (.A2(net220),
    .A1(net115),
    .B1(net110),
    .X(_0795_));
 sg13g2_a22oi_1 _5574_ (.Y(_0796_),
    .B1(_0795_),
    .B2(_3727_),
    .A2(_0794_),
    .A1(net110));
 sg13g2_a21o_1 _5575_ (.A2(net278),
    .A1(_3755_),
    .B1(net290),
    .X(_0797_));
 sg13g2_a21o_1 _5576_ (.A2(net290),
    .A1(_3906_),
    .B1(_0238_),
    .X(_0798_));
 sg13g2_or2_1 _5577_ (.X(_0799_),
    .B(_3908_),
    .A(net292));
 sg13g2_a221oi_1 _5578_ (.B2(net234),
    .C1(_0799_),
    .B1(_0798_),
    .A1(net164),
    .Y(_0800_),
    .A2(_0797_));
 sg13g2_o21ai_1 _5579_ (.B1(net221),
    .Y(_0801_),
    .A1(net292),
    .A2(net267));
 sg13g2_nor2_1 _5580_ (.A(net267),
    .B(_3909_),
    .Y(_0802_));
 sg13g2_a21o_1 _5581_ (.A2(_0801_),
    .A1(_0500_),
    .B1(_0802_),
    .X(_0803_));
 sg13g2_a221oi_1 _5582_ (.B2(net234),
    .C1(_0775_),
    .B1(_0798_),
    .A1(net164),
    .Y(_0804_),
    .A2(_0797_));
 sg13g2_nor2_1 _5583_ (.A(net233),
    .B(_0799_),
    .Y(_0805_));
 sg13g2_nor4_2 _5584_ (.A(_0800_),
    .B(_0803_),
    .C(_0804_),
    .Y(_0806_),
    .D(_0805_));
 sg13g2_nand4_1 _5585_ (.B(_0774_),
    .C(_0806_),
    .A(_0786_),
    .Y(_0807_),
    .D(_0791_));
 sg13g2_o21ai_1 _5586_ (.B1(_0807_),
    .Y(_0808_),
    .A1(_0796_),
    .A2(_0792_));
 sg13g2_nor2_1 _5587_ (.A(_0793_),
    .B(_0808_),
    .Y(_0809_));
 sg13g2_nand3_1 _5588_ (.B(_4143_),
    .C(_0594_),
    .A(_4116_),
    .Y(_0810_));
 sg13g2_nor2_1 _5589_ (.A(net196),
    .B(net298),
    .Y(_0811_));
 sg13g2_nand4_1 _5590_ (.B(net116),
    .C(net230),
    .A(_3932_),
    .Y(_0812_),
    .D(_0811_));
 sg13g2_nand2_1 _5591_ (.Y(_0813_),
    .A(_0810_),
    .B(_0812_));
 sg13g2_nand4_1 _5592_ (.B(_0564_),
    .C(net319),
    .A(net312),
    .Y(_0814_),
    .D(_0546_));
 sg13g2_nand3_1 _5593_ (.B(_0218_),
    .C(_4210_),
    .A(_3893_),
    .Y(_0815_));
 sg13g2_nand2_1 _5594_ (.Y(_0816_),
    .A(_0814_),
    .B(_0815_));
 sg13g2_a21o_1 _5595_ (.A2(net304),
    .A1(_3544_),
    .B1(_3893_),
    .X(_0817_));
 sg13g2_a21o_1 _5596_ (.A2(_3893_),
    .A1(net304),
    .B1(net313),
    .X(_0818_));
 sg13g2_a22oi_1 _5597_ (.Y(_0819_),
    .B1(_0818_),
    .B2(_4209_),
    .A2(_0817_),
    .A1(net313));
 sg13g2_inv_1 _5598_ (.Y(_0820_),
    .A(_0819_));
 sg13g2_a21oi_1 _5599_ (.A1(_3893_),
    .A2(net312),
    .Y(_0821_),
    .B1(net187));
 sg13g2_and2_1 _5600_ (.A(net312),
    .B(net187),
    .X(_0822_));
 sg13g2_o21ai_1 _5601_ (.B1(net185),
    .Y(_0823_),
    .A1(net319),
    .A2(_0822_));
 sg13g2_o21ai_1 _5602_ (.B1(_0823_),
    .Y(_0824_),
    .A1(_0548_),
    .A2(_0821_));
 sg13g2_a21oi_1 _5603_ (.A1(_0816_),
    .A2(_0820_),
    .Y(_0825_),
    .B1(_0824_));
 sg13g2_nand4_1 _5604_ (.B(net320),
    .C(net275),
    .A(_3632_),
    .Y(_0826_),
    .D(_0526_));
 sg13g2_inv_1 _5605_ (.Y(_0827_),
    .A(\collatz.iter[61] ));
 sg13g2_nand4_1 _5606_ (.B(_0827_),
    .C(net299),
    .A(net293),
    .Y(_0828_),
    .D(_3650_));
 sg13g2_nand2_1 _5607_ (.Y(_0829_),
    .A(_0826_),
    .B(_0828_));
 sg13g2_inv_1 _5608_ (.Y(_0830_),
    .A(_3632_));
 sg13g2_nand4_1 _5609_ (.B(_0830_),
    .C(_3820_),
    .A(net302),
    .Y(_0831_),
    .D(_0531_));
 sg13g2_nor2b_1 _5610_ (.A(\collatz.iter[54] ),
    .B_N(net306),
    .Y(_0832_));
 sg13g2_nand4_1 _5611_ (.B(_3632_),
    .C(_0533_),
    .A(net307),
    .Y(_0833_),
    .D(_0832_));
 sg13g2_nand2_1 _5612_ (.Y(_0834_),
    .A(_0831_),
    .B(_0833_));
 sg13g2_and4_1 _5613_ (.A(net318),
    .B(_0582_),
    .C(net303),
    .D(_3882_),
    .X(_0835_));
 sg13g2_nand4_1 _5614_ (.B(net254),
    .C(_0544_),
    .A(_4176_),
    .Y(_0836_),
    .D(_0217_));
 sg13g2_nand2b_1 _5615_ (.Y(_0837_),
    .B(_0836_),
    .A_N(_0835_));
 sg13g2_nand3_1 _5616_ (.B(_0834_),
    .C(_0837_),
    .A(_0829_),
    .Y(_0838_));
 sg13g2_a21oi_1 _5617_ (.A1(net195),
    .A2(net293),
    .Y(_0839_),
    .B1(net275));
 sg13g2_a21oi_1 _5618_ (.A1(net293),
    .A2(net275),
    .Y(_0840_),
    .B1(_3767_));
 sg13g2_nand2b_1 _5619_ (.Y(_0841_),
    .B(_3641_),
    .A_N(_0840_));
 sg13g2_o21ai_1 _5620_ (.B1(_0841_),
    .Y(_0842_),
    .A1(_4117_),
    .A2(_0839_));
 sg13g2_a21oi_1 _5621_ (.A1(net307),
    .A2(net302),
    .Y(_0843_),
    .B1(_3632_));
 sg13g2_nand2b_1 _5622_ (.Y(_0844_),
    .B(net294),
    .A_N(_0843_));
 sg13g2_a21oi_1 _5623_ (.A1(net302),
    .A2(_3632_),
    .Y(_0845_),
    .B1(net294));
 sg13g2_nand2b_1 _5624_ (.Y(_0846_),
    .B(_3730_),
    .A_N(_0845_));
 sg13g2_a22oi_1 _5625_ (.Y(_0847_),
    .B1(_0826_),
    .B2(_0828_),
    .A2(_0846_),
    .A1(_0844_));
 sg13g2_a21o_1 _5626_ (.A2(net318),
    .A1(_3880_),
    .B1(_3728_),
    .X(_0848_));
 sg13g2_a21o_1 _5627_ (.A2(_3728_),
    .A1(net318),
    .B1(_3740_),
    .X(_0849_));
 sg13g2_a22oi_1 _5628_ (.Y(_0850_),
    .B1(_0849_),
    .B2(_3881_),
    .A2(_0848_),
    .A1(_3740_));
 sg13g2_buf_1 _5629_ (.A(_0850_),
    .X(_0851_));
 sg13g2_a221oi_1 _5630_ (.B2(_0833_),
    .C1(_0851_),
    .B1(_0831_),
    .A1(_0826_),
    .Y(_0852_),
    .A2(_0828_));
 sg13g2_nor3_1 _5631_ (.A(_0842_),
    .B(_0847_),
    .C(_0852_),
    .Y(_0853_));
 sg13g2_o21ai_1 _5632_ (.B1(_0853_),
    .Y(_0854_),
    .A1(_0825_),
    .A2(_0838_));
 sg13g2_and2_1 _5633_ (.A(_0780_),
    .B(_0781_),
    .X(_0855_));
 sg13g2_a21o_1 _5634_ (.A2(_3885_),
    .A1(_3927_),
    .B1(_3929_),
    .X(_0856_));
 sg13g2_a21o_1 _5635_ (.A2(_3929_),
    .A1(_3885_),
    .B1(_3840_),
    .X(_0857_));
 sg13g2_a22oi_1 _5636_ (.Y(_0858_),
    .B1(_0857_),
    .B2(_3796_),
    .A2(_0856_),
    .A1(net289));
 sg13g2_buf_1 _5637_ (.A(_0858_),
    .X(_0859_));
 sg13g2_a21o_1 _5638_ (.A2(net291),
    .A1(net277),
    .B1(_3763_),
    .X(_0860_));
 sg13g2_a21o_1 _5639_ (.A2(_3762_),
    .A1(net291),
    .B1(_3826_),
    .X(_0861_));
 sg13g2_a22oi_1 _5640_ (.Y(_0862_),
    .B1(_0861_),
    .B2(net241),
    .A2(_0860_),
    .A1(_0318_));
 sg13g2_a21o_1 _5641_ (.A2(_0784_),
    .A1(_0783_),
    .B1(_0862_),
    .X(_0863_));
 sg13g2_a21o_1 _5642_ (.A2(_3793_),
    .A1(_3762_),
    .B1(net215),
    .X(_0864_));
 sg13g2_a21o_1 _5643_ (.A2(_3928_),
    .A1(_3793_),
    .B1(_3883_),
    .X(_0865_));
 sg13g2_a22oi_1 _5644_ (.Y(_0866_),
    .B1(_0865_),
    .B2(_3765_),
    .A2(_0864_),
    .A1(_3884_));
 sg13g2_and2_1 _5645_ (.A(_0859_),
    .B(_0866_),
    .X(_0867_));
 sg13g2_and2_1 _5646_ (.A(_0787_),
    .B(_0788_),
    .X(_0868_));
 sg13g2_a221oi_1 _5647_ (.B2(_0867_),
    .C1(_0868_),
    .B1(_0863_),
    .A1(_0855_),
    .Y(_0869_),
    .A2(_0859_));
 sg13g2_o21ai_1 _5648_ (.B1(_0575_),
    .Y(_0870_),
    .A1(_0569_),
    .A2(_4196_));
 sg13g2_o21ai_1 _5649_ (.B1(_0538_),
    .Y(_0871_),
    .A1(_4196_),
    .A2(_0575_));
 sg13g2_a22oi_1 _5650_ (.Y(_0872_),
    .B1(_0871_),
    .B2(net161),
    .A2(_0870_),
    .A1(net160));
 sg13g2_a21o_1 _5651_ (.A2(_3768_),
    .A1(net275),
    .B1(net282),
    .X(_0873_));
 sg13g2_a21o_1 _5652_ (.A2(net282),
    .A1(_4115_),
    .B1(_3769_),
    .X(_0874_));
 sg13g2_a22oi_1 _5653_ (.Y(_0875_),
    .B1(_0874_),
    .B2(_3733_),
    .A2(_0873_),
    .A1(_3769_));
 sg13g2_buf_1 _5654_ (.A(_0875_),
    .X(_0876_));
 sg13g2_nand3b_1 _5655_ (.B(_0872_),
    .C(_0876_),
    .Y(_0877_),
    .A_N(_0869_));
 sg13g2_a21oi_1 _5656_ (.A1(_0813_),
    .A2(_0854_),
    .Y(_0878_),
    .B1(_0877_));
 sg13g2_nand2_2 _5657_ (.Y(_0879_),
    .A(_0829_),
    .B(_0834_));
 sg13g2_nor2b_1 _5658_ (.A(_0879_),
    .B_N(_0813_),
    .Y(_0880_));
 sg13g2_nor2b_1 _5659_ (.A(_0835_),
    .B_N(_0836_),
    .Y(_0881_));
 sg13g2_and2_1 _5660_ (.A(_0814_),
    .B(_0815_),
    .X(_0882_));
 sg13g2_buf_1 _5661_ (.A(_0882_),
    .X(_0883_));
 sg13g2_nor2_1 _5662_ (.A(net186),
    .B(_0213_),
    .Y(_0884_));
 sg13g2_nor2_1 _5663_ (.A(net159),
    .B(_0539_),
    .Y(_0885_));
 sg13g2_and2_1 _5664_ (.A(net159),
    .B(_4187_),
    .X(_0886_));
 sg13g2_a22oi_1 _5665_ (.Y(_0887_),
    .B1(_0886_),
    .B2(_4211_),
    .A2(_0885_),
    .A1(_0884_));
 sg13g2_buf_1 _5666_ (.A(_0887_),
    .X(_0888_));
 sg13g2_nor3_1 _5667_ (.A(_0881_),
    .B(_0883_),
    .C(_0888_),
    .Y(_0889_));
 sg13g2_inv_1 _5668_ (.Y(_0890_),
    .A(_0876_));
 sg13g2_a221oi_1 _5669_ (.B2(_0889_),
    .C1(_0890_),
    .B1(_0880_),
    .A1(_0813_),
    .Y(_0891_),
    .A2(_0854_));
 sg13g2_a221oi_1 _5670_ (.B2(_0878_),
    .C1(_0891_),
    .B1(_0809_),
    .A1(_0738_),
    .Y(_0892_),
    .A2(_0739_));
 sg13g2_buf_1 _5671_ (.A(_0892_),
    .X(_0893_));
 sg13g2_buf_1 _5672_ (.A(_3847_),
    .X(_0894_));
 sg13g2_inv_1 _5673_ (.Y(_0895_),
    .A(_4106_));
 sg13g2_nand4_1 _5674_ (.B(_0895_),
    .C(_0604_),
    .A(net148),
    .Y(_0896_),
    .D(_4131_));
 sg13g2_nand2_1 _5675_ (.Y(_0897_),
    .A(net244),
    .B(net197));
 sg13g2_or2_1 _5676_ (.X(_0898_),
    .B(_3693_),
    .A(_3847_));
 sg13g2_buf_1 _5677_ (.A(_0898_),
    .X(_0899_));
 sg13g2_or3_1 _5678_ (.A(net193),
    .B(_0897_),
    .C(_0899_),
    .X(_0900_));
 sg13g2_and2_1 _5679_ (.A(_0896_),
    .B(_0900_),
    .X(_0901_));
 sg13g2_buf_1 _5680_ (.A(_0901_),
    .X(_0902_));
 sg13g2_a22oi_1 _5681_ (.Y(_0903_),
    .B1(_0718_),
    .B2(_0719_),
    .A2(_0715_),
    .A1(_0713_));
 sg13g2_nand2_1 _5682_ (.Y(_0904_),
    .A(_3900_),
    .B(_0651_));
 sg13g2_nand3_1 _5683_ (.B(_4064_),
    .C(_4069_),
    .A(net170),
    .Y(_0905_));
 sg13g2_nand2_1 _5684_ (.Y(_0906_),
    .A(_0904_),
    .B(_0905_));
 sg13g2_nand2_1 _5685_ (.Y(_0907_),
    .A(_0903_),
    .B(_0906_));
 sg13g2_nor3_1 _5686_ (.A(net197),
    .B(net227),
    .C(net269),
    .Y(_0908_));
 sg13g2_nor2_1 _5687_ (.A(net316),
    .B(_3943_),
    .Y(_0909_));
 sg13g2_and3_1 _5688_ (.X(_0910_),
    .A(net197),
    .B(net227),
    .C(_4097_));
 sg13g2_a22oi_1 _5689_ (.Y(_0911_),
    .B1(_0909_),
    .B2(_0910_),
    .A2(_0606_),
    .A1(_0908_));
 sg13g2_nand3_1 _5690_ (.B(_4068_),
    .C(_4078_),
    .A(net171),
    .Y(_0912_));
 sg13g2_nand3_1 _5691_ (.B(_4073_),
    .C(_4081_),
    .A(_0668_),
    .Y(_0913_));
 sg13g2_nand2_1 _5692_ (.Y(_0914_),
    .A(_0912_),
    .B(_0913_));
 sg13g2_nand3b_1 _5693_ (.B(_3835_),
    .C(_0416_),
    .Y(_0915_),
    .A_N(_3915_));
 sg13g2_nor2b_1 _5694_ (.A(_3945_),
    .B_N(_3915_),
    .Y(_0916_));
 sg13g2_nand3_1 _5695_ (.B(_4091_),
    .C(_0916_),
    .A(net269),
    .Y(_0917_));
 sg13g2_or4_1 _5696_ (.A(_3916_),
    .B(_4089_),
    .C(_3853_),
    .D(_0411_),
    .X(_0918_));
 sg13g2_nor2b_1 _5697_ (.A(net314),
    .B_N(_3852_),
    .Y(_0919_));
 sg13g2_nand3_1 _5698_ (.B(_4077_),
    .C(_0919_),
    .A(_3916_),
    .Y(_0920_));
 sg13g2_a22oi_1 _5699_ (.Y(_0921_),
    .B1(_0918_),
    .B2(_0920_),
    .A2(_0917_),
    .A1(_0915_));
 sg13g2_buf_1 _5700_ (.A(_0921_),
    .X(_0922_));
 sg13g2_nand3b_1 _5701_ (.B(_0914_),
    .C(_0922_),
    .Y(_0923_),
    .A_N(_0911_));
 sg13g2_buf_1 _5702_ (.A(_0923_),
    .X(_0924_));
 sg13g2_or2_1 _5703_ (.X(_0925_),
    .B(_0924_),
    .A(_0907_));
 sg13g2_nor2_1 _5704_ (.A(_0902_),
    .B(_0925_),
    .Y(_0926_));
 sg13g2_a21o_1 _5705_ (.A2(net316),
    .A1(net197),
    .B1(_4097_),
    .X(_0927_));
 sg13g2_a21o_1 _5706_ (.A2(net269),
    .A1(net316),
    .B1(_3943_),
    .X(_0928_));
 sg13g2_a22oi_1 _5707_ (.Y(_0929_),
    .B1(_0928_),
    .B2(net227),
    .A2(_0927_),
    .A1(net208));
 sg13g2_a21oi_1 _5708_ (.A1(_0915_),
    .A2(_0917_),
    .Y(_0930_),
    .B1(_0929_));
 sg13g2_a21o_1 _5709_ (.A2(_3945_),
    .A1(net269),
    .B1(net219),
    .X(_0931_));
 sg13g2_a21o_1 _5710_ (.A2(net219),
    .A1(_3945_),
    .B1(net315),
    .X(_0932_));
 sg13g2_a22oi_1 _5711_ (.Y(_0933_),
    .B1(_0932_),
    .B2(net173),
    .A2(_0931_),
    .A1(net155));
 sg13g2_nand3b_1 _5712_ (.B(_0933_),
    .C(_3854_),
    .Y(_0934_),
    .A_N(_0930_));
 sg13g2_a21o_1 _5713_ (.A2(_0934_),
    .A1(_0639_),
    .B1(net111),
    .X(_0935_));
 sg13g2_nor2b_1 _5714_ (.A(_0930_),
    .B_N(_0933_),
    .Y(_0936_));
 sg13g2_o21ai_1 _5715_ (.B1(net218),
    .Y(_0937_),
    .A1(net314),
    .A2(_3853_));
 sg13g2_nor2_1 _5716_ (.A(_0355_),
    .B(net218),
    .Y(_0938_));
 sg13g2_a21o_1 _5717_ (.A2(_0937_),
    .A1(_4086_),
    .B1(_0938_),
    .X(_0939_));
 sg13g2_a221oi_1 _5718_ (.B2(_0413_),
    .C1(_0939_),
    .B1(_0936_),
    .A1(_0912_),
    .Y(_0940_),
    .A2(_0913_));
 sg13g2_a21o_1 _5719_ (.A2(net153),
    .A1(net171),
    .B1(net170),
    .X(_0941_));
 sg13g2_a21o_1 _5720_ (.A2(net170),
    .A1(net153),
    .B1(net154),
    .X(_0942_));
 sg13g2_a22oi_1 _5721_ (.Y(_0943_),
    .B1(_0942_),
    .B2(net206),
    .A2(_0941_),
    .A1(_0659_));
 sg13g2_inv_1 _5722_ (.Y(_0944_),
    .A(_0943_));
 sg13g2_a21oi_1 _5723_ (.A1(_0935_),
    .A2(_0940_),
    .Y(_0945_),
    .B1(_0944_));
 sg13g2_inv_1 _5724_ (.Y(_0946_),
    .A(_4155_));
 sg13g2_inv_1 _5725_ (.Y(_0947_),
    .A(net287));
 sg13g2_o21ai_1 _5726_ (.B1(_0947_),
    .Y(_0948_),
    .A1(_4148_),
    .A2(net193));
 sg13g2_o21ai_1 _5727_ (.B1(net193),
    .Y(_0949_),
    .A1(_0598_),
    .A2(_4148_));
 sg13g2_buf_1 _5728_ (.A(_3846_),
    .X(_0950_));
 sg13g2_a22oi_1 _5729_ (.Y(_0951_),
    .B1(_0949_),
    .B2(net147),
    .A2(_0948_),
    .A1(net238));
 sg13g2_o21ai_1 _5730_ (.B1(_0895_),
    .Y(_0952_),
    .A1(_0946_),
    .A2(_0951_));
 sg13g2_nand2_1 _5731_ (.Y(_0953_),
    .A(net148),
    .B(net96));
 sg13g2_o21ai_1 _5732_ (.B1(_0953_),
    .Y(_0954_),
    .A1(_0897_),
    .A2(_0951_));
 sg13g2_a21oi_1 _5733_ (.A1(net192),
    .A2(net197),
    .Y(_0955_),
    .B1(net157));
 sg13g2_nor2_1 _5734_ (.A(_4112_),
    .B(_0955_),
    .Y(_0956_));
 sg13g2_a221oi_1 _5735_ (.B2(net229),
    .C1(_0956_),
    .B1(_0954_),
    .A1(net96),
    .Y(_0957_),
    .A2(_0952_));
 sg13g2_buf_1 _5736_ (.A(_0957_),
    .X(_0958_));
 sg13g2_or2_1 _5737_ (.X(_0959_),
    .B(_0925_),
    .A(_0958_));
 sg13g2_o21ai_1 _5738_ (.B1(_0959_),
    .Y(_0960_),
    .A1(_0907_),
    .A2(_0945_));
 sg13g2_a21oi_1 _5739_ (.A1(_0893_),
    .A2(_0926_),
    .Y(_0961_),
    .B1(_0960_));
 sg13g2_nand2b_1 _5740_ (.Y(_0962_),
    .B(_0961_),
    .A_N(_0737_));
 sg13g2_xnor2_1 _5741_ (.Y(_0963_),
    .A(_0711_),
    .B(_0962_));
 sg13g2_buf_1 _5742_ (.A(_3447_),
    .X(_0964_));
 sg13g2_nor2_1 _5743_ (.A(net52),
    .B(net146),
    .Y(_0965_));
 sg13g2_a21oi_1 _5744_ (.A1(net50),
    .A2(_0963_),
    .Y(_0966_),
    .B1(_0965_));
 sg13g2_nand2_1 _5745_ (.Y(_0967_),
    .A(net80),
    .B(_0966_));
 sg13g2_o21ai_1 _5746_ (.B1(_0967_),
    .Y(_0968_),
    .A1(net75),
    .A2(_0710_));
 sg13g2_and2_1 _5747_ (.A(_4043_),
    .B(_0968_),
    .X(_0031_));
 sg13g2_xnor2_1 _5748_ (.Y(_0969_),
    .A(net146),
    .B(net150));
 sg13g2_and2_1 _5749_ (.A(_3696_),
    .B(_3697_),
    .X(_0970_));
 sg13g2_o21ai_1 _5750_ (.B1(net242),
    .Y(_0971_),
    .A1(_0733_),
    .A2(_0970_));
 sg13g2_o21ai_1 _5751_ (.B1(_0971_),
    .Y(_0972_),
    .A1(_0701_),
    .A2(_3698_));
 sg13g2_a21oi_1 _5752_ (.A1(net152),
    .A2(net310),
    .Y(_0973_),
    .B1(_0723_));
 sg13g2_o21ai_1 _5753_ (.B1(net149),
    .Y(_0974_),
    .A1(net152),
    .A2(net310));
 sg13g2_o21ai_1 _5754_ (.B1(_0974_),
    .Y(_0975_),
    .A1(_0649_),
    .A2(_0973_));
 sg13g2_buf_1 _5755_ (.A(_0975_),
    .X(_0976_));
 sg13g2_nand3_1 _5756_ (.B(_4059_),
    .C(_0651_),
    .A(net310),
    .Y(_0977_));
 sg13g2_nand3_1 _5757_ (.B(_3722_),
    .C(_4069_),
    .A(_0717_),
    .Y(_0978_));
 sg13g2_a22oi_1 _5758_ (.Y(_0979_),
    .B1(net154),
    .B2(_3786_),
    .A2(_3896_),
    .A1(net153));
 sg13g2_nand2b_1 _5759_ (.Y(_0980_),
    .B(_3948_),
    .A_N(_0979_));
 sg13g2_o21ai_1 _5760_ (.B1(net170),
    .Y(_0981_),
    .A1(net154),
    .A2(net243));
 sg13g2_a22oi_1 _5761_ (.Y(_0982_),
    .B1(_0980_),
    .B2(_0981_),
    .A2(_0978_),
    .A1(_0977_));
 sg13g2_nand3_1 _5762_ (.B(_4056_),
    .C(_0407_),
    .A(_0694_),
    .Y(_0983_));
 sg13g2_nand3_1 _5763_ (.B(_3698_),
    .C(_4052_),
    .A(_3920_),
    .Y(_0984_));
 sg13g2_nand2_1 _5764_ (.Y(_0985_),
    .A(net168),
    .B(_3817_));
 sg13g2_and2_1 _5765_ (.A(_3813_),
    .B(net235),
    .X(_0986_));
 sg13g2_buf_1 _5766_ (.A(_0986_),
    .X(_0987_));
 sg13g2_o21ai_1 _5767_ (.B1(net199),
    .Y(_0988_),
    .A1(_0987_),
    .A2(_0728_));
 sg13g2_a22oi_1 _5768_ (.Y(_0989_),
    .B1(_0985_),
    .B2(_0988_),
    .A2(_0984_),
    .A1(_0983_));
 sg13g2_nor4_2 _5769_ (.A(_0972_),
    .B(_0976_),
    .C(_0982_),
    .Y(_0990_),
    .D(_0989_));
 sg13g2_nand2_1 _5770_ (.Y(_0991_),
    .A(_0977_),
    .B(_0978_));
 sg13g2_nand3_1 _5771_ (.B(_4073_),
    .C(_4081_),
    .A(net243),
    .Y(_0992_));
 sg13g2_nand3b_1 _5772_ (.B(_4068_),
    .C(_4078_),
    .Y(_0993_),
    .A_N(net243));
 sg13g2_nand2_1 _5773_ (.Y(_0994_),
    .A(_0992_),
    .B(_0993_));
 sg13g2_buf_2 _5774_ (.A(_0994_),
    .X(_0995_));
 sg13g2_nand2_1 _5775_ (.Y(_0996_),
    .A(_0991_),
    .B(_0995_));
 sg13g2_nand4_1 _5776_ (.B(net268),
    .C(net181),
    .A(_0235_),
    .Y(_0997_),
    .D(_0765_));
 sg13g2_nand3_1 _5777_ (.B(_3824_),
    .C(_0272_),
    .A(net290),
    .Y(_0998_));
 sg13g2_inv_1 _5778_ (.Y(_0999_),
    .A(net292));
 sg13g2_nand4_1 _5779_ (.B(_0999_),
    .C(_0249_),
    .A(net182),
    .Y(_1000_),
    .D(_0250_));
 sg13g2_nand4_1 _5780_ (.B(_3909_),
    .C(_3760_),
    .A(net181),
    .Y(_1001_),
    .D(_3889_));
 sg13g2_a22oi_1 _5781_ (.Y(_1002_),
    .B1(_1000_),
    .B2(_1001_),
    .A2(_0998_),
    .A1(_0997_));
 sg13g2_a21oi_1 _5782_ (.A1(net180),
    .A2(net222),
    .Y(_1003_),
    .B1(_0759_));
 sg13g2_o21ai_1 _5783_ (.B1(net250),
    .Y(_1004_),
    .A1(_0276_),
    .A2(_3907_));
 sg13g2_o21ai_1 _5784_ (.B1(_1004_),
    .Y(_1005_),
    .A1(_0275_),
    .A2(_1003_));
 sg13g2_a21oi_1 _5785_ (.A1(net236),
    .A2(net177),
    .Y(_1006_),
    .B1(_0745_));
 sg13g2_o21ai_1 _5786_ (.B1(net251),
    .Y(_1007_),
    .A1(net236),
    .A2(net177));
 sg13g2_o21ai_1 _5787_ (.B1(_1007_),
    .Y(_1008_),
    .A1(_0281_),
    .A2(_1006_));
 sg13g2_nand4_1 _5788_ (.B(_3751_),
    .C(_0286_),
    .A(_0284_),
    .Y(_1009_),
    .D(_0754_));
 sg13g2_nor2b_1 _5789_ (.A(_3751_),
    .B_N(_3808_),
    .Y(_1010_));
 sg13g2_nand4_1 _5790_ (.B(_3810_),
    .C(_3667_),
    .A(_0281_),
    .Y(_1011_),
    .D(_1010_));
 sg13g2_nand3b_1 _5791_ (.B(_0293_),
    .C(_0751_),
    .Y(_1012_),
    .A_N(_3709_));
 sg13g2_nand3_1 _5792_ (.B(_0290_),
    .C(_0468_),
    .A(net237),
    .Y(_1013_));
 sg13g2_nor2b_1 _5793_ (.A(_3757_),
    .B_N(_3860_),
    .Y(_1014_));
 sg13g2_a21oi_1 _5794_ (.A1(_0468_),
    .A2(_1014_),
    .Y(_1015_),
    .B1(net284));
 sg13g2_a221oi_1 _5795_ (.B2(_1013_),
    .C1(_1015_),
    .B1(_1012_),
    .A1(_1009_),
    .Y(_1016_),
    .A2(_1011_));
 sg13g2_a22oi_1 _5796_ (.Y(_1017_),
    .B1(net256),
    .B2(net237),
    .A2(_3713_),
    .A1(_3709_));
 sg13g2_nand2b_1 _5797_ (.Y(_1018_),
    .B(_3758_),
    .A_N(_1017_));
 sg13g2_nand2_1 _5798_ (.Y(_1019_),
    .A(net178),
    .B(_0471_));
 sg13g2_a22oi_1 _5799_ (.Y(_1020_),
    .B1(_1018_),
    .B2(_1019_),
    .A2(_1011_),
    .A1(_1009_));
 sg13g2_or3_1 _5800_ (.A(_1008_),
    .B(_1016_),
    .C(_1020_),
    .X(_1021_));
 sg13g2_buf_1 _5801_ (.A(_1021_),
    .X(_1022_));
 sg13g2_or4_1 _5802_ (.A(_0275_),
    .B(_0461_),
    .C(net180),
    .D(net278),
    .X(_1023_));
 sg13g2_nand4_1 _5803_ (.B(net177),
    .C(_3907_),
    .A(_0275_),
    .Y(_1024_),
    .D(_0740_));
 sg13g2_o21ai_1 _5804_ (.B1(_1024_),
    .Y(_1025_),
    .A1(_0303_),
    .A2(_1023_));
 sg13g2_and2_1 _5805_ (.A(_1002_),
    .B(_1025_),
    .X(_1026_));
 sg13g2_a22oi_1 _5806_ (.Y(_1027_),
    .B1(_0238_),
    .B2(_3823_),
    .A2(_3838_),
    .A1(_3906_));
 sg13g2_o21ai_1 _5807_ (.B1(_3838_),
    .Y(_1028_),
    .A1(net268),
    .A2(_3823_));
 sg13g2_o21ai_1 _5808_ (.B1(_1028_),
    .Y(_1029_),
    .A1(_0235_),
    .A2(_1027_));
 sg13g2_inv_1 _5809_ (.Y(_1030_),
    .A(_3889_));
 sg13g2_o21ai_1 _5810_ (.B1(_1030_),
    .Y(_1031_),
    .A1(_0517_),
    .A2(_1029_));
 sg13g2_o21ai_1 _5811_ (.B1(_0517_),
    .Y(_1032_),
    .A1(net165),
    .A2(_1029_));
 sg13g2_a21oi_1 _5812_ (.A1(net112),
    .A2(net115),
    .Y(_1033_),
    .B1(net165));
 sg13g2_a221oi_1 _5813_ (.B2(_0500_),
    .C1(_1033_),
    .B1(_1032_),
    .A1(_0999_),
    .Y(_1034_),
    .A2(_1031_));
 sg13g2_a221oi_1 _5814_ (.B2(_1026_),
    .C1(_1034_),
    .B1(_1022_),
    .A1(_1002_),
    .Y(_1035_),
    .A2(_1005_));
 sg13g2_buf_2 _5815_ (.A(_1035_),
    .X(_1036_));
 sg13g2_nand4_1 _5816_ (.B(net259),
    .C(net258),
    .A(net158),
    .Y(_1037_),
    .D(_0884_));
 sg13g2_nand3_1 _5817_ (.B(_3707_),
    .C(_4187_),
    .A(net184),
    .Y(_1038_));
 sg13g2_nand2_1 _5818_ (.Y(_1039_),
    .A(_1037_),
    .B(_1038_));
 sg13g2_nand3_1 _5819_ (.B(net159),
    .C(_3739_),
    .A(net161),
    .Y(_1040_));
 sg13g2_nand4_1 _5820_ (.B(net160),
    .C(net158),
    .A(net231),
    .Y(_1041_),
    .D(_3555_));
 sg13g2_o21ai_1 _5821_ (.B1(_1041_),
    .Y(_1042_),
    .A1(net231),
    .A2(_1040_));
 sg13g2_nand2_2 _5822_ (.Y(_1043_),
    .A(_1039_),
    .B(_1042_));
 sg13g2_nand3_1 _5823_ (.B(_4194_),
    .C(_0491_),
    .A(net231),
    .Y(_1044_));
 sg13g2_nor2_1 _5824_ (.A(net232),
    .B(net231),
    .Y(_1045_));
 sg13g2_nand3_1 _5825_ (.B(_1045_),
    .C(_0204_),
    .A(net214),
    .Y(_1046_));
 sg13g2_nand2_1 _5826_ (.Y(_1047_),
    .A(_1044_),
    .B(_1046_));
 sg13g2_nand3_1 _5827_ (.B(_0207_),
    .C(_0496_),
    .A(_3886_),
    .Y(_1048_));
 sg13g2_nand3_1 _5828_ (.B(_3887_),
    .C(_0263_),
    .A(net215),
    .Y(_1049_));
 sg13g2_nand2_1 _5829_ (.Y(_1050_),
    .A(_1048_),
    .B(_1049_));
 sg13g2_nand2_1 _5830_ (.Y(_1051_),
    .A(_1047_),
    .B(_1050_));
 sg13g2_nand3b_1 _5831_ (.B(_0244_),
    .C(_0265_),
    .Y(_1052_),
    .A_N(net240));
 sg13g2_nand4_1 _5832_ (.B(net176),
    .C(net240),
    .A(_0256_),
    .Y(_1053_),
    .D(_0259_));
 sg13g2_and3_1 _5833_ (.X(_1054_),
    .A(net115),
    .B(_0770_),
    .C(net110));
 sg13g2_nor3_1 _5834_ (.A(_0252_),
    .B(net176),
    .C(_0771_),
    .Y(_1055_));
 sg13g2_a22oi_1 _5835_ (.Y(_1056_),
    .B1(_1055_),
    .B2(net220),
    .A2(_1054_),
    .A1(_0247_));
 sg13g2_a21o_1 _5836_ (.A2(_1053_),
    .A1(_1052_),
    .B1(_1056_),
    .X(_1057_));
 sg13g2_inv_1 _5837_ (.Y(_1058_),
    .A(_3821_));
 sg13g2_and3_1 _5838_ (.X(_1059_),
    .A(net194),
    .B(_1058_),
    .C(_3931_));
 sg13g2_nor3_1 _5839_ (.A(net194),
    .B(_1058_),
    .C(_4125_),
    .Y(_1060_));
 sg13g2_a22oi_1 _5840_ (.Y(_1061_),
    .B1(_1060_),
    .B2(_0827_),
    .A2(_1059_),
    .A1(_0328_));
 sg13g2_buf_1 _5841_ (.A(_1061_),
    .X(_1062_));
 sg13g2_nand3_1 _5842_ (.B(_3692_),
    .C(_4210_),
    .A(net187),
    .Y(_1063_));
 sg13g2_nand4_1 _5843_ (.B(_0564_),
    .C(net183),
    .A(net258),
    .Y(_1064_),
    .D(_0221_));
 sg13g2_nand2_1 _5844_ (.Y(_1065_),
    .A(_1063_),
    .B(_1064_));
 sg13g2_nand3_1 _5845_ (.B(_3822_),
    .C(_0832_),
    .A(net195),
    .Y(_1066_));
 sg13g2_nand4_1 _5846_ (.B(_0830_),
    .C(_0528_),
    .A(net189),
    .Y(_1067_),
    .D(_0330_));
 sg13g2_nand3_1 _5847_ (.B(_3742_),
    .C(_0217_),
    .A(net254),
    .Y(_1068_));
 sg13g2_nand4_1 _5848_ (.B(net303),
    .C(net302),
    .A(_4173_),
    .Y(_1069_),
    .D(_0224_));
 sg13g2_a22oi_1 _5849_ (.Y(_1070_),
    .B1(_1068_),
    .B2(_1069_),
    .A2(_1067_),
    .A1(_1066_));
 sg13g2_nand3b_1 _5850_ (.B(_1065_),
    .C(_1070_),
    .Y(_1071_),
    .A_N(_1062_));
 sg13g2_nor4_1 _5851_ (.A(_1043_),
    .B(_1051_),
    .C(_1057_),
    .D(_1071_),
    .Y(_1072_));
 sg13g2_nor2b_1 _5852_ (.A(_1036_),
    .B_N(_1072_),
    .Y(_1073_));
 sg13g2_a22oi_1 _5853_ (.Y(_1074_),
    .B1(_3884_),
    .B2(_3886_),
    .A2(_3928_),
    .A1(_3793_));
 sg13g2_nand2b_1 _5854_ (.Y(_1075_),
    .B(_3765_),
    .A_N(_1074_));
 sg13g2_o21ai_1 _5855_ (.B1(_1075_),
    .Y(_1076_),
    .A1(_0485_),
    .A2(_3887_));
 sg13g2_a22oi_1 _5856_ (.Y(_1077_),
    .B1(net232),
    .B2(_3843_),
    .A2(net214),
    .A1(net225));
 sg13g2_o21ai_1 _5857_ (.B1(net214),
    .Y(_1078_),
    .A1(net232),
    .A2(net231));
 sg13g2_o21ai_1 _5858_ (.B1(_1078_),
    .Y(_1079_),
    .A1(_4191_),
    .A2(_1077_));
 sg13g2_a21oi_1 _5859_ (.A1(_1047_),
    .A2(_1076_),
    .Y(_1080_),
    .B1(_1079_));
 sg13g2_a22oi_1 _5860_ (.Y(_1081_),
    .B1(net175),
    .B2(net240),
    .A2(net247),
    .A1(net176));
 sg13g2_o21ai_1 _5861_ (.B1(net247),
    .Y(_1082_),
    .A1(net175),
    .A2(net240));
 sg13g2_o21ai_1 _5862_ (.B1(_1082_),
    .Y(_1083_),
    .A1(_0256_),
    .A2(_1081_));
 sg13g2_o21ai_1 _5863_ (.B1(net220),
    .Y(_1084_),
    .A1(net110),
    .A2(net176));
 sg13g2_a22oi_1 _5864_ (.Y(_1085_),
    .B1(net216),
    .B2(net176),
    .A2(net220),
    .A1(net248));
 sg13g2_nand2b_1 _5865_ (.Y(_1086_),
    .B(net255),
    .A_N(_1085_));
 sg13g2_a22oi_1 _5866_ (.Y(_1087_),
    .B1(_1084_),
    .B2(_1086_),
    .A2(_1053_),
    .A1(_1052_));
 sg13g2_a22oi_1 _5867_ (.Y(_1088_),
    .B1(_1048_),
    .B2(_1049_),
    .A2(_1046_),
    .A1(_1044_));
 sg13g2_o21ai_1 _5868_ (.B1(_1088_),
    .Y(_1089_),
    .A1(_1083_),
    .A2(_1087_));
 sg13g2_a21oi_1 _5869_ (.A1(_1080_),
    .A2(_1089_),
    .Y(_1090_),
    .B1(_1043_));
 sg13g2_inv_1 _5870_ (.Y(_1091_),
    .A(_1071_));
 sg13g2_and2_1 _5871_ (.A(_1090_),
    .B(_1091_),
    .X(_1092_));
 sg13g2_nor2_1 _5872_ (.A(_1073_),
    .B(_1092_),
    .Y(_1093_));
 sg13g2_nand3b_1 _5873_ (.B(_4077_),
    .C(_0919_),
    .Y(_1094_),
    .A_N(_3801_));
 sg13g2_nand4_1 _5874_ (.B(_3919_),
    .C(_3801_),
    .A(net172),
    .Y(_1095_),
    .D(_3854_));
 sg13g2_nand3_1 _5875_ (.B(_3702_),
    .C(_0916_),
    .A(_0345_),
    .Y(_1096_));
 sg13g2_nand3_1 _5876_ (.B(_4087_),
    .C(_0416_),
    .A(net172),
    .Y(_1097_));
 sg13g2_a22oi_1 _5877_ (.Y(_1098_),
    .B1(_1096_),
    .B2(_1097_),
    .A2(_1095_),
    .A1(_1094_));
 sg13g2_buf_1 _5878_ (.A(_1098_),
    .X(_1099_));
 sg13g2_nand3_1 _5879_ (.B(_4096_),
    .C(_4098_),
    .A(net156),
    .Y(_1100_));
 sg13g2_inv_1 _5880_ (.Y(_1101_),
    .A(net316));
 sg13g2_nand4_1 _5881_ (.B(_1101_),
    .C(net167),
    .A(net97),
    .Y(_1102_),
    .D(_4100_));
 sg13g2_nand2_2 _5882_ (.Y(_1103_),
    .A(_1100_),
    .B(_1102_));
 sg13g2_nand4_1 _5883_ (.B(_0946_),
    .C(net98),
    .A(net244),
    .Y(_1104_),
    .D(_3695_));
 sg13g2_nor2_1 _5884_ (.A(_3784_),
    .B(_4106_),
    .Y(_1105_));
 sg13g2_nand4_1 _5885_ (.B(net157),
    .C(net156),
    .A(net148),
    .Y(_1106_),
    .D(_1105_));
 sg13g2_nand2_1 _5886_ (.Y(_1107_),
    .A(_1104_),
    .B(_1106_));
 sg13g2_nand3_1 _5887_ (.B(_3848_),
    .C(_4136_),
    .A(_4148_),
    .Y(_1108_));
 sg13g2_nand4_1 _5888_ (.B(_4154_),
    .C(_3847_),
    .A(net245),
    .Y(_1109_),
    .D(_4133_));
 sg13g2_nand4_1 _5889_ (.B(net196),
    .C(net245),
    .A(_4122_),
    .Y(_1110_),
    .D(_4143_));
 sg13g2_nand4_1 _5890_ (.B(net282),
    .C(_4148_),
    .A(_3733_),
    .Y(_1111_),
    .D(_0811_));
 sg13g2_a22oi_1 _5891_ (.Y(_1112_),
    .B1(_1110_),
    .B2(_1111_),
    .A2(_1109_),
    .A1(_1108_));
 sg13g2_buf_1 _5892_ (.A(_1112_),
    .X(_1113_));
 sg13g2_and3_1 _5893_ (.X(_1114_),
    .A(_1103_),
    .B(_1107_),
    .C(_1113_));
 sg13g2_nand2_1 _5894_ (.Y(_1115_),
    .A(_1099_),
    .B(_1114_));
 sg13g2_and2_1 _5895_ (.A(net156),
    .B(_4096_),
    .X(_1116_));
 sg13g2_and2_1 _5896_ (.A(net97),
    .B(net167),
    .X(_1117_));
 sg13g2_a22oi_1 _5897_ (.Y(_1118_),
    .B1(_0604_),
    .B2(net156),
    .A2(net197),
    .A1(net192));
 sg13g2_o21ai_1 _5898_ (.B1(_0615_),
    .Y(_1119_),
    .A1(net157),
    .A2(_0624_));
 sg13g2_o21ai_1 _5899_ (.B1(_1119_),
    .Y(_1120_),
    .A1(_4112_),
    .A2(_1118_));
 sg13g2_o21ai_1 _5900_ (.B1(_1120_),
    .Y(_1121_),
    .A1(_1116_),
    .A2(_1117_));
 sg13g2_o21ai_1 _5901_ (.B1(net167),
    .Y(_1122_),
    .A1(_3944_),
    .A2(_3946_));
 sg13g2_and2_1 _5902_ (.A(net316),
    .B(_0418_),
    .X(_1123_));
 sg13g2_o21ai_1 _5903_ (.B1(net97),
    .Y(_1124_),
    .A1(_4096_),
    .A2(_1123_));
 sg13g2_and2_1 _5904_ (.A(_1122_),
    .B(_1124_),
    .X(_1125_));
 sg13g2_nand2_1 _5905_ (.Y(_1126_),
    .A(_1121_),
    .B(_1125_));
 sg13g2_nand2_1 _5906_ (.Y(_1127_),
    .A(_1066_),
    .B(_1067_));
 sg13g2_nand2_1 _5907_ (.Y(_1128_),
    .A(_1068_),
    .B(_1069_));
 sg13g2_inv_1 _5908_ (.Y(_1129_),
    .A(net185));
 sg13g2_a21oi_1 _5909_ (.A1(net183),
    .A2(_3691_),
    .Y(_1130_),
    .B1(_0822_));
 sg13g2_o21ai_1 _5910_ (.B1(net187),
    .Y(_1131_),
    .A1(_0220_),
    .A2(net188));
 sg13g2_o21ai_1 _5911_ (.B1(_1131_),
    .Y(_1132_),
    .A1(_1129_),
    .A2(_1130_));
 sg13g2_buf_1 _5912_ (.A(_1132_),
    .X(_1133_));
 sg13g2_a22oi_1 _5913_ (.Y(_1134_),
    .B1(net190),
    .B2(net189),
    .A2(net254),
    .A1(_4173_));
 sg13g2_nand2b_1 _5914_ (.Y(_1135_),
    .B(_4165_),
    .A_N(_1134_));
 sg13g2_o21ai_1 _5915_ (.B1(_1135_),
    .Y(_1136_),
    .A1(_0582_),
    .A2(_3742_));
 sg13g2_a21o_1 _5916_ (.A2(_1133_),
    .A1(_1128_),
    .B1(_1136_),
    .X(_1137_));
 sg13g2_a22oi_1 _5917_ (.Y(_1138_),
    .B1(net160),
    .B2(net158),
    .A2(net159),
    .A1(net231));
 sg13g2_o21ai_1 _5918_ (.B1(_0574_),
    .Y(_1139_),
    .A1(net160),
    .A2(_0577_));
 sg13g2_o21ai_1 _5919_ (.B1(_1139_),
    .Y(_1140_),
    .A1(_4192_),
    .A2(_1138_));
 sg13g2_a22oi_1 _5920_ (.Y(_1141_),
    .B1(net259),
    .B2(_3706_),
    .A2(net184),
    .A1(_0577_));
 sg13g2_o21ai_1 _5921_ (.B1(_0213_),
    .Y(_1142_),
    .A1(net259),
    .A2(_3706_));
 sg13g2_o21ai_1 _5922_ (.B1(_1142_),
    .Y(_1143_),
    .A1(_4185_),
    .A2(_1141_));
 sg13g2_a21o_1 _5923_ (.A2(_1140_),
    .A1(_1039_),
    .B1(_1143_),
    .X(_1144_));
 sg13g2_a22oi_1 _5924_ (.Y(_1145_),
    .B1(_1063_),
    .B2(_1064_),
    .A2(_1069_),
    .A1(_1068_));
 sg13g2_and2_1 _5925_ (.A(_1127_),
    .B(_1145_),
    .X(_1146_));
 sg13g2_a22oi_1 _5926_ (.Y(_1147_),
    .B1(net147),
    .B2(net192),
    .A2(_3866_),
    .A1(net245));
 sg13g2_o21ai_1 _5927_ (.B1(net229),
    .Y(_1148_),
    .A1(net147),
    .A2(_4155_));
 sg13g2_o21ai_1 _5928_ (.B1(_1148_),
    .Y(_1149_),
    .A1(_4142_),
    .A2(_1147_));
 sg13g2_buf_1 _5929_ (.A(_1149_),
    .X(_1150_));
 sg13g2_o21ai_1 _5930_ (.B1(net230),
    .Y(_1151_),
    .A1(_0426_),
    .A2(net114));
 sg13g2_a22oi_1 _5931_ (.Y(_1152_),
    .B1(net166),
    .B2(net114),
    .A2(_3864_),
    .A1(_4115_));
 sg13g2_nand2b_1 _5932_ (.Y(_1153_),
    .B(_3734_),
    .A_N(_1152_));
 sg13g2_a22oi_1 _5933_ (.Y(_1154_),
    .B1(_1151_),
    .B2(_1153_),
    .A2(_1109_),
    .A1(_1108_));
 sg13g2_a22oi_1 _5934_ (.Y(_1155_),
    .B1(_0327_),
    .B2(net101),
    .A2(net213),
    .A1(net163));
 sg13g2_nand2b_1 _5935_ (.Y(_1156_),
    .B(net194),
    .A_N(_1155_));
 sg13g2_o21ai_1 _5936_ (.B1(_1156_),
    .Y(_1157_),
    .A1(_0827_),
    .A2(_0328_));
 sg13g2_buf_1 _5937_ (.A(_1157_),
    .X(_1158_));
 sg13g2_a22oi_1 _5938_ (.Y(_1159_),
    .B1(net162),
    .B2(net163),
    .A2(net195),
    .A1(_4170_));
 sg13g2_o21ai_1 _5939_ (.B1(net195),
    .Y(_1160_),
    .A1(_0530_),
    .A2(_0528_));
 sg13g2_o21ai_1 _5940_ (.B1(_1160_),
    .Y(_1161_),
    .A1(_0223_),
    .A2(_1159_));
 sg13g2_or4_1 _5941_ (.A(_1150_),
    .B(_1154_),
    .C(_1158_),
    .D(_1161_),
    .X(_1162_));
 sg13g2_a221oi_1 _5942_ (.B2(_1146_),
    .C1(_1162_),
    .B1(_1144_),
    .A1(_1127_),
    .Y(_1163_),
    .A2(_1137_));
 sg13g2_nand2_1 _5943_ (.Y(_1164_),
    .A(_1108_),
    .B(_1109_));
 sg13g2_o21ai_1 _5944_ (.B1(_1151_),
    .Y(_1165_),
    .A1(_4122_),
    .A2(_1152_));
 sg13g2_nand2b_1 _5945_ (.Y(_1166_),
    .B(_1062_),
    .A_N(_1158_));
 sg13g2_a221oi_1 _5946_ (.B2(_1166_),
    .C1(_1150_),
    .B1(_1113_),
    .A1(_1164_),
    .Y(_1167_),
    .A2(_1165_));
 sg13g2_nor2_1 _5947_ (.A(_1163_),
    .B(_1167_),
    .Y(_1168_));
 sg13g2_and3_1 _5948_ (.X(_1169_),
    .A(_1099_),
    .B(_1103_),
    .C(_1107_));
 sg13g2_a22oi_1 _5949_ (.Y(_1170_),
    .B1(_1168_),
    .B2(_1169_),
    .A2(_1126_),
    .A1(_1099_));
 sg13g2_o21ai_1 _5950_ (.B1(_1170_),
    .Y(_1171_),
    .A1(_1093_),
    .A2(_1115_));
 sg13g2_a22oi_1 _5951_ (.Y(_1172_),
    .B1(net155),
    .B2(_0347_),
    .A2(net111),
    .A1(_3946_));
 sg13g2_o21ai_1 _5952_ (.B1(net111),
    .Y(_1173_),
    .A1(net155),
    .A2(net172));
 sg13g2_o21ai_1 _5953_ (.B1(_1173_),
    .Y(_1174_),
    .A1(_4094_),
    .A2(_1172_));
 sg13g2_nand2_1 _5954_ (.Y(_1175_),
    .A(_1094_),
    .B(_1095_));
 sg13g2_a22oi_1 _5955_ (.Y(_1176_),
    .B1(net218),
    .B2(_0669_),
    .A2(net171),
    .A1(net172));
 sg13g2_o21ai_1 _5956_ (.B1(_0355_),
    .Y(_1177_),
    .A1(net218),
    .A2(_0669_));
 sg13g2_o21ai_1 _5957_ (.B1(_1177_),
    .Y(_1178_),
    .A1(_4086_),
    .A2(_1176_));
 sg13g2_a21oi_1 _5958_ (.A1(_1174_),
    .A2(_1175_),
    .Y(_1179_),
    .B1(_1178_));
 sg13g2_nand2b_1 _5959_ (.Y(_1180_),
    .B(_1179_),
    .A_N(_1171_));
 sg13g2_nand2b_1 _5960_ (.Y(_1181_),
    .B(_1180_),
    .A_N(_0996_));
 sg13g2_nand2_1 _5961_ (.Y(_1182_),
    .A(_0983_),
    .B(_0984_));
 sg13g2_inv_1 _5962_ (.Y(_1183_),
    .A(net199));
 sg13g2_o21ai_1 _5963_ (.B1(_3817_),
    .Y(_1184_),
    .A1(_0678_),
    .A2(net168));
 sg13g2_nor2_1 _5964_ (.A(net168),
    .B(_0987_),
    .Y(_1185_));
 sg13g2_a21oi_1 _5965_ (.A1(_1183_),
    .A2(_1184_),
    .Y(_1186_),
    .B1(_1185_));
 sg13g2_a21oi_2 _5966_ (.B1(_0972_),
    .Y(_1187_),
    .A2(_1186_),
    .A1(_1182_));
 sg13g2_a21oi_1 _5967_ (.A1(_0990_),
    .A2(_1181_),
    .Y(_1188_),
    .B1(_1187_));
 sg13g2_xnor2_1 _5968_ (.Y(_1189_),
    .A(_0969_),
    .B(_1188_));
 sg13g2_inv_1 _5969_ (.Y(_1190_),
    .A(_3743_));
 sg13g2_o21ai_1 _5970_ (.B1(net80),
    .Y(_1191_),
    .A1(net39),
    .A2(_1190_));
 sg13g2_a21oi_1 _5971_ (.A1(net41),
    .A2(_1189_),
    .Y(_1192_),
    .B1(_1191_));
 sg13g2_inv_1 _5972_ (.Y(_1193_),
    .A(\collatz.iter[103] ));
 sg13g2_buf_1 _5973_ (.A(ui_in[7]),
    .X(_1194_));
 sg13g2_nand2_1 _5974_ (.Y(_1195_),
    .A(net324),
    .B(_0391_));
 sg13g2_o21ai_1 _5975_ (.B1(_1195_),
    .Y(_1196_),
    .A1(_1193_),
    .A2(net20));
 sg13g2_o21ai_1 _5976_ (.B1(net270),
    .Y(_1197_),
    .A1(net82),
    .A2(_1196_));
 sg13g2_nor2_1 _5977_ (.A(_1192_),
    .B(_1197_),
    .Y(_0032_));
 sg13g2_buf_1 _5978_ (.A(net78),
    .X(_1198_));
 sg13g2_buf_1 _5979_ (.A(net51),
    .X(_1199_));
 sg13g2_nand2_1 _5980_ (.Y(_1200_),
    .A(_0362_),
    .B(_0365_));
 sg13g2_inv_1 _5981_ (.Y(_1201_),
    .A(_0360_));
 sg13g2_a21oi_1 _5982_ (.A1(_4066_),
    .A2(_1200_),
    .Y(_1202_),
    .B1(_1201_));
 sg13g2_inv_1 _5983_ (.Y(_1203_),
    .A(_0356_));
 sg13g2_a21oi_1 _5984_ (.A1(_4083_),
    .A2(_0350_),
    .Y(_1204_),
    .B1(_1203_));
 sg13g2_a21oi_1 _5985_ (.A1(_4099_),
    .A2(_4101_),
    .Y(_1205_),
    .B1(_4107_));
 sg13g2_a22oi_1 _5986_ (.Y(_1206_),
    .B1(_4088_),
    .B2(_4092_),
    .A2(_4082_),
    .A1(_4079_));
 sg13g2_o21ai_1 _5987_ (.B1(_1206_),
    .Y(_1207_),
    .A1(_0344_),
    .A2(_1205_));
 sg13g2_nand2_1 _5988_ (.Y(_1208_),
    .A(_4066_),
    .B(_4075_));
 sg13g2_a21o_1 _5989_ (.A2(_1207_),
    .A1(_1204_),
    .B1(_1208_),
    .X(_1209_));
 sg13g2_nor4_1 _5990_ (.A(_3788_),
    .B(_3920_),
    .C(_0397_),
    .D(_0708_),
    .Y(_1210_));
 sg13g2_nor4_1 _5991_ (.A(_0701_),
    .B(_3696_),
    .C(_1193_),
    .D(_3697_),
    .Y(_1211_));
 sg13g2_a22oi_1 _5992_ (.Y(_1212_),
    .B1(_1211_),
    .B2(net242),
    .A2(_1210_),
    .A1(_1193_));
 sg13g2_buf_2 _5993_ (.A(_1212_),
    .X(_1213_));
 sg13g2_a221oi_1 _5994_ (.B2(_1209_),
    .C1(_1213_),
    .B1(_1202_),
    .A1(_4054_),
    .Y(_1214_),
    .A2(_4057_));
 sg13g2_a21o_1 _5995_ (.A2(net200),
    .A1(_3788_),
    .B1(_3447_),
    .X(_1215_));
 sg13g2_a21o_1 _5996_ (.A2(net321),
    .A1(net200),
    .B1(_3697_),
    .X(_1216_));
 sg13g2_a22oi_1 _5997_ (.Y(_1217_),
    .B1(_1216_),
    .B2(net217),
    .A2(_1215_),
    .A1(net150));
 sg13g2_o21ai_1 _5998_ (.B1(_1217_),
    .Y(_1218_),
    .A1(_0376_),
    .A2(_1213_));
 sg13g2_nor2_1 _5999_ (.A(_4163_),
    .B(_0338_),
    .Y(_1219_));
 sg13g2_nand4_1 _6000_ (.B(_4066_),
    .C(_4075_),
    .A(_4058_),
    .Y(_1220_),
    .D(_4083_));
 sg13g2_or2_1 _6001_ (.X(_1221_),
    .B(_4103_),
    .A(_1220_));
 sg13g2_buf_1 _6002_ (.A(_1221_),
    .X(_1222_));
 sg13g2_nor3_1 _6003_ (.A(_1219_),
    .B(_1222_),
    .C(_1213_),
    .Y(_1223_));
 sg13g2_or3_1 _6004_ (.A(_1214_),
    .B(_1218_),
    .C(_1223_),
    .X(_1224_));
 sg13g2_buf_1 _6005_ (.A(_3743_),
    .X(_1225_));
 sg13g2_xor2_1 _6006_ (.B(_1225_),
    .A(net146),
    .X(_1226_));
 sg13g2_xnor2_1 _6007_ (.Y(_1227_),
    .A(_1224_),
    .B(_1226_));
 sg13g2_buf_1 _6008_ (.A(_0692_),
    .X(_1228_));
 sg13g2_buf_1 _6009_ (.A(_3456_),
    .X(_1229_));
 sg13g2_nor2_1 _6010_ (.A(net36),
    .B(net144),
    .Y(_1230_));
 sg13g2_a21oi_1 _6011_ (.A1(net37),
    .A2(_1227_),
    .Y(_1231_),
    .B1(_1230_));
 sg13g2_nand2_1 _6012_ (.Y(_1232_),
    .A(_1198_),
    .B(_1231_));
 sg13g2_and2_1 _6013_ (.A(net1),
    .B(net83),
    .X(_1233_));
 sg13g2_buf_2 _6014_ (.A(_1233_),
    .X(_1234_));
 sg13g2_nand3_1 _6015_ (.B(_0383_),
    .C(net272),
    .A(_3978_),
    .Y(_1235_));
 sg13g2_nand2_1 _6016_ (.Y(_1236_),
    .A(net109),
    .B(_0389_));
 sg13g2_buf_2 _6017_ (.A(_1236_),
    .X(_1237_));
 sg13g2_nor2_1 _6018_ (.A(_1235_),
    .B(_1237_),
    .Y(_1238_));
 sg13g2_buf_2 _6019_ (.A(_1238_),
    .X(_1239_));
 sg13g2_nand2_1 _6020_ (.Y(_1240_),
    .A(_0383_),
    .B(net272));
 sg13g2_nor2_1 _6021_ (.A(_3979_),
    .B(_1240_),
    .Y(_1241_));
 sg13g2_a21oi_1 _6022_ (.A1(net66),
    .A2(_1241_),
    .Y(_1242_),
    .B1(net203));
 sg13g2_buf_2 _6023_ (.A(_1242_),
    .X(_1243_));
 sg13g2_a22oi_1 _6024_ (.Y(_1244_),
    .B1(_1243_),
    .B2(net145),
    .A2(_1239_),
    .A1(_1234_));
 sg13g2_a21oi_1 _6025_ (.A1(_1232_),
    .A2(_1244_),
    .Y(_0033_),
    .B1(_3965_));
 sg13g2_and2_1 _6026_ (.A(_3697_),
    .B(_3743_),
    .X(_1245_));
 sg13g2_buf_2 _6027_ (.A(_1245_),
    .X(_1246_));
 sg13g2_a21o_1 _6028_ (.A2(_0688_),
    .A1(net146),
    .B1(_1246_),
    .X(_1247_));
 sg13g2_and2_1 _6029_ (.A(_0688_),
    .B(_1246_),
    .X(_1248_));
 sg13g2_o21ai_1 _6030_ (.B1(net321),
    .Y(_1249_),
    .A1(net150),
    .A2(net145));
 sg13g2_nand3_1 _6031_ (.B(net200),
    .C(_0964_),
    .A(net217),
    .Y(_1250_));
 sg13g2_nand2_1 _6032_ (.Y(_1251_),
    .A(_1249_),
    .B(_1250_));
 sg13g2_a221oi_1 _6033_ (.B2(net200),
    .C1(_1251_),
    .B1(_1248_),
    .A1(net217),
    .Y(_1252_),
    .A2(_1247_));
 sg13g2_buf_1 _6034_ (.A(_1252_),
    .X(_1253_));
 sg13g2_nand2_1 _6035_ (.Y(_1254_),
    .A(_0532_),
    .B(_0534_));
 sg13g2_and3_1 _6036_ (.X(_1255_),
    .A(_1254_),
    .B(_0542_),
    .C(_0551_));
 sg13g2_nand2_1 _6037_ (.Y(_1256_),
    .A(_0511_),
    .B(_0557_));
 sg13g2_and2_1 _6038_ (.A(_0318_),
    .B(_0496_),
    .X(_1257_));
 sg13g2_a22oi_1 _6039_ (.Y(_1258_),
    .B1(net291),
    .B2(_3826_),
    .A2(net241),
    .A1(net216));
 sg13g2_o21ai_1 _6040_ (.B1(_0442_),
    .Y(_1259_),
    .A1(_0770_),
    .A2(_1258_));
 sg13g2_o21ai_1 _6041_ (.B1(_1259_),
    .Y(_1260_),
    .A1(_0497_),
    .A2(_1257_));
 sg13g2_and3_1 _6042_ (.X(_1261_),
    .A(_0494_),
    .B(_0498_),
    .C(_1260_));
 sg13g2_a21oi_1 _6043_ (.A1(_0489_),
    .A2(_0557_),
    .Y(_1262_),
    .B1(_0573_));
 sg13g2_o21ai_1 _6044_ (.B1(_1262_),
    .Y(_1263_),
    .A1(_1256_),
    .A2(_1261_));
 sg13g2_a21oi_1 _6045_ (.A1(_0503_),
    .A2(_0519_),
    .Y(_1264_),
    .B1(_0444_));
 sg13g2_a22oi_1 _6046_ (.Y(_1265_),
    .B1(_0514_),
    .B2(_0518_),
    .A2(_0452_),
    .A1(_0449_));
 sg13g2_nand3_1 _6047_ (.B(_0464_),
    .C(_1265_),
    .A(_0460_),
    .Y(_1266_));
 sg13g2_nand4_1 _6048_ (.B(_0480_),
    .C(_0483_),
    .A(_0474_),
    .Y(_1267_),
    .D(_1265_));
 sg13g2_nand3_1 _6049_ (.B(_1266_),
    .C(_1267_),
    .A(_1264_),
    .Y(_1268_));
 sg13g2_nand3_1 _6050_ (.B(_0542_),
    .C(_0551_),
    .A(_1254_),
    .Y(_1269_));
 sg13g2_nand2b_1 _6051_ (.Y(_1270_),
    .B(_0522_),
    .A_N(_0509_));
 sg13g2_nor3_1 _6052_ (.A(_1269_),
    .B(_1256_),
    .C(_1270_),
    .Y(_1271_));
 sg13g2_nand2_1 _6053_ (.Y(_1272_),
    .A(_0547_),
    .B(_0549_));
 sg13g2_a21oi_1 _6054_ (.A1(_0579_),
    .A2(_1272_),
    .Y(_1273_),
    .B1(_0563_));
 sg13g2_nand2_1 _6055_ (.Y(_1274_),
    .A(_1254_),
    .B(_0559_));
 sg13g2_a21oi_1 _6056_ (.A1(_1254_),
    .A2(_0567_),
    .Y(_1275_),
    .B1(_0585_));
 sg13g2_o21ai_1 _6057_ (.B1(_1275_),
    .Y(_1276_),
    .A1(_1273_),
    .A2(_1274_));
 sg13g2_a221oi_1 _6058_ (.B2(_1271_),
    .C1(_1276_),
    .B1(_1268_),
    .A1(_1255_),
    .Y(_1277_),
    .A2(_1263_));
 sg13g2_buf_1 _6059_ (.A(_1277_),
    .X(_1278_));
 sg13g2_nand2_1 _6060_ (.Y(_1279_),
    .A(_0595_),
    .B(_0596_));
 sg13g2_nand2_1 _6061_ (.Y(_1280_),
    .A(_0417_),
    .B(_0419_));
 sg13g2_nand2b_1 _6062_ (.Y(_1281_),
    .B(_1280_),
    .A_N(_0633_));
 sg13g2_nand2_1 _6063_ (.Y(_1282_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_inv_1 _6064_ (.Y(_1283_),
    .A(_1282_));
 sg13g2_nor3_1 _6065_ (.A(_1281_),
    .B(_0609_),
    .C(_1283_),
    .Y(_1284_));
 sg13g2_and2_1 _6066_ (.A(_0425_),
    .B(_0613_),
    .X(_1285_));
 sg13g2_buf_1 _6067_ (.A(_1285_),
    .X(_1286_));
 sg13g2_nand4_1 _6068_ (.B(_1279_),
    .C(_1284_),
    .A(_0586_),
    .Y(_1287_),
    .D(_1286_));
 sg13g2_a21oi_1 _6069_ (.A1(net96),
    .A2(net97),
    .Y(_1288_),
    .B1(_0606_));
 sg13g2_o21ai_1 _6070_ (.B1(_0625_),
    .Y(_1289_),
    .A1(_0895_),
    .A2(_1288_));
 sg13g2_nand2_1 _6071_ (.Y(_1290_),
    .A(_0635_),
    .B(_0636_));
 sg13g2_a21oi_1 _6072_ (.A1(_1280_),
    .A2(_1289_),
    .Y(_1291_),
    .B1(_1290_));
 sg13g2_o21ai_1 _6073_ (.B1(_0641_),
    .Y(_1292_),
    .A1(_0633_),
    .A2(_1291_));
 sg13g2_and2_1 _6074_ (.A(_3770_),
    .B(_0587_),
    .X(_1293_));
 sg13g2_nor2_1 _6075_ (.A(_0830_),
    .B(_0588_),
    .Y(_1294_));
 sg13g2_nand2_1 _6076_ (.Y(_1295_),
    .A(_0594_),
    .B(_0587_));
 sg13g2_nand2_1 _6077_ (.Y(_1296_),
    .A(net101),
    .B(net166));
 sg13g2_a22oi_1 _6078_ (.Y(_1297_),
    .B1(_1296_),
    .B2(_4122_),
    .A2(_0811_),
    .A1(_0827_));
 sg13g2_o21ai_1 _6079_ (.B1(_1297_),
    .Y(_1298_),
    .A1(_1294_),
    .A2(_1295_));
 sg13g2_a221oi_1 _6080_ (.B2(_1293_),
    .C1(_1298_),
    .B1(_0589_),
    .A1(_4117_),
    .Y(_1299_),
    .A2(_0594_));
 sg13g2_nand2_1 _6081_ (.Y(_1300_),
    .A(net193),
    .B(_4112_));
 sg13g2_o21ai_1 _6082_ (.B1(_1300_),
    .Y(_1301_),
    .A1(_0899_),
    .A2(_0602_));
 sg13g2_o21ai_1 _6083_ (.B1(_0899_),
    .Y(_1302_),
    .A1(net244),
    .A2(_0602_));
 sg13g2_a21oi_1 _6084_ (.A1(net148),
    .A2(net96),
    .Y(_1303_),
    .B1(net244));
 sg13g2_a221oi_1 _6085_ (.B2(net193),
    .C1(_1303_),
    .B1(_1302_),
    .A1(_0947_),
    .Y(_1304_),
    .A2(_1301_));
 sg13g2_a21o_1 _6086_ (.A2(_1299_),
    .A1(_1286_),
    .B1(_1304_),
    .X(_1305_));
 sg13g2_a221oi_1 _6087_ (.B2(_1305_),
    .C1(_0672_),
    .B1(_1284_),
    .A1(_1282_),
    .Y(_1306_),
    .A2(_1292_));
 sg13g2_o21ai_1 _6088_ (.B1(_1306_),
    .Y(_1307_),
    .A1(_1278_),
    .A2(_1287_));
 sg13g2_buf_2 _6089_ (.A(_1307_),
    .X(_1308_));
 sg13g2_a221oi_1 _6090_ (.B2(_1308_),
    .C1(_0682_),
    .B1(_0655_),
    .A1(_0666_),
    .Y(_1309_),
    .A2(_0676_));
 sg13g2_buf_2 _6091_ (.A(_1309_),
    .X(_1310_));
 sg13g2_nand3b_1 _6092_ (.B(_0407_),
    .C(_1246_),
    .Y(_1311_),
    .A_N(net321));
 sg13g2_nor2_1 _6093_ (.A(_3697_),
    .B(_3743_),
    .Y(_1312_));
 sg13g2_nand3_1 _6094_ (.B(_0408_),
    .C(_1312_),
    .A(net321),
    .Y(_1313_));
 sg13g2_a22oi_1 _6095_ (.Y(_1314_),
    .B1(_1311_),
    .B2(_1313_),
    .A2(_0658_),
    .A1(_0656_));
 sg13g2_nand2b_1 _6096_ (.Y(_1315_),
    .B(_1314_),
    .A_N(_1310_));
 sg13g2_and2_1 _6097_ (.A(_1253_),
    .B(_1315_),
    .X(_1316_));
 sg13g2_xnor2_1 _6098_ (.Y(_1317_),
    .A(net144),
    .B(net145));
 sg13g2_xnor2_1 _6099_ (.Y(_1318_),
    .A(_1316_),
    .B(_1317_));
 sg13g2_buf_1 _6100_ (.A(net301),
    .X(_1319_));
 sg13g2_nor2_1 _6101_ (.A(net36),
    .B(net143),
    .Y(_1320_));
 sg13g2_a21oi_1 _6102_ (.A1(net37),
    .A2(_1318_),
    .Y(_1321_),
    .B1(_1320_));
 sg13g2_nand2_1 _6103_ (.Y(_1322_),
    .A(net64),
    .B(_1321_));
 sg13g2_and2_1 _6104_ (.A(_3973_),
    .B(net83),
    .X(_1323_));
 sg13g2_buf_2 _6105_ (.A(_1323_),
    .X(_1324_));
 sg13g2_a22oi_1 _6106_ (.Y(_1325_),
    .B1(_1324_),
    .B2(_1239_),
    .A2(_1243_),
    .A1(net144));
 sg13g2_buf_1 _6107_ (.A(net204),
    .X(_1326_));
 sg13g2_a21oi_1 _6108_ (.A1(_1322_),
    .A2(_1325_),
    .Y(_0034_),
    .B1(net94));
 sg13g2_and2_1 _6109_ (.A(net321),
    .B(_3456_),
    .X(_1327_));
 sg13g2_buf_1 _6110_ (.A(_1327_),
    .X(_1328_));
 sg13g2_nand3_1 _6111_ (.B(_1312_),
    .C(_1328_),
    .A(net217),
    .Y(_1329_));
 sg13g2_buf_1 _6112_ (.A(_1329_),
    .X(_1330_));
 sg13g2_nand3_1 _6113_ (.B(_3464_),
    .C(_1246_),
    .A(_0701_),
    .Y(_1331_));
 sg13g2_buf_1 _6114_ (.A(_1331_),
    .X(_1332_));
 sg13g2_nand2_1 _6115_ (.Y(_1333_),
    .A(_1330_),
    .B(_1332_));
 sg13g2_a21o_1 _6116_ (.A2(net150),
    .A1(net217),
    .B1(_3456_),
    .X(_1334_));
 sg13g2_nand2_1 _6117_ (.Y(_1335_),
    .A(net145),
    .B(_1334_));
 sg13g2_a21o_1 _6118_ (.A2(_3456_),
    .A1(net150),
    .B1(net145),
    .X(_1336_));
 sg13g2_nand2_1 _6119_ (.Y(_1337_),
    .A(net146),
    .B(_1336_));
 sg13g2_nand2_1 _6120_ (.Y(_1338_),
    .A(_1335_),
    .B(_1337_));
 sg13g2_a21oi_1 _6121_ (.A1(_0962_),
    .A2(_1333_),
    .Y(_1339_),
    .B1(_1338_));
 sg13g2_xnor2_1 _6122_ (.Y(_1340_),
    .A(net144),
    .B(net143));
 sg13g2_xnor2_1 _6123_ (.Y(_1341_),
    .A(_1339_),
    .B(_1340_));
 sg13g2_buf_1 _6124_ (.A(_3566_),
    .X(_1342_));
 sg13g2_nor2_1 _6125_ (.A(net36),
    .B(_1342_),
    .Y(_1343_));
 sg13g2_a21oi_1 _6126_ (.A1(net37),
    .A2(_1341_),
    .Y(_1344_),
    .B1(_1343_));
 sg13g2_nand2_1 _6127_ (.Y(_1345_),
    .A(net64),
    .B(_1344_));
 sg13g2_buf_1 _6128_ (.A(ui_in[2]),
    .X(_1346_));
 sg13g2_and2_1 _6129_ (.A(_1346_),
    .B(net83),
    .X(_1347_));
 sg13g2_buf_2 _6130_ (.A(_1347_),
    .X(_1348_));
 sg13g2_a22oi_1 _6131_ (.Y(_1349_),
    .B1(_1348_),
    .B2(_1239_),
    .A2(_1243_),
    .A1(net143));
 sg13g2_a21oi_1 _6132_ (.A1(_1345_),
    .A2(_1349_),
    .Y(_0035_),
    .B1(_1326_));
 sg13g2_nand2_1 _6133_ (.Y(_1350_),
    .A(_1107_),
    .B(_1164_));
 sg13g2_nand2_1 _6134_ (.Y(_1351_),
    .A(_1110_),
    .B(_1111_));
 sg13g2_inv_1 _6135_ (.Y(_1352_),
    .A(_1062_));
 sg13g2_nand2_1 _6136_ (.Y(_1353_),
    .A(_1351_),
    .B(_1352_));
 sg13g2_nor2_1 _6137_ (.A(_1350_),
    .B(_1353_),
    .Y(_1354_));
 sg13g2_nand2_1 _6138_ (.Y(_1355_),
    .A(_1052_),
    .B(_1053_));
 sg13g2_nand2_1 _6139_ (.Y(_1356_),
    .A(_1050_),
    .B(_1355_));
 sg13g2_or2_1 _6140_ (.X(_1357_),
    .B(_1356_),
    .A(_1056_));
 sg13g2_or2_1 _6141_ (.X(_1358_),
    .B(_1087_),
    .A(_1083_));
 sg13g2_a21oi_1 _6142_ (.A1(_1050_),
    .A2(_1358_),
    .Y(_1359_),
    .B1(_1076_));
 sg13g2_o21ai_1 _6143_ (.B1(_1359_),
    .Y(_1360_),
    .A1(_1036_),
    .A2(_1357_));
 sg13g2_inv_1 _6144_ (.Y(_1361_),
    .A(_1047_));
 sg13g2_nand2_1 _6145_ (.Y(_1362_),
    .A(_1065_),
    .B(_1070_));
 sg13g2_nor3_1 _6146_ (.A(_1043_),
    .B(_1361_),
    .C(_1362_),
    .Y(_1363_));
 sg13g2_a21o_1 _6147_ (.A2(_1079_),
    .A1(_1042_),
    .B1(_1140_),
    .X(_1364_));
 sg13g2_or2_1 _6148_ (.X(_1365_),
    .B(_1143_),
    .A(_1133_));
 sg13g2_a21oi_1 _6149_ (.A1(_1039_),
    .A2(_1364_),
    .Y(_1366_),
    .B1(_1365_));
 sg13g2_o21ai_1 _6150_ (.B1(_1070_),
    .Y(_1367_),
    .A1(_1133_),
    .A2(_1065_));
 sg13g2_a21oi_1 _6151_ (.A1(_1127_),
    .A2(_1136_),
    .Y(_1368_),
    .B1(_1161_));
 sg13g2_o21ai_1 _6152_ (.B1(_1368_),
    .Y(_1369_),
    .A1(_1366_),
    .A2(_1367_));
 sg13g2_a21o_1 _6153_ (.A2(_1363_),
    .A1(_1360_),
    .B1(_1369_),
    .X(_1370_));
 sg13g2_a21oi_1 _6154_ (.A1(_1351_),
    .A2(_1158_),
    .Y(_1371_),
    .B1(_1165_));
 sg13g2_a21oi_1 _6155_ (.A1(_1107_),
    .A2(_1150_),
    .Y(_1372_),
    .B1(_1120_));
 sg13g2_o21ai_1 _6156_ (.B1(_1372_),
    .Y(_1373_),
    .A1(_1350_),
    .A2(_1371_));
 sg13g2_a21o_1 _6157_ (.A2(_1370_),
    .A1(_1354_),
    .B1(_1373_),
    .X(_1374_));
 sg13g2_buf_1 _6158_ (.A(_1374_),
    .X(_1375_));
 sg13g2_and2_1 _6159_ (.A(_3743_),
    .B(_3744_),
    .X(_1376_));
 sg13g2_buf_1 _6160_ (.A(_1376_),
    .X(_1377_));
 sg13g2_nand3_1 _6161_ (.B(_3464_),
    .C(_1377_),
    .A(net150),
    .Y(_1378_));
 sg13g2_nand3_1 _6162_ (.B(_3745_),
    .C(_1328_),
    .A(_0708_),
    .Y(_1379_));
 sg13g2_nand2_1 _6163_ (.Y(_1380_),
    .A(_1378_),
    .B(_1379_));
 sg13g2_nand2_1 _6164_ (.Y(_1381_),
    .A(_1182_),
    .B(_1380_));
 sg13g2_nand4_1 _6165_ (.B(_0644_),
    .C(_0369_),
    .A(net296),
    .Y(_1382_),
    .D(_4063_));
 sg13g2_nand3_1 _6166_ (.B(_3777_),
    .C(_0987_),
    .A(_3721_),
    .Y(_1383_));
 sg13g2_nand2_1 _6167_ (.Y(_1384_),
    .A(_1382_),
    .B(_1383_));
 sg13g2_nand2_1 _6168_ (.Y(_1385_),
    .A(_0991_),
    .B(_1384_));
 sg13g2_nand3_1 _6169_ (.B(_1103_),
    .C(_0995_),
    .A(_1099_),
    .Y(_1386_));
 sg13g2_nor3_2 _6170_ (.A(_1381_),
    .B(_1385_),
    .C(_1386_),
    .Y(_1387_));
 sg13g2_nor2_1 _6171_ (.A(_3817_),
    .B(_0976_),
    .Y(_1388_));
 sg13g2_inv_1 _6172_ (.Y(_1389_),
    .A(_0678_));
 sg13g2_o21ai_1 _6173_ (.B1(_1389_),
    .Y(_1390_),
    .A1(_3777_),
    .A2(_1388_));
 sg13g2_o21ai_1 _6174_ (.B1(_3817_),
    .Y(_1391_),
    .A1(net168),
    .A2(_0976_));
 sg13g2_a21oi_1 _6175_ (.A1(_1183_),
    .A2(_1391_),
    .Y(_1392_),
    .B1(_1185_));
 sg13g2_a22oi_1 _6176_ (.Y(_1393_),
    .B1(_1382_),
    .B2(_1383_),
    .A2(_0978_),
    .A1(_0977_));
 sg13g2_nand2_1 _6177_ (.Y(_1394_),
    .A(_1096_),
    .B(_1097_));
 sg13g2_nand2_1 _6178_ (.Y(_1395_),
    .A(_1122_),
    .B(_1124_));
 sg13g2_a21oi_1 _6179_ (.A1(_1394_),
    .A2(_1395_),
    .Y(_1396_),
    .B1(_1174_));
 sg13g2_nand2_1 _6180_ (.Y(_1397_),
    .A(_1175_),
    .B(_0995_));
 sg13g2_nand2_1 _6181_ (.Y(_1398_),
    .A(_0980_),
    .B(_0981_));
 sg13g2_a21oi_1 _6182_ (.A1(_1178_),
    .A2(_0995_),
    .Y(_1399_),
    .B1(_1398_));
 sg13g2_o21ai_1 _6183_ (.B1(_1399_),
    .Y(_1400_),
    .A1(_1396_),
    .A2(_1397_));
 sg13g2_a22oi_1 _6184_ (.Y(_1401_),
    .B1(_1393_),
    .B2(_1400_),
    .A2(_1392_),
    .A1(_1390_));
 sg13g2_nor2_1 _6185_ (.A(_0701_),
    .B(_3698_),
    .Y(_1402_));
 sg13g2_nand2_1 _6186_ (.Y(_1403_),
    .A(_3743_),
    .B(net301));
 sg13g2_a21oi_1 _6187_ (.A1(net242),
    .A2(_0970_),
    .Y(_1404_),
    .B1(net217));
 sg13g2_nand2_1 _6188_ (.Y(_1405_),
    .A(_0964_),
    .B(_1229_));
 sg13g2_o21ai_1 _6189_ (.B1(_1405_),
    .Y(_1406_),
    .A1(_1403_),
    .A2(_1404_));
 sg13g2_o21ai_1 _6190_ (.B1(_0708_),
    .Y(_1407_),
    .A1(_0971_),
    .A2(_1405_));
 sg13g2_o21ai_1 _6191_ (.B1(_1229_),
    .Y(_1408_),
    .A1(net145),
    .A2(net143));
 sg13g2_nand2_1 _6192_ (.Y(_1409_),
    .A(net321),
    .B(_1377_));
 sg13g2_nand2_1 _6193_ (.Y(_1410_),
    .A(_1408_),
    .B(_1409_));
 sg13g2_a221oi_1 _6194_ (.B2(_1407_),
    .C1(_1410_),
    .B1(_1406_),
    .A1(_1402_),
    .Y(_1411_),
    .A2(_1328_));
 sg13g2_o21ai_1 _6195_ (.B1(_1411_),
    .Y(_1412_),
    .A1(_1381_),
    .A2(_1401_));
 sg13g2_a21oi_2 _6196_ (.B1(_1412_),
    .Y(_1413_),
    .A2(_1387_),
    .A1(_1375_));
 sg13g2_xnor2_1 _6197_ (.Y(_1414_),
    .A(net142),
    .B(net143));
 sg13g2_xnor2_1 _6198_ (.Y(_1415_),
    .A(_1413_),
    .B(_1414_));
 sg13g2_buf_1 _6199_ (.A(_0692_),
    .X(_1416_));
 sg13g2_buf_1 _6200_ (.A(net286),
    .X(_1417_));
 sg13g2_nor2_1 _6201_ (.A(net35),
    .B(net141),
    .Y(_1418_));
 sg13g2_a21oi_1 _6202_ (.A1(net37),
    .A2(_1415_),
    .Y(_1419_),
    .B1(_1418_));
 sg13g2_nand2_1 _6203_ (.Y(_1420_),
    .A(net64),
    .B(_1419_));
 sg13g2_and2_1 _6204_ (.A(net2),
    .B(_3985_),
    .X(_1421_));
 sg13g2_buf_2 _6205_ (.A(_1421_),
    .X(_1422_));
 sg13g2_a22oi_1 _6206_ (.Y(_1423_),
    .B1(_1422_),
    .B2(_1239_),
    .A2(_1243_),
    .A1(net142));
 sg13g2_a21oi_1 _6207_ (.A1(_1420_),
    .A2(_1423_),
    .Y(_0036_),
    .B1(net94));
 sg13g2_inv_1 _6208_ (.Y(_1424_),
    .A(_3577_));
 sg13g2_nor2_1 _6209_ (.A(_1217_),
    .B(_1403_),
    .Y(_1425_));
 sg13g2_a21oi_1 _6210_ (.A1(net145),
    .A2(net142),
    .Y(_1426_),
    .B1(_1319_));
 sg13g2_nor2b_1 _6211_ (.A(_1426_),
    .B_N(net144),
    .Y(_1427_));
 sg13g2_and2_1 _6212_ (.A(net142),
    .B(net143),
    .X(_1428_));
 sg13g2_nand2_1 _6213_ (.Y(_1429_),
    .A(net142),
    .B(_1328_));
 sg13g2_o21ai_1 _6214_ (.B1(_1409_),
    .Y(_1430_),
    .A1(_1217_),
    .A2(_1429_));
 sg13g2_nor4_2 _6215_ (.A(_1425_),
    .B(_1427_),
    .C(_1428_),
    .Y(_1431_),
    .D(_1430_));
 sg13g2_nand2b_1 _6216_ (.Y(_1432_),
    .B(_0375_),
    .A_N(_0372_));
 sg13g2_nor2_1 _6217_ (.A(_3566_),
    .B(_1403_),
    .Y(_1433_));
 sg13g2_nor2b_1 _6218_ (.A(net301),
    .B_N(_3566_),
    .Y(_1434_));
 sg13g2_and2_1 _6219_ (.A(_1190_),
    .B(_1434_),
    .X(_1435_));
 sg13g2_a22oi_1 _6220_ (.Y(_1436_),
    .B1(_1435_),
    .B2(_1328_),
    .A2(_1433_),
    .A1(_3464_));
 sg13g2_nor2_2 _6221_ (.A(_1213_),
    .B(_1436_),
    .Y(_1437_));
 sg13g2_o21ai_1 _6222_ (.B1(_1437_),
    .Y(_1438_),
    .A1(_1432_),
    .A2(_0368_));
 sg13g2_nand3b_1 _6223_ (.B(_1437_),
    .C(_4085_),
    .Y(_1439_),
    .A_N(_0351_));
 sg13g2_and3_1 _6224_ (.X(_1440_),
    .A(_1431_),
    .B(_1438_),
    .C(_1439_));
 sg13g2_nand2_1 _6225_ (.Y(_1441_),
    .A(_4114_),
    .B(_4138_));
 sg13g2_a21o_1 _6226_ (.A2(net299),
    .A1(_3641_),
    .B1(net252),
    .X(_1442_));
 sg13g2_a22oi_1 _6227_ (.Y(_1443_),
    .B1(_4128_),
    .B2(_3931_),
    .A2(_1442_),
    .A1(net196));
 sg13g2_a21oi_1 _6228_ (.A1(_4141_),
    .A2(_4145_),
    .Y(_1444_),
    .B1(_1443_));
 sg13g2_a22oi_1 _6229_ (.Y(_1445_),
    .B1(_0326_),
    .B2(_0329_),
    .A2(_4145_),
    .A1(_4141_));
 sg13g2_nor3_1 _6230_ (.A(_4153_),
    .B(_1444_),
    .C(_1445_),
    .Y(_1446_));
 sg13g2_a21oi_1 _6231_ (.A1(_4114_),
    .A2(_4159_),
    .Y(_1447_),
    .B1(_4108_));
 sg13g2_o21ai_1 _6232_ (.B1(_1447_),
    .Y(_1448_),
    .A1(_1441_),
    .A2(_1446_));
 sg13g2_nand3b_1 _6233_ (.B(_1437_),
    .C(_1448_),
    .Y(_1449_),
    .A_N(_1222_));
 sg13g2_a21o_1 _6234_ (.A2(_4159_),
    .A1(_4114_),
    .B1(_4108_),
    .X(_1450_));
 sg13g2_inv_1 _6235_ (.Y(_1451_),
    .A(_4168_));
 sg13g2_o21ai_1 _6236_ (.B1(_4121_),
    .Y(_1452_),
    .A1(_0335_),
    .A2(_1451_));
 sg13g2_buf_1 _6237_ (.A(_1452_),
    .X(_1453_));
 sg13g2_nor2b_1 _6238_ (.A(_4150_),
    .B_N(_4152_),
    .Y(_1454_));
 sg13g2_a21o_1 _6239_ (.A2(_4145_),
    .A1(_4141_),
    .B1(_1443_),
    .X(_1455_));
 sg13g2_a221oi_1 _6240_ (.B2(_1455_),
    .C1(_0325_),
    .B1(_1454_),
    .A1(_4134_),
    .Y(_1456_),
    .A2(_4137_));
 sg13g2_nor3_1 _6241_ (.A(_1450_),
    .B(_1453_),
    .C(_1456_),
    .Y(_1457_));
 sg13g2_and4_1 _6242_ (.A(_1431_),
    .B(_1438_),
    .C(_1439_),
    .D(_1457_),
    .X(_1458_));
 sg13g2_a21oi_1 _6243_ (.A1(_0245_),
    .A2(_0248_),
    .Y(_1459_),
    .B1(_0311_));
 sg13g2_nand2b_1 _6244_ (.Y(_1460_),
    .B(_0316_),
    .A_N(_1459_));
 sg13g2_a22oi_1 _6245_ (.Y(_1461_),
    .B1(_0261_),
    .B2(_0267_),
    .A2(_0208_),
    .A1(_0206_));
 sg13g2_and2_1 _6246_ (.A(_4216_),
    .B(_1461_),
    .X(_1462_));
 sg13g2_and3_1 _6247_ (.X(_1463_),
    .A(_0255_),
    .B(_4216_),
    .C(_1461_));
 sg13g2_a22oi_1 _6248_ (.Y(_1464_),
    .B1(_1463_),
    .B2(_0242_),
    .A2(_1462_),
    .A1(_1460_));
 sg13g2_and2_1 _6249_ (.A(_0206_),
    .B(_0208_),
    .X(_1465_));
 sg13g2_and2_1 _6250_ (.A(_4206_),
    .B(_4201_),
    .X(_1466_));
 sg13g2_o21ai_1 _6251_ (.B1(_1466_),
    .Y(_1467_),
    .A1(_1465_),
    .A2(_0321_));
 sg13g2_and2_1 _6252_ (.A(_4195_),
    .B(_4198_),
    .X(_1468_));
 sg13g2_a21oi_1 _6253_ (.A1(_4206_),
    .A2(_1468_),
    .Y(_1469_),
    .B1(_4190_));
 sg13g2_and4_1 _6254_ (.A(_0255_),
    .B(_0279_),
    .C(_4216_),
    .D(_1461_),
    .X(_1470_));
 sg13g2_a21o_1 _6255_ (.A2(_0222_),
    .A1(_0219_),
    .B1(_0214_),
    .X(_1471_));
 sg13g2_nand3_1 _6256_ (.B(_1471_),
    .C(_4184_),
    .A(_4178_),
    .Y(_1472_));
 sg13g2_a221oi_1 _6257_ (.B2(_1470_),
    .C1(_1472_),
    .B1(_0308_),
    .A1(_1467_),
    .Y(_1473_),
    .A2(_1469_));
 sg13g2_a21o_1 _6258_ (.A2(_0222_),
    .A1(_0219_),
    .B1(_4213_),
    .X(_1474_));
 sg13g2_and3_1 _6259_ (.X(_1475_),
    .A(_4178_),
    .B(_1471_),
    .C(_1474_));
 sg13g2_a21o_1 _6260_ (.A2(_1473_),
    .A1(_1464_),
    .B1(_1475_),
    .X(_1476_));
 sg13g2_a21oi_1 _6261_ (.A1(_0225_),
    .A2(_0226_),
    .Y(_1477_),
    .B1(_0335_));
 sg13g2_nor4_1 _6262_ (.A(_1450_),
    .B(_1453_),
    .C(_1477_),
    .D(_1456_),
    .Y(_1478_));
 sg13g2_and4_1 _6263_ (.A(_1431_),
    .B(_1438_),
    .C(_1439_),
    .D(_1478_),
    .X(_1479_));
 sg13g2_a221oi_1 _6264_ (.B2(_1476_),
    .C1(_1479_),
    .B1(_1458_),
    .A1(_1440_),
    .Y(_1480_),
    .A2(_1449_));
 sg13g2_buf_2 _6265_ (.A(_1480_),
    .X(_1481_));
 sg13g2_xnor2_1 _6266_ (.Y(_1482_),
    .A(net142),
    .B(net141));
 sg13g2_xnor2_1 _6267_ (.Y(_1483_),
    .A(_1481_),
    .B(_1482_));
 sg13g2_nand2_1 _6268_ (.Y(_1484_),
    .A(net40),
    .B(_1483_));
 sg13g2_o21ai_1 _6269_ (.B1(_1484_),
    .Y(_1485_),
    .A1(net42),
    .A2(_1424_));
 sg13g2_nand2_1 _6270_ (.Y(_1486_),
    .A(net64),
    .B(_1485_));
 sg13g2_buf_1 _6271_ (.A(_0382_),
    .X(_1487_));
 sg13g2_a22oi_1 _6272_ (.Y(_1488_),
    .B1(_1243_),
    .B2(net141),
    .A2(_1239_),
    .A1(net265));
 sg13g2_a21oi_1 _6273_ (.A1(_1486_),
    .A2(_1488_),
    .Y(_0037_),
    .B1(net94));
 sg13g2_nand2_1 _6274_ (.Y(_1489_),
    .A(_0542_),
    .B(_0557_));
 sg13g2_a21oi_1 _6275_ (.A1(_0542_),
    .A2(_0573_),
    .Y(_1490_),
    .B1(_0579_));
 sg13g2_o21ai_1 _6276_ (.B1(_1490_),
    .Y(_1491_),
    .A1(_0506_),
    .A2(_1489_));
 sg13g2_a21o_1 _6277_ (.A2(_1491_),
    .A1(_0551_),
    .B1(_0568_),
    .X(_1492_));
 sg13g2_nor2_1 _6278_ (.A(_0510_),
    .B(_0558_),
    .Y(_1493_));
 sg13g2_nand2_1 _6279_ (.Y(_1494_),
    .A(_0474_),
    .B(_0480_));
 sg13g2_inv_1 _6280_ (.Y(_1495_),
    .A(_0483_));
 sg13g2_nand2_1 _6281_ (.Y(_1496_),
    .A(_0460_),
    .B(_0464_));
 sg13g2_o21ai_1 _6282_ (.B1(_1496_),
    .Y(_1497_),
    .A1(_1494_),
    .A2(_1495_));
 sg13g2_a21oi_1 _6283_ (.A1(_0453_),
    .A2(_1497_),
    .Y(_1498_),
    .B1(_0503_));
 sg13g2_nand2_1 _6284_ (.Y(_1499_),
    .A(_0519_),
    .B(_0522_));
 sg13g2_o21ai_1 _6285_ (.B1(_0447_),
    .Y(_1500_),
    .A1(_1498_),
    .A2(_1499_));
 sg13g2_a21oi_1 _6286_ (.A1(_0585_),
    .A2(_0586_),
    .Y(_1501_),
    .B1(_0590_));
 sg13g2_a22oi_1 _6287_ (.Y(_1502_),
    .B1(_0427_),
    .B2(_0429_),
    .A2(_0424_),
    .A1(_0421_));
 sg13g2_a22oi_1 _6288_ (.Y(_1503_),
    .B1(_0610_),
    .B2(_0612_),
    .A2(_0608_),
    .A1(_0607_));
 sg13g2_o21ai_1 _6289_ (.B1(_1503_),
    .Y(_1504_),
    .A1(_0602_),
    .A2(_1502_));
 sg13g2_nand3_1 _6290_ (.B(_1501_),
    .C(_1504_),
    .A(_0630_),
    .Y(_1505_));
 sg13g2_a221oi_1 _6291_ (.B2(_1500_),
    .C1(_1505_),
    .B1(_1493_),
    .A1(_0536_),
    .Y(_1506_),
    .A2(_1492_));
 sg13g2_nand3_1 _6292_ (.B(_0625_),
    .C(_0629_),
    .A(_0623_),
    .Y(_1507_));
 sg13g2_nor3_1 _6293_ (.A(_0602_),
    .B(_1502_),
    .C(_0597_),
    .Y(_1508_));
 sg13g2_nor2_1 _6294_ (.A(_0614_),
    .B(_1508_),
    .Y(_1509_));
 sg13g2_nor2_1 _6295_ (.A(_1507_),
    .B(_1509_),
    .Y(_1510_));
 sg13g2_inv_1 _6296_ (.Y(_1511_),
    .A(_3566_));
 sg13g2_nor2b_1 _6297_ (.A(_3456_),
    .B_N(net286),
    .Y(_1512_));
 sg13g2_nand3_1 _6298_ (.B(_1377_),
    .C(_1512_),
    .A(_1511_),
    .Y(_1513_));
 sg13g2_buf_1 _6299_ (.A(_1513_),
    .X(_1514_));
 sg13g2_inv_1 _6300_ (.Y(_1515_),
    .A(_3849_));
 sg13g2_nand4_1 _6301_ (.B(_1190_),
    .C(_1515_),
    .A(_3456_),
    .Y(_1516_),
    .D(_1434_));
 sg13g2_buf_1 _6302_ (.A(_1516_),
    .X(_1517_));
 sg13g2_a22oi_1 _6303_ (.Y(_1518_),
    .B1(_1514_),
    .B2(_1517_),
    .A2(_1313_),
    .A1(_1311_));
 sg13g2_buf_2 _6304_ (.A(_1518_),
    .X(_1519_));
 sg13g2_nand3_1 _6305_ (.B(_0663_),
    .C(_1519_),
    .A(_0655_),
    .Y(_1520_));
 sg13g2_or3_1 _6306_ (.A(_1281_),
    .B(_1510_),
    .C(_1520_),
    .X(_1521_));
 sg13g2_nand2_1 _6307_ (.Y(_1522_),
    .A(_1514_),
    .B(_1517_));
 sg13g2_a21oi_1 _6308_ (.A1(net200),
    .A2(net321),
    .Y(_1523_),
    .B1(_1246_));
 sg13g2_o21ai_1 _6309_ (.B1(_1249_),
    .Y(_1524_),
    .A1(_0701_),
    .A2(_1523_));
 sg13g2_nand2b_1 _6310_ (.Y(_1525_),
    .B(_0642_),
    .A_N(_0664_));
 sg13g2_nand2_1 _6311_ (.Y(_1526_),
    .A(_0689_),
    .B(_1525_));
 sg13g2_a22oi_1 _6312_ (.Y(_1527_),
    .B1(net301),
    .B2(_1417_),
    .A2(_1342_),
    .A1(_3743_));
 sg13g2_nand2b_1 _6313_ (.Y(_1528_),
    .B(net144),
    .A_N(_1527_));
 sg13g2_o21ai_1 _6314_ (.B1(net142),
    .Y(_1529_),
    .A1(net143),
    .A2(_1417_));
 sg13g2_nand2_1 _6315_ (.Y(_1530_),
    .A(_1528_),
    .B(_1529_));
 sg13g2_a221oi_1 _6316_ (.B2(_1526_),
    .C1(_1530_),
    .B1(_1519_),
    .A1(_1522_),
    .Y(_1531_),
    .A2(_1524_));
 sg13g2_o21ai_1 _6317_ (.B1(_1531_),
    .Y(_1532_),
    .A1(_1506_),
    .A2(_1521_));
 sg13g2_buf_1 _6318_ (.A(_3577_),
    .X(_1533_));
 sg13g2_xor2_1 _6319_ (.B(net141),
    .A(net140),
    .X(_1534_));
 sg13g2_xnor2_1 _6320_ (.Y(_1535_),
    .A(_1532_),
    .B(_1534_));
 sg13g2_buf_1 _6321_ (.A(net285),
    .X(_1536_));
 sg13g2_nor2_1 _6322_ (.A(net35),
    .B(net139),
    .Y(_1537_));
 sg13g2_a21oi_1 _6323_ (.A1(net37),
    .A2(_1535_),
    .Y(_1538_),
    .B1(_1537_));
 sg13g2_nand2_1 _6324_ (.Y(_1539_),
    .A(net64),
    .B(_1538_));
 sg13g2_a22oi_1 _6325_ (.Y(_1540_),
    .B1(_1243_),
    .B2(net140),
    .A2(_1239_),
    .A1(net266));
 sg13g2_a21oi_1 _6326_ (.A1(_1539_),
    .A2(_1540_),
    .Y(_0038_),
    .B1(net94));
 sg13g2_nand2_1 _6327_ (.Y(_1541_),
    .A(_0755_),
    .B(_0756_));
 sg13g2_a21oi_1 _6328_ (.A1(_0753_),
    .A2(_1541_),
    .Y(_1542_),
    .B1(_0747_));
 sg13g2_xor2_1 _6329_ (.B(net177),
    .A(net251),
    .X(_1543_));
 sg13g2_xnor2_1 _6330_ (.Y(_1544_),
    .A(_1542_),
    .B(_1543_));
 sg13g2_nand2_1 _6331_ (.Y(_1545_),
    .A(net36),
    .B(_1544_));
 sg13g2_o21ai_1 _6332_ (.B1(_1545_),
    .Y(_1546_),
    .A1(net42),
    .A2(_0275_));
 sg13g2_nor2_1 _6333_ (.A(net65),
    .B(_1546_),
    .Y(_1547_));
 sg13g2_nand2_1 _6334_ (.Y(_1548_),
    .A(_3975_),
    .B(_3978_));
 sg13g2_nor4_1 _6335_ (.A(_3977_),
    .B(_3980_),
    .C(_4000_),
    .D(_1548_),
    .Y(_1549_));
 sg13g2_nor2b_1 _6336_ (.A(_3976_),
    .B_N(_1549_),
    .Y(_1550_));
 sg13g2_buf_1 _6337_ (.A(_1550_),
    .X(_1551_));
 sg13g2_buf_1 _6338_ (.A(_1551_),
    .X(_1552_));
 sg13g2_nor2_1 _6339_ (.A(_0286_),
    .B(net63),
    .Y(_1553_));
 sg13g2_a221oi_1 _6340_ (.B2(net18),
    .C1(net76),
    .B1(_1553_),
    .A1(_1348_),
    .Y(_1554_),
    .A2(net63));
 sg13g2_nor3_1 _6341_ (.A(_0403_),
    .B(_1547_),
    .C(_1554_),
    .Y(_0039_));
 sg13g2_nor3_1 _6342_ (.A(_0883_),
    .B(_0872_),
    .C(_0888_),
    .Y(_1555_));
 sg13g2_nand2b_1 _6343_ (.Y(_1556_),
    .B(_0825_),
    .A_N(_1555_));
 sg13g2_nand3_1 _6344_ (.B(_0767_),
    .C(_0778_),
    .A(_0774_),
    .Y(_1557_));
 sg13g2_nand2_1 _6345_ (.Y(_1558_),
    .A(_0774_),
    .B(_0806_));
 sg13g2_o21ai_1 _6346_ (.B1(_1558_),
    .Y(_1559_),
    .A1(_0763_),
    .A2(_1557_));
 sg13g2_nor4_1 _6347_ (.A(_0881_),
    .B(_0883_),
    .C(_0888_),
    .D(_0792_),
    .Y(_1560_));
 sg13g2_or4_1 _6348_ (.A(_0881_),
    .B(_0883_),
    .C(_0888_),
    .D(_0868_),
    .X(_1561_));
 sg13g2_inv_1 _6349_ (.Y(_1562_),
    .A(_0862_));
 sg13g2_a21oi_1 _6350_ (.A1(_0789_),
    .A2(_0790_),
    .Y(_1563_),
    .B1(_0796_));
 sg13g2_o21ai_1 _6351_ (.B1(_0786_),
    .Y(_1564_),
    .A1(_1562_),
    .A2(_1563_));
 sg13g2_a21o_1 _6352_ (.A2(_0781_),
    .A1(_0780_),
    .B1(_0866_),
    .X(_1565_));
 sg13g2_and3_1 _6353_ (.X(_1566_),
    .A(_0851_),
    .B(_0859_),
    .C(_1565_));
 sg13g2_a22oi_1 _6354_ (.Y(_1567_),
    .B1(_1564_),
    .B2(_1566_),
    .A2(_1561_),
    .A1(_0851_));
 sg13g2_a221oi_1 _6355_ (.B2(_1560_),
    .C1(_1567_),
    .B1(_1559_),
    .A1(_0837_),
    .Y(_1568_),
    .A2(_1556_));
 sg13g2_buf_1 _6356_ (.A(_1568_),
    .X(_1569_));
 sg13g2_nor2_1 _6357_ (.A(_0842_),
    .B(_0847_),
    .Y(_1570_));
 sg13g2_o21ai_1 _6358_ (.B1(_1570_),
    .Y(_1571_),
    .A1(_0879_),
    .A2(_1569_));
 sg13g2_a22oi_1 _6359_ (.Y(_1572_),
    .B1(_0738_),
    .B2(_0739_),
    .A2(_0812_),
    .A1(_0810_));
 sg13g2_nand3b_1 _6360_ (.B(net147),
    .C(net114),
    .Y(_1573_),
    .A_N(_0876_));
 sg13g2_a22oi_1 _6361_ (.Y(_1574_),
    .B1(_0948_),
    .B2(net238),
    .A2(net147),
    .A1(net229));
 sg13g2_nand3b_1 _6362_ (.B(_4136_),
    .C(net230),
    .Y(_1575_),
    .A_N(_0876_));
 sg13g2_nand3_1 _6363_ (.B(net114),
    .C(net147),
    .A(net230),
    .Y(_1576_));
 sg13g2_nand4_1 _6364_ (.B(_1574_),
    .C(_1575_),
    .A(_1573_),
    .Y(_1577_),
    .D(_1576_));
 sg13g2_a21o_1 _6365_ (.A2(_1572_),
    .A1(_1571_),
    .B1(_1577_),
    .X(_1578_));
 sg13g2_a21oi_2 _6366_ (.B1(_0911_),
    .Y(_1579_),
    .A2(_0900_),
    .A1(_0896_));
 sg13g2_a21oi_1 _6367_ (.A1(net244),
    .A2(net148),
    .Y(_1580_),
    .B1(net157));
 sg13g2_nand2b_1 _6368_ (.Y(_1581_),
    .B(_0910_),
    .A_N(_1580_));
 sg13g2_nand3b_1 _6369_ (.B(_0606_),
    .C(net244),
    .Y(_1582_),
    .A_N(_0955_));
 sg13g2_a21o_1 _6370_ (.A2(net192),
    .A1(net229),
    .B1(net98),
    .X(_1583_));
 sg13g2_nand3_1 _6371_ (.B(_0606_),
    .C(_1583_),
    .A(net96),
    .Y(_1584_));
 sg13g2_nand4_1 _6372_ (.B(_1581_),
    .C(_1582_),
    .A(_0929_),
    .Y(_1585_),
    .D(_1584_));
 sg13g2_a21oi_1 _6373_ (.A1(_1578_),
    .A2(_1579_),
    .Y(_1586_),
    .B1(_1585_));
 sg13g2_nor2b_1 _6374_ (.A(_1586_),
    .B_N(_0922_),
    .Y(_1587_));
 sg13g2_nand3_1 _6375_ (.B(_0906_),
    .C(_0914_),
    .A(_0903_),
    .Y(_1588_));
 sg13g2_nand3_1 _6376_ (.B(_3588_),
    .C(_1512_),
    .A(net143),
    .Y(_1589_));
 sg13g2_nor2b_1 _6377_ (.A(net286),
    .B_N(_3577_),
    .Y(_1590_));
 sg13g2_nand3_1 _6378_ (.B(_1434_),
    .C(_1590_),
    .A(net144),
    .Y(_1591_));
 sg13g2_a22oi_1 _6379_ (.Y(_1592_),
    .B1(_1589_),
    .B2(_1591_),
    .A2(_1332_),
    .A1(_1330_));
 sg13g2_nor2b_1 _6380_ (.A(_1588_),
    .B_N(_1592_),
    .Y(_1593_));
 sg13g2_a221oi_1 _6381_ (.B2(net173),
    .C1(_0639_),
    .B1(_0932_),
    .A1(net155),
    .Y(_1594_),
    .A2(_0931_));
 sg13g2_or3_1 _6382_ (.A(net219),
    .B(net198),
    .C(net171),
    .X(_1595_));
 sg13g2_a221oi_1 _6383_ (.B2(net173),
    .C1(_1595_),
    .B1(_0932_),
    .A1(net155),
    .Y(_1596_),
    .A2(_0931_));
 sg13g2_nor2_1 _6384_ (.A(net111),
    .B(_0639_),
    .Y(_1597_));
 sg13g2_nor4_2 _6385_ (.A(_0939_),
    .B(_1594_),
    .C(_1596_),
    .Y(_1598_),
    .D(_1597_));
 sg13g2_nand3_1 _6386_ (.B(_1598_),
    .C(_0914_),
    .A(_0906_),
    .Y(_1599_));
 sg13g2_a22oi_1 _6387_ (.Y(_1600_),
    .B1(_0727_),
    .B2(_0729_),
    .A2(_0715_),
    .A1(_0713_));
 sg13g2_a21oi_1 _6388_ (.A1(_0904_),
    .A2(_0905_),
    .Y(_1601_),
    .B1(_0943_));
 sg13g2_nor4_1 _6389_ (.A(_0736_),
    .B(_1600_),
    .C(_0725_),
    .D(_1601_),
    .Y(_1602_));
 sg13g2_o21ai_1 _6390_ (.B1(net169),
    .Y(_1603_),
    .A1(net151),
    .A2(net168));
 sg13g2_o21ai_1 _6391_ (.B1(net168),
    .Y(_1604_),
    .A1(_0717_),
    .A2(net151));
 sg13g2_and2_1 _6392_ (.A(_0644_),
    .B(_1604_),
    .X(_1605_));
 sg13g2_a221oi_1 _6393_ (.B2(_1183_),
    .C1(_1605_),
    .B1(_1603_),
    .A1(_0713_),
    .Y(_1606_),
    .A2(_0715_));
 sg13g2_o21ai_1 _6394_ (.B1(_1592_),
    .Y(_1607_),
    .A1(_0736_),
    .A2(_1606_));
 sg13g2_a21oi_1 _6395_ (.A1(_1599_),
    .A2(_1602_),
    .Y(_1608_),
    .B1(_1607_));
 sg13g2_a21oi_1 _6396_ (.A1(_3456_),
    .A2(net301),
    .Y(_1609_),
    .B1(_1533_));
 sg13g2_and2_1 _6397_ (.A(net301),
    .B(_3577_),
    .X(_1610_));
 sg13g2_o21ai_1 _6398_ (.B1(_3566_),
    .Y(_1611_),
    .A1(net141),
    .A2(_1610_));
 sg13g2_o21ai_1 _6399_ (.B1(_1611_),
    .Y(_1612_),
    .A1(_1515_),
    .A2(_1609_));
 sg13g2_a22oi_1 _6400_ (.Y(_1613_),
    .B1(_1336_),
    .B2(net146),
    .A2(_1334_),
    .A1(_1225_));
 sg13g2_a21oi_1 _6401_ (.A1(_1589_),
    .A2(_1591_),
    .Y(_1614_),
    .B1(_1613_));
 sg13g2_nor2_1 _6402_ (.A(_1612_),
    .B(_1614_),
    .Y(_1615_));
 sg13g2_nand2b_1 _6403_ (.Y(_1616_),
    .B(_1615_),
    .A_N(_1608_));
 sg13g2_a21oi_2 _6404_ (.B1(_1616_),
    .Y(_1617_),
    .A2(_1593_),
    .A1(_1587_));
 sg13g2_xnor2_1 _6405_ (.Y(_1618_),
    .A(net140),
    .B(net139));
 sg13g2_xnor2_1 _6406_ (.Y(_1619_),
    .A(_1617_),
    .B(_1618_));
 sg13g2_nor2_1 _6407_ (.A(net35),
    .B(net223),
    .Y(_1620_));
 sg13g2_a21oi_1 _6408_ (.A1(net37),
    .A2(_1619_),
    .Y(_1621_),
    .B1(_1620_));
 sg13g2_nand2_1 _6409_ (.Y(_1622_),
    .A(net64),
    .B(_1621_));
 sg13g2_buf_1 _6410_ (.A(net325),
    .X(_1623_));
 sg13g2_a22oi_1 _6411_ (.Y(_1624_),
    .B1(_1243_),
    .B2(net139),
    .A2(_1239_),
    .A1(net264));
 sg13g2_a21oi_1 _6412_ (.A1(_1622_),
    .A2(_1624_),
    .Y(_0040_),
    .B1(net94));
 sg13g2_nand2_1 _6413_ (.Y(_1625_),
    .A(_1103_),
    .B(_1107_));
 sg13g2_o21ai_1 _6414_ (.B1(_1113_),
    .Y(_1626_),
    .A1(_1073_),
    .A2(_1092_));
 sg13g2_nor2b_1 _6415_ (.A(_1168_),
    .B_N(_1626_),
    .Y(_1627_));
 sg13g2_and2_1 _6416_ (.A(_1121_),
    .B(_1125_),
    .X(_1628_));
 sg13g2_o21ai_1 _6417_ (.B1(_1628_),
    .Y(_1629_),
    .A1(_1625_),
    .A2(_1627_));
 sg13g2_nand4_1 _6418_ (.B(net141),
    .C(net139),
    .A(net301),
    .Y(_1630_),
    .D(_3588_));
 sg13g2_nand3_1 _6419_ (.B(_3851_),
    .C(_1434_),
    .A(_1533_),
    .Y(_1631_));
 sg13g2_a22oi_1 _6420_ (.Y(_1632_),
    .B1(_1630_),
    .B2(_1631_),
    .A2(_1379_),
    .A1(_1378_));
 sg13g2_a22oi_1 _6421_ (.Y(_1633_),
    .B1(_0992_),
    .B2(_0993_),
    .A2(_0984_),
    .A1(_0983_));
 sg13g2_and4_1 _6422_ (.A(_1099_),
    .B(_1393_),
    .C(_1632_),
    .D(_1633_),
    .X(_1634_));
 sg13g2_buf_1 _6423_ (.A(_1634_),
    .X(_1635_));
 sg13g2_nand2_1 _6424_ (.Y(_1636_),
    .A(_1630_),
    .B(_1631_));
 sg13g2_nand2_1 _6425_ (.Y(_1637_),
    .A(_1380_),
    .B(_1636_));
 sg13g2_nor2_1 _6426_ (.A(_1187_),
    .B(_1637_),
    .Y(_1638_));
 sg13g2_o21ai_1 _6427_ (.B1(_0990_),
    .Y(_1639_),
    .A1(_1179_),
    .A2(_0996_));
 sg13g2_a21oi_1 _6428_ (.A1(net141),
    .A2(_1536_),
    .Y(_1640_),
    .B1(_1610_));
 sg13g2_o21ai_1 _6429_ (.B1(net140),
    .Y(_1641_),
    .A1(net141),
    .A2(_1536_));
 sg13g2_o21ai_1 _6430_ (.B1(_1641_),
    .Y(_1642_),
    .A1(_1511_),
    .A2(_1640_));
 sg13g2_and2_1 _6431_ (.A(net150),
    .B(net144),
    .X(_1643_));
 sg13g2_o21ai_1 _6432_ (.B1(net146),
    .Y(_1644_),
    .A1(_1643_),
    .A2(_1377_));
 sg13g2_a22oi_1 _6433_ (.Y(_1645_),
    .B1(_1644_),
    .B2(_1408_),
    .A2(_1631_),
    .A1(_1630_));
 sg13g2_or2_1 _6434_ (.X(_1646_),
    .B(_1645_),
    .A(_1642_));
 sg13g2_a21o_1 _6435_ (.A2(_1639_),
    .A1(_1638_),
    .B1(_1646_),
    .X(_1647_));
 sg13g2_a21oi_2 _6436_ (.B1(_1647_),
    .Y(_1648_),
    .A2(_1635_),
    .A1(_1629_));
 sg13g2_xnor2_1 _6437_ (.Y(_1649_),
    .A(net223),
    .B(net139));
 sg13g2_xnor2_1 _6438_ (.Y(_1650_),
    .A(_1648_),
    .B(_1649_));
 sg13g2_buf_1 _6439_ (.A(_3804_),
    .X(_1651_));
 sg13g2_nor2_1 _6440_ (.A(net35),
    .B(net138),
    .Y(_1652_));
 sg13g2_a21oi_1 _6441_ (.A1(net37),
    .A2(_1650_),
    .Y(_1653_),
    .B1(_1652_));
 sg13g2_nand2_1 _6442_ (.Y(_1654_),
    .A(net64),
    .B(_1653_));
 sg13g2_buf_1 _6443_ (.A(_1194_),
    .X(_1655_));
 sg13g2_a22oi_1 _6444_ (.Y(_1656_),
    .B1(_1243_),
    .B2(net223),
    .A2(_1239_),
    .A1(net263));
 sg13g2_a21oi_1 _6445_ (.A1(_1654_),
    .A2(_1656_),
    .Y(_0041_),
    .B1(net94));
 sg13g2_buf_1 _6446_ (.A(net80),
    .X(_1657_));
 sg13g2_nor2b_1 _6447_ (.A(net285),
    .B_N(_3901_),
    .Y(_1658_));
 sg13g2_nand3_1 _6448_ (.B(_1590_),
    .C(_1658_),
    .A(_3566_),
    .Y(_1659_));
 sg13g2_inv_1 _6449_ (.Y(_1660_),
    .A(_3901_));
 sg13g2_nand4_1 _6450_ (.B(_1660_),
    .C(net139),
    .A(_3849_),
    .Y(_1661_),
    .D(_3588_));
 sg13g2_and2_1 _6451_ (.A(_1659_),
    .B(_1661_),
    .X(_1662_));
 sg13g2_buf_1 _6452_ (.A(_1662_),
    .X(_1663_));
 sg13g2_nor2_1 _6453_ (.A(_1436_),
    .B(_1663_),
    .Y(_1664_));
 sg13g2_a21o_1 _6454_ (.A2(net145),
    .A1(net146),
    .B1(net142),
    .X(_1665_));
 sg13g2_a21oi_1 _6455_ (.A1(_1319_),
    .A2(_1665_),
    .Y(_1666_),
    .B1(_1427_));
 sg13g2_a21o_1 _6456_ (.A2(net286),
    .A1(_3566_),
    .B1(_3901_),
    .X(_1667_));
 sg13g2_a21o_1 _6457_ (.A2(_3901_),
    .A1(net286),
    .B1(net285),
    .X(_1668_));
 sg13g2_a22oi_1 _6458_ (.Y(_1669_),
    .B1(_1668_),
    .B2(net140),
    .A2(_1667_),
    .A1(net285));
 sg13g2_o21ai_1 _6459_ (.B1(_1669_),
    .Y(_1670_),
    .A1(_1663_),
    .A2(_1666_));
 sg13g2_a21oi_1 _6460_ (.A1(_1224_),
    .A2(_1664_),
    .Y(_1671_),
    .B1(_1670_));
 sg13g2_xnor2_1 _6461_ (.Y(_1672_),
    .A(net223),
    .B(net138));
 sg13g2_xnor2_1 _6462_ (.Y(_1673_),
    .A(_1671_),
    .B(_1672_));
 sg13g2_buf_1 _6463_ (.A(net280),
    .X(_1674_));
 sg13g2_nor2_1 _6464_ (.A(net35),
    .B(net137),
    .Y(_1675_));
 sg13g2_a21oi_1 _6465_ (.A1(net37),
    .A2(_1673_),
    .Y(_1676_),
    .B1(_1675_));
 sg13g2_nand2_1 _6466_ (.Y(_1677_),
    .A(net62),
    .B(_1676_));
 sg13g2_nand3_1 _6467_ (.B(net329),
    .C(net272),
    .A(_3979_),
    .Y(_1678_));
 sg13g2_nor2_1 _6468_ (.A(_1237_),
    .B(_1678_),
    .Y(_1679_));
 sg13g2_buf_2 _6469_ (.A(_1679_),
    .X(_1680_));
 sg13g2_inv_1 _6470_ (.Y(_1681_),
    .A(_1678_));
 sg13g2_a21oi_1 _6471_ (.A1(net66),
    .A2(_1681_),
    .Y(_1682_),
    .B1(net100));
 sg13g2_buf_2 _6472_ (.A(_1682_),
    .X(_1683_));
 sg13g2_a22oi_1 _6473_ (.Y(_1684_),
    .B1(_1683_),
    .B2(net138),
    .A2(_1680_),
    .A1(net328));
 sg13g2_a21oi_1 _6474_ (.A1(_1677_),
    .A2(_1684_),
    .Y(_0042_),
    .B1(_1326_));
 sg13g2_buf_1 _6475_ (.A(_3805_),
    .X(_1685_));
 sg13g2_inv_1 _6476_ (.Y(_1686_),
    .A(net136));
 sg13g2_buf_1 _6477_ (.A(net52),
    .X(_1687_));
 sg13g2_a22oi_1 _6478_ (.Y(_1688_),
    .B1(net285),
    .B2(net138),
    .A2(net223),
    .A1(net286));
 sg13g2_o21ai_1 _6479_ (.B1(net223),
    .Y(_1689_),
    .A1(net285),
    .A2(_3804_));
 sg13g2_o21ai_1 _6480_ (.B1(_1689_),
    .Y(_1690_),
    .A1(_1424_),
    .A2(_1688_));
 sg13g2_and2_1 _6481_ (.A(net285),
    .B(_3804_),
    .X(_1691_));
 sg13g2_nand4_1 _6482_ (.B(net286),
    .C(_1660_),
    .A(_1424_),
    .Y(_1692_),
    .D(_1691_));
 sg13g2_inv_1 _6483_ (.Y(_1693_),
    .A(_3804_));
 sg13g2_nand3_1 _6484_ (.B(_1590_),
    .C(_1658_),
    .A(_1693_),
    .Y(_1694_));
 sg13g2_a22oi_1 _6485_ (.Y(_1695_),
    .B1(_1692_),
    .B2(_1694_),
    .A2(_1529_),
    .A1(_1528_));
 sg13g2_and2_1 _6486_ (.A(_1514_),
    .B(_1517_),
    .X(_1696_));
 sg13g2_a221oi_1 _6487_ (.B2(_1694_),
    .C1(_1696_),
    .B1(_1692_),
    .A1(_1253_),
    .Y(_1697_),
    .A2(_1315_));
 sg13g2_or3_1 _6488_ (.A(_1690_),
    .B(_1695_),
    .C(_1697_),
    .X(_1698_));
 sg13g2_xnor2_1 _6489_ (.Y(_1699_),
    .A(net137),
    .B(net138));
 sg13g2_xnor2_1 _6490_ (.Y(_1700_),
    .A(_1698_),
    .B(_1699_));
 sg13g2_nand2_1 _6491_ (.Y(_1701_),
    .A(net34),
    .B(_1700_));
 sg13g2_o21ai_1 _6492_ (.B1(_1701_),
    .Y(_1702_),
    .A1(net42),
    .A2(_1686_));
 sg13g2_nand2_1 _6493_ (.Y(_1703_),
    .A(net62),
    .B(_1702_));
 sg13g2_a22oi_1 _6494_ (.Y(_1704_),
    .B1(_1683_),
    .B2(net137),
    .A2(_1680_),
    .A1(net274));
 sg13g2_a21oi_1 _6495_ (.A1(_1703_),
    .A2(_1704_),
    .Y(_0043_),
    .B1(net94));
 sg13g2_buf_1 _6496_ (.A(net51),
    .X(_1705_));
 sg13g2_nand2_1 _6497_ (.Y(_1706_),
    .A(_1589_),
    .B(_1591_));
 sg13g2_nor2b_1 _6498_ (.A(_3804_),
    .B_N(net280),
    .Y(_1707_));
 sg13g2_nand3_1 _6499_ (.B(_1658_),
    .C(_1707_),
    .A(net140),
    .Y(_1708_));
 sg13g2_nor2_1 _6500_ (.A(_3901_),
    .B(net280),
    .Y(_1709_));
 sg13g2_nand3b_1 _6501_ (.B(_1709_),
    .C(_1691_),
    .Y(_1710_),
    .A_N(net140));
 sg13g2_nand2_1 _6502_ (.Y(_1711_),
    .A(_1708_),
    .B(_1710_));
 sg13g2_nand2_1 _6503_ (.Y(_1712_),
    .A(_1706_),
    .B(_1711_));
 sg13g2_and2_1 _6504_ (.A(net285),
    .B(net280),
    .X(_1713_));
 sg13g2_o21ai_1 _6505_ (.B1(net223),
    .Y(_1714_),
    .A1(net138),
    .A2(_1713_));
 sg13g2_a21oi_1 _6506_ (.A1(net140),
    .A2(net139),
    .Y(_1715_),
    .B1(net280));
 sg13g2_nand2b_1 _6507_ (.Y(_1716_),
    .B(net138),
    .A_N(_1715_));
 sg13g2_nand2_1 _6508_ (.Y(_1717_),
    .A(_1714_),
    .B(_1716_));
 sg13g2_a21oi_1 _6509_ (.A1(_1612_),
    .A2(_1711_),
    .Y(_1718_),
    .B1(_1717_));
 sg13g2_o21ai_1 _6510_ (.B1(_1718_),
    .Y(_1719_),
    .A1(_1339_),
    .A2(_1712_));
 sg13g2_xor2_1 _6511_ (.B(net136),
    .A(net137),
    .X(_1720_));
 sg13g2_xnor2_1 _6512_ (.Y(_1721_),
    .A(_1719_),
    .B(_1720_));
 sg13g2_buf_1 _6513_ (.A(net279),
    .X(_1722_));
 sg13g2_nor2_1 _6514_ (.A(net35),
    .B(net135),
    .Y(_1723_));
 sg13g2_a21oi_1 _6515_ (.A1(net33),
    .A2(_1721_),
    .Y(_1724_),
    .B1(_1723_));
 sg13g2_nand2_1 _6516_ (.Y(_1725_),
    .A(net62),
    .B(_1724_));
 sg13g2_buf_1 _6517_ (.A(_1346_),
    .X(_1726_));
 sg13g2_a22oi_1 _6518_ (.Y(_1727_),
    .B1(_1683_),
    .B2(net136),
    .A2(_1680_),
    .A1(net262));
 sg13g2_a21oi_1 _6519_ (.A1(_1725_),
    .A2(_1727_),
    .Y(_0044_),
    .B1(net94));
 sg13g2_and2_1 _6520_ (.A(_3804_),
    .B(_3805_),
    .X(_1728_));
 sg13g2_buf_1 _6521_ (.A(_1728_),
    .X(_1729_));
 sg13g2_nand3_1 _6522_ (.B(_1709_),
    .C(_1729_),
    .A(net139),
    .Y(_1730_));
 sg13g2_nand3_1 _6523_ (.B(_3807_),
    .C(_1658_),
    .A(net137),
    .Y(_1731_));
 sg13g2_nand2_1 _6524_ (.Y(_1732_),
    .A(_1730_),
    .B(_1731_));
 sg13g2_nand2_1 _6525_ (.Y(_1733_),
    .A(_1636_),
    .B(_1732_));
 sg13g2_inv_1 _6526_ (.Y(_1734_),
    .A(net137));
 sg13g2_o21ai_1 _6527_ (.B1(_3902_),
    .Y(_1735_),
    .A1(_1713_),
    .A2(_1729_));
 sg13g2_o21ai_1 _6528_ (.B1(_1735_),
    .Y(_1736_),
    .A1(_1734_),
    .A2(_3807_));
 sg13g2_a21oi_1 _6529_ (.A1(_1642_),
    .A2(_1732_),
    .Y(_1737_),
    .B1(_1736_));
 sg13g2_o21ai_1 _6530_ (.B1(_1737_),
    .Y(_1738_),
    .A1(_1413_),
    .A2(_1733_));
 sg13g2_xor2_1 _6531_ (.B(_1685_),
    .A(_1722_),
    .X(_1739_));
 sg13g2_xnor2_1 _6532_ (.Y(_1740_),
    .A(_1738_),
    .B(_1739_));
 sg13g2_buf_1 _6533_ (.A(net322),
    .X(_1741_));
 sg13g2_nor2_1 _6534_ (.A(net35),
    .B(net134),
    .Y(_1742_));
 sg13g2_a21oi_1 _6535_ (.A1(net33),
    .A2(_1740_),
    .Y(_1743_),
    .B1(_1742_));
 sg13g2_nand2_1 _6536_ (.Y(_1744_),
    .A(net62),
    .B(_1743_));
 sg13g2_buf_1 _6537_ (.A(net2),
    .X(_1745_));
 sg13g2_a22oi_1 _6538_ (.Y(_1746_),
    .B1(_1683_),
    .B2(net135),
    .A2(_1680_),
    .A1(net323));
 sg13g2_buf_2 _6539_ (.A(net204),
    .X(_1747_));
 sg13g2_a21oi_1 _6540_ (.A1(_1744_),
    .A2(_1746_),
    .Y(_0045_),
    .B1(_1747_));
 sg13g2_nand3_1 _6541_ (.B(net135),
    .C(_3807_),
    .A(_1674_),
    .Y(_1748_));
 sg13g2_nand2_1 _6542_ (.Y(_1749_),
    .A(_3905_),
    .B(_1729_));
 sg13g2_o21ai_1 _6543_ (.B1(_1749_),
    .Y(_1750_),
    .A1(_1660_),
    .A2(_1748_));
 sg13g2_nor2b_1 _6544_ (.A(_1663_),
    .B_N(_1750_),
    .Y(_1751_));
 sg13g2_inv_1 _6545_ (.Y(_1752_),
    .A(net279));
 sg13g2_a21o_1 _6546_ (.A2(_1669_),
    .A1(_1693_),
    .B1(_1752_),
    .X(_1753_));
 sg13g2_nor2_1 _6547_ (.A(net280),
    .B(net279),
    .Y(_1754_));
 sg13g2_a21o_1 _6548_ (.A2(_1754_),
    .A1(_1669_),
    .B1(_3807_),
    .X(_1755_));
 sg13g2_o21ai_1 _6549_ (.B1(net136),
    .Y(_1756_),
    .A1(net138),
    .A2(net279));
 sg13g2_and2_1 _6550_ (.A(_1734_),
    .B(_1756_),
    .X(_1757_));
 sg13g2_a221oi_1 _6551_ (.B2(_1660_),
    .C1(_1757_),
    .B1(_1755_),
    .A1(_1686_),
    .Y(_1758_),
    .A2(_1753_));
 sg13g2_a21oi_1 _6552_ (.A1(_1481_),
    .A2(_1751_),
    .Y(_1759_),
    .B1(_1758_));
 sg13g2_xnor2_1 _6553_ (.Y(_1760_),
    .A(net135),
    .B(net134));
 sg13g2_xnor2_1 _6554_ (.Y(_1761_),
    .A(_1759_),
    .B(_1760_));
 sg13g2_nor2_1 _6555_ (.A(net35),
    .B(net261),
    .Y(_1762_));
 sg13g2_a21oi_1 _6556_ (.A1(net33),
    .A2(_1761_),
    .Y(_1763_),
    .B1(_1762_));
 sg13g2_nand2_1 _6557_ (.Y(_1764_),
    .A(net62),
    .B(_1763_));
 sg13g2_a22oi_1 _6558_ (.Y(_1765_),
    .B1(_1683_),
    .B2(net134),
    .A2(_1680_),
    .A1(net265));
 sg13g2_a21oi_1 _6559_ (.A1(_1764_),
    .A2(_1765_),
    .Y(_0046_),
    .B1(_1747_));
 sg13g2_nand3_1 _6560_ (.B(_1729_),
    .C(_1754_),
    .A(net322),
    .Y(_1766_));
 sg13g2_nor2_1 _6561_ (.A(_3805_),
    .B(net322),
    .Y(_1767_));
 sg13g2_nand3_1 _6562_ (.B(_1707_),
    .C(_1767_),
    .A(net279),
    .Y(_1768_));
 sg13g2_a22oi_1 _6563_ (.Y(_1769_),
    .B1(_1766_),
    .B2(_1768_),
    .A2(_1694_),
    .A1(_1692_));
 sg13g2_buf_2 _6564_ (.A(_1769_),
    .X(_1770_));
 sg13g2_a21oi_1 _6565_ (.A1(net136),
    .A2(net322),
    .Y(_1771_),
    .B1(net279));
 sg13g2_nor3_1 _6566_ (.A(net280),
    .B(net136),
    .C(net134),
    .Y(_1772_));
 sg13g2_or2_1 _6567_ (.X(_1773_),
    .B(_1772_),
    .A(_1771_));
 sg13g2_inv_1 _6568_ (.Y(_1774_),
    .A(_1689_));
 sg13g2_nor2_1 _6569_ (.A(_1424_),
    .B(_1688_),
    .Y(_1775_));
 sg13g2_nor4_1 _6570_ (.A(net137),
    .B(net135),
    .C(_1774_),
    .D(_1775_),
    .Y(_1776_));
 sg13g2_nor3_1 _6571_ (.A(net137),
    .B(_1651_),
    .C(net135),
    .Y(_1777_));
 sg13g2_nand2_1 _6572_ (.Y(_1778_),
    .A(_1693_),
    .B(_1686_));
 sg13g2_nor4_1 _6573_ (.A(net134),
    .B(_1778_),
    .C(_1774_),
    .D(_1775_),
    .Y(_1779_));
 sg13g2_nor4_1 _6574_ (.A(_1773_),
    .B(_1776_),
    .C(_1777_),
    .D(_1779_),
    .Y(_1780_));
 sg13g2_a21oi_1 _6575_ (.A1(_1532_),
    .A2(_1770_),
    .Y(_1781_),
    .B1(_1780_));
 sg13g2_nor2b_1 _6576_ (.A(_3473_),
    .B_N(net322),
    .Y(_1782_));
 sg13g2_buf_2 _6577_ (.A(_1782_),
    .X(_1783_));
 sg13g2_nor2b_1 _6578_ (.A(net322),
    .B_N(_3473_),
    .Y(_1784_));
 sg13g2_nor2_1 _6579_ (.A(_1783_),
    .B(_1784_),
    .Y(_1785_));
 sg13g2_xnor2_1 _6580_ (.Y(_1786_),
    .A(_1781_),
    .B(_1785_));
 sg13g2_buf_1 _6581_ (.A(_3399_),
    .X(_1787_));
 sg13g2_nor2_1 _6582_ (.A(_1416_),
    .B(net133),
    .Y(_1788_));
 sg13g2_a21oi_1 _6583_ (.A1(net33),
    .A2(_1786_),
    .Y(_1789_),
    .B1(_1788_));
 sg13g2_nand2_1 _6584_ (.Y(_1790_),
    .A(net62),
    .B(_1789_));
 sg13g2_a22oi_1 _6585_ (.Y(_1791_),
    .B1(_1683_),
    .B2(net261),
    .A2(_1680_),
    .A1(net266));
 sg13g2_a21oi_1 _6586_ (.A1(_1790_),
    .A2(_1791_),
    .Y(_0047_),
    .B1(_1747_));
 sg13g2_nand3_1 _6587_ (.B(_1754_),
    .C(_1783_),
    .A(net136),
    .Y(_1792_));
 sg13g2_nand4_1 _6588_ (.B(net279),
    .C(net261),
    .A(net280),
    .Y(_1793_),
    .D(_1767_));
 sg13g2_a22oi_1 _6589_ (.Y(_1794_),
    .B1(_1792_),
    .B2(_1793_),
    .A2(_1710_),
    .A1(_1708_));
 sg13g2_inv_1 _6590_ (.Y(_1795_),
    .A(_1794_));
 sg13g2_inv_1 _6591_ (.Y(_1796_),
    .A(_3389_));
 sg13g2_a21oi_1 _6592_ (.A1(_1674_),
    .A2(net136),
    .Y(_1797_),
    .B1(net261));
 sg13g2_and2_1 _6593_ (.A(_3805_),
    .B(_3473_),
    .X(_1798_));
 sg13g2_o21ai_1 _6594_ (.B1(_1722_),
    .Y(_1799_),
    .A1(net134),
    .A2(_1798_));
 sg13g2_o21ai_1 _6595_ (.B1(_1799_),
    .Y(_1800_),
    .A1(_1796_),
    .A2(_1797_));
 sg13g2_buf_1 _6596_ (.A(_1800_),
    .X(_1801_));
 sg13g2_a22oi_1 _6597_ (.Y(_1802_),
    .B1(_1792_),
    .B2(_1793_),
    .A2(_1716_),
    .A1(_1714_));
 sg13g2_nor2_1 _6598_ (.A(_1801_),
    .B(_1802_),
    .Y(_1803_));
 sg13g2_o21ai_1 _6599_ (.B1(_1803_),
    .Y(_1804_),
    .A1(_1617_),
    .A2(_1795_));
 sg13g2_xor2_1 _6600_ (.B(net133),
    .A(net261),
    .X(_1805_));
 sg13g2_xnor2_1 _6601_ (.Y(_1806_),
    .A(_1804_),
    .B(_1805_));
 sg13g2_nor2_1 _6602_ (.A(_1416_),
    .B(net260),
    .Y(_1807_));
 sg13g2_a21oi_1 _6603_ (.A1(net33),
    .A2(_1806_),
    .Y(_1808_),
    .B1(_1807_));
 sg13g2_nand2_1 _6604_ (.Y(_1809_),
    .A(net62),
    .B(_1808_));
 sg13g2_a22oi_1 _6605_ (.Y(_1810_),
    .B1(_1683_),
    .B2(net133),
    .A2(_1680_),
    .A1(net264));
 sg13g2_a21oi_1 _6606_ (.A1(_1809_),
    .A2(_1810_),
    .Y(_0048_),
    .B1(_1747_));
 sg13g2_nand4_1 _6607_ (.B(_1686_),
    .C(net261),
    .A(net135),
    .Y(_1811_),
    .D(_3409_));
 sg13g2_nand4_1 _6608_ (.B(_1685_),
    .C(net133),
    .A(_1752_),
    .Y(_1812_),
    .D(_1783_));
 sg13g2_nand2_2 _6609_ (.Y(_1813_),
    .A(_1811_),
    .B(_1812_));
 sg13g2_nand2_2 _6610_ (.Y(_1814_),
    .A(_1732_),
    .B(_1813_));
 sg13g2_a21oi_1 _6611_ (.A1(net134),
    .A2(net133),
    .Y(_1815_),
    .B1(_1798_));
 sg13g2_o21ai_1 _6612_ (.B1(net261),
    .Y(_1816_),
    .A1(net134),
    .A2(net133));
 sg13g2_o21ai_1 _6613_ (.B1(_1816_),
    .Y(_1817_),
    .A1(_1752_),
    .A2(_1815_));
 sg13g2_a21oi_1 _6614_ (.A1(_1736_),
    .A2(_1813_),
    .Y(_1818_),
    .B1(_1817_));
 sg13g2_o21ai_1 _6615_ (.B1(_1818_),
    .Y(_1819_),
    .A1(_1648_),
    .A2(_1814_));
 sg13g2_nor2b_1 _6616_ (.A(_3489_),
    .B_N(_3399_),
    .Y(_1820_));
 sg13g2_buf_2 _6617_ (.A(_1820_),
    .X(_1821_));
 sg13g2_nor2b_1 _6618_ (.A(_3399_),
    .B_N(_3489_),
    .Y(_1822_));
 sg13g2_nor2_1 _6619_ (.A(_1821_),
    .B(_1822_),
    .Y(_1823_));
 sg13g2_xor2_1 _6620_ (.B(_1823_),
    .A(_1819_),
    .X(_1824_));
 sg13g2_buf_1 _6621_ (.A(_0692_),
    .X(_1825_));
 sg13g2_nor2_1 _6622_ (.A(net32),
    .B(net211),
    .Y(_1826_));
 sg13g2_a21oi_1 _6623_ (.A1(net33),
    .A2(_1824_),
    .Y(_1827_),
    .B1(_1826_));
 sg13g2_nand2_1 _6624_ (.Y(_1828_),
    .A(net62),
    .B(_1827_));
 sg13g2_a22oi_1 _6625_ (.Y(_1829_),
    .B1(_1683_),
    .B2(net260),
    .A2(_1680_),
    .A1(net263));
 sg13g2_a21oi_1 _6626_ (.A1(_1828_),
    .A2(_1829_),
    .Y(_0049_),
    .B1(_1747_));
 sg13g2_xor2_1 _6627_ (.B(_0303_),
    .A(net300),
    .X(_1830_));
 sg13g2_xnor2_1 _6628_ (.Y(_1831_),
    .A(_1022_),
    .B(_1830_));
 sg13g2_nor2_1 _6629_ (.A(net38),
    .B(net180),
    .Y(_1832_));
 sg13g2_a21oi_1 _6630_ (.A1(net39),
    .A2(_1831_),
    .Y(_1833_),
    .B1(_1832_));
 sg13g2_nor2_1 _6631_ (.A(net65),
    .B(_1833_),
    .Y(_1834_));
 sg13g2_nor2_1 _6632_ (.A(_0275_),
    .B(net63),
    .Y(_1835_));
 sg13g2_a221oi_1 _6633_ (.B2(net18),
    .C1(net76),
    .B1(_1835_),
    .A1(_1422_),
    .Y(_1836_),
    .A2(net63));
 sg13g2_nor3_1 _6634_ (.A(net99),
    .B(_1834_),
    .C(_1836_),
    .Y(_0050_));
 sg13g2_nand2_1 _6635_ (.Y(_1837_),
    .A(_1784_),
    .B(_1822_));
 sg13g2_nand3_1 _6636_ (.B(_1783_),
    .C(_1821_),
    .A(_1752_),
    .Y(_1838_));
 sg13g2_o21ai_1 _6637_ (.B1(_1838_),
    .Y(_1839_),
    .A1(_1752_),
    .A2(_1837_));
 sg13g2_buf_1 _6638_ (.A(_1839_),
    .X(_1840_));
 sg13g2_o21ai_1 _6639_ (.B1(net135),
    .Y(_1841_),
    .A1(_3902_),
    .A2(_1651_));
 sg13g2_a21oi_1 _6640_ (.A1(_1686_),
    .A2(_1841_),
    .Y(_1842_),
    .B1(_1757_));
 sg13g2_and2_1 _6641_ (.A(_1840_),
    .B(_1842_),
    .X(_1843_));
 sg13g2_inv_1 _6642_ (.Y(_1844_),
    .A(_1670_));
 sg13g2_o21ai_1 _6643_ (.B1(_1844_),
    .Y(_1845_),
    .A1(_3807_),
    .A2(_3905_));
 sg13g2_inv_1 _6644_ (.Y(_1846_),
    .A(_3473_));
 sg13g2_a21oi_1 _6645_ (.A1(_1741_),
    .A2(net260),
    .Y(_1847_),
    .B1(_3399_));
 sg13g2_a21oi_1 _6646_ (.A1(_3904_),
    .A2(net322),
    .Y(_1848_),
    .B1(net260));
 sg13g2_nand2b_1 _6647_ (.Y(_1849_),
    .B(net133),
    .A_N(_1848_));
 sg13g2_o21ai_1 _6648_ (.B1(_1849_),
    .Y(_1850_),
    .A1(_1846_),
    .A2(_1847_));
 sg13g2_a21oi_1 _6649_ (.A1(_1843_),
    .A2(_1845_),
    .Y(_1851_),
    .B1(_1850_));
 sg13g2_nor3_1 _6650_ (.A(_1220_),
    .B(_4103_),
    .C(_1213_),
    .Y(_1852_));
 sg13g2_and3_1 _6651_ (.X(_1853_),
    .A(_1664_),
    .B(_1750_),
    .C(_1840_));
 sg13g2_and2_1 _6652_ (.A(_1852_),
    .B(_1853_),
    .X(_1854_));
 sg13g2_o21ai_1 _6653_ (.B1(_1854_),
    .Y(_1855_),
    .A1(_4163_),
    .A2(_0338_));
 sg13g2_o21ai_1 _6654_ (.B1(_1853_),
    .Y(_1856_),
    .A1(_1214_),
    .A2(_1218_));
 sg13g2_nand3_1 _6655_ (.B(_1855_),
    .C(_1856_),
    .A(_1851_),
    .Y(_1857_));
 sg13g2_buf_2 _6656_ (.A(_1857_),
    .X(_1858_));
 sg13g2_xor2_1 _6657_ (.B(net211),
    .A(_3500_),
    .X(_1859_));
 sg13g2_xnor2_1 _6658_ (.Y(_1860_),
    .A(_1858_),
    .B(_1859_));
 sg13g2_nor2_1 _6659_ (.A(net32),
    .B(net212),
    .Y(_1861_));
 sg13g2_a21oi_1 _6660_ (.A1(net33),
    .A2(_1860_),
    .Y(_1862_),
    .B1(_1861_));
 sg13g2_nand2_1 _6661_ (.Y(_1863_),
    .A(_1657_),
    .B(_1862_));
 sg13g2_nand3_1 _6662_ (.B(net329),
    .C(net272),
    .A(_3978_),
    .Y(_1864_));
 sg13g2_buf_1 _6663_ (.A(_1864_),
    .X(_1865_));
 sg13g2_inv_1 _6664_ (.Y(_1866_),
    .A(_1865_));
 sg13g2_a21oi_1 _6665_ (.A1(net66),
    .A2(_1866_),
    .Y(_1867_),
    .B1(net203));
 sg13g2_buf_2 _6666_ (.A(_1867_),
    .X(_1868_));
 sg13g2_nor2_1 _6667_ (.A(_1237_),
    .B(_1865_),
    .Y(_1869_));
 sg13g2_buf_2 _6668_ (.A(_1869_),
    .X(_1870_));
 sg13g2_a22oi_1 _6669_ (.Y(_1871_),
    .B1(_1870_),
    .B2(_1234_),
    .A2(_1868_),
    .A1(net211));
 sg13g2_a21oi_1 _6670_ (.A1(_1863_),
    .A2(_1871_),
    .Y(_0051_),
    .B1(_1747_));
 sg13g2_nand3_1 _6671_ (.B(_1783_),
    .C(_1821_),
    .A(_3936_),
    .Y(_1872_));
 sg13g2_o21ai_1 _6672_ (.B1(_1872_),
    .Y(_1873_),
    .A1(_3936_),
    .A2(_1837_));
 sg13g2_buf_1 _6673_ (.A(_1873_),
    .X(_1874_));
 sg13g2_nand3_1 _6674_ (.B(_1770_),
    .C(_1874_),
    .A(_1522_),
    .Y(_1875_));
 sg13g2_nor3_1 _6675_ (.A(_1771_),
    .B(_1772_),
    .C(_1777_),
    .Y(_1876_));
 sg13g2_and2_1 _6676_ (.A(_1874_),
    .B(_1876_),
    .X(_1877_));
 sg13g2_a21oi_1 _6677_ (.A1(_1796_),
    .A2(_3807_),
    .Y(_1878_),
    .B1(_1754_));
 sg13g2_or3_1 _6678_ (.A(_1690_),
    .B(_1695_),
    .C(_1878_),
    .X(_1879_));
 sg13g2_a22oi_1 _6679_ (.Y(_1880_),
    .B1(net133),
    .B2(net211),
    .A2(net260),
    .A1(_1741_));
 sg13g2_o21ai_1 _6680_ (.B1(net260),
    .Y(_1881_),
    .A1(_1787_),
    .A2(net211));
 sg13g2_o21ai_1 _6681_ (.B1(_1881_),
    .Y(_1882_),
    .A1(_1846_),
    .A2(_1880_));
 sg13g2_a21oi_1 _6682_ (.A1(_1877_),
    .A2(_1879_),
    .Y(_1883_),
    .B1(_1882_));
 sg13g2_o21ai_1 _6683_ (.B1(_1883_),
    .Y(_1884_),
    .A1(_1316_),
    .A2(_1875_));
 sg13g2_nor2b_1 _6684_ (.A(_3934_),
    .B_N(_3936_),
    .Y(_1885_));
 sg13g2_buf_2 _6685_ (.A(_1885_),
    .X(_1886_));
 sg13g2_nor2b_1 _6686_ (.A(_3936_),
    .B_N(_3934_),
    .Y(_1887_));
 sg13g2_buf_2 _6687_ (.A(_1887_),
    .X(_1888_));
 sg13g2_nor2_1 _6688_ (.A(_1886_),
    .B(_1888_),
    .Y(_1889_));
 sg13g2_xor2_1 _6689_ (.B(_1889_),
    .A(_1884_),
    .X(_1890_));
 sg13g2_buf_1 _6690_ (.A(_3599_),
    .X(_1891_));
 sg13g2_nor2_1 _6691_ (.A(net32),
    .B(net132),
    .Y(_1892_));
 sg13g2_a21oi_1 _6692_ (.A1(net33),
    .A2(_1890_),
    .Y(_1893_),
    .B1(_1892_));
 sg13g2_nand2_1 _6693_ (.Y(_1894_),
    .A(_1657_),
    .B(_1893_));
 sg13g2_a22oi_1 _6694_ (.Y(_1895_),
    .B1(_1870_),
    .B2(_1324_),
    .A2(_1868_),
    .A1(_3935_));
 sg13g2_a21oi_1 _6695_ (.A1(_1894_),
    .A2(_1895_),
    .Y(_0052_),
    .B1(_1747_));
 sg13g2_buf_1 _6696_ (.A(net80),
    .X(_1896_));
 sg13g2_nand2_1 _6697_ (.Y(_1897_),
    .A(_1792_),
    .B(_1793_));
 sg13g2_nand3_1 _6698_ (.B(_1821_),
    .C(_1886_),
    .A(_1846_),
    .Y(_1898_));
 sg13g2_nand3_1 _6699_ (.B(_1822_),
    .C(_1888_),
    .A(net261),
    .Y(_1899_));
 sg13g2_nand2_1 _6700_ (.Y(_1900_),
    .A(_1898_),
    .B(_1899_));
 sg13g2_nand2_1 _6701_ (.Y(_1901_),
    .A(_1897_),
    .B(_1900_));
 sg13g2_inv_1 _6702_ (.Y(_1902_),
    .A(_1901_));
 sg13g2_a21oi_1 _6703_ (.A1(_3481_),
    .A2(_3399_),
    .Y(_1903_),
    .B1(_3934_));
 sg13g2_nand2b_1 _6704_ (.Y(_1904_),
    .B(net211),
    .A_N(_1903_));
 sg13g2_a21oi_1 _6705_ (.A1(_3399_),
    .A2(_3934_),
    .Y(_1905_),
    .B1(_3936_));
 sg13g2_nand2b_1 _6706_ (.Y(_1906_),
    .B(net260),
    .A_N(_1905_));
 sg13g2_nand2_1 _6707_ (.Y(_1907_),
    .A(_1904_),
    .B(_1906_));
 sg13g2_a21oi_1 _6708_ (.A1(_1801_),
    .A2(_1900_),
    .Y(_1908_),
    .B1(_1907_));
 sg13g2_inv_1 _6709_ (.Y(_1909_),
    .A(_1908_));
 sg13g2_a21oi_1 _6710_ (.A1(_1719_),
    .A2(_1902_),
    .Y(_1910_),
    .B1(_1909_));
 sg13g2_xnor2_1 _6711_ (.Y(_1911_),
    .A(net212),
    .B(net132));
 sg13g2_xnor2_1 _6712_ (.Y(_1912_),
    .A(_1910_),
    .B(_1911_));
 sg13g2_buf_1 _6713_ (.A(_3419_),
    .X(_1913_));
 sg13g2_nor2_1 _6714_ (.A(net32),
    .B(_1913_),
    .Y(_1914_));
 sg13g2_a21oi_1 _6715_ (.A1(_1705_),
    .A2(_1912_),
    .Y(_1915_),
    .B1(_1914_));
 sg13g2_nand2_1 _6716_ (.Y(_1916_),
    .A(net61),
    .B(_1915_));
 sg13g2_a22oi_1 _6717_ (.Y(_1917_),
    .B1(_1870_),
    .B2(_1348_),
    .A2(_1868_),
    .A1(_1891_));
 sg13g2_a21oi_1 _6718_ (.A1(_1916_),
    .A2(_1917_),
    .Y(_0053_),
    .B1(_1747_));
 sg13g2_buf_1 _6719_ (.A(_3610_),
    .X(_1918_));
 sg13g2_inv_1 _6720_ (.Y(_1919_),
    .A(net130));
 sg13g2_nand3_1 _6721_ (.B(_1821_),
    .C(_1886_),
    .A(net132),
    .Y(_1920_));
 sg13g2_inv_1 _6722_ (.Y(_1921_),
    .A(_3599_));
 sg13g2_nand3_1 _6723_ (.B(_1822_),
    .C(_1888_),
    .A(_1921_),
    .Y(_1922_));
 sg13g2_nand2_2 _6724_ (.Y(_1923_),
    .A(_1920_),
    .B(_1922_));
 sg13g2_nand2_1 _6725_ (.Y(_1924_),
    .A(_1813_),
    .B(_1923_));
 sg13g2_or2_1 _6726_ (.X(_1925_),
    .B(_1924_),
    .A(_1733_));
 sg13g2_buf_1 _6727_ (.A(_1925_),
    .X(_1926_));
 sg13g2_inv_1 _6728_ (.Y(_1927_),
    .A(_1813_));
 sg13g2_inv_1 _6729_ (.Y(_1928_),
    .A(_1817_));
 sg13g2_o21ai_1 _6730_ (.B1(_1928_),
    .Y(_1929_),
    .A1(_1737_),
    .A2(_1927_));
 sg13g2_inv_1 _6731_ (.Y(_1930_),
    .A(_3489_));
 sg13g2_a22oi_1 _6732_ (.Y(_1931_),
    .B1(net211),
    .B2(net132),
    .A2(net212),
    .A1(_1787_));
 sg13g2_o21ai_1 _6733_ (.B1(net212),
    .Y(_1932_),
    .A1(_3937_),
    .A2(net132));
 sg13g2_o21ai_1 _6734_ (.B1(_1932_),
    .Y(_1933_),
    .A1(_1930_),
    .A2(_1931_));
 sg13g2_a21oi_1 _6735_ (.A1(_1923_),
    .A2(_1929_),
    .Y(_1934_),
    .B1(_1933_));
 sg13g2_o21ai_1 _6736_ (.B1(_1934_),
    .Y(_1935_),
    .A1(_1413_),
    .A2(_1926_));
 sg13g2_xnor2_1 _6737_ (.Y(_1936_),
    .A(net131),
    .B(net132));
 sg13g2_xnor2_1 _6738_ (.Y(_1937_),
    .A(_1935_),
    .B(_1936_));
 sg13g2_nand2_1 _6739_ (.Y(_1938_),
    .A(net34),
    .B(_1937_));
 sg13g2_o21ai_1 _6740_ (.B1(_1938_),
    .Y(_1939_),
    .A1(net42),
    .A2(_1919_));
 sg13g2_nand2_1 _6741_ (.Y(_1940_),
    .A(net61),
    .B(_1939_));
 sg13g2_a22oi_1 _6742_ (.Y(_1941_),
    .B1(_1870_),
    .B2(_1422_),
    .A2(_1868_),
    .A1(_1913_));
 sg13g2_a21oi_1 _6743_ (.A1(_1940_),
    .A2(_1941_),
    .Y(_0054_),
    .B1(_1747_));
 sg13g2_nand4_1 _6744_ (.B(_3419_),
    .C(_1921_),
    .A(_3489_),
    .Y(_1942_),
    .D(_1888_));
 sg13g2_inv_1 _6745_ (.Y(_1943_),
    .A(_3419_));
 sg13g2_nand4_1 _6746_ (.B(_1943_),
    .C(_3599_),
    .A(_1930_),
    .Y(_1944_),
    .D(_1886_));
 sg13g2_nand2_1 _6747_ (.Y(_1945_),
    .A(_1942_),
    .B(_1944_));
 sg13g2_nand2_1 _6748_ (.Y(_1946_),
    .A(_1840_),
    .B(_1945_));
 sg13g2_a21o_1 _6749_ (.A2(_3419_),
    .A1(_3936_),
    .B1(_3599_),
    .X(_1947_));
 sg13g2_a21o_1 _6750_ (.A2(_3936_),
    .A1(_3500_),
    .B1(net131),
    .X(_1948_));
 sg13g2_a22oi_1 _6751_ (.Y(_1949_),
    .B1(_1948_),
    .B2(net132),
    .A2(_1947_),
    .A1(net212));
 sg13g2_inv_1 _6752_ (.Y(_1950_),
    .A(_1949_));
 sg13g2_a21oi_1 _6753_ (.A1(_1850_),
    .A2(_1945_),
    .Y(_1951_),
    .B1(_1950_));
 sg13g2_o21ai_1 _6754_ (.B1(_1951_),
    .Y(_1952_),
    .A1(_1759_),
    .A2(_1946_));
 sg13g2_xor2_1 _6755_ (.B(_1918_),
    .A(net131),
    .X(_1953_));
 sg13g2_xnor2_1 _6756_ (.Y(_1954_),
    .A(_1952_),
    .B(_1953_));
 sg13g2_buf_1 _6757_ (.A(_3429_),
    .X(_1955_));
 sg13g2_nor2_1 _6758_ (.A(net32),
    .B(net129),
    .Y(_1956_));
 sg13g2_a21oi_1 _6759_ (.A1(_1705_),
    .A2(_1954_),
    .Y(_1957_),
    .B1(_1956_));
 sg13g2_nand2_1 _6760_ (.Y(_1958_),
    .A(net61),
    .B(_1957_));
 sg13g2_a22oi_1 _6761_ (.Y(_1959_),
    .B1(_1870_),
    .B2(_1487_),
    .A2(_1868_),
    .A1(net130));
 sg13g2_a21oi_1 _6762_ (.A1(_1958_),
    .A2(_1959_),
    .Y(_0055_),
    .B1(_1747_));
 sg13g2_buf_1 _6763_ (.A(net51),
    .X(_1960_));
 sg13g2_and2_1 _6764_ (.A(_3599_),
    .B(_3610_),
    .X(_1961_));
 sg13g2_nand3_1 _6765_ (.B(_1886_),
    .C(_1961_),
    .A(_1943_),
    .Y(_1962_));
 sg13g2_nand3_1 _6766_ (.B(_3621_),
    .C(_1888_),
    .A(net131),
    .Y(_1963_));
 sg13g2_nand2_1 _6767_ (.Y(_1964_),
    .A(_1962_),
    .B(_1963_));
 sg13g2_and2_1 _6768_ (.A(_1874_),
    .B(_1964_),
    .X(_1965_));
 sg13g2_inv_1 _6769_ (.Y(_1966_),
    .A(_1882_));
 sg13g2_and2_1 _6770_ (.A(_1962_),
    .B(_1963_),
    .X(_1967_));
 sg13g2_buf_1 _6771_ (.A(_1967_),
    .X(_1968_));
 sg13g2_inv_1 _6772_ (.Y(_1969_),
    .A(_3621_));
 sg13g2_a22oi_1 _6773_ (.Y(_1970_),
    .B1(net132),
    .B2(net130),
    .A2(net131),
    .A1(_3937_));
 sg13g2_inv_1 _6774_ (.Y(_1971_),
    .A(_1970_));
 sg13g2_a22oi_1 _6775_ (.Y(_1972_),
    .B1(_1971_),
    .B2(net212),
    .A2(_1969_),
    .A1(net131));
 sg13g2_o21ai_1 _6776_ (.B1(_1972_),
    .Y(_1973_),
    .A1(_1966_),
    .A2(_1968_));
 sg13g2_a21oi_1 _6777_ (.A1(_1780_),
    .A2(_1965_),
    .Y(_1974_),
    .B1(_1973_));
 sg13g2_nand4_1 _6778_ (.B(_1770_),
    .C(_1874_),
    .A(_1532_),
    .Y(_1975_),
    .D(_1964_));
 sg13g2_and2_1 _6779_ (.A(_1974_),
    .B(_1975_),
    .X(_1976_));
 sg13g2_xnor2_1 _6780_ (.Y(_1977_),
    .A(net129),
    .B(net130));
 sg13g2_xnor2_1 _6781_ (.Y(_1978_),
    .A(_1976_),
    .B(_1977_));
 sg13g2_nor2_1 _6782_ (.A(_1825_),
    .B(net209),
    .Y(_1979_));
 sg13g2_a21oi_1 _6783_ (.A1(_1960_),
    .A2(_1978_),
    .Y(_1980_),
    .B1(_1979_));
 sg13g2_nand2_1 _6784_ (.Y(_1981_),
    .A(_1896_),
    .B(_1980_));
 sg13g2_a22oi_1 _6785_ (.Y(_1982_),
    .B1(_1870_),
    .B2(_0699_),
    .A2(_1868_),
    .A1(_1955_));
 sg13g2_buf_1 _6786_ (.A(net204),
    .X(_1983_));
 sg13g2_a21oi_1 _6787_ (.A1(_1981_),
    .A2(_1982_),
    .Y(_0056_),
    .B1(net93));
 sg13g2_inv_1 _6788_ (.Y(_1984_),
    .A(_1804_));
 sg13g2_nand4_1 _6789_ (.B(net131),
    .C(net129),
    .A(net212),
    .Y(_1985_),
    .D(_3621_));
 sg13g2_nand3b_1 _6790_ (.B(_3438_),
    .C(_1961_),
    .Y(_1986_),
    .A_N(_3934_));
 sg13g2_buf_1 _6791_ (.A(_1986_),
    .X(_1987_));
 sg13g2_nand2_1 _6792_ (.Y(_1988_),
    .A(_1985_),
    .B(_1987_));
 sg13g2_nand2_1 _6793_ (.Y(_1989_),
    .A(_1900_),
    .B(_1988_));
 sg13g2_a21oi_1 _6794_ (.A1(_3935_),
    .A2(_3599_),
    .Y(_1990_),
    .B1(net129));
 sg13g2_and2_1 _6795_ (.A(_3599_),
    .B(_3429_),
    .X(_1991_));
 sg13g2_o21ai_1 _6796_ (.B1(net131),
    .Y(_1992_),
    .A1(net130),
    .A2(_1991_));
 sg13g2_o21ai_1 _6797_ (.B1(_1992_),
    .Y(_1993_),
    .A1(_1919_),
    .A2(_1990_));
 sg13g2_buf_1 _6798_ (.A(_1993_),
    .X(_1994_));
 sg13g2_a22oi_1 _6799_ (.Y(_1995_),
    .B1(_1985_),
    .B2(_1987_),
    .A2(_1906_),
    .A1(_1904_));
 sg13g2_nor2_1 _6800_ (.A(_1994_),
    .B(_1995_),
    .Y(_1996_));
 sg13g2_o21ai_1 _6801_ (.B1(_1996_),
    .Y(_1997_),
    .A1(_1984_),
    .A2(_1989_));
 sg13g2_xnor2_1 _6802_ (.Y(_1998_),
    .A(net129),
    .B(net209));
 sg13g2_xnor2_1 _6803_ (.Y(_1999_),
    .A(_1997_),
    .B(_1998_));
 sg13g2_inv_2 _6804_ (.Y(_2000_),
    .A(net210));
 sg13g2_nor2_1 _6805_ (.A(_1199_),
    .B(_2000_),
    .Y(_2001_));
 sg13g2_a21oi_1 _6806_ (.A1(net41),
    .A2(_1999_),
    .Y(_2002_),
    .B1(_2001_));
 sg13g2_a22oi_1 _6807_ (.Y(_2003_),
    .B1(_1870_),
    .B2(net325),
    .A2(_1868_),
    .A1(net209));
 sg13g2_nand2b_1 _6808_ (.Y(_2004_),
    .B(net270),
    .A_N(_2003_));
 sg13g2_o21ai_1 _6809_ (.B1(_2004_),
    .Y(_0057_),
    .A1(_0393_),
    .A2(_2002_));
 sg13g2_nor2b_1 _6810_ (.A(_3610_),
    .B_N(_3429_),
    .Y(_2005_));
 sg13g2_nand3_1 _6811_ (.B(_1921_),
    .C(_2005_),
    .A(_3419_),
    .Y(_2006_));
 sg13g2_and2_1 _6812_ (.A(_3610_),
    .B(_3940_),
    .X(_2007_));
 sg13g2_buf_1 _6813_ (.A(_2007_),
    .X(_2008_));
 sg13g2_nand3_1 _6814_ (.B(_3438_),
    .C(_2008_),
    .A(_1891_),
    .Y(_2009_));
 sg13g2_o21ai_1 _6815_ (.B1(_2009_),
    .Y(_2010_),
    .A1(net209),
    .A2(_2006_));
 sg13g2_buf_1 _6816_ (.A(_2010_),
    .X(_2011_));
 sg13g2_nor2_1 _6817_ (.A(_1991_),
    .B(_2008_),
    .Y(_2012_));
 sg13g2_o21ai_1 _6818_ (.B1(net129),
    .Y(_2013_),
    .A1(net130),
    .A2(net209));
 sg13g2_o21ai_1 _6819_ (.B1(_2013_),
    .Y(_2014_),
    .A1(_1943_),
    .A2(_2012_));
 sg13g2_a21o_1 _6820_ (.A2(_2011_),
    .A1(_1933_),
    .B1(_2014_),
    .X(_2015_));
 sg13g2_nand2_2 _6821_ (.Y(_2016_),
    .A(_1923_),
    .B(_2011_));
 sg13g2_nor2b_1 _6822_ (.A(_2016_),
    .B_N(_1819_),
    .Y(_2017_));
 sg13g2_nor2_1 _6823_ (.A(_2015_),
    .B(_2017_),
    .Y(_2018_));
 sg13g2_xnor2_1 _6824_ (.Y(_2019_),
    .A(net210),
    .B(net209));
 sg13g2_xnor2_1 _6825_ (.Y(_2020_),
    .A(_2018_),
    .B(_2019_));
 sg13g2_buf_1 _6826_ (.A(_3723_),
    .X(_2021_));
 sg13g2_nor2_1 _6827_ (.A(_1825_),
    .B(net128),
    .Y(_2022_));
 sg13g2_a21oi_1 _6828_ (.A1(_1960_),
    .A2(_2020_),
    .Y(_2023_),
    .B1(_2022_));
 sg13g2_nand2_1 _6829_ (.Y(_2024_),
    .A(_1896_),
    .B(_2023_));
 sg13g2_a22oi_1 _6830_ (.Y(_2025_),
    .B1(_1870_),
    .B2(_1655_),
    .A2(_1868_),
    .A1(_3939_));
 sg13g2_a21oi_1 _6831_ (.A1(_2024_),
    .A2(_2025_),
    .Y(_0058_),
    .B1(net93));
 sg13g2_xnor2_1 _6832_ (.Y(_2026_),
    .A(net210),
    .B(net128));
 sg13g2_nor2b_1 _6833_ (.A(_3940_),
    .B_N(_3938_),
    .Y(_2027_));
 sg13g2_nand3_1 _6834_ (.B(_2005_),
    .C(_2027_),
    .A(_3419_),
    .Y(_2028_));
 sg13g2_nand3_1 _6835_ (.B(_3438_),
    .C(_2008_),
    .A(_2000_),
    .Y(_2029_));
 sg13g2_and2_1 _6836_ (.A(_2028_),
    .B(_2029_),
    .X(_2030_));
 sg13g2_buf_1 _6837_ (.A(_2030_),
    .X(_2031_));
 sg13g2_a21oi_1 _6838_ (.A1(_1942_),
    .A2(_1944_),
    .Y(_2032_),
    .B1(_2031_));
 sg13g2_a21o_1 _6839_ (.A2(net130),
    .A1(_3419_),
    .B1(net210),
    .X(_2033_));
 sg13g2_a21o_1 _6840_ (.A2(_3939_),
    .A1(net130),
    .B1(_3940_),
    .X(_2034_));
 sg13g2_a22oi_1 _6841_ (.Y(_2035_),
    .B1(_2034_),
    .B2(net129),
    .A2(_2033_),
    .A1(_3940_));
 sg13g2_o21ai_1 _6842_ (.B1(_2035_),
    .Y(_2036_),
    .A1(_1949_),
    .A2(_2031_));
 sg13g2_a21oi_1 _6843_ (.A1(_1858_),
    .A2(_2032_),
    .Y(_2037_),
    .B1(_2036_));
 sg13g2_xnor2_1 _6844_ (.Y(_2038_),
    .A(_2026_),
    .B(_2037_));
 sg13g2_nor2b_1 _6845_ (.A(net81),
    .B_N(_0015_),
    .Y(_2039_));
 sg13g2_a21oi_2 _6846_ (.B1(_2039_),
    .Y(_2040_),
    .A2(_2038_),
    .A1(net67));
 sg13g2_nand2_1 _6847_ (.Y(_2041_),
    .A(net106),
    .B(_2040_));
 sg13g2_nand2_1 _6848_ (.Y(_2042_),
    .A(_0384_),
    .B(net83));
 sg13g2_inv_1 _6849_ (.Y(_2043_),
    .A(_2042_));
 sg13g2_a21oi_1 _6850_ (.A1(net66),
    .A2(_2043_),
    .Y(_2044_),
    .B1(net203));
 sg13g2_buf_2 _6851_ (.A(_2044_),
    .X(_2045_));
 sg13g2_nand2_1 _6852_ (.Y(_2046_),
    .A(net328),
    .B(net83));
 sg13g2_nor3_1 _6853_ (.A(_3983_),
    .B(_2046_),
    .C(_1237_),
    .Y(_2047_));
 sg13g2_a21oi_1 _6854_ (.A1(net128),
    .A2(_2045_),
    .Y(_2048_),
    .B1(_2047_));
 sg13g2_a21oi_1 _6855_ (.A1(_2041_),
    .A2(_2048_),
    .Y(_0059_),
    .B1(net93));
 sg13g2_inv_1 _6856_ (.Y(_2049_),
    .A(_3429_));
 sg13g2_nor2b_1 _6857_ (.A(_3938_),
    .B_N(_3723_),
    .Y(_2050_));
 sg13g2_nand3_1 _6858_ (.B(_2008_),
    .C(_2050_),
    .A(_2049_),
    .Y(_2051_));
 sg13g2_inv_1 _6859_ (.Y(_2052_),
    .A(_3723_));
 sg13g2_nand3_1 _6860_ (.B(_2005_),
    .C(_2027_),
    .A(_2052_),
    .Y(_2053_));
 sg13g2_and2_1 _6861_ (.A(_2051_),
    .B(_2053_),
    .X(_2054_));
 sg13g2_buf_1 _6862_ (.A(_2054_),
    .X(_2055_));
 sg13g2_nand4_1 _6863_ (.B(_1522_),
    .C(_1770_),
    .A(_1314_),
    .Y(_2056_),
    .D(_1874_));
 sg13g2_or3_1 _6864_ (.A(_1968_),
    .B(_2055_),
    .C(_2056_),
    .X(_2057_));
 sg13g2_buf_1 _6865_ (.A(_3746_),
    .X(_2058_));
 sg13g2_xnor2_1 _6866_ (.Y(_2059_),
    .A(net127),
    .B(_2021_));
 sg13g2_nand2b_1 _6867_ (.Y(_2060_),
    .B(net202),
    .A_N(_2059_));
 sg13g2_or3_1 _6868_ (.A(_1310_),
    .B(_2057_),
    .C(_2060_),
    .X(_2061_));
 sg13g2_nor2_1 _6869_ (.A(_1968_),
    .B(_2055_),
    .Y(_2062_));
 sg13g2_o21ai_1 _6870_ (.B1(_1883_),
    .Y(_2063_),
    .A1(_1253_),
    .A2(_1875_));
 sg13g2_a22oi_1 _6871_ (.Y(_2064_),
    .B1(_3941_),
    .B2(net128),
    .A2(net210),
    .A1(_1918_));
 sg13g2_o21ai_1 _6872_ (.B1(net210),
    .Y(_2065_),
    .A1(_3941_),
    .A2(net128));
 sg13g2_o21ai_1 _6873_ (.B1(_2065_),
    .Y(_2066_),
    .A1(_2049_),
    .A2(_2064_));
 sg13g2_inv_1 _6874_ (.Y(_2067_),
    .A(_2066_));
 sg13g2_o21ai_1 _6875_ (.B1(_2067_),
    .Y(_2068_),
    .A1(_1972_),
    .A2(_2055_));
 sg13g2_a21oi_1 _6876_ (.A1(_2062_),
    .A2(_2063_),
    .Y(_2069_),
    .B1(_2068_));
 sg13g2_or2_1 _6877_ (.X(_2070_),
    .B(_2060_),
    .A(_2069_));
 sg13g2_nand4_1 _6878_ (.B(_2059_),
    .C(_2069_),
    .A(net103),
    .Y(_2071_),
    .D(_2057_));
 sg13g2_and3_1 _6879_ (.X(_2072_),
    .A(net103),
    .B(_2059_),
    .C(_2069_));
 sg13g2_a22oi_1 _6880_ (.Y(_2073_),
    .B1(_1310_),
    .B2(_2072_),
    .A2(_0014_),
    .A1(net113));
 sg13g2_nand4_1 _6881_ (.B(_2070_),
    .C(_2071_),
    .A(_2061_),
    .Y(_2074_),
    .D(_2073_));
 sg13g2_inv_1 _6882_ (.Y(_2075_),
    .A(_2074_));
 sg13g2_nand2_1 _6883_ (.Y(_2076_),
    .A(net106),
    .B(_2075_));
 sg13g2_nor2_1 _6884_ (.A(_1237_),
    .B(_2042_),
    .Y(_2077_));
 sg13g2_buf_2 _6885_ (.A(_2077_),
    .X(_2078_));
 sg13g2_a22oi_1 _6886_ (.Y(_2079_),
    .B1(_2078_),
    .B2(net274),
    .A2(_2045_),
    .A1(_2058_));
 sg13g2_a21oi_1 _6887_ (.A1(_2076_),
    .A2(_2079_),
    .Y(_0060_),
    .B1(net93));
 sg13g2_buf_1 _6888_ (.A(_3964_),
    .X(_2080_));
 sg13g2_nand2_1 _6889_ (.Y(_2081_),
    .A(net327),
    .B(_1551_));
 sg13g2_o21ai_1 _6890_ (.B1(_2081_),
    .Y(_2082_),
    .A1(_0454_),
    .A2(net63));
 sg13g2_nor2_1 _6891_ (.A(net82),
    .B(_2082_),
    .Y(_2083_));
 sg13g2_buf_1 _6892_ (.A(net77),
    .X(_2084_));
 sg13g2_xor2_1 _6893_ (.B(net180),
    .A(_3753_),
    .X(_2085_));
 sg13g2_xnor2_1 _6894_ (.Y(_2086_),
    .A(_0308_),
    .B(_2085_));
 sg13g2_nor2_1 _6895_ (.A(net34),
    .B(net250),
    .Y(_2087_));
 sg13g2_a21oi_1 _6896_ (.A1(net41),
    .A2(_2086_),
    .Y(_2088_),
    .B1(_2087_));
 sg13g2_nor2_1 _6897_ (.A(net60),
    .B(_2088_),
    .Y(_2089_));
 sg13g2_nor3_1 _6898_ (.A(net92),
    .B(_2083_),
    .C(_2089_),
    .Y(_0061_));
 sg13g2_buf_1 _6899_ (.A(net309),
    .X(_2090_));
 sg13g2_xor2_1 _6900_ (.B(net126),
    .A(_2058_),
    .X(_2091_));
 sg13g2_and2_1 _6901_ (.A(_0904_),
    .B(_0905_),
    .X(_2092_));
 sg13g2_buf_1 _6902_ (.A(_2092_),
    .X(_2093_));
 sg13g2_nor3_1 _6903_ (.A(_2093_),
    .B(_0902_),
    .C(_0924_),
    .Y(_2094_));
 sg13g2_or3_1 _6904_ (.A(_2093_),
    .B(_0924_),
    .C(_0958_),
    .X(_2095_));
 sg13g2_o21ai_1 _6905_ (.B1(_2095_),
    .Y(_2096_),
    .A1(_2093_),
    .A2(_0945_));
 sg13g2_a21o_1 _6906_ (.A2(_2094_),
    .A1(_0893_),
    .B1(_2096_),
    .X(_2097_));
 sg13g2_nand2_1 _6907_ (.Y(_2098_),
    .A(_2049_),
    .B(_2050_));
 sg13g2_inv_1 _6908_ (.Y(_2099_),
    .A(_3746_));
 sg13g2_nand2_1 _6909_ (.Y(_2100_),
    .A(_3940_),
    .B(_2099_));
 sg13g2_nor2b_1 _6910_ (.A(_3723_),
    .B_N(_3746_),
    .Y(_2101_));
 sg13g2_nand3_1 _6911_ (.B(_2027_),
    .C(_2101_),
    .A(_1955_),
    .Y(_2102_));
 sg13g2_o21ai_1 _6912_ (.B1(_2102_),
    .Y(_2103_),
    .A1(_2098_),
    .A2(_2100_));
 sg13g2_buf_1 _6913_ (.A(_2103_),
    .X(_2104_));
 sg13g2_nand2_1 _6914_ (.Y(_2105_),
    .A(_1988_),
    .B(_2104_));
 sg13g2_a21oi_1 _6915_ (.A1(_0736_),
    .A2(_1333_),
    .Y(_2106_),
    .B1(_1338_));
 sg13g2_o21ai_1 _6916_ (.B1(_1718_),
    .Y(_2107_),
    .A1(_1712_),
    .A2(_2106_));
 sg13g2_a21oi_1 _6917_ (.A1(_1902_),
    .A2(_2107_),
    .Y(_2108_),
    .B1(_1909_));
 sg13g2_a21oi_1 _6918_ (.A1(_3940_),
    .A2(_3746_),
    .Y(_2109_),
    .B1(_3723_));
 sg13g2_a21oi_1 _6919_ (.A1(net129),
    .A2(_3940_),
    .Y(_2110_),
    .B1(_3746_));
 sg13g2_nand2b_1 _6920_ (.Y(_2111_),
    .B(_2021_),
    .A_N(_2110_));
 sg13g2_o21ai_1 _6921_ (.B1(_2111_),
    .Y(_2112_),
    .A1(_2000_),
    .A2(_2109_));
 sg13g2_buf_1 _6922_ (.A(_2112_),
    .X(_2113_));
 sg13g2_a21oi_1 _6923_ (.A1(_1994_),
    .A2(_2104_),
    .Y(_2114_),
    .B1(_2113_));
 sg13g2_o21ai_1 _6924_ (.B1(_2114_),
    .Y(_2115_),
    .A1(_2105_),
    .A2(_2108_));
 sg13g2_or3_1 _6925_ (.A(_0730_),
    .B(_0725_),
    .C(_2115_),
    .X(_2116_));
 sg13g2_nand2_1 _6926_ (.Y(_2117_),
    .A(_1333_),
    .B(_1606_));
 sg13g2_nor4_1 _6927_ (.A(_1712_),
    .B(_1901_),
    .C(_2105_),
    .D(_2117_),
    .Y(_2118_));
 sg13g2_or2_1 _6928_ (.X(_2119_),
    .B(_2118_),
    .A(_2115_));
 sg13g2_buf_1 _6929_ (.A(_2119_),
    .X(_2120_));
 sg13g2_o21ai_1 _6930_ (.B1(_2120_),
    .Y(_2121_),
    .A1(_2097_),
    .A2(_2116_));
 sg13g2_xnor2_1 _6931_ (.Y(_2122_),
    .A(_2091_),
    .B(_2121_));
 sg13g2_nand2_1 _6932_ (.Y(_2123_),
    .A(net67),
    .B(_2122_));
 sg13g2_or2_1 _6933_ (.X(_2124_),
    .B(_0013_),
    .A(_4029_));
 sg13g2_and2_1 _6934_ (.A(_2123_),
    .B(_2124_),
    .X(_2125_));
 sg13g2_nand2b_1 _6935_ (.Y(_2126_),
    .B(net100),
    .A_N(_2125_));
 sg13g2_a22oi_1 _6936_ (.Y(_2127_),
    .B1(_2078_),
    .B2(_1726_),
    .A2(_2045_),
    .A1(net126));
 sg13g2_a21oi_1 _6937_ (.A1(_2126_),
    .A2(_2127_),
    .Y(_0062_),
    .B1(_1983_));
 sg13g2_buf_1 _6938_ (.A(_3747_),
    .X(_2128_));
 sg13g2_xnor2_1 _6939_ (.Y(_2129_),
    .A(net125),
    .B(net126));
 sg13g2_nand2_1 _6940_ (.Y(_2130_),
    .A(net309),
    .B(_2050_));
 sg13g2_nand3_1 _6941_ (.B(_3725_),
    .C(_2027_),
    .A(_3746_),
    .Y(_2131_));
 sg13g2_o21ai_1 _6942_ (.B1(_2131_),
    .Y(_2132_),
    .A1(_2100_),
    .A2(_2130_));
 sg13g2_buf_2 _6943_ (.A(_2132_),
    .X(_2133_));
 sg13g2_nand2_1 _6944_ (.Y(_2134_),
    .A(_2011_),
    .B(_2133_));
 sg13g2_nor3_1 _6945_ (.A(_1381_),
    .B(_1926_),
    .C(_2134_),
    .Y(_2135_));
 sg13g2_nor2b_1 _6946_ (.A(_2129_),
    .B_N(_2135_),
    .Y(_2136_));
 sg13g2_nor2_1 _6947_ (.A(_1924_),
    .B(_2134_),
    .Y(_2137_));
 sg13g2_o21ai_1 _6948_ (.B1(_1737_),
    .Y(_2138_),
    .A1(_1411_),
    .A2(_1733_));
 sg13g2_a21o_1 _6949_ (.A2(_1923_),
    .A1(_1817_),
    .B1(_1933_),
    .X(_2139_));
 sg13g2_a21o_1 _6950_ (.A2(_2139_),
    .A1(_2011_),
    .B1(_2014_),
    .X(_2140_));
 sg13g2_a22oi_1 _6951_ (.Y(_2141_),
    .B1(net128),
    .B2(net126),
    .A2(net127),
    .A1(net209));
 sg13g2_o21ai_1 _6952_ (.B1(net127),
    .Y(_2142_),
    .A1(net128),
    .A2(net126));
 sg13g2_o21ai_1 _6953_ (.B1(_2142_),
    .Y(_2143_),
    .A1(_2000_),
    .A2(_2141_));
 sg13g2_buf_1 _6954_ (.A(_2143_),
    .X(_2144_));
 sg13g2_a221oi_1 _6955_ (.B2(_2133_),
    .C1(_2144_),
    .B1(_2140_),
    .A1(_2137_),
    .Y(_2145_),
    .A2(_2138_));
 sg13g2_nand2_1 _6956_ (.Y(_2146_),
    .A(_2129_),
    .B(_2145_));
 sg13g2_and2_1 _6957_ (.A(_1175_),
    .B(_0995_),
    .X(_2147_));
 sg13g2_nand2_1 _6958_ (.Y(_2148_),
    .A(_1394_),
    .B(_1103_));
 sg13g2_o21ai_1 _6959_ (.B1(_1396_),
    .Y(_2149_),
    .A1(_1372_),
    .A2(_2148_));
 sg13g2_a21o_1 _6960_ (.A2(_0995_),
    .A1(_1178_),
    .B1(_1398_),
    .X(_2150_));
 sg13g2_a21oi_1 _6961_ (.A1(_2147_),
    .A2(_2149_),
    .Y(_2151_),
    .B1(_2150_));
 sg13g2_nand2_1 _6962_ (.Y(_2152_),
    .A(_1390_),
    .B(_1392_));
 sg13g2_o21ai_1 _6963_ (.B1(_2152_),
    .Y(_2153_),
    .A1(_1385_),
    .A2(_2151_));
 sg13g2_nor2_1 _6964_ (.A(_2146_),
    .B(_2153_),
    .Y(_2154_));
 sg13g2_a21oi_1 _6965_ (.A1(_1360_),
    .A2(_1363_),
    .Y(_2155_),
    .B1(_1369_));
 sg13g2_o21ai_1 _6966_ (.B1(_1371_),
    .Y(_2156_),
    .A1(_1353_),
    .A2(_2155_));
 sg13g2_and2_1 _6967_ (.A(_1100_),
    .B(_1102_),
    .X(_2157_));
 sg13g2_nand3_1 _6968_ (.B(_0995_),
    .C(_1393_),
    .A(_1099_),
    .Y(_2158_));
 sg13g2_nor3_1 _6969_ (.A(_2157_),
    .B(_1350_),
    .C(_2158_),
    .Y(_2159_));
 sg13g2_nand2_1 _6970_ (.Y(_2160_),
    .A(_2156_),
    .B(_2159_));
 sg13g2_mux2_1 _6971_ (.A0(_2136_),
    .A1(_2154_),
    .S(_2160_),
    .X(_2161_));
 sg13g2_or2_1 _6972_ (.X(_2162_),
    .B(_0012_),
    .A(net103));
 sg13g2_nand2_1 _6973_ (.Y(_2163_),
    .A(_2135_),
    .B(_2153_));
 sg13g2_a21oi_1 _6974_ (.A1(_2145_),
    .A2(_2163_),
    .Y(_2164_),
    .B1(_2129_));
 sg13g2_o21ai_1 _6975_ (.B1(net103),
    .Y(_2165_),
    .A1(_2135_),
    .A2(_2146_));
 sg13g2_or2_1 _6976_ (.X(_2166_),
    .B(_2165_),
    .A(_2164_));
 sg13g2_a22oi_1 _6977_ (.Y(_2167_),
    .B1(_2162_),
    .B2(_2166_),
    .A2(_2161_),
    .A1(net81));
 sg13g2_nand2_1 _6978_ (.Y(_2168_),
    .A(net106),
    .B(_2167_));
 sg13g2_a22oi_1 _6979_ (.Y(_2169_),
    .B1(_2078_),
    .B2(_1745_),
    .A2(_2045_),
    .A1(_2128_));
 sg13g2_a21oi_1 _6980_ (.A1(_2168_),
    .A2(_2169_),
    .Y(_0063_),
    .B1(_1983_));
 sg13g2_nand3_1 _6981_ (.B(_3749_),
    .C(_2050_),
    .A(net309),
    .Y(_2170_));
 sg13g2_nor2b_1 _6982_ (.A(net309),
    .B_N(_3747_),
    .Y(_2171_));
 sg13g2_nand3_1 _6983_ (.B(_2101_),
    .C(_2171_),
    .A(net210),
    .Y(_2172_));
 sg13g2_a22oi_1 _6984_ (.Y(_2173_),
    .B1(_2170_),
    .B2(_2172_),
    .A2(_2029_),
    .A1(_2028_));
 sg13g2_and3_1 _6985_ (.X(_2174_),
    .A(_1840_),
    .B(_1945_),
    .C(_2173_));
 sg13g2_buf_1 _6986_ (.A(_2174_),
    .X(_2175_));
 sg13g2_and3_1 _6987_ (.X(_2176_),
    .A(_1437_),
    .B(_1751_),
    .C(_2175_));
 sg13g2_nand2b_1 _6988_ (.Y(_2177_),
    .B(_2176_),
    .A_N(_1222_));
 sg13g2_nand2_1 _6989_ (.Y(_2178_),
    .A(_1445_),
    .B(_1477_));
 sg13g2_nor3_1 _6990_ (.A(_1441_),
    .B(_1474_),
    .C(_2178_),
    .Y(_2179_));
 sg13g2_nand2_1 _6991_ (.Y(_2180_),
    .A(_1467_),
    .B(_1469_));
 sg13g2_nand2_1 _6992_ (.Y(_2181_),
    .A(_0308_),
    .B(_1470_));
 sg13g2_nand4_1 _6993_ (.B(_2180_),
    .C(_1464_),
    .A(_4184_),
    .Y(_2182_),
    .D(_2181_));
 sg13g2_buf_1 _6994_ (.A(_2182_),
    .X(_2183_));
 sg13g2_nand3b_1 _6995_ (.B(_2179_),
    .C(_2183_),
    .Y(_2184_),
    .A_N(_2177_));
 sg13g2_a221oi_1 _6996_ (.B2(_0226_),
    .C1(_0335_),
    .B1(_0225_),
    .A1(_4178_),
    .Y(_2185_),
    .A2(_1471_));
 sg13g2_o21ai_1 _6997_ (.B1(_1445_),
    .Y(_2186_),
    .A1(_1453_),
    .A2(_2185_));
 sg13g2_and3_1 _6998_ (.X(_2187_),
    .A(_1454_),
    .B(_1455_),
    .C(_2186_));
 sg13g2_or3_1 _6999_ (.A(_1441_),
    .B(_2187_),
    .C(_2177_),
    .X(_2188_));
 sg13g2_xor2_1 _7000_ (.B(net297),
    .A(net125),
    .X(_2189_));
 sg13g2_nand2_1 _7001_ (.Y(_2190_),
    .A(net202),
    .B(_2189_));
 sg13g2_a21oi_1 _7002_ (.A1(_2184_),
    .A2(_2188_),
    .Y(_2191_),
    .B1(_2190_));
 sg13g2_nand2b_1 _7003_ (.Y(_2192_),
    .B(_1750_),
    .A_N(_1663_));
 sg13g2_nor2_1 _7004_ (.A(_1431_),
    .B(_2192_),
    .Y(_2193_));
 sg13g2_nand2b_1 _7005_ (.Y(_2194_),
    .B(_1951_),
    .A_N(_1758_));
 sg13g2_nand2_1 _7006_ (.Y(_2195_),
    .A(_2170_),
    .B(_2172_));
 sg13g2_nand2b_1 _7007_ (.Y(_2196_),
    .B(_2195_),
    .A_N(_2031_));
 sg13g2_a21oi_1 _7008_ (.A1(_1951_),
    .A2(_1946_),
    .Y(_2197_),
    .B1(_2196_));
 sg13g2_o21ai_1 _7009_ (.B1(_2197_),
    .Y(_2198_),
    .A1(_2193_),
    .A2(_2194_));
 sg13g2_and4_1 _7010_ (.A(_4085_),
    .B(_1437_),
    .C(_1751_),
    .D(_2175_),
    .X(_2199_));
 sg13g2_o21ai_1 _7011_ (.B1(_0351_),
    .Y(_2200_),
    .A1(_4103_),
    .A2(_1447_));
 sg13g2_a21o_1 _7012_ (.A2(_2035_),
    .A1(_3749_),
    .B1(_3725_),
    .X(_2201_));
 sg13g2_or2_1 _7013_ (.X(_2202_),
    .B(_3747_),
    .A(_3723_));
 sg13g2_a21o_1 _7014_ (.A2(_2202_),
    .A1(net126),
    .B1(net127),
    .X(_2203_));
 sg13g2_o21ai_1 _7015_ (.B1(_2203_),
    .Y(_2204_),
    .A1(_2128_),
    .A2(net126));
 sg13g2_a221oi_1 _7016_ (.B2(_2000_),
    .C1(_2204_),
    .B1(_2201_),
    .A1(_3725_),
    .Y(_2205_),
    .A2(_2035_));
 sg13g2_a221oi_1 _7017_ (.B2(_2200_),
    .C1(_2205_),
    .B1(_2199_),
    .A1(_0377_),
    .Y(_2206_),
    .A2(_2176_));
 sg13g2_nor2_1 _7018_ (.A(_3861_),
    .B(_2189_),
    .Y(_2207_));
 sg13g2_and3_1 _7019_ (.X(_2208_),
    .A(_2198_),
    .B(_2206_),
    .C(_2207_));
 sg13g2_and3_1 _7020_ (.X(_2209_),
    .A(_2184_),
    .B(_2188_),
    .C(_2208_));
 sg13g2_nor2_1 _7021_ (.A(_2206_),
    .B(_2190_),
    .Y(_2210_));
 sg13g2_nand2_1 _7022_ (.Y(_2211_),
    .A(net113),
    .B(_0011_));
 sg13g2_o21ai_1 _7023_ (.B1(_2211_),
    .Y(_2212_),
    .A1(_2198_),
    .A2(_2190_));
 sg13g2_nor4_2 _7024_ (.A(_2191_),
    .B(_2209_),
    .C(_2210_),
    .Y(_2213_),
    .D(_2212_));
 sg13g2_nand2_1 _7025_ (.Y(_2214_),
    .A(net106),
    .B(_2213_));
 sg13g2_a22oi_1 _7026_ (.Y(_2215_),
    .B1(_2078_),
    .B2(_1487_),
    .A2(_2045_),
    .A1(_3771_));
 sg13g2_a21oi_1 _7027_ (.A1(_2214_),
    .A2(_2215_),
    .Y(_0064_),
    .B1(net93));
 sg13g2_nand4_1 _7028_ (.B(_0542_),
    .C(_0551_),
    .A(_0536_),
    .Y(_2216_),
    .D(_0557_));
 sg13g2_nand4_1 _7029_ (.B(_0655_),
    .C(_0663_),
    .A(_0420_),
    .Y(_2217_),
    .D(_1519_));
 sg13g2_nand2_1 _7030_ (.Y(_2218_),
    .A(_0597_),
    .B(_1503_));
 sg13g2_inv_1 _7031_ (.Y(_2219_),
    .A(_3724_));
 sg13g2_inv_2 _7032_ (.Y(_2220_),
    .A(net297));
 sg13g2_nand4_1 _7033_ (.B(_2219_),
    .C(_2220_),
    .A(_3747_),
    .Y(_2221_),
    .D(_2101_));
 sg13g2_and2_1 _7034_ (.A(net309),
    .B(\collatz.iter[132] ),
    .X(_2222_));
 sg13g2_buf_1 _7035_ (.A(_2222_),
    .X(_2223_));
 sg13g2_nand3_1 _7036_ (.B(_3749_),
    .C(_2223_),
    .A(_3723_),
    .Y(_2224_));
 sg13g2_a22oi_1 _7037_ (.Y(_2225_),
    .B1(_2221_),
    .B2(_2224_),
    .A2(_2053_),
    .A1(_2051_));
 sg13g2_nand4_1 _7038_ (.B(_1874_),
    .C(_1964_),
    .A(_1770_),
    .Y(_2226_),
    .D(_2225_));
 sg13g2_nor4_2 _7039_ (.A(_2216_),
    .B(_2217_),
    .C(_2218_),
    .Y(_2227_),
    .D(_2226_));
 sg13g2_nor2b_1 _7040_ (.A(_0525_),
    .B_N(_2227_),
    .Y(_2228_));
 sg13g2_buf_1 _7041_ (.A(_3877_),
    .X(_2229_));
 sg13g2_xnor2_1 _7042_ (.Y(_2230_),
    .A(net124),
    .B(net297));
 sg13g2_nor2_1 _7043_ (.A(_3861_),
    .B(_2230_),
    .Y(_2231_));
 sg13g2_buf_1 _7044_ (.A(net283),
    .X(_2232_));
 sg13g2_nand3_1 _7045_ (.B(_0524_),
    .C(_2227_),
    .A(_0505_),
    .Y(_2233_));
 sg13g2_and3_1 _7046_ (.X(_2234_),
    .A(net123),
    .B(_2230_),
    .C(_2233_));
 sg13g2_nand4_1 _7047_ (.B(_1874_),
    .C(_1964_),
    .A(_1770_),
    .Y(_2235_),
    .D(_2225_));
 sg13g2_a21oi_1 _7048_ (.A1(_0420_),
    .A2(_1507_),
    .Y(_2236_),
    .B1(_0642_));
 sg13g2_nor3_1 _7049_ (.A(_1520_),
    .B(_2235_),
    .C(_2236_),
    .Y(_2237_));
 sg13g2_or4_1 _7050_ (.A(_1281_),
    .B(_1520_),
    .C(_2235_),
    .D(_2218_),
    .X(_2238_));
 sg13g2_nand2_1 _7051_ (.Y(_2239_),
    .A(_2219_),
    .B(_2220_));
 sg13g2_nor2_1 _7052_ (.A(_2066_),
    .B(_2239_),
    .Y(_2240_));
 sg13g2_nor2_1 _7053_ (.A(_3749_),
    .B(_2240_),
    .Y(_2241_));
 sg13g2_o21ai_1 _7054_ (.B1(_2239_),
    .Y(_2242_),
    .A1(net125),
    .A2(_2066_));
 sg13g2_nor2_1 _7055_ (.A(net125),
    .B(_2223_),
    .Y(_2243_));
 sg13g2_a21oi_1 _7056_ (.A1(_2099_),
    .A2(_2242_),
    .Y(_2244_),
    .B1(_2243_));
 sg13g2_o21ai_1 _7057_ (.B1(_2244_),
    .Y(_2245_),
    .A1(net128),
    .A2(_2241_));
 sg13g2_o21ai_1 _7058_ (.B1(_2245_),
    .Y(_2246_),
    .A1(_0592_),
    .A2(_2238_));
 sg13g2_a21oi_1 _7059_ (.A1(_1522_),
    .A2(_1524_),
    .Y(_2247_),
    .B1(_1530_));
 sg13g2_nand3b_1 _7060_ (.B(_1770_),
    .C(_1965_),
    .Y(_2248_),
    .A_N(_2247_));
 sg13g2_a221oi_1 _7061_ (.B2(_1974_),
    .C1(_2055_),
    .B1(_2248_),
    .A1(_2221_),
    .Y(_2249_),
    .A2(_2224_));
 sg13g2_and3_1 _7062_ (.X(_2250_),
    .A(_0665_),
    .B(_0666_),
    .C(_1519_));
 sg13g2_and3_1 _7063_ (.X(_2251_),
    .A(_0665_),
    .B(_0682_),
    .C(_1519_));
 sg13g2_a221oi_1 _7064_ (.B2(_0677_),
    .C1(_2251_),
    .B1(_2250_),
    .A1(_0688_),
    .Y(_2252_),
    .A2(_1519_));
 sg13g2_or2_1 _7065_ (.X(_2253_),
    .B(_2217_),
    .A(_1504_));
 sg13g2_a21oi_1 _7066_ (.A1(_2252_),
    .A2(_2253_),
    .Y(_2254_),
    .B1(_2226_));
 sg13g2_nor4_2 _7067_ (.A(_2237_),
    .B(_2246_),
    .C(_2249_),
    .Y(_2255_),
    .D(_2254_));
 sg13g2_mux2_1 _7068_ (.A0(_2231_),
    .A1(_2234_),
    .S(_2255_),
    .X(_2256_));
 sg13g2_a221oi_1 _7069_ (.B2(_2231_),
    .C1(_2256_),
    .B1(_2228_),
    .A1(net113),
    .Y(_2257_),
    .A2(_0010_));
 sg13g2_buf_2 _7070_ (.A(_2257_),
    .X(_2258_));
 sg13g2_nand2_1 _7071_ (.Y(_2259_),
    .A(net106),
    .B(_2258_));
 sg13g2_a22oi_1 _7072_ (.Y(_2260_),
    .B1(_2078_),
    .B2(_0699_),
    .A2(_2045_),
    .A1(_2229_));
 sg13g2_a21oi_1 _7073_ (.A1(_2259_),
    .A2(_2260_),
    .Y(_0065_),
    .B1(net93));
 sg13g2_buf_1 _7074_ (.A(_3772_),
    .X(_2261_));
 sg13g2_xor2_1 _7075_ (.B(net122),
    .A(net124),
    .X(_2262_));
 sg13g2_o21ai_1 _7076_ (.B1(_1794_),
    .Y(_2263_),
    .A1(_1612_),
    .A2(_1614_));
 sg13g2_nor4_1 _7077_ (.A(_1801_),
    .B(_1802_),
    .C(_1994_),
    .D(_1995_),
    .Y(_2264_));
 sg13g2_nand2_1 _7078_ (.Y(_2265_),
    .A(_3749_),
    .B(_2223_));
 sg13g2_nor2b_1 _7079_ (.A(_3771_),
    .B_N(_3877_),
    .Y(_2266_));
 sg13g2_nand3_1 _7080_ (.B(_2171_),
    .C(_2266_),
    .A(net127),
    .Y(_2267_));
 sg13g2_o21ai_1 _7081_ (.B1(_2267_),
    .Y(_2268_),
    .A1(net124),
    .A2(_2265_));
 sg13g2_buf_1 _7082_ (.A(_2268_),
    .X(_2269_));
 sg13g2_nand2_1 _7083_ (.Y(_2270_),
    .A(_2104_),
    .B(_2269_));
 sg13g2_a221oi_1 _7084_ (.B2(_2264_),
    .C1(_2270_),
    .B1(_2263_),
    .A1(_1996_),
    .Y(_2271_),
    .A2(_1989_));
 sg13g2_a21oi_1 _7085_ (.A1(net127),
    .A2(net126),
    .Y(_2272_),
    .B1(net124));
 sg13g2_and2_1 _7086_ (.A(net309),
    .B(net124),
    .X(_2273_));
 sg13g2_o21ai_1 _7087_ (.B1(net125),
    .Y(_2274_),
    .A1(net297),
    .A2(_2273_));
 sg13g2_o21ai_1 _7088_ (.B1(_2274_),
    .Y(_2275_),
    .A1(_2220_),
    .A2(_2272_));
 sg13g2_a21oi_1 _7089_ (.A1(_2113_),
    .A2(_2269_),
    .Y(_2276_),
    .B1(_2275_));
 sg13g2_nand2b_1 _7090_ (.Y(_2277_),
    .B(_2276_),
    .A_N(_2271_));
 sg13g2_nor2_1 _7091_ (.A(_0736_),
    .B(_1600_),
    .Y(_2278_));
 sg13g2_o21ai_1 _7092_ (.B1(_0903_),
    .Y(_2279_),
    .A1(_0725_),
    .A2(_1601_));
 sg13g2_and2_1 _7093_ (.A(_2278_),
    .B(_2279_),
    .X(_2280_));
 sg13g2_and2_1 _7094_ (.A(_0922_),
    .B(_1579_),
    .X(_2281_));
 sg13g2_and3_1 _7095_ (.X(_2282_),
    .A(_0922_),
    .B(_1572_),
    .C(_1579_));
 sg13g2_or2_1 _7096_ (.X(_2283_),
    .B(_0847_),
    .A(_0842_));
 sg13g2_a22oi_1 _7097_ (.Y(_2284_),
    .B1(_2282_),
    .B2(_2283_),
    .A2(_2281_),
    .A1(_1577_));
 sg13g2_a21oi_1 _7098_ (.A1(_0922_),
    .A2(_1585_),
    .Y(_2285_),
    .B1(_1598_));
 sg13g2_and3_1 _7099_ (.X(_2286_),
    .A(_2278_),
    .B(_2279_),
    .C(_2285_));
 sg13g2_a22oi_1 _7100_ (.Y(_2287_),
    .B1(_1985_),
    .B2(_1987_),
    .A2(_1899_),
    .A1(_1898_));
 sg13g2_nand4_1 _7101_ (.B(_2287_),
    .C(_2104_),
    .A(_1794_),
    .Y(_2288_),
    .D(_2269_));
 sg13g2_buf_1 _7102_ (.A(_2288_),
    .X(_2289_));
 sg13g2_nand3b_1 _7103_ (.B(_1706_),
    .C(_1333_),
    .Y(_2290_),
    .A_N(_2289_));
 sg13g2_a221oi_1 _7104_ (.B2(_2286_),
    .C1(_2290_),
    .B1(_2284_),
    .A1(_2280_),
    .Y(_2291_),
    .A2(_1588_));
 sg13g2_or4_1 _7105_ (.A(_3861_),
    .B(_2262_),
    .C(_2277_),
    .D(_2291_),
    .X(_2292_));
 sg13g2_nand2_1 _7106_ (.Y(_2293_),
    .A(net283),
    .B(_2262_));
 sg13g2_nand2_1 _7107_ (.Y(_2294_),
    .A(_1593_),
    .B(_2282_));
 sg13g2_nor4_2 _7108_ (.A(_0879_),
    .B(_1569_),
    .C(_2294_),
    .Y(_2295_),
    .D(_2289_));
 sg13g2_mux2_1 _7109_ (.A0(_2292_),
    .A1(_2293_),
    .S(_2295_),
    .X(_2296_));
 sg13g2_inv_1 _7110_ (.Y(_2297_),
    .A(_2293_));
 sg13g2_nand2_1 _7111_ (.Y(_2298_),
    .A(_2297_),
    .B(_2291_));
 sg13g2_a22oi_1 _7112_ (.Y(_2299_),
    .B1(_2277_),
    .B2(_2297_),
    .A2(_0009_),
    .A1(net113));
 sg13g2_and3_1 _7113_ (.X(_2300_),
    .A(_2296_),
    .B(_2298_),
    .C(_2299_));
 sg13g2_buf_1 _7114_ (.A(_2300_),
    .X(_2301_));
 sg13g2_nand2_1 _7115_ (.Y(_2302_),
    .A(net106),
    .B(_2301_));
 sg13g2_a22oi_1 _7116_ (.Y(_2303_),
    .B1(_2078_),
    .B2(_1623_),
    .A2(_2045_),
    .A1(net122));
 sg13g2_a21oi_1 _7117_ (.A1(_2302_),
    .A2(_2303_),
    .Y(_0066_),
    .B1(net93));
 sg13g2_nand2_1 _7118_ (.Y(_2304_),
    .A(net297),
    .B(_3772_));
 sg13g2_nor4_1 _7119_ (.A(_3747_),
    .B(_2219_),
    .C(net124),
    .D(_2304_),
    .Y(_2305_));
 sg13g2_inv_1 _7120_ (.Y(_2306_),
    .A(_3747_));
 sg13g2_inv_1 _7121_ (.Y(_2307_),
    .A(_3877_));
 sg13g2_nor4_1 _7122_ (.A(_2306_),
    .B(net309),
    .C(_2307_),
    .D(_3774_),
    .Y(_2308_));
 sg13g2_o21ai_1 _7123_ (.B1(_2133_),
    .Y(_2309_),
    .A1(_2305_),
    .A2(_2308_));
 sg13g2_buf_1 _7124_ (.A(_2309_),
    .X(_2310_));
 sg13g2_or4_1 _7125_ (.A(_1637_),
    .B(_1814_),
    .C(_2016_),
    .D(_2310_),
    .X(_2311_));
 sg13g2_buf_1 _7126_ (.A(_2311_),
    .X(_2312_));
 sg13g2_nor3_1 _7127_ (.A(_1187_),
    .B(_0996_),
    .C(_2312_),
    .Y(_2313_));
 sg13g2_nor4_1 _7128_ (.A(_1187_),
    .B(_1179_),
    .C(_0996_),
    .D(_2312_),
    .Y(_2314_));
 sg13g2_nor3_1 _7129_ (.A(_1187_),
    .B(_0990_),
    .C(_2312_),
    .Y(_2315_));
 sg13g2_or2_1 _7130_ (.X(_2316_),
    .B(_2315_),
    .A(_2314_));
 sg13g2_a21oi_1 _7131_ (.A1(_1171_),
    .A2(_2313_),
    .Y(_2317_),
    .B1(_2316_));
 sg13g2_buf_1 _7132_ (.A(_3878_),
    .X(_2318_));
 sg13g2_xnor2_1 _7133_ (.Y(_2319_),
    .A(_2318_),
    .B(_2261_));
 sg13g2_nand2b_1 _7134_ (.Y(_2320_),
    .B(net103),
    .A_N(_2319_));
 sg13g2_nor2_1 _7135_ (.A(_2317_),
    .B(_2320_),
    .Y(_2321_));
 sg13g2_inv_1 _7136_ (.Y(_2322_),
    .A(_2144_));
 sg13g2_nor2_1 _7137_ (.A(_2305_),
    .B(_2308_),
    .Y(_2323_));
 sg13g2_nand2b_1 _7138_ (.Y(_2324_),
    .B(_2304_),
    .A_N(_2273_));
 sg13g2_a22oi_1 _7139_ (.Y(_2325_),
    .B1(_2324_),
    .B2(net125),
    .A2(_3774_),
    .A1(net124));
 sg13g2_o21ai_1 _7140_ (.B1(_2325_),
    .Y(_2326_),
    .A1(_2322_),
    .A2(_2323_));
 sg13g2_nand2b_1 _7141_ (.Y(_2327_),
    .B(_1646_),
    .A_N(_1814_));
 sg13g2_a21oi_1 _7142_ (.A1(_1818_),
    .A2(_2327_),
    .Y(_2328_),
    .B1(_2016_));
 sg13g2_nor2_1 _7143_ (.A(_2015_),
    .B(_2328_),
    .Y(_2329_));
 sg13g2_nor2_1 _7144_ (.A(_2310_),
    .B(_2329_),
    .Y(_2330_));
 sg13g2_nor2_1 _7145_ (.A(_2326_),
    .B(_2330_),
    .Y(_2331_));
 sg13g2_and4_1 _7146_ (.A(net81),
    .B(_2319_),
    .C(_2331_),
    .D(_2317_),
    .X(_2332_));
 sg13g2_nand2_1 _7147_ (.Y(_2333_),
    .A(net113),
    .B(_0008_));
 sg13g2_o21ai_1 _7148_ (.B1(_2333_),
    .Y(_2334_),
    .A1(_2331_),
    .A2(_2320_));
 sg13g2_nor3_1 _7149_ (.A(_2321_),
    .B(_2332_),
    .C(_2334_),
    .Y(_2335_));
 sg13g2_nand2_1 _7150_ (.Y(_2336_),
    .A(net100),
    .B(_2335_));
 sg13g2_a22oi_1 _7151_ (.Y(_2337_),
    .B1(_2078_),
    .B2(_1655_),
    .A2(_2045_),
    .A1(net121));
 sg13g2_a21oi_1 _7152_ (.A1(_2336_),
    .A2(_2337_),
    .Y(_0067_),
    .B1(net93));
 sg13g2_xor2_1 _7153_ (.B(net205),
    .A(net121),
    .X(_2338_));
 sg13g2_inv_2 _7154_ (.Y(_2339_),
    .A(_3878_));
 sg13g2_o21ai_1 _7155_ (.B1(_2339_),
    .Y(_2340_),
    .A1(_2306_),
    .A2(_2220_));
 sg13g2_inv_1 _7156_ (.Y(_2341_),
    .A(_3772_));
 sg13g2_o21ai_1 _7157_ (.B1(_2341_),
    .Y(_2342_),
    .A1(_2220_),
    .A2(_2339_));
 sg13g2_a22oi_1 _7158_ (.Y(_2343_),
    .B1(_2342_),
    .B2(_2229_),
    .A2(_2340_),
    .A1(_2261_));
 sg13g2_a21oi_1 _7159_ (.A1(_2000_),
    .A2(_3749_),
    .Y(_2344_),
    .B1(_3725_));
 sg13g2_a21oi_1 _7160_ (.A1(_2000_),
    .A2(_2052_),
    .Y(_2345_),
    .B1(_2306_));
 sg13g2_o21ai_1 _7161_ (.B1(_2203_),
    .Y(_2346_),
    .A1(_2090_),
    .A2(_2345_));
 sg13g2_nand3_1 _7162_ (.B(net122),
    .C(_3879_),
    .A(net297),
    .Y(_2347_));
 sg13g2_nor2b_1 _7163_ (.A(_3772_),
    .B_N(net121),
    .Y(_2348_));
 sg13g2_nand3_1 _7164_ (.B(_2266_),
    .C(_2348_),
    .A(net125),
    .Y(_2349_));
 sg13g2_o21ai_1 _7165_ (.B1(_2349_),
    .Y(_2350_),
    .A1(net125),
    .A2(_2347_));
 sg13g2_nor2b_1 _7166_ (.A(_2346_),
    .B_N(_2350_),
    .Y(_2351_));
 sg13g2_o21ai_1 _7167_ (.B1(_2351_),
    .Y(_2352_),
    .A1(_2036_),
    .A2(_2344_));
 sg13g2_nand2_1 _7168_ (.Y(_2353_),
    .A(_2343_),
    .B(_2352_));
 sg13g2_nor3_1 _7169_ (.A(net113),
    .B(_2338_),
    .C(_2353_),
    .Y(_2354_));
 sg13g2_and3_1 _7170_ (.X(_2355_),
    .A(_2032_),
    .B(_2195_),
    .C(_2350_));
 sg13g2_and3_1 _7171_ (.X(_2356_),
    .A(net202),
    .B(_2338_),
    .C(_2355_));
 sg13g2_mux2_1 _7172_ (.A0(_2354_),
    .A1(_2356_),
    .S(_1858_),
    .X(_2357_));
 sg13g2_nor2_1 _7173_ (.A(_2338_),
    .B(_2355_),
    .Y(_2358_));
 sg13g2_mux2_1 _7174_ (.A0(_2358_),
    .A1(_2338_),
    .S(_2353_),
    .X(_2359_));
 sg13g2_mux2_1 _7175_ (.A0(_0007_),
    .A1(_2359_),
    .S(_4029_),
    .X(_2360_));
 sg13g2_nor2_1 _7176_ (.A(_2357_),
    .B(_2360_),
    .Y(_2361_));
 sg13g2_nand2_1 _7177_ (.Y(_2362_),
    .A(net100),
    .B(_2361_));
 sg13g2_buf_1 _7178_ (.A(net77),
    .X(_2363_));
 sg13g2_inv_2 _7179_ (.Y(_2364_),
    .A(net205));
 sg13g2_and2_1 _7180_ (.A(_3976_),
    .B(_1549_),
    .X(_2365_));
 sg13g2_buf_2 _7181_ (.A(_2365_),
    .X(_2366_));
 sg13g2_buf_1 _7182_ (.A(_2366_),
    .X(_2367_));
 sg13g2_nand2_1 _7183_ (.Y(_2368_),
    .A(_4028_),
    .B(_2367_));
 sg13g2_o21ai_1 _7184_ (.B1(_2368_),
    .Y(_2369_),
    .A1(_2364_),
    .A2(net58));
 sg13g2_nand2_1 _7185_ (.Y(_2370_),
    .A(net59),
    .B(_2369_));
 sg13g2_buf_1 _7186_ (.A(net204),
    .X(_2371_));
 sg13g2_a21oi_1 _7187_ (.A1(_2362_),
    .A2(_2370_),
    .Y(_0068_),
    .B1(net91));
 sg13g2_nand2_1 _7188_ (.Y(_2372_),
    .A(_0666_),
    .B(_0667_));
 sg13g2_nand2_1 _7189_ (.Y(_2373_),
    .A(_2221_),
    .B(_2224_));
 sg13g2_nand3_1 _7190_ (.B(_2266_),
    .C(_2348_),
    .A(_2364_),
    .Y(_2374_));
 sg13g2_o21ai_1 _7191_ (.B1(_2374_),
    .Y(_2375_),
    .A1(_2364_),
    .A2(_2347_));
 sg13g2_nand3_1 _7192_ (.B(_2373_),
    .C(_2375_),
    .A(_2062_),
    .Y(_2376_));
 sg13g2_nor3_1 _7193_ (.A(_2372_),
    .B(_2056_),
    .C(_2376_),
    .Y(_2377_));
 sg13g2_buf_1 _7194_ (.A(_3855_),
    .X(_2378_));
 sg13g2_xnor2_1 _7195_ (.Y(_2379_),
    .A(net120),
    .B(net205));
 sg13g2_nor2_1 _7196_ (.A(_3861_),
    .B(_2379_),
    .Y(_2380_));
 sg13g2_nand3_1 _7197_ (.B(_2377_),
    .C(_2380_),
    .A(_1308_),
    .Y(_2381_));
 sg13g2_a22oi_1 _7198_ (.Y(_2382_),
    .B1(_0674_),
    .B2(_0675_),
    .A2(_0648_),
    .A1(_0645_));
 sg13g2_o21ai_1 _7199_ (.B1(_1314_),
    .Y(_2383_),
    .A1(_0682_),
    .A2(_2382_));
 sg13g2_a21o_1 _7200_ (.A2(_2383_),
    .A1(_1253_),
    .B1(_1875_),
    .X(_2384_));
 sg13g2_a21o_1 _7201_ (.A2(_2384_),
    .A1(_1883_),
    .B1(_2376_),
    .X(_2385_));
 sg13g2_inv_1 _7202_ (.Y(_2386_),
    .A(_2375_));
 sg13g2_a21oi_1 _7203_ (.A1(_2202_),
    .A2(_2239_),
    .Y(_2387_),
    .B1(net127));
 sg13g2_nor3_1 _7204_ (.A(_2243_),
    .B(_2386_),
    .C(_2387_),
    .Y(_2388_));
 sg13g2_a21oi_1 _7205_ (.A1(_2220_),
    .A2(_3725_),
    .Y(_2389_),
    .B1(_3749_));
 sg13g2_or2_1 _7206_ (.X(_2390_),
    .B(_2389_),
    .A(_2068_));
 sg13g2_a22oi_1 _7207_ (.Y(_2391_),
    .B1(net122),
    .B2(_3949_),
    .A2(net121),
    .A1(net297));
 sg13g2_o21ai_1 _7208_ (.B1(net121),
    .Y(_2392_),
    .A1(net122),
    .A2(net205));
 sg13g2_o21ai_1 _7209_ (.B1(_2392_),
    .Y(_2393_),
    .A1(_2307_),
    .A2(_2391_));
 sg13g2_a21oi_1 _7210_ (.A1(_2388_),
    .A2(_2390_),
    .Y(_2394_),
    .B1(_2393_));
 sg13g2_nand4_1 _7211_ (.B(_2379_),
    .C(_2385_),
    .A(net123),
    .Y(_2395_),
    .D(_2394_));
 sg13g2_a21o_1 _7212_ (.A2(_2377_),
    .A1(_1308_),
    .B1(_2395_),
    .X(_2396_));
 sg13g2_nand2_1 _7213_ (.Y(_2397_),
    .A(_2385_),
    .B(_2394_));
 sg13g2_a22oi_1 _7214_ (.Y(_2398_),
    .B1(_2397_),
    .B2(_2380_),
    .A2(_0006_),
    .A1(net113));
 sg13g2_nand3_1 _7215_ (.B(_2396_),
    .C(_2398_),
    .A(_2381_),
    .Y(_2399_));
 sg13g2_buf_1 _7216_ (.A(_2399_),
    .X(_2400_));
 sg13g2_or2_1 _7217_ (.X(_2401_),
    .B(_2400_),
    .A(_3958_));
 sg13g2_inv_1 _7218_ (.Y(_2402_),
    .A(_3855_));
 sg13g2_nand2_1 _7219_ (.Y(_2403_),
    .A(net274),
    .B(_2366_));
 sg13g2_o21ai_1 _7220_ (.B1(_2403_),
    .Y(_2404_),
    .A1(_2402_),
    .A2(net58));
 sg13g2_nand2_1 _7221_ (.Y(_2405_),
    .A(net59),
    .B(_2404_));
 sg13g2_a21oi_1 _7222_ (.A1(_2401_),
    .A2(_2405_),
    .Y(_0069_),
    .B1(net91));
 sg13g2_nand2_1 _7223_ (.Y(_2406_),
    .A(_3862_),
    .B(_0005_));
 sg13g2_xor2_1 _7224_ (.B(net228),
    .A(net120),
    .X(_2407_));
 sg13g2_or2_1 _7225_ (.X(_2408_),
    .B(_2407_),
    .A(_3861_));
 sg13g2_nand2_1 _7226_ (.Y(_2409_),
    .A(net202),
    .B(_2407_));
 sg13g2_inv_1 _7227_ (.Y(_2410_),
    .A(_2105_));
 sg13g2_o21ai_1 _7228_ (.B1(_1908_),
    .Y(_2411_),
    .A1(_1718_),
    .A2(_1901_));
 sg13g2_a221oi_1 _7229_ (.B2(_2411_),
    .C1(_2113_),
    .B1(_2410_),
    .A1(_1994_),
    .Y(_2412_),
    .A2(_2104_));
 sg13g2_nand3_1 _7230_ (.B(_3949_),
    .C(_3879_),
    .A(net122),
    .Y(_2413_));
 sg13g2_nor2b_1 _7231_ (.A(_3949_),
    .B_N(_3855_),
    .Y(_2414_));
 sg13g2_nand3_1 _7232_ (.B(_2348_),
    .C(_2414_),
    .A(net124),
    .Y(_2415_));
 sg13g2_o21ai_1 _7233_ (.B1(_2415_),
    .Y(_2416_),
    .A1(_3855_),
    .A2(_2413_));
 sg13g2_nand2_1 _7234_ (.Y(_2417_),
    .A(_2269_),
    .B(_2416_));
 sg13g2_o21ai_1 _7235_ (.B1(_2402_),
    .Y(_2418_),
    .A1(_2307_),
    .A2(_2341_));
 sg13g2_o21ai_1 _7236_ (.B1(_2364_),
    .Y(_2419_),
    .A1(_2341_),
    .A2(_2402_));
 sg13g2_a22oi_1 _7237_ (.Y(_2420_),
    .B1(_2419_),
    .B2(net121),
    .A2(_2418_),
    .A1(net205));
 sg13g2_inv_1 _7238_ (.Y(_2421_),
    .A(_2420_));
 sg13g2_a21oi_1 _7239_ (.A1(_2275_),
    .A2(_2416_),
    .Y(_2422_),
    .B1(_2421_));
 sg13g2_o21ai_1 _7240_ (.B1(_2422_),
    .Y(_2423_),
    .A1(_2412_),
    .A2(_2417_));
 sg13g2_nor3_1 _7241_ (.A(_0737_),
    .B(_1338_),
    .C(_2423_),
    .Y(_2424_));
 sg13g2_nor4_1 _7242_ (.A(_1712_),
    .B(_1901_),
    .C(_2105_),
    .D(_2417_),
    .Y(_2425_));
 sg13g2_nand3_1 _7243_ (.B(_1330_),
    .C(_1332_),
    .A(_1613_),
    .Y(_2426_));
 sg13g2_a21oi_1 _7244_ (.A1(_2425_),
    .A2(_2426_),
    .Y(_2427_),
    .B1(_2423_));
 sg13g2_a21oi_1 _7245_ (.A1(_0961_),
    .A2(_2424_),
    .Y(_2428_),
    .B1(_2427_));
 sg13g2_mux2_1 _7246_ (.A0(_2408_),
    .A1(_2409_),
    .S(_2428_),
    .X(_2429_));
 sg13g2_buf_1 _7247_ (.A(_2429_),
    .X(_2430_));
 sg13g2_nand3_1 _7248_ (.B(_2406_),
    .C(_2430_),
    .A(net100),
    .Y(_2431_));
 sg13g2_inv_1 _7249_ (.Y(_2432_),
    .A(net228));
 sg13g2_nand2_1 _7250_ (.Y(_2433_),
    .A(net262),
    .B(_2366_));
 sg13g2_o21ai_1 _7251_ (.B1(_2433_),
    .Y(_2434_),
    .A1(_2432_),
    .A2(net58));
 sg13g2_nand2_1 _7252_ (.Y(_2435_),
    .A(net59),
    .B(_2434_));
 sg13g2_a21oi_1 _7253_ (.A1(_2431_),
    .A2(_2435_),
    .Y(_0070_),
    .B1(net91));
 sg13g2_nor4_1 _7254_ (.A(_2339_),
    .B(net122),
    .C(_3949_),
    .D(net228),
    .Y(_2436_));
 sg13g2_nand2_1 _7255_ (.Y(_2437_),
    .A(_3949_),
    .B(_3868_));
 sg13g2_nor4_1 _7256_ (.A(net121),
    .B(_2341_),
    .C(_3855_),
    .D(_2437_),
    .Y(_2438_));
 sg13g2_a21oi_1 _7257_ (.A1(net120),
    .A2(_2436_),
    .Y(_2439_),
    .B1(_2438_));
 sg13g2_or3_1 _7258_ (.A(_2134_),
    .B(_2323_),
    .C(_2439_),
    .X(_2440_));
 sg13g2_nor2_1 _7259_ (.A(_1926_),
    .B(_2440_),
    .Y(_2441_));
 sg13g2_nand3_1 _7260_ (.B(_1387_),
    .C(_2441_),
    .A(_1373_),
    .Y(_2442_));
 sg13g2_inv_1 _7261_ (.Y(_2443_),
    .A(_2439_));
 sg13g2_a21oi_1 _7262_ (.A1(_2014_),
    .A2(_2133_),
    .Y(_2444_),
    .B1(_2144_));
 sg13g2_o21ai_1 _7263_ (.B1(_2325_),
    .Y(_2445_),
    .A1(_2323_),
    .A2(_2444_));
 sg13g2_a22oi_1 _7264_ (.Y(_2446_),
    .B1(net205),
    .B2(net228),
    .A2(net120),
    .A1(net122));
 sg13g2_o21ai_1 _7265_ (.B1(_2378_),
    .Y(_2447_),
    .A1(net205),
    .A2(net228));
 sg13g2_o21ai_1 _7266_ (.B1(_2447_),
    .Y(_2448_),
    .A1(_2339_),
    .A2(_2446_));
 sg13g2_a21oi_1 _7267_ (.A1(_2443_),
    .A2(_2445_),
    .Y(_2449_),
    .B1(_2448_));
 sg13g2_o21ai_1 _7268_ (.B1(_2449_),
    .Y(_2450_),
    .A1(_1934_),
    .A2(_2440_));
 sg13g2_a21oi_1 _7269_ (.A1(_1412_),
    .A2(_2441_),
    .Y(_2451_),
    .B1(_2450_));
 sg13g2_nand4_1 _7270_ (.B(_1370_),
    .C(_1387_),
    .A(_1354_),
    .Y(_2452_),
    .D(_2441_));
 sg13g2_nand3_1 _7271_ (.B(_2451_),
    .C(_2452_),
    .A(_2442_),
    .Y(_2453_));
 sg13g2_buf_1 _7272_ (.A(_2453_),
    .X(_2454_));
 sg13g2_buf_1 _7273_ (.A(_3856_),
    .X(_2455_));
 sg13g2_xor2_1 _7274_ (.B(net228),
    .A(_2455_),
    .X(_2456_));
 sg13g2_xnor2_1 _7275_ (.Y(_2457_),
    .A(_2454_),
    .B(_2456_));
 sg13g2_nor2b_1 _7276_ (.A(net103),
    .B_N(_0004_),
    .Y(_2458_));
 sg13g2_a21oi_1 _7277_ (.A1(net67),
    .A2(_2457_),
    .Y(_2459_),
    .B1(_2458_));
 sg13g2_nand2_1 _7278_ (.Y(_2460_),
    .A(net100),
    .B(_2459_));
 sg13g2_inv_1 _7279_ (.Y(_2461_),
    .A(net119));
 sg13g2_nand2_1 _7280_ (.Y(_2462_),
    .A(_1745_),
    .B(_2366_));
 sg13g2_o21ai_1 _7281_ (.B1(_2462_),
    .Y(_2463_),
    .A1(_2461_),
    .A2(net58));
 sg13g2_nand2_1 _7282_ (.Y(_2464_),
    .A(net59),
    .B(_2463_));
 sg13g2_a21oi_1 _7283_ (.A1(_2460_),
    .A2(_2464_),
    .Y(_0071_),
    .B1(net91));
 sg13g2_buf_1 _7284_ (.A(net204),
    .X(_2465_));
 sg13g2_buf_1 _7285_ (.A(net78),
    .X(_2466_));
 sg13g2_or2_1 _7286_ (.X(_2467_),
    .B(_0740_),
    .A(_0273_));
 sg13g2_nand3_1 _7287_ (.B(_0458_),
    .C(_1494_),
    .A(_0456_),
    .Y(_2468_));
 sg13g2_xnor2_1 _7288_ (.Y(_2469_),
    .A(_2467_),
    .B(_2468_));
 sg13g2_buf_1 _7289_ (.A(_0692_),
    .X(_2470_));
 sg13g2_nor2_1 _7290_ (.A(_2470_),
    .B(net222),
    .Y(_2471_));
 sg13g2_a21oi_1 _7291_ (.A1(net39),
    .A2(_2469_),
    .Y(_2472_),
    .B1(_2471_));
 sg13g2_nand2_1 _7292_ (.Y(_2473_),
    .A(net326),
    .B(net63));
 sg13g2_nand2b_1 _7293_ (.Y(_2474_),
    .B(net250),
    .A_N(_1551_));
 sg13g2_a21oi_1 _7294_ (.A1(_2473_),
    .A2(_2474_),
    .Y(_2475_),
    .B1(_4039_));
 sg13g2_a21oi_1 _7295_ (.A1(_2466_),
    .A2(_2472_),
    .Y(_2476_),
    .B1(_2475_));
 sg13g2_nor2_1 _7296_ (.A(net90),
    .B(_2476_),
    .Y(_0072_));
 sg13g2_or2_1 _7297_ (.X(_2477_),
    .B(_0003_),
    .A(net123));
 sg13g2_xnor2_1 _7298_ (.Y(_2478_),
    .A(net119),
    .B(_3830_));
 sg13g2_nor4_1 _7299_ (.A(net121),
    .B(_2378_),
    .C(net119),
    .D(_2437_),
    .Y(_2479_));
 sg13g2_nand2_1 _7300_ (.Y(_2480_),
    .A(_3855_),
    .B(_3856_));
 sg13g2_nor4_1 _7301_ (.A(_2339_),
    .B(net205),
    .C(net228),
    .D(_2480_),
    .Y(_2481_));
 sg13g2_o21ai_1 _7302_ (.B1(_2350_),
    .Y(_2482_),
    .A1(_2479_),
    .A2(_2481_));
 sg13g2_or4_1 _7303_ (.A(_2192_),
    .B(_1946_),
    .C(_2196_),
    .D(_2482_),
    .X(_2483_));
 sg13g2_buf_1 _7304_ (.A(_2483_),
    .X(_2484_));
 sg13g2_nand2_1 _7305_ (.Y(_2485_),
    .A(_2478_),
    .B(_2484_));
 sg13g2_a21o_1 _7306_ (.A2(_1945_),
    .A1(_1850_),
    .B1(_1950_),
    .X(_2486_));
 sg13g2_a221oi_1 _7307_ (.B2(_1758_),
    .C1(_2205_),
    .B1(_2175_),
    .A1(_2486_),
    .Y(_2487_),
    .A2(_2173_));
 sg13g2_o21ai_1 _7308_ (.B1(_2461_),
    .Y(_2488_),
    .A1(_2364_),
    .A2(_2343_));
 sg13g2_o21ai_1 _7309_ (.B1(_2437_),
    .Y(_2489_),
    .A1(_2343_),
    .A2(_2480_));
 sg13g2_a21oi_1 _7310_ (.A1(_3950_),
    .A2(_2455_),
    .Y(_2490_),
    .B1(_3869_));
 sg13g2_nor2_1 _7311_ (.A(_2402_),
    .B(_2490_),
    .Y(_2491_));
 sg13g2_a221oi_1 _7312_ (.B2(_2318_),
    .C1(_2491_),
    .B1(_2489_),
    .A1(_3869_),
    .Y(_2492_),
    .A2(_2488_));
 sg13g2_o21ai_1 _7313_ (.B1(_2492_),
    .Y(_2493_),
    .A1(_2482_),
    .A2(_2487_));
 sg13g2_mux2_1 _7314_ (.A0(_2485_),
    .A1(_2478_),
    .S(_2493_),
    .X(_2494_));
 sg13g2_nand2_1 _7315_ (.Y(_2495_),
    .A(net202),
    .B(_2494_));
 sg13g2_nor3_1 _7316_ (.A(_3861_),
    .B(_2478_),
    .C(_2484_),
    .Y(_2496_));
 sg13g2_nand2_1 _7317_ (.Y(_2497_),
    .A(net123),
    .B(_2478_));
 sg13g2_nor3_1 _7318_ (.A(_1481_),
    .B(_2493_),
    .C(_2497_),
    .Y(_2498_));
 sg13g2_a221oi_1 _7319_ (.B2(_1481_),
    .C1(_2498_),
    .B1(_2496_),
    .A1(_2477_),
    .Y(_2499_),
    .A2(_2495_));
 sg13g2_nand2_1 _7320_ (.Y(_2500_),
    .A(_0399_),
    .B(_2499_));
 sg13g2_nand2_1 _7321_ (.Y(_2501_),
    .A(net327),
    .B(_2366_));
 sg13g2_o21ai_1 _7322_ (.B1(_2501_),
    .Y(_2502_),
    .A1(_3831_),
    .A2(_2367_));
 sg13g2_nand2_1 _7323_ (.Y(_2503_),
    .A(net59),
    .B(_2502_));
 sg13g2_a21oi_1 _7324_ (.A1(_2500_),
    .A2(_2503_),
    .Y(_0073_),
    .B1(net91));
 sg13g2_or2_1 _7325_ (.X(_2504_),
    .B(_0001_),
    .A(net123));
 sg13g2_nor2_1 _7326_ (.A(_3868_),
    .B(_3830_),
    .Y(_2505_));
 sg13g2_and2_1 _7327_ (.A(_3868_),
    .B(_3830_),
    .X(_2506_));
 sg13g2_buf_1 _7328_ (.A(_2506_),
    .X(_2507_));
 sg13g2_a21o_1 _7329_ (.A2(_2393_),
    .A1(net119),
    .B1(_2507_),
    .X(_2508_));
 sg13g2_nand2_1 _7330_ (.Y(_2509_),
    .A(_2393_),
    .B(_2507_));
 sg13g2_a21oi_1 _7331_ (.A1(_2480_),
    .A2(_2509_),
    .Y(_2510_),
    .B1(_2364_));
 sg13g2_a21oi_1 _7332_ (.A1(net120),
    .A2(_2508_),
    .Y(_2511_),
    .B1(_2510_));
 sg13g2_o21ai_1 _7333_ (.B1(_2511_),
    .Y(_2512_),
    .A1(_2461_),
    .A2(_2505_));
 sg13g2_buf_1 _7334_ (.A(_2512_),
    .X(_2513_));
 sg13g2_xor2_1 _7335_ (.B(_3830_),
    .A(net281),
    .X(_2514_));
 sg13g2_buf_1 _7336_ (.A(_2514_),
    .X(_2515_));
 sg13g2_nand2_1 _7337_ (.Y(_2516_),
    .A(_3857_),
    .B(_2507_));
 sg13g2_nand3_1 _7338_ (.B(_2505_),
    .C(_2414_),
    .A(net119),
    .Y(_2517_));
 sg13g2_o21ai_1 _7339_ (.B1(_2517_),
    .Y(_2518_),
    .A1(_2364_),
    .A2(_2516_));
 sg13g2_nand2_1 _7340_ (.Y(_2519_),
    .A(_2375_),
    .B(_2518_));
 sg13g2_inv_1 _7341_ (.Y(_2520_),
    .A(_2519_));
 sg13g2_nor3_1 _7342_ (.A(_2513_),
    .B(_2515_),
    .C(_2520_),
    .Y(_2521_));
 sg13g2_nand2_1 _7343_ (.Y(_2522_),
    .A(_2513_),
    .B(_2515_));
 sg13g2_nand3b_1 _7344_ (.B(net123),
    .C(_2522_),
    .Y(_2523_),
    .A_N(_2521_));
 sg13g2_nor4_1 _7345_ (.A(_3861_),
    .B(_2228_),
    .C(_2513_),
    .D(_2515_),
    .Y(_2524_));
 sg13g2_nand3_1 _7346_ (.B(_2515_),
    .C(_2520_),
    .A(net123),
    .Y(_2525_));
 sg13g2_a21oi_1 _7347_ (.A1(_2255_),
    .A2(_2233_),
    .Y(_2526_),
    .B1(_2525_));
 sg13g2_a221oi_1 _7348_ (.B2(_2255_),
    .C1(_2526_),
    .B1(_2524_),
    .A1(_2504_),
    .Y(_2527_),
    .A2(_2523_));
 sg13g2_nand2_1 _7349_ (.Y(_2528_),
    .A(net100),
    .B(_2527_));
 sg13g2_inv_1 _7350_ (.Y(_2529_),
    .A(_3870_));
 sg13g2_nand2_1 _7351_ (.Y(_2530_),
    .A(net326),
    .B(_2366_));
 sg13g2_o21ai_1 _7352_ (.B1(_2530_),
    .Y(_2531_),
    .A1(_2529_),
    .A2(net58));
 sg13g2_nand2_1 _7353_ (.Y(_2532_),
    .A(net60),
    .B(_2531_));
 sg13g2_a21oi_1 _7354_ (.A1(_2528_),
    .A2(_2532_),
    .Y(_0074_),
    .B1(net91));
 sg13g2_nor2_1 _7355_ (.A(_3833_),
    .B(net58),
    .Y(_2533_));
 sg13g2_a21oi_1 _7356_ (.A1(_1623_),
    .A2(net58),
    .Y(_2534_),
    .B1(_2533_));
 sg13g2_inv_1 _7357_ (.Y(_2535_),
    .A(_0000_));
 sg13g2_xnor2_1 _7358_ (.Y(_2536_),
    .A(net281),
    .B(_3832_));
 sg13g2_inv_1 _7359_ (.Y(_2537_),
    .A(_2275_));
 sg13g2_o21ai_1 _7360_ (.B1(_2269_),
    .Y(_2538_),
    .A1(_2113_),
    .A2(_2104_));
 sg13g2_nand4_1 _7361_ (.B(_3856_),
    .C(net281),
    .A(net120),
    .Y(_2539_),
    .D(_2505_));
 sg13g2_o21ai_1 _7362_ (.B1(_2539_),
    .Y(_2540_),
    .A1(net281),
    .A2(_2516_));
 sg13g2_nand2_1 _7363_ (.Y(_2541_),
    .A(_2416_),
    .B(_2540_));
 sg13g2_a21oi_1 _7364_ (.A1(_2537_),
    .A2(_2538_),
    .Y(_2542_),
    .B1(_2541_));
 sg13g2_o21ai_1 _7365_ (.B1(_2287_),
    .Y(_2543_),
    .A1(_1801_),
    .A2(_1802_));
 sg13g2_nand3_1 _7366_ (.B(_2276_),
    .C(_2543_),
    .A(_1996_),
    .Y(_2544_));
 sg13g2_o21ai_1 _7367_ (.B1(_2529_),
    .Y(_2545_),
    .A1(_2432_),
    .A2(_2420_));
 sg13g2_nand3_1 _7368_ (.B(net119),
    .C(net281),
    .A(net120),
    .Y(_2546_));
 sg13g2_o21ai_1 _7369_ (.B1(_3831_),
    .Y(_2547_),
    .A1(_2432_),
    .A2(_2529_));
 sg13g2_a22oi_1 _7370_ (.Y(_2548_),
    .B1(_2547_),
    .B2(net119),
    .A2(_2507_),
    .A1(net120));
 sg13g2_o21ai_1 _7371_ (.B1(_2548_),
    .Y(_2549_),
    .A1(_2420_),
    .A2(_2546_));
 sg13g2_a221oi_1 _7372_ (.B2(_3830_),
    .C1(_2549_),
    .B1(_2545_),
    .A1(_2542_),
    .Y(_2550_),
    .A2(_2544_));
 sg13g2_a21o_1 _7373_ (.A2(_1579_),
    .A1(_1577_),
    .B1(_1585_),
    .X(_2551_));
 sg13g2_nand3_1 _7374_ (.B(_1593_),
    .C(_2551_),
    .A(_0922_),
    .Y(_2552_));
 sg13g2_inv_1 _7375_ (.Y(_2553_),
    .A(_1615_));
 sg13g2_nor2_1 _7376_ (.A(_2289_),
    .B(_2541_),
    .Y(_2554_));
 sg13g2_o21ai_1 _7377_ (.B1(_2554_),
    .Y(_2555_),
    .A1(_2553_),
    .A2(_1608_));
 sg13g2_nand4_1 _7378_ (.B(_2550_),
    .C(_2552_),
    .A(_2536_),
    .Y(_2556_),
    .D(_2555_));
 sg13g2_nand2b_1 _7379_ (.Y(_2557_),
    .B(_2554_),
    .A_N(_2536_));
 sg13g2_nand2_1 _7380_ (.Y(_2558_),
    .A(_1559_),
    .B(_1560_));
 sg13g2_nand2_1 _7381_ (.Y(_2559_),
    .A(_0851_),
    .B(_1561_));
 sg13g2_nand2_1 _7382_ (.Y(_2560_),
    .A(_1564_),
    .B(_1566_));
 sg13g2_a221oi_1 _7383_ (.B2(_2560_),
    .C1(_2283_),
    .B1(_2559_),
    .A1(_0837_),
    .Y(_2561_),
    .A2(_1556_));
 sg13g2_a221oi_1 _7384_ (.B2(_2561_),
    .C1(_2294_),
    .B1(_2558_),
    .A1(_1570_),
    .Y(_2562_),
    .A2(_0879_));
 sg13g2_mux2_1 _7385_ (.A0(_2556_),
    .A1(_2557_),
    .S(_2562_),
    .X(_2563_));
 sg13g2_nor2_1 _7386_ (.A(_2553_),
    .B(_1608_),
    .Y(_2564_));
 sg13g2_a21o_1 _7387_ (.A2(_2552_),
    .A1(_2564_),
    .B1(_2557_),
    .X(_2565_));
 sg13g2_o21ai_1 _7388_ (.B1(_2536_),
    .Y(_2566_),
    .A1(_2289_),
    .A2(_2541_));
 sg13g2_mux2_1 _7389_ (.A0(_2536_),
    .A1(_2566_),
    .S(_2550_),
    .X(_2567_));
 sg13g2_and3_1 _7390_ (.X(_2568_),
    .A(net103),
    .B(_2565_),
    .C(_2567_));
 sg13g2_a22oi_1 _7391_ (.Y(_2569_),
    .B1(_2563_),
    .B2(_2568_),
    .A2(_2535_),
    .A1(net84));
 sg13g2_a21o_1 _7392_ (.A2(_2569_),
    .A1(_3971_),
    .B1(_3963_),
    .X(_2570_));
 sg13g2_a21oi_1 _7393_ (.A1(net59),
    .A2(_2534_),
    .Y(_0075_),
    .B1(_2570_));
 sg13g2_nor2b_1 _7394_ (.A(_1062_),
    .B_N(_1127_),
    .Y(_2571_));
 sg13g2_a221oi_1 _7395_ (.B2(_1137_),
    .C1(_1158_),
    .B1(_2571_),
    .A1(_1352_),
    .Y(_2572_),
    .A2(_1161_));
 sg13g2_nand2_1 _7396_ (.Y(_2573_),
    .A(_1114_),
    .B(_1635_));
 sg13g2_inv_1 _7397_ (.Y(_2574_),
    .A(_1150_));
 sg13g2_and3_1 _7398_ (.X(_2575_),
    .A(_4148_),
    .B(_3848_),
    .C(_4136_));
 sg13g2_and4_1 _7399_ (.A(net114),
    .B(_4154_),
    .C(net148),
    .D(_4133_),
    .X(_2576_));
 sg13g2_o21ai_1 _7400_ (.B1(_1165_),
    .Y(_2577_),
    .A1(_2575_),
    .A2(_2576_));
 sg13g2_a221oi_1 _7401_ (.B2(_2577_),
    .C1(_2157_),
    .B1(_2574_),
    .A1(_1104_),
    .Y(_2578_),
    .A2(_1106_));
 sg13g2_o21ai_1 _7402_ (.B1(_1635_),
    .Y(_2579_),
    .A1(_1126_),
    .A2(_2578_));
 sg13g2_o21ai_1 _7403_ (.B1(_2579_),
    .Y(_2580_),
    .A1(_2572_),
    .A2(_2573_));
 sg13g2_nand4_1 _7404_ (.B(net281),
    .C(_3833_),
    .A(net119),
    .Y(_2581_),
    .D(_2505_));
 sg13g2_nor2_1 _7405_ (.A(_3856_),
    .B(net281),
    .Y(_2582_));
 sg13g2_nand3_1 _7406_ (.B(_2507_),
    .C(_2582_),
    .A(_3832_),
    .Y(_2583_));
 sg13g2_a21o_1 _7407_ (.A2(_2583_),
    .A1(_2581_),
    .B1(_2439_),
    .X(_2584_));
 sg13g2_nor4_1 _7408_ (.A(_1814_),
    .B(_2016_),
    .C(_2310_),
    .D(_2584_),
    .Y(_2585_));
 sg13g2_o21ai_1 _7409_ (.B1(_2585_),
    .Y(_2586_),
    .A1(_1647_),
    .A2(_2580_));
 sg13g2_nor2_1 _7410_ (.A(_2015_),
    .B(_2326_),
    .Y(_2587_));
 sg13g2_o21ai_1 _7411_ (.B1(_2587_),
    .Y(_2588_),
    .A1(_1818_),
    .A2(_2016_));
 sg13g2_nor2_1 _7412_ (.A(_2133_),
    .B(_2144_),
    .Y(_2589_));
 sg13g2_o21ai_1 _7413_ (.B1(_2325_),
    .Y(_2590_),
    .A1(_2323_),
    .A2(_2589_));
 sg13g2_nor2b_1 _7414_ (.A(_2584_),
    .B_N(_2590_),
    .Y(_2591_));
 sg13g2_nand2_1 _7415_ (.Y(_2592_),
    .A(_3831_),
    .B(_3833_));
 sg13g2_o21ai_1 _7416_ (.B1(_2592_),
    .Y(_2593_),
    .A1(net281),
    .A2(_2448_));
 sg13g2_nand2_1 _7417_ (.Y(_2594_),
    .A(_3830_),
    .B(_3832_));
 sg13g2_a22oi_1 _7418_ (.Y(_2595_),
    .B1(_2594_),
    .B2(_2529_),
    .A2(_2593_),
    .A1(_2461_));
 sg13g2_nor2_1 _7419_ (.A(_2592_),
    .B(_2448_),
    .Y(_2596_));
 sg13g2_o21ai_1 _7420_ (.B1(_2432_),
    .Y(_2597_),
    .A1(_2582_),
    .A2(_2596_));
 sg13g2_a22oi_1 _7421_ (.Y(_2598_),
    .B1(_2595_),
    .B2(_2597_),
    .A2(_2591_),
    .A1(_2588_));
 sg13g2_nor4_2 _7422_ (.A(_1043_),
    .B(_1051_),
    .C(_1036_),
    .Y(_2599_),
    .D(_1057_));
 sg13g2_or2_1 _7423_ (.X(_2600_),
    .B(_1090_),
    .A(_1144_));
 sg13g2_nor3_1 _7424_ (.A(_1150_),
    .B(_1154_),
    .C(_1113_),
    .Y(_2601_));
 sg13g2_o21ai_1 _7425_ (.B1(_1628_),
    .Y(_2602_),
    .A1(_1625_),
    .A2(_2601_));
 sg13g2_nor4_1 _7426_ (.A(_1814_),
    .B(_2016_),
    .C(_2310_),
    .D(_2584_),
    .Y(_2603_));
 sg13g2_and4_1 _7427_ (.A(_1091_),
    .B(_1635_),
    .C(_2602_),
    .D(_2603_),
    .X(_2604_));
 sg13g2_o21ai_1 _7428_ (.B1(_2604_),
    .Y(_2605_),
    .A1(_2599_),
    .A2(_2600_));
 sg13g2_nand3_1 _7429_ (.B(_2598_),
    .C(_2605_),
    .A(_2586_),
    .Y(_2606_));
 sg13g2_xnor2_1 _7430_ (.Y(_2607_),
    .A(_3922_),
    .B(_3832_));
 sg13g2_xnor2_1 _7431_ (.Y(_2608_),
    .A(_2606_),
    .B(_2607_));
 sg13g2_nand3_1 _7432_ (.B(_3970_),
    .C(_2608_),
    .A(net52),
    .Y(_2609_));
 sg13g2_inv_1 _7433_ (.Y(_2610_),
    .A(_3922_));
 sg13g2_nand2_1 _7434_ (.Y(_2611_),
    .A(net324),
    .B(_2366_));
 sg13g2_o21ai_1 _7435_ (.B1(_2611_),
    .Y(_2612_),
    .A1(_2610_),
    .A2(net58));
 sg13g2_nand2_1 _7436_ (.Y(_2613_),
    .A(net60),
    .B(_2612_));
 sg13g2_a21oi_1 _7437_ (.A1(_2609_),
    .A2(_2613_),
    .Y(_0076_),
    .B1(_2371_));
 sg13g2_mux2_1 _7438_ (.A0(net222),
    .A1(net325),
    .S(_1552_),
    .X(_2614_));
 sg13g2_nor2_1 _7439_ (.A(net82),
    .B(_2614_),
    .Y(_2615_));
 sg13g2_xnor2_1 _7440_ (.Y(_2616_),
    .A(net250),
    .B(net222));
 sg13g2_xnor2_1 _7441_ (.Y(_2617_),
    .A(_0763_),
    .B(_2616_));
 sg13g2_nor2_1 _7442_ (.A(net34),
    .B(net234),
    .Y(_2618_));
 sg13g2_a21oi_1 _7443_ (.A1(net41),
    .A2(_2617_),
    .Y(_2619_),
    .B1(_2618_));
 sg13g2_nor2_1 _7444_ (.A(net60),
    .B(_2619_),
    .Y(_2620_));
 sg13g2_nor3_1 _7445_ (.A(_2080_),
    .B(_2615_),
    .C(_2620_),
    .Y(_0077_));
 sg13g2_buf_1 _7446_ (.A(net51),
    .X(_2621_));
 sg13g2_a21oi_1 _7447_ (.A1(_1022_),
    .A2(_1025_),
    .Y(_2622_),
    .B1(_1005_));
 sg13g2_xnor2_1 _7448_ (.Y(_2623_),
    .A(net234),
    .B(net222));
 sg13g2_xnor2_1 _7449_ (.Y(_2624_),
    .A(_2622_),
    .B(_2623_));
 sg13g2_nor2_1 _7450_ (.A(net38),
    .B(net164),
    .Y(_2625_));
 sg13g2_a21oi_1 _7451_ (.A1(net29),
    .A2(_2624_),
    .Y(_2626_),
    .B1(_2625_));
 sg13g2_nor2_1 _7452_ (.A(net65),
    .B(_2626_),
    .Y(_2627_));
 sg13g2_buf_1 _7453_ (.A(net78),
    .X(_2628_));
 sg13g2_nand2_1 _7454_ (.Y(_2629_),
    .A(net324),
    .B(net63));
 sg13g2_o21ai_1 _7455_ (.B1(_2629_),
    .Y(_2630_),
    .A1(_0235_),
    .A2(_1552_));
 sg13g2_nor2_1 _7456_ (.A(net56),
    .B(_2630_),
    .Y(_2631_));
 sg13g2_nor3_1 _7457_ (.A(_2080_),
    .B(_2627_),
    .C(_2631_),
    .Y(_0078_));
 sg13g2_nand2_1 _7458_ (.Y(_2632_),
    .A(_0274_),
    .B(_0278_));
 sg13g2_nand2_1 _7459_ (.Y(_2633_),
    .A(_0308_),
    .B(_2632_));
 sg13g2_nand2_1 _7460_ (.Y(_2634_),
    .A(_0232_),
    .B(_2633_));
 sg13g2_xor2_1 _7461_ (.B(_0448_),
    .A(net234),
    .X(_2635_));
 sg13g2_xnor2_1 _7462_ (.Y(_2636_),
    .A(_2634_),
    .B(_2635_));
 sg13g2_nor2_1 _7463_ (.A(net38),
    .B(net233),
    .Y(_2637_));
 sg13g2_a21oi_1 _7464_ (.A1(net29),
    .A2(_2636_),
    .Y(_2638_),
    .B1(_2637_));
 sg13g2_nor2_1 _7465_ (.A(net65),
    .B(_2638_),
    .Y(_2639_));
 sg13g2_xnor2_1 _7466_ (.Y(_2640_),
    .A(_3977_),
    .B(_0384_));
 sg13g2_nand3b_1 _7467_ (.B(_2640_),
    .C(_3975_),
    .Y(_2641_),
    .A_N(_3976_));
 sg13g2_buf_2 _7468_ (.A(_2641_),
    .X(_2642_));
 sg13g2_nor3_1 _7469_ (.A(_3978_),
    .B(_0383_),
    .C(net272),
    .Y(_2643_));
 sg13g2_nor2b_1 _7470_ (.A(_2642_),
    .B_N(_2643_),
    .Y(_2644_));
 sg13g2_buf_1 _7471_ (.A(_2644_),
    .X(_2645_));
 sg13g2_inv_2 _7472_ (.Y(_2646_),
    .A(_0395_));
 sg13g2_nor2_2 _7473_ (.A(_2646_),
    .B(_2644_),
    .Y(_2647_));
 sg13g2_a221oi_1 _7474_ (.B2(net164),
    .C1(net76),
    .B1(_2647_),
    .A1(net328),
    .Y(_2648_),
    .A2(net49));
 sg13g2_nor3_1 _7475_ (.A(net92),
    .B(_2639_),
    .C(_2648_),
    .Y(_0079_));
 sg13g2_xor2_1 _7476_ (.B(net164),
    .A(net233),
    .X(_2649_));
 sg13g2_xnor2_1 _7477_ (.Y(_2650_),
    .A(_1497_),
    .B(_2649_));
 sg13g2_nor2_1 _7478_ (.A(net38),
    .B(net181),
    .Y(_2651_));
 sg13g2_a21oi_1 _7479_ (.A1(net29),
    .A2(_2650_),
    .Y(_2652_),
    .B1(_2651_));
 sg13g2_nor2_1 _7480_ (.A(net65),
    .B(_2652_),
    .Y(_2653_));
 sg13g2_a221oi_1 _7481_ (.B2(net233),
    .C1(net76),
    .B1(_2647_),
    .A1(net274),
    .Y(_2654_),
    .A2(net49));
 sg13g2_nor3_1 _7482_ (.A(net92),
    .B(_2653_),
    .C(_2654_),
    .Y(_0080_));
 sg13g2_a22oi_1 _7483_ (.Y(_2655_),
    .B1(_0798_),
    .B2(_3837_),
    .A2(_0797_),
    .A1(_0448_));
 sg13g2_o21ai_1 _7484_ (.B1(_2655_),
    .Y(_2656_),
    .A1(_0763_),
    .A2(_0768_));
 sg13g2_xor2_1 _7485_ (.B(_0237_),
    .A(_3839_),
    .X(_2657_));
 sg13g2_xnor2_1 _7486_ (.Y(_2658_),
    .A(_2656_),
    .B(_2657_));
 sg13g2_nor2_1 _7487_ (.A(_0693_),
    .B(_0236_),
    .Y(_2659_));
 sg13g2_a21oi_1 _7488_ (.A1(_2621_),
    .A2(_2658_),
    .Y(_2660_),
    .B1(_2659_));
 sg13g2_nor2_1 _7489_ (.A(_0405_),
    .B(_2660_),
    .Y(_2661_));
 sg13g2_a221oi_1 _7490_ (.B2(net181),
    .C1(net76),
    .B1(_2647_),
    .A1(net262),
    .Y(_2662_),
    .A2(net49));
 sg13g2_nor3_1 _7491_ (.A(net92),
    .B(_2661_),
    .C(_2662_),
    .Y(_0081_));
 sg13g2_nor2_1 _7492_ (.A(_0500_),
    .B(net49),
    .Y(_2663_));
 sg13g2_a221oi_1 _7493_ (.B2(_0700_),
    .C1(_0706_),
    .B1(_2663_),
    .A1(net323),
    .Y(_2664_),
    .A2(_2645_));
 sg13g2_xor2_1 _7494_ (.B(_0237_),
    .A(net182),
    .X(_2665_));
 sg13g2_a21oi_1 _7495_ (.A1(_0997_),
    .A2(_0998_),
    .Y(_2666_),
    .B1(_2622_));
 sg13g2_nor2_1 _7496_ (.A(_1029_),
    .B(_2666_),
    .Y(_2667_));
 sg13g2_xnor2_1 _7497_ (.Y(_2668_),
    .A(_2665_),
    .B(_2667_));
 sg13g2_mux2_1 _7498_ (.A0(net112),
    .A1(_2668_),
    .S(_4046_),
    .X(_2669_));
 sg13g2_nor2_1 _7499_ (.A(_2084_),
    .B(_2669_),
    .Y(_2670_));
 sg13g2_nor3_1 _7500_ (.A(net92),
    .B(_2664_),
    .C(_2670_),
    .Y(_0082_));
 sg13g2_a21o_1 _7501_ (.A2(_0279_),
    .A1(_0308_),
    .B1(_0242_),
    .X(_2671_));
 sg13g2_buf_1 _7502_ (.A(_2671_),
    .X(_2672_));
 sg13g2_xor2_1 _7503_ (.B(_3910_),
    .A(_0236_),
    .X(_2673_));
 sg13g2_xnor2_1 _7504_ (.Y(_2674_),
    .A(_2672_),
    .B(_2673_));
 sg13g2_nor2_1 _7505_ (.A(_0693_),
    .B(_0432_),
    .Y(_2675_));
 sg13g2_a21oi_1 _7506_ (.A1(_2621_),
    .A2(_2674_),
    .Y(_2676_),
    .B1(_2675_));
 sg13g2_nor2_1 _7507_ (.A(_0405_),
    .B(_2676_),
    .Y(_2677_));
 sg13g2_a221oi_1 _7508_ (.B2(_3910_),
    .C1(net76),
    .B1(_2647_),
    .A1(net265),
    .Y(_2678_),
    .A2(net49));
 sg13g2_nor3_1 _7509_ (.A(net92),
    .B(_2677_),
    .C(_2678_),
    .Y(_0083_));
 sg13g2_buf_1 _7510_ (.A(_0404_),
    .X(_2679_));
 sg13g2_xnor2_1 _7511_ (.Y(_2680_),
    .A(net165),
    .B(net112));
 sg13g2_xnor2_1 _7512_ (.Y(_2681_),
    .A(_1498_),
    .B(_2680_));
 sg13g2_nor2_1 _7513_ (.A(net38),
    .B(net115),
    .Y(_2682_));
 sg13g2_a21oi_1 _7514_ (.A1(net29),
    .A2(_2681_),
    .Y(_2683_),
    .B1(_2682_));
 sg13g2_nor2_1 _7515_ (.A(_2679_),
    .B(_2683_),
    .Y(_2684_));
 sg13g2_a221oi_1 _7516_ (.B2(net165),
    .C1(_0704_),
    .B1(_2647_),
    .A1(net266),
    .Y(_2685_),
    .A2(net49));
 sg13g2_nor3_1 _7517_ (.A(net92),
    .B(_2684_),
    .C(_2685_),
    .Y(_0084_));
 sg13g2_nor2b_1 _7518_ (.A(net49),
    .B_N(_3761_),
    .Y(_2686_));
 sg13g2_a221oi_1 _7519_ (.B2(net18),
    .C1(_0706_),
    .B1(_2686_),
    .A1(net325),
    .Y(_2687_),
    .A2(_2645_));
 sg13g2_nor2_1 _7520_ (.A(_0763_),
    .B(_0768_),
    .Y(_2688_));
 sg13g2_a21o_1 _7521_ (.A2(_2688_),
    .A1(_0778_),
    .B1(_0806_),
    .X(_2689_));
 sg13g2_xor2_1 _7522_ (.B(net115),
    .A(_0432_),
    .X(_2690_));
 sg13g2_xnor2_1 _7523_ (.Y(_2691_),
    .A(_2689_),
    .B(_2690_));
 sg13g2_nor2_1 _7524_ (.A(net34),
    .B(net255),
    .Y(_2692_));
 sg13g2_a21oi_1 _7525_ (.A1(net41),
    .A2(_2691_),
    .Y(_2693_),
    .B1(_2692_));
 sg13g2_nor2_1 _7526_ (.A(_2084_),
    .B(_2693_),
    .Y(_2694_));
 sg13g2_nor3_1 _7527_ (.A(net92),
    .B(_2687_),
    .C(_2694_),
    .Y(_0085_));
 sg13g2_buf_1 _7528_ (.A(_3964_),
    .X(_2695_));
 sg13g2_xnor2_1 _7529_ (.Y(_2696_),
    .A(net255),
    .B(net115));
 sg13g2_xnor2_1 _7530_ (.Y(_2697_),
    .A(_1036_),
    .B(_2696_));
 sg13g2_nor2_1 _7531_ (.A(net38),
    .B(net110),
    .Y(_2698_));
 sg13g2_a21oi_1 _7532_ (.A1(net29),
    .A2(_2697_),
    .Y(_2699_),
    .B1(_2698_));
 sg13g2_nor2_1 _7533_ (.A(_2679_),
    .B(_2699_),
    .Y(_2700_));
 sg13g2_a221oi_1 _7534_ (.B2(net255),
    .C1(_0704_),
    .B1(_2647_),
    .A1(net263),
    .Y(_2701_),
    .A2(net49));
 sg13g2_nor3_1 _7535_ (.A(net89),
    .B(_2700_),
    .C(_2701_),
    .Y(_0086_));
 sg13g2_a21o_1 _7536_ (.A2(_2672_),
    .A1(net112),
    .B1(net255),
    .X(_2702_));
 sg13g2_nand2_1 _7537_ (.Y(_2703_),
    .A(net112),
    .B(_3761_));
 sg13g2_nand2b_1 _7538_ (.Y(_2704_),
    .B(_2672_),
    .A_N(_0515_));
 sg13g2_a21oi_1 _7539_ (.A1(_2703_),
    .A2(_2704_),
    .Y(_2705_),
    .B1(_0500_));
 sg13g2_a221oi_1 _7540_ (.B2(net115),
    .C1(_2705_),
    .B1(_2702_),
    .A1(net165),
    .Y(_2706_),
    .A2(_0310_));
 sg13g2_xor2_1 _7541_ (.B(_3926_),
    .A(net255),
    .X(_2707_));
 sg13g2_xnor2_1 _7542_ (.Y(_2708_),
    .A(_2706_),
    .B(_2707_));
 sg13g2_nand2_1 _7543_ (.Y(_2709_),
    .A(net34),
    .B(_2708_));
 sg13g2_o21ai_1 _7544_ (.B1(_2709_),
    .Y(_2710_),
    .A1(_4034_),
    .A2(_0770_));
 sg13g2_nand2_1 _7545_ (.Y(_2711_),
    .A(net61),
    .B(_2710_));
 sg13g2_nand3b_1 _7546_ (.B(net329),
    .C(_3978_),
    .Y(_2712_),
    .A_N(net272));
 sg13g2_nor2_1 _7547_ (.A(_2642_),
    .B(_2712_),
    .Y(_2713_));
 sg13g2_buf_1 _7548_ (.A(_2713_),
    .X(_2714_));
 sg13g2_mux2_1 _7549_ (.A0(_3926_),
    .A1(_1234_),
    .S(net48),
    .X(_2715_));
 sg13g2_nand2_1 _7550_ (.Y(_2716_),
    .A(net60),
    .B(_2715_));
 sg13g2_a21oi_1 _7551_ (.A1(_2711_),
    .A2(_2716_),
    .Y(_0087_),
    .B1(_2371_));
 sg13g2_and3_1 _7552_ (.X(_2717_),
    .A(_1264_),
    .B(_1266_),
    .C(_1267_));
 sg13g2_xnor2_1 _7553_ (.Y(_2718_),
    .A(net220),
    .B(net110));
 sg13g2_xnor2_1 _7554_ (.Y(_2719_),
    .A(_2717_),
    .B(_2718_));
 sg13g2_nor2_1 _7555_ (.A(net38),
    .B(_0313_),
    .Y(_2720_));
 sg13g2_a21oi_1 _7556_ (.A1(net29),
    .A2(_2719_),
    .Y(_2721_),
    .B1(_2720_));
 sg13g2_nor2_1 _7557_ (.A(net55),
    .B(_2721_),
    .Y(_2722_));
 sg13g2_nor2_2 _7558_ (.A(_2646_),
    .B(_2714_),
    .Y(_2723_));
 sg13g2_buf_1 _7559_ (.A(net104),
    .X(_2724_));
 sg13g2_a221oi_1 _7560_ (.B2(net220),
    .C1(net74),
    .B1(_2723_),
    .A1(_1324_),
    .Y(_2725_),
    .A2(net48));
 sg13g2_nor3_1 _7561_ (.A(_2695_),
    .B(_2722_),
    .C(_2725_),
    .Y(_0088_));
 sg13g2_nand2b_1 _7562_ (.Y(_2726_),
    .B(_0796_),
    .A_N(_1559_));
 sg13g2_xor2_1 _7563_ (.B(net176),
    .A(net220),
    .X(_2727_));
 sg13g2_xnor2_1 _7564_ (.Y(_2728_),
    .A(_2726_),
    .B(_2727_));
 sg13g2_buf_1 _7565_ (.A(_0692_),
    .X(_2729_));
 sg13g2_nor2_1 _7566_ (.A(net28),
    .B(net241),
    .Y(_2730_));
 sg13g2_a21oi_1 _7567_ (.A1(net29),
    .A2(_2728_),
    .Y(_2731_),
    .B1(_2730_));
 sg13g2_nor2_1 _7568_ (.A(net55),
    .B(_2731_),
    .Y(_2732_));
 sg13g2_a221oi_1 _7569_ (.B2(_0313_),
    .C1(net74),
    .B1(_2723_),
    .A1(_1348_),
    .Y(_2733_),
    .A2(net48));
 sg13g2_nor3_1 _7570_ (.A(net89),
    .B(_2732_),
    .C(_2733_),
    .Y(_0089_));
 sg13g2_nand2_1 _7571_ (.Y(_2734_),
    .A(_1084_),
    .B(_1086_));
 sg13g2_nor2_1 _7572_ (.A(_1036_),
    .B(_1056_),
    .Y(_2735_));
 sg13g2_nor2_1 _7573_ (.A(_2734_),
    .B(_2735_),
    .Y(_2736_));
 sg13g2_xor2_1 _7574_ (.B(net176),
    .A(net241),
    .X(_2737_));
 sg13g2_xnor2_1 _7575_ (.Y(_2738_),
    .A(_2736_),
    .B(_2737_));
 sg13g2_mux2_1 _7576_ (.A0(net175),
    .A1(_2738_),
    .S(_1687_),
    .X(_2739_));
 sg13g2_nor2_1 _7577_ (.A(net55),
    .B(_2739_),
    .Y(_2740_));
 sg13g2_a221oi_1 _7578_ (.B2(net241),
    .C1(net74),
    .B1(_2723_),
    .A1(_1422_),
    .Y(_2741_),
    .A2(net48));
 sg13g2_nor3_1 _7579_ (.A(net89),
    .B(_2740_),
    .C(_2741_),
    .Y(_0090_));
 sg13g2_mux2_1 _7580_ (.A0(net175),
    .A1(net327),
    .S(net48),
    .X(_2742_));
 sg13g2_nor2_1 _7581_ (.A(net82),
    .B(_2742_),
    .Y(_2743_));
 sg13g2_a21oi_1 _7582_ (.A1(_0255_),
    .A2(_2672_),
    .Y(_2744_),
    .B1(_1460_));
 sg13g2_xnor2_1 _7583_ (.Y(_2745_),
    .A(_3792_),
    .B(net175));
 sg13g2_xnor2_1 _7584_ (.Y(_2746_),
    .A(_2744_),
    .B(_2745_));
 sg13g2_nor2_1 _7585_ (.A(net36),
    .B(net247),
    .Y(_2747_));
 sg13g2_a21oi_1 _7586_ (.A1(net41),
    .A2(_2746_),
    .Y(_2748_),
    .B1(_2747_));
 sg13g2_nor2_1 _7587_ (.A(net60),
    .B(_2748_),
    .Y(_2749_));
 sg13g2_nor3_1 _7588_ (.A(_2695_),
    .B(_2743_),
    .C(_2749_),
    .Y(_0091_));
 sg13g2_or2_1 _7589_ (.X(_2750_),
    .B(_0265_),
    .A(_0259_));
 sg13g2_xnor2_1 _7590_ (.Y(_2751_),
    .A(_1500_),
    .B(_2750_));
 sg13g2_nor2_1 _7591_ (.A(net28),
    .B(net240),
    .Y(_2752_));
 sg13g2_a21oi_1 _7592_ (.A1(net29),
    .A2(_2751_),
    .Y(_2753_),
    .B1(_2752_));
 sg13g2_nor2_1 _7593_ (.A(net55),
    .B(_2753_),
    .Y(_2754_));
 sg13g2_a221oi_1 _7594_ (.B2(net247),
    .C1(net74),
    .B1(_2723_),
    .A1(net266),
    .Y(_2755_),
    .A2(net48));
 sg13g2_nor3_1 _7595_ (.A(net89),
    .B(_2754_),
    .C(_2755_),
    .Y(_0092_));
 sg13g2_mux2_1 _7596_ (.A0(net262),
    .A1(net257),
    .S(_3988_),
    .X(_2756_));
 sg13g2_nor2b_1 _7597_ (.A(net284),
    .B_N(net257),
    .Y(_2757_));
 sg13g2_nor2_1 _7598_ (.A(_4036_),
    .B(net257),
    .Y(_2758_));
 sg13g2_nor3_1 _7599_ (.A(net84),
    .B(_2757_),
    .C(_2758_),
    .Y(_2759_));
 sg13g2_a21oi_1 _7600_ (.A1(_3969_),
    .A2(net249),
    .Y(_2760_),
    .B1(_2759_));
 sg13g2_nor2_1 _7601_ (.A(net77),
    .B(_2760_),
    .Y(_2761_));
 sg13g2_a21oi_1 _7602_ (.A1(net59),
    .A2(_2756_),
    .Y(_2762_),
    .B1(_2761_));
 sg13g2_nor2_1 _7603_ (.A(net90),
    .B(_2762_),
    .Y(_0093_));
 sg13g2_buf_1 _7604_ (.A(net51),
    .X(_2763_));
 sg13g2_nand2_1 _7605_ (.Y(_2764_),
    .A(_0789_),
    .B(_0790_));
 sg13g2_a21o_1 _7606_ (.A2(_2726_),
    .A1(_2764_),
    .B1(_1562_),
    .X(_2765_));
 sg13g2_buf_1 _7607_ (.A(_2765_),
    .X(_2766_));
 sg13g2_xor2_1 _7608_ (.B(net240),
    .A(net247),
    .X(_2767_));
 sg13g2_xnor2_1 _7609_ (.Y(_2768_),
    .A(_2766_),
    .B(_2767_));
 sg13g2_nor2_1 _7610_ (.A(net28),
    .B(net246),
    .Y(_2769_));
 sg13g2_a21oi_1 _7611_ (.A1(net27),
    .A2(_2768_),
    .Y(_2770_),
    .B1(_2769_));
 sg13g2_nor2_1 _7612_ (.A(net55),
    .B(_2770_),
    .Y(_2771_));
 sg13g2_a221oi_1 _7613_ (.B2(net240),
    .C1(_2724_),
    .B1(_2723_),
    .A1(net264),
    .Y(_2772_),
    .A2(net48));
 sg13g2_nor3_1 _7614_ (.A(net89),
    .B(_2771_),
    .C(_2772_),
    .Y(_0094_));
 sg13g2_a21o_1 _7615_ (.A2(_2735_),
    .A1(_1355_),
    .B1(_1358_),
    .X(_2773_));
 sg13g2_nor2_1 _7616_ (.A(_0257_),
    .B(_0263_),
    .Y(_2774_));
 sg13g2_xor2_1 _7617_ (.B(_2774_),
    .A(_2773_),
    .X(_2775_));
 sg13g2_nor2_1 _7618_ (.A(_2729_),
    .B(net226),
    .Y(_2776_));
 sg13g2_a21oi_1 _7619_ (.A1(net27),
    .A2(_2775_),
    .Y(_2777_),
    .B1(_2776_));
 sg13g2_nor2_1 _7620_ (.A(net55),
    .B(_2777_),
    .Y(_2778_));
 sg13g2_a221oi_1 _7621_ (.B2(net246),
    .C1(_2724_),
    .B1(_2723_),
    .A1(net263),
    .Y(_2779_),
    .A2(net48));
 sg13g2_nor3_1 _7622_ (.A(net89),
    .B(_2778_),
    .C(_2779_),
    .Y(_0095_));
 sg13g2_xnor2_1 _7623_ (.Y(_2780_),
    .A(net246),
    .B(net226));
 sg13g2_xnor2_1 _7624_ (.Y(_2781_),
    .A(_0324_),
    .B(_2780_));
 sg13g2_nor2_1 _7625_ (.A(_2729_),
    .B(net215),
    .Y(_2782_));
 sg13g2_a21oi_1 _7626_ (.A1(_2763_),
    .A2(_2781_),
    .Y(_2783_),
    .B1(_2782_));
 sg13g2_nor2_1 _7627_ (.A(net55),
    .B(_2783_),
    .Y(_2784_));
 sg13g2_nor3_1 _7628_ (.A(net273),
    .B(_1240_),
    .C(_2642_),
    .Y(_2785_));
 sg13g2_buf_1 _7629_ (.A(_2785_),
    .X(_2786_));
 sg13g2_mux2_1 _7630_ (.A0(net226),
    .A1(_4028_),
    .S(_2786_),
    .X(_2787_));
 sg13g2_nor2_1 _7631_ (.A(net56),
    .B(_2787_),
    .Y(_2788_));
 sg13g2_nor3_1 _7632_ (.A(net89),
    .B(_2784_),
    .C(_2788_),
    .Y(_0096_));
 sg13g2_o21ai_1 _7633_ (.B1(_1261_),
    .Y(_2789_),
    .A1(_2717_),
    .A2(_1270_));
 sg13g2_nor2_1 _7634_ (.A(_0205_),
    .B(_0490_),
    .Y(_2790_));
 sg13g2_xor2_1 _7635_ (.B(_2790_),
    .A(_2789_),
    .X(_2791_));
 sg13g2_nor2_1 _7636_ (.A(net28),
    .B(net225),
    .Y(_2792_));
 sg13g2_a21oi_1 _7637_ (.A1(_2763_),
    .A2(_2791_),
    .Y(_2793_),
    .B1(_2792_));
 sg13g2_nor2_1 _7638_ (.A(net55),
    .B(_2793_),
    .Y(_2794_));
 sg13g2_nor2_1 _7639_ (.A(_2646_),
    .B(_2785_),
    .Y(_2795_));
 sg13g2_a221oi_1 _7640_ (.B2(net215),
    .C1(net74),
    .B1(_2795_),
    .A1(net274),
    .Y(_2796_),
    .A2(net47));
 sg13g2_nor3_1 _7641_ (.A(net89),
    .B(_2794_),
    .C(_2796_),
    .Y(_0097_));
 sg13g2_xnor2_1 _7642_ (.Y(_2797_),
    .A(net215),
    .B(net225));
 sg13g2_nand2_1 _7643_ (.Y(_2798_),
    .A(_0783_),
    .B(_0784_));
 sg13g2_inv_1 _7644_ (.Y(_2799_),
    .A(_0866_));
 sg13g2_a21oi_1 _7645_ (.A1(_2798_),
    .A2(_2766_),
    .Y(_2800_),
    .B1(_2799_));
 sg13g2_xnor2_1 _7646_ (.Y(_2801_),
    .A(_2797_),
    .B(_2800_));
 sg13g2_nor2_1 _7647_ (.A(net68),
    .B(_2801_),
    .Y(_2802_));
 sg13g2_a21oi_1 _7648_ (.A1(net68),
    .A2(net239),
    .Y(_2803_),
    .B1(_2802_));
 sg13g2_nor2b_1 _7649_ (.A(_2785_),
    .B_N(net225),
    .Y(_2804_));
 sg13g2_a221oi_1 _7650_ (.B2(_0396_),
    .C1(net78),
    .B1(_2804_),
    .A1(net262),
    .Y(_2805_),
    .A2(net47));
 sg13g2_a21oi_1 _7651_ (.A1(_4045_),
    .A2(_2803_),
    .Y(_2806_),
    .B1(_2805_));
 sg13g2_and2_1 _7652_ (.A(net201),
    .B(_2806_),
    .X(_0098_));
 sg13g2_buf_1 _7653_ (.A(_3964_),
    .X(_2807_));
 sg13g2_buf_1 _7654_ (.A(net109),
    .X(_2808_));
 sg13g2_nor2_1 _7655_ (.A(_0204_),
    .B(_0491_),
    .Y(_2809_));
 sg13g2_xnor2_1 _7656_ (.Y(_2810_),
    .A(_1360_),
    .B(_2809_));
 sg13g2_mux2_1 _7657_ (.A0(net232),
    .A1(_2810_),
    .S(net34),
    .X(_2811_));
 sg13g2_nor2_1 _7658_ (.A(net73),
    .B(_2811_),
    .Y(_2812_));
 sg13g2_a221oi_1 _7659_ (.B2(net239),
    .C1(net74),
    .B1(_2795_),
    .A1(net323),
    .Y(_2813_),
    .A2(_2786_));
 sg13g2_nor3_1 _7660_ (.A(_2807_),
    .B(_2812_),
    .C(_2813_),
    .Y(_0099_));
 sg13g2_o21ai_1 _7661_ (.B1(_4201_),
    .Y(_2814_),
    .A1(_1465_),
    .A2(_0324_));
 sg13g2_xor2_1 _7662_ (.B(net232),
    .A(_3796_),
    .X(_2815_));
 sg13g2_xnor2_1 _7663_ (.Y(_2816_),
    .A(_2814_),
    .B(_2815_));
 sg13g2_nor2_1 _7664_ (.A(net28),
    .B(_3930_),
    .Y(_2817_));
 sg13g2_a21oi_1 _7665_ (.A1(net27),
    .A2(_2816_),
    .Y(_2818_),
    .B1(_2817_));
 sg13g2_nor2_1 _7666_ (.A(_2808_),
    .B(_2818_),
    .Y(_2819_));
 sg13g2_a221oi_1 _7667_ (.B2(net232),
    .C1(net74),
    .B1(_2795_),
    .A1(net265),
    .Y(_2820_),
    .A2(net47));
 sg13g2_nor3_1 _7668_ (.A(_2807_),
    .B(_2819_),
    .C(_2820_),
    .Y(_0100_));
 sg13g2_or2_1 _7669_ (.X(_2821_),
    .B(_4197_),
    .A(_4194_));
 sg13g2_xnor2_1 _7670_ (.Y(_2822_),
    .A(_0525_),
    .B(_2821_));
 sg13g2_nand2_1 _7671_ (.Y(_2823_),
    .A(net34),
    .B(_2822_));
 sg13g2_o21ai_1 _7672_ (.B1(_2823_),
    .Y(_2824_),
    .A1(net42),
    .A2(_4196_));
 sg13g2_a22oi_1 _7673_ (.Y(_2825_),
    .B1(_2795_),
    .B2(net214),
    .A2(net47),
    .A1(net326));
 sg13g2_nor2_1 _7674_ (.A(net75),
    .B(_2825_),
    .Y(_2826_));
 sg13g2_a21oi_1 _7675_ (.A1(_2466_),
    .A2(_2824_),
    .Y(_2827_),
    .B1(_2826_));
 sg13g2_nor2_1 _7676_ (.A(net90),
    .B(_2827_),
    .Y(_0101_));
 sg13g2_xnor2_1 _7677_ (.Y(_2828_),
    .A(net214),
    .B(_3843_));
 sg13g2_nand2_1 _7678_ (.Y(_2829_),
    .A(_0859_),
    .B(_1565_));
 sg13g2_a21oi_1 _7679_ (.A1(_0786_),
    .A2(_2766_),
    .Y(_2830_),
    .B1(_2829_));
 sg13g2_xnor2_1 _7680_ (.Y(_2831_),
    .A(_2828_),
    .B(_2830_));
 sg13g2_nor2_1 _7681_ (.A(net28),
    .B(net161),
    .Y(_2832_));
 sg13g2_a21oi_1 _7682_ (.A1(net27),
    .A2(_2831_),
    .Y(_2833_),
    .B1(_2832_));
 sg13g2_nor2_1 _7683_ (.A(_2808_),
    .B(_2833_),
    .Y(_2834_));
 sg13g2_nor2_1 _7684_ (.A(_4196_),
    .B(net47),
    .Y(_2835_));
 sg13g2_a221oi_1 _7685_ (.B2(_0700_),
    .C1(net74),
    .B1(_2835_),
    .A1(net264),
    .Y(_2836_),
    .A2(net47));
 sg13g2_nor3_1 _7686_ (.A(net88),
    .B(_2834_),
    .C(_2836_),
    .Y(_0102_));
 sg13g2_xor2_1 _7687_ (.B(net231),
    .A(net161),
    .X(_2837_));
 sg13g2_inv_1 _7688_ (.Y(_2838_),
    .A(_2773_));
 sg13g2_o21ai_1 _7689_ (.B1(_1080_),
    .Y(_2839_),
    .A1(_1051_),
    .A2(_2838_));
 sg13g2_xnor2_1 _7690_ (.Y(_2840_),
    .A(_2837_),
    .B(_2839_));
 sg13g2_nand2_1 _7691_ (.Y(_2841_),
    .A(net50),
    .B(_2840_));
 sg13g2_o21ai_1 _7692_ (.B1(_2841_),
    .Y(_2842_),
    .A1(net40),
    .A2(net160));
 sg13g2_nor2_1 _7693_ (.A(_4192_),
    .B(net47),
    .Y(_2843_));
 sg13g2_a221oi_1 _7694_ (.B2(net19),
    .C1(net78),
    .B1(_2843_),
    .A1(net324),
    .Y(_2844_),
    .A2(net47));
 sg13g2_a21oi_1 _7695_ (.A1(net79),
    .A2(_2842_),
    .Y(_2845_),
    .B1(_2844_));
 sg13g2_and2_1 _7696_ (.A(net201),
    .B(_2845_),
    .X(_0103_));
 sg13g2_xnor2_1 _7697_ (.Y(_2846_),
    .A(net249),
    .B(_2758_));
 sg13g2_nor2_1 _7698_ (.A(net28),
    .B(_3711_),
    .Y(_2847_));
 sg13g2_a21oi_1 _7699_ (.A1(net27),
    .A2(_2846_),
    .Y(_2848_),
    .B1(_2847_));
 sg13g2_nor2_1 _7700_ (.A(net73),
    .B(_2848_),
    .Y(_2849_));
 sg13g2_mux2_1 _7701_ (.A0(net323),
    .A1(_3758_),
    .S(_3988_),
    .X(_2850_));
 sg13g2_nor2_1 _7702_ (.A(net56),
    .B(_2850_),
    .Y(_2851_));
 sg13g2_nor3_1 _7703_ (.A(net88),
    .B(_2849_),
    .C(_2851_),
    .Y(_0104_));
 sg13g2_xor2_1 _7704_ (.B(net160),
    .A(net161),
    .X(_2852_));
 sg13g2_inv_1 _7705_ (.Y(_2853_),
    .A(_2814_));
 sg13g2_o21ai_1 _7706_ (.B1(_4206_),
    .Y(_2854_),
    .A1(_1468_),
    .A2(_2853_));
 sg13g2_xnor2_1 _7707_ (.Y(_2855_),
    .A(_2852_),
    .B(_2854_));
 sg13g2_nand2_1 _7708_ (.Y(_2856_),
    .A(net50),
    .B(_2855_));
 sg13g2_o21ai_1 _7709_ (.B1(_2856_),
    .Y(_2857_),
    .A1(net40),
    .A2(net159));
 sg13g2_nor2_1 _7710_ (.A(_1235_),
    .B(_2642_),
    .Y(_2858_));
 sg13g2_buf_1 _7711_ (.A(_2858_),
    .X(_2859_));
 sg13g2_nor2_1 _7712_ (.A(_0538_),
    .B(net46),
    .Y(_2860_));
 sg13g2_a221oi_1 _7713_ (.B2(_0396_),
    .C1(net78),
    .B1(_2860_),
    .A1(_1234_),
    .Y(_2861_),
    .A2(net46));
 sg13g2_a21oi_1 _7714_ (.A1(net79),
    .A2(_2857_),
    .Y(_2862_),
    .B1(_2861_));
 sg13g2_and2_1 _7715_ (.A(net201),
    .B(_2862_),
    .X(_0105_));
 sg13g2_xor2_1 _7716_ (.B(_0570_),
    .A(_0574_),
    .X(_2863_));
 sg13g2_inv_1 _7717_ (.Y(_2864_),
    .A(_2789_));
 sg13g2_o21ai_1 _7718_ (.B1(_1262_),
    .Y(_2865_),
    .A1(_1256_),
    .A2(_2864_));
 sg13g2_xnor2_1 _7719_ (.Y(_2866_),
    .A(_2863_),
    .B(_2865_));
 sg13g2_nor2_1 _7720_ (.A(net28),
    .B(net158),
    .Y(_2867_));
 sg13g2_a21oi_1 _7721_ (.A1(net27),
    .A2(_2866_),
    .Y(_2868_),
    .B1(_2867_));
 sg13g2_nor2_1 _7722_ (.A(net73),
    .B(_2868_),
    .Y(_2869_));
 sg13g2_nor2_1 _7723_ (.A(_0575_),
    .B(net46),
    .Y(_2870_));
 sg13g2_buf_1 _7724_ (.A(net104),
    .X(_2871_));
 sg13g2_a221oi_1 _7725_ (.B2(net18),
    .C1(net72),
    .B1(_2870_),
    .A1(_1324_),
    .Y(_2872_),
    .A2(_2859_));
 sg13g2_nor3_1 _7726_ (.A(net88),
    .B(_2869_),
    .C(_2872_),
    .Y(_0106_));
 sg13g2_nand2b_1 _7727_ (.Y(_2873_),
    .B(_0872_),
    .A_N(_0869_));
 sg13g2_nor3_2 _7728_ (.A(_2873_),
    .B(_0793_),
    .C(_0808_),
    .Y(_2874_));
 sg13g2_xnor2_1 _7729_ (.Y(_2875_),
    .A(net159),
    .B(net158));
 sg13g2_xnor2_1 _7730_ (.Y(_2876_),
    .A(_2874_),
    .B(_2875_));
 sg13g2_buf_1 _7731_ (.A(net67),
    .X(_2877_));
 sg13g2_nor2_1 _7732_ (.A(net45),
    .B(net186),
    .Y(_2878_));
 sg13g2_a21oi_1 _7733_ (.A1(net27),
    .A2(_2876_),
    .Y(_2879_),
    .B1(_2878_));
 sg13g2_nor2_1 _7734_ (.A(net73),
    .B(_2879_),
    .Y(_2880_));
 sg13g2_nor2_2 _7735_ (.A(_2646_),
    .B(_2858_),
    .Y(_2881_));
 sg13g2_a221oi_1 _7736_ (.B2(net158),
    .C1(net72),
    .B1(_2881_),
    .A1(_1348_),
    .Y(_2882_),
    .A2(_2859_));
 sg13g2_nor3_1 _7737_ (.A(net88),
    .B(_2880_),
    .C(_2882_),
    .Y(_0107_));
 sg13g2_a21oi_1 _7738_ (.A1(_1050_),
    .A2(_1083_),
    .Y(_2883_),
    .B1(_1076_));
 sg13g2_nand2_1 _7739_ (.Y(_2884_),
    .A(_2883_),
    .B(_1356_));
 sg13g2_nand3_1 _7740_ (.B(_1047_),
    .C(_2884_),
    .A(_1042_),
    .Y(_2885_));
 sg13g2_a21oi_1 _7741_ (.A1(_2883_),
    .A2(_2736_),
    .Y(_2886_),
    .B1(_2885_));
 sg13g2_nor2_1 _7742_ (.A(_1364_),
    .B(_2886_),
    .Y(_2887_));
 sg13g2_xnor2_1 _7743_ (.Y(_2888_),
    .A(net186),
    .B(net158));
 sg13g2_xnor2_1 _7744_ (.Y(_2889_),
    .A(_2887_),
    .B(_2888_));
 sg13g2_nor2_1 _7745_ (.A(net45),
    .B(_3704_),
    .Y(_2890_));
 sg13g2_a21oi_1 _7746_ (.A1(net27),
    .A2(_2889_),
    .Y(_2891_),
    .B1(_2890_));
 sg13g2_nor2_1 _7747_ (.A(net73),
    .B(_2891_),
    .Y(_2892_));
 sg13g2_a221oi_1 _7748_ (.B2(net186),
    .C1(_2871_),
    .B1(_2881_),
    .A1(_1422_),
    .Y(_2893_),
    .A2(net46));
 sg13g2_nor3_1 _7749_ (.A(net88),
    .B(_2892_),
    .C(_2893_),
    .Y(_0108_));
 sg13g2_buf_1 _7750_ (.A(net52),
    .X(_2894_));
 sg13g2_xor2_1 _7751_ (.B(net259),
    .A(net186),
    .X(_2895_));
 sg13g2_xnor2_1 _7752_ (.Y(_2896_),
    .A(_2183_),
    .B(_2895_));
 sg13g2_nor2_1 _7753_ (.A(_2877_),
    .B(net184),
    .Y(_2897_));
 sg13g2_a21oi_1 _7754_ (.A1(_2894_),
    .A2(_2896_),
    .Y(_2898_),
    .B1(_2897_));
 sg13g2_nor2_1 _7755_ (.A(net73),
    .B(_2898_),
    .Y(_2899_));
 sg13g2_a221oi_1 _7756_ (.B2(net259),
    .C1(net72),
    .B1(_2881_),
    .A1(net265),
    .Y(_2900_),
    .A2(net46));
 sg13g2_nor3_1 _7757_ (.A(net88),
    .B(_2899_),
    .C(_2900_),
    .Y(_0109_));
 sg13g2_o21ai_1 _7758_ (.B1(_1490_),
    .Y(_2901_),
    .A1(_0525_),
    .A2(_1489_));
 sg13g2_xor2_1 _7759_ (.B(net259),
    .A(net184),
    .X(_2902_));
 sg13g2_xnor2_1 _7760_ (.Y(_2903_),
    .A(_2901_),
    .B(_2902_));
 sg13g2_nor2_1 _7761_ (.A(_2877_),
    .B(net258),
    .Y(_2904_));
 sg13g2_a21oi_1 _7762_ (.A1(_2894_),
    .A2(_2903_),
    .Y(_2905_),
    .B1(_2904_));
 sg13g2_nor2_1 _7763_ (.A(net73),
    .B(_2905_),
    .Y(_2906_));
 sg13g2_a221oi_1 _7764_ (.B2(net184),
    .C1(net72),
    .B1(_2881_),
    .A1(net326),
    .Y(_2907_),
    .A2(net46));
 sg13g2_nor3_1 _7765_ (.A(net88),
    .B(_2906_),
    .C(_2907_),
    .Y(_0110_));
 sg13g2_o21ai_1 _7766_ (.B1(_0819_),
    .Y(_2908_),
    .A1(_0888_),
    .A2(_2874_));
 sg13g2_xor2_1 _7767_ (.B(net258),
    .A(net184),
    .X(_2909_));
 sg13g2_xnor2_1 _7768_ (.Y(_2910_),
    .A(_2908_),
    .B(_2909_));
 sg13g2_nor2_1 _7769_ (.A(net84),
    .B(_2910_),
    .Y(_2911_));
 sg13g2_a21oi_1 _7770_ (.A1(net68),
    .A2(net185),
    .Y(_2912_),
    .B1(_2911_));
 sg13g2_a221oi_1 _7771_ (.B2(net258),
    .C1(net78),
    .B1(_2881_),
    .A1(net325),
    .Y(_2913_),
    .A2(net46));
 sg13g2_a21oi_1 _7772_ (.A1(net79),
    .A2(_2912_),
    .Y(_2914_),
    .B1(_2913_));
 sg13g2_and2_1 _7773_ (.A(net201),
    .B(_2914_),
    .X(_0111_));
 sg13g2_nor2_2 _7774_ (.A(_2599_),
    .B(_2600_),
    .Y(_2915_));
 sg13g2_xnor2_1 _7775_ (.Y(_2916_),
    .A(net185),
    .B(net258));
 sg13g2_xnor2_1 _7776_ (.Y(_2917_),
    .A(_2915_),
    .B(_2916_));
 sg13g2_nor2_1 _7777_ (.A(net45),
    .B(net183),
    .Y(_2918_));
 sg13g2_a21oi_1 _7778_ (.A1(net26),
    .A2(_2917_),
    .Y(_2919_),
    .B1(_2918_));
 sg13g2_nor2_1 _7779_ (.A(net73),
    .B(_2919_),
    .Y(_2920_));
 sg13g2_a221oi_1 _7780_ (.B2(net185),
    .C1(_2871_),
    .B1(_2881_),
    .A1(net263),
    .Y(_2921_),
    .A2(net46));
 sg13g2_nor3_1 _7781_ (.A(net88),
    .B(_2920_),
    .C(_2921_),
    .Y(_0112_));
 sg13g2_buf_1 _7782_ (.A(_3963_),
    .X(_2922_));
 sg13g2_buf_1 _7783_ (.A(net109),
    .X(_2923_));
 sg13g2_xnor2_1 _7784_ (.Y(_2924_),
    .A(net185),
    .B(net183));
 sg13g2_and2_1 _7785_ (.A(_4216_),
    .B(_0209_),
    .X(_2925_));
 sg13g2_nor2b_1 _7786_ (.A(_0324_),
    .B_N(_2925_),
    .Y(_2926_));
 sg13g2_nor3_1 _7787_ (.A(_0215_),
    .B(_4214_),
    .C(_2926_),
    .Y(_2927_));
 sg13g2_xnor2_1 _7788_ (.Y(_2928_),
    .A(_2924_),
    .B(_2927_));
 sg13g2_nor2_1 _7789_ (.A(net45),
    .B(net187),
    .Y(_2929_));
 sg13g2_a21oi_1 _7790_ (.A1(net26),
    .A2(_2928_),
    .Y(_2930_),
    .B1(_2929_));
 sg13g2_nor2_1 _7791_ (.A(net71),
    .B(_2930_),
    .Y(_2931_));
 sg13g2_nor2_1 _7792_ (.A(_1678_),
    .B(_2642_),
    .Y(_2932_));
 sg13g2_buf_1 _7793_ (.A(_2932_),
    .X(_2933_));
 sg13g2_buf_1 _7794_ (.A(_2933_),
    .X(_2934_));
 sg13g2_nor2_1 _7795_ (.A(_0548_),
    .B(net25),
    .Y(_2935_));
 sg13g2_a221oi_1 _7796_ (.B2(net18),
    .C1(net72),
    .B1(_2935_),
    .A1(net328),
    .Y(_2936_),
    .A2(net25));
 sg13g2_nor3_1 _7797_ (.A(net118),
    .B(_2931_),
    .C(_2936_),
    .Y(_0113_));
 sg13g2_xnor2_1 _7798_ (.Y(_2937_),
    .A(net187),
    .B(net183));
 sg13g2_a21oi_1 _7799_ (.A1(_1272_),
    .A2(_2901_),
    .Y(_2938_),
    .B1(_0563_));
 sg13g2_xnor2_1 _7800_ (.Y(_2939_),
    .A(_2937_),
    .B(_2938_));
 sg13g2_nand2_1 _7801_ (.Y(_2940_),
    .A(net50),
    .B(_2939_));
 sg13g2_o21ai_1 _7802_ (.B1(_2940_),
    .Y(_2941_),
    .A1(net40),
    .A2(net188));
 sg13g2_nor2_1 _7803_ (.A(_0564_),
    .B(_2933_),
    .Y(_2942_));
 sg13g2_a221oi_1 _7804_ (.B2(net19),
    .C1(net104),
    .B1(_2942_),
    .A1(net274),
    .Y(_2943_),
    .A2(net25));
 sg13g2_a21oi_1 _7805_ (.A1(net79),
    .A2(_2941_),
    .Y(_2944_),
    .B1(_2943_));
 sg13g2_and2_1 _7806_ (.A(net201),
    .B(_2944_),
    .X(_0114_));
 sg13g2_mux2_1 _7807_ (.A0(net327),
    .A1(net256),
    .S(_3988_),
    .X(_2945_));
 sg13g2_xnor2_1 _7808_ (.Y(_2946_),
    .A(net249),
    .B(net256));
 sg13g2_xnor2_1 _7809_ (.Y(_2947_),
    .A(_0297_),
    .B(_2946_));
 sg13g2_nor2_1 _7810_ (.A(_3863_),
    .B(_2947_),
    .Y(_2948_));
 sg13g2_a21oi_1 _7811_ (.A1(net68),
    .A2(net178),
    .Y(_2949_),
    .B1(_2948_));
 sg13g2_nor2_1 _7812_ (.A(net77),
    .B(_2949_),
    .Y(_2950_));
 sg13g2_a21oi_1 _7813_ (.A1(net59),
    .A2(_2945_),
    .Y(_2951_),
    .B1(_2950_));
 sg13g2_nor2_1 _7814_ (.A(net90),
    .B(_2951_),
    .Y(_0115_));
 sg13g2_xnor2_1 _7815_ (.Y(_2952_),
    .A(net187),
    .B(net188));
 sg13g2_a21oi_1 _7816_ (.A1(_0816_),
    .A2(_2908_),
    .Y(_2953_),
    .B1(_0824_));
 sg13g2_xnor2_1 _7817_ (.Y(_2954_),
    .A(_2952_),
    .B(_2953_));
 sg13g2_nor2_1 _7818_ (.A(net45),
    .B(net191),
    .Y(_2955_));
 sg13g2_a21oi_1 _7819_ (.A1(net26),
    .A2(_2954_),
    .Y(_2956_),
    .B1(_2955_));
 sg13g2_nor2_1 _7820_ (.A(net71),
    .B(_2956_),
    .Y(_2957_));
 sg13g2_nor2b_1 _7821_ (.A(net25),
    .B_N(net188),
    .Y(_2958_));
 sg13g2_a221oi_1 _7822_ (.B2(net18),
    .C1(net72),
    .B1(_2958_),
    .A1(net262),
    .Y(_2959_),
    .A2(_2934_));
 sg13g2_nor3_1 _7823_ (.A(net118),
    .B(_2957_),
    .C(_2959_),
    .Y(_0116_));
 sg13g2_inv_1 _7824_ (.Y(_2960_),
    .A(_2915_));
 sg13g2_a21o_1 _7825_ (.A2(_2960_),
    .A1(_1065_),
    .B1(_1133_),
    .X(_2961_));
 sg13g2_xor2_1 _7826_ (.B(net188),
    .A(net191),
    .X(_2962_));
 sg13g2_xnor2_1 _7827_ (.Y(_2963_),
    .A(_2961_),
    .B(_2962_));
 sg13g2_nor2_1 _7828_ (.A(net45),
    .B(net190),
    .Y(_2964_));
 sg13g2_a21oi_1 _7829_ (.A1(net26),
    .A2(_2963_),
    .Y(_2965_),
    .B1(_2964_));
 sg13g2_nor2_1 _7830_ (.A(_2923_),
    .B(_2965_),
    .Y(_2966_));
 sg13g2_nor2_1 _7831_ (.A(_2646_),
    .B(_2933_),
    .Y(_2967_));
 sg13g2_a221oi_1 _7832_ (.B2(net191),
    .C1(net72),
    .B1(_2967_),
    .A1(net323),
    .Y(_2968_),
    .A2(_2934_));
 sg13g2_nor3_1 _7833_ (.A(_2922_),
    .B(_2966_),
    .C(_2968_),
    .Y(_0117_));
 sg13g2_xnor2_1 _7834_ (.Y(_2969_),
    .A(net191),
    .B(net190));
 sg13g2_xnor2_1 _7835_ (.Y(_2970_),
    .A(_1476_),
    .B(_2969_));
 sg13g2_nor2_1 _7836_ (.A(net45),
    .B(net254),
    .Y(_2971_));
 sg13g2_a21oi_1 _7837_ (.A1(net26),
    .A2(_2970_),
    .Y(_2972_),
    .B1(_2971_));
 sg13g2_nor2_1 _7838_ (.A(_2923_),
    .B(_2972_),
    .Y(_2973_));
 sg13g2_a221oi_1 _7839_ (.B2(net190),
    .C1(net72),
    .B1(_2967_),
    .A1(net327),
    .Y(_2974_),
    .A2(net25));
 sg13g2_nor3_1 _7840_ (.A(net118),
    .B(_2973_),
    .C(_2974_),
    .Y(_0118_));
 sg13g2_xnor2_1 _7841_ (.Y(_2975_),
    .A(net254),
    .B(net190));
 sg13g2_a21oi_1 _7842_ (.A1(_0551_),
    .A2(_2901_),
    .Y(_2976_),
    .B1(_0568_));
 sg13g2_xnor2_1 _7843_ (.Y(_2977_),
    .A(_2975_),
    .B(_2976_));
 sg13g2_nand2_1 _7844_ (.Y(_2978_),
    .A(net50),
    .B(_2977_));
 sg13g2_o21ai_1 _7845_ (.B1(_2978_),
    .Y(_2979_),
    .A1(net40),
    .A2(net189));
 sg13g2_nor2_1 _7846_ (.A(_0582_),
    .B(_2933_),
    .Y(_2980_));
 sg13g2_a221oi_1 _7847_ (.B2(net19),
    .C1(net104),
    .B1(_2980_),
    .A1(net326),
    .Y(_2981_),
    .A2(net25));
 sg13g2_a21oi_1 _7848_ (.A1(net79),
    .A2(_2979_),
    .Y(_2982_),
    .B1(_2981_));
 sg13g2_and2_1 _7849_ (.A(net201),
    .B(_2982_),
    .X(_0119_));
 sg13g2_xnor2_1 _7850_ (.Y(_2983_),
    .A(net254),
    .B(net189));
 sg13g2_xnor2_1 _7851_ (.Y(_2984_),
    .A(_1569_),
    .B(_2983_));
 sg13g2_nor2_1 _7852_ (.A(net45),
    .B(net253),
    .Y(_2985_));
 sg13g2_a21oi_1 _7853_ (.A1(net26),
    .A2(_2984_),
    .Y(_2986_),
    .B1(_2985_));
 sg13g2_nor2_1 _7854_ (.A(net71),
    .B(_2986_),
    .Y(_2987_));
 sg13g2_buf_1 _7855_ (.A(net95),
    .X(_2988_));
 sg13g2_a221oi_1 _7856_ (.B2(net189),
    .C1(net70),
    .B1(_2967_),
    .A1(net264),
    .Y(_2989_),
    .A2(net25));
 sg13g2_nor3_1 _7857_ (.A(_2922_),
    .B(_2987_),
    .C(_2989_),
    .Y(_0120_));
 sg13g2_xnor2_1 _7858_ (.Y(_2990_),
    .A(net253),
    .B(_4170_));
 sg13g2_a21oi_1 _7859_ (.A1(_1145_),
    .A2(_2960_),
    .Y(_2991_),
    .B1(_1137_));
 sg13g2_xnor2_1 _7860_ (.Y(_2992_),
    .A(_2990_),
    .B(_2991_));
 sg13g2_nand2_1 _7861_ (.Y(_2993_),
    .A(net50),
    .B(_2992_));
 sg13g2_o21ai_1 _7862_ (.B1(_2993_),
    .Y(_2994_),
    .A1(_4046_),
    .A2(net162));
 sg13g2_nor2_1 _7863_ (.A(_0223_),
    .B(_2933_),
    .Y(_2995_));
 sg13g2_a221oi_1 _7864_ (.B2(net19),
    .C1(net104),
    .B1(_2995_),
    .A1(net324),
    .Y(_2996_),
    .A2(net25));
 sg13g2_a21oi_1 _7865_ (.A1(net79),
    .A2(_2994_),
    .Y(_2997_),
    .B1(_2996_));
 sg13g2_and2_1 _7866_ (.A(net201),
    .B(_2997_),
    .X(_0121_));
 sg13g2_and2_1 _7867_ (.A(_4180_),
    .B(_0228_),
    .X(_2998_));
 sg13g2_and2_1 _7868_ (.A(_0229_),
    .B(_0324_),
    .X(_2999_));
 sg13g2_nor2_1 _7869_ (.A(_2998_),
    .B(_2999_),
    .Y(_3000_));
 sg13g2_xor2_1 _7870_ (.B(_0530_),
    .A(net253),
    .X(_3001_));
 sg13g2_xnor2_1 _7871_ (.Y(_3002_),
    .A(_3000_),
    .B(_3001_));
 sg13g2_nor2_1 _7872_ (.A(net68),
    .B(_3002_),
    .Y(_3003_));
 sg13g2_a21oi_1 _7873_ (.A1(net68),
    .A2(net195),
    .Y(_3004_),
    .B1(_3003_));
 sg13g2_nand2_1 _7874_ (.Y(_3005_),
    .A(net82),
    .B(_3004_));
 sg13g2_buf_1 _7875_ (.A(net109),
    .X(_3006_));
 sg13g2_nor2_1 _7876_ (.A(_1865_),
    .B(_2642_),
    .Y(_3007_));
 sg13g2_buf_1 _7877_ (.A(_3007_),
    .X(_3008_));
 sg13g2_nand2_1 _7878_ (.Y(_3009_),
    .A(_1234_),
    .B(_3008_));
 sg13g2_o21ai_1 _7879_ (.B1(net162),
    .Y(_3010_),
    .A1(_1865_),
    .A2(_2642_));
 sg13g2_nand3_1 _7880_ (.B(_3009_),
    .C(_3010_),
    .A(net69),
    .Y(_3011_));
 sg13g2_and3_1 _7881_ (.X(_0122_),
    .A(net270),
    .B(_3005_),
    .C(_3011_));
 sg13g2_xnor2_1 _7882_ (.Y(_3012_),
    .A(_4120_),
    .B(net162));
 sg13g2_xnor2_1 _7883_ (.Y(_3013_),
    .A(_1278_),
    .B(_3012_));
 sg13g2_buf_1 _7884_ (.A(net67),
    .X(_3014_));
 sg13g2_nor2_1 _7885_ (.A(net43),
    .B(net163),
    .Y(_3015_));
 sg13g2_a21oi_1 _7886_ (.A1(net26),
    .A2(_3013_),
    .Y(_3016_),
    .B1(_3015_));
 sg13g2_nor2_1 _7887_ (.A(net71),
    .B(_3016_),
    .Y(_3017_));
 sg13g2_nor2_2 _7888_ (.A(_2646_),
    .B(net44),
    .Y(_3018_));
 sg13g2_a221oi_1 _7889_ (.B2(net195),
    .C1(net70),
    .B1(_3018_),
    .A1(_1324_),
    .Y(_3019_),
    .A2(net44));
 sg13g2_nor3_1 _7890_ (.A(net118),
    .B(_3017_),
    .C(_3019_),
    .Y(_0123_));
 sg13g2_xnor2_1 _7891_ (.Y(_3020_),
    .A(_4120_),
    .B(net163));
 sg13g2_nand2_1 _7892_ (.Y(_3021_),
    .A(_0844_),
    .B(_0846_));
 sg13g2_a21oi_1 _7893_ (.A1(_0831_),
    .A2(_0833_),
    .Y(_3022_),
    .B1(_1569_));
 sg13g2_nor2_1 _7894_ (.A(_3021_),
    .B(_3022_),
    .Y(_3023_));
 sg13g2_xnor2_1 _7895_ (.Y(_3024_),
    .A(_3020_),
    .B(_3023_));
 sg13g2_nor2_1 _7896_ (.A(net84),
    .B(_3024_),
    .Y(_3025_));
 sg13g2_a21oi_1 _7897_ (.A1(net68),
    .A2(net194),
    .Y(_3026_),
    .B1(_3025_));
 sg13g2_nor2_1 _7898_ (.A(_1058_),
    .B(net44),
    .Y(_3027_));
 sg13g2_a221oi_1 _7899_ (.B2(net19),
    .C1(net104),
    .B1(_3027_),
    .A1(_1348_),
    .Y(_3028_),
    .A2(net44));
 sg13g2_a21oi_1 _7900_ (.A1(net79),
    .A2(_3026_),
    .Y(_3029_),
    .B1(_3028_));
 sg13g2_and2_1 _7901_ (.A(net201),
    .B(_3029_),
    .X(_0124_));
 sg13g2_xnor2_1 _7902_ (.Y(_3030_),
    .A(net194),
    .B(net163));
 sg13g2_xnor2_1 _7903_ (.Y(_3031_),
    .A(_2155_),
    .B(_3030_));
 sg13g2_nor2_1 _7904_ (.A(net43),
    .B(net174),
    .Y(_3032_));
 sg13g2_a21oi_1 _7905_ (.A1(net26),
    .A2(_3031_),
    .Y(_3033_),
    .B1(_3032_));
 sg13g2_nor2_1 _7906_ (.A(net71),
    .B(_3033_),
    .Y(_3034_));
 sg13g2_a221oi_1 _7907_ (.B2(net194),
    .C1(net70),
    .B1(_3018_),
    .A1(_1422_),
    .Y(_3035_),
    .A2(net44));
 sg13g2_nor3_1 _7908_ (.A(net118),
    .B(_3034_),
    .C(_3035_),
    .Y(_0125_));
 sg13g2_mux2_1 _7909_ (.A0(net326),
    .A1(net178),
    .S(_3988_),
    .X(_3036_));
 sg13g2_inv_1 _7910_ (.Y(_3037_),
    .A(net237));
 sg13g2_nand2_1 _7911_ (.Y(_3038_),
    .A(_0469_),
    .B(_0470_));
 sg13g2_xor2_1 _7912_ (.B(net256),
    .A(net178),
    .X(_3039_));
 sg13g2_xnor2_1 _7913_ (.Y(_3040_),
    .A(_3038_),
    .B(_3039_));
 sg13g2_mux2_1 _7914_ (.A0(_3037_),
    .A1(_3040_),
    .S(net52),
    .X(_3041_));
 sg13g2_nor2_1 _7915_ (.A(net77),
    .B(_3041_),
    .Y(_3042_));
 sg13g2_a21oi_1 _7916_ (.A1(_2363_),
    .A2(_3036_),
    .Y(_3043_),
    .B1(_3042_));
 sg13g2_nor2_1 _7917_ (.A(net90),
    .B(_3043_),
    .Y(_0126_));
 sg13g2_a21oi_1 _7918_ (.A1(_1464_),
    .A2(_1473_),
    .Y(_3044_),
    .B1(_1475_));
 sg13g2_a21oi_1 _7919_ (.A1(_1477_),
    .A2(_3044_),
    .Y(_3045_),
    .B1(_1453_));
 sg13g2_xor2_1 _7920_ (.B(net174),
    .A(_4127_),
    .X(_3046_));
 sg13g2_xnor2_1 _7921_ (.Y(_3047_),
    .A(_3045_),
    .B(_3046_));
 sg13g2_nor2_1 _7922_ (.A(_4037_),
    .B(_0827_),
    .Y(_3048_));
 sg13g2_a21oi_1 _7923_ (.A1(net42),
    .A2(_3047_),
    .Y(_3049_),
    .B1(_3048_));
 sg13g2_nor2_1 _7924_ (.A(_4117_),
    .B(_3007_),
    .Y(_3050_));
 sg13g2_a221oi_1 _7925_ (.B2(net19),
    .C1(net104),
    .B1(_3050_),
    .A1(net327),
    .Y(_3051_),
    .A2(_3008_));
 sg13g2_a21oi_1 _7926_ (.A1(net79),
    .A2(_3049_),
    .Y(_3052_),
    .B1(_3051_));
 sg13g2_and2_1 _7927_ (.A(net270),
    .B(_3052_),
    .X(_0127_));
 sg13g2_buf_1 _7928_ (.A(net52),
    .X(_3053_));
 sg13g2_xor2_1 _7929_ (.B(net174),
    .A(net213),
    .X(_3054_));
 sg13g2_xnor2_1 _7930_ (.Y(_3055_),
    .A(_0593_),
    .B(_3054_));
 sg13g2_nor2_1 _7931_ (.A(net43),
    .B(net101),
    .Y(_3056_));
 sg13g2_a21oi_1 _7932_ (.A1(net24),
    .A2(_3055_),
    .Y(_3057_),
    .B1(_3056_));
 sg13g2_nor2_1 _7933_ (.A(net71),
    .B(_3057_),
    .Y(_3058_));
 sg13g2_a221oi_1 _7934_ (.B2(net213),
    .C1(net70),
    .B1(_3018_),
    .A1(net326),
    .Y(_3059_),
    .A2(net44));
 sg13g2_nor3_1 _7935_ (.A(net118),
    .B(_3058_),
    .C(_3059_),
    .Y(_0128_));
 sg13g2_xor2_1 _7936_ (.B(net101),
    .A(net213),
    .X(_3060_));
 sg13g2_xnor2_1 _7937_ (.Y(_3061_),
    .A(_1571_),
    .B(_3060_));
 sg13g2_nor2_1 _7938_ (.A(net43),
    .B(net116),
    .Y(_3062_));
 sg13g2_a21oi_1 _7939_ (.A1(net24),
    .A2(_3061_),
    .Y(_3063_),
    .B1(_3062_));
 sg13g2_nor2_1 _7940_ (.A(net71),
    .B(_3063_),
    .Y(_3064_));
 sg13g2_a221oi_1 _7941_ (.B2(net101),
    .C1(net70),
    .B1(_3018_),
    .A1(net325),
    .Y(_3065_),
    .A2(net44));
 sg13g2_nor3_1 _7942_ (.A(net118),
    .B(_3064_),
    .C(_3065_),
    .Y(_0129_));
 sg13g2_o21ai_1 _7943_ (.B1(_2572_),
    .Y(_3066_),
    .A1(_1071_),
    .A2(_2915_));
 sg13g2_xor2_1 _7944_ (.B(net101),
    .A(net116),
    .X(_3067_));
 sg13g2_xnor2_1 _7945_ (.Y(_3068_),
    .A(_3066_),
    .B(_3067_));
 sg13g2_nor2_1 _7946_ (.A(net43),
    .B(net166),
    .Y(_3069_));
 sg13g2_a21oi_1 _7947_ (.A1(net24),
    .A2(_3068_),
    .Y(_3070_),
    .B1(_3069_));
 sg13g2_nor2_1 _7948_ (.A(net71),
    .B(_3070_),
    .Y(_3071_));
 sg13g2_a221oi_1 _7949_ (.B2(net116),
    .C1(net70),
    .B1(_3018_),
    .A1(net324),
    .Y(_3072_),
    .A2(net44));
 sg13g2_nor3_1 _7950_ (.A(net118),
    .B(_3071_),
    .C(_3072_),
    .Y(_0130_));
 sg13g2_buf_1 _7951_ (.A(_3963_),
    .X(_3073_));
 sg13g2_or3_1 _7952_ (.A(_2998_),
    .B(_2999_),
    .C(_0336_),
    .X(_3074_));
 sg13g2_and2_1 _7953_ (.A(_4130_),
    .B(_3074_),
    .X(_3075_));
 sg13g2_xnor2_1 _7954_ (.Y(_3076_),
    .A(_3734_),
    .B(_0426_));
 sg13g2_xnor2_1 _7955_ (.Y(_3077_),
    .A(_3075_),
    .B(_3076_));
 sg13g2_nor2_1 _7956_ (.A(_3014_),
    .B(net230),
    .Y(_3078_));
 sg13g2_a21oi_1 _7957_ (.A1(net24),
    .A2(_3077_),
    .Y(_3079_),
    .B1(_3078_));
 sg13g2_nor2_1 _7958_ (.A(net69),
    .B(_3079_),
    .Y(_3080_));
 sg13g2_nor2_1 _7959_ (.A(_2042_),
    .B(_2642_),
    .Y(_3081_));
 sg13g2_buf_1 _7960_ (.A(_3081_),
    .X(_3082_));
 sg13g2_nor2_2 _7961_ (.A(_2646_),
    .B(_3081_),
    .Y(_3083_));
 sg13g2_a221oi_1 _7962_ (.B2(net166),
    .C1(net70),
    .B1(_3083_),
    .A1(net328),
    .Y(_3084_),
    .A2(net23));
 sg13g2_nor3_1 _7963_ (.A(net117),
    .B(_3080_),
    .C(_3084_),
    .Y(_0131_));
 sg13g2_nand2_1 _7964_ (.Y(_3085_),
    .A(_0586_),
    .B(_1279_));
 sg13g2_nor2_1 _7965_ (.A(_1278_),
    .B(_3085_),
    .Y(_3086_));
 sg13g2_or2_1 _7966_ (.X(_3087_),
    .B(_3086_),
    .A(_1299_));
 sg13g2_xnor2_1 _7967_ (.Y(_3088_),
    .A(net230),
    .B(net166));
 sg13g2_xnor2_1 _7968_ (.Y(_3089_),
    .A(_3087_),
    .B(_3088_));
 sg13g2_nand2_1 _7969_ (.Y(_3090_),
    .A(net36),
    .B(_3089_));
 sg13g2_o21ai_1 _7970_ (.B1(_3090_),
    .Y(_3091_),
    .A1(net42),
    .A2(_4148_));
 sg13g2_nor2_1 _7971_ (.A(net69),
    .B(_3091_),
    .Y(_3092_));
 sg13g2_a221oi_1 _7972_ (.B2(_3865_),
    .C1(net70),
    .B1(_3083_),
    .A1(_3974_),
    .Y(_3093_),
    .A2(net23));
 sg13g2_nor3_1 _7973_ (.A(net117),
    .B(_3092_),
    .C(_3093_),
    .Y(_0132_));
 sg13g2_a221oi_1 _7974_ (.B2(net114),
    .C1(net75),
    .B1(_3083_),
    .A1(net262),
    .Y(_3094_),
    .A2(net23));
 sg13g2_nand2_1 _7975_ (.Y(_3095_),
    .A(_0889_),
    .B(_0880_));
 sg13g2_a21oi_1 _7976_ (.A1(_0813_),
    .A2(_0854_),
    .Y(_3096_),
    .B1(_0890_));
 sg13g2_o21ai_1 _7977_ (.B1(_3096_),
    .Y(_3097_),
    .A1(_3095_),
    .A2(_2874_));
 sg13g2_xor2_1 _7978_ (.B(net114),
    .A(net230),
    .X(_3098_));
 sg13g2_xnor2_1 _7979_ (.Y(_3099_),
    .A(_3097_),
    .B(_3098_));
 sg13g2_nor2_1 _7980_ (.A(_1228_),
    .B(net238),
    .Y(_3100_));
 sg13g2_a21oi_1 _7981_ (.A1(net41),
    .A2(_3099_),
    .Y(_3101_),
    .B1(_3100_));
 sg13g2_nor2_1 _7982_ (.A(net60),
    .B(_3101_),
    .Y(_3102_));
 sg13g2_nor3_1 _7983_ (.A(_3073_),
    .B(_3094_),
    .C(_3102_),
    .Y(_0133_));
 sg13g2_nand2_1 _7984_ (.Y(_3103_),
    .A(net323),
    .B(net23));
 sg13g2_o21ai_1 _7985_ (.B1(_3103_),
    .Y(_3104_),
    .A1(_4142_),
    .A2(_3082_));
 sg13g2_nor2_1 _7986_ (.A(net82),
    .B(_3104_),
    .Y(_3105_));
 sg13g2_xor2_1 _7987_ (.B(_3783_),
    .A(net238),
    .X(_3106_));
 sg13g2_xnor2_1 _7988_ (.Y(_3107_),
    .A(_2156_),
    .B(_3106_));
 sg13g2_nor2_1 _7989_ (.A(net36),
    .B(net147),
    .Y(_3108_));
 sg13g2_a21oi_1 _7990_ (.A1(_4038_),
    .A2(_3107_),
    .Y(_3109_),
    .B1(_3108_));
 sg13g2_nor2_1 _7991_ (.A(net65),
    .B(_3109_),
    .Y(_3110_));
 sg13g2_nor3_1 _7992_ (.A(net117),
    .B(_3105_),
    .C(_3110_),
    .Y(_0134_));
 sg13g2_nor2_1 _7993_ (.A(_1474_),
    .B(_2178_),
    .Y(_3111_));
 sg13g2_nand2_1 _7994_ (.Y(_3112_),
    .A(_2183_),
    .B(_3111_));
 sg13g2_nand2_1 _7995_ (.Y(_3113_),
    .A(_2187_),
    .B(_3112_));
 sg13g2_xor2_1 _7996_ (.B(_0950_),
    .A(_3798_),
    .X(_3114_));
 sg13g2_xnor2_1 _7997_ (.Y(_3115_),
    .A(_3113_),
    .B(_3114_));
 sg13g2_nand2_1 _7998_ (.Y(_3116_),
    .A(_4047_),
    .B(_3115_));
 sg13g2_o21ai_1 _7999_ (.B1(_3116_),
    .Y(_3117_),
    .A1(net40),
    .A2(_3867_));
 sg13g2_a221oi_1 _8000_ (.B2(_0950_),
    .C1(_4026_),
    .B1(_3083_),
    .A1(net327),
    .Y(_3118_),
    .A2(net23));
 sg13g2_a21oi_1 _8001_ (.A1(net75),
    .A2(_3117_),
    .Y(_3119_),
    .B1(_3118_));
 sg13g2_and2_1 _8002_ (.A(net270),
    .B(_3119_),
    .X(_0135_));
 sg13g2_xnor2_1 _8003_ (.Y(_3120_),
    .A(net229),
    .B(net147));
 sg13g2_xnor2_1 _8004_ (.Y(_3121_),
    .A(_0603_),
    .B(_3120_));
 sg13g2_nor2_1 _8005_ (.A(_3863_),
    .B(_3121_),
    .Y(_3122_));
 sg13g2_a21oi_1 _8006_ (.A1(net68),
    .A2(net148),
    .Y(_3123_),
    .B1(_3122_));
 sg13g2_a221oi_1 _8007_ (.B2(net229),
    .C1(_4026_),
    .B1(_3083_),
    .A1(net326),
    .Y(_3124_),
    .A2(_3082_));
 sg13g2_a21oi_1 _8008_ (.A1(net75),
    .A2(_3123_),
    .Y(_3125_),
    .B1(_3124_));
 sg13g2_and2_1 _8009_ (.A(_4042_),
    .B(_3125_),
    .X(_0136_));
 sg13g2_mux2_1 _8010_ (.A0(net325),
    .A1(net237),
    .S(_3988_),
    .X(_3126_));
 sg13g2_xnor2_1 _8011_ (.Y(_3127_),
    .A(_0292_),
    .B(net237));
 sg13g2_xnor2_1 _8012_ (.Y(_3128_),
    .A(_0753_),
    .B(_3127_));
 sg13g2_nor2_1 _8013_ (.A(net52),
    .B(_0281_),
    .Y(_3129_));
 sg13g2_a21oi_1 _8014_ (.A1(_1687_),
    .A2(_3128_),
    .Y(_3130_),
    .B1(_3129_));
 sg13g2_nor2_1 _8015_ (.A(_0404_),
    .B(_3130_),
    .Y(_3131_));
 sg13g2_a21oi_1 _8016_ (.A1(_2363_),
    .A2(_3126_),
    .Y(_3132_),
    .B1(_3131_));
 sg13g2_nor2_1 _8017_ (.A(_2465_),
    .B(_3132_),
    .Y(_0137_));
 sg13g2_xnor2_1 _8018_ (.Y(_3133_),
    .A(net229),
    .B(_0894_));
 sg13g2_xnor2_1 _8019_ (.Y(_3134_),
    .A(_1578_),
    .B(_3133_));
 sg13g2_nand2_1 _8020_ (.Y(_3135_),
    .A(_1228_),
    .B(_3134_));
 sg13g2_o21ai_1 _8021_ (.B1(_3135_),
    .Y(_3136_),
    .A1(_4034_),
    .A2(_4112_));
 sg13g2_nor2_1 _8022_ (.A(net69),
    .B(_3136_),
    .Y(_3137_));
 sg13g2_a221oi_1 _8023_ (.B2(net148),
    .C1(_2988_),
    .B1(_3083_),
    .A1(_0707_),
    .Y(_3138_),
    .A2(net23));
 sg13g2_nor3_1 _8024_ (.A(net117),
    .B(_3137_),
    .C(_3138_),
    .Y(_0138_));
 sg13g2_xnor2_1 _8025_ (.Y(_3139_),
    .A(_3785_),
    .B(_0894_));
 sg13g2_xnor2_1 _8026_ (.Y(_3140_),
    .A(_1627_),
    .B(_3139_));
 sg13g2_nor2_1 _8027_ (.A(net43),
    .B(_0627_),
    .Y(_3141_));
 sg13g2_a21oi_1 _8028_ (.A1(net24),
    .A2(_3140_),
    .Y(_3142_),
    .B1(_3141_));
 sg13g2_nor2_1 _8029_ (.A(_3006_),
    .B(_3142_),
    .Y(_3143_));
 sg13g2_nor2_1 _8030_ (.A(_4112_),
    .B(net23),
    .Y(_3144_));
 sg13g2_a221oi_1 _8031_ (.B2(net18),
    .C1(_2988_),
    .B1(_3144_),
    .A1(net324),
    .Y(_3145_),
    .A2(net23));
 sg13g2_nor3_1 _8032_ (.A(net117),
    .B(_3143_),
    .C(_3145_),
    .Y(_0139_));
 sg13g2_nand3_1 _8033_ (.B(_3982_),
    .C(net66),
    .A(net273),
    .Y(_3146_));
 sg13g2_buf_2 _8034_ (.A(_3146_),
    .X(_3147_));
 sg13g2_nand3_1 _8035_ (.B(_0395_),
    .C(_3147_),
    .A(net96),
    .Y(_3148_));
 sg13g2_o21ai_1 _8036_ (.B1(_3148_),
    .Y(_3149_),
    .A1(_2046_),
    .A2(_3147_));
 sg13g2_nor2_1 _8037_ (.A(net76),
    .B(_3149_),
    .Y(_3150_));
 sg13g2_xor2_1 _8038_ (.B(_0627_),
    .A(net244),
    .X(_3151_));
 sg13g2_o21ai_1 _8039_ (.B1(_4160_),
    .Y(_3152_),
    .A1(_4147_),
    .A2(_3075_));
 sg13g2_xnor2_1 _8040_ (.Y(_3153_),
    .A(_3151_),
    .B(_3152_));
 sg13g2_nor2_1 _8041_ (.A(net36),
    .B(_0615_),
    .Y(_3154_));
 sg13g2_a21oi_1 _8042_ (.A1(_1199_),
    .A2(_3153_),
    .Y(_3155_),
    .B1(_3154_));
 sg13g2_nor2_1 _8043_ (.A(net65),
    .B(_3155_),
    .Y(_3156_));
 sg13g2_nor3_1 _8044_ (.A(net117),
    .B(_3150_),
    .C(_3156_),
    .Y(_0140_));
 sg13g2_a21oi_1 _8045_ (.A1(_1286_),
    .A2(_3087_),
    .Y(_3157_),
    .B1(_1304_));
 sg13g2_xnor2_1 _8046_ (.Y(_3158_),
    .A(net98),
    .B(net96));
 sg13g2_xnor2_1 _8047_ (.Y(_3159_),
    .A(_3157_),
    .B(_3158_));
 sg13g2_nor2_1 _8048_ (.A(net30),
    .B(net156),
    .Y(_3160_));
 sg13g2_a21oi_1 _8049_ (.A1(net39),
    .A2(_3159_),
    .Y(_3162_),
    .B1(_3160_));
 sg13g2_nand2_1 _8050_ (.Y(_3163_),
    .A(_3973_),
    .B(net83));
 sg13g2_nor2_1 _8051_ (.A(_3163_),
    .B(_3147_),
    .Y(_3164_));
 sg13g2_a21oi_1 _8052_ (.A1(net98),
    .A2(_3147_),
    .Y(_3165_),
    .B1(_3164_));
 sg13g2_nor2_1 _8053_ (.A(net75),
    .B(_3165_),
    .Y(_3166_));
 sg13g2_a21oi_1 _8054_ (.A1(net57),
    .A2(_3162_),
    .Y(_3167_),
    .B1(_3166_));
 sg13g2_nor2_1 _8055_ (.A(net90),
    .B(_3167_),
    .Y(_0141_));
 sg13g2_nand2b_1 _8056_ (.Y(_3168_),
    .B(_0893_),
    .A_N(_0902_));
 sg13g2_and2_1 _8057_ (.A(_0958_),
    .B(_3168_),
    .X(_3169_));
 sg13g2_xnor2_1 _8058_ (.Y(_3170_),
    .A(net98),
    .B(net156));
 sg13g2_xnor2_1 _8059_ (.Y(_3172_),
    .A(_3169_),
    .B(_3170_));
 sg13g2_nor2_1 _8060_ (.A(net30),
    .B(net97),
    .Y(_3173_));
 sg13g2_a21oi_1 _8061_ (.A1(net39),
    .A2(_3172_),
    .Y(_3174_),
    .B1(_3173_));
 sg13g2_nand2_1 _8062_ (.Y(_3175_),
    .A(_1346_),
    .B(net83));
 sg13g2_nor2_1 _8063_ (.A(_3175_),
    .B(_3147_),
    .Y(_3176_));
 sg13g2_a21oi_1 _8064_ (.A1(net156),
    .A2(_3147_),
    .Y(_3177_),
    .B1(_3176_));
 sg13g2_nor2_1 _8065_ (.A(net75),
    .B(_3177_),
    .Y(_3178_));
 sg13g2_a21oi_1 _8066_ (.A1(net57),
    .A2(_3174_),
    .Y(_3179_),
    .B1(_3178_));
 sg13g2_nor2_1 _8067_ (.A(net90),
    .B(_3179_),
    .Y(_0142_));
 sg13g2_xor2_1 _8068_ (.B(_0624_),
    .A(_0620_),
    .X(_3180_));
 sg13g2_xnor2_1 _8069_ (.Y(_3182_),
    .A(_1375_),
    .B(_3180_));
 sg13g2_nor2_1 _8070_ (.A(net43),
    .B(net208),
    .Y(_3183_));
 sg13g2_a21oi_1 _8071_ (.A1(_3053_),
    .A2(_3182_),
    .Y(_3184_),
    .B1(_3183_));
 sg13g2_nor2_1 _8072_ (.A(net69),
    .B(_3184_),
    .Y(_3185_));
 sg13g2_mux2_1 _8073_ (.A0(_1422_),
    .A1(_0620_),
    .S(_3147_),
    .X(_3186_));
 sg13g2_nor2_1 _8074_ (.A(net56),
    .B(_3186_),
    .Y(_3187_));
 sg13g2_nor3_1 _8075_ (.A(net117),
    .B(_3185_),
    .C(_3187_),
    .Y(_0143_));
 sg13g2_xnor2_1 _8076_ (.Y(_3188_),
    .A(net97),
    .B(_3944_));
 sg13g2_xnor2_1 _8077_ (.Y(_3189_),
    .A(_0339_),
    .B(_3188_));
 sg13g2_nor2_1 _8078_ (.A(net32),
    .B(net167),
    .Y(_3190_));
 sg13g2_a21oi_1 _8079_ (.A1(net31),
    .A2(_3189_),
    .Y(_3192_),
    .B1(_3190_));
 sg13g2_nand2_1 _8080_ (.Y(_3193_),
    .A(net61),
    .B(_3192_));
 sg13g2_nor4_2 _8081_ (.A(_3979_),
    .B(net329),
    .C(net272),
    .Y(_3194_),
    .D(_1237_));
 sg13g2_and2_1 _8082_ (.A(net109),
    .B(_3147_),
    .X(_3195_));
 sg13g2_buf_1 _8083_ (.A(_3195_),
    .X(_3196_));
 sg13g2_a22oi_1 _8084_ (.Y(_3197_),
    .B1(_3196_),
    .B2(net208),
    .A2(_3194_),
    .A1(net265));
 sg13g2_a21oi_1 _8085_ (.A1(_3193_),
    .A2(_3197_),
    .Y(_0144_),
    .B1(net91));
 sg13g2_xor2_1 _8086_ (.B(net208),
    .A(net167),
    .X(_3198_));
 sg13g2_xnor2_1 _8087_ (.Y(_3199_),
    .A(_0631_),
    .B(_3198_));
 sg13g2_nor2_1 _8088_ (.A(net32),
    .B(net207),
    .Y(_3200_));
 sg13g2_a21oi_1 _8089_ (.A1(net31),
    .A2(_3199_),
    .Y(_3202_),
    .B1(_3200_));
 sg13g2_nand2_1 _8090_ (.Y(_3203_),
    .A(net61),
    .B(_3202_));
 sg13g2_a22oi_1 _8091_ (.Y(_3204_),
    .B1(_3196_),
    .B2(net167),
    .A2(_3194_),
    .A1(net266));
 sg13g2_a21oi_1 _8092_ (.A1(_3203_),
    .A2(_3204_),
    .Y(_0145_),
    .B1(net91));
 sg13g2_xnor2_1 _8093_ (.Y(_3205_),
    .A(_0418_),
    .B(net207));
 sg13g2_xnor2_1 _8094_ (.Y(_3206_),
    .A(_1586_),
    .B(_3205_));
 sg13g2_nor2_1 _8095_ (.A(net32),
    .B(net173),
    .Y(_3207_));
 sg13g2_a21oi_1 _8096_ (.A1(net31),
    .A2(_3206_),
    .Y(_3208_),
    .B1(_3207_));
 sg13g2_nand2_1 _8097_ (.Y(_3209_),
    .A(net61),
    .B(_3208_));
 sg13g2_a22oi_1 _8098_ (.Y(_3210_),
    .B1(_3196_),
    .B2(net207),
    .A2(_3194_),
    .A1(net264));
 sg13g2_buf_1 _8099_ (.A(net204),
    .X(_3212_));
 sg13g2_a21oi_1 _8100_ (.A1(_3209_),
    .A2(_3210_),
    .Y(_0146_),
    .B1(_3212_));
 sg13g2_xor2_1 _8101_ (.B(net207),
    .A(net173),
    .X(_3213_));
 sg13g2_xnor2_1 _8102_ (.Y(_3214_),
    .A(_1629_),
    .B(_3213_));
 sg13g2_buf_1 _8103_ (.A(_0692_),
    .X(_3215_));
 sg13g2_nor2_1 _8104_ (.A(_3215_),
    .B(net155),
    .Y(_3216_));
 sg13g2_a21oi_1 _8105_ (.A1(net31),
    .A2(_3214_),
    .Y(_3217_),
    .B1(_3216_));
 sg13g2_nand2_1 _8106_ (.Y(_3218_),
    .A(net61),
    .B(_3217_));
 sg13g2_a22oi_1 _8107_ (.Y(_3219_),
    .B1(_3196_),
    .B2(net173),
    .A2(_3194_),
    .A1(net263));
 sg13g2_a21oi_1 _8108_ (.A1(_3218_),
    .A2(_3219_),
    .Y(_0147_),
    .B1(_3212_));
 sg13g2_nand2_1 _8109_ (.Y(_3221_),
    .A(_1018_),
    .B(_1019_));
 sg13g2_a21oi_1 _8110_ (.A1(_1012_),
    .A2(_1013_),
    .Y(_3222_),
    .B1(_1015_));
 sg13g2_nor2_1 _8111_ (.A(_3221_),
    .B(_3222_),
    .Y(_3223_));
 sg13g2_xnor2_1 _8112_ (.Y(_3224_),
    .A(net179),
    .B(net237));
 sg13g2_xnor2_1 _8113_ (.Y(_3225_),
    .A(_3223_),
    .B(_3224_));
 sg13g2_nor2_1 _8114_ (.A(_3014_),
    .B(net236),
    .Y(_3226_));
 sg13g2_a21oi_1 _8115_ (.A1(_3053_),
    .A2(_3225_),
    .Y(_3227_),
    .B1(_3226_));
 sg13g2_nor2_1 _8116_ (.A(net69),
    .B(_3227_),
    .Y(_3228_));
 sg13g2_mux2_1 _8117_ (.A0(net324),
    .A1(net179),
    .S(_3988_),
    .X(_3229_));
 sg13g2_nor2_1 _8118_ (.A(net56),
    .B(_3229_),
    .Y(_3230_));
 sg13g2_nor3_1 _8119_ (.A(_3073_),
    .B(_3228_),
    .C(_3230_),
    .Y(_0148_));
 sg13g2_buf_1 _8120_ (.A(net78),
    .X(_3232_));
 sg13g2_nand2_1 _8121_ (.Y(_3233_),
    .A(_4107_),
    .B(_1219_));
 sg13g2_a21oi_1 _8122_ (.A1(_4102_),
    .A2(_3233_),
    .Y(_3234_),
    .B1(_0344_));
 sg13g2_xor2_1 _8123_ (.B(_0634_),
    .A(net173),
    .X(_3235_));
 sg13g2_xnor2_1 _8124_ (.Y(_3236_),
    .A(_3234_),
    .B(_3235_));
 sg13g2_mux2_1 _8125_ (.A0(_3917_),
    .A1(_3236_),
    .S(net40),
    .X(_3237_));
 sg13g2_nand2_1 _8126_ (.Y(_3238_),
    .A(net54),
    .B(_3237_));
 sg13g2_nor2b_1 _8127_ (.A(_1237_),
    .B_N(_2643_),
    .Y(_3239_));
 sg13g2_buf_2 _8128_ (.A(_3239_),
    .X(_3240_));
 sg13g2_a21oi_1 _8129_ (.A1(net66),
    .A2(_2643_),
    .Y(_3242_),
    .B1(net100));
 sg13g2_buf_2 _8130_ (.A(_3242_),
    .X(_3243_));
 sg13g2_a22oi_1 _8131_ (.Y(_3244_),
    .B1(_3243_),
    .B2(net155),
    .A2(_3240_),
    .A1(net328));
 sg13g2_a21oi_1 _8132_ (.A1(_3238_),
    .A2(_3244_),
    .Y(_0149_),
    .B1(net87));
 sg13g2_a21oi_1 _8133_ (.A1(_1280_),
    .A2(_0631_),
    .Y(_3245_),
    .B1(_1290_));
 sg13g2_xnor2_1 _8134_ (.Y(_3246_),
    .A(net111),
    .B(net155));
 sg13g2_xnor2_1 _8135_ (.Y(_3247_),
    .A(_3245_),
    .B(_3246_));
 sg13g2_nor2_1 _8136_ (.A(net22),
    .B(net172),
    .Y(_3248_));
 sg13g2_a21oi_1 _8137_ (.A1(net31),
    .A2(_3247_),
    .Y(_3249_),
    .B1(_3248_));
 sg13g2_nand2_1 _8138_ (.Y(_3250_),
    .A(net54),
    .B(_3249_));
 sg13g2_a22oi_1 _8139_ (.Y(_3252_),
    .B1(_3243_),
    .B2(net111),
    .A2(_3240_),
    .A1(net274));
 sg13g2_a21oi_1 _8140_ (.A1(_3250_),
    .A2(_3252_),
    .Y(_0150_),
    .B1(net87));
 sg13g2_xor2_1 _8141_ (.B(net172),
    .A(net111),
    .X(_3253_));
 sg13g2_nand2_1 _8142_ (.Y(_3254_),
    .A(_0915_),
    .B(_0917_));
 sg13g2_nand2_1 _8143_ (.Y(_3255_),
    .A(_1579_),
    .B(_0893_));
 sg13g2_o21ai_1 _8144_ (.B1(_3255_),
    .Y(_3256_),
    .A1(_0911_),
    .A2(_0958_));
 sg13g2_nand2_1 _8145_ (.Y(_3257_),
    .A(_3254_),
    .B(_3256_));
 sg13g2_nand2_1 _8146_ (.Y(_3258_),
    .A(_0936_),
    .B(_3257_));
 sg13g2_xnor2_1 _8147_ (.Y(_3259_),
    .A(_3253_),
    .B(_3258_));
 sg13g2_nor2_1 _8148_ (.A(net22),
    .B(net198),
    .Y(_3260_));
 sg13g2_a21oi_1 _8149_ (.A1(net31),
    .A2(_3259_),
    .Y(_3262_),
    .B1(_3260_));
 sg13g2_nand2_1 _8150_ (.Y(_3263_),
    .A(net54),
    .B(_3262_));
 sg13g2_a22oi_1 _8151_ (.Y(_3264_),
    .B1(_3243_),
    .B2(net172),
    .A2(_3240_),
    .A1(net262));
 sg13g2_a21oi_1 _8152_ (.A1(_3263_),
    .A2(_3264_),
    .Y(_0151_),
    .B1(net87));
 sg13g2_nand2b_1 _8153_ (.Y(_3265_),
    .B(_1375_),
    .A_N(_2148_));
 sg13g2_nand2_1 _8154_ (.Y(_3266_),
    .A(_1396_),
    .B(_3265_));
 sg13g2_xor2_1 _8155_ (.B(net172),
    .A(net198),
    .X(_3267_));
 sg13g2_xnor2_1 _8156_ (.Y(_3268_),
    .A(_3266_),
    .B(_3267_));
 sg13g2_nor2_1 _8157_ (.A(_3215_),
    .B(net218),
    .Y(_3269_));
 sg13g2_a21oi_1 _8158_ (.A1(net31),
    .A2(_3268_),
    .Y(_3270_),
    .B1(_3269_));
 sg13g2_nand2_1 _8159_ (.Y(_3272_),
    .A(_3232_),
    .B(_3270_));
 sg13g2_a22oi_1 _8160_ (.Y(_3273_),
    .B1(_3243_),
    .B2(net198),
    .A2(_3240_),
    .A1(net323));
 sg13g2_a21oi_1 _8161_ (.A1(_3272_),
    .A2(_3273_),
    .Y(_0152_),
    .B1(net87));
 sg13g2_xor2_1 _8162_ (.B(net218),
    .A(net198),
    .X(_3274_));
 sg13g2_xnor2_1 _8163_ (.Y(_3275_),
    .A(_0352_),
    .B(_3274_));
 sg13g2_nor2_1 _8164_ (.A(net22),
    .B(net171),
    .Y(_3276_));
 sg13g2_a21oi_1 _8165_ (.A1(net31),
    .A2(_3275_),
    .Y(_3277_),
    .B1(_3276_));
 sg13g2_nand2_1 _8166_ (.Y(_3278_),
    .A(_3232_),
    .B(_3277_));
 sg13g2_a22oi_1 _8167_ (.Y(_3279_),
    .B1(_3243_),
    .B2(net218),
    .A2(_3240_),
    .A1(net265));
 sg13g2_a21oi_1 _8168_ (.A1(_3278_),
    .A2(_3279_),
    .Y(_0153_),
    .B1(net87));
 sg13g2_buf_1 _8169_ (.A(net51),
    .X(_3281_));
 sg13g2_nor2_1 _8170_ (.A(_4077_),
    .B(_0660_),
    .Y(_3282_));
 sg13g2_xnor2_1 _8171_ (.Y(_3283_),
    .A(_0643_),
    .B(_3282_));
 sg13g2_nor2_1 _8172_ (.A(net22),
    .B(net153),
    .Y(_3284_));
 sg13g2_a21oi_1 _8173_ (.A1(net21),
    .A2(_3283_),
    .Y(_3285_),
    .B1(_3284_));
 sg13g2_nand2_1 _8174_ (.Y(_3286_),
    .A(net54),
    .B(_3285_));
 sg13g2_a22oi_1 _8175_ (.Y(_3287_),
    .B1(_3243_),
    .B2(net171),
    .A2(_3240_),
    .A1(net266));
 sg13g2_a21oi_1 _8176_ (.A1(_3286_),
    .A2(_3287_),
    .Y(_0154_),
    .B1(net87));
 sg13g2_nor2_1 _8177_ (.A(_1598_),
    .B(_1587_),
    .Y(_3288_));
 sg13g2_xnor2_1 _8178_ (.Y(_3289_),
    .A(net171),
    .B(net153));
 sg13g2_xnor2_1 _8179_ (.Y(_3291_),
    .A(_3288_),
    .B(_3289_));
 sg13g2_nor2_1 _8180_ (.A(net22),
    .B(net206),
    .Y(_3292_));
 sg13g2_a21oi_1 _8181_ (.A1(net21),
    .A2(_3291_),
    .Y(_3293_),
    .B1(_3292_));
 sg13g2_nand2_1 _8182_ (.Y(_3294_),
    .A(net54),
    .B(_3293_));
 sg13g2_a22oi_1 _8183_ (.Y(_3295_),
    .B1(_3243_),
    .B2(net153),
    .A2(_3240_),
    .A1(net264));
 sg13g2_a21oi_1 _8184_ (.A1(_3294_),
    .A2(_3295_),
    .Y(_0155_),
    .B1(net87));
 sg13g2_nor2_1 _8185_ (.A(_4078_),
    .B(_4081_),
    .Y(_3296_));
 sg13g2_xor2_1 _8186_ (.B(_3296_),
    .A(_1180_),
    .X(_3297_));
 sg13g2_nor2_1 _8187_ (.A(net22),
    .B(_0659_),
    .Y(_3298_));
 sg13g2_a21oi_1 _8188_ (.A1(net21),
    .A2(_3297_),
    .Y(_3299_),
    .B1(_3298_));
 sg13g2_nand2_1 _8189_ (.Y(_3301_),
    .A(net54),
    .B(_3299_));
 sg13g2_a22oi_1 _8190_ (.Y(_3302_),
    .B1(_3243_),
    .B2(net206),
    .A2(_3240_),
    .A1(net263));
 sg13g2_a21oi_1 _8191_ (.A1(_3301_),
    .A2(_3302_),
    .Y(_0156_),
    .B1(net87));
 sg13g2_nand2_1 _8192_ (.Y(_3303_),
    .A(_4083_),
    .B(_4093_));
 sg13g2_o21ai_1 _8193_ (.B1(_1204_),
    .Y(_3304_),
    .A1(_3303_),
    .A2(_3234_));
 sg13g2_xor2_1 _8194_ (.B(net154),
    .A(net206),
    .X(_3305_));
 sg13g2_xnor2_1 _8195_ (.Y(_3306_),
    .A(_3304_),
    .B(_3305_));
 sg13g2_nor2_1 _8196_ (.A(net22),
    .B(net170),
    .Y(_3307_));
 sg13g2_a21oi_1 _8197_ (.A1(net21),
    .A2(_3306_),
    .Y(_3308_),
    .B1(_3307_));
 sg13g2_nand2_1 _8198_ (.Y(_3309_),
    .A(net54),
    .B(_3308_));
 sg13g2_inv_1 _8199_ (.Y(_3311_),
    .A(_2712_));
 sg13g2_a21oi_1 _8200_ (.A1(net66),
    .A2(_3311_),
    .Y(_3312_),
    .B1(net203));
 sg13g2_buf_2 _8201_ (.A(_3312_),
    .X(_3313_));
 sg13g2_nor2_1 _8202_ (.A(_1237_),
    .B(_2712_),
    .Y(_3314_));
 sg13g2_buf_2 _8203_ (.A(_3314_),
    .X(_3315_));
 sg13g2_a22oi_1 _8204_ (.Y(_3316_),
    .B1(_3315_),
    .B2(_1234_),
    .A2(_3313_),
    .A1(net154));
 sg13g2_buf_1 _8205_ (.A(_3964_),
    .X(_3317_));
 sg13g2_a21oi_1 _8206_ (.A1(_3309_),
    .A2(_3316_),
    .Y(_0157_),
    .B1(net86));
 sg13g2_nor2_1 _8207_ (.A(_4068_),
    .B(_4073_),
    .Y(_3318_));
 sg13g2_xor2_1 _8208_ (.B(_3318_),
    .A(_1308_),
    .X(_3319_));
 sg13g2_nor2_1 _8209_ (.A(net22),
    .B(net243),
    .Y(_3321_));
 sg13g2_a21oi_1 _8210_ (.A1(net21),
    .A2(_3319_),
    .Y(_3322_),
    .B1(_3321_));
 sg13g2_nand2_1 _8211_ (.Y(_3323_),
    .A(net54),
    .B(_3322_));
 sg13g2_a22oi_1 _8212_ (.Y(_3324_),
    .B1(_3315_),
    .B2(_1324_),
    .A2(_3313_),
    .A1(net170));
 sg13g2_a21oi_1 _8213_ (.A1(_3323_),
    .A2(_3324_),
    .Y(_0158_),
    .B1(net86));
 sg13g2_a21oi_1 _8214_ (.A1(_0291_),
    .A2(_0294_),
    .Y(_3325_),
    .B1(_0297_));
 sg13g2_nor2b_1 _8215_ (.A(_3325_),
    .B_N(_0301_),
    .Y(_3326_));
 sg13g2_xnor2_1 _8216_ (.Y(_3327_),
    .A(_0284_),
    .B(_3811_));
 sg13g2_xnor2_1 _8217_ (.Y(_3328_),
    .A(_3326_),
    .B(_3327_));
 sg13g2_nor2_1 _8218_ (.A(_2470_),
    .B(net251),
    .Y(_3329_));
 sg13g2_a21oi_1 _8219_ (.A1(_0406_),
    .A2(_3328_),
    .Y(_3331_),
    .B1(_3329_));
 sg13g2_mux2_1 _8220_ (.A0(_0285_),
    .A1(_2046_),
    .S(_1551_),
    .X(_3332_));
 sg13g2_nor2_1 _8221_ (.A(net75),
    .B(_3332_),
    .Y(_3333_));
 sg13g2_a21oi_1 _8222_ (.A1(net56),
    .A2(_3331_),
    .Y(_3334_),
    .B1(_3333_));
 sg13g2_nor2_1 _8223_ (.A(_2465_),
    .B(_3334_),
    .Y(_0159_));
 sg13g2_o21ai_1 _8224_ (.B1(_0945_),
    .Y(_3335_),
    .A1(_0924_),
    .A2(_3169_));
 sg13g2_xor2_1 _8225_ (.B(net243),
    .A(net170),
    .X(_3336_));
 sg13g2_xnor2_1 _8226_ (.Y(_3337_),
    .A(_3335_),
    .B(_3336_));
 sg13g2_nor2_1 _8227_ (.A(net30),
    .B(net224),
    .Y(_3338_));
 sg13g2_a21oi_1 _8228_ (.A1(net21),
    .A2(_3337_),
    .Y(_3339_),
    .B1(_3338_));
 sg13g2_nand2_1 _8229_ (.Y(_3341_),
    .A(net57),
    .B(_3339_));
 sg13g2_a22oi_1 _8230_ (.Y(_3342_),
    .B1(_3315_),
    .B2(_1348_),
    .A2(_3313_),
    .A1(net243));
 sg13g2_a21oi_1 _8231_ (.A1(_3341_),
    .A2(_3342_),
    .Y(_0160_),
    .B1(net86));
 sg13g2_a21oi_1 _8232_ (.A1(_2147_),
    .A2(_3266_),
    .Y(_3343_),
    .B1(_2150_));
 sg13g2_xnor2_1 _8233_ (.Y(_3344_),
    .A(net224),
    .B(_3787_));
 sg13g2_xnor2_1 _8234_ (.Y(_3345_),
    .A(_3343_),
    .B(_3344_));
 sg13g2_o21ai_1 _8235_ (.B1(net102),
    .Y(_3346_),
    .A1(net51),
    .A2(net152));
 sg13g2_a21oi_1 _8236_ (.A1(net39),
    .A2(_3345_),
    .Y(_3347_),
    .B1(_3346_));
 sg13g2_a221oi_1 _8237_ (.B2(_1422_),
    .C1(_3347_),
    .B1(_3315_),
    .A1(net224),
    .Y(_3348_),
    .A2(_3313_));
 sg13g2_nor2_1 _8238_ (.A(net90),
    .B(_3348_),
    .Y(_0161_));
 sg13g2_a21oi_1 _8239_ (.A1(_4075_),
    .A2(_3304_),
    .Y(_3350_),
    .B1(_1200_));
 sg13g2_xnor2_1 _8240_ (.Y(_3351_),
    .A(net224),
    .B(net152));
 sg13g2_xnor2_1 _8241_ (.Y(_3352_),
    .A(_3350_),
    .B(_3351_));
 sg13g2_nor2_1 _8242_ (.A(net30),
    .B(net149),
    .Y(_3353_));
 sg13g2_a21oi_1 _8243_ (.A1(net21),
    .A2(_3352_),
    .Y(_3354_),
    .B1(_3353_));
 sg13g2_nand2_1 _8244_ (.Y(_3355_),
    .A(net57),
    .B(_3354_));
 sg13g2_a22oi_1 _8245_ (.Y(_3356_),
    .B1(_3315_),
    .B2(net265),
    .A2(_3313_),
    .A1(net152));
 sg13g2_a21oi_1 _8246_ (.A1(_3355_),
    .A2(_3356_),
    .Y(_0162_),
    .B1(net86));
 sg13g2_a21oi_1 _8247_ (.A1(_0667_),
    .A2(_1308_),
    .Y(_3357_),
    .B1(_0676_));
 sg13g2_xnor2_1 _8248_ (.Y(_3358_),
    .A(net149),
    .B(_0673_));
 sg13g2_xnor2_1 _8249_ (.Y(_3360_),
    .A(_3357_),
    .B(_3358_));
 sg13g2_nor2_1 _8250_ (.A(net30),
    .B(net151),
    .Y(_3361_));
 sg13g2_a21oi_1 _8251_ (.A1(_3281_),
    .A2(_3360_),
    .Y(_3362_),
    .B1(_3361_));
 sg13g2_nand2_1 _8252_ (.Y(_3363_),
    .A(net57),
    .B(_3362_));
 sg13g2_a22oi_1 _8253_ (.Y(_3364_),
    .B1(_3315_),
    .B2(net266),
    .A2(_3313_),
    .A1(net149));
 sg13g2_a21oi_1 _8254_ (.A1(_3363_),
    .A2(_3364_),
    .Y(_0163_),
    .B1(net86));
 sg13g2_nor2b_1 _8255_ (.A(_0722_),
    .B_N(_0724_),
    .Y(_3365_));
 sg13g2_nand2b_1 _8256_ (.Y(_3366_),
    .B(_3365_),
    .A_N(_2097_));
 sg13g2_xor2_1 _8257_ (.B(net151),
    .A(net149),
    .X(_3367_));
 sg13g2_xnor2_1 _8258_ (.Y(_3368_),
    .A(_3366_),
    .B(_3367_));
 sg13g2_nor2_1 _8259_ (.A(net30),
    .B(net199),
    .Y(_3370_));
 sg13g2_a21oi_1 _8260_ (.A1(net21),
    .A2(_3368_),
    .Y(_3371_),
    .B1(_3370_));
 sg13g2_nand2_1 _8261_ (.Y(_3372_),
    .A(net57),
    .B(_3371_));
 sg13g2_a22oi_1 _8262_ (.Y(_3373_),
    .B1(_3315_),
    .B2(net264),
    .A2(_3313_),
    .A1(net151));
 sg13g2_a21oi_1 _8263_ (.A1(_3372_),
    .A2(_3373_),
    .Y(_0164_),
    .B1(net86));
 sg13g2_nor2_1 _8264_ (.A(_4060_),
    .B(_4063_),
    .Y(_3374_));
 sg13g2_nor2_1 _8265_ (.A(_0976_),
    .B(_0982_),
    .Y(_3375_));
 sg13g2_nand2_1 _8266_ (.Y(_3376_),
    .A(_3375_),
    .B(_1181_));
 sg13g2_xor2_1 _8267_ (.B(_3376_),
    .A(_3374_),
    .X(_3377_));
 sg13g2_nor2_1 _8268_ (.A(net30),
    .B(net169),
    .Y(_3378_));
 sg13g2_a21oi_1 _8269_ (.A1(_3281_),
    .A2(_3377_),
    .Y(_3380_),
    .B1(_3378_));
 sg13g2_nand2_1 _8270_ (.Y(_3381_),
    .A(net57),
    .B(_3380_));
 sg13g2_a22oi_1 _8271_ (.Y(_3382_),
    .B1(_3315_),
    .B2(net263),
    .A2(_3313_),
    .A1(net199));
 sg13g2_a21oi_1 _8272_ (.A1(_3381_),
    .A2(_3382_),
    .Y(_0165_),
    .B1(net86));
 sg13g2_inv_1 _8273_ (.Y(_3383_),
    .A(_3304_));
 sg13g2_o21ai_1 _8274_ (.B1(_1202_),
    .Y(_3384_),
    .A1(_1208_),
    .A2(_3383_));
 sg13g2_xor2_1 _8275_ (.B(net169),
    .A(net199),
    .X(_3385_));
 sg13g2_xnor2_1 _8276_ (.Y(_3386_),
    .A(_3384_),
    .B(_3385_));
 sg13g2_nor2_1 _8277_ (.A(net43),
    .B(net168),
    .Y(_3387_));
 sg13g2_a21oi_1 _8278_ (.A1(net24),
    .A2(_3386_),
    .Y(_3388_),
    .B1(_3387_));
 sg13g2_nor2_1 _8279_ (.A(net69),
    .B(_3388_),
    .Y(_3390_));
 sg13g2_nand2_1 _8280_ (.Y(_3391_),
    .A(net328),
    .B(net20));
 sg13g2_o21ai_1 _8281_ (.B1(_3391_),
    .Y(_3392_),
    .A1(_0644_),
    .A2(net20));
 sg13g2_nor2_1 _8282_ (.A(net56),
    .B(_3392_),
    .Y(_3393_));
 sg13g2_nor3_1 _8283_ (.A(net117),
    .B(_3390_),
    .C(_3393_),
    .Y(_0166_));
 sg13g2_nor2_1 _8284_ (.A(_4053_),
    .B(_0657_),
    .Y(_3394_));
 sg13g2_xnor2_1 _8285_ (.Y(_3395_),
    .A(_1310_),
    .B(_3394_));
 sg13g2_nor2_1 _8286_ (.A(net30),
    .B(_3815_),
    .Y(_3396_));
 sg13g2_a21oi_1 _8287_ (.A1(net39),
    .A2(_3395_),
    .Y(_3397_),
    .B1(_3396_));
 sg13g2_nand2_1 _8288_ (.Y(_3398_),
    .A(net57),
    .B(_3397_));
 sg13g2_nand2_1 _8289_ (.Y(_3400_),
    .A(_3974_),
    .B(_0391_));
 sg13g2_o21ai_1 _8290_ (.B1(_3400_),
    .Y(_3401_),
    .A1(_0684_),
    .A2(_0392_));
 sg13g2_nand2_1 _8291_ (.Y(_3402_),
    .A(net60),
    .B(_3401_));
 sg13g2_a21oi_1 _8292_ (.A1(_3398_),
    .A2(_3402_),
    .Y(_0167_),
    .B1(net86));
 sg13g2_a21oi_1 _8293_ (.A1(_0720_),
    .A2(_3366_),
    .Y(_3403_),
    .B1(_0730_));
 sg13g2_xnor2_1 _8294_ (.Y(_3404_),
    .A(_0374_),
    .B(net235));
 sg13g2_xnor2_1 _8295_ (.Y(_3405_),
    .A(_3403_),
    .B(_3404_));
 sg13g2_nor2_1 _8296_ (.A(net50),
    .B(net242),
    .Y(_3406_));
 sg13g2_a21oi_1 _8297_ (.A1(net24),
    .A2(_3405_),
    .Y(_3407_),
    .B1(_3406_));
 sg13g2_nor2_1 _8298_ (.A(_3006_),
    .B(_3407_),
    .Y(_3408_));
 sg13g2_nand2_1 _8299_ (.Y(_3410_),
    .A(_1726_),
    .B(_0391_));
 sg13g2_o21ai_1 _8300_ (.B1(_3410_),
    .Y(_3411_),
    .A1(_0369_),
    .A2(net20));
 sg13g2_nor2_1 _8301_ (.A(net82),
    .B(_3411_),
    .Y(_3412_));
 sg13g2_nor3_1 _8302_ (.A(net204),
    .B(_3408_),
    .C(_3412_),
    .Y(_0168_));
 sg13g2_o21ai_1 _8303_ (.B1(_2152_),
    .Y(_3413_),
    .A1(_1385_),
    .A2(_3343_));
 sg13g2_or2_1 _8304_ (.X(_3414_),
    .B(_4056_),
    .A(_4052_));
 sg13g2_xnor2_1 _8305_ (.Y(_3415_),
    .A(_3413_),
    .B(_3414_));
 sg13g2_nor2_1 _8306_ (.A(_4047_),
    .B(net200),
    .Y(_3416_));
 sg13g2_a21oi_1 _8307_ (.A1(net24),
    .A2(_3415_),
    .Y(_3417_),
    .B1(_3416_));
 sg13g2_nor2_1 _8308_ (.A(net69),
    .B(_3417_),
    .Y(_3418_));
 sg13g2_mux2_1 _8309_ (.A0(_3789_),
    .A1(net323),
    .S(net20),
    .X(_3420_));
 sg13g2_nor2_1 _8310_ (.A(net82),
    .B(_3420_),
    .Y(_3421_));
 sg13g2_nor3_1 _8311_ (.A(_3966_),
    .B(_3418_),
    .C(_3421_),
    .Y(_0169_));
 sg13g2_a21oi_1 _8312_ (.A1(_0281_),
    .A2(_0477_),
    .Y(_3422_),
    .B1(_0479_));
 sg13g2_nand2_1 _8313_ (.Y(_3423_),
    .A(_0474_),
    .B(_3422_));
 sg13g2_xor2_1 _8314_ (.B(_3811_),
    .A(net251),
    .X(_3424_));
 sg13g2_xnor2_1 _8315_ (.Y(_3425_),
    .A(_3423_),
    .B(_3424_));
 sg13g2_o21ai_1 _8316_ (.B1(_4039_),
    .Y(_3426_),
    .A1(_0406_),
    .A2(_0286_));
 sg13g2_a21oi_1 _8317_ (.A1(net41),
    .A2(_3425_),
    .Y(_3427_),
    .B1(_3426_));
 sg13g2_mux2_1 _8318_ (.A0(net251),
    .A1(_1324_),
    .S(net63),
    .X(_3428_));
 sg13g2_o21ai_1 _8319_ (.B1(net270),
    .Y(_3430_),
    .A1(_4027_),
    .A2(_3428_));
 sg13g2_nor2_1 _8320_ (.A(_3427_),
    .B(_3430_),
    .Y(_0170_));
 sg13g2_nor2_1 _8321_ (.A(net102),
    .B(_3959_),
    .Y(_3431_));
 sg13g2_nor2_1 _8322_ (.A(net77),
    .B(_3201_),
    .Y(_3432_));
 sg13g2_a21oi_1 _8323_ (.A1(_3201_),
    .A2(_3431_),
    .Y(_3433_),
    .B1(_3432_));
 sg13g2_nor2_1 _8324_ (.A(_3965_),
    .B(_3433_),
    .Y(_0171_));
 sg13g2_and3_1 _8325_ (.X(_3434_),
    .A(_3161_),
    .B(_3300_),
    .C(_3251_));
 sg13g2_buf_1 _8326_ (.A(_3434_),
    .X(_3435_));
 sg13g2_nand2_1 _8327_ (.Y(_3436_),
    .A(_3290_),
    .B(_3435_));
 sg13g2_nand3_1 _8328_ (.B(net53),
    .C(_3436_),
    .A(_3310_),
    .Y(_3437_));
 sg13g2_or2_1 _8329_ (.X(_3439_),
    .B(_3436_),
    .A(_3310_));
 sg13g2_a21oi_1 _8330_ (.A1(_3437_),
    .A2(_3439_),
    .Y(_0172_),
    .B1(_3317_));
 sg13g2_nand3_1 _8331_ (.B(_3290_),
    .C(_3435_),
    .A(_3310_),
    .Y(_3440_));
 sg13g2_nand3_1 _8332_ (.B(net53),
    .C(_3440_),
    .A(_3340_),
    .Y(_3441_));
 sg13g2_and3_1 _8333_ (.X(_3442_),
    .A(_3310_),
    .B(_3290_),
    .C(_3435_));
 sg13g2_buf_1 _8334_ (.A(_3442_),
    .X(_3443_));
 sg13g2_nand2b_1 _8335_ (.Y(_3444_),
    .B(_3443_),
    .A_N(_3340_));
 sg13g2_a21oi_1 _8336_ (.A1(_3441_),
    .A2(_3444_),
    .Y(_0173_),
    .B1(_3317_));
 sg13g2_nand2_1 _8337_ (.Y(_3445_),
    .A(_4042_),
    .B(net53));
 sg13g2_nand2_1 _8338_ (.Y(_3446_),
    .A(_3340_),
    .B(_3443_));
 sg13g2_xor2_1 _8339_ (.B(_3446_),
    .A(_3349_),
    .X(_3448_));
 sg13g2_nor2_1 _8340_ (.A(_3445_),
    .B(_3448_),
    .Y(_0174_));
 sg13g2_nand2_1 _8341_ (.Y(_3449_),
    .A(\collatz.orbit_len[13] ),
    .B(net53));
 sg13g2_nand3_1 _8342_ (.B(_3349_),
    .C(_3443_),
    .A(_3340_),
    .Y(_3450_));
 sg13g2_mux2_1 _8343_ (.A0(\collatz.orbit_len[13] ),
    .A1(_3449_),
    .S(_3450_),
    .X(_3451_));
 sg13g2_nor2_1 _8344_ (.A(net108),
    .B(_3451_),
    .Y(_0175_));
 sg13g2_nor2_1 _8345_ (.A(_3359_),
    .B(_3440_),
    .Y(_3452_));
 sg13g2_nand3b_1 _8346_ (.B(_3320_),
    .C(net53),
    .Y(_3453_),
    .A_N(_3452_));
 sg13g2_nand2b_1 _8347_ (.Y(_3454_),
    .B(_3452_),
    .A_N(_3320_));
 sg13g2_buf_1 _8348_ (.A(_3964_),
    .X(_3455_));
 sg13g2_a21oi_1 _8349_ (.A1(_3453_),
    .A2(_3454_),
    .Y(_0176_),
    .B1(net85));
 sg13g2_nand2_1 _8350_ (.Y(_3457_),
    .A(_3320_),
    .B(_3452_));
 sg13g2_nand3_1 _8351_ (.B(net53),
    .C(_3457_),
    .A(\collatz.orbit_len[15] ),
    .Y(_3458_));
 sg13g2_or2_1 _8352_ (.X(_3459_),
    .B(_3457_),
    .A(\collatz.orbit_len[15] ));
 sg13g2_a21oi_1 _8353_ (.A1(_3458_),
    .A2(_3459_),
    .Y(_0177_),
    .B1(net85));
 sg13g2_xor2_1 _8354_ (.B(_3201_),
    .A(_3191_),
    .X(_3460_));
 sg13g2_a22oi_1 _8355_ (.Y(_3461_),
    .B1(_3460_),
    .B2(net64),
    .A2(_3431_),
    .A1(_3191_));
 sg13g2_nor2_1 _8356_ (.A(net108),
    .B(_3461_),
    .Y(_0178_));
 sg13g2_nand2_1 _8357_ (.Y(_3462_),
    .A(_3191_),
    .B(_3201_));
 sg13g2_xnor2_1 _8358_ (.Y(_3463_),
    .A(_3211_),
    .B(_3462_));
 sg13g2_a22oi_1 _8359_ (.Y(_3465_),
    .B1(_3463_),
    .B2(_1198_),
    .A2(_3431_),
    .A1(_3211_));
 sg13g2_nor2_1 _8360_ (.A(net108),
    .B(_3465_),
    .Y(_0179_));
 sg13g2_xnor2_1 _8361_ (.Y(_3466_),
    .A(\collatz.orbit_len[3] ),
    .B(_3220_));
 sg13g2_nor3_1 _8362_ (.A(net80),
    .B(_3181_),
    .C(_3959_),
    .Y(_3467_));
 sg13g2_a21oi_1 _8363_ (.A1(net56),
    .A2(_3466_),
    .Y(_3468_),
    .B1(_3467_));
 sg13g2_nor2_1 _8364_ (.A(net108),
    .B(_3468_),
    .Y(_0180_));
 sg13g2_inv_1 _8365_ (.Y(_3469_),
    .A(\collatz.orbit_len[4] ));
 sg13g2_xnor2_1 _8366_ (.Y(_3470_),
    .A(_3469_),
    .B(_3231_));
 sg13g2_nor3_1 _8367_ (.A(net80),
    .B(_3469_),
    .C(_3959_),
    .Y(_3471_));
 sg13g2_a21oi_1 _8368_ (.A1(_2628_),
    .A2(_3470_),
    .Y(_3472_),
    .B1(_3471_));
 sg13g2_nor2_1 _8369_ (.A(net108),
    .B(_3472_),
    .Y(_0181_));
 sg13g2_xnor2_1 _8370_ (.Y(_3474_),
    .A(\collatz.orbit_len[5] ),
    .B(_3241_));
 sg13g2_nor3_1 _8371_ (.A(net80),
    .B(_3171_),
    .C(_3959_),
    .Y(_3475_));
 sg13g2_a21oi_1 _8372_ (.A1(_2628_),
    .A2(_3474_),
    .Y(_3476_),
    .B1(_3475_));
 sg13g2_nor2_1 _8373_ (.A(net108),
    .B(_3476_),
    .Y(_0182_));
 sg13g2_nand2_1 _8374_ (.Y(_3477_),
    .A(_0400_),
    .B(_3251_));
 sg13g2_xor2_1 _8375_ (.B(_3477_),
    .A(_3300_),
    .X(_3478_));
 sg13g2_nor2_1 _8376_ (.A(_3445_),
    .B(_3478_),
    .Y(_0183_));
 sg13g2_nand2_1 _8377_ (.Y(_3479_),
    .A(_3261_),
    .B(net53));
 sg13g2_mux2_1 _8378_ (.A0(_3479_),
    .A1(_3261_),
    .S(_3435_),
    .X(_3480_));
 sg13g2_nor2_1 _8379_ (.A(net108),
    .B(_3480_),
    .Y(_0184_));
 sg13g2_nand2_1 _8380_ (.Y(_3482_),
    .A(_3261_),
    .B(_3435_));
 sg13g2_xor2_1 _8381_ (.B(_3482_),
    .A(_3271_),
    .X(_3483_));
 sg13g2_nor2_1 _8382_ (.A(_3445_),
    .B(_3483_),
    .Y(_0185_));
 sg13g2_nand3_1 _8383_ (.B(_3271_),
    .C(_3435_),
    .A(_3261_),
    .Y(_3484_));
 sg13g2_nand3_1 _8384_ (.B(_3962_),
    .C(_3484_),
    .A(\collatz.orbit_len[9] ),
    .Y(_3485_));
 sg13g2_o21ai_1 _8385_ (.B1(_3485_),
    .Y(_3486_),
    .A1(\collatz.orbit_len[9] ),
    .A2(_3484_));
 sg13g2_and2_1 _8386_ (.A(net270),
    .B(_3486_),
    .X(_0186_));
 sg13g2_xnor2_1 _8387_ (.Y(_3487_),
    .A(net271),
    .B(_2527_));
 sg13g2_nand2b_1 _8388_ (.Y(_3488_),
    .B(net123),
    .A_N(_4020_));
 sg13g2_nand4_1 _8389_ (.B(_4020_),
    .C(_2565_),
    .A(net202),
    .Y(_3490_),
    .D(_2567_));
 sg13g2_mux2_1 _8390_ (.A0(_3488_),
    .A1(_3490_),
    .S(_2563_),
    .X(_3491_));
 sg13g2_xor2_1 _8391_ (.B(_4020_),
    .A(_0000_),
    .X(_3492_));
 sg13g2_a21oi_1 _8392_ (.A1(_2565_),
    .A2(_2567_),
    .Y(_3493_),
    .B1(_3488_));
 sg13g2_a21oi_1 _8393_ (.A1(net113),
    .A2(_3492_),
    .Y(_3494_),
    .B1(_3493_));
 sg13g2_xor2_1 _8394_ (.B(_3832_),
    .A(_3922_),
    .X(_3495_));
 sg13g2_nand3_1 _8395_ (.B(_2605_),
    .C(_3495_),
    .A(net202),
    .Y(_3496_));
 sg13g2_nand2_1 _8396_ (.Y(_3497_),
    .A(_2232_),
    .B(_2607_));
 sg13g2_nand2_1 _8397_ (.Y(_3498_),
    .A(_2586_),
    .B(_2598_));
 sg13g2_mux2_1 _8398_ (.A0(_3496_),
    .A1(_3497_),
    .S(_3498_),
    .X(_3499_));
 sg13g2_o21ai_1 _8399_ (.B1(\collatz.path_record_h16[15] ),
    .Y(_3501_),
    .A1(_2605_),
    .A2(_3497_));
 sg13g2_inv_1 _8400_ (.Y(_3502_),
    .A(_3501_));
 sg13g2_nand2b_1 _8401_ (.Y(_3503_),
    .B(_2232_),
    .A_N(\collatz.path_record_h16[15] ));
 sg13g2_nor2_1 _8402_ (.A(_2607_),
    .B(_3503_),
    .Y(_3504_));
 sg13g2_nor2_1 _8403_ (.A(_3495_),
    .B(_3503_),
    .Y(_3505_));
 sg13g2_mux2_1 _8404_ (.A0(_3504_),
    .A1(_3505_),
    .S(_2606_),
    .X(_3506_));
 sg13g2_a221oi_1 _8405_ (.B2(_3502_),
    .C1(_3506_),
    .B1(_3499_),
    .A1(_3491_),
    .Y(_3507_),
    .A2(_3494_));
 sg13g2_inv_1 _8406_ (.Y(_3508_),
    .A(_0002_));
 sg13g2_xnor2_1 _8407_ (.Y(_3509_),
    .A(_3508_),
    .B(_2499_));
 sg13g2_and3_1 _8408_ (.X(_3510_),
    .A(_3487_),
    .B(_3507_),
    .C(_3509_));
 sg13g2_nand2_1 _8409_ (.Y(_3512_),
    .A(_4009_),
    .B(_2458_));
 sg13g2_nand4_1 _8410_ (.B(_4009_),
    .C(_2454_),
    .A(net81),
    .Y(_3513_),
    .D(_2456_));
 sg13g2_nand2_1 _8411_ (.Y(_3514_),
    .A(_4030_),
    .B(_4009_));
 sg13g2_or3_1 _8412_ (.A(_2454_),
    .B(_2456_),
    .C(_3514_),
    .X(_3515_));
 sg13g2_nand3_1 _8413_ (.B(_3513_),
    .C(_3515_),
    .A(_3512_),
    .Y(_3516_));
 sg13g2_nand2_1 _8414_ (.Y(_3517_),
    .A(_2406_),
    .B(_2430_));
 sg13g2_inv_1 _8415_ (.Y(_3518_),
    .A(\collatz.path_record_h16[9] ));
 sg13g2_or2_1 _8416_ (.X(_3519_),
    .B(_2360_),
    .A(_3996_));
 sg13g2_nor3_1 _8417_ (.A(_2357_),
    .B(_2400_),
    .C(_3519_),
    .Y(_3520_));
 sg13g2_o21ai_1 _8418_ (.B1(_2400_),
    .Y(_3521_),
    .A1(_2357_),
    .A2(_3519_));
 sg13g2_o21ai_1 _8419_ (.B1(_3521_),
    .Y(_3523_),
    .A1(_3518_),
    .A2(_3520_));
 sg13g2_nor2_1 _8420_ (.A(_3517_),
    .B(_3523_),
    .Y(_3524_));
 sg13g2_a21oi_1 _8421_ (.A1(_3517_),
    .A2(_3523_),
    .Y(_3525_),
    .B1(\collatz.path_record_h16[10] ));
 sg13g2_nor2_1 _8422_ (.A(_3524_),
    .B(_3525_),
    .Y(_3526_));
 sg13g2_nand2b_1 _8423_ (.Y(_3527_),
    .B(_2459_),
    .A_N(_4009_));
 sg13g2_o21ai_1 _8424_ (.B1(_3527_),
    .Y(_3528_),
    .A1(_3516_),
    .A2(_3526_));
 sg13g2_or2_1 _8425_ (.X(_3529_),
    .B(_2458_),
    .A(_4009_));
 sg13g2_a21oi_1 _8426_ (.A1(net81),
    .A2(_2457_),
    .Y(_3530_),
    .B1(_3529_));
 sg13g2_xor2_1 _8427_ (.B(_2361_),
    .A(_3996_),
    .X(_3531_));
 sg13g2_nor3_1 _8428_ (.A(_3530_),
    .B(_3516_),
    .C(_3531_),
    .Y(_3532_));
 sg13g2_inv_1 _8429_ (.Y(_3534_),
    .A(\collatz.path_record_h16[10] ));
 sg13g2_nand3_1 _8430_ (.B(_2406_),
    .C(_2430_),
    .A(_3534_),
    .Y(_3535_));
 sg13g2_a21o_1 _8431_ (.A2(_2430_),
    .A1(_2406_),
    .B1(_3534_),
    .X(_3536_));
 sg13g2_xnor2_1 _8432_ (.Y(_3537_),
    .A(_3518_),
    .B(_2400_));
 sg13g2_and4_1 _8433_ (.A(_3510_),
    .B(_3535_),
    .C(_3536_),
    .D(_3537_),
    .X(_3538_));
 sg13g2_nand2_1 _8434_ (.Y(_3539_),
    .A(_3532_),
    .B(_3538_));
 sg13g2_nor2b_1 _8435_ (.A(_2335_),
    .B_N(_4023_),
    .Y(_3540_));
 sg13g2_nor4_1 _8436_ (.A(_4023_),
    .B(_2321_),
    .C(_2332_),
    .D(_2334_),
    .Y(_3541_));
 sg13g2_nand2b_1 _8437_ (.Y(_3542_),
    .B(\collatz.path_record_h16[3] ),
    .A_N(_2167_));
 sg13g2_xnor2_1 _8438_ (.Y(_3543_),
    .A(_4015_),
    .B(_2258_));
 sg13g2_xnor2_1 _8439_ (.Y(_3545_),
    .A(_4019_),
    .B(_2301_));
 sg13g2_xnor2_1 _8440_ (.Y(_3546_),
    .A(_4012_),
    .B(_2213_));
 sg13g2_nand4_1 _8441_ (.B(_3543_),
    .C(_3545_),
    .A(_3542_),
    .Y(_3547_),
    .D(_3546_));
 sg13g2_nor4_2 _8442_ (.A(_3539_),
    .B(_3540_),
    .C(_3541_),
    .Y(_3548_),
    .D(_3547_));
 sg13g2_nand2b_1 _8443_ (.Y(_3549_),
    .B(_2167_),
    .A_N(\collatz.path_record_h16[3] ));
 sg13g2_nand2_1 _8444_ (.Y(_3550_),
    .A(_3995_),
    .B(_2074_));
 sg13g2_inv_1 _8445_ (.Y(_3551_),
    .A(\collatz.path_record_h16[1] ));
 sg13g2_o21ai_1 _8446_ (.B1(_3551_),
    .Y(_3552_),
    .A1(_2040_),
    .A2(_3550_));
 sg13g2_inv_1 _8447_ (.Y(_3553_),
    .A(_3995_));
 sg13g2_o21ai_1 _8448_ (.B1(_2075_),
    .Y(_3554_),
    .A1(_3553_),
    .A2(_2040_));
 sg13g2_and2_1 _8449_ (.A(_4006_),
    .B(_2124_),
    .X(_3556_));
 sg13g2_buf_1 _8450_ (.A(_3556_),
    .X(_3557_));
 sg13g2_and2_1 _8451_ (.A(_2123_),
    .B(_3557_),
    .X(_3558_));
 sg13g2_a21o_1 _8452_ (.A2(_3554_),
    .A1(_3552_),
    .B1(_3558_),
    .X(_3559_));
 sg13g2_or2_1 _8453_ (.X(_3560_),
    .B(_2125_),
    .A(_4006_));
 sg13g2_nand3_1 _8454_ (.B(_3559_),
    .C(_3560_),
    .A(_3549_),
    .Y(_3561_));
 sg13g2_nand2b_1 _8455_ (.Y(_3562_),
    .B(_4023_),
    .A_N(_2335_));
 sg13g2_inv_1 _8456_ (.Y(_3563_),
    .A(_2258_));
 sg13g2_inv_1 _8457_ (.Y(_3564_),
    .A(_2301_));
 sg13g2_nand2b_1 _8458_ (.Y(_3565_),
    .B(_2213_),
    .A_N(_4012_));
 sg13g2_a221oi_1 _8459_ (.B2(_4019_),
    .C1(_3565_),
    .B1(_3564_),
    .A1(_4015_),
    .Y(_3567_),
    .A2(_3563_));
 sg13g2_nor3_1 _8460_ (.A(_4019_),
    .B(_4015_),
    .C(_3563_),
    .Y(_3568_));
 sg13g2_nand2b_1 _8461_ (.Y(_3569_),
    .B(_2258_),
    .A_N(_4015_));
 sg13g2_a21oi_1 _8462_ (.A1(_4019_),
    .A2(_3569_),
    .Y(_3570_),
    .B1(_3564_));
 sg13g2_or4_1 _8463_ (.A(_3541_),
    .B(_3567_),
    .C(_3568_),
    .D(_3570_),
    .X(_3571_));
 sg13g2_nand4_1 _8464_ (.B(_3538_),
    .C(_3562_),
    .A(_3532_),
    .Y(_3572_),
    .D(_3571_));
 sg13g2_inv_1 _8465_ (.Y(_3573_),
    .A(_2515_));
 sg13g2_nand2_1 _8466_ (.Y(_3574_),
    .A(_3573_),
    .B(_2520_));
 sg13g2_a21oi_1 _8467_ (.A1(_2255_),
    .A2(_2233_),
    .Y(_3575_),
    .B1(_3574_));
 sg13g2_or4_1 _8468_ (.A(_2237_),
    .B(_2246_),
    .C(_2249_),
    .D(_2254_),
    .X(_3576_));
 sg13g2_nor4_1 _8469_ (.A(_3576_),
    .B(_2228_),
    .C(_2513_),
    .D(_3573_),
    .Y(_3578_));
 sg13g2_o21ai_1 _8470_ (.B1(net81),
    .Y(_3579_),
    .A1(_3575_),
    .A2(_3578_));
 sg13g2_nand2_1 _8471_ (.Y(_3580_),
    .A(_2515_),
    .B(_2519_));
 sg13g2_mux2_1 _8472_ (.A0(_3580_),
    .A1(_2515_),
    .S(_2513_),
    .X(_3581_));
 sg13g2_nand2b_1 _8473_ (.Y(_3582_),
    .B(_0002_),
    .A_N(_0003_));
 sg13g2_a21oi_1 _8474_ (.A1(_0001_),
    .A2(net271),
    .Y(_3583_),
    .B1(_3582_));
 sg13g2_nor2_1 _8475_ (.A(_0001_),
    .B(net271),
    .Y(_3584_));
 sg13g2_nor3_1 _8476_ (.A(_4030_),
    .B(_3583_),
    .C(_3584_),
    .Y(_3585_));
 sg13g2_a21o_1 _8477_ (.A2(_3581_),
    .A1(net81),
    .B1(_3585_),
    .X(_3586_));
 sg13g2_or3_1 _8478_ (.A(_4031_),
    .B(_0001_),
    .C(_3582_),
    .X(_3587_));
 sg13g2_a22oi_1 _8479_ (.Y(_3589_),
    .B1(_3587_),
    .B2(net271),
    .A2(_3586_),
    .A1(_3579_));
 sg13g2_inv_1 _8480_ (.Y(_3590_),
    .A(_2484_));
 sg13g2_a21oi_1 _8481_ (.A1(_1481_),
    .A2(_3590_),
    .Y(_3591_),
    .B1(_2493_));
 sg13g2_xor2_1 _8482_ (.B(_3591_),
    .A(_2478_),
    .X(_3592_));
 sg13g2_nand2b_1 _8483_ (.Y(_3593_),
    .B(_0002_),
    .A_N(net271));
 sg13g2_nand3_1 _8484_ (.B(_3581_),
    .C(_3593_),
    .A(_4031_),
    .Y(_3594_));
 sg13g2_nand2b_1 _8485_ (.Y(_3595_),
    .B(_3594_),
    .A_N(_3585_));
 sg13g2_a221oi_1 _8486_ (.B2(_3595_),
    .C1(_2569_),
    .B1(_3579_),
    .A1(net271),
    .Y(_3596_),
    .A2(_3508_));
 sg13g2_o21ai_1 _8487_ (.B1(_3596_),
    .Y(_3597_),
    .A1(_3589_),
    .A2(_3592_));
 sg13g2_a22oi_1 _8488_ (.Y(_3598_),
    .B1(_3579_),
    .B2(_3595_),
    .A2(_3508_),
    .A1(net271));
 sg13g2_o21ai_1 _8489_ (.B1(_3598_),
    .Y(_3600_),
    .A1(_3589_),
    .A2(_3592_));
 sg13g2_a22oi_1 _8490_ (.Y(_3601_),
    .B1(_3600_),
    .B2(_2569_),
    .A2(_3597_),
    .A1(_4020_));
 sg13g2_nand2_1 _8491_ (.Y(_3602_),
    .A(_3499_),
    .B(_3502_));
 sg13g2_o21ai_1 _8492_ (.B1(_3602_),
    .Y(_3603_),
    .A1(_3506_),
    .A2(_3601_));
 sg13g2_nand3_1 _8493_ (.B(_3572_),
    .C(_3603_),
    .A(_3962_),
    .Y(_3604_));
 sg13g2_a221oi_1 _8494_ (.B2(_3561_),
    .C1(_3604_),
    .B1(_3548_),
    .A1(_3510_),
    .Y(_3605_),
    .A2(_3528_));
 sg13g2_buf_8 _8495_ (.A(_3605_),
    .X(_3606_));
 sg13g2_buf_8 _8496_ (.A(_3606_),
    .X(_3607_));
 sg13g2_xnor2_1 _8497_ (.Y(_3608_),
    .A(net127),
    .B(_2090_));
 sg13g2_nor2_1 _8498_ (.A(net84),
    .B(_4006_),
    .Y(_3609_));
 sg13g2_nand3_1 _8499_ (.B(_2120_),
    .C(_3609_),
    .A(_3608_),
    .Y(_3611_));
 sg13g2_nand2_1 _8500_ (.Y(_3612_),
    .A(_2091_),
    .B(_3609_));
 sg13g2_nor2_1 _8501_ (.A(_2097_),
    .B(_2116_),
    .Y(_3613_));
 sg13g2_mux2_1 _8502_ (.A0(_3611_),
    .A1(_3612_),
    .S(_3613_),
    .X(_3614_));
 sg13g2_nand3_1 _8503_ (.B(_2120_),
    .C(_3557_),
    .A(_2091_),
    .Y(_3615_));
 sg13g2_nand2_1 _8504_ (.Y(_3616_),
    .A(_3608_),
    .B(_3557_));
 sg13g2_mux2_1 _8505_ (.A0(_3615_),
    .A1(_3616_),
    .S(_3613_),
    .X(_3617_));
 sg13g2_xnor2_1 _8506_ (.Y(_3618_),
    .A(_3551_),
    .B(_2074_));
 sg13g2_xnor2_1 _8507_ (.Y(_3619_),
    .A(_0013_),
    .B(_4006_));
 sg13g2_a21oi_1 _8508_ (.A1(_3612_),
    .A2(_3616_),
    .Y(_3620_),
    .B1(_2120_));
 sg13g2_a21oi_1 _8509_ (.A1(net84),
    .A2(_3619_),
    .Y(_3622_),
    .B1(_3620_));
 sg13g2_and4_1 _8510_ (.A(_3961_),
    .B(_3549_),
    .C(_3618_),
    .D(_3622_),
    .X(_3623_));
 sg13g2_xnor2_1 _8511_ (.Y(_3624_),
    .A(_3995_),
    .B(_2040_));
 sg13g2_and4_1 _8512_ (.A(_3614_),
    .B(_3617_),
    .C(_3623_),
    .D(_3624_),
    .X(_3625_));
 sg13g2_a21oi_1 _8513_ (.A1(_3956_),
    .A2(_3959_),
    .Y(_3626_),
    .B1(_3161_));
 sg13g2_a21o_1 _8514_ (.A2(_3625_),
    .A1(_3548_),
    .B1(_3626_),
    .X(_3627_));
 sg13g2_buf_8 _8515_ (.A(_3627_),
    .X(_3628_));
 sg13g2_buf_1 _8516_ (.A(_3628_),
    .X(_3629_));
 sg13g2_o21ai_1 _8517_ (.B1(_3995_),
    .Y(_3630_),
    .A1(net17),
    .A2(net16));
 sg13g2_buf_8 _8518_ (.A(_3606_),
    .X(_3631_));
 sg13g2_a21oi_1 _8519_ (.A1(_3548_),
    .A2(_3625_),
    .Y(_3633_),
    .B1(_3626_));
 sg13g2_buf_2 _8520_ (.A(_3633_),
    .X(_3634_));
 sg13g2_buf_1 _8521_ (.A(_3634_),
    .X(_3635_));
 sg13g2_o21ai_1 _8522_ (.B1(_2041_),
    .Y(_3636_),
    .A1(_2052_),
    .A2(net95));
 sg13g2_nand3b_1 _8523_ (.B(net14),
    .C(_3636_),
    .Y(_3637_),
    .A_N(net15));
 sg13g2_a21oi_1 _8524_ (.A1(_3630_),
    .A2(_3637_),
    .Y(_0187_),
    .B1(net85));
 sg13g2_o21ai_1 _8525_ (.B1(\collatz.path_record_h16[10] ),
    .Y(_3638_),
    .A1(_3607_),
    .A2(_3629_));
 sg13g2_o21ai_1 _8526_ (.B1(_2431_),
    .Y(_3639_),
    .A1(_2432_),
    .A2(_0703_));
 sg13g2_nand3b_1 _8527_ (.B(net14),
    .C(_3639_),
    .Y(_3640_),
    .A_N(net15));
 sg13g2_a21oi_1 _8528_ (.A1(_3638_),
    .A2(_3640_),
    .Y(_0188_),
    .B1(net85));
 sg13g2_o21ai_1 _8529_ (.B1(_4009_),
    .Y(_3642_),
    .A1(_3607_),
    .A2(_3629_));
 sg13g2_o21ai_1 _8530_ (.B1(_2460_),
    .Y(_3643_),
    .A1(_2461_),
    .A2(net95));
 sg13g2_nand3b_1 _8531_ (.B(_3635_),
    .C(_3643_),
    .Y(_3644_),
    .A_N(net15));
 sg13g2_a21oi_1 _8532_ (.A1(_3642_),
    .A2(_3644_),
    .Y(_0189_),
    .B1(net85));
 sg13g2_o21ai_1 _8533_ (.B1(\collatz.path_record_h16[12] ),
    .Y(_3645_),
    .A1(net17),
    .A2(net16));
 sg13g2_o21ai_1 _8534_ (.B1(_2500_),
    .Y(_3646_),
    .A1(_3831_),
    .A2(_0703_));
 sg13g2_nand3b_1 _8535_ (.B(net14),
    .C(_3646_),
    .Y(_3647_),
    .A_N(net15));
 sg13g2_a21oi_1 _8536_ (.A1(_3645_),
    .A2(_3647_),
    .Y(_0190_),
    .B1(net85));
 sg13g2_o21ai_1 _8537_ (.B1(net271),
    .Y(_3648_),
    .A1(net17),
    .A2(net16));
 sg13g2_o21ai_1 _8538_ (.B1(_2528_),
    .Y(_3649_),
    .A1(_2529_),
    .A2(net95));
 sg13g2_nand3b_1 _8539_ (.B(_3635_),
    .C(_3649_),
    .Y(_3651_),
    .A_N(_3631_));
 sg13g2_a21oi_1 _8540_ (.A1(_3648_),
    .A2(_3651_),
    .Y(_0191_),
    .B1(_3455_));
 sg13g2_and2_1 _8541_ (.A(_3956_),
    .B(_4020_),
    .X(_3652_));
 sg13g2_a21oi_1 _8542_ (.A1(_3833_),
    .A2(net77),
    .Y(_3653_),
    .B1(_2570_));
 sg13g2_nor2_1 _8543_ (.A(_3606_),
    .B(_3628_),
    .Y(_3654_));
 sg13g2_mux2_1 _8544_ (.A0(_3652_),
    .A1(_3653_),
    .S(_3654_),
    .X(_0192_));
 sg13g2_o21ai_1 _8545_ (.B1(\collatz.path_record_h16[15] ),
    .Y(_3655_),
    .A1(net17),
    .A2(net16));
 sg13g2_buf_8 _8546_ (.A(_3606_),
    .X(_3656_));
 sg13g2_o21ai_1 _8547_ (.B1(_2609_),
    .Y(_3657_),
    .A1(_2610_),
    .A2(net95));
 sg13g2_nand3b_1 _8548_ (.B(net14),
    .C(_3657_),
    .Y(_3658_),
    .A_N(_3656_));
 sg13g2_a21oi_1 _8549_ (.A1(_3655_),
    .A2(_3658_),
    .Y(_0193_),
    .B1(_3455_));
 sg13g2_o21ai_1 _8550_ (.B1(\collatz.path_record_h16[1] ),
    .Y(_3660_),
    .A1(net17),
    .A2(net16));
 sg13g2_o21ai_1 _8551_ (.B1(_2076_),
    .Y(_3661_),
    .A1(_2099_),
    .A2(net95));
 sg13g2_nand3b_1 _8552_ (.B(net14),
    .C(_3661_),
    .Y(_3662_),
    .A_N(net13));
 sg13g2_a21oi_1 _8553_ (.A1(_3660_),
    .A2(_3662_),
    .Y(_0194_),
    .B1(net85));
 sg13g2_o21ai_1 _8554_ (.B1(_4006_),
    .Y(_3663_),
    .A1(net17),
    .A2(net16));
 sg13g2_o21ai_1 _8555_ (.B1(_2126_),
    .Y(_3664_),
    .A1(_2219_),
    .A2(net95));
 sg13g2_nand3b_1 _8556_ (.B(net14),
    .C(_3664_),
    .Y(_3665_),
    .A_N(net13));
 sg13g2_a21oi_1 _8557_ (.A1(_3663_),
    .A2(_3665_),
    .Y(_0195_),
    .B1(net85));
 sg13g2_o21ai_1 _8558_ (.B1(\collatz.path_record_h16[3] ),
    .Y(_3666_),
    .A1(net17),
    .A2(net16));
 sg13g2_o21ai_1 _8559_ (.B1(_2168_),
    .Y(_3668_),
    .A1(_2306_),
    .A2(net102));
 sg13g2_nand3b_1 _8560_ (.B(net14),
    .C(_3668_),
    .Y(_3669_),
    .A_N(net13));
 sg13g2_a21oi_1 _8561_ (.A1(_3666_),
    .A2(_3669_),
    .Y(_0196_),
    .B1(net99));
 sg13g2_o21ai_1 _8562_ (.B1(_4012_),
    .Y(_3670_),
    .A1(net17),
    .A2(net16));
 sg13g2_o21ai_1 _8563_ (.B1(_2214_),
    .Y(_3671_),
    .A1(_2220_),
    .A2(net102));
 sg13g2_nand3b_1 _8564_ (.B(net14),
    .C(_3671_),
    .Y(_3672_),
    .A_N(net13));
 sg13g2_a21oi_1 _8565_ (.A1(_3670_),
    .A2(_3672_),
    .Y(_0197_),
    .B1(net99));
 sg13g2_o21ai_1 _8566_ (.B1(_4015_),
    .Y(_3673_),
    .A1(net15),
    .A2(_3628_));
 sg13g2_o21ai_1 _8567_ (.B1(_2259_),
    .Y(_3674_),
    .A1(_2307_),
    .A2(net102));
 sg13g2_nand3b_1 _8568_ (.B(_3634_),
    .C(_3674_),
    .Y(_3675_),
    .A_N(net13));
 sg13g2_a21oi_1 _8569_ (.A1(_3673_),
    .A2(_3675_),
    .Y(_0198_),
    .B1(net99));
 sg13g2_o21ai_1 _8570_ (.B1(_4019_),
    .Y(_3677_),
    .A1(net15),
    .A2(_3628_));
 sg13g2_o21ai_1 _8571_ (.B1(_2302_),
    .Y(_3678_),
    .A1(_2341_),
    .A2(net102));
 sg13g2_nand3b_1 _8572_ (.B(_3634_),
    .C(_3678_),
    .Y(_3679_),
    .A_N(net13));
 sg13g2_a21oi_1 _8573_ (.A1(_3677_),
    .A2(_3679_),
    .Y(_0199_),
    .B1(net99));
 sg13g2_o21ai_1 _8574_ (.B1(_4023_),
    .Y(_3680_),
    .A1(net15),
    .A2(_3628_));
 sg13g2_o21ai_1 _8575_ (.B1(_2336_),
    .Y(_3681_),
    .A1(_2339_),
    .A2(net102));
 sg13g2_nand3b_1 _8576_ (.B(_3634_),
    .C(_3681_),
    .Y(_3682_),
    .A_N(net13));
 sg13g2_a21oi_1 _8577_ (.A1(_3680_),
    .A2(_3682_),
    .Y(_0200_),
    .B1(net99));
 sg13g2_o21ai_1 _8578_ (.B1(_3996_),
    .Y(_3683_),
    .A1(net15),
    .A2(_3628_));
 sg13g2_o21ai_1 _8579_ (.B1(_2362_),
    .Y(_3685_),
    .A1(_2364_),
    .A2(_4044_));
 sg13g2_nand3b_1 _8580_ (.B(_3634_),
    .C(_3685_),
    .Y(_3686_),
    .A_N(net13));
 sg13g2_a21oi_1 _8581_ (.A1(_3683_),
    .A2(_3686_),
    .Y(_0201_),
    .B1(net99));
 sg13g2_o21ai_1 _8582_ (.B1(\collatz.path_record_h16[9] ),
    .Y(_3687_),
    .A1(_3631_),
    .A2(_3628_));
 sg13g2_o21ai_1 _8583_ (.B1(_2401_),
    .Y(_3688_),
    .A1(_2402_),
    .A2(_4044_));
 sg13g2_nand3b_1 _8584_ (.B(_3634_),
    .C(_3688_),
    .Y(_3689_),
    .A_N(_3656_));
 sg13g2_a21oi_1 _8585_ (.A1(_3687_),
    .A2(_3689_),
    .Y(_0202_),
    .B1(net99));
 sg13g2_dfrbp_1 _8586_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net344),
    .D(_0018_),
    .Q_N(_4383_),
    .Q(\collatz.iter[1] ));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _8586__344 (.L_HI(net344));
 sg13g2_buf_1 _8589_ (.A(net330),
    .X(uio_oe[0]));
 sg13g2_buf_1 _8590_ (.A(net331),
    .X(uio_oe[1]));
 sg13g2_buf_1 _8591_ (.A(net332),
    .X(uio_oe[2]));
 sg13g2_buf_1 _8592_ (.A(net333),
    .X(uio_oe[3]));
 sg13g2_buf_1 _8593_ (.A(net334),
    .X(uio_oe[4]));
 sg13g2_buf_1 _8594_ (.A(net335),
    .X(uio_oe[5]));
 sg13g2_buf_1 _8595_ (.A(net336),
    .X(uio_oe[6]));
 sg13g2_buf_1 _8596_ (.A(\collatz.comp ),
    .X(net3));
 sg13g2_buf_1 _8597_ (.A(net337),
    .X(uio_out[0]));
 sg13g2_buf_1 _8598_ (.A(net338),
    .X(uio_out[1]));
 sg13g2_buf_1 _8599_ (.A(net339),
    .X(uio_out[2]));
 sg13g2_buf_1 _8600_ (.A(net340),
    .X(uio_out[3]));
 sg13g2_buf_1 _8601_ (.A(net341),
    .X(uio_out[4]));
 sg13g2_buf_1 _8602_ (.A(net342),
    .X(uio_out[5]));
 sg13g2_buf_1 _8603_ (.A(net343),
    .X(uio_out[6]));
 sg13g2_buf_1 _8604_ (.A(\collatz.busy ),
    .X(net4));
 sg13g2_dfrbp_1 \data_out[0]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net345),
    .D(_0019_),
    .Q_N(_4382_),
    .Q(net5));
 sg13g2_dfrbp_1 \data_out[1]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net346),
    .D(_0020_),
    .Q_N(_4381_),
    .Q(net6));
 sg13g2_dfrbp_1 \data_out[2]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net347),
    .D(_0021_),
    .Q_N(_4380_),
    .Q(net7));
 sg13g2_dfrbp_1 \data_out[3]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net348),
    .D(_0022_),
    .Q_N(_4379_),
    .Q(net8));
 sg13g2_dfrbp_1 \data_out[4]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net349),
    .D(_0023_),
    .Q_N(_4378_),
    .Q(net9));
 sg13g2_dfrbp_1 \data_out[5]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net350),
    .D(_0024_),
    .Q_N(_4377_),
    .Q(net10));
 sg13g2_dfrbp_1 \data_out[6]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net351),
    .D(_0025_),
    .Q_N(_4376_),
    .Q(net11));
 sg13g2_dfrbp_1 \data_out[7]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net352),
    .D(_0026_),
    .Q_N(_4375_),
    .Q(net12));
 sg13g2_dfrbp_1 \ioctl[7]$_SDFFE_PP0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net353),
    .D(_0027_),
    .Q_N(_0017_),
    .Q(\collatz.comp ));
 sg13g2_dfrbp_1 \iter[0]$_SDFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net354),
    .D(_0028_),
    .Q_N(_0016_),
    .Q(\collatz.iter[0] ));
 sg13g2_dfrbp_1 \iter[100]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net355),
    .D(_0029_),
    .Q_N(_4374_),
    .Q(\collatz.iter[100] ));
 sg13g2_dfrbp_1 \iter[101]$_SDFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net356),
    .D(_0030_),
    .Q_N(_4373_),
    .Q(\collatz.iter[101] ));
 sg13g2_dfrbp_1 \iter[102]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net357),
    .D(_0031_),
    .Q_N(_4372_),
    .Q(\collatz.iter[102] ));
 sg13g2_dfrbp_1 \iter[103]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net358),
    .D(_0032_),
    .Q_N(_4371_),
    .Q(\collatz.iter[103] ));
 sg13g2_dfrbp_1 \iter[104]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net359),
    .D(_0033_),
    .Q_N(_4370_),
    .Q(\collatz.iter[104] ));
 sg13g2_dfrbp_1 \iter[105]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net360),
    .D(_0034_),
    .Q_N(_4369_),
    .Q(\collatz.iter[105] ));
 sg13g2_dfrbp_1 \iter[106]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net361),
    .D(_0035_),
    .Q_N(_4368_),
    .Q(\collatz.iter[106] ));
 sg13g2_dfrbp_1 \iter[107]$_SDFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net362),
    .D(_0036_),
    .Q_N(_4367_),
    .Q(\collatz.iter[107] ));
 sg13g2_dfrbp_1 \iter[108]$_SDFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net363),
    .D(_0037_),
    .Q_N(_4366_),
    .Q(\collatz.iter[108] ));
 sg13g2_dfrbp_1 \iter[109]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net364),
    .D(_0038_),
    .Q_N(_4365_),
    .Q(\collatz.iter[109] ));
 sg13g2_dfrbp_1 \iter[10]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net365),
    .D(_0039_),
    .Q_N(_4364_),
    .Q(\collatz.iter[10] ));
 sg13g2_dfrbp_1 \iter[110]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net366),
    .D(_0040_),
    .Q_N(_4363_),
    .Q(\collatz.iter[110] ));
 sg13g2_dfrbp_1 \iter[111]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net367),
    .D(_0041_),
    .Q_N(_4362_),
    .Q(\collatz.iter[111] ));
 sg13g2_dfrbp_1 \iter[112]$_SDFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net368),
    .D(_0042_),
    .Q_N(_4361_),
    .Q(\collatz.iter[112] ));
 sg13g2_dfrbp_1 \iter[113]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net369),
    .D(_0043_),
    .Q_N(_4360_),
    .Q(\collatz.iter[113] ));
 sg13g2_dfrbp_1 \iter[114]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net370),
    .D(_0044_),
    .Q_N(_4359_),
    .Q(\collatz.iter[114] ));
 sg13g2_dfrbp_1 \iter[115]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net371),
    .D(_0045_),
    .Q_N(_4358_),
    .Q(\collatz.iter[115] ));
 sg13g2_dfrbp_1 \iter[116]$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net372),
    .D(_0046_),
    .Q_N(_4357_),
    .Q(\collatz.iter[116] ));
 sg13g2_dfrbp_1 \iter[117]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net373),
    .D(_0047_),
    .Q_N(_4356_),
    .Q(\collatz.iter[117] ));
 sg13g2_dfrbp_1 \iter[118]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net374),
    .D(_0048_),
    .Q_N(_4355_),
    .Q(\collatz.iter[118] ));
 sg13g2_dfrbp_1 \iter[119]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net375),
    .D(_0049_),
    .Q_N(_4354_),
    .Q(\collatz.iter[119] ));
 sg13g2_dfrbp_1 \iter[11]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net376),
    .D(_0050_),
    .Q_N(_4353_),
    .Q(\collatz.iter[11] ));
 sg13g2_dfrbp_1 \iter[120]$_SDFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net377),
    .D(_0051_),
    .Q_N(_4352_),
    .Q(\collatz.iter[120] ));
 sg13g2_dfrbp_1 \iter[121]$_SDFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net378),
    .D(_0052_),
    .Q_N(_4351_),
    .Q(\collatz.iter[121] ));
 sg13g2_dfrbp_1 \iter[122]$_SDFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net379),
    .D(_0053_),
    .Q_N(_4350_),
    .Q(\collatz.iter[122] ));
 sg13g2_dfrbp_1 \iter[123]$_SDFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net380),
    .D(_0054_),
    .Q_N(_4349_),
    .Q(\collatz.iter[123] ));
 sg13g2_dfrbp_1 \iter[124]$_SDFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net381),
    .D(_0055_),
    .Q_N(_4348_),
    .Q(\collatz.iter[124] ));
 sg13g2_dfrbp_1 \iter[125]$_SDFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net382),
    .D(_0056_),
    .Q_N(_4347_),
    .Q(\collatz.iter[125] ));
 sg13g2_dfrbp_1 \iter[126]$_SDFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net383),
    .D(_0057_),
    .Q_N(_4346_),
    .Q(\collatz.iter[126] ));
 sg13g2_dfrbp_1 \iter[127]$_SDFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net384),
    .D(_0058_),
    .Q_N(_4345_),
    .Q(\collatz.iter[127] ));
 sg13g2_dfrbp_1 \iter[128]$_SDFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net385),
    .D(_0059_),
    .Q_N(_4344_),
    .Q(\collatz.iter[128] ));
 sg13g2_dfrbp_1 \iter[129]$_SDFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net386),
    .D(_0060_),
    .Q_N(_0015_),
    .Q(\collatz.iter[129] ));
 sg13g2_dfrbp_1 \iter[12]$_SDFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net387),
    .D(_0061_),
    .Q_N(_4343_),
    .Q(\collatz.iter[12] ));
 sg13g2_dfrbp_1 \iter[130]$_SDFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net388),
    .D(_0062_),
    .Q_N(_0014_),
    .Q(\collatz.iter[130] ));
 sg13g2_dfrbp_1 \iter[131]$_SDFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net389),
    .D(_0063_),
    .Q_N(_0013_),
    .Q(\collatz.iter[131] ));
 sg13g2_dfrbp_1 \iter[132]$_SDFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net390),
    .D(_0064_),
    .Q_N(_0012_),
    .Q(\collatz.iter[132] ));
 sg13g2_dfrbp_1 \iter[133]$_SDFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net391),
    .D(_0065_),
    .Q_N(_0011_),
    .Q(\collatz.iter[133] ));
 sg13g2_dfrbp_1 \iter[134]$_SDFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net392),
    .D(_0066_),
    .Q_N(_0010_),
    .Q(\collatz.iter[134] ));
 sg13g2_dfrbp_1 \iter[135]$_SDFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net393),
    .D(_0067_),
    .Q_N(_0009_),
    .Q(\collatz.iter[135] ));
 sg13g2_dfrbp_1 \iter[136]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net394),
    .D(_0068_),
    .Q_N(_0008_),
    .Q(\collatz.iter[136] ));
 sg13g2_dfrbp_1 \iter[137]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net395),
    .D(_0069_),
    .Q_N(_0007_),
    .Q(\collatz.iter[137] ));
 sg13g2_dfrbp_1 \iter[138]$_SDFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net396),
    .D(_0070_),
    .Q_N(_0006_),
    .Q(\collatz.iter[138] ));
 sg13g2_dfrbp_1 \iter[139]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net397),
    .D(_0071_),
    .Q_N(_0005_),
    .Q(\collatz.iter[139] ));
 sg13g2_dfrbp_1 \iter[13]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net398),
    .D(_0072_),
    .Q_N(_4342_),
    .Q(\collatz.iter[13] ));
 sg13g2_dfrbp_1 \iter[140]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net399),
    .D(_0073_),
    .Q_N(_0004_),
    .Q(\collatz.iter[140] ));
 sg13g2_dfrbp_1 \iter[141]$_SDFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net400),
    .D(_0074_),
    .Q_N(_0003_),
    .Q(\collatz.iter[141] ));
 sg13g2_dfrbp_1 \iter[142]$_SDFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net401),
    .D(_0075_),
    .Q_N(_0001_),
    .Q(\collatz.iter[142] ));
 sg13g2_dfrbp_1 \iter[143]$_SDFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net402),
    .D(_0076_),
    .Q_N(_0000_),
    .Q(\collatz.iter[143] ));
 sg13g2_dfrbp_1 \iter[14]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net403),
    .D(_0077_),
    .Q_N(_4341_),
    .Q(\collatz.iter[14] ));
 sg13g2_dfrbp_1 \iter[15]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net404),
    .D(_0078_),
    .Q_N(_4340_),
    .Q(\collatz.iter[15] ));
 sg13g2_dfrbp_1 \iter[16]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net405),
    .D(_0079_),
    .Q_N(_4339_),
    .Q(\collatz.iter[16] ));
 sg13g2_dfrbp_1 \iter[17]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net406),
    .D(_0080_),
    .Q_N(_4338_),
    .Q(\collatz.iter[17] ));
 sg13g2_dfrbp_1 \iter[18]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net407),
    .D(_0081_),
    .Q_N(_4337_),
    .Q(\collatz.iter[18] ));
 sg13g2_dfrbp_1 \iter[19]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net408),
    .D(_0082_),
    .Q_N(_4336_),
    .Q(\collatz.iter[19] ));
 sg13g2_dfrbp_1 \iter[20]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net409),
    .D(_0083_),
    .Q_N(_4335_),
    .Q(\collatz.iter[20] ));
 sg13g2_dfrbp_1 \iter[21]$_SDFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net410),
    .D(_0084_),
    .Q_N(_4334_),
    .Q(\collatz.iter[21] ));
 sg13g2_dfrbp_1 \iter[22]$_SDFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net411),
    .D(_0085_),
    .Q_N(_4333_),
    .Q(\collatz.iter[22] ));
 sg13g2_dfrbp_1 \iter[23]$_SDFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net412),
    .D(_0086_),
    .Q_N(_4332_),
    .Q(\collatz.iter[23] ));
 sg13g2_dfrbp_1 \iter[24]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net413),
    .D(_0087_),
    .Q_N(_4331_),
    .Q(\collatz.iter[24] ));
 sg13g2_dfrbp_1 \iter[25]$_SDFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net414),
    .D(_0088_),
    .Q_N(_4330_),
    .Q(\collatz.iter[25] ));
 sg13g2_dfrbp_1 \iter[26]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net415),
    .D(_0089_),
    .Q_N(_4329_),
    .Q(\collatz.iter[26] ));
 sg13g2_dfrbp_1 \iter[27]$_SDFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net416),
    .D(_0090_),
    .Q_N(_4328_),
    .Q(\collatz.iter[27] ));
 sg13g2_dfrbp_1 \iter[28]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net417),
    .D(_0091_),
    .Q_N(_4327_),
    .Q(\collatz.iter[28] ));
 sg13g2_dfrbp_1 \iter[29]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net418),
    .D(_0092_),
    .Q_N(_4326_),
    .Q(\collatz.iter[29] ));
 sg13g2_dfrbp_1 \iter[2]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net419),
    .D(_0093_),
    .Q_N(_4325_),
    .Q(\collatz.iter[2] ));
 sg13g2_dfrbp_1 \iter[30]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net420),
    .D(_0094_),
    .Q_N(_4324_),
    .Q(\collatz.iter[30] ));
 sg13g2_dfrbp_1 \iter[31]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net421),
    .D(_0095_),
    .Q_N(_4323_),
    .Q(\collatz.iter[31] ));
 sg13g2_dfrbp_1 \iter[32]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net422),
    .D(_0096_),
    .Q_N(_4322_),
    .Q(\collatz.iter[32] ));
 sg13g2_dfrbp_1 \iter[33]$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net423),
    .D(_0097_),
    .Q_N(_4321_),
    .Q(\collatz.iter[33] ));
 sg13g2_dfrbp_1 \iter[34]$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net424),
    .D(_0098_),
    .Q_N(_4320_),
    .Q(\collatz.iter[34] ));
 sg13g2_dfrbp_1 \iter[35]$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net425),
    .D(_0099_),
    .Q_N(_4319_),
    .Q(\collatz.iter[35] ));
 sg13g2_dfrbp_1 \iter[36]$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net426),
    .D(_0100_),
    .Q_N(_4318_),
    .Q(\collatz.iter[36] ));
 sg13g2_dfrbp_1 \iter[37]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net427),
    .D(_0101_),
    .Q_N(_4317_),
    .Q(\collatz.iter[37] ));
 sg13g2_dfrbp_1 \iter[38]$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net428),
    .D(_0102_),
    .Q_N(_4316_),
    .Q(\collatz.iter[38] ));
 sg13g2_dfrbp_1 \iter[39]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net429),
    .D(_0103_),
    .Q_N(_4315_),
    .Q(\collatz.iter[39] ));
 sg13g2_dfrbp_1 \iter[3]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net430),
    .D(_0104_),
    .Q_N(_4314_),
    .Q(\collatz.iter[3] ));
 sg13g2_dfrbp_1 \iter[40]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net431),
    .D(_0105_),
    .Q_N(_4313_),
    .Q(\collatz.iter[40] ));
 sg13g2_dfrbp_1 \iter[41]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net432),
    .D(_0106_),
    .Q_N(_4312_),
    .Q(\collatz.iter[41] ));
 sg13g2_dfrbp_1 \iter[42]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net433),
    .D(_0107_),
    .Q_N(_4311_),
    .Q(\collatz.iter[42] ));
 sg13g2_dfrbp_1 \iter[43]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net434),
    .D(_0108_),
    .Q_N(_4310_),
    .Q(\collatz.iter[43] ));
 sg13g2_dfrbp_1 \iter[44]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net435),
    .D(_0109_),
    .Q_N(_4309_),
    .Q(\collatz.iter[44] ));
 sg13g2_dfrbp_1 \iter[45]$_SDFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net436),
    .D(_0110_),
    .Q_N(_4308_),
    .Q(\collatz.iter[45] ));
 sg13g2_dfrbp_1 \iter[46]$_SDFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net437),
    .D(_0111_),
    .Q_N(_4307_),
    .Q(\collatz.iter[46] ));
 sg13g2_dfrbp_1 \iter[47]$_SDFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net438),
    .D(_0112_),
    .Q_N(_4306_),
    .Q(\collatz.iter[47] ));
 sg13g2_dfrbp_1 \iter[48]$_SDFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net439),
    .D(_0113_),
    .Q_N(_4305_),
    .Q(\collatz.iter[48] ));
 sg13g2_dfrbp_1 \iter[49]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net440),
    .D(_0114_),
    .Q_N(_4304_),
    .Q(\collatz.iter[49] ));
 sg13g2_dfrbp_1 \iter[4]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net441),
    .D(_0115_),
    .Q_N(_4303_),
    .Q(\collatz.iter[4] ));
 sg13g2_dfrbp_1 \iter[50]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net442),
    .D(_0116_),
    .Q_N(_4302_),
    .Q(\collatz.iter[50] ));
 sg13g2_dfrbp_1 \iter[51]$_SDFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net443),
    .D(_0117_),
    .Q_N(_4301_),
    .Q(\collatz.iter[51] ));
 sg13g2_dfrbp_1 \iter[52]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net444),
    .D(_0118_),
    .Q_N(_4300_),
    .Q(\collatz.iter[52] ));
 sg13g2_dfrbp_1 \iter[53]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net445),
    .D(_0119_),
    .Q_N(_4299_),
    .Q(\collatz.iter[53] ));
 sg13g2_dfrbp_1 \iter[54]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net446),
    .D(_0120_),
    .Q_N(_4298_),
    .Q(\collatz.iter[54] ));
 sg13g2_dfrbp_1 \iter[55]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net447),
    .D(_0121_),
    .Q_N(_4297_),
    .Q(\collatz.iter[55] ));
 sg13g2_dfrbp_1 \iter[56]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net448),
    .D(_0122_),
    .Q_N(_4296_),
    .Q(\collatz.iter[56] ));
 sg13g2_dfrbp_1 \iter[57]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net449),
    .D(_0123_),
    .Q_N(_4295_),
    .Q(\collatz.iter[57] ));
 sg13g2_dfrbp_1 \iter[58]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net450),
    .D(_0124_),
    .Q_N(_4294_),
    .Q(\collatz.iter[58] ));
 sg13g2_dfrbp_1 \iter[59]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net451),
    .D(_0125_),
    .Q_N(_4293_),
    .Q(\collatz.iter[59] ));
 sg13g2_dfrbp_1 \iter[5]$_SDFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net452),
    .D(_0126_),
    .Q_N(_4292_),
    .Q(\collatz.iter[5] ));
 sg13g2_dfrbp_1 \iter[60]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net453),
    .D(_0127_),
    .Q_N(_4291_),
    .Q(\collatz.iter[60] ));
 sg13g2_dfrbp_1 \iter[61]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net454),
    .D(_0128_),
    .Q_N(_4290_),
    .Q(\collatz.iter[61] ));
 sg13g2_dfrbp_1 \iter[62]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net455),
    .D(_0129_),
    .Q_N(_4289_),
    .Q(\collatz.iter[62] ));
 sg13g2_dfrbp_1 \iter[63]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net456),
    .D(_0130_),
    .Q_N(_4288_),
    .Q(\collatz.iter[63] ));
 sg13g2_dfrbp_1 \iter[64]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net457),
    .D(_0131_),
    .Q_N(_4287_),
    .Q(\collatz.iter[64] ));
 sg13g2_dfrbp_1 \iter[65]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net458),
    .D(_0132_),
    .Q_N(_4286_),
    .Q(\collatz.iter[65] ));
 sg13g2_dfrbp_1 \iter[66]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net459),
    .D(_0133_),
    .Q_N(_4285_),
    .Q(\collatz.iter[66] ));
 sg13g2_dfrbp_1 \iter[67]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net460),
    .D(_0134_),
    .Q_N(_4284_),
    .Q(\collatz.iter[67] ));
 sg13g2_dfrbp_1 \iter[68]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net461),
    .D(_0135_),
    .Q_N(_4283_),
    .Q(\collatz.iter[68] ));
 sg13g2_dfrbp_1 \iter[69]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net462),
    .D(_0136_),
    .Q_N(_4282_),
    .Q(\collatz.iter[69] ));
 sg13g2_dfrbp_1 \iter[6]$_SDFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net463),
    .D(_0137_),
    .Q_N(_4281_),
    .Q(\collatz.iter[6] ));
 sg13g2_dfrbp_1 \iter[70]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net464),
    .D(_0138_),
    .Q_N(_4280_),
    .Q(\collatz.iter[70] ));
 sg13g2_dfrbp_1 \iter[71]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net465),
    .D(_0139_),
    .Q_N(_4279_),
    .Q(\collatz.iter[71] ));
 sg13g2_dfrbp_1 \iter[72]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net466),
    .D(_0140_),
    .Q_N(_4278_),
    .Q(\collatz.iter[72] ));
 sg13g2_dfrbp_1 \iter[73]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net467),
    .D(_0141_),
    .Q_N(_4277_),
    .Q(\collatz.iter[73] ));
 sg13g2_dfrbp_1 \iter[74]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net468),
    .D(_0142_),
    .Q_N(_4276_),
    .Q(\collatz.iter[74] ));
 sg13g2_dfrbp_1 \iter[75]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net469),
    .D(_0143_),
    .Q_N(_4275_),
    .Q(\collatz.iter[75] ));
 sg13g2_dfrbp_1 \iter[76]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net470),
    .D(_0144_),
    .Q_N(_4274_),
    .Q(\collatz.iter[76] ));
 sg13g2_dfrbp_1 \iter[77]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net471),
    .D(_0145_),
    .Q_N(_4273_),
    .Q(\collatz.iter[77] ));
 sg13g2_dfrbp_1 \iter[78]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net472),
    .D(_0146_),
    .Q_N(_4272_),
    .Q(\collatz.iter[78] ));
 sg13g2_dfrbp_1 \iter[79]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net473),
    .D(_0147_),
    .Q_N(_4271_),
    .Q(\collatz.iter[79] ));
 sg13g2_dfrbp_1 \iter[7]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net474),
    .D(_0148_),
    .Q_N(_4270_),
    .Q(\collatz.iter[7] ));
 sg13g2_dfrbp_1 \iter[80]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net475),
    .D(_0149_),
    .Q_N(_4269_),
    .Q(\collatz.iter[80] ));
 sg13g2_dfrbp_1 \iter[81]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net476),
    .D(_0150_),
    .Q_N(_4268_),
    .Q(\collatz.iter[81] ));
 sg13g2_dfrbp_1 \iter[82]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net477),
    .D(_0151_),
    .Q_N(_4267_),
    .Q(\collatz.iter[82] ));
 sg13g2_dfrbp_1 \iter[83]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net478),
    .D(_0152_),
    .Q_N(_4266_),
    .Q(\collatz.iter[83] ));
 sg13g2_dfrbp_1 \iter[84]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net479),
    .D(_0153_),
    .Q_N(_4265_),
    .Q(\collatz.iter[84] ));
 sg13g2_dfrbp_1 \iter[85]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net480),
    .D(_0154_),
    .Q_N(_4264_),
    .Q(\collatz.iter[85] ));
 sg13g2_dfrbp_1 \iter[86]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net481),
    .D(_0155_),
    .Q_N(_4263_),
    .Q(\collatz.iter[86] ));
 sg13g2_dfrbp_1 \iter[87]$_SDFF_PN0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net482),
    .D(_0156_),
    .Q_N(_4262_),
    .Q(\collatz.iter[87] ));
 sg13g2_dfrbp_1 \iter[88]$_SDFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net483),
    .D(_0157_),
    .Q_N(_4261_),
    .Q(\collatz.iter[88] ));
 sg13g2_dfrbp_1 \iter[89]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net484),
    .D(_0158_),
    .Q_N(_4260_),
    .Q(\collatz.iter[89] ));
 sg13g2_dfrbp_1 \iter[8]$_SDFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net485),
    .D(_0159_),
    .Q_N(_4259_),
    .Q(\collatz.iter[8] ));
 sg13g2_dfrbp_1 \iter[90]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net486),
    .D(_0160_),
    .Q_N(_4258_),
    .Q(\collatz.iter[90] ));
 sg13g2_dfrbp_1 \iter[91]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net487),
    .D(_0161_),
    .Q_N(_4257_),
    .Q(\collatz.iter[91] ));
 sg13g2_dfrbp_1 \iter[92]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net488),
    .D(_0162_),
    .Q_N(_4256_),
    .Q(\collatz.iter[92] ));
 sg13g2_dfrbp_1 \iter[93]$_SDFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net489),
    .D(_0163_),
    .Q_N(_4255_),
    .Q(\collatz.iter[93] ));
 sg13g2_dfrbp_1 \iter[94]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net490),
    .D(_0164_),
    .Q_N(_4254_),
    .Q(\collatz.iter[94] ));
 sg13g2_dfrbp_1 \iter[95]$_SDFF_PN0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net491),
    .D(_0165_),
    .Q_N(_4253_),
    .Q(\collatz.iter[95] ));
 sg13g2_dfrbp_1 \iter[96]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net492),
    .D(_0166_),
    .Q_N(_4252_),
    .Q(\collatz.iter[96] ));
 sg13g2_dfrbp_1 \iter[97]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net493),
    .D(_0167_),
    .Q_N(_4251_),
    .Q(\collatz.iter[97] ));
 sg13g2_dfrbp_1 \iter[98]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net494),
    .D(_0168_),
    .Q_N(_4250_),
    .Q(\collatz.iter[98] ));
 sg13g2_dfrbp_1 \iter[99]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net495),
    .D(_0169_),
    .Q_N(_4249_),
    .Q(\collatz.iter[99] ));
 sg13g2_dfrbp_1 \iter[9]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net496),
    .D(_0170_),
    .Q_N(_4248_),
    .Q(\collatz.iter[9] ));
 sg13g2_dfrbp_1 \orbit_len[0]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net497),
    .D(_0171_),
    .Q_N(_4247_),
    .Q(\collatz.orbit_len[0] ));
 sg13g2_dfrbp_1 \orbit_len[10]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net498),
    .D(_0172_),
    .Q_N(_4246_),
    .Q(\collatz.orbit_len[10] ));
 sg13g2_dfrbp_1 \orbit_len[11]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net499),
    .D(_0173_),
    .Q_N(_4245_),
    .Q(\collatz.orbit_len[11] ));
 sg13g2_dfrbp_1 \orbit_len[12]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net500),
    .D(_0174_),
    .Q_N(_4244_),
    .Q(\collatz.orbit_len[12] ));
 sg13g2_dfrbp_1 \orbit_len[13]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net501),
    .D(_0175_),
    .Q_N(_4243_),
    .Q(\collatz.orbit_len[13] ));
 sg13g2_dfrbp_1 \orbit_len[14]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net502),
    .D(_0176_),
    .Q_N(_4242_),
    .Q(\collatz.orbit_len[14] ));
 sg13g2_dfrbp_1 \orbit_len[15]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net503),
    .D(_0177_),
    .Q_N(_4241_),
    .Q(\collatz.orbit_len[15] ));
 sg13g2_dfrbp_1 \orbit_len[1]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net504),
    .D(_0178_),
    .Q_N(_4240_),
    .Q(\collatz.orbit_len[1] ));
 sg13g2_dfrbp_1 \orbit_len[2]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net505),
    .D(_0179_),
    .Q_N(_4239_),
    .Q(\collatz.orbit_len[2] ));
 sg13g2_dfrbp_1 \orbit_len[3]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net506),
    .D(_0180_),
    .Q_N(_4238_),
    .Q(\collatz.orbit_len[3] ));
 sg13g2_dfrbp_1 \orbit_len[4]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net507),
    .D(_0181_),
    .Q_N(_4237_),
    .Q(\collatz.orbit_len[4] ));
 sg13g2_dfrbp_1 \orbit_len[5]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net508),
    .D(_0182_),
    .Q_N(_4236_),
    .Q(\collatz.orbit_len[5] ));
 sg13g2_dfrbp_1 \orbit_len[6]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net509),
    .D(_0183_),
    .Q_N(_4235_),
    .Q(\collatz.orbit_len[6] ));
 sg13g2_dfrbp_1 \orbit_len[7]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net510),
    .D(_0184_),
    .Q_N(_4234_),
    .Q(\collatz.orbit_len[7] ));
 sg13g2_dfrbp_1 \orbit_len[8]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net511),
    .D(_0185_),
    .Q_N(_4233_),
    .Q(\collatz.orbit_len[8] ));
 sg13g2_dfrbp_1 \orbit_len[9]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net512),
    .D(_0186_),
    .Q_N(_4232_),
    .Q(\collatz.orbit_len[9] ));
 sg13g2_dfrbp_1 \path_record_h16[0]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net513),
    .D(_0187_),
    .Q_N(_4231_),
    .Q(\collatz.path_record_h16[0] ));
 sg13g2_dfrbp_1 \path_record_h16[10]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net514),
    .D(_0188_),
    .Q_N(_4230_),
    .Q(\collatz.path_record_h16[10] ));
 sg13g2_dfrbp_1 \path_record_h16[11]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net515),
    .D(_0189_),
    .Q_N(_4229_),
    .Q(\collatz.path_record_h16[11] ));
 sg13g2_dfrbp_1 \path_record_h16[12]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net516),
    .D(_0190_),
    .Q_N(_0002_),
    .Q(\collatz.path_record_h16[12] ));
 sg13g2_dfrbp_1 \path_record_h16[13]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net517),
    .D(_0191_),
    .Q_N(_4228_),
    .Q(\collatz.path_record_h16[13] ));
 sg13g2_dfrbp_1 \path_record_h16[14]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net518),
    .D(_0192_),
    .Q_N(_4227_),
    .Q(\collatz.path_record_h16[14] ));
 sg13g2_dfrbp_1 \path_record_h16[15]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net519),
    .D(_0193_),
    .Q_N(_4226_),
    .Q(\collatz.path_record_h16[15] ));
 sg13g2_dfrbp_1 \path_record_h16[1]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net520),
    .D(_0194_),
    .Q_N(_4225_),
    .Q(\collatz.path_record_h16[1] ));
 sg13g2_dfrbp_1 \path_record_h16[2]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net521),
    .D(_0195_),
    .Q_N(_4224_),
    .Q(\collatz.path_record_h16[2] ));
 sg13g2_dfrbp_1 \path_record_h16[3]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net522),
    .D(_0196_),
    .Q_N(_4223_),
    .Q(\collatz.path_record_h16[3] ));
 sg13g2_dfrbp_1 \path_record_h16[4]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net523),
    .D(_0197_),
    .Q_N(_4222_),
    .Q(\collatz.path_record_h16[4] ));
 sg13g2_dfrbp_1 \path_record_h16[5]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net524),
    .D(_0198_),
    .Q_N(_4221_),
    .Q(\collatz.path_record_h16[5] ));
 sg13g2_dfrbp_1 \path_record_h16[6]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net525),
    .D(_0199_),
    .Q_N(_4220_),
    .Q(\collatz.path_record_h16[6] ));
 sg13g2_dfrbp_1 \path_record_h16[7]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net526),
    .D(_0200_),
    .Q_N(_4219_),
    .Q(\collatz.path_record_h16[7] ));
 sg13g2_dfrbp_1 \path_record_h16[8]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net527),
    .D(_0201_),
    .Q_N(_4218_),
    .Q(\collatz.path_record_h16[8] ));
 sg13g2_dfrbp_1 \path_record_h16[9]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net528),
    .D(_0202_),
    .Q_N(_4217_),
    .Q(\collatz.path_record_h16[9] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_oe[7]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_out[7]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[0]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[1]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[2]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[3]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[4]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[5]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[6]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[7]));
 sg13g2_buf_1 fanout13 (.A(_3656_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_3635_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_3631_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_3629_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_3607_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0700_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0396_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0392_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_3281_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_3215_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_3082_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_3053_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_2934_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_2894_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_2763_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_2729_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_2621_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_2470_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1960_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_1825_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1705_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1687_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1416_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1228_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1199_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0693_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0406_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_4046_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_4038_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_4034_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_3014_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_3008_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_2877_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_2859_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_2786_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_2714_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_2645_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_4047_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_4037_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_4033_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_3962_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_3232_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_2679_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_2628_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_2466_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_2367_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_2363_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_2084_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1896_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1657_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1552_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1198_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0405_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0389_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_4032_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_3969_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_3006_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_2988_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_2923_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_2871_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_2808_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_2724_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0706_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0704_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0404_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0400_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_4045_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_4039_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_4031_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_4027_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_3985_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_3863_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_3455_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_3317_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_3212_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_2807_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_2695_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_2465_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_2371_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_2080_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_1983_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_1326_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_0703_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0627_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_0620_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_0615_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_0403_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_0399_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_4116_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_4044_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_4030_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_4026_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_3994_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_3971_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_3967_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_3965_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_3958_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_3926_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_3917_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_3910_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_3862_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_3783_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_3761_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_3734_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_3073_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_2922_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_2455_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_2378_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_2318_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_2261_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_2232_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_2229_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_2128_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_2090_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_2058_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_2021_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_1955_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_1918_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_1913_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_1891_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_1787_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_1741_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_1722_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_1685_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_1674_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_1651_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_1536_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_1533_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_1417_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_1342_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_1319_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_1229_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_1225_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_0964_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_0950_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_0894_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_0717_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_0694_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_0678_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_0673_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_0669_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_0659_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_0634_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_0624_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_0604_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_0577_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_0574_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_0570_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_0552_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_0530_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_0528_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_0448_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_0432_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_0426_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_0418_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_0374_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_0370_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_0364_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_0355_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_0347_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_0345_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_0327_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_0318_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_0313_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_0303_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_0292_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_0284_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_0276_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_0237_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_0236_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_0220_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_0213_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_0210_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_4209_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_4176_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_4173_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_4170_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_4169_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_4165_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_4155_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_4154_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_4127_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_4120_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_4115_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_4106_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_4089_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_4050_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_4048_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_4043_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_4029_),
    .X(net202));
 sg13g2_buf_1 fanout203 (.A(_3970_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_3966_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_3950_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_3948_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_3946_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_3944_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_3941_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_3939_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_3937_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_3935_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_3932_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_3930_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_3928_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_3925_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_3921_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_3919_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_3916_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_3912_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_3909_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_3907_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_3902_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_3898_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_3886_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_3884_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_3874_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_3869_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_3867_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_3865_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_3843_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_3841_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_3839_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_3837_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_3815_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_3811_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_3809_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_3798_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_3796_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_3794_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_3792_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_3789_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_3787_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_3785_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_3782_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_3765_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_3763_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_3760_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_3758_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_3755_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_3752_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_3733_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_3731_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_3729_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_3727_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_3711_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_3709_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_3706_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_3704_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_3500_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_3481_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_1726_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_1655_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_1623_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_1487_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_0699_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_0249_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_0238_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_4097_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_4042_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_4016_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_4000_),
    .X(net272));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(_3997_));
 sg13g2_buf_2 fanout274 (.A(_3974_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_3931_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_3918_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_3911_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_3906_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_3904_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_3903_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_3870_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_3864_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_3860_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_3859_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_3850_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_3849_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_3846_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_3842_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_3840_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_3838_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_3825_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_3823_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_3821_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_3820_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_3784_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_3776_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_3771_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_3769_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_3767_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_3753_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_3744_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_3741_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_3740_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_3738_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_3737_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_3730_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_3728_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_3726_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_3724_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_3721_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_3720_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_3705_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_3703_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_3701_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_3700_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_3694_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_3693_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_3691_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_3690_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_3641_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_3447_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_3389_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_1745_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_1194_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_0707_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_0698_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_0382_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_4028_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_3980_),
    .X(net329));
 sg13g2_tielo _8589__330 (.L_LO(net330));
 sg13g2_tielo _8590__331 (.L_LO(net331));
 sg13g2_tielo _8591__332 (.L_LO(net332));
 sg13g2_tielo _8592__333 (.L_LO(net333));
 sg13g2_tielo _8593__334 (.L_LO(net334));
 sg13g2_tielo _8594__335 (.L_LO(net335));
 sg13g2_tielo _8595__336 (.L_LO(net336));
 sg13g2_tielo _8597__337 (.L_LO(net337));
 sg13g2_tielo _8598__338 (.L_LO(net338));
 sg13g2_tielo _8599__339 (.L_LO(net339));
 sg13g2_tielo _8600__340 (.L_LO(net340));
 sg13g2_tielo _8601__341 (.L_LO(net341));
 sg13g2_tielo _8602__342 (.L_LO(net342));
 sg13g2_tielo _8603__343 (.L_LO(net343));
 sg13g2_tiehi \data_out[0]$_SDFFE_PN0P__345  (.L_HI(net345));
 sg13g2_tiehi \data_out[1]$_SDFFE_PN0P__346  (.L_HI(net346));
 sg13g2_tiehi \data_out[2]$_SDFFE_PN0P__347  (.L_HI(net347));
 sg13g2_tiehi \data_out[3]$_SDFFE_PN0P__348  (.L_HI(net348));
 sg13g2_tiehi \data_out[4]$_SDFFE_PN0P__349  (.L_HI(net349));
 sg13g2_tiehi \data_out[5]$_SDFFE_PN0P__350  (.L_HI(net350));
 sg13g2_tiehi \data_out[6]$_SDFFE_PN0P__351  (.L_HI(net351));
 sg13g2_tiehi \data_out[7]$_SDFFE_PN0P__352  (.L_HI(net352));
 sg13g2_tiehi \ioctl[7]$_SDFFE_PP0P__353  (.L_HI(net353));
 sg13g2_tiehi \iter[0]$_SDFF_PN0__354  (.L_HI(net354));
 sg13g2_tiehi \iter[100]$_SDFF_PN0__355  (.L_HI(net355));
 sg13g2_tiehi \iter[101]$_SDFF_PN0__356  (.L_HI(net356));
 sg13g2_tiehi \iter[102]$_SDFF_PN0__357  (.L_HI(net357));
 sg13g2_tiehi \iter[103]$_SDFF_PN0__358  (.L_HI(net358));
 sg13g2_tiehi \iter[104]$_SDFF_PN0__359  (.L_HI(net359));
 sg13g2_tiehi \iter[105]$_SDFF_PN0__360  (.L_HI(net360));
 sg13g2_tiehi \iter[106]$_SDFF_PN0__361  (.L_HI(net361));
 sg13g2_tiehi \iter[107]$_SDFF_PN0__362  (.L_HI(net362));
 sg13g2_tiehi \iter[108]$_SDFF_PN0__363  (.L_HI(net363));
 sg13g2_tiehi \iter[109]$_SDFF_PN0__364  (.L_HI(net364));
 sg13g2_tiehi \iter[10]$_SDFF_PN0__365  (.L_HI(net365));
 sg13g2_tiehi \iter[110]$_SDFF_PN0__366  (.L_HI(net366));
 sg13g2_tiehi \iter[111]$_SDFF_PN0__367  (.L_HI(net367));
 sg13g2_tiehi \iter[112]$_SDFF_PN0__368  (.L_HI(net368));
 sg13g2_tiehi \iter[113]$_SDFF_PN0__369  (.L_HI(net369));
 sg13g2_tiehi \iter[114]$_SDFF_PN0__370  (.L_HI(net370));
 sg13g2_tiehi \iter[115]$_SDFF_PN0__371  (.L_HI(net371));
 sg13g2_tiehi \iter[116]$_SDFF_PN0__372  (.L_HI(net372));
 sg13g2_tiehi \iter[117]$_SDFF_PN0__373  (.L_HI(net373));
 sg13g2_tiehi \iter[118]$_SDFF_PN0__374  (.L_HI(net374));
 sg13g2_tiehi \iter[119]$_SDFF_PN0__375  (.L_HI(net375));
 sg13g2_tiehi \iter[11]$_SDFF_PN0__376  (.L_HI(net376));
 sg13g2_tiehi \iter[120]$_SDFF_PN0__377  (.L_HI(net377));
 sg13g2_tiehi \iter[121]$_SDFF_PN0__378  (.L_HI(net378));
 sg13g2_tiehi \iter[122]$_SDFF_PN0__379  (.L_HI(net379));
 sg13g2_tiehi \iter[123]$_SDFF_PN0__380  (.L_HI(net380));
 sg13g2_tiehi \iter[124]$_SDFF_PN0__381  (.L_HI(net381));
 sg13g2_tiehi \iter[125]$_SDFF_PN0__382  (.L_HI(net382));
 sg13g2_tiehi \iter[126]$_SDFF_PN0__383  (.L_HI(net383));
 sg13g2_tiehi \iter[127]$_SDFF_PN0__384  (.L_HI(net384));
 sg13g2_tiehi \iter[128]$_SDFF_PN0__385  (.L_HI(net385));
 sg13g2_tiehi \iter[129]$_SDFF_PN0__386  (.L_HI(net386));
 sg13g2_tiehi \iter[12]$_SDFF_PN0__387  (.L_HI(net387));
 sg13g2_tiehi \iter[130]$_SDFF_PN0__388  (.L_HI(net388));
 sg13g2_tiehi \iter[131]$_SDFF_PN0__389  (.L_HI(net389));
 sg13g2_tiehi \iter[132]$_SDFF_PN0__390  (.L_HI(net390));
 sg13g2_tiehi \iter[133]$_SDFF_PN0__391  (.L_HI(net391));
 sg13g2_tiehi \iter[134]$_SDFF_PN0__392  (.L_HI(net392));
 sg13g2_tiehi \iter[135]$_SDFF_PN0__393  (.L_HI(net393));
 sg13g2_tiehi \iter[136]$_SDFF_PN0__394  (.L_HI(net394));
 sg13g2_tiehi \iter[137]$_SDFF_PN0__395  (.L_HI(net395));
 sg13g2_tiehi \iter[138]$_SDFF_PN0__396  (.L_HI(net396));
 sg13g2_tiehi \iter[139]$_SDFF_PN0__397  (.L_HI(net397));
 sg13g2_tiehi \iter[13]$_SDFF_PN0__398  (.L_HI(net398));
 sg13g2_tiehi \iter[140]$_SDFF_PN0__399  (.L_HI(net399));
 sg13g2_tiehi \iter[141]$_SDFF_PN0__400  (.L_HI(net400));
 sg13g2_tiehi \iter[142]$_SDFF_PN0__401  (.L_HI(net401));
 sg13g2_tiehi \iter[143]$_SDFF_PN0__402  (.L_HI(net402));
 sg13g2_tiehi \iter[14]$_SDFF_PN0__403  (.L_HI(net403));
 sg13g2_tiehi \iter[15]$_SDFF_PN0__404  (.L_HI(net404));
 sg13g2_tiehi \iter[16]$_SDFF_PN0__405  (.L_HI(net405));
 sg13g2_tiehi \iter[17]$_SDFF_PN0__406  (.L_HI(net406));
 sg13g2_tiehi \iter[18]$_SDFF_PN0__407  (.L_HI(net407));
 sg13g2_tiehi \iter[19]$_SDFF_PN0__408  (.L_HI(net408));
 sg13g2_tiehi \iter[20]$_SDFF_PN0__409  (.L_HI(net409));
 sg13g2_tiehi \iter[21]$_SDFF_PN0__410  (.L_HI(net410));
 sg13g2_tiehi \iter[22]$_SDFF_PN0__411  (.L_HI(net411));
 sg13g2_tiehi \iter[23]$_SDFF_PN0__412  (.L_HI(net412));
 sg13g2_tiehi \iter[24]$_SDFF_PN0__413  (.L_HI(net413));
 sg13g2_tiehi \iter[25]$_SDFF_PN0__414  (.L_HI(net414));
 sg13g2_tiehi \iter[26]$_SDFF_PN0__415  (.L_HI(net415));
 sg13g2_tiehi \iter[27]$_SDFF_PN0__416  (.L_HI(net416));
 sg13g2_tiehi \iter[28]$_SDFF_PN0__417  (.L_HI(net417));
 sg13g2_tiehi \iter[29]$_SDFF_PN0__418  (.L_HI(net418));
 sg13g2_tiehi \iter[2]$_SDFF_PN0__419  (.L_HI(net419));
 sg13g2_tiehi \iter[30]$_SDFF_PN0__420  (.L_HI(net420));
 sg13g2_tiehi \iter[31]$_SDFF_PN0__421  (.L_HI(net421));
 sg13g2_tiehi \iter[32]$_SDFF_PN0__422  (.L_HI(net422));
 sg13g2_tiehi \iter[33]$_SDFF_PN0__423  (.L_HI(net423));
 sg13g2_tiehi \iter[34]$_SDFF_PN0__424  (.L_HI(net424));
 sg13g2_tiehi \iter[35]$_SDFF_PN0__425  (.L_HI(net425));
 sg13g2_tiehi \iter[36]$_SDFF_PN0__426  (.L_HI(net426));
 sg13g2_tiehi \iter[37]$_SDFF_PN0__427  (.L_HI(net427));
 sg13g2_tiehi \iter[38]$_SDFF_PN0__428  (.L_HI(net428));
 sg13g2_tiehi \iter[39]$_SDFF_PN0__429  (.L_HI(net429));
 sg13g2_tiehi \iter[3]$_SDFF_PN0__430  (.L_HI(net430));
 sg13g2_tiehi \iter[40]$_SDFF_PN0__431  (.L_HI(net431));
 sg13g2_tiehi \iter[41]$_SDFF_PN0__432  (.L_HI(net432));
 sg13g2_tiehi \iter[42]$_SDFF_PN0__433  (.L_HI(net433));
 sg13g2_tiehi \iter[43]$_SDFF_PN0__434  (.L_HI(net434));
 sg13g2_tiehi \iter[44]$_SDFF_PN0__435  (.L_HI(net435));
 sg13g2_tiehi \iter[45]$_SDFF_PN0__436  (.L_HI(net436));
 sg13g2_tiehi \iter[46]$_SDFF_PN0__437  (.L_HI(net437));
 sg13g2_tiehi \iter[47]$_SDFF_PN0__438  (.L_HI(net438));
 sg13g2_tiehi \iter[48]$_SDFF_PN0__439  (.L_HI(net439));
 sg13g2_tiehi \iter[49]$_SDFF_PN0__440  (.L_HI(net440));
 sg13g2_tiehi \iter[4]$_SDFF_PN0__441  (.L_HI(net441));
 sg13g2_tiehi \iter[50]$_SDFF_PN0__442  (.L_HI(net442));
 sg13g2_tiehi \iter[51]$_SDFF_PN0__443  (.L_HI(net443));
 sg13g2_tiehi \iter[52]$_SDFF_PN0__444  (.L_HI(net444));
 sg13g2_tiehi \iter[53]$_SDFF_PN0__445  (.L_HI(net445));
 sg13g2_tiehi \iter[54]$_SDFF_PN0__446  (.L_HI(net446));
 sg13g2_tiehi \iter[55]$_SDFF_PN0__447  (.L_HI(net447));
 sg13g2_tiehi \iter[56]$_SDFF_PN0__448  (.L_HI(net448));
 sg13g2_tiehi \iter[57]$_SDFF_PN0__449  (.L_HI(net449));
 sg13g2_tiehi \iter[58]$_SDFF_PN0__450  (.L_HI(net450));
 sg13g2_tiehi \iter[59]$_SDFF_PN0__451  (.L_HI(net451));
 sg13g2_tiehi \iter[5]$_SDFF_PN0__452  (.L_HI(net452));
 sg13g2_tiehi \iter[60]$_SDFF_PN0__453  (.L_HI(net453));
 sg13g2_tiehi \iter[61]$_SDFF_PN0__454  (.L_HI(net454));
 sg13g2_tiehi \iter[62]$_SDFF_PN0__455  (.L_HI(net455));
 sg13g2_tiehi \iter[63]$_SDFF_PN0__456  (.L_HI(net456));
 sg13g2_tiehi \iter[64]$_SDFF_PN0__457  (.L_HI(net457));
 sg13g2_tiehi \iter[65]$_SDFF_PN0__458  (.L_HI(net458));
 sg13g2_tiehi \iter[66]$_SDFF_PN0__459  (.L_HI(net459));
 sg13g2_tiehi \iter[67]$_SDFF_PN0__460  (.L_HI(net460));
 sg13g2_tiehi \iter[68]$_SDFF_PN0__461  (.L_HI(net461));
 sg13g2_tiehi \iter[69]$_SDFF_PN0__462  (.L_HI(net462));
 sg13g2_tiehi \iter[6]$_SDFF_PN0__463  (.L_HI(net463));
 sg13g2_tiehi \iter[70]$_SDFF_PN0__464  (.L_HI(net464));
 sg13g2_tiehi \iter[71]$_SDFF_PN0__465  (.L_HI(net465));
 sg13g2_tiehi \iter[72]$_SDFF_PN0__466  (.L_HI(net466));
 sg13g2_tiehi \iter[73]$_SDFF_PN0__467  (.L_HI(net467));
 sg13g2_tiehi \iter[74]$_SDFF_PN0__468  (.L_HI(net468));
 sg13g2_tiehi \iter[75]$_SDFF_PN0__469  (.L_HI(net469));
 sg13g2_tiehi \iter[76]$_SDFF_PN0__470  (.L_HI(net470));
 sg13g2_tiehi \iter[77]$_SDFF_PN0__471  (.L_HI(net471));
 sg13g2_tiehi \iter[78]$_SDFF_PN0__472  (.L_HI(net472));
 sg13g2_tiehi \iter[79]$_SDFF_PN0__473  (.L_HI(net473));
 sg13g2_tiehi \iter[7]$_SDFF_PN0__474  (.L_HI(net474));
 sg13g2_tiehi \iter[80]$_SDFF_PN0__475  (.L_HI(net475));
 sg13g2_tiehi \iter[81]$_SDFF_PN0__476  (.L_HI(net476));
 sg13g2_tiehi \iter[82]$_SDFF_PN0__477  (.L_HI(net477));
 sg13g2_tiehi \iter[83]$_SDFF_PN0__478  (.L_HI(net478));
 sg13g2_tiehi \iter[84]$_SDFF_PN0__479  (.L_HI(net479));
 sg13g2_tiehi \iter[85]$_SDFF_PN0__480  (.L_HI(net480));
 sg13g2_tiehi \iter[86]$_SDFF_PN0__481  (.L_HI(net481));
 sg13g2_tiehi \iter[87]$_SDFF_PN0__482  (.L_HI(net482));
 sg13g2_tiehi \iter[88]$_SDFF_PN0__483  (.L_HI(net483));
 sg13g2_tiehi \iter[89]$_SDFF_PN0__484  (.L_HI(net484));
 sg13g2_tiehi \iter[8]$_SDFF_PN0__485  (.L_HI(net485));
 sg13g2_tiehi \iter[90]$_SDFF_PN0__486  (.L_HI(net486));
 sg13g2_tiehi \iter[91]$_SDFF_PN0__487  (.L_HI(net487));
 sg13g2_tiehi \iter[92]$_SDFF_PN0__488  (.L_HI(net488));
 sg13g2_tiehi \iter[93]$_SDFF_PN0__489  (.L_HI(net489));
 sg13g2_tiehi \iter[94]$_SDFF_PN0__490  (.L_HI(net490));
 sg13g2_tiehi \iter[95]$_SDFF_PN0__491  (.L_HI(net491));
 sg13g2_tiehi \iter[96]$_SDFF_PN0__492  (.L_HI(net492));
 sg13g2_tiehi \iter[97]$_SDFF_PN0__493  (.L_HI(net493));
 sg13g2_tiehi \iter[98]$_SDFF_PN0__494  (.L_HI(net494));
 sg13g2_tiehi \iter[99]$_SDFF_PN0__495  (.L_HI(net495));
 sg13g2_tiehi \iter[9]$_SDFF_PN0__496  (.L_HI(net496));
 sg13g2_tiehi \orbit_len[0]$_SDFFE_PN0P__497  (.L_HI(net497));
 sg13g2_tiehi \orbit_len[10]$_SDFFE_PN0P__498  (.L_HI(net498));
 sg13g2_tiehi \orbit_len[11]$_SDFFE_PN0P__499  (.L_HI(net499));
 sg13g2_tiehi \orbit_len[12]$_SDFFE_PN0P__500  (.L_HI(net500));
 sg13g2_tiehi \orbit_len[13]$_SDFFE_PN0P__501  (.L_HI(net501));
 sg13g2_tiehi \orbit_len[14]$_SDFFE_PN0P__502  (.L_HI(net502));
 sg13g2_tiehi \orbit_len[15]$_SDFFE_PN0P__503  (.L_HI(net503));
 sg13g2_tiehi \orbit_len[1]$_SDFFE_PN0P__504  (.L_HI(net504));
 sg13g2_tiehi \orbit_len[2]$_SDFFE_PN0P__505  (.L_HI(net505));
 sg13g2_tiehi \orbit_len[3]$_SDFFE_PN0P__506  (.L_HI(net506));
 sg13g2_tiehi \orbit_len[4]$_SDFFE_PN0P__507  (.L_HI(net507));
 sg13g2_tiehi \orbit_len[5]$_SDFFE_PN0P__508  (.L_HI(net508));
 sg13g2_tiehi \orbit_len[6]$_SDFFE_PN0P__509  (.L_HI(net509));
 sg13g2_tiehi \orbit_len[7]$_SDFFE_PN0P__510  (.L_HI(net510));
 sg13g2_tiehi \orbit_len[8]$_SDFFE_PN0P__511  (.L_HI(net511));
 sg13g2_tiehi \orbit_len[9]$_SDFFE_PN0P__512  (.L_HI(net512));
 sg13g2_tiehi \path_record_h16[0]$_SDFFE_PN0P__513  (.L_HI(net513));
 sg13g2_tiehi \path_record_h16[10]$_SDFFE_PN0P__514  (.L_HI(net514));
 sg13g2_tiehi \path_record_h16[11]$_SDFFE_PN0P__515  (.L_HI(net515));
 sg13g2_tiehi \path_record_h16[12]$_SDFFE_PN0P__516  (.L_HI(net516));
 sg13g2_tiehi \path_record_h16[13]$_SDFFE_PN0P__517  (.L_HI(net517));
 sg13g2_tiehi \path_record_h16[14]$_SDFFE_PN0P__518  (.L_HI(net518));
 sg13g2_tiehi \path_record_h16[15]$_SDFFE_PN0P__519  (.L_HI(net519));
 sg13g2_tiehi \path_record_h16[1]$_SDFFE_PN0P__520  (.L_HI(net520));
 sg13g2_tiehi \path_record_h16[2]$_SDFFE_PN0P__521  (.L_HI(net521));
 sg13g2_tiehi \path_record_h16[3]$_SDFFE_PN0P__522  (.L_HI(net522));
 sg13g2_tiehi \path_record_h16[4]$_SDFFE_PN0P__523  (.L_HI(net523));
 sg13g2_tiehi \path_record_h16[5]$_SDFFE_PN0P__524  (.L_HI(net524));
 sg13g2_tiehi \path_record_h16[6]$_SDFFE_PN0P__525  (.L_HI(net525));
 sg13g2_tiehi \path_record_h16[7]$_SDFFE_PN0P__526  (.L_HI(net526));
 sg13g2_tiehi \path_record_h16[8]$_SDFFE_PN0P__527  (.L_HI(net527));
 sg13g2_tiehi \path_record_h16[9]$_SDFFE_PN0P__528  (.L_HI(net528));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_31__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0143_));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(_0143_));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_antennanp ANTENNA_6 (.A(clk));
 sg13g2_antennanp ANTENNA_7 (.A(_0143_));
 sg13g2_antennanp ANTENNA_8 (.A(clk));
 sg13g2_antennanp ANTENNA_9 (.A(clk));
 sg13g2_antennanp ANTENNA_10 (.A(_0143_));
 sg13g2_antennanp ANTENNA_11 (.A(clk));
 sg13g2_antennanp ANTENNA_12 (.A(clk));
 sg13g2_antennanp ANTENNA_13 (.A(clk));
 sg13g2_antennanp ANTENNA_14 (.A(_0143_));
 sg13g2_antennanp ANTENNA_15 (.A(clk));
 sg13g2_antennanp ANTENNA_16 (.A(clk));
 sg13g2_antennanp ANTENNA_17 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_4 FILLER_0_7 ();
 sg13g2_fill_1 FILLER_0_11 ();
 sg13g2_fill_1 FILLER_0_16 ();
 sg13g2_fill_1 FILLER_0_43 ();
 sg13g2_fill_1 FILLER_0_52 ();
 sg13g2_fill_2 FILLER_0_83 ();
 sg13g2_fill_1 FILLER_0_85 ();
 sg13g2_fill_2 FILLER_0_116 ();
 sg13g2_fill_2 FILLER_0_200 ();
 sg13g2_fill_2 FILLER_0_228 ();
 sg13g2_fill_1 FILLER_0_260 ();
 sg13g2_fill_2 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_423 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_33 ();
 sg13g2_fill_2 FILLER_1_39 ();
 sg13g2_fill_2 FILLER_1_67 ();
 sg13g2_fill_1 FILLER_1_69 ();
 sg13g2_decap_4 FILLER_1_74 ();
 sg13g2_fill_1 FILLER_1_78 ();
 sg13g2_fill_2 FILLER_1_92 ();
 sg13g2_decap_4 FILLER_1_107 ();
 sg13g2_fill_1 FILLER_1_111 ();
 sg13g2_fill_1 FILLER_1_125 ();
 sg13g2_fill_2 FILLER_1_130 ();
 sg13g2_fill_2 FILLER_1_158 ();
 sg13g2_fill_2 FILLER_1_173 ();
 sg13g2_fill_1 FILLER_1_175 ();
 sg13g2_fill_2 FILLER_1_180 ();
 sg13g2_fill_1 FILLER_1_208 ();
 sg13g2_fill_1 FILLER_1_217 ();
 sg13g2_decap_4 FILLER_1_222 ();
 sg13g2_fill_2 FILLER_1_265 ();
 sg13g2_decap_8 FILLER_1_274 ();
 sg13g2_decap_4 FILLER_1_281 ();
 sg13g2_fill_1 FILLER_1_315 ();
 sg13g2_fill_1 FILLER_1_329 ();
 sg13g2_fill_2 FILLER_1_343 ();
 sg13g2_fill_1 FILLER_1_350 ();
 sg13g2_fill_1 FILLER_1_355 ();
 sg13g2_fill_1 FILLER_1_360 ();
 sg13g2_fill_1 FILLER_1_365 ();
 sg13g2_fill_2 FILLER_1_374 ();
 sg13g2_fill_1 FILLER_1_380 ();
 sg13g2_fill_1 FILLER_1_385 ();
 sg13g2_fill_2 FILLER_1_389 ();
 sg13g2_fill_2 FILLER_1_395 ();
 sg13g2_fill_2 FILLER_1_401 ();
 sg13g2_fill_1 FILLER_1_403 ();
 sg13g2_decap_8 FILLER_1_408 ();
 sg13g2_fill_2 FILLER_1_415 ();
 sg13g2_fill_1 FILLER_1_417 ();
 sg13g2_decap_8 FILLER_1_423 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_fill_2 FILLER_2_18 ();
 sg13g2_fill_1 FILLER_2_20 ();
 sg13g2_fill_1 FILLER_2_26 ();
 sg13g2_fill_1 FILLER_2_31 ();
 sg13g2_fill_1 FILLER_2_36 ();
 sg13g2_fill_2 FILLER_2_63 ();
 sg13g2_fill_1 FILLER_2_91 ();
 sg13g2_fill_1 FILLER_2_131 ();
 sg13g2_fill_2 FILLER_2_136 ();
 sg13g2_fill_2 FILLER_2_184 ();
 sg13g2_decap_4 FILLER_2_190 ();
 sg13g2_fill_2 FILLER_2_194 ();
 sg13g2_fill_2 FILLER_2_200 ();
 sg13g2_fill_1 FILLER_2_236 ();
 sg13g2_fill_1 FILLER_2_245 ();
 sg13g2_fill_2 FILLER_2_289 ();
 sg13g2_fill_2 FILLER_2_295 ();
 sg13g2_fill_1 FILLER_2_297 ();
 sg13g2_decap_4 FILLER_2_302 ();
 sg13g2_fill_2 FILLER_2_306 ();
 sg13g2_fill_2 FILLER_2_313 ();
 sg13g2_fill_2 FILLER_2_324 ();
 sg13g2_fill_1 FILLER_2_326 ();
 sg13g2_fill_1 FILLER_2_377 ();
 sg13g2_fill_2 FILLER_2_383 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_7 ();
 sg13g2_fill_1 FILLER_3_9 ();
 sg13g2_fill_1 FILLER_3_31 ();
 sg13g2_fill_1 FILLER_3_42 ();
 sg13g2_fill_1 FILLER_3_47 ();
 sg13g2_fill_1 FILLER_3_57 ();
 sg13g2_fill_2 FILLER_3_62 ();
 sg13g2_fill_1 FILLER_3_64 ();
 sg13g2_fill_2 FILLER_3_78 ();
 sg13g2_fill_1 FILLER_3_80 ();
 sg13g2_decap_8 FILLER_3_85 ();
 sg13g2_decap_4 FILLER_3_96 ();
 sg13g2_fill_1 FILLER_3_100 ();
 sg13g2_decap_4 FILLER_3_105 ();
 sg13g2_fill_1 FILLER_3_109 ();
 sg13g2_fill_2 FILLER_3_114 ();
 sg13g2_fill_1 FILLER_3_124 ();
 sg13g2_fill_2 FILLER_3_156 ();
 sg13g2_fill_1 FILLER_3_163 ();
 sg13g2_fill_2 FILLER_3_168 ();
 sg13g2_fill_1 FILLER_3_174 ();
 sg13g2_fill_1 FILLER_3_189 ();
 sg13g2_fill_1 FILLER_3_199 ();
 sg13g2_fill_1 FILLER_3_205 ();
 sg13g2_fill_1 FILLER_3_210 ();
 sg13g2_fill_1 FILLER_3_215 ();
 sg13g2_fill_1 FILLER_3_220 ();
 sg13g2_fill_1 FILLER_3_226 ();
 sg13g2_fill_1 FILLER_3_236 ();
 sg13g2_fill_2 FILLER_3_289 ();
 sg13g2_fill_1 FILLER_3_321 ();
 sg13g2_fill_1 FILLER_3_370 ();
 sg13g2_fill_2 FILLER_3_376 ();
 sg13g2_fill_2 FILLER_3_383 ();
 sg13g2_fill_2 FILLER_3_389 ();
 sg13g2_fill_2 FILLER_3_396 ();
 sg13g2_fill_1 FILLER_3_398 ();
 sg13g2_fill_2 FILLER_3_403 ();
 sg13g2_decap_4 FILLER_3_409 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_4 FILLER_3_424 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_4 FILLER_4_7 ();
 sg13g2_fill_1 FILLER_4_11 ();
 sg13g2_fill_2 FILLER_4_43 ();
 sg13g2_fill_2 FILLER_4_51 ();
 sg13g2_fill_1 FILLER_4_53 ();
 sg13g2_fill_2 FILLER_4_59 ();
 sg13g2_fill_1 FILLER_4_65 ();
 sg13g2_fill_1 FILLER_4_92 ();
 sg13g2_fill_1 FILLER_4_129 ();
 sg13g2_fill_1 FILLER_4_136 ();
 sg13g2_fill_1 FILLER_4_151 ();
 sg13g2_fill_2 FILLER_4_173 ();
 sg13g2_fill_2 FILLER_4_195 ();
 sg13g2_fill_1 FILLER_4_202 ();
 sg13g2_fill_1 FILLER_4_219 ();
 sg13g2_fill_2 FILLER_4_224 ();
 sg13g2_fill_1 FILLER_4_243 ();
 sg13g2_fill_2 FILLER_4_249 ();
 sg13g2_fill_2 FILLER_4_255 ();
 sg13g2_fill_1 FILLER_4_257 ();
 sg13g2_fill_2 FILLER_4_263 ();
 sg13g2_fill_1 FILLER_4_265 ();
 sg13g2_fill_2 FILLER_4_270 ();
 sg13g2_fill_1 FILLER_4_327 ();
 sg13g2_fill_1 FILLER_4_333 ();
 sg13g2_fill_1 FILLER_4_339 ();
 sg13g2_fill_1 FILLER_4_349 ();
 sg13g2_fill_2 FILLER_4_375 ();
 sg13g2_fill_1 FILLER_4_391 ();
 sg13g2_fill_2 FILLER_4_418 ();
 sg13g2_fill_1 FILLER_4_420 ();
 sg13g2_decap_4 FILLER_4_425 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_fill_1 FILLER_5_55 ();
 sg13g2_fill_1 FILLER_5_136 ();
 sg13g2_fill_1 FILLER_5_147 ();
 sg13g2_fill_1 FILLER_5_166 ();
 sg13g2_fill_1 FILLER_5_177 ();
 sg13g2_fill_1 FILLER_5_182 ();
 sg13g2_fill_1 FILLER_5_246 ();
 sg13g2_fill_1 FILLER_5_251 ();
 sg13g2_fill_1 FILLER_5_257 ();
 sg13g2_fill_2 FILLER_5_263 ();
 sg13g2_fill_1 FILLER_5_269 ();
 sg13g2_fill_1 FILLER_5_275 ();
 sg13g2_fill_2 FILLER_5_314 ();
 sg13g2_fill_1 FILLER_5_316 ();
 sg13g2_fill_2 FILLER_5_338 ();
 sg13g2_fill_1 FILLER_5_364 ();
 sg13g2_fill_2 FILLER_5_391 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_7 ();
 sg13g2_fill_1 FILLER_6_12 ();
 sg13g2_fill_1 FILLER_6_19 ();
 sg13g2_fill_1 FILLER_6_25 ();
 sg13g2_fill_2 FILLER_6_30 ();
 sg13g2_fill_2 FILLER_6_53 ();
 sg13g2_fill_1 FILLER_6_55 ();
 sg13g2_fill_2 FILLER_6_65 ();
 sg13g2_fill_2 FILLER_6_91 ();
 sg13g2_fill_2 FILLER_6_131 ();
 sg13g2_fill_1 FILLER_6_147 ();
 sg13g2_fill_2 FILLER_6_177 ();
 sg13g2_fill_1 FILLER_6_201 ();
 sg13g2_fill_2 FILLER_6_213 ();
 sg13g2_fill_1 FILLER_6_219 ();
 sg13g2_fill_1 FILLER_6_225 ();
 sg13g2_fill_1 FILLER_6_235 ();
 sg13g2_fill_2 FILLER_6_267 ();
 sg13g2_fill_1 FILLER_6_269 ();
 sg13g2_decap_8 FILLER_6_275 ();
 sg13g2_fill_2 FILLER_6_296 ();
 sg13g2_fill_1 FILLER_6_298 ();
 sg13g2_fill_2 FILLER_6_340 ();
 sg13g2_fill_1 FILLER_6_347 ();
 sg13g2_fill_2 FILLER_6_356 ();
 sg13g2_fill_2 FILLER_6_363 ();
 sg13g2_fill_1 FILLER_6_377 ();
 sg13g2_fill_1 FILLER_6_383 ();
 sg13g2_fill_2 FILLER_6_401 ();
 sg13g2_fill_2 FILLER_6_421 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_fill_1 FILLER_7_40 ();
 sg13g2_fill_2 FILLER_7_63 ();
 sg13g2_fill_1 FILLER_7_65 ();
 sg13g2_fill_2 FILLER_7_105 ();
 sg13g2_fill_2 FILLER_7_128 ();
 sg13g2_fill_1 FILLER_7_130 ();
 sg13g2_fill_1 FILLER_7_152 ();
 sg13g2_fill_1 FILLER_7_166 ();
 sg13g2_fill_1 FILLER_7_208 ();
 sg13g2_fill_2 FILLER_7_218 ();
 sg13g2_fill_1 FILLER_7_225 ();
 sg13g2_decap_4 FILLER_7_253 ();
 sg13g2_fill_1 FILLER_7_257 ();
 sg13g2_fill_2 FILLER_7_264 ();
 sg13g2_fill_1 FILLER_7_266 ();
 sg13g2_fill_1 FILLER_7_275 ();
 sg13g2_fill_1 FILLER_7_297 ();
 sg13g2_fill_1 FILLER_7_311 ();
 sg13g2_fill_1 FILLER_7_328 ();
 sg13g2_fill_2 FILLER_7_372 ();
 sg13g2_fill_1 FILLER_7_383 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_47 ();
 sg13g2_decap_4 FILLER_8_54 ();
 sg13g2_fill_1 FILLER_8_87 ();
 sg13g2_fill_2 FILLER_8_114 ();
 sg13g2_fill_1 FILLER_8_116 ();
 sg13g2_fill_2 FILLER_8_121 ();
 sg13g2_fill_1 FILLER_8_123 ();
 sg13g2_fill_1 FILLER_8_208 ();
 sg13g2_fill_1 FILLER_8_213 ();
 sg13g2_fill_1 FILLER_8_218 ();
 sg13g2_fill_1 FILLER_8_231 ();
 sg13g2_fill_1 FILLER_8_294 ();
 sg13g2_fill_2 FILLER_8_300 ();
 sg13g2_fill_1 FILLER_8_307 ();
 sg13g2_fill_2 FILLER_8_314 ();
 sg13g2_fill_1 FILLER_8_322 ();
 sg13g2_fill_1 FILLER_8_328 ();
 sg13g2_fill_1 FILLER_8_338 ();
 sg13g2_fill_2 FILLER_8_351 ();
 sg13g2_fill_1 FILLER_8_361 ();
 sg13g2_fill_1 FILLER_8_367 ();
 sg13g2_fill_1 FILLER_8_372 ();
 sg13g2_fill_1 FILLER_8_378 ();
 sg13g2_fill_1 FILLER_8_393 ();
 sg13g2_fill_2 FILLER_8_414 ();
 sg13g2_fill_1 FILLER_8_416 ();
 sg13g2_decap_4 FILLER_8_425 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_fill_1 FILLER_9_34 ();
 sg13g2_fill_2 FILLER_9_40 ();
 sg13g2_fill_2 FILLER_9_68 ();
 sg13g2_fill_1 FILLER_9_103 ();
 sg13g2_decap_4 FILLER_9_112 ();
 sg13g2_fill_1 FILLER_9_126 ();
 sg13g2_decap_4 FILLER_9_134 ();
 sg13g2_decap_4 FILLER_9_142 ();
 sg13g2_fill_1 FILLER_9_146 ();
 sg13g2_fill_1 FILLER_9_153 ();
 sg13g2_fill_2 FILLER_9_187 ();
 sg13g2_fill_1 FILLER_9_189 ();
 sg13g2_fill_1 FILLER_9_200 ();
 sg13g2_fill_2 FILLER_9_223 ();
 sg13g2_fill_1 FILLER_9_225 ();
 sg13g2_fill_1 FILLER_9_234 ();
 sg13g2_fill_2 FILLER_9_245 ();
 sg13g2_fill_1 FILLER_9_247 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_fill_2 FILLER_9_259 ();
 sg13g2_fill_1 FILLER_9_261 ();
 sg13g2_fill_1 FILLER_9_266 ();
 sg13g2_fill_2 FILLER_9_311 ();
 sg13g2_fill_1 FILLER_9_313 ();
 sg13g2_fill_2 FILLER_9_320 ();
 sg13g2_fill_1 FILLER_9_342 ();
 sg13g2_fill_1 FILLER_9_347 ();
 sg13g2_fill_1 FILLER_9_370 ();
 sg13g2_fill_1 FILLER_9_399 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_fill_1 FILLER_9_415 ();
 sg13g2_decap_8 FILLER_9_421 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_2 ();
 sg13g2_fill_1 FILLER_10_8 ();
 sg13g2_fill_1 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_21 ();
 sg13g2_fill_1 FILLER_10_31 ();
 sg13g2_fill_2 FILLER_10_53 ();
 sg13g2_fill_1 FILLER_10_55 ();
 sg13g2_fill_2 FILLER_10_65 ();
 sg13g2_fill_1 FILLER_10_84 ();
 sg13g2_fill_2 FILLER_10_106 ();
 sg13g2_fill_2 FILLER_10_127 ();
 sg13g2_decap_4 FILLER_10_135 ();
 sg13g2_fill_2 FILLER_10_165 ();
 sg13g2_fill_1 FILLER_10_167 ();
 sg13g2_fill_1 FILLER_10_173 ();
 sg13g2_fill_2 FILLER_10_182 ();
 sg13g2_fill_2 FILLER_10_196 ();
 sg13g2_fill_1 FILLER_10_198 ();
 sg13g2_fill_1 FILLER_10_211 ();
 sg13g2_fill_1 FILLER_10_217 ();
 sg13g2_fill_1 FILLER_10_223 ();
 sg13g2_fill_1 FILLER_10_229 ();
 sg13g2_fill_1 FILLER_10_235 ();
 sg13g2_fill_2 FILLER_10_240 ();
 sg13g2_decap_4 FILLER_10_255 ();
 sg13g2_fill_1 FILLER_10_259 ();
 sg13g2_fill_1 FILLER_10_323 ();
 sg13g2_fill_1 FILLER_10_328 ();
 sg13g2_fill_1 FILLER_10_335 ();
 sg13g2_fill_1 FILLER_10_353 ();
 sg13g2_fill_1 FILLER_10_406 ();
 sg13g2_fill_2 FILLER_10_411 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_23 ();
 sg13g2_fill_1 FILLER_11_29 ();
 sg13g2_decap_4 FILLER_11_38 ();
 sg13g2_fill_2 FILLER_11_49 ();
 sg13g2_fill_2 FILLER_11_59 ();
 sg13g2_fill_1 FILLER_11_61 ();
 sg13g2_fill_1 FILLER_11_97 ();
 sg13g2_decap_8 FILLER_11_103 ();
 sg13g2_fill_1 FILLER_11_123 ();
 sg13g2_decap_8 FILLER_11_163 ();
 sg13g2_fill_1 FILLER_11_180 ();
 sg13g2_decap_4 FILLER_11_185 ();
 sg13g2_fill_1 FILLER_11_194 ();
 sg13g2_fill_1 FILLER_11_199 ();
 sg13g2_fill_1 FILLER_11_204 ();
 sg13g2_fill_1 FILLER_11_210 ();
 sg13g2_fill_2 FILLER_11_224 ();
 sg13g2_fill_1 FILLER_11_231 ();
 sg13g2_fill_1 FILLER_11_258 ();
 sg13g2_decap_4 FILLER_11_272 ();
 sg13g2_fill_2 FILLER_11_276 ();
 sg13g2_decap_4 FILLER_11_283 ();
 sg13g2_fill_1 FILLER_11_287 ();
 sg13g2_fill_2 FILLER_11_342 ();
 sg13g2_fill_1 FILLER_11_390 ();
 sg13g2_decap_4 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_12_31 ();
 sg13g2_fill_2 FILLER_12_46 ();
 sg13g2_fill_1 FILLER_12_48 ();
 sg13g2_fill_2 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_66 ();
 sg13g2_fill_1 FILLER_12_73 ();
 sg13g2_fill_1 FILLER_12_80 ();
 sg13g2_fill_1 FILLER_12_85 ();
 sg13g2_fill_2 FILLER_12_99 ();
 sg13g2_fill_1 FILLER_12_120 ();
 sg13g2_fill_2 FILLER_12_125 ();
 sg13g2_fill_1 FILLER_12_135 ();
 sg13g2_fill_2 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_fill_2 FILLER_12_154 ();
 sg13g2_fill_1 FILLER_12_156 ();
 sg13g2_fill_1 FILLER_12_195 ();
 sg13g2_fill_1 FILLER_12_206 ();
 sg13g2_fill_1 FILLER_12_212 ();
 sg13g2_fill_1 FILLER_12_218 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_fill_2 FILLER_12_271 ();
 sg13g2_fill_1 FILLER_12_301 ();
 sg13g2_fill_2 FILLER_12_342 ();
 sg13g2_fill_1 FILLER_12_344 ();
 sg13g2_fill_1 FILLER_12_355 ();
 sg13g2_fill_1 FILLER_12_360 ();
 sg13g2_fill_1 FILLER_12_367 ();
 sg13g2_fill_1 FILLER_12_373 ();
 sg13g2_fill_2 FILLER_12_379 ();
 sg13g2_fill_1 FILLER_12_385 ();
 sg13g2_fill_1 FILLER_12_392 ();
 sg13g2_fill_1 FILLER_12_397 ();
 sg13g2_fill_1 FILLER_12_402 ();
 sg13g2_fill_1 FILLER_12_415 ();
 sg13g2_decap_4 FILLER_12_421 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_11 ();
 sg13g2_fill_1 FILLER_13_13 ();
 sg13g2_decap_4 FILLER_13_20 ();
 sg13g2_fill_1 FILLER_13_40 ();
 sg13g2_fill_2 FILLER_13_60 ();
 sg13g2_decap_8 FILLER_13_66 ();
 sg13g2_fill_1 FILLER_13_73 ();
 sg13g2_fill_1 FILLER_13_114 ();
 sg13g2_fill_2 FILLER_13_121 ();
 sg13g2_fill_1 FILLER_13_123 ();
 sg13g2_fill_1 FILLER_13_129 ();
 sg13g2_decap_4 FILLER_13_146 ();
 sg13g2_fill_2 FILLER_13_154 ();
 sg13g2_fill_2 FILLER_13_161 ();
 sg13g2_fill_2 FILLER_13_168 ();
 sg13g2_fill_1 FILLER_13_170 ();
 sg13g2_decap_4 FILLER_13_174 ();
 sg13g2_decap_4 FILLER_13_183 ();
 sg13g2_fill_2 FILLER_13_193 ();
 sg13g2_fill_1 FILLER_13_195 ();
 sg13g2_fill_1 FILLER_13_223 ();
 sg13g2_fill_1 FILLER_13_230 ();
 sg13g2_fill_1 FILLER_13_238 ();
 sg13g2_fill_1 FILLER_13_265 ();
 sg13g2_fill_2 FILLER_13_278 ();
 sg13g2_fill_2 FILLER_13_285 ();
 sg13g2_fill_2 FILLER_13_292 ();
 sg13g2_fill_1 FILLER_13_294 ();
 sg13g2_fill_2 FILLER_13_306 ();
 sg13g2_fill_1 FILLER_13_308 ();
 sg13g2_fill_2 FILLER_13_324 ();
 sg13g2_fill_1 FILLER_13_350 ();
 sg13g2_fill_1 FILLER_13_356 ();
 sg13g2_fill_1 FILLER_13_389 ();
 sg13g2_fill_2 FILLER_13_421 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_decap_4 FILLER_14_16 ();
 sg13g2_fill_2 FILLER_14_34 ();
 sg13g2_fill_1 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_82 ();
 sg13g2_fill_1 FILLER_14_88 ();
 sg13g2_fill_1 FILLER_14_107 ();
 sg13g2_fill_2 FILLER_14_125 ();
 sg13g2_fill_2 FILLER_14_140 ();
 sg13g2_fill_2 FILLER_14_147 ();
 sg13g2_fill_1 FILLER_14_149 ();
 sg13g2_fill_1 FILLER_14_157 ();
 sg13g2_fill_2 FILLER_14_168 ();
 sg13g2_fill_1 FILLER_14_176 ();
 sg13g2_fill_1 FILLER_14_182 ();
 sg13g2_fill_1 FILLER_14_197 ();
 sg13g2_fill_1 FILLER_14_227 ();
 sg13g2_fill_2 FILLER_14_248 ();
 sg13g2_fill_2 FILLER_14_254 ();
 sg13g2_fill_2 FILLER_14_260 ();
 sg13g2_fill_1 FILLER_14_262 ();
 sg13g2_fill_1 FILLER_14_275 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_293 ();
 sg13g2_fill_2 FILLER_14_313 ();
 sg13g2_fill_2 FILLER_14_320 ();
 sg13g2_fill_1 FILLER_14_322 ();
 sg13g2_fill_1 FILLER_14_328 ();
 sg13g2_fill_2 FILLER_14_335 ();
 sg13g2_fill_1 FILLER_14_337 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_4 FILLER_14_357 ();
 sg13g2_fill_2 FILLER_14_373 ();
 sg13g2_fill_2 FILLER_14_405 ();
 sg13g2_fill_2 FILLER_14_416 ();
 sg13g2_fill_1 FILLER_14_418 ();
 sg13g2_fill_2 FILLER_14_428 ();
 sg13g2_fill_2 FILLER_15_30 ();
 sg13g2_decap_4 FILLER_15_46 ();
 sg13g2_fill_1 FILLER_15_50 ();
 sg13g2_fill_2 FILLER_15_63 ();
 sg13g2_fill_1 FILLER_15_70 ();
 sg13g2_fill_2 FILLER_15_79 ();
 sg13g2_fill_1 FILLER_15_91 ();
 sg13g2_decap_4 FILLER_15_97 ();
 sg13g2_fill_1 FILLER_15_101 ();
 sg13g2_fill_2 FILLER_15_106 ();
 sg13g2_fill_2 FILLER_15_113 ();
 sg13g2_decap_4 FILLER_15_143 ();
 sg13g2_fill_2 FILLER_15_161 ();
 sg13g2_fill_1 FILLER_15_163 ();
 sg13g2_decap_4 FILLER_15_168 ();
 sg13g2_fill_1 FILLER_15_172 ();
 sg13g2_fill_2 FILLER_15_191 ();
 sg13g2_fill_1 FILLER_15_193 ();
 sg13g2_decap_4 FILLER_15_234 ();
 sg13g2_decap_8 FILLER_15_251 ();
 sg13g2_decap_8 FILLER_15_258 ();
 sg13g2_fill_1 FILLER_15_269 ();
 sg13g2_fill_1 FILLER_15_274 ();
 sg13g2_fill_1 FILLER_15_280 ();
 sg13g2_fill_1 FILLER_15_286 ();
 sg13g2_fill_2 FILLER_15_309 ();
 sg13g2_fill_1 FILLER_15_337 ();
 sg13g2_fill_2 FILLER_15_352 ();
 sg13g2_fill_2 FILLER_15_385 ();
 sg13g2_fill_2 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_403 ();
 sg13g2_fill_1 FILLER_16_35 ();
 sg13g2_fill_1 FILLER_16_39 ();
 sg13g2_fill_1 FILLER_16_45 ();
 sg13g2_fill_1 FILLER_16_51 ();
 sg13g2_fill_2 FILLER_16_64 ();
 sg13g2_fill_2 FILLER_16_86 ();
 sg13g2_fill_1 FILLER_16_88 ();
 sg13g2_fill_2 FILLER_16_116 ();
 sg13g2_fill_2 FILLER_16_138 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_fill_2 FILLER_16_167 ();
 sg13g2_decap_4 FILLER_16_176 ();
 sg13g2_fill_2 FILLER_16_204 ();
 sg13g2_decap_4 FILLER_16_216 ();
 sg13g2_fill_1 FILLER_16_220 ();
 sg13g2_decap_4 FILLER_16_229 ();
 sg13g2_fill_1 FILLER_16_233 ();
 sg13g2_fill_1 FILLER_16_250 ();
 sg13g2_decap_8 FILLER_16_256 ();
 sg13g2_fill_2 FILLER_16_277 ();
 sg13g2_fill_1 FILLER_16_279 ();
 sg13g2_fill_2 FILLER_16_286 ();
 sg13g2_fill_2 FILLER_16_301 ();
 sg13g2_decap_4 FILLER_16_317 ();
 sg13g2_decap_4 FILLER_16_328 ();
 sg13g2_fill_2 FILLER_16_336 ();
 sg13g2_fill_1 FILLER_16_338 ();
 sg13g2_fill_2 FILLER_16_353 ();
 sg13g2_fill_1 FILLER_16_355 ();
 sg13g2_fill_2 FILLER_16_366 ();
 sg13g2_fill_1 FILLER_16_368 ();
 sg13g2_decap_4 FILLER_16_374 ();
 sg13g2_fill_1 FILLER_16_378 ();
 sg13g2_fill_1 FILLER_16_382 ();
 sg13g2_fill_2 FILLER_16_388 ();
 sg13g2_fill_2 FILLER_16_395 ();
 sg13g2_fill_2 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_18 ();
 sg13g2_fill_1 FILLER_17_49 ();
 sg13g2_fill_1 FILLER_17_54 ();
 sg13g2_fill_2 FILLER_17_76 ();
 sg13g2_fill_1 FILLER_17_78 ();
 sg13g2_fill_1 FILLER_17_95 ();
 sg13g2_fill_1 FILLER_17_114 ();
 sg13g2_fill_1 FILLER_17_120 ();
 sg13g2_fill_1 FILLER_17_126 ();
 sg13g2_fill_2 FILLER_17_131 ();
 sg13g2_fill_2 FILLER_17_141 ();
 sg13g2_fill_1 FILLER_17_156 ();
 sg13g2_fill_2 FILLER_17_161 ();
 sg13g2_fill_1 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_175 ();
 sg13g2_fill_2 FILLER_17_183 ();
 sg13g2_fill_1 FILLER_17_185 ();
 sg13g2_fill_1 FILLER_17_194 ();
 sg13g2_fill_2 FILLER_17_200 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_212 ();
 sg13g2_fill_1 FILLER_17_214 ();
 sg13g2_fill_1 FILLER_17_223 ();
 sg13g2_fill_1 FILLER_17_229 ();
 sg13g2_fill_1 FILLER_17_234 ();
 sg13g2_fill_2 FILLER_17_240 ();
 sg13g2_fill_2 FILLER_17_247 ();
 sg13g2_fill_1 FILLER_17_249 ();
 sg13g2_fill_2 FILLER_17_255 ();
 sg13g2_fill_1 FILLER_17_257 ();
 sg13g2_fill_1 FILLER_17_285 ();
 sg13g2_fill_1 FILLER_17_290 ();
 sg13g2_fill_1 FILLER_17_296 ();
 sg13g2_fill_1 FILLER_17_308 ();
 sg13g2_decap_4 FILLER_17_318 ();
 sg13g2_fill_1 FILLER_17_333 ();
 sg13g2_fill_1 FILLER_17_348 ();
 sg13g2_fill_2 FILLER_17_354 ();
 sg13g2_fill_1 FILLER_17_360 ();
 sg13g2_fill_1 FILLER_17_366 ();
 sg13g2_fill_1 FILLER_17_371 ();
 sg13g2_fill_1 FILLER_17_377 ();
 sg13g2_fill_2 FILLER_17_409 ();
 sg13g2_fill_1 FILLER_17_416 ();
 sg13g2_fill_2 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_6 ();
 sg13g2_fill_2 FILLER_18_20 ();
 sg13g2_fill_1 FILLER_18_22 ();
 sg13g2_fill_2 FILLER_18_55 ();
 sg13g2_fill_1 FILLER_18_62 ();
 sg13g2_fill_1 FILLER_18_66 ();
 sg13g2_fill_2 FILLER_18_80 ();
 sg13g2_fill_1 FILLER_18_82 ();
 sg13g2_fill_1 FILLER_18_88 ();
 sg13g2_fill_1 FILLER_18_94 ();
 sg13g2_fill_1 FILLER_18_100 ();
 sg13g2_fill_1 FILLER_18_107 ();
 sg13g2_fill_1 FILLER_18_114 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_137 ();
 sg13g2_fill_1 FILLER_18_144 ();
 sg13g2_fill_1 FILLER_18_156 ();
 sg13g2_decap_8 FILLER_18_162 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_fill_2 FILLER_18_179 ();
 sg13g2_fill_2 FILLER_18_185 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_1 FILLER_18_192 ();
 sg13g2_fill_2 FILLER_18_198 ();
 sg13g2_fill_1 FILLER_18_200 ();
 sg13g2_decap_4 FILLER_18_210 ();
 sg13g2_fill_2 FILLER_18_268 ();
 sg13g2_fill_1 FILLER_18_270 ();
 sg13g2_decap_4 FILLER_18_277 ();
 sg13g2_fill_1 FILLER_18_292 ();
 sg13g2_fill_1 FILLER_18_304 ();
 sg13g2_fill_2 FILLER_18_313 ();
 sg13g2_fill_2 FILLER_18_323 ();
 sg13g2_fill_1 FILLER_18_325 ();
 sg13g2_fill_2 FILLER_18_331 ();
 sg13g2_fill_2 FILLER_18_338 ();
 sg13g2_fill_1 FILLER_18_340 ();
 sg13g2_fill_1 FILLER_18_379 ();
 sg13g2_fill_2 FILLER_18_385 ();
 sg13g2_fill_1 FILLER_18_401 ();
 sg13g2_fill_2 FILLER_18_420 ();
 sg13g2_fill_1 FILLER_18_422 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_fill_1 FILLER_19_4 ();
 sg13g2_fill_1 FILLER_19_19 ();
 sg13g2_fill_1 FILLER_19_29 ();
 sg13g2_fill_1 FILLER_19_35 ();
 sg13g2_fill_1 FILLER_19_43 ();
 sg13g2_fill_1 FILLER_19_49 ();
 sg13g2_decap_4 FILLER_19_61 ();
 sg13g2_fill_2 FILLER_19_70 ();
 sg13g2_decap_4 FILLER_19_77 ();
 sg13g2_fill_2 FILLER_19_90 ();
 sg13g2_fill_1 FILLER_19_92 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_fill_1 FILLER_19_120 ();
 sg13g2_fill_2 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_128 ();
 sg13g2_fill_1 FILLER_19_147 ();
 sg13g2_fill_1 FILLER_19_158 ();
 sg13g2_fill_2 FILLER_19_192 ();
 sg13g2_decap_8 FILLER_19_199 ();
 sg13g2_decap_8 FILLER_19_215 ();
 sg13g2_decap_4 FILLER_19_222 ();
 sg13g2_fill_1 FILLER_19_226 ();
 sg13g2_fill_2 FILLER_19_252 ();
 sg13g2_fill_1 FILLER_19_254 ();
 sg13g2_fill_2 FILLER_19_265 ();
 sg13g2_fill_2 FILLER_19_276 ();
 sg13g2_fill_2 FILLER_19_284 ();
 sg13g2_fill_1 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_294 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_327 ();
 sg13g2_fill_2 FILLER_19_331 ();
 sg13g2_fill_2 FILLER_19_338 ();
 sg13g2_fill_2 FILLER_19_344 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_fill_2 FILLER_19_353 ();
 sg13g2_fill_1 FILLER_19_355 ();
 sg13g2_fill_1 FILLER_19_374 ();
 sg13g2_fill_2 FILLER_19_379 ();
 sg13g2_fill_1 FILLER_19_392 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_6 ();
 sg13g2_fill_2 FILLER_20_12 ();
 sg13g2_fill_1 FILLER_20_22 ();
 sg13g2_fill_2 FILLER_20_29 ();
 sg13g2_fill_1 FILLER_20_55 ();
 sg13g2_fill_1 FILLER_20_61 ();
 sg13g2_fill_1 FILLER_20_66 ();
 sg13g2_fill_1 FILLER_20_78 ();
 sg13g2_fill_1 FILLER_20_84 ();
 sg13g2_fill_1 FILLER_20_90 ();
 sg13g2_decap_4 FILLER_20_97 ();
 sg13g2_fill_1 FILLER_20_101 ();
 sg13g2_fill_1 FILLER_20_109 ();
 sg13g2_fill_2 FILLER_20_115 ();
 sg13g2_fill_1 FILLER_20_117 ();
 sg13g2_fill_1 FILLER_20_126 ();
 sg13g2_decap_4 FILLER_20_149 ();
 sg13g2_fill_1 FILLER_20_167 ();
 sg13g2_fill_2 FILLER_20_173 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_190 ();
 sg13g2_fill_2 FILLER_20_199 ();
 sg13g2_fill_1 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_222 ();
 sg13g2_fill_2 FILLER_20_248 ();
 sg13g2_fill_1 FILLER_20_250 ();
 sg13g2_fill_1 FILLER_20_256 ();
 sg13g2_fill_1 FILLER_20_261 ();
 sg13g2_fill_2 FILLER_20_279 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_decap_4 FILLER_20_292 ();
 sg13g2_fill_1 FILLER_20_304 ();
 sg13g2_fill_1 FILLER_20_311 ();
 sg13g2_fill_1 FILLER_20_318 ();
 sg13g2_fill_1 FILLER_20_327 ();
 sg13g2_fill_1 FILLER_20_333 ();
 sg13g2_fill_2 FILLER_20_338 ();
 sg13g2_fill_2 FILLER_20_359 ();
 sg13g2_fill_1 FILLER_20_361 ();
 sg13g2_fill_2 FILLER_20_391 ();
 sg13g2_fill_2 FILLER_20_408 ();
 sg13g2_fill_1 FILLER_20_424 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_10 ();
 sg13g2_fill_1 FILLER_21_16 ();
 sg13g2_fill_1 FILLER_21_21 ();
 sg13g2_fill_1 FILLER_21_34 ();
 sg13g2_fill_1 FILLER_21_39 ();
 sg13g2_fill_1 FILLER_21_45 ();
 sg13g2_fill_1 FILLER_21_51 ();
 sg13g2_decap_4 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_66 ();
 sg13g2_fill_1 FILLER_21_72 ();
 sg13g2_fill_1 FILLER_21_83 ();
 sg13g2_fill_2 FILLER_21_114 ();
 sg13g2_fill_2 FILLER_21_122 ();
 sg13g2_fill_1 FILLER_21_124 ();
 sg13g2_fill_1 FILLER_21_129 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_fill_1 FILLER_21_163 ();
 sg13g2_fill_1 FILLER_21_174 ();
 sg13g2_fill_1 FILLER_21_179 ();
 sg13g2_fill_2 FILLER_21_189 ();
 sg13g2_fill_1 FILLER_21_196 ();
 sg13g2_fill_1 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_209 ();
 sg13g2_fill_2 FILLER_21_219 ();
 sg13g2_fill_1 FILLER_21_221 ();
 sg13g2_fill_2 FILLER_21_236 ();
 sg13g2_fill_2 FILLER_21_260 ();
 sg13g2_fill_1 FILLER_21_266 ();
 sg13g2_fill_1 FILLER_21_272 ();
 sg13g2_fill_1 FILLER_21_297 ();
 sg13g2_fill_2 FILLER_21_307 ();
 sg13g2_fill_1 FILLER_21_314 ();
 sg13g2_decap_4 FILLER_21_331 ();
 sg13g2_fill_2 FILLER_21_348 ();
 sg13g2_fill_2 FILLER_21_368 ();
 sg13g2_fill_1 FILLER_21_370 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_32 ();
 sg13g2_fill_1 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_69 ();
 sg13g2_fill_2 FILLER_22_75 ();
 sg13g2_fill_2 FILLER_22_84 ();
 sg13g2_fill_1 FILLER_22_91 ();
 sg13g2_fill_2 FILLER_22_97 ();
 sg13g2_fill_1 FILLER_22_106 ();
 sg13g2_fill_2 FILLER_22_111 ();
 sg13g2_fill_1 FILLER_22_113 ();
 sg13g2_decap_4 FILLER_22_119 ();
 sg13g2_fill_2 FILLER_22_123 ();
 sg13g2_fill_1 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_fill_2 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_200 ();
 sg13g2_fill_2 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_212 ();
 sg13g2_fill_1 FILLER_22_218 ();
 sg13g2_fill_1 FILLER_22_225 ();
 sg13g2_fill_2 FILLER_22_238 ();
 sg13g2_fill_2 FILLER_22_260 ();
 sg13g2_fill_1 FILLER_22_267 ();
 sg13g2_fill_1 FILLER_22_273 ();
 sg13g2_fill_1 FILLER_22_280 ();
 sg13g2_fill_1 FILLER_22_286 ();
 sg13g2_fill_1 FILLER_22_291 ();
 sg13g2_fill_1 FILLER_22_297 ();
 sg13g2_fill_1 FILLER_22_303 ();
 sg13g2_fill_1 FILLER_22_312 ();
 sg13g2_fill_1 FILLER_22_320 ();
 sg13g2_fill_2 FILLER_22_325 ();
 sg13g2_fill_1 FILLER_22_359 ();
 sg13g2_fill_2 FILLER_22_422 ();
 sg13g2_fill_1 FILLER_22_424 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_fill_1 FILLER_23_9 ();
 sg13g2_fill_1 FILLER_23_15 ();
 sg13g2_fill_1 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_27 ();
 sg13g2_fill_1 FILLER_23_33 ();
 sg13g2_fill_2 FILLER_23_39 ();
 sg13g2_fill_1 FILLER_23_41 ();
 sg13g2_fill_1 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_55 ();
 sg13g2_fill_1 FILLER_23_61 ();
 sg13g2_decap_8 FILLER_23_67 ();
 sg13g2_fill_2 FILLER_23_74 ();
 sg13g2_fill_2 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_93 ();
 sg13g2_fill_1 FILLER_23_114 ();
 sg13g2_fill_1 FILLER_23_120 ();
 sg13g2_fill_1 FILLER_23_125 ();
 sg13g2_fill_2 FILLER_23_131 ();
 sg13g2_fill_2 FILLER_23_144 ();
 sg13g2_fill_1 FILLER_23_155 ();
 sg13g2_fill_1 FILLER_23_171 ();
 sg13g2_fill_1 FILLER_23_177 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_fill_1 FILLER_23_198 ();
 sg13g2_fill_1 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_252 ();
 sg13g2_fill_1 FILLER_23_258 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_277 ();
 sg13g2_fill_2 FILLER_23_282 ();
 sg13g2_fill_1 FILLER_23_314 ();
 sg13g2_fill_1 FILLER_23_322 ();
 sg13g2_fill_1 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_343 ();
 sg13g2_decap_4 FILLER_23_353 ();
 sg13g2_fill_2 FILLER_23_357 ();
 sg13g2_fill_1 FILLER_23_374 ();
 sg13g2_fill_2 FILLER_23_379 ();
 sg13g2_fill_1 FILLER_23_386 ();
 sg13g2_fill_2 FILLER_23_398 ();
 sg13g2_fill_2 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_418 ();
 sg13g2_decap_4 FILLER_23_425 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_fill_1 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_28 ();
 sg13g2_fill_1 FILLER_24_35 ();
 sg13g2_fill_2 FILLER_24_41 ();
 sg13g2_fill_1 FILLER_24_43 ();
 sg13g2_fill_1 FILLER_24_70 ();
 sg13g2_fill_2 FILLER_24_81 ();
 sg13g2_fill_2 FILLER_24_95 ();
 sg13g2_fill_1 FILLER_24_97 ();
 sg13g2_decap_4 FILLER_24_110 ();
 sg13g2_decap_4 FILLER_24_118 ();
 sg13g2_fill_2 FILLER_24_134 ();
 sg13g2_fill_2 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_191 ();
 sg13g2_decap_8 FILLER_24_197 ();
 sg13g2_fill_2 FILLER_24_204 ();
 sg13g2_fill_1 FILLER_24_206 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_240 ();
 sg13g2_decap_8 FILLER_24_249 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_decap_4 FILLER_24_270 ();
 sg13g2_fill_1 FILLER_24_274 ();
 sg13g2_fill_1 FILLER_24_290 ();
 sg13g2_fill_1 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_317 ();
 sg13g2_fill_1 FILLER_24_328 ();
 sg13g2_decap_8 FILLER_24_334 ();
 sg13g2_fill_2 FILLER_24_341 ();
 sg13g2_fill_1 FILLER_24_354 ();
 sg13g2_fill_2 FILLER_24_395 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_decap_4 FILLER_25_11 ();
 sg13g2_fill_2 FILLER_25_15 ();
 sg13g2_fill_1 FILLER_25_29 ();
 sg13g2_fill_1 FILLER_25_36 ();
 sg13g2_fill_1 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_58 ();
 sg13g2_fill_2 FILLER_25_68 ();
 sg13g2_fill_1 FILLER_25_79 ();
 sg13g2_fill_1 FILLER_25_85 ();
 sg13g2_fill_1 FILLER_25_90 ();
 sg13g2_fill_2 FILLER_25_95 ();
 sg13g2_fill_1 FILLER_25_102 ();
 sg13g2_fill_1 FILLER_25_121 ();
 sg13g2_fill_1 FILLER_25_142 ();
 sg13g2_fill_1 FILLER_25_148 ();
 sg13g2_fill_1 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_162 ();
 sg13g2_decap_8 FILLER_25_169 ();
 sg13g2_fill_1 FILLER_25_176 ();
 sg13g2_fill_2 FILLER_25_182 ();
 sg13g2_fill_1 FILLER_25_196 ();
 sg13g2_fill_2 FILLER_25_202 ();
 sg13g2_fill_1 FILLER_25_212 ();
 sg13g2_fill_1 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_fill_1 FILLER_25_245 ();
 sg13g2_fill_1 FILLER_25_251 ();
 sg13g2_fill_1 FILLER_25_259 ();
 sg13g2_fill_2 FILLER_25_267 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_fill_2 FILLER_25_282 ();
 sg13g2_decap_4 FILLER_25_313 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_fill_2 FILLER_25_329 ();
 sg13g2_fill_2 FILLER_25_335 ();
 sg13g2_fill_1 FILLER_25_337 ();
 sg13g2_fill_2 FILLER_25_347 ();
 sg13g2_fill_2 FILLER_25_383 ();
 sg13g2_fill_1 FILLER_25_390 ();
 sg13g2_fill_2 FILLER_25_395 ();
 sg13g2_fill_1 FILLER_25_402 ();
 sg13g2_fill_2 FILLER_25_408 ();
 sg13g2_fill_2 FILLER_25_414 ();
 sg13g2_fill_2 FILLER_25_420 ();
 sg13g2_fill_2 FILLER_25_427 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_fill_2 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_51 ();
 sg13g2_fill_1 FILLER_26_81 ();
 sg13g2_fill_1 FILLER_26_88 ();
 sg13g2_fill_1 FILLER_26_94 ();
 sg13g2_fill_2 FILLER_26_106 ();
 sg13g2_fill_1 FILLER_26_122 ();
 sg13g2_fill_1 FILLER_26_136 ();
 sg13g2_fill_1 FILLER_26_145 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_fill_2 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_199 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_fill_1 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_244 ();
 sg13g2_fill_2 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_260 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_fill_1 FILLER_26_284 ();
 sg13g2_fill_1 FILLER_26_307 ();
 sg13g2_fill_1 FILLER_26_320 ();
 sg13g2_fill_1 FILLER_26_329 ();
 sg13g2_fill_2 FILLER_26_346 ();
 sg13g2_fill_1 FILLER_26_380 ();
 sg13g2_fill_1 FILLER_26_391 ();
 sg13g2_decap_4 FILLER_26_396 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_6 ();
 sg13g2_decap_4 FILLER_27_11 ();
 sg13g2_fill_2 FILLER_27_15 ();
 sg13g2_fill_1 FILLER_27_22 ();
 sg13g2_fill_1 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_37 ();
 sg13g2_fill_1 FILLER_27_45 ();
 sg13g2_fill_2 FILLER_27_60 ();
 sg13g2_fill_2 FILLER_27_67 ();
 sg13g2_fill_1 FILLER_27_69 ();
 sg13g2_fill_1 FILLER_27_75 ();
 sg13g2_fill_2 FILLER_27_80 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_decap_4 FILLER_27_103 ();
 sg13g2_fill_2 FILLER_27_107 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_131 ();
 sg13g2_fill_1 FILLER_27_137 ();
 sg13g2_fill_1 FILLER_27_142 ();
 sg13g2_fill_1 FILLER_27_148 ();
 sg13g2_fill_2 FILLER_27_154 ();
 sg13g2_fill_2 FILLER_27_164 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_174 ();
 sg13g2_fill_1 FILLER_27_180 ();
 sg13g2_fill_2 FILLER_27_195 ();
 sg13g2_fill_1 FILLER_27_197 ();
 sg13g2_fill_2 FILLER_27_223 ();
 sg13g2_fill_2 FILLER_27_236 ();
 sg13g2_fill_2 FILLER_27_242 ();
 sg13g2_fill_1 FILLER_27_244 ();
 sg13g2_fill_1 FILLER_27_251 ();
 sg13g2_decap_4 FILLER_27_261 ();
 sg13g2_fill_1 FILLER_27_265 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_312 ();
 sg13g2_fill_2 FILLER_27_318 ();
 sg13g2_decap_8 FILLER_27_324 ();
 sg13g2_fill_1 FILLER_27_335 ();
 sg13g2_fill_2 FILLER_27_352 ();
 sg13g2_fill_1 FILLER_27_354 ();
 sg13g2_fill_1 FILLER_27_380 ();
 sg13g2_decap_4 FILLER_27_386 ();
 sg13g2_fill_2 FILLER_27_395 ();
 sg13g2_fill_2 FILLER_27_401 ();
 sg13g2_fill_2 FILLER_27_408 ();
 sg13g2_fill_1 FILLER_27_410 ();
 sg13g2_decap_4 FILLER_27_419 ();
 sg13g2_fill_2 FILLER_27_423 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_fill_2 FILLER_28_9 ();
 sg13g2_fill_1 FILLER_28_11 ();
 sg13g2_fill_2 FILLER_28_59 ();
 sg13g2_fill_1 FILLER_28_61 ();
 sg13g2_fill_2 FILLER_28_67 ();
 sg13g2_fill_1 FILLER_28_69 ();
 sg13g2_fill_1 FILLER_28_93 ();
 sg13g2_fill_1 FILLER_28_104 ();
 sg13g2_fill_1 FILLER_28_110 ();
 sg13g2_fill_2 FILLER_28_121 ();
 sg13g2_fill_2 FILLER_28_128 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_fill_1 FILLER_28_136 ();
 sg13g2_fill_2 FILLER_28_142 ();
 sg13g2_fill_1 FILLER_28_149 ();
 sg13g2_fill_2 FILLER_28_155 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_decap_8 FILLER_28_163 ();
 sg13g2_decap_4 FILLER_28_175 ();
 sg13g2_fill_1 FILLER_28_179 ();
 sg13g2_decap_4 FILLER_28_184 ();
 sg13g2_fill_2 FILLER_28_188 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_4 FILLER_28_203 ();
 sg13g2_fill_1 FILLER_28_221 ();
 sg13g2_fill_1 FILLER_28_239 ();
 sg13g2_fill_1 FILLER_28_263 ();
 sg13g2_fill_2 FILLER_28_269 ();
 sg13g2_fill_2 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_307 ();
 sg13g2_fill_2 FILLER_28_330 ();
 sg13g2_fill_1 FILLER_28_341 ();
 sg13g2_fill_1 FILLER_28_362 ();
 sg13g2_fill_2 FILLER_28_367 ();
 sg13g2_fill_1 FILLER_28_378 ();
 sg13g2_fill_1 FILLER_28_384 ();
 sg13g2_fill_1 FILLER_28_403 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_25 ();
 sg13g2_fill_1 FILLER_29_32 ();
 sg13g2_fill_2 FILLER_29_39 ();
 sg13g2_fill_1 FILLER_29_46 ();
 sg13g2_fill_2 FILLER_29_51 ();
 sg13g2_fill_1 FILLER_29_58 ();
 sg13g2_fill_1 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_69 ();
 sg13g2_decap_4 FILLER_29_75 ();
 sg13g2_decap_4 FILLER_29_86 ();
 sg13g2_fill_2 FILLER_29_95 ();
 sg13g2_fill_1 FILLER_29_97 ();
 sg13g2_fill_1 FILLER_29_102 ();
 sg13g2_fill_1 FILLER_29_111 ();
 sg13g2_fill_1 FILLER_29_120 ();
 sg13g2_fill_2 FILLER_29_126 ();
 sg13g2_fill_2 FILLER_29_134 ();
 sg13g2_fill_2 FILLER_29_141 ();
 sg13g2_fill_1 FILLER_29_143 ();
 sg13g2_fill_1 FILLER_29_173 ();
 sg13g2_fill_1 FILLER_29_188 ();
 sg13g2_fill_2 FILLER_29_193 ();
 sg13g2_fill_2 FILLER_29_235 ();
 sg13g2_fill_1 FILLER_29_237 ();
 sg13g2_fill_1 FILLER_29_264 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_fill_1 FILLER_29_282 ();
 sg13g2_fill_1 FILLER_29_287 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_309 ();
 sg13g2_fill_2 FILLER_29_318 ();
 sg13g2_fill_1 FILLER_29_320 ();
 sg13g2_fill_1 FILLER_29_353 ();
 sg13g2_fill_1 FILLER_29_359 ();
 sg13g2_fill_1 FILLER_29_365 ();
 sg13g2_fill_1 FILLER_29_371 ();
 sg13g2_fill_1 FILLER_29_420 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_fill_2 FILLER_30_13 ();
 sg13g2_fill_1 FILLER_30_20 ();
 sg13g2_fill_2 FILLER_30_26 ();
 sg13g2_fill_2 FILLER_30_39 ();
 sg13g2_fill_1 FILLER_30_41 ();
 sg13g2_decap_4 FILLER_30_47 ();
 sg13g2_fill_2 FILLER_30_51 ();
 sg13g2_fill_2 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_65 ();
 sg13g2_fill_2 FILLER_30_70 ();
 sg13g2_fill_1 FILLER_30_72 ();
 sg13g2_fill_2 FILLER_30_78 ();
 sg13g2_fill_1 FILLER_30_91 ();
 sg13g2_fill_1 FILLER_30_98 ();
 sg13g2_fill_1 FILLER_30_108 ();
 sg13g2_fill_2 FILLER_30_155 ();
 sg13g2_decap_4 FILLER_30_166 ();
 sg13g2_fill_2 FILLER_30_170 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_decap_8 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_206 ();
 sg13g2_fill_2 FILLER_30_213 ();
 sg13g2_fill_1 FILLER_30_220 ();
 sg13g2_fill_1 FILLER_30_226 ();
 sg13g2_fill_1 FILLER_30_232 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_fill_1 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_249 ();
 sg13g2_fill_2 FILLER_30_255 ();
 sg13g2_fill_2 FILLER_30_268 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_fill_1 FILLER_30_281 ();
 sg13g2_fill_1 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_323 ();
 sg13g2_fill_1 FILLER_30_325 ();
 sg13g2_fill_1 FILLER_30_331 ();
 sg13g2_decap_4 FILLER_30_337 ();
 sg13g2_fill_2 FILLER_30_375 ();
 sg13g2_fill_1 FILLER_30_381 ();
 sg13g2_fill_1 FILLER_30_386 ();
 sg13g2_fill_2 FILLER_30_390 ();
 sg13g2_fill_2 FILLER_30_398 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_16 ();
 sg13g2_fill_1 FILLER_31_22 ();
 sg13g2_fill_1 FILLER_31_28 ();
 sg13g2_fill_1 FILLER_31_34 ();
 sg13g2_fill_2 FILLER_31_39 ();
 sg13g2_fill_1 FILLER_31_57 ();
 sg13g2_decap_4 FILLER_31_67 ();
 sg13g2_fill_1 FILLER_31_71 ();
 sg13g2_fill_1 FILLER_31_78 ();
 sg13g2_fill_1 FILLER_31_83 ();
 sg13g2_fill_1 FILLER_31_101 ();
 sg13g2_fill_2 FILLER_31_108 ();
 sg13g2_fill_1 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_157 ();
 sg13g2_decap_4 FILLER_31_176 ();
 sg13g2_fill_2 FILLER_31_225 ();
 sg13g2_fill_1 FILLER_31_241 ();
 sg13g2_fill_2 FILLER_31_248 ();
 sg13g2_fill_1 FILLER_31_255 ();
 sg13g2_fill_1 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_295 ();
 sg13g2_fill_2 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_324 ();
 sg13g2_fill_1 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_356 ();
 sg13g2_fill_2 FILLER_31_372 ();
 sg13g2_fill_2 FILLER_31_400 ();
 sg13g2_fill_1 FILLER_31_407 ();
 sg13g2_fill_1 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_419 ();
 sg13g2_decap_4 FILLER_31_426 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_20 ();
 sg13g2_decap_4 FILLER_32_26 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_fill_1 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_57 ();
 sg13g2_decap_4 FILLER_32_63 ();
 sg13g2_fill_1 FILLER_32_99 ();
 sg13g2_decap_4 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_133 ();
 sg13g2_fill_2 FILLER_32_149 ();
 sg13g2_fill_1 FILLER_32_160 ();
 sg13g2_fill_1 FILLER_32_165 ();
 sg13g2_fill_1 FILLER_32_171 ();
 sg13g2_fill_1 FILLER_32_176 ();
 sg13g2_fill_1 FILLER_32_183 ();
 sg13g2_fill_2 FILLER_32_189 ();
 sg13g2_fill_2 FILLER_32_196 ();
 sg13g2_fill_2 FILLER_32_202 ();
 sg13g2_fill_1 FILLER_32_204 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_fill_1 FILLER_32_216 ();
 sg13g2_fill_1 FILLER_32_240 ();
 sg13g2_fill_2 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_252 ();
 sg13g2_fill_2 FILLER_32_259 ();
 sg13g2_fill_2 FILLER_32_311 ();
 sg13g2_fill_2 FILLER_32_329 ();
 sg13g2_fill_2 FILLER_32_336 ();
 sg13g2_fill_1 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_351 ();
 sg13g2_fill_2 FILLER_32_357 ();
 sg13g2_fill_1 FILLER_32_359 ();
 sg13g2_fill_2 FILLER_32_363 ();
 sg13g2_fill_1 FILLER_32_373 ();
 sg13g2_fill_1 FILLER_32_387 ();
 sg13g2_fill_1 FILLER_32_392 ();
 sg13g2_fill_1 FILLER_32_402 ();
 sg13g2_decap_4 FILLER_32_426 ();
 sg13g2_fill_1 FILLER_33_41 ();
 sg13g2_fill_2 FILLER_33_48 ();
 sg13g2_fill_1 FILLER_33_50 ();
 sg13g2_fill_1 FILLER_33_63 ();
 sg13g2_fill_2 FILLER_33_75 ();
 sg13g2_fill_2 FILLER_33_82 ();
 sg13g2_fill_1 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_89 ();
 sg13g2_fill_1 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_97 ();
 sg13g2_fill_1 FILLER_33_99 ();
 sg13g2_fill_2 FILLER_33_128 ();
 sg13g2_decap_4 FILLER_33_134 ();
 sg13g2_fill_1 FILLER_33_163 ();
 sg13g2_fill_2 FILLER_33_184 ();
 sg13g2_fill_1 FILLER_33_186 ();
 sg13g2_fill_2 FILLER_33_191 ();
 sg13g2_fill_2 FILLER_33_204 ();
 sg13g2_fill_1 FILLER_33_206 ();
 sg13g2_fill_2 FILLER_33_216 ();
 sg13g2_decap_4 FILLER_33_227 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_fill_2 FILLER_33_246 ();
 sg13g2_fill_2 FILLER_33_259 ();
 sg13g2_fill_2 FILLER_33_269 ();
 sg13g2_fill_2 FILLER_33_274 ();
 sg13g2_fill_1 FILLER_33_282 ();
 sg13g2_fill_2 FILLER_33_339 ();
 sg13g2_fill_2 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_fill_2 FILLER_33_376 ();
 sg13g2_fill_2 FILLER_33_387 ();
 sg13g2_fill_1 FILLER_33_398 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_2 FILLER_33_421 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_39 ();
 sg13g2_decap_4 FILLER_34_60 ();
 sg13g2_fill_1 FILLER_34_76 ();
 sg13g2_fill_2 FILLER_34_83 ();
 sg13g2_fill_1 FILLER_34_85 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_fill_2 FILLER_34_95 ();
 sg13g2_fill_1 FILLER_34_97 ();
 sg13g2_decap_4 FILLER_34_103 ();
 sg13g2_fill_1 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_fill_1 FILLER_34_142 ();
 sg13g2_fill_1 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_172 ();
 sg13g2_fill_1 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_224 ();
 sg13g2_fill_1 FILLER_34_235 ();
 sg13g2_fill_2 FILLER_34_250 ();
 sg13g2_fill_2 FILLER_34_286 ();
 sg13g2_fill_1 FILLER_34_293 ();
 sg13g2_decap_8 FILLER_34_310 ();
 sg13g2_decap_4 FILLER_34_317 ();
 sg13g2_fill_1 FILLER_34_321 ();
 sg13g2_fill_2 FILLER_34_330 ();
 sg13g2_fill_1 FILLER_34_336 ();
 sg13g2_fill_1 FILLER_34_345 ();
 sg13g2_fill_2 FILLER_34_375 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_decap_4 FILLER_34_392 ();
 sg13g2_fill_2 FILLER_34_402 ();
 sg13g2_fill_2 FILLER_35_5 ();
 sg13g2_fill_2 FILLER_35_34 ();
 sg13g2_fill_1 FILLER_35_36 ();
 sg13g2_fill_1 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_53 ();
 sg13g2_decap_4 FILLER_35_60 ();
 sg13g2_fill_1 FILLER_35_64 ();
 sg13g2_fill_2 FILLER_35_70 ();
 sg13g2_fill_1 FILLER_35_107 ();
 sg13g2_fill_1 FILLER_35_130 ();
 sg13g2_fill_1 FILLER_35_141 ();
 sg13g2_fill_1 FILLER_35_160 ();
 sg13g2_fill_1 FILLER_35_166 ();
 sg13g2_fill_2 FILLER_35_196 ();
 sg13g2_fill_1 FILLER_35_198 ();
 sg13g2_decap_4 FILLER_35_205 ();
 sg13g2_fill_2 FILLER_35_215 ();
 sg13g2_fill_1 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_234 ();
 sg13g2_fill_2 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_271 ();
 sg13g2_fill_2 FILLER_35_281 ();
 sg13g2_fill_1 FILLER_35_283 ();
 sg13g2_fill_2 FILLER_35_293 ();
 sg13g2_fill_2 FILLER_35_303 ();
 sg13g2_fill_1 FILLER_35_319 ();
 sg13g2_decap_4 FILLER_35_341 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_383 ();
 sg13g2_fill_1 FILLER_35_389 ();
 sg13g2_fill_1 FILLER_35_396 ();
 sg13g2_fill_1 FILLER_35_414 ();
 sg13g2_decap_8 FILLER_35_419 ();
 sg13g2_decap_4 FILLER_35_426 ();
 sg13g2_fill_1 FILLER_36_16 ();
 sg13g2_fill_2 FILLER_36_36 ();
 sg13g2_fill_1 FILLER_36_50 ();
 sg13g2_fill_1 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_77 ();
 sg13g2_fill_2 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_fill_2 FILLER_36_103 ();
 sg13g2_fill_2 FILLER_36_124 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_132 ();
 sg13g2_fill_1 FILLER_36_138 ();
 sg13g2_fill_1 FILLER_36_159 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_fill_2 FILLER_36_192 ();
 sg13g2_fill_2 FILLER_36_198 ();
 sg13g2_fill_2 FILLER_36_204 ();
 sg13g2_fill_1 FILLER_36_206 ();
 sg13g2_decap_4 FILLER_36_220 ();
 sg13g2_fill_1 FILLER_36_224 ();
 sg13g2_fill_2 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_286 ();
 sg13g2_fill_1 FILLER_36_288 ();
 sg13g2_fill_2 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_295 ();
 sg13g2_fill_2 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_315 ();
 sg13g2_fill_1 FILLER_36_320 ();
 sg13g2_fill_1 FILLER_36_325 ();
 sg13g2_fill_1 FILLER_36_332 ();
 sg13g2_fill_2 FILLER_36_338 ();
 sg13g2_fill_1 FILLER_36_345 ();
 sg13g2_fill_1 FILLER_36_395 ();
 sg13g2_fill_2 FILLER_36_411 ();
 sg13g2_fill_1 FILLER_36_418 ();
 sg13g2_decap_8 FILLER_36_423 ();
 sg13g2_fill_1 FILLER_37_45 ();
 sg13g2_fill_2 FILLER_37_59 ();
 sg13g2_fill_1 FILLER_37_66 ();
 sg13g2_fill_1 FILLER_37_72 ();
 sg13g2_fill_1 FILLER_37_77 ();
 sg13g2_fill_1 FILLER_37_98 ();
 sg13g2_fill_1 FILLER_37_104 ();
 sg13g2_fill_2 FILLER_37_112 ();
 sg13g2_decap_4 FILLER_37_124 ();
 sg13g2_fill_1 FILLER_37_128 ();
 sg13g2_fill_1 FILLER_37_134 ();
 sg13g2_fill_2 FILLER_37_140 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_fill_2 FILLER_37_155 ();
 sg13g2_fill_2 FILLER_37_183 ();
 sg13g2_fill_2 FILLER_37_224 ();
 sg13g2_fill_1 FILLER_37_226 ();
 sg13g2_fill_2 FILLER_37_260 ();
 sg13g2_fill_2 FILLER_37_270 ();
 sg13g2_fill_2 FILLER_37_315 ();
 sg13g2_fill_2 FILLER_37_346 ();
 sg13g2_fill_1 FILLER_37_383 ();
 sg13g2_fill_1 FILLER_37_387 ();
 sg13g2_fill_1 FILLER_37_393 ();
 sg13g2_fill_1 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_12 ();
 sg13g2_fill_1 FILLER_38_32 ();
 sg13g2_fill_2 FILLER_38_37 ();
 sg13g2_decap_4 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_53 ();
 sg13g2_fill_2 FILLER_38_58 ();
 sg13g2_fill_1 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_81 ();
 sg13g2_fill_2 FILLER_38_85 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_fill_2 FILLER_38_104 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_fill_1 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_153 ();
 sg13g2_fill_1 FILLER_38_232 ();
 sg13g2_fill_2 FILLER_38_288 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_309 ();
 sg13g2_decap_4 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_fill_2 FILLER_38_380 ();
 sg13g2_fill_1 FILLER_38_387 ();
 sg13g2_fill_2 FILLER_38_401 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_2 FILLER_38_412 ();
 sg13g2_fill_2 FILLER_38_418 ();
 sg13g2_fill_1 FILLER_38_420 ();
 sg13g2_decap_4 FILLER_38_426 ();
 sg13g2_fill_1 FILLER_39_16 ();
 sg13g2_fill_1 FILLER_39_22 ();
 sg13g2_fill_2 FILLER_39_40 ();
 sg13g2_fill_1 FILLER_39_42 ();
 sg13g2_fill_1 FILLER_39_48 ();
 sg13g2_decap_4 FILLER_39_59 ();
 sg13g2_fill_2 FILLER_39_71 ();
 sg13g2_fill_1 FILLER_39_73 ();
 sg13g2_fill_1 FILLER_39_87 ();
 sg13g2_fill_1 FILLER_39_96 ();
 sg13g2_fill_2 FILLER_39_102 ();
 sg13g2_fill_1 FILLER_39_112 ();
 sg13g2_fill_1 FILLER_39_127 ();
 sg13g2_fill_2 FILLER_39_132 ();
 sg13g2_fill_2 FILLER_39_148 ();
 sg13g2_fill_1 FILLER_39_154 ();
 sg13g2_fill_2 FILLER_39_164 ();
 sg13g2_fill_2 FILLER_39_170 ();
 sg13g2_fill_1 FILLER_39_176 ();
 sg13g2_fill_1 FILLER_39_201 ();
 sg13g2_fill_1 FILLER_39_235 ();
 sg13g2_fill_1 FILLER_39_241 ();
 sg13g2_fill_1 FILLER_39_246 ();
 sg13g2_fill_1 FILLER_39_251 ();
 sg13g2_fill_2 FILLER_39_261 ();
 sg13g2_fill_1 FILLER_39_284 ();
 sg13g2_decap_4 FILLER_39_315 ();
 sg13g2_fill_2 FILLER_39_332 ();
 sg13g2_fill_1 FILLER_39_334 ();
 sg13g2_fill_1 FILLER_39_368 ();
 sg13g2_fill_2 FILLER_39_394 ();
 sg13g2_fill_1 FILLER_39_396 ();
 sg13g2_fill_2 FILLER_39_402 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_7 ();
 sg13g2_fill_2 FILLER_40_13 ();
 sg13g2_fill_1 FILLER_40_20 ();
 sg13g2_fill_2 FILLER_40_26 ();
 sg13g2_fill_1 FILLER_40_32 ();
 sg13g2_fill_2 FILLER_40_66 ();
 sg13g2_fill_2 FILLER_40_93 ();
 sg13g2_fill_1 FILLER_40_95 ();
 sg13g2_fill_2 FILLER_40_101 ();
 sg13g2_fill_1 FILLER_40_103 ();
 sg13g2_fill_1 FILLER_40_110 ();
 sg13g2_fill_2 FILLER_40_117 ();
 sg13g2_fill_1 FILLER_40_127 ();
 sg13g2_fill_1 FILLER_40_132 ();
 sg13g2_fill_2 FILLER_40_137 ();
 sg13g2_fill_1 FILLER_40_139 ();
 sg13g2_fill_2 FILLER_40_152 ();
 sg13g2_fill_2 FILLER_40_162 ();
 sg13g2_fill_1 FILLER_40_173 ();
 sg13g2_fill_2 FILLER_40_179 ();
 sg13g2_fill_2 FILLER_40_214 ();
 sg13g2_fill_2 FILLER_40_220 ();
 sg13g2_fill_1 FILLER_40_242 ();
 sg13g2_fill_1 FILLER_40_266 ();
 sg13g2_fill_1 FILLER_40_272 ();
 sg13g2_fill_1 FILLER_40_281 ();
 sg13g2_fill_1 FILLER_40_290 ();
 sg13g2_fill_1 FILLER_40_295 ();
 sg13g2_fill_2 FILLER_40_300 ();
 sg13g2_fill_2 FILLER_40_311 ();
 sg13g2_fill_2 FILLER_40_324 ();
 sg13g2_fill_1 FILLER_40_326 ();
 sg13g2_fill_1 FILLER_40_366 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_fill_2 FILLER_40_377 ();
 sg13g2_fill_1 FILLER_40_390 ();
 sg13g2_fill_2 FILLER_40_398 ();
 sg13g2_decap_8 FILLER_40_405 ();
 sg13g2_decap_4 FILLER_40_412 ();
 sg13g2_fill_1 FILLER_40_416 ();
 sg13g2_decap_4 FILLER_41_8 ();
 sg13g2_fill_2 FILLER_41_12 ();
 sg13g2_fill_1 FILLER_41_40 ();
 sg13g2_fill_1 FILLER_41_46 ();
 sg13g2_fill_1 FILLER_41_55 ();
 sg13g2_fill_1 FILLER_41_61 ();
 sg13g2_fill_1 FILLER_41_72 ();
 sg13g2_fill_1 FILLER_41_81 ();
 sg13g2_fill_1 FILLER_41_86 ();
 sg13g2_fill_2 FILLER_41_92 ();
 sg13g2_fill_2 FILLER_41_103 ();
 sg13g2_decap_8 FILLER_41_110 ();
 sg13g2_fill_2 FILLER_41_125 ();
 sg13g2_fill_1 FILLER_41_127 ();
 sg13g2_fill_1 FILLER_41_133 ();
 sg13g2_fill_2 FILLER_41_160 ();
 sg13g2_fill_2 FILLER_41_189 ();
 sg13g2_fill_1 FILLER_41_200 ();
 sg13g2_fill_2 FILLER_41_216 ();
 sg13g2_decap_8 FILLER_41_223 ();
 sg13g2_fill_1 FILLER_41_290 ();
 sg13g2_fill_1 FILLER_41_295 ();
 sg13g2_decap_4 FILLER_41_335 ();
 sg13g2_fill_1 FILLER_41_339 ();
 sg13g2_fill_2 FILLER_41_350 ();
 sg13g2_fill_2 FILLER_41_356 ();
 sg13g2_fill_2 FILLER_41_366 ();
 sg13g2_fill_1 FILLER_41_368 ();
 sg13g2_fill_2 FILLER_41_381 ();
 sg13g2_fill_1 FILLER_41_396 ();
 sg13g2_fill_1 FILLER_41_423 ();
 sg13g2_fill_2 FILLER_41_428 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_13 ();
 sg13g2_fill_1 FILLER_42_19 ();
 sg13g2_decap_8 FILLER_42_31 ();
 sg13g2_decap_8 FILLER_42_38 ();
 sg13g2_fill_1 FILLER_42_45 ();
 sg13g2_fill_2 FILLER_42_55 ();
 sg13g2_fill_1 FILLER_42_57 ();
 sg13g2_decap_4 FILLER_42_67 ();
 sg13g2_fill_1 FILLER_42_83 ();
 sg13g2_fill_1 FILLER_42_113 ();
 sg13g2_fill_2 FILLER_42_130 ();
 sg13g2_fill_1 FILLER_42_160 ();
 sg13g2_fill_1 FILLER_42_165 ();
 sg13g2_fill_1 FILLER_42_176 ();
 sg13g2_fill_1 FILLER_42_182 ();
 sg13g2_fill_1 FILLER_42_232 ();
 sg13g2_fill_1 FILLER_42_259 ();
 sg13g2_fill_1 FILLER_42_273 ();
 sg13g2_fill_1 FILLER_42_278 ();
 sg13g2_fill_1 FILLER_42_283 ();
 sg13g2_fill_1 FILLER_42_304 ();
 sg13g2_fill_2 FILLER_42_309 ();
 sg13g2_decap_4 FILLER_42_317 ();
 sg13g2_fill_2 FILLER_42_321 ();
 sg13g2_fill_2 FILLER_42_335 ();
 sg13g2_fill_1 FILLER_42_337 ();
 sg13g2_fill_2 FILLER_42_348 ();
 sg13g2_fill_2 FILLER_42_359 ();
 sg13g2_decap_4 FILLER_42_366 ();
 sg13g2_fill_1 FILLER_42_370 ();
 sg13g2_fill_1 FILLER_42_410 ();
 sg13g2_decap_4 FILLER_42_424 ();
 sg13g2_fill_2 FILLER_42_428 ();
 sg13g2_fill_1 FILLER_43_44 ();
 sg13g2_fill_1 FILLER_43_58 ();
 sg13g2_fill_1 FILLER_43_63 ();
 sg13g2_fill_1 FILLER_43_76 ();
 sg13g2_fill_1 FILLER_43_82 ();
 sg13g2_fill_2 FILLER_43_92 ();
 sg13g2_fill_1 FILLER_43_99 ();
 sg13g2_fill_2 FILLER_43_105 ();
 sg13g2_fill_1 FILLER_43_107 ();
 sg13g2_fill_2 FILLER_43_113 ();
 sg13g2_fill_1 FILLER_43_115 ();
 sg13g2_fill_1 FILLER_43_167 ();
 sg13g2_fill_1 FILLER_43_189 ();
 sg13g2_fill_1 FILLER_43_228 ();
 sg13g2_fill_1 FILLER_43_242 ();
 sg13g2_fill_1 FILLER_43_267 ();
 sg13g2_decap_4 FILLER_43_304 ();
 sg13g2_fill_1 FILLER_43_308 ();
 sg13g2_fill_2 FILLER_43_313 ();
 sg13g2_fill_1 FILLER_43_320 ();
 sg13g2_fill_1 FILLER_43_335 ();
 sg13g2_fill_2 FILLER_43_345 ();
 sg13g2_fill_1 FILLER_43_347 ();
 sg13g2_decap_4 FILLER_43_373 ();
 sg13g2_fill_2 FILLER_43_377 ();
 sg13g2_fill_1 FILLER_43_395 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_4 FILLER_43_414 ();
 sg13g2_fill_1 FILLER_43_418 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_11 ();
 sg13g2_fill_1 FILLER_44_16 ();
 sg13g2_fill_1 FILLER_44_27 ();
 sg13g2_fill_2 FILLER_44_31 ();
 sg13g2_fill_2 FILLER_44_37 ();
 sg13g2_fill_1 FILLER_44_39 ();
 sg13g2_fill_1 FILLER_44_47 ();
 sg13g2_fill_2 FILLER_44_55 ();
 sg13g2_fill_1 FILLER_44_57 ();
 sg13g2_fill_2 FILLER_44_71 ();
 sg13g2_fill_2 FILLER_44_83 ();
 sg13g2_fill_1 FILLER_44_85 ();
 sg13g2_fill_1 FILLER_44_90 ();
 sg13g2_fill_1 FILLER_44_95 ();
 sg13g2_fill_1 FILLER_44_100 ();
 sg13g2_fill_1 FILLER_44_117 ();
 sg13g2_fill_1 FILLER_44_125 ();
 sg13g2_fill_1 FILLER_44_131 ();
 sg13g2_fill_1 FILLER_44_136 ();
 sg13g2_fill_2 FILLER_44_142 ();
 sg13g2_fill_2 FILLER_44_148 ();
 sg13g2_fill_1 FILLER_44_171 ();
 sg13g2_fill_2 FILLER_44_184 ();
 sg13g2_fill_2 FILLER_44_190 ();
 sg13g2_fill_2 FILLER_44_200 ();
 sg13g2_fill_2 FILLER_44_207 ();
 sg13g2_fill_1 FILLER_44_209 ();
 sg13g2_fill_1 FILLER_44_215 ();
 sg13g2_fill_2 FILLER_44_222 ();
 sg13g2_fill_1 FILLER_44_224 ();
 sg13g2_fill_2 FILLER_44_281 ();
 sg13g2_fill_1 FILLER_44_288 ();
 sg13g2_decap_4 FILLER_44_315 ();
 sg13g2_fill_2 FILLER_44_319 ();
 sg13g2_fill_1 FILLER_44_340 ();
 sg13g2_fill_1 FILLER_44_346 ();
 sg13g2_fill_1 FILLER_44_352 ();
 sg13g2_decap_4 FILLER_44_367 ();
 sg13g2_fill_1 FILLER_44_378 ();
 sg13g2_fill_1 FILLER_44_384 ();
 sg13g2_fill_1 FILLER_44_391 ();
 sg13g2_fill_1 FILLER_44_397 ();
 sg13g2_fill_1 FILLER_44_403 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_10 ();
 sg13g2_fill_1 FILLER_45_23 ();
 sg13g2_fill_1 FILLER_45_34 ();
 sg13g2_fill_2 FILLER_45_47 ();
 sg13g2_fill_1 FILLER_45_49 ();
 sg13g2_fill_1 FILLER_45_54 ();
 sg13g2_fill_2 FILLER_45_63 ();
 sg13g2_fill_1 FILLER_45_84 ();
 sg13g2_fill_2 FILLER_45_103 ();
 sg13g2_fill_1 FILLER_45_105 ();
 sg13g2_fill_1 FILLER_45_111 ();
 sg13g2_fill_1 FILLER_45_126 ();
 sg13g2_fill_1 FILLER_45_132 ();
 sg13g2_fill_2 FILLER_45_141 ();
 sg13g2_fill_1 FILLER_45_143 ();
 sg13g2_fill_1 FILLER_45_153 ();
 sg13g2_fill_1 FILLER_45_164 ();
 sg13g2_fill_1 FILLER_45_177 ();
 sg13g2_fill_1 FILLER_45_204 ();
 sg13g2_fill_2 FILLER_45_218 ();
 sg13g2_fill_2 FILLER_45_225 ();
 sg13g2_fill_1 FILLER_45_227 ();
 sg13g2_fill_2 FILLER_45_251 ();
 sg13g2_fill_2 FILLER_45_263 ();
 sg13g2_fill_1 FILLER_45_270 ();
 sg13g2_fill_2 FILLER_45_275 ();
 sg13g2_fill_1 FILLER_45_277 ();
 sg13g2_fill_1 FILLER_45_283 ();
 sg13g2_fill_1 FILLER_45_297 ();
 sg13g2_fill_1 FILLER_45_303 ();
 sg13g2_decap_8 FILLER_45_309 ();
 sg13g2_decap_4 FILLER_45_338 ();
 sg13g2_fill_1 FILLER_45_342 ();
 sg13g2_fill_2 FILLER_45_363 ();
 sg13g2_fill_2 FILLER_45_377 ();
 sg13g2_fill_1 FILLER_45_391 ();
 sg13g2_fill_1 FILLER_45_399 ();
 sg13g2_fill_1 FILLER_45_413 ();
 sg13g2_fill_1 FILLER_45_418 ();
 sg13g2_fill_1 FILLER_45_424 ();
 sg13g2_fill_1 FILLER_45_429 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_17 ();
 sg13g2_fill_2 FILLER_46_40 ();
 sg13g2_fill_2 FILLER_46_61 ();
 sg13g2_fill_1 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_71 ();
 sg13g2_decap_4 FILLER_46_87 ();
 sg13g2_fill_1 FILLER_46_106 ();
 sg13g2_fill_1 FILLER_46_111 ();
 sg13g2_fill_1 FILLER_46_116 ();
 sg13g2_fill_1 FILLER_46_122 ();
 sg13g2_fill_1 FILLER_46_127 ();
 sg13g2_fill_2 FILLER_46_131 ();
 sg13g2_fill_2 FILLER_46_138 ();
 sg13g2_fill_1 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_149 ();
 sg13g2_fill_2 FILLER_46_156 ();
 sg13g2_fill_2 FILLER_46_174 ();
 sg13g2_fill_2 FILLER_46_181 ();
 sg13g2_fill_1 FILLER_46_187 ();
 sg13g2_fill_1 FILLER_46_197 ();
 sg13g2_decap_4 FILLER_46_203 ();
 sg13g2_decap_4 FILLER_46_268 ();
 sg13g2_fill_2 FILLER_46_282 ();
 sg13g2_fill_1 FILLER_46_310 ();
 sg13g2_fill_1 FILLER_46_315 ();
 sg13g2_fill_1 FILLER_46_320 ();
 sg13g2_fill_1 FILLER_46_326 ();
 sg13g2_fill_1 FILLER_46_332 ();
 sg13g2_fill_1 FILLER_46_340 ();
 sg13g2_fill_1 FILLER_46_371 ();
 sg13g2_fill_2 FILLER_46_382 ();
 sg13g2_fill_1 FILLER_46_384 ();
 sg13g2_fill_2 FILLER_46_401 ();
 sg13g2_fill_1 FILLER_46_429 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_2 ();
 sg13g2_fill_2 FILLER_47_8 ();
 sg13g2_fill_2 FILLER_47_34 ();
 sg13g2_fill_2 FILLER_47_55 ();
 sg13g2_fill_1 FILLER_47_57 ();
 sg13g2_fill_2 FILLER_47_67 ();
 sg13g2_fill_1 FILLER_47_74 ();
 sg13g2_fill_2 FILLER_47_127 ();
 sg13g2_fill_2 FILLER_47_144 ();
 sg13g2_decap_8 FILLER_47_149 ();
 sg13g2_decap_4 FILLER_47_156 ();
 sg13g2_fill_2 FILLER_47_160 ();
 sg13g2_fill_1 FILLER_47_172 ();
 sg13g2_fill_2 FILLER_47_182 ();
 sg13g2_fill_1 FILLER_47_184 ();
 sg13g2_decap_4 FILLER_47_189 ();
 sg13g2_fill_2 FILLER_47_209 ();
 sg13g2_fill_1 FILLER_47_211 ();
 sg13g2_fill_1 FILLER_47_217 ();
 sg13g2_fill_1 FILLER_47_227 ();
 sg13g2_fill_1 FILLER_47_236 ();
 sg13g2_fill_1 FILLER_47_282 ();
 sg13g2_fill_2 FILLER_47_287 ();
 sg13g2_fill_2 FILLER_47_302 ();
 sg13g2_fill_2 FILLER_47_308 ();
 sg13g2_fill_1 FILLER_47_315 ();
 sg13g2_fill_1 FILLER_47_320 ();
 sg13g2_fill_1 FILLER_47_329 ();
 sg13g2_fill_1 FILLER_47_335 ();
 sg13g2_fill_1 FILLER_47_340 ();
 sg13g2_fill_1 FILLER_47_345 ();
 sg13g2_fill_2 FILLER_47_350 ();
 sg13g2_fill_1 FILLER_47_352 ();
 sg13g2_fill_1 FILLER_47_370 ();
 sg13g2_decap_4 FILLER_47_377 ();
 sg13g2_fill_2 FILLER_47_381 ();
 sg13g2_decap_4 FILLER_47_391 ();
 sg13g2_fill_1 FILLER_47_395 ();
 sg13g2_fill_2 FILLER_47_415 ();
 sg13g2_fill_2 FILLER_48_13 ();
 sg13g2_fill_1 FILLER_48_37 ();
 sg13g2_fill_2 FILLER_48_43 ();
 sg13g2_fill_1 FILLER_48_45 ();
 sg13g2_decap_4 FILLER_48_51 ();
 sg13g2_fill_2 FILLER_48_55 ();
 sg13g2_fill_2 FILLER_48_78 ();
 sg13g2_fill_1 FILLER_48_84 ();
 sg13g2_fill_1 FILLER_48_95 ();
 sg13g2_fill_1 FILLER_48_112 ();
 sg13g2_fill_1 FILLER_48_127 ();
 sg13g2_fill_1 FILLER_48_134 ();
 sg13g2_fill_2 FILLER_48_147 ();
 sg13g2_fill_2 FILLER_48_158 ();
 sg13g2_fill_1 FILLER_48_160 ();
 sg13g2_fill_1 FILLER_48_176 ();
 sg13g2_fill_2 FILLER_48_194 ();
 sg13g2_decap_4 FILLER_48_208 ();
 sg13g2_fill_1 FILLER_48_212 ();
 sg13g2_fill_2 FILLER_48_218 ();
 sg13g2_fill_1 FILLER_48_251 ();
 sg13g2_fill_2 FILLER_48_260 ();
 sg13g2_fill_1 FILLER_48_266 ();
 sg13g2_fill_1 FILLER_48_272 ();
 sg13g2_fill_1 FILLER_48_282 ();
 sg13g2_fill_1 FILLER_48_288 ();
 sg13g2_fill_1 FILLER_48_315 ();
 sg13g2_fill_1 FILLER_48_320 ();
 sg13g2_fill_1 FILLER_48_329 ();
 sg13g2_fill_1 FILLER_48_348 ();
 sg13g2_fill_2 FILLER_48_366 ();
 sg13g2_fill_1 FILLER_48_368 ();
 sg13g2_fill_1 FILLER_48_374 ();
 sg13g2_fill_2 FILLER_48_382 ();
 sg13g2_fill_1 FILLER_48_389 ();
 sg13g2_fill_1 FILLER_48_394 ();
 sg13g2_fill_2 FILLER_48_400 ();
 sg13g2_fill_2 FILLER_48_428 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_6 ();
 sg13g2_fill_1 FILLER_49_13 ();
 sg13g2_fill_1 FILLER_49_25 ();
 sg13g2_fill_1 FILLER_49_53 ();
 sg13g2_fill_2 FILLER_49_75 ();
 sg13g2_fill_2 FILLER_49_82 ();
 sg13g2_fill_2 FILLER_49_100 ();
 sg13g2_fill_1 FILLER_49_110 ();
 sg13g2_fill_2 FILLER_49_115 ();
 sg13g2_fill_1 FILLER_49_117 ();
 sg13g2_fill_1 FILLER_49_128 ();
 sg13g2_fill_2 FILLER_49_133 ();
 sg13g2_fill_1 FILLER_49_144 ();
 sg13g2_fill_1 FILLER_49_170 ();
 sg13g2_fill_1 FILLER_49_176 ();
 sg13g2_fill_1 FILLER_49_185 ();
 sg13g2_fill_2 FILLER_49_212 ();
 sg13g2_fill_2 FILLER_49_223 ();
 sg13g2_fill_1 FILLER_49_225 ();
 sg13g2_fill_1 FILLER_49_247 ();
 sg13g2_fill_1 FILLER_49_257 ();
 sg13g2_fill_1 FILLER_49_295 ();
 sg13g2_fill_2 FILLER_49_312 ();
 sg13g2_fill_1 FILLER_49_314 ();
 sg13g2_fill_2 FILLER_49_340 ();
 sg13g2_fill_2 FILLER_49_354 ();
 sg13g2_fill_2 FILLER_49_361 ();
 sg13g2_fill_2 FILLER_49_368 ();
 sg13g2_fill_1 FILLER_49_412 ();
 sg13g2_decap_4 FILLER_49_417 ();
 sg13g2_decap_4 FILLER_49_426 ();
 sg13g2_fill_1 FILLER_50_30 ();
 sg13g2_decap_8 FILLER_50_45 ();
 sg13g2_fill_1 FILLER_50_52 ();
 sg13g2_fill_2 FILLER_50_57 ();
 sg13g2_decap_4 FILLER_50_64 ();
 sg13g2_fill_1 FILLER_50_68 ();
 sg13g2_fill_2 FILLER_50_79 ();
 sg13g2_fill_1 FILLER_50_86 ();
 sg13g2_fill_2 FILLER_50_91 ();
 sg13g2_fill_2 FILLER_50_99 ();
 sg13g2_fill_1 FILLER_50_105 ();
 sg13g2_fill_1 FILLER_50_116 ();
 sg13g2_fill_2 FILLER_50_124 ();
 sg13g2_decap_4 FILLER_50_131 ();
 sg13g2_fill_2 FILLER_50_158 ();
 sg13g2_fill_1 FILLER_50_202 ();
 sg13g2_fill_1 FILLER_50_211 ();
 sg13g2_fill_2 FILLER_50_229 ();
 sg13g2_fill_1 FILLER_50_239 ();
 sg13g2_fill_2 FILLER_50_253 ();
 sg13g2_fill_1 FILLER_50_298 ();
 sg13g2_fill_2 FILLER_50_303 ();
 sg13g2_fill_1 FILLER_50_310 ();
 sg13g2_fill_2 FILLER_50_315 ();
 sg13g2_fill_1 FILLER_50_317 ();
 sg13g2_fill_2 FILLER_50_345 ();
 sg13g2_fill_2 FILLER_50_353 ();
 sg13g2_fill_1 FILLER_50_355 ();
 sg13g2_fill_1 FILLER_50_371 ();
 sg13g2_fill_1 FILLER_50_396 ();
 sg13g2_fill_2 FILLER_50_402 ();
 sg13g2_fill_2 FILLER_51_26 ();
 sg13g2_decap_4 FILLER_51_43 ();
 sg13g2_fill_1 FILLER_51_47 ();
 sg13g2_fill_1 FILLER_51_59 ();
 sg13g2_decap_4 FILLER_51_66 ();
 sg13g2_fill_1 FILLER_51_74 ();
 sg13g2_fill_2 FILLER_51_84 ();
 sg13g2_fill_2 FILLER_51_107 ();
 sg13g2_fill_1 FILLER_51_124 ();
 sg13g2_fill_1 FILLER_51_151 ();
 sg13g2_fill_2 FILLER_51_163 ();
 sg13g2_fill_1 FILLER_51_169 ();
 sg13g2_fill_1 FILLER_51_175 ();
 sg13g2_fill_1 FILLER_51_186 ();
 sg13g2_fill_1 FILLER_51_195 ();
 sg13g2_fill_1 FILLER_51_201 ();
 sg13g2_fill_1 FILLER_51_206 ();
 sg13g2_fill_2 FILLER_51_266 ();
 sg13g2_fill_1 FILLER_51_298 ();
 sg13g2_fill_1 FILLER_51_303 ();
 sg13g2_fill_1 FILLER_51_309 ();
 sg13g2_fill_1 FILLER_51_320 ();
 sg13g2_fill_1 FILLER_51_331 ();
 sg13g2_fill_1 FILLER_51_364 ();
 sg13g2_fill_1 FILLER_51_392 ();
 sg13g2_fill_1 FILLER_51_412 ();
 sg13g2_decap_8 FILLER_51_421 ();
 sg13g2_fill_2 FILLER_51_428 ();
 sg13g2_fill_1 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_9 ();
 sg13g2_fill_1 FILLER_52_14 ();
 sg13g2_fill_2 FILLER_52_25 ();
 sg13g2_fill_1 FILLER_52_27 ();
 sg13g2_fill_2 FILLER_52_48 ();
 sg13g2_fill_2 FILLER_52_55 ();
 sg13g2_fill_1 FILLER_52_62 ();
 sg13g2_fill_1 FILLER_52_89 ();
 sg13g2_fill_1 FILLER_52_96 ();
 sg13g2_fill_1 FILLER_52_113 ();
 sg13g2_decap_4 FILLER_52_119 ();
 sg13g2_fill_2 FILLER_52_163 ();
 sg13g2_fill_1 FILLER_52_165 ();
 sg13g2_fill_1 FILLER_52_186 ();
 sg13g2_fill_1 FILLER_52_192 ();
 sg13g2_fill_2 FILLER_52_198 ();
 sg13g2_fill_1 FILLER_52_212 ();
 sg13g2_fill_2 FILLER_52_226 ();
 sg13g2_fill_1 FILLER_52_238 ();
 sg13g2_fill_1 FILLER_52_243 ();
 sg13g2_fill_2 FILLER_52_254 ();
 sg13g2_fill_1 FILLER_52_279 ();
 sg13g2_fill_2 FILLER_52_298 ();
 sg13g2_fill_1 FILLER_52_305 ();
 sg13g2_fill_2 FILLER_52_311 ();
 sg13g2_fill_1 FILLER_52_330 ();
 sg13g2_fill_2 FILLER_52_371 ();
 sg13g2_fill_1 FILLER_52_373 ();
 sg13g2_fill_1 FILLER_52_392 ();
 sg13g2_fill_2 FILLER_52_398 ();
 sg13g2_decap_4 FILLER_53_0 ();
 sg13g2_decap_4 FILLER_53_12 ();
 sg13g2_fill_1 FILLER_53_16 ();
 sg13g2_fill_1 FILLER_53_22 ();
 sg13g2_fill_1 FILLER_53_28 ();
 sg13g2_fill_1 FILLER_53_34 ();
 sg13g2_fill_1 FILLER_53_46 ();
 sg13g2_fill_2 FILLER_53_52 ();
 sg13g2_fill_1 FILLER_53_54 ();
 sg13g2_fill_2 FILLER_53_60 ();
 sg13g2_fill_2 FILLER_53_67 ();
 sg13g2_fill_1 FILLER_53_69 ();
 sg13g2_fill_1 FILLER_53_75 ();
 sg13g2_fill_2 FILLER_53_84 ();
 sg13g2_fill_1 FILLER_53_86 ();
 sg13g2_decap_4 FILLER_53_100 ();
 sg13g2_fill_1 FILLER_53_132 ();
 sg13g2_fill_1 FILLER_53_161 ();
 sg13g2_fill_2 FILLER_53_174 ();
 sg13g2_fill_1 FILLER_53_176 ();
 sg13g2_fill_2 FILLER_53_199 ();
 sg13g2_decap_8 FILLER_53_206 ();
 sg13g2_fill_1 FILLER_53_246 ();
 sg13g2_decap_4 FILLER_53_273 ();
 sg13g2_fill_1 FILLER_53_277 ();
 sg13g2_fill_1 FILLER_53_320 ();
 sg13g2_fill_1 FILLER_53_330 ();
 sg13g2_fill_1 FILLER_53_339 ();
 sg13g2_fill_1 FILLER_53_348 ();
 sg13g2_fill_1 FILLER_53_354 ();
 sg13g2_fill_1 FILLER_53_370 ();
 sg13g2_fill_2 FILLER_53_376 ();
 sg13g2_fill_2 FILLER_53_383 ();
 sg13g2_decap_4 FILLER_53_392 ();
 sg13g2_fill_2 FILLER_53_401 ();
 sg13g2_fill_1 FILLER_53_403 ();
 sg13g2_fill_1 FILLER_54_32 ();
 sg13g2_fill_2 FILLER_54_59 ();
 sg13g2_fill_1 FILLER_54_71 ();
 sg13g2_fill_2 FILLER_54_77 ();
 sg13g2_fill_1 FILLER_54_79 ();
 sg13g2_fill_2 FILLER_54_106 ();
 sg13g2_fill_1 FILLER_54_108 ();
 sg13g2_fill_2 FILLER_54_125 ();
 sg13g2_fill_1 FILLER_54_127 ();
 sg13g2_fill_1 FILLER_54_136 ();
 sg13g2_fill_1 FILLER_54_147 ();
 sg13g2_fill_1 FILLER_54_193 ();
 sg13g2_decap_4 FILLER_54_215 ();
 sg13g2_fill_2 FILLER_54_219 ();
 sg13g2_fill_2 FILLER_54_225 ();
 sg13g2_fill_1 FILLER_54_227 ();
 sg13g2_fill_1 FILLER_54_231 ();
 sg13g2_fill_1 FILLER_54_236 ();
 sg13g2_fill_1 FILLER_54_242 ();
 sg13g2_fill_2 FILLER_54_257 ();
 sg13g2_decap_8 FILLER_54_274 ();
 sg13g2_fill_2 FILLER_54_359 ();
 sg13g2_fill_2 FILLER_54_393 ();
 sg13g2_decap_4 FILLER_54_403 ();
 sg13g2_fill_2 FILLER_54_412 ();
 sg13g2_fill_1 FILLER_54_414 ();
 sg13g2_decap_8 FILLER_54_419 ();
 sg13g2_decap_4 FILLER_54_426 ();
 sg13g2_fill_1 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_6 ();
 sg13g2_fill_1 FILLER_55_12 ();
 sg13g2_fill_2 FILLER_55_18 ();
 sg13g2_fill_1 FILLER_55_37 ();
 sg13g2_fill_1 FILLER_55_43 ();
 sg13g2_fill_1 FILLER_55_48 ();
 sg13g2_fill_1 FILLER_55_59 ();
 sg13g2_fill_1 FILLER_55_64 ();
 sg13g2_fill_2 FILLER_55_71 ();
 sg13g2_fill_1 FILLER_55_78 ();
 sg13g2_fill_1 FILLER_55_85 ();
 sg13g2_fill_1 FILLER_55_90 ();
 sg13g2_decap_4 FILLER_55_95 ();
 sg13g2_fill_1 FILLER_55_99 ();
 sg13g2_fill_2 FILLER_55_104 ();
 sg13g2_fill_1 FILLER_55_111 ();
 sg13g2_fill_1 FILLER_55_117 ();
 sg13g2_fill_1 FILLER_55_123 ();
 sg13g2_fill_2 FILLER_55_129 ();
 sg13g2_decap_8 FILLER_55_135 ();
 sg13g2_fill_2 FILLER_55_149 ();
 sg13g2_fill_2 FILLER_55_158 ();
 sg13g2_fill_2 FILLER_55_202 ();
 sg13g2_fill_1 FILLER_55_230 ();
 sg13g2_decap_4 FILLER_55_236 ();
 sg13g2_fill_1 FILLER_55_245 ();
 sg13g2_fill_2 FILLER_55_259 ();
 sg13g2_fill_2 FILLER_55_267 ();
 sg13g2_fill_1 FILLER_55_269 ();
 sg13g2_fill_1 FILLER_55_294 ();
 sg13g2_fill_2 FILLER_55_308 ();
 sg13g2_fill_1 FILLER_55_328 ();
 sg13g2_fill_1 FILLER_55_344 ();
 sg13g2_fill_2 FILLER_55_366 ();
 sg13g2_fill_2 FILLER_55_372 ();
 sg13g2_fill_1 FILLER_55_379 ();
 sg13g2_fill_1 FILLER_55_385 ();
 sg13g2_fill_1 FILLER_55_395 ();
 sg13g2_fill_1 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_5 ();
 sg13g2_fill_2 FILLER_56_12 ();
 sg13g2_fill_2 FILLER_56_18 ();
 sg13g2_fill_2 FILLER_56_25 ();
 sg13g2_fill_1 FILLER_56_76 ();
 sg13g2_fill_1 FILLER_56_86 ();
 sg13g2_fill_1 FILLER_56_93 ();
 sg13g2_fill_1 FILLER_56_104 ();
 sg13g2_fill_1 FILLER_56_122 ();
 sg13g2_fill_1 FILLER_56_135 ();
 sg13g2_fill_1 FILLER_56_141 ();
 sg13g2_fill_1 FILLER_56_147 ();
 sg13g2_fill_2 FILLER_56_152 ();
 sg13g2_fill_2 FILLER_56_158 ();
 sg13g2_fill_2 FILLER_56_165 ();
 sg13g2_fill_2 FILLER_56_232 ();
 sg13g2_fill_1 FILLER_56_239 ();
 sg13g2_fill_1 FILLER_56_290 ();
 sg13g2_fill_1 FILLER_56_295 ();
 sg13g2_fill_1 FILLER_56_306 ();
 sg13g2_decap_8 FILLER_56_311 ();
 sg13g2_fill_2 FILLER_56_318 ();
 sg13g2_fill_1 FILLER_56_320 ();
 sg13g2_fill_2 FILLER_56_329 ();
 sg13g2_fill_1 FILLER_56_361 ();
 sg13g2_fill_1 FILLER_56_367 ();
 sg13g2_fill_1 FILLER_56_373 ();
 sg13g2_fill_1 FILLER_56_390 ();
 sg13g2_fill_2 FILLER_56_400 ();
 sg13g2_fill_2 FILLER_57_47 ();
 sg13g2_fill_2 FILLER_57_74 ();
 sg13g2_fill_1 FILLER_57_99 ();
 sg13g2_fill_1 FILLER_57_105 ();
 sg13g2_fill_2 FILLER_57_123 ();
 sg13g2_fill_1 FILLER_57_134 ();
 sg13g2_fill_2 FILLER_57_140 ();
 sg13g2_fill_2 FILLER_57_146 ();
 sg13g2_fill_2 FILLER_57_158 ();
 sg13g2_fill_1 FILLER_57_160 ();
 sg13g2_fill_2 FILLER_57_214 ();
 sg13g2_decap_4 FILLER_57_230 ();
 sg13g2_fill_1 FILLER_57_234 ();
 sg13g2_fill_1 FILLER_57_262 ();
 sg13g2_fill_1 FILLER_57_268 ();
 sg13g2_fill_2 FILLER_57_297 ();
 sg13g2_fill_2 FILLER_57_306 ();
 sg13g2_decap_4 FILLER_57_322 ();
 sg13g2_fill_2 FILLER_57_326 ();
 sg13g2_fill_1 FILLER_57_333 ();
 sg13g2_fill_1 FILLER_57_381 ();
 sg13g2_fill_1 FILLER_57_387 ();
 sg13g2_fill_2 FILLER_57_393 ();
 sg13g2_fill_1 FILLER_57_395 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_fill_2 FILLER_57_416 ();
 sg13g2_fill_2 FILLER_57_423 ();
 sg13g2_fill_1 FILLER_57_425 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_6 ();
 sg13g2_decap_4 FILLER_58_11 ();
 sg13g2_fill_1 FILLER_58_15 ();
 sg13g2_fill_1 FILLER_58_20 ();
 sg13g2_fill_2 FILLER_58_32 ();
 sg13g2_fill_2 FILLER_58_39 ();
 sg13g2_fill_2 FILLER_58_51 ();
 sg13g2_fill_1 FILLER_58_67 ();
 sg13g2_decap_4 FILLER_58_72 ();
 sg13g2_fill_1 FILLER_58_86 ();
 sg13g2_fill_2 FILLER_58_93 ();
 sg13g2_fill_1 FILLER_58_100 ();
 sg13g2_fill_2 FILLER_58_106 ();
 sg13g2_fill_1 FILLER_58_118 ();
 sg13g2_fill_1 FILLER_58_123 ();
 sg13g2_fill_1 FILLER_58_128 ();
 sg13g2_fill_1 FILLER_58_134 ();
 sg13g2_fill_1 FILLER_58_139 ();
 sg13g2_fill_1 FILLER_58_144 ();
 sg13g2_fill_2 FILLER_58_150 ();
 sg13g2_decap_4 FILLER_58_160 ();
 sg13g2_decap_4 FILLER_58_170 ();
 sg13g2_fill_1 FILLER_58_179 ();
 sg13g2_fill_2 FILLER_58_185 ();
 sg13g2_fill_2 FILLER_58_191 ();
 sg13g2_fill_1 FILLER_58_197 ();
 sg13g2_fill_1 FILLER_58_211 ();
 sg13g2_fill_1 FILLER_58_221 ();
 sg13g2_fill_2 FILLER_58_257 ();
 sg13g2_fill_1 FILLER_58_259 ();
 sg13g2_fill_1 FILLER_58_265 ();
 sg13g2_fill_2 FILLER_58_271 ();
 sg13g2_fill_1 FILLER_58_273 ();
 sg13g2_decap_4 FILLER_58_302 ();
 sg13g2_fill_2 FILLER_58_306 ();
 sg13g2_fill_1 FILLER_58_313 ();
 sg13g2_fill_1 FILLER_58_340 ();
 sg13g2_fill_1 FILLER_58_356 ();
 sg13g2_fill_1 FILLER_58_382 ();
 sg13g2_fill_1 FILLER_58_388 ();
 sg13g2_fill_1 FILLER_58_394 ();
 sg13g2_fill_1 FILLER_58_400 ();
 sg13g2_fill_1 FILLER_58_409 ();
 sg13g2_fill_2 FILLER_58_414 ();
 sg13g2_fill_1 FILLER_58_416 ();
 sg13g2_fill_1 FILLER_59_16 ();
 sg13g2_fill_1 FILLER_59_25 ();
 sg13g2_fill_1 FILLER_59_34 ();
 sg13g2_fill_2 FILLER_59_40 ();
 sg13g2_fill_2 FILLER_59_49 ();
 sg13g2_decap_4 FILLER_59_62 ();
 sg13g2_fill_1 FILLER_59_74 ();
 sg13g2_fill_1 FILLER_59_86 ();
 sg13g2_fill_1 FILLER_59_93 ();
 sg13g2_fill_1 FILLER_59_99 ();
 sg13g2_fill_1 FILLER_59_104 ();
 sg13g2_fill_1 FILLER_59_109 ();
 sg13g2_fill_2 FILLER_59_116 ();
 sg13g2_fill_1 FILLER_59_123 ();
 sg13g2_fill_1 FILLER_59_150 ();
 sg13g2_fill_1 FILLER_59_159 ();
 sg13g2_fill_1 FILLER_59_167 ();
 sg13g2_decap_4 FILLER_59_212 ();
 sg13g2_fill_1 FILLER_59_216 ();
 sg13g2_fill_2 FILLER_59_225 ();
 sg13g2_fill_1 FILLER_59_227 ();
 sg13g2_decap_4 FILLER_59_237 ();
 sg13g2_fill_1 FILLER_59_245 ();
 sg13g2_fill_2 FILLER_59_266 ();
 sg13g2_fill_1 FILLER_59_268 ();
 sg13g2_fill_1 FILLER_59_299 ();
 sg13g2_fill_1 FILLER_59_308 ();
 sg13g2_fill_2 FILLER_59_313 ();
 sg13g2_fill_1 FILLER_59_315 ();
 sg13g2_fill_1 FILLER_59_321 ();
 sg13g2_fill_2 FILLER_59_326 ();
 sg13g2_fill_2 FILLER_59_333 ();
 sg13g2_fill_2 FILLER_59_340 ();
 sg13g2_fill_1 FILLER_59_342 ();
 sg13g2_fill_2 FILLER_59_347 ();
 sg13g2_fill_1 FILLER_59_349 ();
 sg13g2_fill_2 FILLER_59_402 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_15 ();
 sg13g2_fill_2 FILLER_60_33 ();
 sg13g2_fill_1 FILLER_60_39 ();
 sg13g2_fill_1 FILLER_60_55 ();
 sg13g2_fill_2 FILLER_60_68 ();
 sg13g2_fill_1 FILLER_60_70 ();
 sg13g2_decap_4 FILLER_60_80 ();
 sg13g2_fill_2 FILLER_60_114 ();
 sg13g2_fill_1 FILLER_60_116 ();
 sg13g2_fill_2 FILLER_60_130 ();
 sg13g2_fill_1 FILLER_60_140 ();
 sg13g2_fill_1 FILLER_60_145 ();
 sg13g2_fill_2 FILLER_60_150 ();
 sg13g2_fill_1 FILLER_60_177 ();
 sg13g2_fill_1 FILLER_60_182 ();
 sg13g2_decap_4 FILLER_60_188 ();
 sg13g2_fill_1 FILLER_60_192 ();
 sg13g2_fill_2 FILLER_60_207 ();
 sg13g2_fill_1 FILLER_60_209 ();
 sg13g2_decap_4 FILLER_60_218 ();
 sg13g2_fill_2 FILLER_60_266 ();
 sg13g2_fill_1 FILLER_60_268 ();
 sg13g2_fill_2 FILLER_60_280 ();
 sg13g2_fill_2 FILLER_60_307 ();
 sg13g2_fill_1 FILLER_60_309 ();
 sg13g2_fill_2 FILLER_60_314 ();
 sg13g2_fill_2 FILLER_60_321 ();
 sg13g2_fill_2 FILLER_60_327 ();
 sg13g2_fill_2 FILLER_60_339 ();
 sg13g2_fill_1 FILLER_60_341 ();
 sg13g2_fill_1 FILLER_60_347 ();
 sg13g2_fill_1 FILLER_60_352 ();
 sg13g2_fill_1 FILLER_60_386 ();
 sg13g2_fill_1 FILLER_60_398 ();
 sg13g2_fill_2 FILLER_60_406 ();
 sg13g2_fill_2 FILLER_60_414 ();
 sg13g2_fill_2 FILLER_60_420 ();
 sg13g2_decap_4 FILLER_60_426 ();
 sg13g2_decap_4 FILLER_61_13 ();
 sg13g2_fill_2 FILLER_61_17 ();
 sg13g2_fill_2 FILLER_61_28 ();
 sg13g2_fill_2 FILLER_61_34 ();
 sg13g2_decap_4 FILLER_61_61 ();
 sg13g2_fill_2 FILLER_61_71 ();
 sg13g2_fill_1 FILLER_61_73 ();
 sg13g2_fill_1 FILLER_61_79 ();
 sg13g2_decap_4 FILLER_61_100 ();
 sg13g2_fill_2 FILLER_61_104 ();
 sg13g2_fill_2 FILLER_61_118 ();
 sg13g2_fill_2 FILLER_61_138 ();
 sg13g2_fill_1 FILLER_61_145 ();
 sg13g2_fill_1 FILLER_61_154 ();
 sg13g2_fill_1 FILLER_61_162 ();
 sg13g2_fill_1 FILLER_61_168 ();
 sg13g2_fill_1 FILLER_61_174 ();
 sg13g2_fill_1 FILLER_61_201 ();
 sg13g2_fill_2 FILLER_61_228 ();
 sg13g2_fill_1 FILLER_61_234 ();
 sg13g2_fill_1 FILLER_61_240 ();
 sg13g2_fill_2 FILLER_61_267 ();
 sg13g2_fill_1 FILLER_61_269 ();
 sg13g2_fill_1 FILLER_61_286 ();
 sg13g2_fill_1 FILLER_61_299 ();
 sg13g2_fill_1 FILLER_61_345 ();
 sg13g2_fill_1 FILLER_61_351 ();
 sg13g2_fill_2 FILLER_61_362 ();
 sg13g2_fill_2 FILLER_61_428 ();
 sg13g2_fill_1 FILLER_62_5 ();
 sg13g2_fill_1 FILLER_62_12 ();
 sg13g2_fill_2 FILLER_62_42 ();
 sg13g2_fill_1 FILLER_62_44 ();
 sg13g2_fill_2 FILLER_62_81 ();
 sg13g2_fill_2 FILLER_62_113 ();
 sg13g2_fill_1 FILLER_62_124 ();
 sg13g2_fill_1 FILLER_62_168 ();
 sg13g2_fill_1 FILLER_62_191 ();
 sg13g2_fill_2 FILLER_62_200 ();
 sg13g2_fill_2 FILLER_62_237 ();
 sg13g2_fill_2 FILLER_62_266 ();
 sg13g2_fill_1 FILLER_62_290 ();
 sg13g2_fill_2 FILLER_62_314 ();
 sg13g2_fill_2 FILLER_62_328 ();
 sg13g2_fill_1 FILLER_62_330 ();
 sg13g2_fill_1 FILLER_62_350 ();
 sg13g2_fill_2 FILLER_62_358 ();
 sg13g2_fill_1 FILLER_62_365 ();
 sg13g2_fill_1 FILLER_62_375 ();
 sg13g2_decap_4 FILLER_62_421 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_6 ();
 sg13g2_fill_1 FILLER_63_12 ();
 sg13g2_fill_2 FILLER_63_24 ();
 sg13g2_fill_1 FILLER_63_53 ();
 sg13g2_fill_1 FILLER_63_96 ();
 sg13g2_fill_2 FILLER_63_110 ();
 sg13g2_fill_2 FILLER_63_116 ();
 sg13g2_fill_2 FILLER_63_122 ();
 sg13g2_fill_1 FILLER_63_129 ();
 sg13g2_fill_1 FILLER_63_139 ();
 sg13g2_fill_2 FILLER_63_170 ();
 sg13g2_fill_2 FILLER_63_180 ();
 sg13g2_decap_4 FILLER_63_186 ();
 sg13g2_fill_2 FILLER_63_195 ();
 sg13g2_fill_1 FILLER_63_197 ();
 sg13g2_fill_1 FILLER_63_202 ();
 sg13g2_fill_1 FILLER_63_207 ();
 sg13g2_fill_1 FILLER_63_259 ();
 sg13g2_fill_1 FILLER_63_263 ();
 sg13g2_decap_8 FILLER_63_272 ();
 sg13g2_fill_1 FILLER_63_279 ();
 sg13g2_fill_1 FILLER_63_293 ();
 sg13g2_fill_1 FILLER_63_315 ();
 sg13g2_fill_2 FILLER_63_321 ();
 sg13g2_fill_1 FILLER_63_339 ();
 sg13g2_fill_2 FILLER_63_378 ();
 sg13g2_fill_1 FILLER_63_384 ();
 sg13g2_fill_1 FILLER_63_390 ();
 sg13g2_fill_1 FILLER_63_403 ();
 sg13g2_fill_1 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_6 ();
 sg13g2_fill_1 FILLER_64_8 ();
 sg13g2_fill_1 FILLER_64_36 ();
 sg13g2_fill_1 FILLER_64_54 ();
 sg13g2_fill_2 FILLER_64_63 ();
 sg13g2_fill_2 FILLER_64_87 ();
 sg13g2_fill_2 FILLER_64_116 ();
 sg13g2_fill_2 FILLER_64_147 ();
 sg13g2_decap_4 FILLER_64_158 ();
 sg13g2_fill_1 FILLER_64_162 ();
 sg13g2_fill_2 FILLER_64_197 ();
 sg13g2_decap_4 FILLER_64_220 ();
 sg13g2_decap_4 FILLER_64_266 ();
 sg13g2_fill_2 FILLER_64_274 ();
 sg13g2_fill_1 FILLER_64_276 ();
 sg13g2_fill_1 FILLER_64_281 ();
 sg13g2_decap_4 FILLER_64_312 ();
 sg13g2_fill_1 FILLER_64_321 ();
 sg13g2_decap_4 FILLER_64_326 ();
 sg13g2_fill_1 FILLER_64_330 ();
 sg13g2_fill_1 FILLER_64_336 ();
 sg13g2_fill_1 FILLER_64_341 ();
 sg13g2_fill_2 FILLER_64_347 ();
 sg13g2_fill_1 FILLER_64_354 ();
 sg13g2_fill_2 FILLER_64_384 ();
 sg13g2_fill_1 FILLER_64_393 ();
 sg13g2_fill_1 FILLER_64_402 ();
 sg13g2_fill_2 FILLER_64_415 ();
 sg13g2_fill_1 FILLER_64_417 ();
 sg13g2_fill_2 FILLER_64_422 ();
 sg13g2_fill_1 FILLER_64_424 ();
 sg13g2_fill_1 FILLER_64_429 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_12 ();
 sg13g2_fill_1 FILLER_65_14 ();
 sg13g2_fill_1 FILLER_65_57 ();
 sg13g2_fill_1 FILLER_65_74 ();
 sg13g2_fill_2 FILLER_65_153 ();
 sg13g2_fill_1 FILLER_65_164 ();
 sg13g2_decap_4 FILLER_65_175 ();
 sg13g2_fill_1 FILLER_65_187 ();
 sg13g2_fill_1 FILLER_65_193 ();
 sg13g2_decap_8 FILLER_65_236 ();
 sg13g2_decap_4 FILLER_65_243 ();
 sg13g2_fill_2 FILLER_65_255 ();
 sg13g2_decap_4 FILLER_65_266 ();
 sg13g2_decap_4 FILLER_65_274 ();
 sg13g2_fill_1 FILLER_65_278 ();
 sg13g2_fill_2 FILLER_65_296 ();
 sg13g2_fill_1 FILLER_65_328 ();
 sg13g2_fill_2 FILLER_65_337 ();
 sg13g2_fill_1 FILLER_65_364 ();
 sg13g2_fill_2 FILLER_65_373 ();
 sg13g2_fill_2 FILLER_65_398 ();
 sg13g2_fill_1 FILLER_65_406 ();
 sg13g2_fill_1 FILLER_65_414 ();
 sg13g2_fill_2 FILLER_65_419 ();
 sg13g2_fill_2 FILLER_65_427 ();
 sg13g2_fill_1 FILLER_65_429 ();
 sg13g2_fill_1 FILLER_66_47 ();
 sg13g2_fill_1 FILLER_66_54 ();
 sg13g2_fill_1 FILLER_66_60 ();
 sg13g2_fill_1 FILLER_66_66 ();
 sg13g2_fill_2 FILLER_66_80 ();
 sg13g2_fill_2 FILLER_66_92 ();
 sg13g2_fill_1 FILLER_66_94 ();
 sg13g2_fill_2 FILLER_66_99 ();
 sg13g2_fill_1 FILLER_66_101 ();
 sg13g2_fill_2 FILLER_66_106 ();
 sg13g2_fill_1 FILLER_66_108 ();
 sg13g2_decap_4 FILLER_66_125 ();
 sg13g2_fill_1 FILLER_66_129 ();
 sg13g2_fill_1 FILLER_66_139 ();
 sg13g2_fill_1 FILLER_66_157 ();
 sg13g2_decap_4 FILLER_66_167 ();
 sg13g2_fill_1 FILLER_66_181 ();
 sg13g2_fill_1 FILLER_66_195 ();
 sg13g2_fill_1 FILLER_66_204 ();
 sg13g2_fill_2 FILLER_66_209 ();
 sg13g2_fill_2 FILLER_66_248 ();
 sg13g2_fill_2 FILLER_66_289 ();
 sg13g2_decap_8 FILLER_66_322 ();
 sg13g2_fill_1 FILLER_66_329 ();
 sg13g2_fill_1 FILLER_66_361 ();
 sg13g2_fill_2 FILLER_66_367 ();
 sg13g2_fill_1 FILLER_66_369 ();
 sg13g2_fill_1 FILLER_66_377 ();
 sg13g2_fill_1 FILLER_66_390 ();
 sg13g2_fill_2 FILLER_66_402 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_42 ();
 sg13g2_fill_1 FILLER_67_50 ();
 sg13g2_fill_1 FILLER_67_77 ();
 sg13g2_fill_1 FILLER_67_84 ();
 sg13g2_fill_2 FILLER_67_111 ();
 sg13g2_fill_1 FILLER_67_118 ();
 sg13g2_fill_1 FILLER_67_137 ();
 sg13g2_fill_2 FILLER_67_159 ();
 sg13g2_fill_1 FILLER_67_217 ();
 sg13g2_fill_1 FILLER_67_222 ();
 sg13g2_fill_2 FILLER_67_227 ();
 sg13g2_fill_1 FILLER_67_229 ();
 sg13g2_fill_1 FILLER_67_234 ();
 sg13g2_decap_4 FILLER_67_239 ();
 sg13g2_fill_1 FILLER_67_243 ();
 sg13g2_fill_2 FILLER_67_254 ();
 sg13g2_fill_1 FILLER_67_256 ();
 sg13g2_fill_2 FILLER_67_261 ();
 sg13g2_fill_1 FILLER_67_263 ();
 sg13g2_fill_2 FILLER_67_272 ();
 sg13g2_fill_1 FILLER_67_274 ();
 sg13g2_fill_2 FILLER_67_280 ();
 sg13g2_fill_1 FILLER_67_287 ();
 sg13g2_fill_1 FILLER_67_293 ();
 sg13g2_fill_1 FILLER_67_300 ();
 sg13g2_fill_2 FILLER_67_320 ();
 sg13g2_decap_4 FILLER_67_330 ();
 sg13g2_fill_1 FILLER_67_380 ();
 sg13g2_fill_2 FILLER_67_404 ();
 sg13g2_fill_2 FILLER_67_421 ();
 sg13g2_fill_2 FILLER_67_427 ();
 sg13g2_fill_1 FILLER_67_429 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_40 ();
 sg13g2_fill_1 FILLER_68_51 ();
 sg13g2_fill_1 FILLER_68_57 ();
 sg13g2_decap_4 FILLER_68_70 ();
 sg13g2_decap_4 FILLER_68_78 ();
 sg13g2_fill_2 FILLER_68_82 ();
 sg13g2_fill_2 FILLER_68_88 ();
 sg13g2_fill_1 FILLER_68_121 ();
 sg13g2_fill_1 FILLER_68_127 ();
 sg13g2_fill_1 FILLER_68_177 ();
 sg13g2_fill_2 FILLER_68_182 ();
 sg13g2_fill_1 FILLER_68_184 ();
 sg13g2_fill_2 FILLER_68_193 ();
 sg13g2_decap_8 FILLER_68_203 ();
 sg13g2_fill_1 FILLER_68_215 ();
 sg13g2_fill_1 FILLER_68_242 ();
 sg13g2_fill_1 FILLER_68_248 ();
 sg13g2_fill_1 FILLER_68_254 ();
 sg13g2_fill_2 FILLER_68_303 ();
 sg13g2_fill_1 FILLER_68_311 ();
 sg13g2_fill_2 FILLER_68_318 ();
 sg13g2_fill_1 FILLER_68_320 ();
 sg13g2_fill_2 FILLER_68_401 ();
 sg13g2_fill_1 FILLER_68_403 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_10 ();
 sg13g2_decap_4 FILLER_69_16 ();
 sg13g2_fill_2 FILLER_69_20 ();
 sg13g2_decap_8 FILLER_69_27 ();
 sg13g2_fill_1 FILLER_69_34 ();
 sg13g2_fill_2 FILLER_69_44 ();
 sg13g2_fill_2 FILLER_69_51 ();
 sg13g2_fill_2 FILLER_69_73 ();
 sg13g2_fill_2 FILLER_69_80 ();
 sg13g2_fill_1 FILLER_69_82 ();
 sg13g2_fill_2 FILLER_69_105 ();
 sg13g2_fill_2 FILLER_69_117 ();
 sg13g2_fill_2 FILLER_69_146 ();
 sg13g2_fill_1 FILLER_69_148 ();
 sg13g2_fill_2 FILLER_69_209 ();
 sg13g2_fill_1 FILLER_69_216 ();
 sg13g2_fill_1 FILLER_69_222 ();
 sg13g2_fill_1 FILLER_69_227 ();
 sg13g2_fill_1 FILLER_69_236 ();
 sg13g2_decap_4 FILLER_69_241 ();
 sg13g2_fill_2 FILLER_69_245 ();
 sg13g2_fill_2 FILLER_69_252 ();
 sg13g2_fill_1 FILLER_69_254 ();
 sg13g2_fill_2 FILLER_69_259 ();
 sg13g2_decap_4 FILLER_69_346 ();
 sg13g2_fill_1 FILLER_69_350 ();
 sg13g2_fill_1 FILLER_69_363 ();
 sg13g2_fill_1 FILLER_69_388 ();
 sg13g2_fill_1 FILLER_69_425 ();
 sg13g2_fill_1 FILLER_70_31 ();
 sg13g2_fill_1 FILLER_70_44 ();
 sg13g2_fill_2 FILLER_70_55 ();
 sg13g2_fill_1 FILLER_70_57 ();
 sg13g2_fill_2 FILLER_70_62 ();
 sg13g2_decap_8 FILLER_70_80 ();
 sg13g2_decap_8 FILLER_70_87 ();
 sg13g2_decap_4 FILLER_70_94 ();
 sg13g2_fill_2 FILLER_70_98 ();
 sg13g2_fill_1 FILLER_70_111 ();
 sg13g2_fill_2 FILLER_70_127 ();
 sg13g2_fill_2 FILLER_70_184 ();
 sg13g2_fill_1 FILLER_70_186 ();
 sg13g2_fill_2 FILLER_70_202 ();
 sg13g2_fill_1 FILLER_70_208 ();
 sg13g2_fill_2 FILLER_70_267 ();
 sg13g2_fill_1 FILLER_70_269 ();
 sg13g2_fill_1 FILLER_70_283 ();
 sg13g2_decap_4 FILLER_70_301 ();
 sg13g2_fill_2 FILLER_70_333 ();
 sg13g2_fill_1 FILLER_70_371 ();
 sg13g2_decap_8 FILLER_70_421 ();
 sg13g2_fill_2 FILLER_70_428 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_4 FILLER_71_15 ();
 sg13g2_fill_1 FILLER_71_19 ();
 sg13g2_fill_2 FILLER_71_60 ();
 sg13g2_decap_4 FILLER_71_67 ();
 sg13g2_decap_4 FILLER_71_103 ();
 sg13g2_fill_1 FILLER_71_118 ();
 sg13g2_fill_2 FILLER_71_127 ();
 sg13g2_fill_1 FILLER_71_134 ();
 sg13g2_decap_4 FILLER_71_154 ();
 sg13g2_fill_1 FILLER_71_158 ();
 sg13g2_fill_1 FILLER_71_164 ();
 sg13g2_fill_2 FILLER_71_183 ();
 sg13g2_fill_1 FILLER_71_185 ();
 sg13g2_fill_1 FILLER_71_208 ();
 sg13g2_fill_1 FILLER_71_214 ();
 sg13g2_decap_4 FILLER_71_269 ();
 sg13g2_fill_1 FILLER_71_278 ();
 sg13g2_fill_1 FILLER_71_283 ();
 sg13g2_fill_2 FILLER_71_288 ();
 sg13g2_fill_1 FILLER_71_307 ();
 sg13g2_fill_2 FILLER_71_346 ();
 sg13g2_fill_1 FILLER_71_391 ();
 sg13g2_decap_8 FILLER_71_422 ();
 sg13g2_fill_1 FILLER_71_429 ();
 sg13g2_fill_1 FILLER_72_43 ();
 sg13g2_fill_1 FILLER_72_52 ();
 sg13g2_fill_1 FILLER_72_58 ();
 sg13g2_fill_2 FILLER_72_69 ();
 sg13g2_fill_1 FILLER_72_79 ();
 sg13g2_fill_2 FILLER_72_94 ();
 sg13g2_fill_2 FILLER_72_104 ();
 sg13g2_fill_2 FILLER_72_111 ();
 sg13g2_decap_4 FILLER_72_117 ();
 sg13g2_fill_2 FILLER_72_144 ();
 sg13g2_fill_1 FILLER_72_151 ();
 sg13g2_fill_2 FILLER_72_156 ();
 sg13g2_fill_1 FILLER_72_158 ();
 sg13g2_fill_2 FILLER_72_184 ();
 sg13g2_decap_8 FILLER_72_190 ();
 sg13g2_fill_2 FILLER_72_205 ();
 sg13g2_fill_2 FILLER_72_241 ();
 sg13g2_fill_1 FILLER_72_243 ();
 sg13g2_decap_8 FILLER_72_305 ();
 sg13g2_fill_2 FILLER_72_320 ();
 sg13g2_decap_4 FILLER_72_344 ();
 sg13g2_fill_2 FILLER_72_358 ();
 sg13g2_fill_1 FILLER_72_398 ();
 sg13g2_fill_2 FILLER_72_404 ();
 sg13g2_fill_2 FILLER_72_427 ();
 sg13g2_fill_1 FILLER_72_429 ();
 sg13g2_decap_4 FILLER_73_42 ();
 sg13g2_fill_2 FILLER_73_101 ();
 sg13g2_decap_4 FILLER_73_123 ();
 sg13g2_fill_1 FILLER_73_127 ();
 sg13g2_fill_2 FILLER_73_176 ();
 sg13g2_fill_1 FILLER_73_178 ();
 sg13g2_fill_2 FILLER_73_200 ();
 sg13g2_fill_2 FILLER_73_212 ();
 sg13g2_fill_1 FILLER_73_240 ();
 sg13g2_fill_1 FILLER_73_246 ();
 sg13g2_fill_1 FILLER_73_251 ();
 sg13g2_fill_2 FILLER_73_261 ();
 sg13g2_fill_1 FILLER_73_263 ();
 sg13g2_fill_1 FILLER_73_292 ();
 sg13g2_fill_1 FILLER_73_306 ();
 sg13g2_fill_1 FILLER_73_312 ();
 sg13g2_fill_2 FILLER_73_317 ();
 sg13g2_fill_1 FILLER_73_332 ();
 sg13g2_fill_1 FILLER_73_352 ();
 sg13g2_fill_1 FILLER_73_358 ();
 sg13g2_fill_1 FILLER_73_372 ();
 sg13g2_fill_1 FILLER_73_378 ();
 sg13g2_fill_1 FILLER_73_385 ();
 sg13g2_fill_1 FILLER_73_391 ();
 sg13g2_fill_1 FILLER_73_396 ();
 sg13g2_fill_1 FILLER_73_403 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_27 ();
 sg13g2_fill_2 FILLER_74_34 ();
 sg13g2_fill_2 FILLER_74_56 ();
 sg13g2_fill_2 FILLER_74_77 ();
 sg13g2_decap_4 FILLER_74_86 ();
 sg13g2_fill_1 FILLER_74_90 ();
 sg13g2_fill_2 FILLER_74_95 ();
 sg13g2_fill_1 FILLER_74_97 ();
 sg13g2_fill_1 FILLER_74_128 ();
 sg13g2_fill_1 FILLER_74_160 ();
 sg13g2_fill_2 FILLER_74_166 ();
 sg13g2_fill_1 FILLER_74_194 ();
 sg13g2_decap_8 FILLER_74_220 ();
 sg13g2_decap_8 FILLER_74_287 ();
 sg13g2_fill_1 FILLER_74_327 ();
 sg13g2_fill_1 FILLER_74_337 ();
 sg13g2_fill_1 FILLER_74_348 ();
 sg13g2_fill_2 FILLER_74_381 ();
 sg13g2_fill_2 FILLER_74_387 ();
 sg13g2_fill_1 FILLER_74_389 ();
 sg13g2_fill_1 FILLER_74_402 ();
 sg13g2_fill_1 FILLER_74_411 ();
 sg13g2_fill_2 FILLER_74_427 ();
 sg13g2_fill_1 FILLER_74_429 ();
 sg13g2_fill_1 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_5 ();
 sg13g2_fill_1 FILLER_75_20 ();
 sg13g2_fill_2 FILLER_75_26 ();
 sg13g2_fill_2 FILLER_75_32 ();
 sg13g2_fill_2 FILLER_75_39 ();
 sg13g2_fill_1 FILLER_75_53 ();
 sg13g2_fill_2 FILLER_75_58 ();
 sg13g2_fill_1 FILLER_75_68 ();
 sg13g2_fill_1 FILLER_75_77 ();
 sg13g2_decap_4 FILLER_75_113 ();
 sg13g2_fill_1 FILLER_75_117 ();
 sg13g2_fill_1 FILLER_75_122 ();
 sg13g2_fill_1 FILLER_75_135 ();
 sg13g2_fill_2 FILLER_75_143 ();
 sg13g2_fill_2 FILLER_75_149 ();
 sg13g2_fill_1 FILLER_75_151 ();
 sg13g2_fill_1 FILLER_75_178 ();
 sg13g2_fill_2 FILLER_75_184 ();
 sg13g2_fill_1 FILLER_75_191 ();
 sg13g2_fill_2 FILLER_75_197 ();
 sg13g2_decap_4 FILLER_75_210 ();
 sg13g2_fill_1 FILLER_75_235 ();
 sg13g2_fill_1 FILLER_75_242 ();
 sg13g2_fill_1 FILLER_75_275 ();
 sg13g2_fill_2 FILLER_75_307 ();
 sg13g2_fill_1 FILLER_75_314 ();
 sg13g2_fill_1 FILLER_75_357 ();
 sg13g2_fill_1 FILLER_75_363 ();
 sg13g2_fill_2 FILLER_75_372 ();
 sg13g2_fill_1 FILLER_75_379 ();
 sg13g2_fill_1 FILLER_75_388 ();
 sg13g2_fill_2 FILLER_75_401 ();
 sg13g2_fill_1 FILLER_75_403 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_11 ();
 sg13g2_fill_2 FILLER_76_18 ();
 sg13g2_fill_1 FILLER_76_20 ();
 sg13g2_fill_1 FILLER_76_45 ();
 sg13g2_fill_1 FILLER_76_62 ();
 sg13g2_fill_2 FILLER_76_72 ();
 sg13g2_fill_1 FILLER_76_124 ();
 sg13g2_fill_1 FILLER_76_169 ();
 sg13g2_fill_1 FILLER_76_191 ();
 sg13g2_fill_2 FILLER_76_197 ();
 sg13g2_fill_1 FILLER_76_199 ();
 sg13g2_fill_2 FILLER_76_205 ();
 sg13g2_fill_1 FILLER_76_237 ();
 sg13g2_decap_4 FILLER_76_268 ();
 sg13g2_fill_1 FILLER_76_272 ();
 sg13g2_fill_1 FILLER_76_277 ();
 sg13g2_fill_2 FILLER_76_282 ();
 sg13g2_fill_2 FILLER_76_288 ();
 sg13g2_fill_2 FILLER_76_295 ();
 sg13g2_fill_1 FILLER_76_311 ();
 sg13g2_fill_2 FILLER_76_336 ();
 sg13g2_fill_2 FILLER_76_343 ();
 sg13g2_fill_1 FILLER_76_376 ();
 sg13g2_fill_2 FILLER_76_385 ();
 sg13g2_fill_1 FILLER_76_387 ();
 sg13g2_fill_2 FILLER_76_427 ();
 sg13g2_fill_1 FILLER_76_429 ();
 sg13g2_decap_4 FILLER_77_26 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_fill_1 FILLER_77_49 ();
 sg13g2_fill_2 FILLER_77_62 ();
 sg13g2_fill_1 FILLER_77_64 ();
 sg13g2_decap_4 FILLER_77_72 ();
 sg13g2_fill_2 FILLER_77_85 ();
 sg13g2_decap_4 FILLER_77_117 ();
 sg13g2_decap_8 FILLER_77_135 ();
 sg13g2_fill_2 FILLER_77_142 ();
 sg13g2_fill_2 FILLER_77_153 ();
 sg13g2_fill_1 FILLER_77_155 ();
 sg13g2_fill_1 FILLER_77_160 ();
 sg13g2_fill_2 FILLER_77_168 ();
 sg13g2_fill_1 FILLER_77_210 ();
 sg13g2_fill_2 FILLER_77_214 ();
 sg13g2_fill_1 FILLER_77_220 ();
 sg13g2_fill_2 FILLER_77_229 ();
 sg13g2_fill_1 FILLER_77_237 ();
 sg13g2_fill_2 FILLER_77_242 ();
 sg13g2_fill_2 FILLER_77_258 ();
 sg13g2_fill_1 FILLER_77_260 ();
 sg13g2_decap_8 FILLER_77_266 ();
 sg13g2_fill_2 FILLER_77_273 ();
 sg13g2_fill_2 FILLER_77_336 ();
 sg13g2_fill_1 FILLER_77_344 ();
 sg13g2_fill_2 FILLER_77_377 ();
 sg13g2_fill_1 FILLER_77_383 ();
 sg13g2_fill_1 FILLER_77_394 ();
 sg13g2_fill_2 FILLER_77_414 ();
 sg13g2_fill_1 FILLER_77_416 ();
 sg13g2_fill_2 FILLER_77_428 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_31 ();
 sg13g2_fill_1 FILLER_78_43 ();
 sg13g2_fill_1 FILLER_78_49 ();
 sg13g2_fill_1 FILLER_78_55 ();
 sg13g2_fill_1 FILLER_78_60 ();
 sg13g2_fill_1 FILLER_78_66 ();
 sg13g2_decap_4 FILLER_78_72 ();
 sg13g2_fill_2 FILLER_78_76 ();
 sg13g2_fill_1 FILLER_78_100 ();
 sg13g2_fill_2 FILLER_78_106 ();
 sg13g2_decap_4 FILLER_78_118 ();
 sg13g2_fill_1 FILLER_78_153 ();
 sg13g2_fill_1 FILLER_78_210 ();
 sg13g2_fill_1 FILLER_78_249 ();
 sg13g2_fill_2 FILLER_78_402 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_4 FILLER_79_14 ();
 sg13g2_fill_1 FILLER_79_18 ();
 sg13g2_fill_1 FILLER_79_45 ();
 sg13g2_decap_8 FILLER_79_102 ();
 sg13g2_fill_1 FILLER_79_113 ();
 sg13g2_fill_2 FILLER_79_144 ();
 sg13g2_fill_1 FILLER_79_146 ();
 sg13g2_fill_1 FILLER_79_171 ();
 sg13g2_fill_1 FILLER_79_176 ();
 sg13g2_fill_1 FILLER_79_185 ();
 sg13g2_fill_2 FILLER_79_296 ();
 sg13g2_fill_1 FILLER_79_302 ();
 sg13g2_fill_2 FILLER_79_350 ();
 sg13g2_fill_1 FILLER_79_365 ();
 sg13g2_fill_2 FILLER_79_388 ();
 sg13g2_fill_1 FILLER_79_390 ();
 sg13g2_fill_1 FILLER_79_396 ();
 sg13g2_fill_2 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_4 FILLER_80_14 ();
 sg13g2_fill_2 FILLER_80_18 ();
 sg13g2_fill_1 FILLER_80_73 ();
 sg13g2_fill_1 FILLER_80_79 ();
 sg13g2_fill_2 FILLER_80_174 ();
 sg13g2_fill_1 FILLER_80_176 ();
 sg13g2_fill_1 FILLER_80_288 ();
 sg13g2_fill_1 FILLER_80_332 ();
 sg13g2_fill_1 FILLER_80_371 ();
 sg13g2_fill_1 FILLER_80_376 ();
 sg13g2_fill_1 FILLER_80_403 ();
 sg13g2_fill_2 FILLER_80_420 ();
 sg13g2_fill_1 FILLER_80_422 ();
 sg13g2_fill_2 FILLER_80_427 ();
 sg13g2_fill_1 FILLER_80_429 ();
endmodule
