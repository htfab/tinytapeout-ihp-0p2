module tt_um_froith_goldcrest (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire clknet_leaf_0_clk;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire net2016;
 wire _13604_;
 wire _13605_;
 wire \top_ihp.gpio_o_1 ;
 wire \top_ihp.gpio_o_2 ;
 wire \top_ihp.gpio_o_3 ;
 wire \top_ihp.gpio_o_4 ;
 wire \top_ihp.oisc.decoder.decoded[0] ;
 wire \top_ihp.oisc.decoder.decoded[10] ;
 wire \top_ihp.oisc.decoder.decoded[11] ;
 wire \top_ihp.oisc.decoder.decoded[12] ;
 wire \top_ihp.oisc.decoder.decoded[13] ;
 wire \top_ihp.oisc.decoder.decoded[14] ;
 wire \top_ihp.oisc.decoder.decoded[15] ;
 wire \top_ihp.oisc.decoder.decoded[1] ;
 wire \top_ihp.oisc.decoder.decoded[2] ;
 wire \top_ihp.oisc.decoder.decoded[3] ;
 wire \top_ihp.oisc.decoder.decoded[4] ;
 wire \top_ihp.oisc.decoder.decoded[5] ;
 wire \top_ihp.oisc.decoder.decoded[6] ;
 wire \top_ihp.oisc.decoder.decoded[7] ;
 wire \top_ihp.oisc.decoder.instruction[10] ;
 wire \top_ihp.oisc.decoder.instruction[11] ;
 wire \top_ihp.oisc.decoder.instruction[12] ;
 wire \top_ihp.oisc.decoder.instruction[13] ;
 wire \top_ihp.oisc.decoder.instruction[14] ;
 wire \top_ihp.oisc.decoder.instruction[15] ;
 wire \top_ihp.oisc.decoder.instruction[16] ;
 wire \top_ihp.oisc.decoder.instruction[17] ;
 wire \top_ihp.oisc.decoder.instruction[18] ;
 wire \top_ihp.oisc.decoder.instruction[19] ;
 wire \top_ihp.oisc.decoder.instruction[20] ;
 wire \top_ihp.oisc.decoder.instruction[21] ;
 wire \top_ihp.oisc.decoder.instruction[22] ;
 wire \top_ihp.oisc.decoder.instruction[23] ;
 wire \top_ihp.oisc.decoder.instruction[24] ;
 wire \top_ihp.oisc.decoder.instruction[25] ;
 wire \top_ihp.oisc.decoder.instruction[26] ;
 wire \top_ihp.oisc.decoder.instruction[27] ;
 wire \top_ihp.oisc.decoder.instruction[28] ;
 wire \top_ihp.oisc.decoder.instruction[29] ;
 wire \top_ihp.oisc.decoder.instruction[30] ;
 wire \top_ihp.oisc.decoder.instruction[31] ;
 wire \top_ihp.oisc.decoder.instruction[7] ;
 wire \top_ihp.oisc.decoder.instruction[8] ;
 wire \top_ihp.oisc.decoder.instruction[9] ;
 wire \top_ihp.oisc.mem_addr_lowbits[0] ;
 wire \top_ihp.oisc.mem_addr_lowbits[1] ;
 wire \top_ihp.oisc.micro_op[0] ;
 wire \top_ihp.oisc.micro_op[10] ;
 wire \top_ihp.oisc.micro_op[11] ;
 wire \top_ihp.oisc.micro_op[12] ;
 wire \top_ihp.oisc.micro_op[13] ;
 wire \top_ihp.oisc.micro_op[14] ;
 wire \top_ihp.oisc.micro_op[15] ;
 wire \top_ihp.oisc.micro_op[1] ;
 wire \top_ihp.oisc.micro_op[2] ;
 wire \top_ihp.oisc.micro_op[3] ;
 wire \top_ihp.oisc.micro_op[4] ;
 wire \top_ihp.oisc.micro_op[5] ;
 wire \top_ihp.oisc.micro_op[8] ;
 wire \top_ihp.oisc.micro_op[9] ;
 wire \top_ihp.oisc.micro_pc[0] ;
 wire \top_ihp.oisc.micro_pc[1] ;
 wire \top_ihp.oisc.micro_pc[2] ;
 wire \top_ihp.oisc.micro_pc[3] ;
 wire \top_ihp.oisc.micro_pc[4] ;
 wire \top_ihp.oisc.micro_pc[5] ;
 wire \top_ihp.oisc.micro_pc[6] ;
 wire \top_ihp.oisc.micro_pc[7] ;
 wire \top_ihp.oisc.micro_res_addr[0] ;
 wire \top_ihp.oisc.micro_res_addr[1] ;
 wire \top_ihp.oisc.micro_res_addr[2] ;
 wire \top_ihp.oisc.micro_res_addr[3] ;
 wire \top_ihp.oisc.micro_state[0] ;
 wire \top_ihp.oisc.micro_state[1] ;
 wire \top_ihp.oisc.micro_state[2] ;
 wire \top_ihp.oisc.op_a[0] ;
 wire \top_ihp.oisc.op_a[10] ;
 wire \top_ihp.oisc.op_a[11] ;
 wire \top_ihp.oisc.op_a[12] ;
 wire \top_ihp.oisc.op_a[13] ;
 wire \top_ihp.oisc.op_a[14] ;
 wire \top_ihp.oisc.op_a[15] ;
 wire \top_ihp.oisc.op_a[16] ;
 wire \top_ihp.oisc.op_a[17] ;
 wire \top_ihp.oisc.op_a[18] ;
 wire \top_ihp.oisc.op_a[19] ;
 wire \top_ihp.oisc.op_a[1] ;
 wire \top_ihp.oisc.op_a[20] ;
 wire \top_ihp.oisc.op_a[21] ;
 wire \top_ihp.oisc.op_a[22] ;
 wire \top_ihp.oisc.op_a[23] ;
 wire \top_ihp.oisc.op_a[24] ;
 wire \top_ihp.oisc.op_a[25] ;
 wire \top_ihp.oisc.op_a[26] ;
 wire \top_ihp.oisc.op_a[27] ;
 wire \top_ihp.oisc.op_a[28] ;
 wire \top_ihp.oisc.op_a[29] ;
 wire \top_ihp.oisc.op_a[2] ;
 wire \top_ihp.oisc.op_a[30] ;
 wire \top_ihp.oisc.op_a[31] ;
 wire \top_ihp.oisc.op_a[3] ;
 wire \top_ihp.oisc.op_a[4] ;
 wire \top_ihp.oisc.op_a[5] ;
 wire \top_ihp.oisc.op_a[6] ;
 wire \top_ihp.oisc.op_a[7] ;
 wire \top_ihp.oisc.op_a[8] ;
 wire \top_ihp.oisc.op_a[9] ;
 wire \top_ihp.oisc.op_b[0] ;
 wire \top_ihp.oisc.op_b[10] ;
 wire \top_ihp.oisc.op_b[11] ;
 wire \top_ihp.oisc.op_b[12] ;
 wire \top_ihp.oisc.op_b[13] ;
 wire \top_ihp.oisc.op_b[14] ;
 wire \top_ihp.oisc.op_b[15] ;
 wire \top_ihp.oisc.op_b[16] ;
 wire \top_ihp.oisc.op_b[17] ;
 wire \top_ihp.oisc.op_b[18] ;
 wire \top_ihp.oisc.op_b[19] ;
 wire \top_ihp.oisc.op_b[1] ;
 wire \top_ihp.oisc.op_b[20] ;
 wire \top_ihp.oisc.op_b[21] ;
 wire \top_ihp.oisc.op_b[22] ;
 wire \top_ihp.oisc.op_b[23] ;
 wire \top_ihp.oisc.op_b[24] ;
 wire \top_ihp.oisc.op_b[25] ;
 wire \top_ihp.oisc.op_b[26] ;
 wire \top_ihp.oisc.op_b[27] ;
 wire \top_ihp.oisc.op_b[28] ;
 wire \top_ihp.oisc.op_b[29] ;
 wire \top_ihp.oisc.op_b[2] ;
 wire \top_ihp.oisc.op_b[30] ;
 wire \top_ihp.oisc.op_b[31] ;
 wire \top_ihp.oisc.op_b[3] ;
 wire \top_ihp.oisc.op_b[4] ;
 wire \top_ihp.oisc.op_b[5] ;
 wire \top_ihp.oisc.op_b[6] ;
 wire \top_ihp.oisc.op_b[7] ;
 wire \top_ihp.oisc.op_b[8] ;
 wire \top_ihp.oisc.op_b[9] ;
 wire \top_ihp.oisc.reg_rb[0] ;
 wire \top_ihp.oisc.reg_rb[1] ;
 wire \top_ihp.oisc.reg_rb[2] ;
 wire \top_ihp.oisc.reg_rb[3] ;
 wire \top_ihp.oisc.regs[0][0] ;
 wire \top_ihp.oisc.regs[0][10] ;
 wire \top_ihp.oisc.regs[0][11] ;
 wire \top_ihp.oisc.regs[0][12] ;
 wire \top_ihp.oisc.regs[0][13] ;
 wire \top_ihp.oisc.regs[0][14] ;
 wire \top_ihp.oisc.regs[0][15] ;
 wire \top_ihp.oisc.regs[0][16] ;
 wire \top_ihp.oisc.regs[0][17] ;
 wire \top_ihp.oisc.regs[0][18] ;
 wire \top_ihp.oisc.regs[0][19] ;
 wire \top_ihp.oisc.regs[0][1] ;
 wire \top_ihp.oisc.regs[0][20] ;
 wire \top_ihp.oisc.regs[0][21] ;
 wire \top_ihp.oisc.regs[0][22] ;
 wire \top_ihp.oisc.regs[0][23] ;
 wire \top_ihp.oisc.regs[0][24] ;
 wire \top_ihp.oisc.regs[0][25] ;
 wire \top_ihp.oisc.regs[0][26] ;
 wire \top_ihp.oisc.regs[0][27] ;
 wire \top_ihp.oisc.regs[0][28] ;
 wire \top_ihp.oisc.regs[0][29] ;
 wire \top_ihp.oisc.regs[0][2] ;
 wire \top_ihp.oisc.regs[0][30] ;
 wire \top_ihp.oisc.regs[0][31] ;
 wire \top_ihp.oisc.regs[0][3] ;
 wire \top_ihp.oisc.regs[0][4] ;
 wire \top_ihp.oisc.regs[0][5] ;
 wire \top_ihp.oisc.regs[0][6] ;
 wire \top_ihp.oisc.regs[0][7] ;
 wire \top_ihp.oisc.regs[0][8] ;
 wire \top_ihp.oisc.regs[0][9] ;
 wire \top_ihp.oisc.regs[10][0] ;
 wire \top_ihp.oisc.regs[10][10] ;
 wire \top_ihp.oisc.regs[10][11] ;
 wire \top_ihp.oisc.regs[10][12] ;
 wire \top_ihp.oisc.regs[10][13] ;
 wire \top_ihp.oisc.regs[10][14] ;
 wire \top_ihp.oisc.regs[10][15] ;
 wire \top_ihp.oisc.regs[10][16] ;
 wire \top_ihp.oisc.regs[10][17] ;
 wire \top_ihp.oisc.regs[10][18] ;
 wire \top_ihp.oisc.regs[10][19] ;
 wire \top_ihp.oisc.regs[10][1] ;
 wire \top_ihp.oisc.regs[10][20] ;
 wire \top_ihp.oisc.regs[10][21] ;
 wire \top_ihp.oisc.regs[10][22] ;
 wire \top_ihp.oisc.regs[10][23] ;
 wire \top_ihp.oisc.regs[10][24] ;
 wire \top_ihp.oisc.regs[10][25] ;
 wire \top_ihp.oisc.regs[10][26] ;
 wire \top_ihp.oisc.regs[10][27] ;
 wire \top_ihp.oisc.regs[10][28] ;
 wire \top_ihp.oisc.regs[10][29] ;
 wire \top_ihp.oisc.regs[10][2] ;
 wire \top_ihp.oisc.regs[10][30] ;
 wire \top_ihp.oisc.regs[10][31] ;
 wire \top_ihp.oisc.regs[10][3] ;
 wire \top_ihp.oisc.regs[10][4] ;
 wire \top_ihp.oisc.regs[10][5] ;
 wire \top_ihp.oisc.regs[10][6] ;
 wire \top_ihp.oisc.regs[10][7] ;
 wire \top_ihp.oisc.regs[10][8] ;
 wire \top_ihp.oisc.regs[10][9] ;
 wire \top_ihp.oisc.regs[11][0] ;
 wire \top_ihp.oisc.regs[11][10] ;
 wire \top_ihp.oisc.regs[11][11] ;
 wire \top_ihp.oisc.regs[11][12] ;
 wire \top_ihp.oisc.regs[11][13] ;
 wire \top_ihp.oisc.regs[11][14] ;
 wire \top_ihp.oisc.regs[11][15] ;
 wire \top_ihp.oisc.regs[11][16] ;
 wire \top_ihp.oisc.regs[11][17] ;
 wire \top_ihp.oisc.regs[11][18] ;
 wire \top_ihp.oisc.regs[11][19] ;
 wire \top_ihp.oisc.regs[11][1] ;
 wire \top_ihp.oisc.regs[11][20] ;
 wire \top_ihp.oisc.regs[11][21] ;
 wire \top_ihp.oisc.regs[11][22] ;
 wire \top_ihp.oisc.regs[11][23] ;
 wire \top_ihp.oisc.regs[11][24] ;
 wire \top_ihp.oisc.regs[11][25] ;
 wire \top_ihp.oisc.regs[11][26] ;
 wire \top_ihp.oisc.regs[11][27] ;
 wire \top_ihp.oisc.regs[11][28] ;
 wire \top_ihp.oisc.regs[11][29] ;
 wire \top_ihp.oisc.regs[11][2] ;
 wire \top_ihp.oisc.regs[11][30] ;
 wire \top_ihp.oisc.regs[11][31] ;
 wire \top_ihp.oisc.regs[11][3] ;
 wire \top_ihp.oisc.regs[11][4] ;
 wire \top_ihp.oisc.regs[11][5] ;
 wire \top_ihp.oisc.regs[11][6] ;
 wire \top_ihp.oisc.regs[11][7] ;
 wire \top_ihp.oisc.regs[11][8] ;
 wire \top_ihp.oisc.regs[11][9] ;
 wire \top_ihp.oisc.regs[12][0] ;
 wire \top_ihp.oisc.regs[12][10] ;
 wire \top_ihp.oisc.regs[12][11] ;
 wire \top_ihp.oisc.regs[12][12] ;
 wire \top_ihp.oisc.regs[12][13] ;
 wire \top_ihp.oisc.regs[12][14] ;
 wire \top_ihp.oisc.regs[12][15] ;
 wire \top_ihp.oisc.regs[12][16] ;
 wire \top_ihp.oisc.regs[12][17] ;
 wire \top_ihp.oisc.regs[12][18] ;
 wire \top_ihp.oisc.regs[12][19] ;
 wire \top_ihp.oisc.regs[12][1] ;
 wire \top_ihp.oisc.regs[12][20] ;
 wire \top_ihp.oisc.regs[12][21] ;
 wire \top_ihp.oisc.regs[12][22] ;
 wire \top_ihp.oisc.regs[12][23] ;
 wire \top_ihp.oisc.regs[12][24] ;
 wire \top_ihp.oisc.regs[12][25] ;
 wire \top_ihp.oisc.regs[12][26] ;
 wire \top_ihp.oisc.regs[12][27] ;
 wire \top_ihp.oisc.regs[12][28] ;
 wire \top_ihp.oisc.regs[12][29] ;
 wire \top_ihp.oisc.regs[12][2] ;
 wire \top_ihp.oisc.regs[12][30] ;
 wire \top_ihp.oisc.regs[12][31] ;
 wire \top_ihp.oisc.regs[12][3] ;
 wire \top_ihp.oisc.regs[12][4] ;
 wire \top_ihp.oisc.regs[12][5] ;
 wire \top_ihp.oisc.regs[12][6] ;
 wire \top_ihp.oisc.regs[12][7] ;
 wire \top_ihp.oisc.regs[12][8] ;
 wire \top_ihp.oisc.regs[12][9] ;
 wire \top_ihp.oisc.regs[13][0] ;
 wire \top_ihp.oisc.regs[13][10] ;
 wire \top_ihp.oisc.regs[13][11] ;
 wire \top_ihp.oisc.regs[13][12] ;
 wire \top_ihp.oisc.regs[13][13] ;
 wire \top_ihp.oisc.regs[13][14] ;
 wire \top_ihp.oisc.regs[13][15] ;
 wire \top_ihp.oisc.regs[13][16] ;
 wire \top_ihp.oisc.regs[13][17] ;
 wire \top_ihp.oisc.regs[13][18] ;
 wire \top_ihp.oisc.regs[13][19] ;
 wire \top_ihp.oisc.regs[13][1] ;
 wire \top_ihp.oisc.regs[13][20] ;
 wire \top_ihp.oisc.regs[13][21] ;
 wire \top_ihp.oisc.regs[13][22] ;
 wire \top_ihp.oisc.regs[13][23] ;
 wire \top_ihp.oisc.regs[13][24] ;
 wire \top_ihp.oisc.regs[13][25] ;
 wire \top_ihp.oisc.regs[13][26] ;
 wire \top_ihp.oisc.regs[13][27] ;
 wire \top_ihp.oisc.regs[13][28] ;
 wire \top_ihp.oisc.regs[13][29] ;
 wire \top_ihp.oisc.regs[13][2] ;
 wire \top_ihp.oisc.regs[13][30] ;
 wire \top_ihp.oisc.regs[13][31] ;
 wire \top_ihp.oisc.regs[13][3] ;
 wire \top_ihp.oisc.regs[13][4] ;
 wire \top_ihp.oisc.regs[13][5] ;
 wire \top_ihp.oisc.regs[13][6] ;
 wire \top_ihp.oisc.regs[13][7] ;
 wire \top_ihp.oisc.regs[13][8] ;
 wire \top_ihp.oisc.regs[13][9] ;
 wire \top_ihp.oisc.regs[14][0] ;
 wire \top_ihp.oisc.regs[14][10] ;
 wire \top_ihp.oisc.regs[14][11] ;
 wire \top_ihp.oisc.regs[14][12] ;
 wire \top_ihp.oisc.regs[14][13] ;
 wire \top_ihp.oisc.regs[14][14] ;
 wire \top_ihp.oisc.regs[14][15] ;
 wire \top_ihp.oisc.regs[14][16] ;
 wire \top_ihp.oisc.regs[14][17] ;
 wire \top_ihp.oisc.regs[14][18] ;
 wire \top_ihp.oisc.regs[14][19] ;
 wire \top_ihp.oisc.regs[14][1] ;
 wire \top_ihp.oisc.regs[14][20] ;
 wire \top_ihp.oisc.regs[14][21] ;
 wire \top_ihp.oisc.regs[14][22] ;
 wire \top_ihp.oisc.regs[14][23] ;
 wire \top_ihp.oisc.regs[14][24] ;
 wire \top_ihp.oisc.regs[14][25] ;
 wire \top_ihp.oisc.regs[14][26] ;
 wire \top_ihp.oisc.regs[14][27] ;
 wire \top_ihp.oisc.regs[14][28] ;
 wire \top_ihp.oisc.regs[14][29] ;
 wire \top_ihp.oisc.regs[14][2] ;
 wire \top_ihp.oisc.regs[14][30] ;
 wire \top_ihp.oisc.regs[14][31] ;
 wire \top_ihp.oisc.regs[14][3] ;
 wire \top_ihp.oisc.regs[14][4] ;
 wire \top_ihp.oisc.regs[14][5] ;
 wire \top_ihp.oisc.regs[14][6] ;
 wire \top_ihp.oisc.regs[14][7] ;
 wire \top_ihp.oisc.regs[14][8] ;
 wire \top_ihp.oisc.regs[14][9] ;
 wire \top_ihp.oisc.regs[15][0] ;
 wire \top_ihp.oisc.regs[15][10] ;
 wire \top_ihp.oisc.regs[15][11] ;
 wire \top_ihp.oisc.regs[15][12] ;
 wire \top_ihp.oisc.regs[15][13] ;
 wire \top_ihp.oisc.regs[15][14] ;
 wire \top_ihp.oisc.regs[15][15] ;
 wire \top_ihp.oisc.regs[15][16] ;
 wire \top_ihp.oisc.regs[15][17] ;
 wire \top_ihp.oisc.regs[15][18] ;
 wire \top_ihp.oisc.regs[15][19] ;
 wire \top_ihp.oisc.regs[15][1] ;
 wire \top_ihp.oisc.regs[15][20] ;
 wire \top_ihp.oisc.regs[15][21] ;
 wire \top_ihp.oisc.regs[15][22] ;
 wire \top_ihp.oisc.regs[15][23] ;
 wire \top_ihp.oisc.regs[15][24] ;
 wire \top_ihp.oisc.regs[15][25] ;
 wire \top_ihp.oisc.regs[15][26] ;
 wire \top_ihp.oisc.regs[15][27] ;
 wire \top_ihp.oisc.regs[15][28] ;
 wire \top_ihp.oisc.regs[15][29] ;
 wire \top_ihp.oisc.regs[15][2] ;
 wire \top_ihp.oisc.regs[15][30] ;
 wire \top_ihp.oisc.regs[15][31] ;
 wire \top_ihp.oisc.regs[15][3] ;
 wire \top_ihp.oisc.regs[15][4] ;
 wire \top_ihp.oisc.regs[15][5] ;
 wire \top_ihp.oisc.regs[15][6] ;
 wire \top_ihp.oisc.regs[15][7] ;
 wire \top_ihp.oisc.regs[15][8] ;
 wire \top_ihp.oisc.regs[15][9] ;
 wire \top_ihp.oisc.regs[16][0] ;
 wire \top_ihp.oisc.regs[16][10] ;
 wire \top_ihp.oisc.regs[16][11] ;
 wire \top_ihp.oisc.regs[16][12] ;
 wire \top_ihp.oisc.regs[16][13] ;
 wire \top_ihp.oisc.regs[16][14] ;
 wire \top_ihp.oisc.regs[16][15] ;
 wire \top_ihp.oisc.regs[16][16] ;
 wire \top_ihp.oisc.regs[16][17] ;
 wire \top_ihp.oisc.regs[16][18] ;
 wire \top_ihp.oisc.regs[16][19] ;
 wire \top_ihp.oisc.regs[16][1] ;
 wire \top_ihp.oisc.regs[16][20] ;
 wire \top_ihp.oisc.regs[16][21] ;
 wire \top_ihp.oisc.regs[16][22] ;
 wire \top_ihp.oisc.regs[16][23] ;
 wire \top_ihp.oisc.regs[16][24] ;
 wire \top_ihp.oisc.regs[16][25] ;
 wire \top_ihp.oisc.regs[16][26] ;
 wire \top_ihp.oisc.regs[16][27] ;
 wire \top_ihp.oisc.regs[16][28] ;
 wire \top_ihp.oisc.regs[16][29] ;
 wire \top_ihp.oisc.regs[16][2] ;
 wire \top_ihp.oisc.regs[16][30] ;
 wire \top_ihp.oisc.regs[16][31] ;
 wire \top_ihp.oisc.regs[16][3] ;
 wire \top_ihp.oisc.regs[16][4] ;
 wire \top_ihp.oisc.regs[16][5] ;
 wire \top_ihp.oisc.regs[16][6] ;
 wire \top_ihp.oisc.regs[16][7] ;
 wire \top_ihp.oisc.regs[16][8] ;
 wire \top_ihp.oisc.regs[16][9] ;
 wire \top_ihp.oisc.regs[17][0] ;
 wire \top_ihp.oisc.regs[17][10] ;
 wire \top_ihp.oisc.regs[17][11] ;
 wire \top_ihp.oisc.regs[17][12] ;
 wire \top_ihp.oisc.regs[17][13] ;
 wire \top_ihp.oisc.regs[17][14] ;
 wire \top_ihp.oisc.regs[17][15] ;
 wire \top_ihp.oisc.regs[17][16] ;
 wire \top_ihp.oisc.regs[17][17] ;
 wire \top_ihp.oisc.regs[17][18] ;
 wire \top_ihp.oisc.regs[17][19] ;
 wire \top_ihp.oisc.regs[17][1] ;
 wire \top_ihp.oisc.regs[17][20] ;
 wire \top_ihp.oisc.regs[17][21] ;
 wire \top_ihp.oisc.regs[17][22] ;
 wire \top_ihp.oisc.regs[17][23] ;
 wire \top_ihp.oisc.regs[17][24] ;
 wire \top_ihp.oisc.regs[17][25] ;
 wire \top_ihp.oisc.regs[17][26] ;
 wire \top_ihp.oisc.regs[17][27] ;
 wire \top_ihp.oisc.regs[17][28] ;
 wire \top_ihp.oisc.regs[17][29] ;
 wire \top_ihp.oisc.regs[17][2] ;
 wire \top_ihp.oisc.regs[17][30] ;
 wire \top_ihp.oisc.regs[17][31] ;
 wire \top_ihp.oisc.regs[17][3] ;
 wire \top_ihp.oisc.regs[17][4] ;
 wire \top_ihp.oisc.regs[17][5] ;
 wire \top_ihp.oisc.regs[17][6] ;
 wire \top_ihp.oisc.regs[17][7] ;
 wire \top_ihp.oisc.regs[17][8] ;
 wire \top_ihp.oisc.regs[17][9] ;
 wire \top_ihp.oisc.regs[18][0] ;
 wire \top_ihp.oisc.regs[18][10] ;
 wire \top_ihp.oisc.regs[18][11] ;
 wire \top_ihp.oisc.regs[18][12] ;
 wire \top_ihp.oisc.regs[18][13] ;
 wire \top_ihp.oisc.regs[18][14] ;
 wire \top_ihp.oisc.regs[18][15] ;
 wire \top_ihp.oisc.regs[18][16] ;
 wire \top_ihp.oisc.regs[18][17] ;
 wire \top_ihp.oisc.regs[18][18] ;
 wire \top_ihp.oisc.regs[18][19] ;
 wire \top_ihp.oisc.regs[18][1] ;
 wire \top_ihp.oisc.regs[18][20] ;
 wire \top_ihp.oisc.regs[18][21] ;
 wire \top_ihp.oisc.regs[18][22] ;
 wire \top_ihp.oisc.regs[18][23] ;
 wire \top_ihp.oisc.regs[18][24] ;
 wire \top_ihp.oisc.regs[18][25] ;
 wire \top_ihp.oisc.regs[18][26] ;
 wire \top_ihp.oisc.regs[18][27] ;
 wire \top_ihp.oisc.regs[18][28] ;
 wire \top_ihp.oisc.regs[18][29] ;
 wire \top_ihp.oisc.regs[18][2] ;
 wire \top_ihp.oisc.regs[18][30] ;
 wire \top_ihp.oisc.regs[18][31] ;
 wire \top_ihp.oisc.regs[18][3] ;
 wire \top_ihp.oisc.regs[18][4] ;
 wire \top_ihp.oisc.regs[18][5] ;
 wire \top_ihp.oisc.regs[18][6] ;
 wire \top_ihp.oisc.regs[18][7] ;
 wire \top_ihp.oisc.regs[18][8] ;
 wire \top_ihp.oisc.regs[18][9] ;
 wire \top_ihp.oisc.regs[19][0] ;
 wire \top_ihp.oisc.regs[19][10] ;
 wire \top_ihp.oisc.regs[19][11] ;
 wire \top_ihp.oisc.regs[19][12] ;
 wire \top_ihp.oisc.regs[19][13] ;
 wire \top_ihp.oisc.regs[19][14] ;
 wire \top_ihp.oisc.regs[19][15] ;
 wire \top_ihp.oisc.regs[19][16] ;
 wire \top_ihp.oisc.regs[19][17] ;
 wire \top_ihp.oisc.regs[19][18] ;
 wire \top_ihp.oisc.regs[19][19] ;
 wire \top_ihp.oisc.regs[19][1] ;
 wire \top_ihp.oisc.regs[19][20] ;
 wire \top_ihp.oisc.regs[19][21] ;
 wire \top_ihp.oisc.regs[19][22] ;
 wire \top_ihp.oisc.regs[19][23] ;
 wire \top_ihp.oisc.regs[19][24] ;
 wire \top_ihp.oisc.regs[19][25] ;
 wire \top_ihp.oisc.regs[19][26] ;
 wire \top_ihp.oisc.regs[19][27] ;
 wire \top_ihp.oisc.regs[19][28] ;
 wire \top_ihp.oisc.regs[19][29] ;
 wire \top_ihp.oisc.regs[19][2] ;
 wire \top_ihp.oisc.regs[19][30] ;
 wire \top_ihp.oisc.regs[19][31] ;
 wire \top_ihp.oisc.regs[19][3] ;
 wire \top_ihp.oisc.regs[19][4] ;
 wire \top_ihp.oisc.regs[19][5] ;
 wire \top_ihp.oisc.regs[19][6] ;
 wire \top_ihp.oisc.regs[19][7] ;
 wire \top_ihp.oisc.regs[19][8] ;
 wire \top_ihp.oisc.regs[19][9] ;
 wire \top_ihp.oisc.regs[1][0] ;
 wire \top_ihp.oisc.regs[1][10] ;
 wire \top_ihp.oisc.regs[1][11] ;
 wire \top_ihp.oisc.regs[1][12] ;
 wire \top_ihp.oisc.regs[1][13] ;
 wire \top_ihp.oisc.regs[1][14] ;
 wire \top_ihp.oisc.regs[1][15] ;
 wire \top_ihp.oisc.regs[1][16] ;
 wire \top_ihp.oisc.regs[1][17] ;
 wire \top_ihp.oisc.regs[1][18] ;
 wire \top_ihp.oisc.regs[1][19] ;
 wire \top_ihp.oisc.regs[1][1] ;
 wire \top_ihp.oisc.regs[1][20] ;
 wire \top_ihp.oisc.regs[1][21] ;
 wire \top_ihp.oisc.regs[1][22] ;
 wire \top_ihp.oisc.regs[1][23] ;
 wire \top_ihp.oisc.regs[1][24] ;
 wire \top_ihp.oisc.regs[1][25] ;
 wire \top_ihp.oisc.regs[1][26] ;
 wire \top_ihp.oisc.regs[1][27] ;
 wire \top_ihp.oisc.regs[1][28] ;
 wire \top_ihp.oisc.regs[1][29] ;
 wire \top_ihp.oisc.regs[1][2] ;
 wire \top_ihp.oisc.regs[1][30] ;
 wire \top_ihp.oisc.regs[1][31] ;
 wire \top_ihp.oisc.regs[1][3] ;
 wire \top_ihp.oisc.regs[1][4] ;
 wire \top_ihp.oisc.regs[1][5] ;
 wire \top_ihp.oisc.regs[1][6] ;
 wire \top_ihp.oisc.regs[1][7] ;
 wire \top_ihp.oisc.regs[1][8] ;
 wire \top_ihp.oisc.regs[1][9] ;
 wire \top_ihp.oisc.regs[20][0] ;
 wire \top_ihp.oisc.regs[20][10] ;
 wire \top_ihp.oisc.regs[20][11] ;
 wire \top_ihp.oisc.regs[20][12] ;
 wire \top_ihp.oisc.regs[20][13] ;
 wire \top_ihp.oisc.regs[20][14] ;
 wire \top_ihp.oisc.regs[20][15] ;
 wire \top_ihp.oisc.regs[20][16] ;
 wire \top_ihp.oisc.regs[20][17] ;
 wire \top_ihp.oisc.regs[20][18] ;
 wire \top_ihp.oisc.regs[20][19] ;
 wire \top_ihp.oisc.regs[20][1] ;
 wire \top_ihp.oisc.regs[20][20] ;
 wire \top_ihp.oisc.regs[20][21] ;
 wire \top_ihp.oisc.regs[20][22] ;
 wire \top_ihp.oisc.regs[20][23] ;
 wire \top_ihp.oisc.regs[20][24] ;
 wire \top_ihp.oisc.regs[20][25] ;
 wire \top_ihp.oisc.regs[20][26] ;
 wire \top_ihp.oisc.regs[20][27] ;
 wire \top_ihp.oisc.regs[20][28] ;
 wire \top_ihp.oisc.regs[20][29] ;
 wire \top_ihp.oisc.regs[20][2] ;
 wire \top_ihp.oisc.regs[20][30] ;
 wire \top_ihp.oisc.regs[20][31] ;
 wire \top_ihp.oisc.regs[20][3] ;
 wire \top_ihp.oisc.regs[20][4] ;
 wire \top_ihp.oisc.regs[20][5] ;
 wire \top_ihp.oisc.regs[20][6] ;
 wire \top_ihp.oisc.regs[20][7] ;
 wire \top_ihp.oisc.regs[20][8] ;
 wire \top_ihp.oisc.regs[20][9] ;
 wire \top_ihp.oisc.regs[21][0] ;
 wire \top_ihp.oisc.regs[21][10] ;
 wire \top_ihp.oisc.regs[21][11] ;
 wire \top_ihp.oisc.regs[21][12] ;
 wire \top_ihp.oisc.regs[21][13] ;
 wire \top_ihp.oisc.regs[21][14] ;
 wire \top_ihp.oisc.regs[21][15] ;
 wire \top_ihp.oisc.regs[21][16] ;
 wire \top_ihp.oisc.regs[21][17] ;
 wire \top_ihp.oisc.regs[21][18] ;
 wire \top_ihp.oisc.regs[21][19] ;
 wire \top_ihp.oisc.regs[21][1] ;
 wire \top_ihp.oisc.regs[21][20] ;
 wire \top_ihp.oisc.regs[21][21] ;
 wire \top_ihp.oisc.regs[21][22] ;
 wire \top_ihp.oisc.regs[21][23] ;
 wire \top_ihp.oisc.regs[21][24] ;
 wire \top_ihp.oisc.regs[21][25] ;
 wire \top_ihp.oisc.regs[21][26] ;
 wire \top_ihp.oisc.regs[21][27] ;
 wire \top_ihp.oisc.regs[21][28] ;
 wire \top_ihp.oisc.regs[21][29] ;
 wire \top_ihp.oisc.regs[21][2] ;
 wire \top_ihp.oisc.regs[21][30] ;
 wire \top_ihp.oisc.regs[21][31] ;
 wire \top_ihp.oisc.regs[21][3] ;
 wire \top_ihp.oisc.regs[21][4] ;
 wire \top_ihp.oisc.regs[21][5] ;
 wire \top_ihp.oisc.regs[21][6] ;
 wire \top_ihp.oisc.regs[21][7] ;
 wire \top_ihp.oisc.regs[21][8] ;
 wire \top_ihp.oisc.regs[21][9] ;
 wire \top_ihp.oisc.regs[22][0] ;
 wire \top_ihp.oisc.regs[22][10] ;
 wire \top_ihp.oisc.regs[22][11] ;
 wire \top_ihp.oisc.regs[22][12] ;
 wire \top_ihp.oisc.regs[22][13] ;
 wire \top_ihp.oisc.regs[22][14] ;
 wire \top_ihp.oisc.regs[22][15] ;
 wire \top_ihp.oisc.regs[22][16] ;
 wire \top_ihp.oisc.regs[22][17] ;
 wire \top_ihp.oisc.regs[22][18] ;
 wire \top_ihp.oisc.regs[22][19] ;
 wire \top_ihp.oisc.regs[22][1] ;
 wire \top_ihp.oisc.regs[22][20] ;
 wire \top_ihp.oisc.regs[22][21] ;
 wire \top_ihp.oisc.regs[22][22] ;
 wire \top_ihp.oisc.regs[22][23] ;
 wire \top_ihp.oisc.regs[22][24] ;
 wire \top_ihp.oisc.regs[22][25] ;
 wire \top_ihp.oisc.regs[22][26] ;
 wire \top_ihp.oisc.regs[22][27] ;
 wire \top_ihp.oisc.regs[22][28] ;
 wire \top_ihp.oisc.regs[22][29] ;
 wire \top_ihp.oisc.regs[22][2] ;
 wire \top_ihp.oisc.regs[22][30] ;
 wire \top_ihp.oisc.regs[22][31] ;
 wire \top_ihp.oisc.regs[22][3] ;
 wire \top_ihp.oisc.regs[22][4] ;
 wire \top_ihp.oisc.regs[22][5] ;
 wire \top_ihp.oisc.regs[22][6] ;
 wire \top_ihp.oisc.regs[22][7] ;
 wire \top_ihp.oisc.regs[22][8] ;
 wire \top_ihp.oisc.regs[22][9] ;
 wire \top_ihp.oisc.regs[23][0] ;
 wire \top_ihp.oisc.regs[23][10] ;
 wire \top_ihp.oisc.regs[23][11] ;
 wire \top_ihp.oisc.regs[23][12] ;
 wire \top_ihp.oisc.regs[23][13] ;
 wire \top_ihp.oisc.regs[23][14] ;
 wire \top_ihp.oisc.regs[23][15] ;
 wire \top_ihp.oisc.regs[23][16] ;
 wire \top_ihp.oisc.regs[23][17] ;
 wire \top_ihp.oisc.regs[23][18] ;
 wire \top_ihp.oisc.regs[23][19] ;
 wire \top_ihp.oisc.regs[23][1] ;
 wire \top_ihp.oisc.regs[23][20] ;
 wire \top_ihp.oisc.regs[23][21] ;
 wire \top_ihp.oisc.regs[23][22] ;
 wire \top_ihp.oisc.regs[23][23] ;
 wire \top_ihp.oisc.regs[23][24] ;
 wire \top_ihp.oisc.regs[23][25] ;
 wire \top_ihp.oisc.regs[23][26] ;
 wire \top_ihp.oisc.regs[23][27] ;
 wire \top_ihp.oisc.regs[23][28] ;
 wire \top_ihp.oisc.regs[23][29] ;
 wire \top_ihp.oisc.regs[23][2] ;
 wire \top_ihp.oisc.regs[23][30] ;
 wire \top_ihp.oisc.regs[23][31] ;
 wire \top_ihp.oisc.regs[23][3] ;
 wire \top_ihp.oisc.regs[23][4] ;
 wire \top_ihp.oisc.regs[23][5] ;
 wire \top_ihp.oisc.regs[23][6] ;
 wire \top_ihp.oisc.regs[23][7] ;
 wire \top_ihp.oisc.regs[23][8] ;
 wire \top_ihp.oisc.regs[23][9] ;
 wire \top_ihp.oisc.regs[24][0] ;
 wire \top_ihp.oisc.regs[24][10] ;
 wire \top_ihp.oisc.regs[24][11] ;
 wire \top_ihp.oisc.regs[24][12] ;
 wire \top_ihp.oisc.regs[24][13] ;
 wire \top_ihp.oisc.regs[24][14] ;
 wire \top_ihp.oisc.regs[24][15] ;
 wire \top_ihp.oisc.regs[24][16] ;
 wire \top_ihp.oisc.regs[24][17] ;
 wire \top_ihp.oisc.regs[24][18] ;
 wire \top_ihp.oisc.regs[24][19] ;
 wire \top_ihp.oisc.regs[24][1] ;
 wire \top_ihp.oisc.regs[24][20] ;
 wire \top_ihp.oisc.regs[24][21] ;
 wire \top_ihp.oisc.regs[24][22] ;
 wire \top_ihp.oisc.regs[24][23] ;
 wire \top_ihp.oisc.regs[24][24] ;
 wire \top_ihp.oisc.regs[24][25] ;
 wire \top_ihp.oisc.regs[24][26] ;
 wire \top_ihp.oisc.regs[24][27] ;
 wire \top_ihp.oisc.regs[24][28] ;
 wire \top_ihp.oisc.regs[24][29] ;
 wire \top_ihp.oisc.regs[24][2] ;
 wire \top_ihp.oisc.regs[24][30] ;
 wire \top_ihp.oisc.regs[24][31] ;
 wire \top_ihp.oisc.regs[24][3] ;
 wire \top_ihp.oisc.regs[24][4] ;
 wire \top_ihp.oisc.regs[24][5] ;
 wire \top_ihp.oisc.regs[24][6] ;
 wire \top_ihp.oisc.regs[24][7] ;
 wire \top_ihp.oisc.regs[24][8] ;
 wire \top_ihp.oisc.regs[24][9] ;
 wire \top_ihp.oisc.regs[25][0] ;
 wire \top_ihp.oisc.regs[25][10] ;
 wire \top_ihp.oisc.regs[25][11] ;
 wire \top_ihp.oisc.regs[25][12] ;
 wire \top_ihp.oisc.regs[25][13] ;
 wire \top_ihp.oisc.regs[25][14] ;
 wire \top_ihp.oisc.regs[25][15] ;
 wire \top_ihp.oisc.regs[25][16] ;
 wire \top_ihp.oisc.regs[25][17] ;
 wire \top_ihp.oisc.regs[25][18] ;
 wire \top_ihp.oisc.regs[25][19] ;
 wire \top_ihp.oisc.regs[25][1] ;
 wire \top_ihp.oisc.regs[25][20] ;
 wire \top_ihp.oisc.regs[25][21] ;
 wire \top_ihp.oisc.regs[25][22] ;
 wire \top_ihp.oisc.regs[25][23] ;
 wire \top_ihp.oisc.regs[25][24] ;
 wire \top_ihp.oisc.regs[25][25] ;
 wire \top_ihp.oisc.regs[25][26] ;
 wire \top_ihp.oisc.regs[25][27] ;
 wire \top_ihp.oisc.regs[25][28] ;
 wire \top_ihp.oisc.regs[25][29] ;
 wire \top_ihp.oisc.regs[25][2] ;
 wire \top_ihp.oisc.regs[25][30] ;
 wire \top_ihp.oisc.regs[25][31] ;
 wire \top_ihp.oisc.regs[25][3] ;
 wire \top_ihp.oisc.regs[25][4] ;
 wire \top_ihp.oisc.regs[25][5] ;
 wire \top_ihp.oisc.regs[25][6] ;
 wire \top_ihp.oisc.regs[25][7] ;
 wire \top_ihp.oisc.regs[25][8] ;
 wire \top_ihp.oisc.regs[25][9] ;
 wire \top_ihp.oisc.regs[26][0] ;
 wire \top_ihp.oisc.regs[26][10] ;
 wire \top_ihp.oisc.regs[26][11] ;
 wire \top_ihp.oisc.regs[26][12] ;
 wire \top_ihp.oisc.regs[26][13] ;
 wire \top_ihp.oisc.regs[26][14] ;
 wire \top_ihp.oisc.regs[26][15] ;
 wire \top_ihp.oisc.regs[26][16] ;
 wire \top_ihp.oisc.regs[26][17] ;
 wire \top_ihp.oisc.regs[26][18] ;
 wire \top_ihp.oisc.regs[26][19] ;
 wire \top_ihp.oisc.regs[26][1] ;
 wire \top_ihp.oisc.regs[26][20] ;
 wire \top_ihp.oisc.regs[26][21] ;
 wire \top_ihp.oisc.regs[26][22] ;
 wire \top_ihp.oisc.regs[26][23] ;
 wire \top_ihp.oisc.regs[26][24] ;
 wire \top_ihp.oisc.regs[26][25] ;
 wire \top_ihp.oisc.regs[26][26] ;
 wire \top_ihp.oisc.regs[26][27] ;
 wire \top_ihp.oisc.regs[26][28] ;
 wire \top_ihp.oisc.regs[26][29] ;
 wire \top_ihp.oisc.regs[26][2] ;
 wire \top_ihp.oisc.regs[26][30] ;
 wire \top_ihp.oisc.regs[26][31] ;
 wire \top_ihp.oisc.regs[26][3] ;
 wire \top_ihp.oisc.regs[26][4] ;
 wire \top_ihp.oisc.regs[26][5] ;
 wire \top_ihp.oisc.regs[26][6] ;
 wire \top_ihp.oisc.regs[26][7] ;
 wire \top_ihp.oisc.regs[26][8] ;
 wire \top_ihp.oisc.regs[26][9] ;
 wire \top_ihp.oisc.regs[27][0] ;
 wire \top_ihp.oisc.regs[27][10] ;
 wire \top_ihp.oisc.regs[27][11] ;
 wire \top_ihp.oisc.regs[27][12] ;
 wire \top_ihp.oisc.regs[27][13] ;
 wire \top_ihp.oisc.regs[27][14] ;
 wire \top_ihp.oisc.regs[27][15] ;
 wire \top_ihp.oisc.regs[27][16] ;
 wire \top_ihp.oisc.regs[27][17] ;
 wire \top_ihp.oisc.regs[27][18] ;
 wire \top_ihp.oisc.regs[27][19] ;
 wire \top_ihp.oisc.regs[27][1] ;
 wire \top_ihp.oisc.regs[27][20] ;
 wire \top_ihp.oisc.regs[27][21] ;
 wire \top_ihp.oisc.regs[27][22] ;
 wire \top_ihp.oisc.regs[27][23] ;
 wire \top_ihp.oisc.regs[27][24] ;
 wire \top_ihp.oisc.regs[27][25] ;
 wire \top_ihp.oisc.regs[27][26] ;
 wire \top_ihp.oisc.regs[27][27] ;
 wire \top_ihp.oisc.regs[27][28] ;
 wire \top_ihp.oisc.regs[27][29] ;
 wire \top_ihp.oisc.regs[27][2] ;
 wire \top_ihp.oisc.regs[27][30] ;
 wire \top_ihp.oisc.regs[27][31] ;
 wire \top_ihp.oisc.regs[27][3] ;
 wire \top_ihp.oisc.regs[27][4] ;
 wire \top_ihp.oisc.regs[27][5] ;
 wire \top_ihp.oisc.regs[27][6] ;
 wire \top_ihp.oisc.regs[27][7] ;
 wire \top_ihp.oisc.regs[27][8] ;
 wire \top_ihp.oisc.regs[27][9] ;
 wire \top_ihp.oisc.regs[28][0] ;
 wire \top_ihp.oisc.regs[28][10] ;
 wire \top_ihp.oisc.regs[28][11] ;
 wire \top_ihp.oisc.regs[28][12] ;
 wire \top_ihp.oisc.regs[28][13] ;
 wire \top_ihp.oisc.regs[28][14] ;
 wire \top_ihp.oisc.regs[28][15] ;
 wire \top_ihp.oisc.regs[28][16] ;
 wire \top_ihp.oisc.regs[28][17] ;
 wire \top_ihp.oisc.regs[28][18] ;
 wire \top_ihp.oisc.regs[28][19] ;
 wire \top_ihp.oisc.regs[28][1] ;
 wire \top_ihp.oisc.regs[28][20] ;
 wire \top_ihp.oisc.regs[28][21] ;
 wire \top_ihp.oisc.regs[28][22] ;
 wire \top_ihp.oisc.regs[28][23] ;
 wire \top_ihp.oisc.regs[28][24] ;
 wire \top_ihp.oisc.regs[28][25] ;
 wire \top_ihp.oisc.regs[28][26] ;
 wire \top_ihp.oisc.regs[28][27] ;
 wire \top_ihp.oisc.regs[28][28] ;
 wire \top_ihp.oisc.regs[28][29] ;
 wire \top_ihp.oisc.regs[28][2] ;
 wire \top_ihp.oisc.regs[28][30] ;
 wire \top_ihp.oisc.regs[28][31] ;
 wire \top_ihp.oisc.regs[28][3] ;
 wire \top_ihp.oisc.regs[28][4] ;
 wire \top_ihp.oisc.regs[28][5] ;
 wire \top_ihp.oisc.regs[28][6] ;
 wire \top_ihp.oisc.regs[28][7] ;
 wire \top_ihp.oisc.regs[28][8] ;
 wire \top_ihp.oisc.regs[28][9] ;
 wire \top_ihp.oisc.regs[29][0] ;
 wire \top_ihp.oisc.regs[29][10] ;
 wire \top_ihp.oisc.regs[29][11] ;
 wire \top_ihp.oisc.regs[29][12] ;
 wire \top_ihp.oisc.regs[29][13] ;
 wire \top_ihp.oisc.regs[29][14] ;
 wire \top_ihp.oisc.regs[29][15] ;
 wire \top_ihp.oisc.regs[29][16] ;
 wire \top_ihp.oisc.regs[29][17] ;
 wire \top_ihp.oisc.regs[29][18] ;
 wire \top_ihp.oisc.regs[29][19] ;
 wire \top_ihp.oisc.regs[29][1] ;
 wire \top_ihp.oisc.regs[29][20] ;
 wire \top_ihp.oisc.regs[29][21] ;
 wire \top_ihp.oisc.regs[29][22] ;
 wire \top_ihp.oisc.regs[29][23] ;
 wire \top_ihp.oisc.regs[29][24] ;
 wire \top_ihp.oisc.regs[29][25] ;
 wire \top_ihp.oisc.regs[29][26] ;
 wire \top_ihp.oisc.regs[29][27] ;
 wire \top_ihp.oisc.regs[29][28] ;
 wire \top_ihp.oisc.regs[29][29] ;
 wire \top_ihp.oisc.regs[29][2] ;
 wire \top_ihp.oisc.regs[29][30] ;
 wire \top_ihp.oisc.regs[29][31] ;
 wire \top_ihp.oisc.regs[29][3] ;
 wire \top_ihp.oisc.regs[29][4] ;
 wire \top_ihp.oisc.regs[29][5] ;
 wire \top_ihp.oisc.regs[29][6] ;
 wire \top_ihp.oisc.regs[29][7] ;
 wire \top_ihp.oisc.regs[29][8] ;
 wire \top_ihp.oisc.regs[29][9] ;
 wire \top_ihp.oisc.regs[2][0] ;
 wire \top_ihp.oisc.regs[2][10] ;
 wire \top_ihp.oisc.regs[2][11] ;
 wire \top_ihp.oisc.regs[2][12] ;
 wire \top_ihp.oisc.regs[2][13] ;
 wire \top_ihp.oisc.regs[2][14] ;
 wire \top_ihp.oisc.regs[2][15] ;
 wire \top_ihp.oisc.regs[2][16] ;
 wire \top_ihp.oisc.regs[2][17] ;
 wire \top_ihp.oisc.regs[2][18] ;
 wire \top_ihp.oisc.regs[2][19] ;
 wire \top_ihp.oisc.regs[2][1] ;
 wire \top_ihp.oisc.regs[2][20] ;
 wire \top_ihp.oisc.regs[2][21] ;
 wire \top_ihp.oisc.regs[2][22] ;
 wire \top_ihp.oisc.regs[2][23] ;
 wire \top_ihp.oisc.regs[2][24] ;
 wire \top_ihp.oisc.regs[2][25] ;
 wire \top_ihp.oisc.regs[2][26] ;
 wire \top_ihp.oisc.regs[2][27] ;
 wire \top_ihp.oisc.regs[2][28] ;
 wire \top_ihp.oisc.regs[2][29] ;
 wire \top_ihp.oisc.regs[2][2] ;
 wire \top_ihp.oisc.regs[2][30] ;
 wire \top_ihp.oisc.regs[2][31] ;
 wire \top_ihp.oisc.regs[2][3] ;
 wire \top_ihp.oisc.regs[2][4] ;
 wire \top_ihp.oisc.regs[2][5] ;
 wire \top_ihp.oisc.regs[2][6] ;
 wire \top_ihp.oisc.regs[2][7] ;
 wire \top_ihp.oisc.regs[2][8] ;
 wire \top_ihp.oisc.regs[2][9] ;
 wire \top_ihp.oisc.regs[30][0] ;
 wire \top_ihp.oisc.regs[30][10] ;
 wire \top_ihp.oisc.regs[30][11] ;
 wire \top_ihp.oisc.regs[30][12] ;
 wire \top_ihp.oisc.regs[30][13] ;
 wire \top_ihp.oisc.regs[30][14] ;
 wire \top_ihp.oisc.regs[30][15] ;
 wire \top_ihp.oisc.regs[30][16] ;
 wire \top_ihp.oisc.regs[30][17] ;
 wire \top_ihp.oisc.regs[30][18] ;
 wire \top_ihp.oisc.regs[30][19] ;
 wire \top_ihp.oisc.regs[30][1] ;
 wire \top_ihp.oisc.regs[30][20] ;
 wire \top_ihp.oisc.regs[30][21] ;
 wire \top_ihp.oisc.regs[30][22] ;
 wire \top_ihp.oisc.regs[30][23] ;
 wire \top_ihp.oisc.regs[30][24] ;
 wire \top_ihp.oisc.regs[30][25] ;
 wire \top_ihp.oisc.regs[30][26] ;
 wire \top_ihp.oisc.regs[30][27] ;
 wire \top_ihp.oisc.regs[30][28] ;
 wire \top_ihp.oisc.regs[30][29] ;
 wire \top_ihp.oisc.regs[30][2] ;
 wire \top_ihp.oisc.regs[30][30] ;
 wire \top_ihp.oisc.regs[30][31] ;
 wire \top_ihp.oisc.regs[30][3] ;
 wire \top_ihp.oisc.regs[30][4] ;
 wire \top_ihp.oisc.regs[30][5] ;
 wire \top_ihp.oisc.regs[30][6] ;
 wire \top_ihp.oisc.regs[30][7] ;
 wire \top_ihp.oisc.regs[30][8] ;
 wire \top_ihp.oisc.regs[30][9] ;
 wire \top_ihp.oisc.regs[31][0] ;
 wire \top_ihp.oisc.regs[31][10] ;
 wire \top_ihp.oisc.regs[31][11] ;
 wire \top_ihp.oisc.regs[31][12] ;
 wire \top_ihp.oisc.regs[31][13] ;
 wire \top_ihp.oisc.regs[31][14] ;
 wire \top_ihp.oisc.regs[31][15] ;
 wire \top_ihp.oisc.regs[31][16] ;
 wire \top_ihp.oisc.regs[31][17] ;
 wire \top_ihp.oisc.regs[31][18] ;
 wire \top_ihp.oisc.regs[31][19] ;
 wire \top_ihp.oisc.regs[31][1] ;
 wire \top_ihp.oisc.regs[31][20] ;
 wire \top_ihp.oisc.regs[31][21] ;
 wire \top_ihp.oisc.regs[31][22] ;
 wire \top_ihp.oisc.regs[31][23] ;
 wire \top_ihp.oisc.regs[31][24] ;
 wire \top_ihp.oisc.regs[31][25] ;
 wire \top_ihp.oisc.regs[31][26] ;
 wire \top_ihp.oisc.regs[31][27] ;
 wire \top_ihp.oisc.regs[31][28] ;
 wire \top_ihp.oisc.regs[31][29] ;
 wire \top_ihp.oisc.regs[31][2] ;
 wire \top_ihp.oisc.regs[31][30] ;
 wire \top_ihp.oisc.regs[31][31] ;
 wire \top_ihp.oisc.regs[31][3] ;
 wire \top_ihp.oisc.regs[31][4] ;
 wire \top_ihp.oisc.regs[31][5] ;
 wire \top_ihp.oisc.regs[31][6] ;
 wire \top_ihp.oisc.regs[31][7] ;
 wire \top_ihp.oisc.regs[31][8] ;
 wire \top_ihp.oisc.regs[31][9] ;
 wire \top_ihp.oisc.regs[32][0] ;
 wire \top_ihp.oisc.regs[32][10] ;
 wire \top_ihp.oisc.regs[32][11] ;
 wire \top_ihp.oisc.regs[32][12] ;
 wire \top_ihp.oisc.regs[32][13] ;
 wire \top_ihp.oisc.regs[32][14] ;
 wire \top_ihp.oisc.regs[32][15] ;
 wire \top_ihp.oisc.regs[32][16] ;
 wire \top_ihp.oisc.regs[32][17] ;
 wire \top_ihp.oisc.regs[32][18] ;
 wire \top_ihp.oisc.regs[32][19] ;
 wire \top_ihp.oisc.regs[32][1] ;
 wire \top_ihp.oisc.regs[32][20] ;
 wire \top_ihp.oisc.regs[32][21] ;
 wire \top_ihp.oisc.regs[32][22] ;
 wire \top_ihp.oisc.regs[32][23] ;
 wire \top_ihp.oisc.regs[32][24] ;
 wire \top_ihp.oisc.regs[32][25] ;
 wire \top_ihp.oisc.regs[32][26] ;
 wire \top_ihp.oisc.regs[32][27] ;
 wire \top_ihp.oisc.regs[32][28] ;
 wire \top_ihp.oisc.regs[32][29] ;
 wire \top_ihp.oisc.regs[32][2] ;
 wire \top_ihp.oisc.regs[32][30] ;
 wire \top_ihp.oisc.regs[32][31] ;
 wire \top_ihp.oisc.regs[32][3] ;
 wire \top_ihp.oisc.regs[32][4] ;
 wire \top_ihp.oisc.regs[32][5] ;
 wire \top_ihp.oisc.regs[32][6] ;
 wire \top_ihp.oisc.regs[32][7] ;
 wire \top_ihp.oisc.regs[32][8] ;
 wire \top_ihp.oisc.regs[32][9] ;
 wire \top_ihp.oisc.regs[33][0] ;
 wire \top_ihp.oisc.regs[33][10] ;
 wire \top_ihp.oisc.regs[33][11] ;
 wire \top_ihp.oisc.regs[33][12] ;
 wire \top_ihp.oisc.regs[33][13] ;
 wire \top_ihp.oisc.regs[33][14] ;
 wire \top_ihp.oisc.regs[33][15] ;
 wire \top_ihp.oisc.regs[33][16] ;
 wire \top_ihp.oisc.regs[33][17] ;
 wire \top_ihp.oisc.regs[33][18] ;
 wire \top_ihp.oisc.regs[33][19] ;
 wire \top_ihp.oisc.regs[33][1] ;
 wire \top_ihp.oisc.regs[33][20] ;
 wire \top_ihp.oisc.regs[33][21] ;
 wire \top_ihp.oisc.regs[33][22] ;
 wire \top_ihp.oisc.regs[33][23] ;
 wire \top_ihp.oisc.regs[33][24] ;
 wire \top_ihp.oisc.regs[33][25] ;
 wire \top_ihp.oisc.regs[33][26] ;
 wire \top_ihp.oisc.regs[33][27] ;
 wire \top_ihp.oisc.regs[33][28] ;
 wire \top_ihp.oisc.regs[33][29] ;
 wire \top_ihp.oisc.regs[33][2] ;
 wire \top_ihp.oisc.regs[33][30] ;
 wire \top_ihp.oisc.regs[33][31] ;
 wire \top_ihp.oisc.regs[33][3] ;
 wire \top_ihp.oisc.regs[33][4] ;
 wire \top_ihp.oisc.regs[33][5] ;
 wire \top_ihp.oisc.regs[33][6] ;
 wire \top_ihp.oisc.regs[33][7] ;
 wire \top_ihp.oisc.regs[33][8] ;
 wire \top_ihp.oisc.regs[33][9] ;
 wire \top_ihp.oisc.regs[34][0] ;
 wire \top_ihp.oisc.regs[34][10] ;
 wire \top_ihp.oisc.regs[34][11] ;
 wire \top_ihp.oisc.regs[34][12] ;
 wire \top_ihp.oisc.regs[34][13] ;
 wire \top_ihp.oisc.regs[34][14] ;
 wire \top_ihp.oisc.regs[34][15] ;
 wire \top_ihp.oisc.regs[34][16] ;
 wire \top_ihp.oisc.regs[34][17] ;
 wire \top_ihp.oisc.regs[34][18] ;
 wire \top_ihp.oisc.regs[34][19] ;
 wire \top_ihp.oisc.regs[34][1] ;
 wire \top_ihp.oisc.regs[34][20] ;
 wire \top_ihp.oisc.regs[34][21] ;
 wire \top_ihp.oisc.regs[34][22] ;
 wire \top_ihp.oisc.regs[34][23] ;
 wire \top_ihp.oisc.regs[34][24] ;
 wire \top_ihp.oisc.regs[34][25] ;
 wire \top_ihp.oisc.regs[34][26] ;
 wire \top_ihp.oisc.regs[34][27] ;
 wire \top_ihp.oisc.regs[34][28] ;
 wire \top_ihp.oisc.regs[34][29] ;
 wire \top_ihp.oisc.regs[34][2] ;
 wire \top_ihp.oisc.regs[34][30] ;
 wire \top_ihp.oisc.regs[34][31] ;
 wire \top_ihp.oisc.regs[34][3] ;
 wire \top_ihp.oisc.regs[34][4] ;
 wire \top_ihp.oisc.regs[34][5] ;
 wire \top_ihp.oisc.regs[34][6] ;
 wire \top_ihp.oisc.regs[34][7] ;
 wire \top_ihp.oisc.regs[34][8] ;
 wire \top_ihp.oisc.regs[34][9] ;
 wire \top_ihp.oisc.regs[35][0] ;
 wire \top_ihp.oisc.regs[35][10] ;
 wire \top_ihp.oisc.regs[35][11] ;
 wire \top_ihp.oisc.regs[35][12] ;
 wire \top_ihp.oisc.regs[35][13] ;
 wire \top_ihp.oisc.regs[35][14] ;
 wire \top_ihp.oisc.regs[35][15] ;
 wire \top_ihp.oisc.regs[35][16] ;
 wire \top_ihp.oisc.regs[35][17] ;
 wire \top_ihp.oisc.regs[35][18] ;
 wire \top_ihp.oisc.regs[35][19] ;
 wire \top_ihp.oisc.regs[35][1] ;
 wire \top_ihp.oisc.regs[35][20] ;
 wire \top_ihp.oisc.regs[35][21] ;
 wire \top_ihp.oisc.regs[35][22] ;
 wire \top_ihp.oisc.regs[35][23] ;
 wire \top_ihp.oisc.regs[35][24] ;
 wire \top_ihp.oisc.regs[35][25] ;
 wire \top_ihp.oisc.regs[35][26] ;
 wire \top_ihp.oisc.regs[35][27] ;
 wire \top_ihp.oisc.regs[35][28] ;
 wire \top_ihp.oisc.regs[35][29] ;
 wire \top_ihp.oisc.regs[35][2] ;
 wire \top_ihp.oisc.regs[35][30] ;
 wire \top_ihp.oisc.regs[35][31] ;
 wire \top_ihp.oisc.regs[35][3] ;
 wire \top_ihp.oisc.regs[35][4] ;
 wire \top_ihp.oisc.regs[35][5] ;
 wire \top_ihp.oisc.regs[35][6] ;
 wire \top_ihp.oisc.regs[35][7] ;
 wire \top_ihp.oisc.regs[35][8] ;
 wire \top_ihp.oisc.regs[35][9] ;
 wire \top_ihp.oisc.regs[36][0] ;
 wire \top_ihp.oisc.regs[36][10] ;
 wire \top_ihp.oisc.regs[36][11] ;
 wire \top_ihp.oisc.regs[36][12] ;
 wire \top_ihp.oisc.regs[36][13] ;
 wire \top_ihp.oisc.regs[36][14] ;
 wire \top_ihp.oisc.regs[36][15] ;
 wire \top_ihp.oisc.regs[36][16] ;
 wire \top_ihp.oisc.regs[36][17] ;
 wire \top_ihp.oisc.regs[36][18] ;
 wire \top_ihp.oisc.regs[36][19] ;
 wire \top_ihp.oisc.regs[36][1] ;
 wire \top_ihp.oisc.regs[36][20] ;
 wire \top_ihp.oisc.regs[36][21] ;
 wire \top_ihp.oisc.regs[36][22] ;
 wire \top_ihp.oisc.regs[36][23] ;
 wire \top_ihp.oisc.regs[36][24] ;
 wire \top_ihp.oisc.regs[36][25] ;
 wire \top_ihp.oisc.regs[36][26] ;
 wire \top_ihp.oisc.regs[36][27] ;
 wire \top_ihp.oisc.regs[36][28] ;
 wire \top_ihp.oisc.regs[36][29] ;
 wire \top_ihp.oisc.regs[36][2] ;
 wire \top_ihp.oisc.regs[36][30] ;
 wire \top_ihp.oisc.regs[36][31] ;
 wire \top_ihp.oisc.regs[36][3] ;
 wire \top_ihp.oisc.regs[36][4] ;
 wire \top_ihp.oisc.regs[36][5] ;
 wire \top_ihp.oisc.regs[36][6] ;
 wire \top_ihp.oisc.regs[36][7] ;
 wire \top_ihp.oisc.regs[36][8] ;
 wire \top_ihp.oisc.regs[36][9] ;
 wire \top_ihp.oisc.regs[37][0] ;
 wire \top_ihp.oisc.regs[37][10] ;
 wire \top_ihp.oisc.regs[37][11] ;
 wire \top_ihp.oisc.regs[37][12] ;
 wire \top_ihp.oisc.regs[37][13] ;
 wire \top_ihp.oisc.regs[37][14] ;
 wire \top_ihp.oisc.regs[37][15] ;
 wire \top_ihp.oisc.regs[37][16] ;
 wire \top_ihp.oisc.regs[37][17] ;
 wire \top_ihp.oisc.regs[37][18] ;
 wire \top_ihp.oisc.regs[37][19] ;
 wire \top_ihp.oisc.regs[37][1] ;
 wire \top_ihp.oisc.regs[37][20] ;
 wire \top_ihp.oisc.regs[37][21] ;
 wire \top_ihp.oisc.regs[37][22] ;
 wire \top_ihp.oisc.regs[37][23] ;
 wire \top_ihp.oisc.regs[37][24] ;
 wire \top_ihp.oisc.regs[37][25] ;
 wire \top_ihp.oisc.regs[37][26] ;
 wire \top_ihp.oisc.regs[37][27] ;
 wire \top_ihp.oisc.regs[37][28] ;
 wire \top_ihp.oisc.regs[37][29] ;
 wire \top_ihp.oisc.regs[37][2] ;
 wire \top_ihp.oisc.regs[37][30] ;
 wire \top_ihp.oisc.regs[37][31] ;
 wire \top_ihp.oisc.regs[37][3] ;
 wire \top_ihp.oisc.regs[37][4] ;
 wire \top_ihp.oisc.regs[37][5] ;
 wire \top_ihp.oisc.regs[37][6] ;
 wire \top_ihp.oisc.regs[37][7] ;
 wire \top_ihp.oisc.regs[37][8] ;
 wire \top_ihp.oisc.regs[37][9] ;
 wire \top_ihp.oisc.regs[38][0] ;
 wire \top_ihp.oisc.regs[38][10] ;
 wire \top_ihp.oisc.regs[38][11] ;
 wire \top_ihp.oisc.regs[38][12] ;
 wire \top_ihp.oisc.regs[38][13] ;
 wire \top_ihp.oisc.regs[38][14] ;
 wire \top_ihp.oisc.regs[38][15] ;
 wire \top_ihp.oisc.regs[38][16] ;
 wire \top_ihp.oisc.regs[38][17] ;
 wire \top_ihp.oisc.regs[38][18] ;
 wire \top_ihp.oisc.regs[38][19] ;
 wire \top_ihp.oisc.regs[38][1] ;
 wire \top_ihp.oisc.regs[38][20] ;
 wire \top_ihp.oisc.regs[38][21] ;
 wire \top_ihp.oisc.regs[38][22] ;
 wire \top_ihp.oisc.regs[38][23] ;
 wire \top_ihp.oisc.regs[38][24] ;
 wire \top_ihp.oisc.regs[38][25] ;
 wire \top_ihp.oisc.regs[38][26] ;
 wire \top_ihp.oisc.regs[38][27] ;
 wire \top_ihp.oisc.regs[38][28] ;
 wire \top_ihp.oisc.regs[38][29] ;
 wire \top_ihp.oisc.regs[38][2] ;
 wire \top_ihp.oisc.regs[38][30] ;
 wire \top_ihp.oisc.regs[38][31] ;
 wire \top_ihp.oisc.regs[38][3] ;
 wire \top_ihp.oisc.regs[38][4] ;
 wire \top_ihp.oisc.regs[38][5] ;
 wire \top_ihp.oisc.regs[38][6] ;
 wire \top_ihp.oisc.regs[38][7] ;
 wire \top_ihp.oisc.regs[38][8] ;
 wire \top_ihp.oisc.regs[38][9] ;
 wire \top_ihp.oisc.regs[39][0] ;
 wire \top_ihp.oisc.regs[39][10] ;
 wire \top_ihp.oisc.regs[39][11] ;
 wire \top_ihp.oisc.regs[39][12] ;
 wire \top_ihp.oisc.regs[39][13] ;
 wire \top_ihp.oisc.regs[39][14] ;
 wire \top_ihp.oisc.regs[39][15] ;
 wire \top_ihp.oisc.regs[39][16] ;
 wire \top_ihp.oisc.regs[39][17] ;
 wire \top_ihp.oisc.regs[39][18] ;
 wire \top_ihp.oisc.regs[39][19] ;
 wire \top_ihp.oisc.regs[39][1] ;
 wire \top_ihp.oisc.regs[39][20] ;
 wire \top_ihp.oisc.regs[39][21] ;
 wire \top_ihp.oisc.regs[39][22] ;
 wire \top_ihp.oisc.regs[39][23] ;
 wire \top_ihp.oisc.regs[39][24] ;
 wire \top_ihp.oisc.regs[39][25] ;
 wire \top_ihp.oisc.regs[39][26] ;
 wire \top_ihp.oisc.regs[39][27] ;
 wire \top_ihp.oisc.regs[39][28] ;
 wire \top_ihp.oisc.regs[39][29] ;
 wire \top_ihp.oisc.regs[39][2] ;
 wire \top_ihp.oisc.regs[39][30] ;
 wire \top_ihp.oisc.regs[39][31] ;
 wire \top_ihp.oisc.regs[39][3] ;
 wire \top_ihp.oisc.regs[39][4] ;
 wire \top_ihp.oisc.regs[39][5] ;
 wire \top_ihp.oisc.regs[39][6] ;
 wire \top_ihp.oisc.regs[39][7] ;
 wire \top_ihp.oisc.regs[39][8] ;
 wire \top_ihp.oisc.regs[39][9] ;
 wire \top_ihp.oisc.regs[3][0] ;
 wire \top_ihp.oisc.regs[3][10] ;
 wire \top_ihp.oisc.regs[3][11] ;
 wire \top_ihp.oisc.regs[3][12] ;
 wire \top_ihp.oisc.regs[3][13] ;
 wire \top_ihp.oisc.regs[3][14] ;
 wire \top_ihp.oisc.regs[3][15] ;
 wire \top_ihp.oisc.regs[3][16] ;
 wire \top_ihp.oisc.regs[3][17] ;
 wire \top_ihp.oisc.regs[3][18] ;
 wire \top_ihp.oisc.regs[3][19] ;
 wire \top_ihp.oisc.regs[3][1] ;
 wire \top_ihp.oisc.regs[3][20] ;
 wire \top_ihp.oisc.regs[3][21] ;
 wire \top_ihp.oisc.regs[3][22] ;
 wire \top_ihp.oisc.regs[3][23] ;
 wire \top_ihp.oisc.regs[3][24] ;
 wire \top_ihp.oisc.regs[3][25] ;
 wire \top_ihp.oisc.regs[3][26] ;
 wire \top_ihp.oisc.regs[3][27] ;
 wire \top_ihp.oisc.regs[3][28] ;
 wire \top_ihp.oisc.regs[3][29] ;
 wire \top_ihp.oisc.regs[3][2] ;
 wire \top_ihp.oisc.regs[3][30] ;
 wire \top_ihp.oisc.regs[3][31] ;
 wire \top_ihp.oisc.regs[3][3] ;
 wire \top_ihp.oisc.regs[3][4] ;
 wire \top_ihp.oisc.regs[3][5] ;
 wire \top_ihp.oisc.regs[3][6] ;
 wire \top_ihp.oisc.regs[3][7] ;
 wire \top_ihp.oisc.regs[3][8] ;
 wire \top_ihp.oisc.regs[3][9] ;
 wire \top_ihp.oisc.regs[40][0] ;
 wire \top_ihp.oisc.regs[40][10] ;
 wire \top_ihp.oisc.regs[40][11] ;
 wire \top_ihp.oisc.regs[40][12] ;
 wire \top_ihp.oisc.regs[40][13] ;
 wire \top_ihp.oisc.regs[40][14] ;
 wire \top_ihp.oisc.regs[40][15] ;
 wire \top_ihp.oisc.regs[40][16] ;
 wire \top_ihp.oisc.regs[40][17] ;
 wire \top_ihp.oisc.regs[40][18] ;
 wire \top_ihp.oisc.regs[40][19] ;
 wire \top_ihp.oisc.regs[40][1] ;
 wire \top_ihp.oisc.regs[40][20] ;
 wire \top_ihp.oisc.regs[40][21] ;
 wire \top_ihp.oisc.regs[40][22] ;
 wire \top_ihp.oisc.regs[40][23] ;
 wire \top_ihp.oisc.regs[40][24] ;
 wire \top_ihp.oisc.regs[40][25] ;
 wire \top_ihp.oisc.regs[40][26] ;
 wire \top_ihp.oisc.regs[40][27] ;
 wire \top_ihp.oisc.regs[40][28] ;
 wire \top_ihp.oisc.regs[40][29] ;
 wire \top_ihp.oisc.regs[40][2] ;
 wire \top_ihp.oisc.regs[40][30] ;
 wire \top_ihp.oisc.regs[40][31] ;
 wire \top_ihp.oisc.regs[40][3] ;
 wire \top_ihp.oisc.regs[40][4] ;
 wire \top_ihp.oisc.regs[40][5] ;
 wire \top_ihp.oisc.regs[40][6] ;
 wire \top_ihp.oisc.regs[40][7] ;
 wire \top_ihp.oisc.regs[40][8] ;
 wire \top_ihp.oisc.regs[40][9] ;
 wire \top_ihp.oisc.regs[41][0] ;
 wire \top_ihp.oisc.regs[41][10] ;
 wire \top_ihp.oisc.regs[41][11] ;
 wire \top_ihp.oisc.regs[41][12] ;
 wire \top_ihp.oisc.regs[41][13] ;
 wire \top_ihp.oisc.regs[41][14] ;
 wire \top_ihp.oisc.regs[41][15] ;
 wire \top_ihp.oisc.regs[41][16] ;
 wire \top_ihp.oisc.regs[41][17] ;
 wire \top_ihp.oisc.regs[41][18] ;
 wire \top_ihp.oisc.regs[41][19] ;
 wire \top_ihp.oisc.regs[41][1] ;
 wire \top_ihp.oisc.regs[41][20] ;
 wire \top_ihp.oisc.regs[41][21] ;
 wire \top_ihp.oisc.regs[41][22] ;
 wire \top_ihp.oisc.regs[41][23] ;
 wire \top_ihp.oisc.regs[41][24] ;
 wire \top_ihp.oisc.regs[41][25] ;
 wire \top_ihp.oisc.regs[41][26] ;
 wire \top_ihp.oisc.regs[41][27] ;
 wire \top_ihp.oisc.regs[41][28] ;
 wire \top_ihp.oisc.regs[41][29] ;
 wire \top_ihp.oisc.regs[41][2] ;
 wire \top_ihp.oisc.regs[41][30] ;
 wire \top_ihp.oisc.regs[41][31] ;
 wire \top_ihp.oisc.regs[41][3] ;
 wire \top_ihp.oisc.regs[41][4] ;
 wire \top_ihp.oisc.regs[41][5] ;
 wire \top_ihp.oisc.regs[41][6] ;
 wire \top_ihp.oisc.regs[41][7] ;
 wire \top_ihp.oisc.regs[41][8] ;
 wire \top_ihp.oisc.regs[41][9] ;
 wire \top_ihp.oisc.regs[42][0] ;
 wire \top_ihp.oisc.regs[42][10] ;
 wire \top_ihp.oisc.regs[42][11] ;
 wire \top_ihp.oisc.regs[42][12] ;
 wire \top_ihp.oisc.regs[42][13] ;
 wire \top_ihp.oisc.regs[42][14] ;
 wire \top_ihp.oisc.regs[42][15] ;
 wire \top_ihp.oisc.regs[42][16] ;
 wire \top_ihp.oisc.regs[42][17] ;
 wire \top_ihp.oisc.regs[42][18] ;
 wire \top_ihp.oisc.regs[42][19] ;
 wire \top_ihp.oisc.regs[42][1] ;
 wire \top_ihp.oisc.regs[42][20] ;
 wire \top_ihp.oisc.regs[42][21] ;
 wire \top_ihp.oisc.regs[42][22] ;
 wire \top_ihp.oisc.regs[42][23] ;
 wire \top_ihp.oisc.regs[42][24] ;
 wire \top_ihp.oisc.regs[42][25] ;
 wire \top_ihp.oisc.regs[42][26] ;
 wire \top_ihp.oisc.regs[42][27] ;
 wire \top_ihp.oisc.regs[42][28] ;
 wire \top_ihp.oisc.regs[42][29] ;
 wire \top_ihp.oisc.regs[42][2] ;
 wire \top_ihp.oisc.regs[42][30] ;
 wire \top_ihp.oisc.regs[42][31] ;
 wire \top_ihp.oisc.regs[42][3] ;
 wire \top_ihp.oisc.regs[42][4] ;
 wire \top_ihp.oisc.regs[42][5] ;
 wire \top_ihp.oisc.regs[42][6] ;
 wire \top_ihp.oisc.regs[42][7] ;
 wire \top_ihp.oisc.regs[42][8] ;
 wire \top_ihp.oisc.regs[42][9] ;
 wire \top_ihp.oisc.regs[43][0] ;
 wire \top_ihp.oisc.regs[43][10] ;
 wire \top_ihp.oisc.regs[43][11] ;
 wire \top_ihp.oisc.regs[43][12] ;
 wire \top_ihp.oisc.regs[43][13] ;
 wire \top_ihp.oisc.regs[43][14] ;
 wire \top_ihp.oisc.regs[43][15] ;
 wire \top_ihp.oisc.regs[43][16] ;
 wire \top_ihp.oisc.regs[43][17] ;
 wire \top_ihp.oisc.regs[43][18] ;
 wire \top_ihp.oisc.regs[43][19] ;
 wire \top_ihp.oisc.regs[43][1] ;
 wire \top_ihp.oisc.regs[43][20] ;
 wire \top_ihp.oisc.regs[43][21] ;
 wire \top_ihp.oisc.regs[43][22] ;
 wire \top_ihp.oisc.regs[43][23] ;
 wire \top_ihp.oisc.regs[43][24] ;
 wire \top_ihp.oisc.regs[43][25] ;
 wire \top_ihp.oisc.regs[43][26] ;
 wire \top_ihp.oisc.regs[43][27] ;
 wire \top_ihp.oisc.regs[43][28] ;
 wire \top_ihp.oisc.regs[43][29] ;
 wire \top_ihp.oisc.regs[43][2] ;
 wire \top_ihp.oisc.regs[43][30] ;
 wire \top_ihp.oisc.regs[43][31] ;
 wire \top_ihp.oisc.regs[43][3] ;
 wire \top_ihp.oisc.regs[43][4] ;
 wire \top_ihp.oisc.regs[43][5] ;
 wire \top_ihp.oisc.regs[43][6] ;
 wire \top_ihp.oisc.regs[43][7] ;
 wire \top_ihp.oisc.regs[43][8] ;
 wire \top_ihp.oisc.regs[43][9] ;
 wire \top_ihp.oisc.regs[44][0] ;
 wire \top_ihp.oisc.regs[44][10] ;
 wire \top_ihp.oisc.regs[44][11] ;
 wire \top_ihp.oisc.regs[44][12] ;
 wire \top_ihp.oisc.regs[44][13] ;
 wire \top_ihp.oisc.regs[44][14] ;
 wire \top_ihp.oisc.regs[44][15] ;
 wire \top_ihp.oisc.regs[44][16] ;
 wire \top_ihp.oisc.regs[44][17] ;
 wire \top_ihp.oisc.regs[44][18] ;
 wire \top_ihp.oisc.regs[44][19] ;
 wire \top_ihp.oisc.regs[44][1] ;
 wire \top_ihp.oisc.regs[44][20] ;
 wire \top_ihp.oisc.regs[44][21] ;
 wire \top_ihp.oisc.regs[44][22] ;
 wire \top_ihp.oisc.regs[44][23] ;
 wire \top_ihp.oisc.regs[44][24] ;
 wire \top_ihp.oisc.regs[44][25] ;
 wire \top_ihp.oisc.regs[44][26] ;
 wire \top_ihp.oisc.regs[44][27] ;
 wire \top_ihp.oisc.regs[44][28] ;
 wire \top_ihp.oisc.regs[44][29] ;
 wire \top_ihp.oisc.regs[44][2] ;
 wire \top_ihp.oisc.regs[44][30] ;
 wire \top_ihp.oisc.regs[44][31] ;
 wire \top_ihp.oisc.regs[44][3] ;
 wire \top_ihp.oisc.regs[44][4] ;
 wire \top_ihp.oisc.regs[44][5] ;
 wire \top_ihp.oisc.regs[44][6] ;
 wire \top_ihp.oisc.regs[44][7] ;
 wire \top_ihp.oisc.regs[44][8] ;
 wire \top_ihp.oisc.regs[44][9] ;
 wire \top_ihp.oisc.regs[45][0] ;
 wire \top_ihp.oisc.regs[45][10] ;
 wire \top_ihp.oisc.regs[45][11] ;
 wire \top_ihp.oisc.regs[45][12] ;
 wire \top_ihp.oisc.regs[45][13] ;
 wire \top_ihp.oisc.regs[45][14] ;
 wire \top_ihp.oisc.regs[45][15] ;
 wire \top_ihp.oisc.regs[45][16] ;
 wire \top_ihp.oisc.regs[45][17] ;
 wire \top_ihp.oisc.regs[45][18] ;
 wire \top_ihp.oisc.regs[45][19] ;
 wire \top_ihp.oisc.regs[45][1] ;
 wire \top_ihp.oisc.regs[45][20] ;
 wire \top_ihp.oisc.regs[45][21] ;
 wire \top_ihp.oisc.regs[45][22] ;
 wire \top_ihp.oisc.regs[45][23] ;
 wire \top_ihp.oisc.regs[45][24] ;
 wire \top_ihp.oisc.regs[45][25] ;
 wire \top_ihp.oisc.regs[45][26] ;
 wire \top_ihp.oisc.regs[45][27] ;
 wire \top_ihp.oisc.regs[45][28] ;
 wire \top_ihp.oisc.regs[45][29] ;
 wire \top_ihp.oisc.regs[45][2] ;
 wire \top_ihp.oisc.regs[45][30] ;
 wire \top_ihp.oisc.regs[45][31] ;
 wire \top_ihp.oisc.regs[45][3] ;
 wire \top_ihp.oisc.regs[45][4] ;
 wire \top_ihp.oisc.regs[45][5] ;
 wire \top_ihp.oisc.regs[45][6] ;
 wire \top_ihp.oisc.regs[45][7] ;
 wire \top_ihp.oisc.regs[45][8] ;
 wire \top_ihp.oisc.regs[45][9] ;
 wire \top_ihp.oisc.regs[46][0] ;
 wire \top_ihp.oisc.regs[46][10] ;
 wire \top_ihp.oisc.regs[46][11] ;
 wire \top_ihp.oisc.regs[46][12] ;
 wire \top_ihp.oisc.regs[46][13] ;
 wire \top_ihp.oisc.regs[46][14] ;
 wire \top_ihp.oisc.regs[46][15] ;
 wire \top_ihp.oisc.regs[46][16] ;
 wire \top_ihp.oisc.regs[46][17] ;
 wire \top_ihp.oisc.regs[46][18] ;
 wire \top_ihp.oisc.regs[46][19] ;
 wire \top_ihp.oisc.regs[46][1] ;
 wire \top_ihp.oisc.regs[46][20] ;
 wire \top_ihp.oisc.regs[46][21] ;
 wire \top_ihp.oisc.regs[46][22] ;
 wire \top_ihp.oisc.regs[46][23] ;
 wire \top_ihp.oisc.regs[46][24] ;
 wire \top_ihp.oisc.regs[46][25] ;
 wire \top_ihp.oisc.regs[46][26] ;
 wire \top_ihp.oisc.regs[46][27] ;
 wire \top_ihp.oisc.regs[46][28] ;
 wire \top_ihp.oisc.regs[46][29] ;
 wire \top_ihp.oisc.regs[46][2] ;
 wire \top_ihp.oisc.regs[46][30] ;
 wire \top_ihp.oisc.regs[46][31] ;
 wire \top_ihp.oisc.regs[46][3] ;
 wire \top_ihp.oisc.regs[46][4] ;
 wire \top_ihp.oisc.regs[46][5] ;
 wire \top_ihp.oisc.regs[46][6] ;
 wire \top_ihp.oisc.regs[46][7] ;
 wire \top_ihp.oisc.regs[46][8] ;
 wire \top_ihp.oisc.regs[46][9] ;
 wire \top_ihp.oisc.regs[47][0] ;
 wire \top_ihp.oisc.regs[47][10] ;
 wire \top_ihp.oisc.regs[47][11] ;
 wire \top_ihp.oisc.regs[47][12] ;
 wire \top_ihp.oisc.regs[47][13] ;
 wire \top_ihp.oisc.regs[47][14] ;
 wire \top_ihp.oisc.regs[47][15] ;
 wire \top_ihp.oisc.regs[47][16] ;
 wire \top_ihp.oisc.regs[47][17] ;
 wire \top_ihp.oisc.regs[47][18] ;
 wire \top_ihp.oisc.regs[47][19] ;
 wire \top_ihp.oisc.regs[47][1] ;
 wire \top_ihp.oisc.regs[47][20] ;
 wire \top_ihp.oisc.regs[47][21] ;
 wire \top_ihp.oisc.regs[47][22] ;
 wire \top_ihp.oisc.regs[47][23] ;
 wire \top_ihp.oisc.regs[47][24] ;
 wire \top_ihp.oisc.regs[47][25] ;
 wire \top_ihp.oisc.regs[47][26] ;
 wire \top_ihp.oisc.regs[47][27] ;
 wire \top_ihp.oisc.regs[47][28] ;
 wire \top_ihp.oisc.regs[47][29] ;
 wire \top_ihp.oisc.regs[47][2] ;
 wire \top_ihp.oisc.regs[47][30] ;
 wire \top_ihp.oisc.regs[47][31] ;
 wire \top_ihp.oisc.regs[47][3] ;
 wire \top_ihp.oisc.regs[47][4] ;
 wire \top_ihp.oisc.regs[47][5] ;
 wire \top_ihp.oisc.regs[47][6] ;
 wire \top_ihp.oisc.regs[47][7] ;
 wire \top_ihp.oisc.regs[47][8] ;
 wire \top_ihp.oisc.regs[47][9] ;
 wire \top_ihp.oisc.regs[48][0] ;
 wire \top_ihp.oisc.regs[48][10] ;
 wire \top_ihp.oisc.regs[48][11] ;
 wire \top_ihp.oisc.regs[48][12] ;
 wire \top_ihp.oisc.regs[48][13] ;
 wire \top_ihp.oisc.regs[48][14] ;
 wire \top_ihp.oisc.regs[48][15] ;
 wire \top_ihp.oisc.regs[48][16] ;
 wire \top_ihp.oisc.regs[48][17] ;
 wire \top_ihp.oisc.regs[48][18] ;
 wire \top_ihp.oisc.regs[48][19] ;
 wire \top_ihp.oisc.regs[48][1] ;
 wire \top_ihp.oisc.regs[48][20] ;
 wire \top_ihp.oisc.regs[48][21] ;
 wire \top_ihp.oisc.regs[48][22] ;
 wire \top_ihp.oisc.regs[48][23] ;
 wire \top_ihp.oisc.regs[48][24] ;
 wire \top_ihp.oisc.regs[48][25] ;
 wire \top_ihp.oisc.regs[48][26] ;
 wire \top_ihp.oisc.regs[48][27] ;
 wire \top_ihp.oisc.regs[48][28] ;
 wire \top_ihp.oisc.regs[48][29] ;
 wire \top_ihp.oisc.regs[48][2] ;
 wire \top_ihp.oisc.regs[48][30] ;
 wire \top_ihp.oisc.regs[48][31] ;
 wire \top_ihp.oisc.regs[48][3] ;
 wire \top_ihp.oisc.regs[48][4] ;
 wire \top_ihp.oisc.regs[48][5] ;
 wire \top_ihp.oisc.regs[48][6] ;
 wire \top_ihp.oisc.regs[48][7] ;
 wire \top_ihp.oisc.regs[48][8] ;
 wire \top_ihp.oisc.regs[48][9] ;
 wire \top_ihp.oisc.regs[49][0] ;
 wire \top_ihp.oisc.regs[49][10] ;
 wire \top_ihp.oisc.regs[49][11] ;
 wire \top_ihp.oisc.regs[49][12] ;
 wire \top_ihp.oisc.regs[49][13] ;
 wire \top_ihp.oisc.regs[49][14] ;
 wire \top_ihp.oisc.regs[49][15] ;
 wire \top_ihp.oisc.regs[49][16] ;
 wire \top_ihp.oisc.regs[49][17] ;
 wire \top_ihp.oisc.regs[49][18] ;
 wire \top_ihp.oisc.regs[49][19] ;
 wire \top_ihp.oisc.regs[49][1] ;
 wire \top_ihp.oisc.regs[49][20] ;
 wire \top_ihp.oisc.regs[49][21] ;
 wire \top_ihp.oisc.regs[49][22] ;
 wire \top_ihp.oisc.regs[49][23] ;
 wire \top_ihp.oisc.regs[49][24] ;
 wire \top_ihp.oisc.regs[49][25] ;
 wire \top_ihp.oisc.regs[49][26] ;
 wire \top_ihp.oisc.regs[49][27] ;
 wire \top_ihp.oisc.regs[49][28] ;
 wire \top_ihp.oisc.regs[49][29] ;
 wire \top_ihp.oisc.regs[49][2] ;
 wire \top_ihp.oisc.regs[49][30] ;
 wire \top_ihp.oisc.regs[49][31] ;
 wire \top_ihp.oisc.regs[49][3] ;
 wire \top_ihp.oisc.regs[49][4] ;
 wire \top_ihp.oisc.regs[49][5] ;
 wire \top_ihp.oisc.regs[49][6] ;
 wire \top_ihp.oisc.regs[49][7] ;
 wire \top_ihp.oisc.regs[49][8] ;
 wire \top_ihp.oisc.regs[49][9] ;
 wire \top_ihp.oisc.regs[4][0] ;
 wire \top_ihp.oisc.regs[4][10] ;
 wire \top_ihp.oisc.regs[4][11] ;
 wire \top_ihp.oisc.regs[4][12] ;
 wire \top_ihp.oisc.regs[4][13] ;
 wire \top_ihp.oisc.regs[4][14] ;
 wire \top_ihp.oisc.regs[4][15] ;
 wire \top_ihp.oisc.regs[4][16] ;
 wire \top_ihp.oisc.regs[4][17] ;
 wire \top_ihp.oisc.regs[4][18] ;
 wire \top_ihp.oisc.regs[4][19] ;
 wire \top_ihp.oisc.regs[4][1] ;
 wire \top_ihp.oisc.regs[4][20] ;
 wire \top_ihp.oisc.regs[4][21] ;
 wire \top_ihp.oisc.regs[4][22] ;
 wire \top_ihp.oisc.regs[4][23] ;
 wire \top_ihp.oisc.regs[4][24] ;
 wire \top_ihp.oisc.regs[4][25] ;
 wire \top_ihp.oisc.regs[4][26] ;
 wire \top_ihp.oisc.regs[4][27] ;
 wire \top_ihp.oisc.regs[4][28] ;
 wire \top_ihp.oisc.regs[4][29] ;
 wire \top_ihp.oisc.regs[4][2] ;
 wire \top_ihp.oisc.regs[4][30] ;
 wire \top_ihp.oisc.regs[4][31] ;
 wire \top_ihp.oisc.regs[4][3] ;
 wire \top_ihp.oisc.regs[4][4] ;
 wire \top_ihp.oisc.regs[4][5] ;
 wire \top_ihp.oisc.regs[4][6] ;
 wire \top_ihp.oisc.regs[4][7] ;
 wire \top_ihp.oisc.regs[4][8] ;
 wire \top_ihp.oisc.regs[4][9] ;
 wire \top_ihp.oisc.regs[50][0] ;
 wire \top_ihp.oisc.regs[50][10] ;
 wire \top_ihp.oisc.regs[50][11] ;
 wire \top_ihp.oisc.regs[50][12] ;
 wire \top_ihp.oisc.regs[50][13] ;
 wire \top_ihp.oisc.regs[50][14] ;
 wire \top_ihp.oisc.regs[50][15] ;
 wire \top_ihp.oisc.regs[50][16] ;
 wire \top_ihp.oisc.regs[50][17] ;
 wire \top_ihp.oisc.regs[50][18] ;
 wire \top_ihp.oisc.regs[50][19] ;
 wire \top_ihp.oisc.regs[50][1] ;
 wire \top_ihp.oisc.regs[50][20] ;
 wire \top_ihp.oisc.regs[50][21] ;
 wire \top_ihp.oisc.regs[50][22] ;
 wire \top_ihp.oisc.regs[50][23] ;
 wire \top_ihp.oisc.regs[50][24] ;
 wire \top_ihp.oisc.regs[50][25] ;
 wire \top_ihp.oisc.regs[50][26] ;
 wire \top_ihp.oisc.regs[50][27] ;
 wire \top_ihp.oisc.regs[50][28] ;
 wire \top_ihp.oisc.regs[50][29] ;
 wire \top_ihp.oisc.regs[50][2] ;
 wire \top_ihp.oisc.regs[50][30] ;
 wire \top_ihp.oisc.regs[50][31] ;
 wire \top_ihp.oisc.regs[50][3] ;
 wire \top_ihp.oisc.regs[50][4] ;
 wire \top_ihp.oisc.regs[50][5] ;
 wire \top_ihp.oisc.regs[50][6] ;
 wire \top_ihp.oisc.regs[50][7] ;
 wire \top_ihp.oisc.regs[50][8] ;
 wire \top_ihp.oisc.regs[50][9] ;
 wire \top_ihp.oisc.regs[51][0] ;
 wire \top_ihp.oisc.regs[51][10] ;
 wire \top_ihp.oisc.regs[51][11] ;
 wire \top_ihp.oisc.regs[51][12] ;
 wire \top_ihp.oisc.regs[51][13] ;
 wire \top_ihp.oisc.regs[51][14] ;
 wire \top_ihp.oisc.regs[51][15] ;
 wire \top_ihp.oisc.regs[51][16] ;
 wire \top_ihp.oisc.regs[51][17] ;
 wire \top_ihp.oisc.regs[51][18] ;
 wire \top_ihp.oisc.regs[51][19] ;
 wire \top_ihp.oisc.regs[51][1] ;
 wire \top_ihp.oisc.regs[51][20] ;
 wire \top_ihp.oisc.regs[51][21] ;
 wire \top_ihp.oisc.regs[51][22] ;
 wire \top_ihp.oisc.regs[51][23] ;
 wire \top_ihp.oisc.regs[51][24] ;
 wire \top_ihp.oisc.regs[51][25] ;
 wire \top_ihp.oisc.regs[51][26] ;
 wire \top_ihp.oisc.regs[51][27] ;
 wire \top_ihp.oisc.regs[51][28] ;
 wire \top_ihp.oisc.regs[51][29] ;
 wire \top_ihp.oisc.regs[51][2] ;
 wire \top_ihp.oisc.regs[51][30] ;
 wire \top_ihp.oisc.regs[51][31] ;
 wire \top_ihp.oisc.regs[51][3] ;
 wire \top_ihp.oisc.regs[51][4] ;
 wire \top_ihp.oisc.regs[51][5] ;
 wire \top_ihp.oisc.regs[51][6] ;
 wire \top_ihp.oisc.regs[51][7] ;
 wire \top_ihp.oisc.regs[51][8] ;
 wire \top_ihp.oisc.regs[51][9] ;
 wire \top_ihp.oisc.regs[52][0] ;
 wire \top_ihp.oisc.regs[52][10] ;
 wire \top_ihp.oisc.regs[52][11] ;
 wire \top_ihp.oisc.regs[52][12] ;
 wire \top_ihp.oisc.regs[52][13] ;
 wire \top_ihp.oisc.regs[52][14] ;
 wire \top_ihp.oisc.regs[52][15] ;
 wire \top_ihp.oisc.regs[52][16] ;
 wire \top_ihp.oisc.regs[52][17] ;
 wire \top_ihp.oisc.regs[52][18] ;
 wire \top_ihp.oisc.regs[52][19] ;
 wire \top_ihp.oisc.regs[52][1] ;
 wire \top_ihp.oisc.regs[52][20] ;
 wire \top_ihp.oisc.regs[52][21] ;
 wire \top_ihp.oisc.regs[52][22] ;
 wire \top_ihp.oisc.regs[52][23] ;
 wire \top_ihp.oisc.regs[52][24] ;
 wire \top_ihp.oisc.regs[52][25] ;
 wire \top_ihp.oisc.regs[52][26] ;
 wire \top_ihp.oisc.regs[52][27] ;
 wire \top_ihp.oisc.regs[52][28] ;
 wire \top_ihp.oisc.regs[52][29] ;
 wire \top_ihp.oisc.regs[52][2] ;
 wire \top_ihp.oisc.regs[52][30] ;
 wire \top_ihp.oisc.regs[52][31] ;
 wire \top_ihp.oisc.regs[52][3] ;
 wire \top_ihp.oisc.regs[52][4] ;
 wire \top_ihp.oisc.regs[52][5] ;
 wire \top_ihp.oisc.regs[52][6] ;
 wire \top_ihp.oisc.regs[52][7] ;
 wire \top_ihp.oisc.regs[52][8] ;
 wire \top_ihp.oisc.regs[52][9] ;
 wire \top_ihp.oisc.regs[53][0] ;
 wire \top_ihp.oisc.regs[53][10] ;
 wire \top_ihp.oisc.regs[53][11] ;
 wire \top_ihp.oisc.regs[53][12] ;
 wire \top_ihp.oisc.regs[53][13] ;
 wire \top_ihp.oisc.regs[53][14] ;
 wire \top_ihp.oisc.regs[53][15] ;
 wire \top_ihp.oisc.regs[53][16] ;
 wire \top_ihp.oisc.regs[53][17] ;
 wire \top_ihp.oisc.regs[53][18] ;
 wire \top_ihp.oisc.regs[53][19] ;
 wire \top_ihp.oisc.regs[53][1] ;
 wire \top_ihp.oisc.regs[53][20] ;
 wire \top_ihp.oisc.regs[53][21] ;
 wire \top_ihp.oisc.regs[53][22] ;
 wire \top_ihp.oisc.regs[53][23] ;
 wire \top_ihp.oisc.regs[53][24] ;
 wire \top_ihp.oisc.regs[53][25] ;
 wire \top_ihp.oisc.regs[53][26] ;
 wire \top_ihp.oisc.regs[53][27] ;
 wire \top_ihp.oisc.regs[53][28] ;
 wire \top_ihp.oisc.regs[53][29] ;
 wire \top_ihp.oisc.regs[53][2] ;
 wire \top_ihp.oisc.regs[53][30] ;
 wire \top_ihp.oisc.regs[53][31] ;
 wire \top_ihp.oisc.regs[53][3] ;
 wire \top_ihp.oisc.regs[53][4] ;
 wire \top_ihp.oisc.regs[53][5] ;
 wire \top_ihp.oisc.regs[53][6] ;
 wire \top_ihp.oisc.regs[53][7] ;
 wire \top_ihp.oisc.regs[53][8] ;
 wire \top_ihp.oisc.regs[53][9] ;
 wire \top_ihp.oisc.regs[54][0] ;
 wire \top_ihp.oisc.regs[54][10] ;
 wire \top_ihp.oisc.regs[54][11] ;
 wire \top_ihp.oisc.regs[54][12] ;
 wire \top_ihp.oisc.regs[54][13] ;
 wire \top_ihp.oisc.regs[54][14] ;
 wire \top_ihp.oisc.regs[54][15] ;
 wire \top_ihp.oisc.regs[54][16] ;
 wire \top_ihp.oisc.regs[54][17] ;
 wire \top_ihp.oisc.regs[54][18] ;
 wire \top_ihp.oisc.regs[54][19] ;
 wire \top_ihp.oisc.regs[54][1] ;
 wire \top_ihp.oisc.regs[54][20] ;
 wire \top_ihp.oisc.regs[54][21] ;
 wire \top_ihp.oisc.regs[54][22] ;
 wire \top_ihp.oisc.regs[54][23] ;
 wire \top_ihp.oisc.regs[54][24] ;
 wire \top_ihp.oisc.regs[54][25] ;
 wire \top_ihp.oisc.regs[54][26] ;
 wire \top_ihp.oisc.regs[54][27] ;
 wire \top_ihp.oisc.regs[54][28] ;
 wire \top_ihp.oisc.regs[54][29] ;
 wire \top_ihp.oisc.regs[54][2] ;
 wire \top_ihp.oisc.regs[54][30] ;
 wire \top_ihp.oisc.regs[54][31] ;
 wire \top_ihp.oisc.regs[54][3] ;
 wire \top_ihp.oisc.regs[54][4] ;
 wire \top_ihp.oisc.regs[54][5] ;
 wire \top_ihp.oisc.regs[54][6] ;
 wire \top_ihp.oisc.regs[54][7] ;
 wire \top_ihp.oisc.regs[54][8] ;
 wire \top_ihp.oisc.regs[54][9] ;
 wire \top_ihp.oisc.regs[55][0] ;
 wire \top_ihp.oisc.regs[55][10] ;
 wire \top_ihp.oisc.regs[55][11] ;
 wire \top_ihp.oisc.regs[55][12] ;
 wire \top_ihp.oisc.regs[55][13] ;
 wire \top_ihp.oisc.regs[55][14] ;
 wire \top_ihp.oisc.regs[55][15] ;
 wire \top_ihp.oisc.regs[55][16] ;
 wire \top_ihp.oisc.regs[55][17] ;
 wire \top_ihp.oisc.regs[55][18] ;
 wire \top_ihp.oisc.regs[55][19] ;
 wire \top_ihp.oisc.regs[55][1] ;
 wire \top_ihp.oisc.regs[55][20] ;
 wire \top_ihp.oisc.regs[55][21] ;
 wire \top_ihp.oisc.regs[55][22] ;
 wire \top_ihp.oisc.regs[55][23] ;
 wire \top_ihp.oisc.regs[55][24] ;
 wire \top_ihp.oisc.regs[55][25] ;
 wire \top_ihp.oisc.regs[55][26] ;
 wire \top_ihp.oisc.regs[55][27] ;
 wire \top_ihp.oisc.regs[55][28] ;
 wire \top_ihp.oisc.regs[55][29] ;
 wire \top_ihp.oisc.regs[55][2] ;
 wire \top_ihp.oisc.regs[55][30] ;
 wire \top_ihp.oisc.regs[55][31] ;
 wire \top_ihp.oisc.regs[55][3] ;
 wire \top_ihp.oisc.regs[55][4] ;
 wire \top_ihp.oisc.regs[55][5] ;
 wire \top_ihp.oisc.regs[55][6] ;
 wire \top_ihp.oisc.regs[55][7] ;
 wire \top_ihp.oisc.regs[55][8] ;
 wire \top_ihp.oisc.regs[55][9] ;
 wire \top_ihp.oisc.regs[56][0] ;
 wire \top_ihp.oisc.regs[56][10] ;
 wire \top_ihp.oisc.regs[56][11] ;
 wire \top_ihp.oisc.regs[56][12] ;
 wire \top_ihp.oisc.regs[56][13] ;
 wire \top_ihp.oisc.regs[56][14] ;
 wire \top_ihp.oisc.regs[56][15] ;
 wire \top_ihp.oisc.regs[56][16] ;
 wire \top_ihp.oisc.regs[56][17] ;
 wire \top_ihp.oisc.regs[56][18] ;
 wire \top_ihp.oisc.regs[56][19] ;
 wire \top_ihp.oisc.regs[56][1] ;
 wire \top_ihp.oisc.regs[56][20] ;
 wire \top_ihp.oisc.regs[56][21] ;
 wire \top_ihp.oisc.regs[56][22] ;
 wire \top_ihp.oisc.regs[56][23] ;
 wire \top_ihp.oisc.regs[56][24] ;
 wire \top_ihp.oisc.regs[56][25] ;
 wire \top_ihp.oisc.regs[56][26] ;
 wire \top_ihp.oisc.regs[56][27] ;
 wire \top_ihp.oisc.regs[56][28] ;
 wire \top_ihp.oisc.regs[56][29] ;
 wire \top_ihp.oisc.regs[56][2] ;
 wire \top_ihp.oisc.regs[56][30] ;
 wire \top_ihp.oisc.regs[56][31] ;
 wire \top_ihp.oisc.regs[56][3] ;
 wire \top_ihp.oisc.regs[56][4] ;
 wire \top_ihp.oisc.regs[56][5] ;
 wire \top_ihp.oisc.regs[56][6] ;
 wire \top_ihp.oisc.regs[56][7] ;
 wire \top_ihp.oisc.regs[56][8] ;
 wire \top_ihp.oisc.regs[56][9] ;
 wire \top_ihp.oisc.regs[57][0] ;
 wire \top_ihp.oisc.regs[57][10] ;
 wire \top_ihp.oisc.regs[57][11] ;
 wire \top_ihp.oisc.regs[57][12] ;
 wire \top_ihp.oisc.regs[57][13] ;
 wire \top_ihp.oisc.regs[57][14] ;
 wire \top_ihp.oisc.regs[57][15] ;
 wire \top_ihp.oisc.regs[57][16] ;
 wire \top_ihp.oisc.regs[57][17] ;
 wire \top_ihp.oisc.regs[57][18] ;
 wire \top_ihp.oisc.regs[57][19] ;
 wire \top_ihp.oisc.regs[57][1] ;
 wire \top_ihp.oisc.regs[57][20] ;
 wire \top_ihp.oisc.regs[57][21] ;
 wire \top_ihp.oisc.regs[57][22] ;
 wire \top_ihp.oisc.regs[57][23] ;
 wire \top_ihp.oisc.regs[57][24] ;
 wire \top_ihp.oisc.regs[57][25] ;
 wire \top_ihp.oisc.regs[57][26] ;
 wire \top_ihp.oisc.regs[57][27] ;
 wire \top_ihp.oisc.regs[57][28] ;
 wire \top_ihp.oisc.regs[57][29] ;
 wire \top_ihp.oisc.regs[57][2] ;
 wire \top_ihp.oisc.regs[57][30] ;
 wire \top_ihp.oisc.regs[57][31] ;
 wire \top_ihp.oisc.regs[57][3] ;
 wire \top_ihp.oisc.regs[57][4] ;
 wire \top_ihp.oisc.regs[57][5] ;
 wire \top_ihp.oisc.regs[57][6] ;
 wire \top_ihp.oisc.regs[57][7] ;
 wire \top_ihp.oisc.regs[57][8] ;
 wire \top_ihp.oisc.regs[57][9] ;
 wire \top_ihp.oisc.regs[58][0] ;
 wire \top_ihp.oisc.regs[58][10] ;
 wire \top_ihp.oisc.regs[58][11] ;
 wire \top_ihp.oisc.regs[58][12] ;
 wire \top_ihp.oisc.regs[58][13] ;
 wire \top_ihp.oisc.regs[58][14] ;
 wire \top_ihp.oisc.regs[58][15] ;
 wire \top_ihp.oisc.regs[58][16] ;
 wire \top_ihp.oisc.regs[58][17] ;
 wire \top_ihp.oisc.regs[58][18] ;
 wire \top_ihp.oisc.regs[58][19] ;
 wire \top_ihp.oisc.regs[58][1] ;
 wire \top_ihp.oisc.regs[58][20] ;
 wire \top_ihp.oisc.regs[58][21] ;
 wire \top_ihp.oisc.regs[58][22] ;
 wire \top_ihp.oisc.regs[58][23] ;
 wire \top_ihp.oisc.regs[58][24] ;
 wire \top_ihp.oisc.regs[58][25] ;
 wire \top_ihp.oisc.regs[58][26] ;
 wire \top_ihp.oisc.regs[58][27] ;
 wire \top_ihp.oisc.regs[58][28] ;
 wire \top_ihp.oisc.regs[58][29] ;
 wire \top_ihp.oisc.regs[58][2] ;
 wire \top_ihp.oisc.regs[58][30] ;
 wire \top_ihp.oisc.regs[58][31] ;
 wire \top_ihp.oisc.regs[58][3] ;
 wire \top_ihp.oisc.regs[58][4] ;
 wire \top_ihp.oisc.regs[58][5] ;
 wire \top_ihp.oisc.regs[58][6] ;
 wire \top_ihp.oisc.regs[58][7] ;
 wire \top_ihp.oisc.regs[58][8] ;
 wire \top_ihp.oisc.regs[58][9] ;
 wire \top_ihp.oisc.regs[59][0] ;
 wire \top_ihp.oisc.regs[59][10] ;
 wire \top_ihp.oisc.regs[59][11] ;
 wire \top_ihp.oisc.regs[59][12] ;
 wire \top_ihp.oisc.regs[59][13] ;
 wire \top_ihp.oisc.regs[59][14] ;
 wire \top_ihp.oisc.regs[59][15] ;
 wire \top_ihp.oisc.regs[59][16] ;
 wire \top_ihp.oisc.regs[59][17] ;
 wire \top_ihp.oisc.regs[59][18] ;
 wire \top_ihp.oisc.regs[59][19] ;
 wire \top_ihp.oisc.regs[59][1] ;
 wire \top_ihp.oisc.regs[59][20] ;
 wire \top_ihp.oisc.regs[59][21] ;
 wire \top_ihp.oisc.regs[59][22] ;
 wire \top_ihp.oisc.regs[59][23] ;
 wire \top_ihp.oisc.regs[59][24] ;
 wire \top_ihp.oisc.regs[59][25] ;
 wire \top_ihp.oisc.regs[59][26] ;
 wire \top_ihp.oisc.regs[59][27] ;
 wire \top_ihp.oisc.regs[59][28] ;
 wire \top_ihp.oisc.regs[59][29] ;
 wire \top_ihp.oisc.regs[59][2] ;
 wire \top_ihp.oisc.regs[59][30] ;
 wire \top_ihp.oisc.regs[59][31] ;
 wire \top_ihp.oisc.regs[59][3] ;
 wire \top_ihp.oisc.regs[59][4] ;
 wire \top_ihp.oisc.regs[59][5] ;
 wire \top_ihp.oisc.regs[59][6] ;
 wire \top_ihp.oisc.regs[59][7] ;
 wire \top_ihp.oisc.regs[59][8] ;
 wire \top_ihp.oisc.regs[59][9] ;
 wire \top_ihp.oisc.regs[5][0] ;
 wire \top_ihp.oisc.regs[5][10] ;
 wire \top_ihp.oisc.regs[5][11] ;
 wire \top_ihp.oisc.regs[5][12] ;
 wire \top_ihp.oisc.regs[5][13] ;
 wire \top_ihp.oisc.regs[5][14] ;
 wire \top_ihp.oisc.regs[5][15] ;
 wire \top_ihp.oisc.regs[5][16] ;
 wire \top_ihp.oisc.regs[5][17] ;
 wire \top_ihp.oisc.regs[5][18] ;
 wire \top_ihp.oisc.regs[5][19] ;
 wire \top_ihp.oisc.regs[5][1] ;
 wire \top_ihp.oisc.regs[5][20] ;
 wire \top_ihp.oisc.regs[5][21] ;
 wire \top_ihp.oisc.regs[5][22] ;
 wire \top_ihp.oisc.regs[5][23] ;
 wire \top_ihp.oisc.regs[5][24] ;
 wire \top_ihp.oisc.regs[5][25] ;
 wire \top_ihp.oisc.regs[5][26] ;
 wire \top_ihp.oisc.regs[5][27] ;
 wire \top_ihp.oisc.regs[5][28] ;
 wire \top_ihp.oisc.regs[5][29] ;
 wire \top_ihp.oisc.regs[5][2] ;
 wire \top_ihp.oisc.regs[5][30] ;
 wire \top_ihp.oisc.regs[5][31] ;
 wire \top_ihp.oisc.regs[5][3] ;
 wire \top_ihp.oisc.regs[5][4] ;
 wire \top_ihp.oisc.regs[5][5] ;
 wire \top_ihp.oisc.regs[5][6] ;
 wire \top_ihp.oisc.regs[5][7] ;
 wire \top_ihp.oisc.regs[5][8] ;
 wire \top_ihp.oisc.regs[5][9] ;
 wire \top_ihp.oisc.regs[60][0] ;
 wire \top_ihp.oisc.regs[60][10] ;
 wire \top_ihp.oisc.regs[60][11] ;
 wire \top_ihp.oisc.regs[60][12] ;
 wire \top_ihp.oisc.regs[60][13] ;
 wire \top_ihp.oisc.regs[60][14] ;
 wire \top_ihp.oisc.regs[60][15] ;
 wire \top_ihp.oisc.regs[60][16] ;
 wire \top_ihp.oisc.regs[60][17] ;
 wire \top_ihp.oisc.regs[60][18] ;
 wire \top_ihp.oisc.regs[60][19] ;
 wire \top_ihp.oisc.regs[60][1] ;
 wire \top_ihp.oisc.regs[60][20] ;
 wire \top_ihp.oisc.regs[60][21] ;
 wire \top_ihp.oisc.regs[60][22] ;
 wire \top_ihp.oisc.regs[60][23] ;
 wire \top_ihp.oisc.regs[60][24] ;
 wire \top_ihp.oisc.regs[60][25] ;
 wire \top_ihp.oisc.regs[60][26] ;
 wire \top_ihp.oisc.regs[60][27] ;
 wire \top_ihp.oisc.regs[60][28] ;
 wire \top_ihp.oisc.regs[60][29] ;
 wire \top_ihp.oisc.regs[60][2] ;
 wire \top_ihp.oisc.regs[60][30] ;
 wire \top_ihp.oisc.regs[60][31] ;
 wire \top_ihp.oisc.regs[60][3] ;
 wire \top_ihp.oisc.regs[60][4] ;
 wire \top_ihp.oisc.regs[60][5] ;
 wire \top_ihp.oisc.regs[60][6] ;
 wire \top_ihp.oisc.regs[60][7] ;
 wire \top_ihp.oisc.regs[60][8] ;
 wire \top_ihp.oisc.regs[60][9] ;
 wire \top_ihp.oisc.regs[61][0] ;
 wire \top_ihp.oisc.regs[61][10] ;
 wire \top_ihp.oisc.regs[61][11] ;
 wire \top_ihp.oisc.regs[61][12] ;
 wire \top_ihp.oisc.regs[61][13] ;
 wire \top_ihp.oisc.regs[61][14] ;
 wire \top_ihp.oisc.regs[61][15] ;
 wire \top_ihp.oisc.regs[61][16] ;
 wire \top_ihp.oisc.regs[61][17] ;
 wire \top_ihp.oisc.regs[61][18] ;
 wire \top_ihp.oisc.regs[61][19] ;
 wire \top_ihp.oisc.regs[61][1] ;
 wire \top_ihp.oisc.regs[61][20] ;
 wire \top_ihp.oisc.regs[61][21] ;
 wire \top_ihp.oisc.regs[61][22] ;
 wire \top_ihp.oisc.regs[61][23] ;
 wire \top_ihp.oisc.regs[61][24] ;
 wire \top_ihp.oisc.regs[61][25] ;
 wire \top_ihp.oisc.regs[61][26] ;
 wire \top_ihp.oisc.regs[61][27] ;
 wire \top_ihp.oisc.regs[61][28] ;
 wire \top_ihp.oisc.regs[61][29] ;
 wire \top_ihp.oisc.regs[61][2] ;
 wire \top_ihp.oisc.regs[61][30] ;
 wire \top_ihp.oisc.regs[61][31] ;
 wire \top_ihp.oisc.regs[61][3] ;
 wire \top_ihp.oisc.regs[61][4] ;
 wire \top_ihp.oisc.regs[61][5] ;
 wire \top_ihp.oisc.regs[61][6] ;
 wire \top_ihp.oisc.regs[61][7] ;
 wire \top_ihp.oisc.regs[61][8] ;
 wire \top_ihp.oisc.regs[61][9] ;
 wire \top_ihp.oisc.regs[62][0] ;
 wire \top_ihp.oisc.regs[62][10] ;
 wire \top_ihp.oisc.regs[62][11] ;
 wire \top_ihp.oisc.regs[62][12] ;
 wire \top_ihp.oisc.regs[62][13] ;
 wire \top_ihp.oisc.regs[62][14] ;
 wire \top_ihp.oisc.regs[62][15] ;
 wire \top_ihp.oisc.regs[62][16] ;
 wire \top_ihp.oisc.regs[62][17] ;
 wire \top_ihp.oisc.regs[62][18] ;
 wire \top_ihp.oisc.regs[62][19] ;
 wire \top_ihp.oisc.regs[62][1] ;
 wire \top_ihp.oisc.regs[62][20] ;
 wire \top_ihp.oisc.regs[62][21] ;
 wire \top_ihp.oisc.regs[62][22] ;
 wire \top_ihp.oisc.regs[62][23] ;
 wire \top_ihp.oisc.regs[62][24] ;
 wire \top_ihp.oisc.regs[62][25] ;
 wire \top_ihp.oisc.regs[62][26] ;
 wire \top_ihp.oisc.regs[62][27] ;
 wire \top_ihp.oisc.regs[62][28] ;
 wire \top_ihp.oisc.regs[62][29] ;
 wire \top_ihp.oisc.regs[62][2] ;
 wire \top_ihp.oisc.regs[62][30] ;
 wire \top_ihp.oisc.regs[62][31] ;
 wire \top_ihp.oisc.regs[62][3] ;
 wire \top_ihp.oisc.regs[62][4] ;
 wire \top_ihp.oisc.regs[62][5] ;
 wire \top_ihp.oisc.regs[62][6] ;
 wire \top_ihp.oisc.regs[62][7] ;
 wire \top_ihp.oisc.regs[62][8] ;
 wire \top_ihp.oisc.regs[62][9] ;
 wire \top_ihp.oisc.regs[63][0] ;
 wire \top_ihp.oisc.regs[63][10] ;
 wire \top_ihp.oisc.regs[63][11] ;
 wire \top_ihp.oisc.regs[63][12] ;
 wire \top_ihp.oisc.regs[63][13] ;
 wire \top_ihp.oisc.regs[63][14] ;
 wire \top_ihp.oisc.regs[63][15] ;
 wire \top_ihp.oisc.regs[63][16] ;
 wire \top_ihp.oisc.regs[63][17] ;
 wire \top_ihp.oisc.regs[63][18] ;
 wire \top_ihp.oisc.regs[63][19] ;
 wire \top_ihp.oisc.regs[63][1] ;
 wire \top_ihp.oisc.regs[63][20] ;
 wire \top_ihp.oisc.regs[63][21] ;
 wire \top_ihp.oisc.regs[63][22] ;
 wire \top_ihp.oisc.regs[63][23] ;
 wire \top_ihp.oisc.regs[63][24] ;
 wire \top_ihp.oisc.regs[63][25] ;
 wire \top_ihp.oisc.regs[63][26] ;
 wire \top_ihp.oisc.regs[63][27] ;
 wire \top_ihp.oisc.regs[63][28] ;
 wire \top_ihp.oisc.regs[63][29] ;
 wire \top_ihp.oisc.regs[63][2] ;
 wire \top_ihp.oisc.regs[63][30] ;
 wire \top_ihp.oisc.regs[63][31] ;
 wire \top_ihp.oisc.regs[63][3] ;
 wire \top_ihp.oisc.regs[63][4] ;
 wire \top_ihp.oisc.regs[63][5] ;
 wire \top_ihp.oisc.regs[63][6] ;
 wire \top_ihp.oisc.regs[63][7] ;
 wire \top_ihp.oisc.regs[63][8] ;
 wire \top_ihp.oisc.regs[63][9] ;
 wire \top_ihp.oisc.regs[6][0] ;
 wire \top_ihp.oisc.regs[6][10] ;
 wire \top_ihp.oisc.regs[6][11] ;
 wire \top_ihp.oisc.regs[6][12] ;
 wire \top_ihp.oisc.regs[6][13] ;
 wire \top_ihp.oisc.regs[6][14] ;
 wire \top_ihp.oisc.regs[6][15] ;
 wire \top_ihp.oisc.regs[6][16] ;
 wire \top_ihp.oisc.regs[6][17] ;
 wire \top_ihp.oisc.regs[6][18] ;
 wire \top_ihp.oisc.regs[6][19] ;
 wire \top_ihp.oisc.regs[6][1] ;
 wire \top_ihp.oisc.regs[6][20] ;
 wire \top_ihp.oisc.regs[6][21] ;
 wire \top_ihp.oisc.regs[6][22] ;
 wire \top_ihp.oisc.regs[6][23] ;
 wire \top_ihp.oisc.regs[6][24] ;
 wire \top_ihp.oisc.regs[6][25] ;
 wire \top_ihp.oisc.regs[6][26] ;
 wire \top_ihp.oisc.regs[6][27] ;
 wire \top_ihp.oisc.regs[6][28] ;
 wire \top_ihp.oisc.regs[6][29] ;
 wire \top_ihp.oisc.regs[6][2] ;
 wire \top_ihp.oisc.regs[6][30] ;
 wire \top_ihp.oisc.regs[6][31] ;
 wire \top_ihp.oisc.regs[6][3] ;
 wire \top_ihp.oisc.regs[6][4] ;
 wire \top_ihp.oisc.regs[6][5] ;
 wire \top_ihp.oisc.regs[6][6] ;
 wire \top_ihp.oisc.regs[6][7] ;
 wire \top_ihp.oisc.regs[6][8] ;
 wire \top_ihp.oisc.regs[6][9] ;
 wire \top_ihp.oisc.regs[7][0] ;
 wire \top_ihp.oisc.regs[7][10] ;
 wire \top_ihp.oisc.regs[7][11] ;
 wire \top_ihp.oisc.regs[7][12] ;
 wire \top_ihp.oisc.regs[7][13] ;
 wire \top_ihp.oisc.regs[7][14] ;
 wire \top_ihp.oisc.regs[7][15] ;
 wire \top_ihp.oisc.regs[7][16] ;
 wire \top_ihp.oisc.regs[7][17] ;
 wire \top_ihp.oisc.regs[7][18] ;
 wire \top_ihp.oisc.regs[7][19] ;
 wire \top_ihp.oisc.regs[7][1] ;
 wire \top_ihp.oisc.regs[7][20] ;
 wire \top_ihp.oisc.regs[7][21] ;
 wire \top_ihp.oisc.regs[7][22] ;
 wire \top_ihp.oisc.regs[7][23] ;
 wire \top_ihp.oisc.regs[7][24] ;
 wire \top_ihp.oisc.regs[7][25] ;
 wire \top_ihp.oisc.regs[7][26] ;
 wire \top_ihp.oisc.regs[7][27] ;
 wire \top_ihp.oisc.regs[7][28] ;
 wire \top_ihp.oisc.regs[7][29] ;
 wire \top_ihp.oisc.regs[7][2] ;
 wire \top_ihp.oisc.regs[7][30] ;
 wire \top_ihp.oisc.regs[7][31] ;
 wire \top_ihp.oisc.regs[7][3] ;
 wire \top_ihp.oisc.regs[7][4] ;
 wire \top_ihp.oisc.regs[7][5] ;
 wire \top_ihp.oisc.regs[7][6] ;
 wire \top_ihp.oisc.regs[7][7] ;
 wire \top_ihp.oisc.regs[7][8] ;
 wire \top_ihp.oisc.regs[7][9] ;
 wire \top_ihp.oisc.regs[8][0] ;
 wire \top_ihp.oisc.regs[8][10] ;
 wire \top_ihp.oisc.regs[8][11] ;
 wire \top_ihp.oisc.regs[8][12] ;
 wire \top_ihp.oisc.regs[8][13] ;
 wire \top_ihp.oisc.regs[8][14] ;
 wire \top_ihp.oisc.regs[8][15] ;
 wire \top_ihp.oisc.regs[8][16] ;
 wire \top_ihp.oisc.regs[8][17] ;
 wire \top_ihp.oisc.regs[8][18] ;
 wire \top_ihp.oisc.regs[8][19] ;
 wire \top_ihp.oisc.regs[8][1] ;
 wire \top_ihp.oisc.regs[8][20] ;
 wire \top_ihp.oisc.regs[8][21] ;
 wire \top_ihp.oisc.regs[8][22] ;
 wire \top_ihp.oisc.regs[8][23] ;
 wire \top_ihp.oisc.regs[8][24] ;
 wire \top_ihp.oisc.regs[8][25] ;
 wire \top_ihp.oisc.regs[8][26] ;
 wire \top_ihp.oisc.regs[8][27] ;
 wire \top_ihp.oisc.regs[8][28] ;
 wire \top_ihp.oisc.regs[8][29] ;
 wire \top_ihp.oisc.regs[8][2] ;
 wire \top_ihp.oisc.regs[8][30] ;
 wire \top_ihp.oisc.regs[8][31] ;
 wire \top_ihp.oisc.regs[8][3] ;
 wire \top_ihp.oisc.regs[8][4] ;
 wire \top_ihp.oisc.regs[8][5] ;
 wire \top_ihp.oisc.regs[8][6] ;
 wire \top_ihp.oisc.regs[8][7] ;
 wire \top_ihp.oisc.regs[8][8] ;
 wire \top_ihp.oisc.regs[8][9] ;
 wire \top_ihp.oisc.regs[9][0] ;
 wire \top_ihp.oisc.regs[9][10] ;
 wire \top_ihp.oisc.regs[9][11] ;
 wire \top_ihp.oisc.regs[9][12] ;
 wire \top_ihp.oisc.regs[9][13] ;
 wire \top_ihp.oisc.regs[9][14] ;
 wire \top_ihp.oisc.regs[9][15] ;
 wire \top_ihp.oisc.regs[9][16] ;
 wire \top_ihp.oisc.regs[9][17] ;
 wire \top_ihp.oisc.regs[9][18] ;
 wire \top_ihp.oisc.regs[9][19] ;
 wire \top_ihp.oisc.regs[9][1] ;
 wire \top_ihp.oisc.regs[9][20] ;
 wire \top_ihp.oisc.regs[9][21] ;
 wire \top_ihp.oisc.regs[9][22] ;
 wire \top_ihp.oisc.regs[9][23] ;
 wire \top_ihp.oisc.regs[9][24] ;
 wire \top_ihp.oisc.regs[9][25] ;
 wire \top_ihp.oisc.regs[9][26] ;
 wire \top_ihp.oisc.regs[9][27] ;
 wire \top_ihp.oisc.regs[9][28] ;
 wire \top_ihp.oisc.regs[9][29] ;
 wire \top_ihp.oisc.regs[9][2] ;
 wire \top_ihp.oisc.regs[9][30] ;
 wire \top_ihp.oisc.regs[9][31] ;
 wire \top_ihp.oisc.regs[9][3] ;
 wire \top_ihp.oisc.regs[9][4] ;
 wire \top_ihp.oisc.regs[9][5] ;
 wire \top_ihp.oisc.regs[9][6] ;
 wire \top_ihp.oisc.regs[9][7] ;
 wire \top_ihp.oisc.regs[9][8] ;
 wire \top_ihp.oisc.regs[9][9] ;
 wire \top_ihp.oisc.state[0] ;
 wire \top_ihp.oisc.state[1] ;
 wire \top_ihp.oisc.state[2] ;
 wire \top_ihp.oisc.state[3] ;
 wire \top_ihp.oisc.state[4] ;
 wire \top_ihp.oisc.state[5] ;
 wire \top_ihp.oisc.state[6] ;
 wire \top_ihp.oisc.wb_adr_o[0] ;
 wire \top_ihp.oisc.wb_adr_o[1] ;
 wire \top_ihp.oisc.wb_dat_o[0] ;
 wire \top_ihp.oisc.wb_dat_o[10] ;
 wire \top_ihp.oisc.wb_dat_o[11] ;
 wire \top_ihp.oisc.wb_dat_o[12] ;
 wire \top_ihp.oisc.wb_dat_o[13] ;
 wire \top_ihp.oisc.wb_dat_o[14] ;
 wire \top_ihp.oisc.wb_dat_o[15] ;
 wire \top_ihp.oisc.wb_dat_o[16] ;
 wire \top_ihp.oisc.wb_dat_o[17] ;
 wire \top_ihp.oisc.wb_dat_o[18] ;
 wire \top_ihp.oisc.wb_dat_o[19] ;
 wire \top_ihp.oisc.wb_dat_o[1] ;
 wire \top_ihp.oisc.wb_dat_o[20] ;
 wire \top_ihp.oisc.wb_dat_o[21] ;
 wire \top_ihp.oisc.wb_dat_o[22] ;
 wire \top_ihp.oisc.wb_dat_o[23] ;
 wire \top_ihp.oisc.wb_dat_o[24] ;
 wire \top_ihp.oisc.wb_dat_o[25] ;
 wire \top_ihp.oisc.wb_dat_o[26] ;
 wire \top_ihp.oisc.wb_dat_o[27] ;
 wire \top_ihp.oisc.wb_dat_o[28] ;
 wire \top_ihp.oisc.wb_dat_o[29] ;
 wire \top_ihp.oisc.wb_dat_o[2] ;
 wire \top_ihp.oisc.wb_dat_o[30] ;
 wire \top_ihp.oisc.wb_dat_o[31] ;
 wire \top_ihp.oisc.wb_dat_o[3] ;
 wire \top_ihp.oisc.wb_dat_o[4] ;
 wire \top_ihp.oisc.wb_dat_o[5] ;
 wire \top_ihp.oisc.wb_dat_o[6] ;
 wire \top_ihp.oisc.wb_dat_o[7] ;
 wire \top_ihp.oisc.wb_dat_o[8] ;
 wire \top_ihp.oisc.wb_dat_o[9] ;
 wire \top_ihp.ram_clk_o ;
 wire \top_ihp.ram_cs_o ;
 wire \top_ihp.ram_data_o ;
 wire \top_ihp.rom_clk_o ;
 wire \top_ihp.rom_cs_o ;
 wire \top_ihp.rom_data_o ;
 wire \top_ihp.spi_clk_o ;
 wire \top_ihp.spi_cs_o_1 ;
 wire \top_ihp.spi_cs_o_2 ;
 wire \top_ihp.spi_cs_o_3 ;
 wire \top_ihp.spi_data_o ;
 wire \top_ihp.tx ;
 wire \top_ihp.wb_ack_coproc ;
 wire \top_ihp.wb_ack_gpio ;
 wire \top_ihp.wb_ack_spi ;
 wire \top_ihp.wb_ack_uart ;
 wire \top_ihp.wb_coproc.dat_o[0] ;
 wire \top_ihp.wb_coproc.dat_o[10] ;
 wire \top_ihp.wb_coproc.dat_o[11] ;
 wire \top_ihp.wb_coproc.dat_o[12] ;
 wire \top_ihp.wb_coproc.dat_o[13] ;
 wire \top_ihp.wb_coproc.dat_o[14] ;
 wire \top_ihp.wb_coproc.dat_o[15] ;
 wire \top_ihp.wb_coproc.dat_o[16] ;
 wire \top_ihp.wb_coproc.dat_o[17] ;
 wire \top_ihp.wb_coproc.dat_o[18] ;
 wire \top_ihp.wb_coproc.dat_o[19] ;
 wire \top_ihp.wb_coproc.dat_o[1] ;
 wire \top_ihp.wb_coproc.dat_o[20] ;
 wire \top_ihp.wb_coproc.dat_o[21] ;
 wire \top_ihp.wb_coproc.dat_o[22] ;
 wire \top_ihp.wb_coproc.dat_o[23] ;
 wire \top_ihp.wb_coproc.dat_o[24] ;
 wire \top_ihp.wb_coproc.dat_o[25] ;
 wire \top_ihp.wb_coproc.dat_o[26] ;
 wire \top_ihp.wb_coproc.dat_o[27] ;
 wire \top_ihp.wb_coproc.dat_o[28] ;
 wire \top_ihp.wb_coproc.dat_o[29] ;
 wire \top_ihp.wb_coproc.dat_o[2] ;
 wire \top_ihp.wb_coproc.dat_o[30] ;
 wire \top_ihp.wb_coproc.dat_o[31] ;
 wire \top_ihp.wb_coproc.dat_o[3] ;
 wire \top_ihp.wb_coproc.dat_o[4] ;
 wire \top_ihp.wb_coproc.dat_o[5] ;
 wire \top_ihp.wb_coproc.dat_o[6] ;
 wire \top_ihp.wb_coproc.dat_o[7] ;
 wire \top_ihp.wb_coproc.dat_o[8] ;
 wire \top_ihp.wb_coproc.dat_o[9] ;
 wire \top_ihp.wb_coproc.opa[0] ;
 wire \top_ihp.wb_coproc.opa[10] ;
 wire \top_ihp.wb_coproc.opa[11] ;
 wire \top_ihp.wb_coproc.opa[12] ;
 wire \top_ihp.wb_coproc.opa[13] ;
 wire \top_ihp.wb_coproc.opa[14] ;
 wire \top_ihp.wb_coproc.opa[15] ;
 wire \top_ihp.wb_coproc.opa[16] ;
 wire \top_ihp.wb_coproc.opa[17] ;
 wire \top_ihp.wb_coproc.opa[18] ;
 wire \top_ihp.wb_coproc.opa[19] ;
 wire \top_ihp.wb_coproc.opa[1] ;
 wire \top_ihp.wb_coproc.opa[20] ;
 wire \top_ihp.wb_coproc.opa[21] ;
 wire \top_ihp.wb_coproc.opa[22] ;
 wire \top_ihp.wb_coproc.opa[23] ;
 wire \top_ihp.wb_coproc.opa[24] ;
 wire \top_ihp.wb_coproc.opa[25] ;
 wire \top_ihp.wb_coproc.opa[26] ;
 wire \top_ihp.wb_coproc.opa[27] ;
 wire \top_ihp.wb_coproc.opa[28] ;
 wire \top_ihp.wb_coproc.opa[29] ;
 wire \top_ihp.wb_coproc.opa[2] ;
 wire \top_ihp.wb_coproc.opa[30] ;
 wire \top_ihp.wb_coproc.opa[31] ;
 wire \top_ihp.wb_coproc.opa[3] ;
 wire \top_ihp.wb_coproc.opa[4] ;
 wire \top_ihp.wb_coproc.opa[5] ;
 wire \top_ihp.wb_coproc.opa[6] ;
 wire \top_ihp.wb_coproc.opa[7] ;
 wire \top_ihp.wb_coproc.opa[8] ;
 wire \top_ihp.wb_coproc.opa[9] ;
 wire \top_ihp.wb_coproc.opb[0] ;
 wire \top_ihp.wb_coproc.opb[10] ;
 wire \top_ihp.wb_coproc.opb[11] ;
 wire \top_ihp.wb_coproc.opb[12] ;
 wire \top_ihp.wb_coproc.opb[13] ;
 wire \top_ihp.wb_coproc.opb[14] ;
 wire \top_ihp.wb_coproc.opb[15] ;
 wire \top_ihp.wb_coproc.opb[16] ;
 wire \top_ihp.wb_coproc.opb[17] ;
 wire \top_ihp.wb_coproc.opb[18] ;
 wire \top_ihp.wb_coproc.opb[19] ;
 wire \top_ihp.wb_coproc.opb[1] ;
 wire \top_ihp.wb_coproc.opb[20] ;
 wire \top_ihp.wb_coproc.opb[21] ;
 wire \top_ihp.wb_coproc.opb[22] ;
 wire \top_ihp.wb_coproc.opb[23] ;
 wire \top_ihp.wb_coproc.opb[24] ;
 wire \top_ihp.wb_coproc.opb[25] ;
 wire \top_ihp.wb_coproc.opb[26] ;
 wire \top_ihp.wb_coproc.opb[27] ;
 wire \top_ihp.wb_coproc.opb[28] ;
 wire \top_ihp.wb_coproc.opb[29] ;
 wire \top_ihp.wb_coproc.opb[2] ;
 wire \top_ihp.wb_coproc.opb[30] ;
 wire \top_ihp.wb_coproc.opb[31] ;
 wire \top_ihp.wb_coproc.opb[3] ;
 wire \top_ihp.wb_coproc.opb[4] ;
 wire \top_ihp.wb_coproc.opb[5] ;
 wire \top_ihp.wb_coproc.opb[6] ;
 wire \top_ihp.wb_coproc.opb[7] ;
 wire \top_ihp.wb_coproc.opb[8] ;
 wire \top_ihp.wb_coproc.opb[9] ;
 wire \top_ihp.wb_dati_gpio[0] ;
 wire \top_ihp.wb_dati_ram[0] ;
 wire \top_ihp.wb_dati_ram[10] ;
 wire \top_ihp.wb_dati_ram[11] ;
 wire \top_ihp.wb_dati_ram[12] ;
 wire \top_ihp.wb_dati_ram[13] ;
 wire \top_ihp.wb_dati_ram[14] ;
 wire \top_ihp.wb_dati_ram[15] ;
 wire \top_ihp.wb_dati_ram[16] ;
 wire \top_ihp.wb_dati_ram[17] ;
 wire \top_ihp.wb_dati_ram[18] ;
 wire \top_ihp.wb_dati_ram[19] ;
 wire \top_ihp.wb_dati_ram[1] ;
 wire \top_ihp.wb_dati_ram[20] ;
 wire \top_ihp.wb_dati_ram[21] ;
 wire \top_ihp.wb_dati_ram[22] ;
 wire \top_ihp.wb_dati_ram[23] ;
 wire \top_ihp.wb_dati_ram[24] ;
 wire \top_ihp.wb_dati_ram[25] ;
 wire \top_ihp.wb_dati_ram[26] ;
 wire \top_ihp.wb_dati_ram[27] ;
 wire \top_ihp.wb_dati_ram[28] ;
 wire \top_ihp.wb_dati_ram[29] ;
 wire \top_ihp.wb_dati_ram[2] ;
 wire \top_ihp.wb_dati_ram[30] ;
 wire \top_ihp.wb_dati_ram[31] ;
 wire \top_ihp.wb_dati_ram[3] ;
 wire \top_ihp.wb_dati_ram[4] ;
 wire \top_ihp.wb_dati_ram[5] ;
 wire \top_ihp.wb_dati_ram[6] ;
 wire \top_ihp.wb_dati_ram[7] ;
 wire \top_ihp.wb_dati_ram[8] ;
 wire \top_ihp.wb_dati_ram[9] ;
 wire \top_ihp.wb_dati_rom[0] ;
 wire \top_ihp.wb_dati_rom[10] ;
 wire \top_ihp.wb_dati_rom[11] ;
 wire \top_ihp.wb_dati_rom[12] ;
 wire \top_ihp.wb_dati_rom[13] ;
 wire \top_ihp.wb_dati_rom[14] ;
 wire \top_ihp.wb_dati_rom[15] ;
 wire \top_ihp.wb_dati_rom[16] ;
 wire \top_ihp.wb_dati_rom[17] ;
 wire \top_ihp.wb_dati_rom[18] ;
 wire \top_ihp.wb_dati_rom[19] ;
 wire \top_ihp.wb_dati_rom[1] ;
 wire \top_ihp.wb_dati_rom[20] ;
 wire \top_ihp.wb_dati_rom[21] ;
 wire \top_ihp.wb_dati_rom[22] ;
 wire \top_ihp.wb_dati_rom[23] ;
 wire \top_ihp.wb_dati_rom[24] ;
 wire \top_ihp.wb_dati_rom[25] ;
 wire \top_ihp.wb_dati_rom[26] ;
 wire \top_ihp.wb_dati_rom[27] ;
 wire \top_ihp.wb_dati_rom[28] ;
 wire \top_ihp.wb_dati_rom[29] ;
 wire \top_ihp.wb_dati_rom[2] ;
 wire \top_ihp.wb_dati_rom[30] ;
 wire \top_ihp.wb_dati_rom[31] ;
 wire \top_ihp.wb_dati_rom[3] ;
 wire \top_ihp.wb_dati_rom[4] ;
 wire \top_ihp.wb_dati_rom[5] ;
 wire \top_ihp.wb_dati_rom[6] ;
 wire \top_ihp.wb_dati_rom[7] ;
 wire \top_ihp.wb_dati_rom[8] ;
 wire \top_ihp.wb_dati_rom[9] ;
 wire \top_ihp.wb_dati_spi[0] ;
 wire \top_ihp.wb_dati_spi[10] ;
 wire \top_ihp.wb_dati_spi[11] ;
 wire \top_ihp.wb_dati_spi[12] ;
 wire \top_ihp.wb_dati_spi[13] ;
 wire \top_ihp.wb_dati_spi[14] ;
 wire \top_ihp.wb_dati_spi[15] ;
 wire \top_ihp.wb_dati_spi[16] ;
 wire \top_ihp.wb_dati_spi[17] ;
 wire \top_ihp.wb_dati_spi[18] ;
 wire \top_ihp.wb_dati_spi[19] ;
 wire \top_ihp.wb_dati_spi[1] ;
 wire \top_ihp.wb_dati_spi[20] ;
 wire \top_ihp.wb_dati_spi[21] ;
 wire \top_ihp.wb_dati_spi[22] ;
 wire \top_ihp.wb_dati_spi[23] ;
 wire \top_ihp.wb_dati_spi[24] ;
 wire \top_ihp.wb_dati_spi[25] ;
 wire \top_ihp.wb_dati_spi[26] ;
 wire \top_ihp.wb_dati_spi[27] ;
 wire \top_ihp.wb_dati_spi[28] ;
 wire \top_ihp.wb_dati_spi[29] ;
 wire \top_ihp.wb_dati_spi[2] ;
 wire \top_ihp.wb_dati_spi[30] ;
 wire \top_ihp.wb_dati_spi[31] ;
 wire \top_ihp.wb_dati_spi[3] ;
 wire \top_ihp.wb_dati_spi[4] ;
 wire \top_ihp.wb_dati_spi[5] ;
 wire \top_ihp.wb_dati_spi[6] ;
 wire \top_ihp.wb_dati_spi[7] ;
 wire \top_ihp.wb_dati_spi[8] ;
 wire \top_ihp.wb_dati_spi[9] ;
 wire \top_ihp.wb_dati_uart[0] ;
 wire \top_ihp.wb_dati_uart[1] ;
 wire \top_ihp.wb_dati_uart[2] ;
 wire \top_ihp.wb_dati_uart[3] ;
 wire \top_ihp.wb_dati_uart[4] ;
 wire \top_ihp.wb_dati_uart[5] ;
 wire \top_ihp.wb_dati_uart[6] ;
 wire \top_ihp.wb_dati_uart[7] ;
 wire \top_ihp.wb_emem.bit_counter[0] ;
 wire \top_ihp.wb_emem.bit_counter[1] ;
 wire \top_ihp.wb_emem.bit_counter[2] ;
 wire \top_ihp.wb_emem.bit_counter[3] ;
 wire \top_ihp.wb_emem.bit_counter[4] ;
 wire \top_ihp.wb_emem.bit_counter[5] ;
 wire \top_ihp.wb_emem.bit_counter[6] ;
 wire \top_ihp.wb_emem.bit_counter[7] ;
 wire \top_ihp.wb_emem.cmd[32] ;
 wire \top_ihp.wb_emem.cmd[33] ;
 wire \top_ihp.wb_emem.cmd[34] ;
 wire \top_ihp.wb_emem.cmd[35] ;
 wire \top_ihp.wb_emem.cmd[36] ;
 wire \top_ihp.wb_emem.cmd[37] ;
 wire \top_ihp.wb_emem.cmd[38] ;
 wire \top_ihp.wb_emem.cmd[39] ;
 wire \top_ihp.wb_emem.cmd[40] ;
 wire \top_ihp.wb_emem.cmd[41] ;
 wire \top_ihp.wb_emem.cmd[42] ;
 wire \top_ihp.wb_emem.cmd[43] ;
 wire \top_ihp.wb_emem.cmd[44] ;
 wire \top_ihp.wb_emem.cmd[45] ;
 wire \top_ihp.wb_emem.cmd[46] ;
 wire \top_ihp.wb_emem.cmd[47] ;
 wire \top_ihp.wb_emem.cmd[48] ;
 wire \top_ihp.wb_emem.cmd[49] ;
 wire \top_ihp.wb_emem.cmd[50] ;
 wire \top_ihp.wb_emem.cmd[51] ;
 wire \top_ihp.wb_emem.cmd[52] ;
 wire \top_ihp.wb_emem.cmd[53] ;
 wire \top_ihp.wb_emem.cmd[54] ;
 wire \top_ihp.wb_emem.cmd[55] ;
 wire \top_ihp.wb_emem.cmd[56] ;
 wire \top_ihp.wb_emem.cmd[57] ;
 wire \top_ihp.wb_emem.cmd[58] ;
 wire \top_ihp.wb_emem.cmd[59] ;
 wire \top_ihp.wb_emem.cmd[60] ;
 wire \top_ihp.wb_emem.cmd[61] ;
 wire \top_ihp.wb_emem.cmd[62] ;
 wire \top_ihp.wb_emem.cmd[63] ;
 wire \top_ihp.wb_emem.last_bit ;
 wire \top_ihp.wb_emem.last_wait ;
 wire \top_ihp.wb_emem.nbits[3] ;
 wire \top_ihp.wb_emem.nbits[4] ;
 wire \top_ihp.wb_emem.nbits[5] ;
 wire \top_ihp.wb_emem.nbits[6] ;
 wire \top_ihp.wb_emem.state[0] ;
 wire \top_ihp.wb_emem.state[1] ;
 wire \top_ihp.wb_emem.state[2] ;
 wire \top_ihp.wb_emem.state[3] ;
 wire \top_ihp.wb_emem.wait_counter[0] ;
 wire \top_ihp.wb_emem.wait_counter[1] ;
 wire \top_ihp.wb_emem.wait_counter[2] ;
 wire \top_ihp.wb_emem.wait_counter[3] ;
 wire \top_ihp.wb_emem.wait_counter[4] ;
 wire \top_ihp.wb_emem.wait_counter[5] ;
 wire \top_ihp.wb_emem.wait_counter[6] ;
 wire \top_ihp.wb_emem.wait_counter[7] ;
 wire \top_ihp.wb_imem.bits_left[0] ;
 wire \top_ihp.wb_imem.bits_left[1] ;
 wire \top_ihp.wb_imem.bits_left[2] ;
 wire \top_ihp.wb_imem.bits_left[3] ;
 wire \top_ihp.wb_imem.bits_left[4] ;
 wire \top_ihp.wb_imem.bits_left[5] ;
 wire \top_ihp.wb_imem.state[0] ;
 wire \top_ihp.wb_imem.state[1] ;
 wire \top_ihp.wb_imem.state[2] ;
 wire \top_ihp.wb_spi.bits_left[0] ;
 wire \top_ihp.wb_spi.bits_left[1] ;
 wire \top_ihp.wb_spi.bits_left[2] ;
 wire \top_ihp.wb_spi.bits_left[3] ;
 wire \top_ihp.wb_spi.bits_left[4] ;
 wire \top_ihp.wb_spi.bits_left[5] ;
 wire \top_ihp.wb_spi.spi_clk_cnt[0] ;
 wire \top_ihp.wb_spi.state ;
 wire \top_ihp.wb_uart.rx_ready ;
 wire \top_ihp.wb_uart.state[0] ;
 wire \top_ihp.wb_uart.state[1] ;
 wire \top_ihp.wb_uart.tx_ready ;
 wire \top_ihp.wb_uart.uart_rx.bit_cnt[0] ;
 wire \top_ihp.wb_uart.uart_rx.bit_cnt[1] ;
 wire \top_ihp.wb_uart.uart_rx.bit_cnt[2] ;
 wire \top_ihp.wb_uart.uart_rx.bit_cnt[3] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[0] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[10] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[11] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[12] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[13] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[14] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[15] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[16] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[17] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[18] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[19] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[1] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[20] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[21] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[22] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[23] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[24] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[25] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[26] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[27] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[28] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[29] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[2] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[30] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[31] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[3] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[4] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[5] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[6] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[7] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[8] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[9] ;
 wire \top_ihp.wb_uart.uart_rx.next_state[0] ;
 wire \top_ihp.wb_uart.uart_rx.next_state[1] ;
 wire \top_ihp.wb_uart.uart_rx.next_state[2] ;
 wire \top_ihp.wb_uart.uart_rx.state[0] ;
 wire \top_ihp.wb_uart.uart_rx.state[1] ;
 wire \top_ihp.wb_uart.uart_rx.state[2] ;
 wire \top_ihp.wb_uart.uart_tx.bit_cnt[0] ;
 wire \top_ihp.wb_uart.uart_tx.bit_cnt[1] ;
 wire \top_ihp.wb_uart.uart_tx.bit_cnt[2] ;
 wire \top_ihp.wb_uart.uart_tx.bit_cnt[3] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[0] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[10] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[11] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[12] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[13] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[14] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[15] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[16] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[17] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[18] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[19] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[1] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[20] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[21] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[22] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[23] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[24] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[25] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[26] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[27] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[28] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[29] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[2] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[30] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[31] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[3] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[4] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[5] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[6] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[7] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[8] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[9] ;
 wire \top_ihp.wb_uart.uart_tx.next_state[0] ;
 wire \top_ihp.wb_uart.uart_tx.next_state[1] ;
 wire \top_ihp.wb_uart.uart_tx.state[0] ;
 wire \top_ihp.wb_uart.uart_tx.state[1] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[0] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[1] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[2] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[3] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[4] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[5] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[6] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_314_clk;
 wire clknet_leaf_315_clk;
 wire clknet_leaf_316_clk;
 wire clknet_leaf_317_clk;
 wire clknet_leaf_318_clk;
 wire clknet_leaf_319_clk;
 wire clknet_leaf_320_clk;
 wire clknet_leaf_321_clk;
 wire clknet_leaf_322_clk;
 wire clknet_leaf_323_clk;
 wire clknet_leaf_324_clk;
 wire clknet_leaf_325_clk;
 wire clknet_leaf_326_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;

 sg13g2_buf_2 _13606_ (.A(\top_ihp.oisc.decoder.decoded[10] ),
    .X(_07958_));
 sg13g2_buf_2 _13607_ (.A(\top_ihp.oisc.state[5] ),
    .X(_07959_));
 sg13g2_buf_1 _13608_ (.A(_07959_),
    .X(_07960_));
 sg13g2_inv_2 _13609_ (.Y(_07961_),
    .A(net1049));
 sg13g2_buf_2 _13610_ (.A(\top_ihp.oisc.micro_op[1] ),
    .X(_07962_));
 sg13g2_buf_2 _13611_ (.A(\top_ihp.oisc.micro_op[0] ),
    .X(_07963_));
 sg13g2_buf_2 _13612_ (.A(\top_ihp.oisc.micro_op[3] ),
    .X(_07964_));
 sg13g2_and4_1 _13613_ (.A(_07962_),
    .B(_07963_),
    .C(_07964_),
    .D(\top_ihp.oisc.micro_state[2] ),
    .X(_07965_));
 sg13g2_buf_1 _13614_ (.A(_07965_),
    .X(_07966_));
 sg13g2_buf_2 _13615_ (.A(\top_ihp.oisc.micro_op[2] ),
    .X(_07967_));
 sg13g2_buf_2 _13616_ (.A(\top_ihp.oisc.micro_op[4] ),
    .X(_07968_));
 sg13g2_buf_1 _13617_ (.A(\top_ihp.oisc.micro_op[5] ),
    .X(_07969_));
 sg13g2_and3_1 _13618_ (.X(_07970_),
    .A(_07967_),
    .B(_07968_),
    .C(_07969_));
 sg13g2_buf_1 _13619_ (.A(_07970_),
    .X(_07971_));
 sg13g2_nand2_1 _13620_ (.Y(_07972_),
    .A(_07966_),
    .B(_07971_));
 sg13g2_buf_2 _13621_ (.A(_07972_),
    .X(_07973_));
 sg13g2_nor2_2 _13622_ (.A(_07961_),
    .B(_07973_),
    .Y(_07974_));
 sg13g2_and2_1 _13623_ (.A(_07958_),
    .B(_07974_),
    .X(_07975_));
 sg13g2_buf_1 _13624_ (.A(_07975_),
    .X(_07976_));
 sg13g2_buf_1 _13625_ (.A(_07976_),
    .X(_07977_));
 sg13g2_buf_1 _13626_ (.A(net857),
    .X(_07978_));
 sg13g2_buf_1 _13627_ (.A(\top_ihp.oisc.op_a[26] ),
    .X(_07979_));
 sg13g2_buf_2 _13628_ (.A(_07979_),
    .X(_07980_));
 sg13g2_inv_1 _13629_ (.Y(_07981_),
    .A(net1048));
 sg13g2_buf_1 _13630_ (.A(_07981_),
    .X(_07982_));
 sg13g2_buf_1 _13631_ (.A(\top_ihp.oisc.state[1] ),
    .X(_07983_));
 sg13g2_buf_1 _13632_ (.A(_07983_),
    .X(_07984_));
 sg13g2_buf_1 _13633_ (.A(net1047),
    .X(_07985_));
 sg13g2_buf_1 _13634_ (.A(net1019),
    .X(_07986_));
 sg13g2_buf_1 _13635_ (.A(_07986_),
    .X(_07987_));
 sg13g2_buf_2 _13636_ (.A(\top_ihp.oisc.op_b[26] ),
    .X(_07988_));
 sg13g2_inv_1 _13637_ (.Y(_07989_),
    .A(_07988_));
 sg13g2_buf_2 _13638_ (.A(\top_ihp.oisc.op_a[20] ),
    .X(_07990_));
 sg13g2_inv_1 _13639_ (.Y(_07991_),
    .A(\top_ihp.oisc.op_b[20] ));
 sg13g2_nor2_1 _13640_ (.A(_07990_),
    .B(_07991_),
    .Y(_07992_));
 sg13g2_buf_1 _13641_ (.A(_07992_),
    .X(_07993_));
 sg13g2_buf_1 _13642_ (.A(\top_ihp.oisc.op_b[19] ),
    .X(_07994_));
 sg13g2_buf_1 _13643_ (.A(\top_ihp.oisc.op_a[18] ),
    .X(_07995_));
 sg13g2_buf_2 _13644_ (.A(\top_ihp.oisc.op_b[18] ),
    .X(_07996_));
 sg13g2_nor2b_1 _13645_ (.A(net1070),
    .B_N(_07996_),
    .Y(_07997_));
 sg13g2_nand2_1 _13646_ (.Y(_07998_),
    .A(net1071),
    .B(_07997_));
 sg13g2_buf_2 _13647_ (.A(\top_ihp.oisc.op_a[19] ),
    .X(_07999_));
 sg13g2_inv_1 _13648_ (.Y(_08000_),
    .A(_07999_));
 sg13g2_o21ai_1 _13649_ (.B1(_08000_),
    .Y(_08001_),
    .A1(\top_ihp.oisc.op_b[19] ),
    .A2(_07997_));
 sg13g2_nor2b_1 _13650_ (.A(\top_ihp.oisc.op_b[20] ),
    .B_N(_07990_),
    .Y(_08002_));
 sg13g2_buf_1 _13651_ (.A(_08002_),
    .X(_08003_));
 sg13g2_a21oi_1 _13652_ (.A1(_07998_),
    .A2(_08001_),
    .Y(_08004_),
    .B1(_08003_));
 sg13g2_buf_8 _13653_ (.A(\top_ihp.oisc.op_a[17] ),
    .X(_08005_));
 sg13g2_buf_8 _13654_ (.A(\top_ihp.oisc.op_b[17] ),
    .X(_08006_));
 sg13g2_nor2b_1 _13655_ (.A(_08005_),
    .B_N(_08006_),
    .Y(_08007_));
 sg13g2_nand2b_1 _13656_ (.Y(_08008_),
    .B(_08005_),
    .A_N(_08006_));
 sg13g2_buf_8 _13657_ (.A(\top_ihp.oisc.op_b[15] ),
    .X(_08009_));
 sg13g2_buf_8 _13658_ (.A(\top_ihp.oisc.op_a[16] ),
    .X(_08010_));
 sg13g2_nor2b_1 _13659_ (.A(_08009_),
    .B_N(net1069),
    .Y(_08011_));
 sg13g2_buf_8 _13660_ (.A(\top_ihp.oisc.op_a[15] ),
    .X(_08012_));
 sg13g2_and2_1 _13661_ (.A(net1069),
    .B(net1068),
    .X(_08013_));
 sg13g2_buf_8 _13662_ (.A(\top_ihp.oisc.op_a[14] ),
    .X(_08014_));
 sg13g2_nand2b_1 _13663_ (.Y(_08015_),
    .B(\top_ihp.oisc.op_b[14] ),
    .A_N(net1067));
 sg13g2_buf_2 _13664_ (.A(_08015_),
    .X(_08016_));
 sg13g2_o21ai_1 _13665_ (.B1(_08016_),
    .Y(_08017_),
    .A1(_08011_),
    .A2(_08013_));
 sg13g2_nor2b_1 _13666_ (.A(_08009_),
    .B_N(net1068),
    .Y(_08018_));
 sg13g2_buf_1 _13667_ (.A(\top_ihp.oisc.op_b[16] ),
    .X(_08019_));
 sg13g2_nor2_1 _13668_ (.A(net1066),
    .B(_08009_),
    .Y(_08020_));
 sg13g2_a22oi_1 _13669_ (.Y(_08021_),
    .B1(_08020_),
    .B2(_08016_),
    .A2(_08018_),
    .A1(net1069));
 sg13g2_inv_1 _13670_ (.Y(_08022_),
    .A(net1066));
 sg13g2_nor2b_1 _13671_ (.A(_08019_),
    .B_N(net1068),
    .Y(_08023_));
 sg13g2_nor2b_1 _13672_ (.A(net1066),
    .B_N(net1069),
    .Y(_08024_));
 sg13g2_a221oi_1 _13673_ (.B2(_08016_),
    .C1(_08024_),
    .B1(_08023_),
    .A1(_08022_),
    .Y(_08025_),
    .A2(_08018_));
 sg13g2_and4_1 _13674_ (.A(_08008_),
    .B(_08017_),
    .C(_08021_),
    .D(_08025_),
    .X(_08026_));
 sg13g2_or4_1 _13675_ (.A(_07993_),
    .B(_08004_),
    .C(_08007_),
    .D(_08026_),
    .X(_08027_));
 sg13g2_buf_8 _13676_ (.A(\top_ihp.oisc.op_b[11] ),
    .X(_08028_));
 sg13g2_buf_1 _13677_ (.A(\top_ihp.oisc.op_a[10] ),
    .X(_08029_));
 sg13g2_buf_2 _13678_ (.A(\top_ihp.oisc.op_b[10] ),
    .X(_08030_));
 sg13g2_nor2b_1 _13679_ (.A(net1065),
    .B_N(_08030_),
    .Y(_08031_));
 sg13g2_buf_8 _13680_ (.A(\top_ihp.oisc.op_b[12] ),
    .X(_08032_));
 sg13g2_buf_8 _13681_ (.A(\top_ihp.oisc.op_a[12] ),
    .X(_08033_));
 sg13g2_nand2b_1 _13682_ (.Y(_08034_),
    .B(net1064),
    .A_N(_08032_));
 sg13g2_o21ai_1 _13683_ (.B1(_08034_),
    .Y(_08035_),
    .A1(_08028_),
    .A2(_08031_));
 sg13g2_buf_8 _13684_ (.A(\top_ihp.oisc.op_a[11] ),
    .X(_08036_));
 sg13g2_nand3b_1 _13685_ (.B(_08030_),
    .C(_08028_),
    .Y(_08037_),
    .A_N(net1065));
 sg13g2_buf_1 _13686_ (.A(_08037_),
    .X(_08038_));
 sg13g2_nand2_1 _13687_ (.Y(_08039_),
    .A(net1063),
    .B(_08038_));
 sg13g2_nand2b_1 _13688_ (.Y(_08040_),
    .B(_08039_),
    .A_N(_08035_));
 sg13g2_xnor2_1 _13689_ (.Y(_08041_),
    .A(net1063),
    .B(_08028_));
 sg13g2_buf_2 _13690_ (.A(_08041_),
    .X(_08042_));
 sg13g2_xnor2_1 _13691_ (.Y(_08043_),
    .A(net1065),
    .B(_08030_));
 sg13g2_xnor2_1 _13692_ (.Y(_08044_),
    .A(net1064),
    .B(_08032_));
 sg13g2_buf_2 _13693_ (.A(_08044_),
    .X(_08045_));
 sg13g2_buf_8 _13694_ (.A(\top_ihp.oisc.op_a[13] ),
    .X(_08046_));
 sg13g2_buf_1 _13695_ (.A(\top_ihp.oisc.op_b[13] ),
    .X(_08047_));
 sg13g2_xnor2_1 _13696_ (.Y(_08048_),
    .A(_08046_),
    .B(_08047_));
 sg13g2_nand4_1 _13697_ (.B(_08043_),
    .C(_08045_),
    .A(_08042_),
    .Y(_08049_),
    .D(_08048_));
 sg13g2_buf_1 _13698_ (.A(_08047_),
    .X(_08050_));
 sg13g2_nor2b_1 _13699_ (.A(net1064),
    .B_N(_08032_),
    .Y(_08051_));
 sg13g2_nor2_1 _13700_ (.A(net1046),
    .B(_08051_),
    .Y(_08052_));
 sg13g2_and2_1 _13701_ (.A(_08049_),
    .B(_08052_),
    .X(_08053_));
 sg13g2_nand2b_1 _13702_ (.Y(_08054_),
    .B(_08032_),
    .A_N(net1064));
 sg13g2_and3_1 _13703_ (.X(_08055_),
    .A(net1063),
    .B(_08038_),
    .C(_08054_));
 sg13g2_nor3_1 _13704_ (.A(_08028_),
    .B(_08031_),
    .C(_08051_),
    .Y(_08056_));
 sg13g2_nand2_1 _13705_ (.Y(_08057_),
    .A(net1046),
    .B(_08034_));
 sg13g2_or3_1 _13706_ (.A(_08055_),
    .B(_08056_),
    .C(_08057_),
    .X(_08058_));
 sg13g2_and2_1 _13707_ (.A(_08046_),
    .B(_08049_),
    .X(_08059_));
 sg13g2_xnor2_1 _13708_ (.Y(_08060_),
    .A(net1068),
    .B(_08009_));
 sg13g2_nand2b_1 _13709_ (.Y(_08061_),
    .B(_08014_),
    .A_N(\top_ihp.oisc.op_b[14] ));
 sg13g2_nand3_1 _13710_ (.B(_08060_),
    .C(_08061_),
    .A(_08016_),
    .Y(_08062_));
 sg13g2_buf_2 _13711_ (.A(_08062_),
    .X(_08063_));
 sg13g2_xor2_1 _13712_ (.B(_08006_),
    .A(_08005_),
    .X(_08064_));
 sg13g2_nor2b_1 _13713_ (.A(net1069),
    .B_N(net1066),
    .Y(_08065_));
 sg13g2_buf_1 _13714_ (.A(_08065_),
    .X(_08066_));
 sg13g2_nor3_1 _13715_ (.A(_08024_),
    .B(_08064_),
    .C(_08066_),
    .Y(_08067_));
 sg13g2_nand2b_1 _13716_ (.Y(_08068_),
    .B(_08067_),
    .A_N(_08063_));
 sg13g2_a221oi_1 _13717_ (.B2(_08059_),
    .C1(_08068_),
    .B1(_08058_),
    .A1(_08040_),
    .Y(_08069_),
    .A2(_08053_));
 sg13g2_nand2b_1 _13718_ (.Y(_08070_),
    .B(net1070),
    .A_N(_07996_));
 sg13g2_buf_1 _13719_ (.A(_08070_),
    .X(_08071_));
 sg13g2_nor2_1 _13720_ (.A(net1071),
    .B(_08071_),
    .Y(_08072_));
 sg13g2_a21oi_1 _13721_ (.A1(net1071),
    .A2(_08071_),
    .Y(_08073_),
    .B1(_08000_));
 sg13g2_nor3_1 _13722_ (.A(_08003_),
    .B(_08072_),
    .C(_08073_),
    .Y(_08074_));
 sg13g2_or2_1 _13723_ (.X(_08075_),
    .B(_08074_),
    .A(_07993_));
 sg13g2_o21ai_1 _13724_ (.B1(_08075_),
    .Y(_08076_),
    .A1(_08027_),
    .A2(_08069_));
 sg13g2_buf_1 _13725_ (.A(_08076_),
    .X(_08077_));
 sg13g2_buf_2 _13726_ (.A(\top_ihp.oisc.op_a[1] ),
    .X(_08078_));
 sg13g2_inv_2 _13727_ (.Y(_08079_),
    .A(_08078_));
 sg13g2_buf_1 _13728_ (.A(\top_ihp.oisc.op_b[1] ),
    .X(_08080_));
 sg13g2_buf_1 _13729_ (.A(\top_ihp.oisc.op_b[0] ),
    .X(_08081_));
 sg13g2_buf_2 _13730_ (.A(\top_ihp.oisc.op_a[0] ),
    .X(_08082_));
 sg13g2_nand2b_1 _13731_ (.Y(_08083_),
    .B(_08082_),
    .A_N(_08081_));
 sg13g2_buf_1 _13732_ (.A(_08083_),
    .X(_08084_));
 sg13g2_o21ai_1 _13733_ (.B1(_08084_),
    .Y(_08085_),
    .A1(_08079_),
    .A2(_08080_));
 sg13g2_buf_2 _13734_ (.A(\top_ihp.oisc.op_a[3] ),
    .X(_08086_));
 sg13g2_buf_2 _13735_ (.A(\top_ihp.oisc.op_b[3] ),
    .X(_08087_));
 sg13g2_nor2b_1 _13736_ (.A(_08086_),
    .B_N(_08087_),
    .Y(_08088_));
 sg13g2_nor2b_1 _13737_ (.A(_08078_),
    .B_N(_08080_),
    .Y(_08089_));
 sg13g2_buf_2 _13738_ (.A(\top_ihp.oisc.op_a[2] ),
    .X(_08090_));
 sg13g2_buf_2 _13739_ (.A(\top_ihp.oisc.op_b[2] ),
    .X(_08091_));
 sg13g2_nor2b_1 _13740_ (.A(_08090_),
    .B_N(_08091_),
    .Y(_08092_));
 sg13g2_nor3_1 _13741_ (.A(_08088_),
    .B(_08089_),
    .C(_08092_),
    .Y(_08093_));
 sg13g2_nand2b_1 _13742_ (.Y(_08094_),
    .B(_08090_),
    .A_N(_08091_));
 sg13g2_buf_1 _13743_ (.A(_08094_),
    .X(_08095_));
 sg13g2_nand2_1 _13744_ (.Y(_08096_),
    .A(_08087_),
    .B(_08095_));
 sg13g2_nor2_1 _13745_ (.A(_08087_),
    .B(_08095_),
    .Y(_08097_));
 sg13g2_a221oi_1 _13746_ (.B2(_08086_),
    .C1(_08097_),
    .B1(_08096_),
    .A1(_08085_),
    .Y(_08098_),
    .A2(_08093_));
 sg13g2_buf_1 _13747_ (.A(_08098_),
    .X(_08099_));
 sg13g2_buf_2 _13748_ (.A(\top_ihp.oisc.op_a[8] ),
    .X(_08100_));
 sg13g2_buf_2 _13749_ (.A(\top_ihp.oisc.op_b[8] ),
    .X(_08101_));
 sg13g2_xnor2_1 _13750_ (.Y(_08102_),
    .A(_08100_),
    .B(_08101_));
 sg13g2_buf_8 _13751_ (.A(\top_ihp.oisc.op_a[9] ),
    .X(_08103_));
 sg13g2_nand2b_1 _13752_ (.Y(_08104_),
    .B(_08103_),
    .A_N(\top_ihp.oisc.op_b[9] ));
 sg13g2_buf_2 _13753_ (.A(_08104_),
    .X(_08105_));
 sg13g2_nand2b_1 _13754_ (.Y(_08106_),
    .B(\top_ihp.oisc.op_b[9] ),
    .A_N(_08103_));
 sg13g2_buf_2 _13755_ (.A(_08106_),
    .X(_08107_));
 sg13g2_nand3_1 _13756_ (.B(_08105_),
    .C(_08107_),
    .A(_08102_),
    .Y(_08108_));
 sg13g2_buf_2 _13757_ (.A(\top_ihp.oisc.op_a[4] ),
    .X(_08109_));
 sg13g2_buf_2 _13758_ (.A(\top_ihp.oisc.op_b[4] ),
    .X(_08110_));
 sg13g2_nor2b_1 _13759_ (.A(_08109_),
    .B_N(_08110_),
    .Y(_08111_));
 sg13g2_buf_2 _13760_ (.A(_08111_),
    .X(_08112_));
 sg13g2_nand2b_1 _13761_ (.Y(_08113_),
    .B(_08109_),
    .A_N(_08110_));
 sg13g2_nand2b_1 _13762_ (.Y(_08114_),
    .B(_08113_),
    .A_N(_08112_));
 sg13g2_buf_1 _13763_ (.A(\top_ihp.oisc.op_b[7] ),
    .X(_08115_));
 sg13g2_buf_2 _13764_ (.A(\top_ihp.oisc.op_a[7] ),
    .X(_08116_));
 sg13g2_nor2b_1 _13765_ (.A(_08115_),
    .B_N(_08116_),
    .Y(_08117_));
 sg13g2_nor2b_1 _13766_ (.A(_08116_),
    .B_N(_08115_),
    .Y(_08118_));
 sg13g2_buf_2 _13767_ (.A(_08118_),
    .X(_08119_));
 sg13g2_or2_1 _13768_ (.X(_08120_),
    .B(_08119_),
    .A(_08117_));
 sg13g2_buf_1 _13769_ (.A(\top_ihp.oisc.op_a[6] ),
    .X(_08121_));
 sg13g2_buf_8 _13770_ (.A(_08121_),
    .X(_08122_));
 sg13g2_buf_1 _13771_ (.A(\top_ihp.oisc.op_b[6] ),
    .X(_08123_));
 sg13g2_nand2b_1 _13772_ (.Y(_08124_),
    .B(net1062),
    .A_N(net1045));
 sg13g2_nand2b_1 _13773_ (.Y(_08125_),
    .B(_08121_),
    .A_N(net1062));
 sg13g2_buf_2 _13774_ (.A(\top_ihp.oisc.op_a[5] ),
    .X(_08126_));
 sg13g2_buf_2 _13775_ (.A(\top_ihp.oisc.op_b[5] ),
    .X(_08127_));
 sg13g2_nand2b_1 _13776_ (.Y(_08128_),
    .B(_08127_),
    .A_N(_08126_));
 sg13g2_buf_1 _13777_ (.A(_08128_),
    .X(_08129_));
 sg13g2_nand2b_1 _13778_ (.Y(_08130_),
    .B(_08126_),
    .A_N(_08127_));
 sg13g2_nand4_1 _13779_ (.B(_08125_),
    .C(_08129_),
    .A(_08124_),
    .Y(_08131_),
    .D(_08130_));
 sg13g2_nor4_1 _13780_ (.A(_08108_),
    .B(_08114_),
    .C(_08120_),
    .D(_08131_),
    .Y(_08132_));
 sg13g2_inv_1 _13781_ (.Y(_08133_),
    .A(_08100_));
 sg13g2_a21oi_1 _13782_ (.A1(_08101_),
    .A2(_08119_),
    .Y(_08134_),
    .B1(_08133_));
 sg13g2_nor2_1 _13783_ (.A(_08101_),
    .B(_08119_),
    .Y(_08135_));
 sg13g2_o21ai_1 _13784_ (.B1(_08107_),
    .Y(_08136_),
    .A1(_08134_),
    .A2(_08135_));
 sg13g2_nor2b_1 _13785_ (.A(net1045),
    .B_N(net1062),
    .Y(_08137_));
 sg13g2_nor3_1 _13786_ (.A(_08127_),
    .B(_08137_),
    .C(_08112_),
    .Y(_08138_));
 sg13g2_inv_1 _13787_ (.Y(_08139_),
    .A(net1045));
 sg13g2_inv_1 _13788_ (.Y(_08140_),
    .A(_08126_));
 sg13g2_a221oi_1 _13789_ (.B2(_08112_),
    .C1(_08140_),
    .B1(_08127_),
    .A1(_08139_),
    .Y(_08141_),
    .A2(net1062));
 sg13g2_nand4_1 _13790_ (.B(_08105_),
    .C(_08107_),
    .A(_08102_),
    .Y(_08142_),
    .D(_08125_));
 sg13g2_nor4_1 _13791_ (.A(_08117_),
    .B(_08138_),
    .C(_08141_),
    .D(_08142_),
    .Y(_08143_));
 sg13g2_a221oi_1 _13792_ (.B2(_08105_),
    .C1(_08143_),
    .B1(_08136_),
    .A1(_08099_),
    .Y(_08144_),
    .A2(_08132_));
 sg13g2_buf_2 _13793_ (.A(_08144_),
    .X(_08145_));
 sg13g2_and2_1 _13794_ (.A(net1063),
    .B(_08038_),
    .X(_08146_));
 sg13g2_o21ai_1 _13795_ (.B1(_08052_),
    .Y(_08147_),
    .A1(_08146_),
    .A2(_08035_));
 sg13g2_nor2_1 _13796_ (.A(_08046_),
    .B(_08063_),
    .Y(_08148_));
 sg13g2_nor4_1 _13797_ (.A(_08055_),
    .B(_08056_),
    .C(_08057_),
    .D(_08063_),
    .Y(_08149_));
 sg13g2_a21oi_1 _13798_ (.A1(_08147_),
    .A2(_08148_),
    .Y(_08150_),
    .B1(_08149_));
 sg13g2_nand3b_1 _13799_ (.B(_08145_),
    .C(_08150_),
    .Y(_08151_),
    .A_N(_08027_));
 sg13g2_buf_1 _13800_ (.A(_08151_),
    .X(_08152_));
 sg13g2_buf_2 _13801_ (.A(\top_ihp.oisc.op_b[21] ),
    .X(_08153_));
 sg13g2_buf_2 _13802_ (.A(\top_ihp.oisc.op_a[24] ),
    .X(_08154_));
 sg13g2_buf_2 _13803_ (.A(\top_ihp.oisc.op_b[24] ),
    .X(_08155_));
 sg13g2_xor2_1 _13804_ (.B(_08155_),
    .A(_08154_),
    .X(_08156_));
 sg13g2_buf_2 _13805_ (.A(\top_ihp.oisc.op_a[25] ),
    .X(_08157_));
 sg13g2_buf_2 _13806_ (.A(\top_ihp.oisc.op_b[25] ),
    .X(_08158_));
 sg13g2_xor2_1 _13807_ (.B(_08158_),
    .A(_08157_),
    .X(_08159_));
 sg13g2_buf_2 _13808_ (.A(\top_ihp.oisc.op_a[22] ),
    .X(_08160_));
 sg13g2_buf_2 _13809_ (.A(\top_ihp.oisc.op_b[22] ),
    .X(_08161_));
 sg13g2_xor2_1 _13810_ (.B(_08161_),
    .A(_08160_),
    .X(_08162_));
 sg13g2_buf_1 _13811_ (.A(\top_ihp.oisc.op_a[23] ),
    .X(_08163_));
 sg13g2_buf_2 _13812_ (.A(\top_ihp.oisc.op_b[23] ),
    .X(_08164_));
 sg13g2_xor2_1 _13813_ (.B(_08164_),
    .A(net1061),
    .X(_08165_));
 sg13g2_nor4_1 _13814_ (.A(_08156_),
    .B(_08159_),
    .C(_08162_),
    .D(_08165_),
    .Y(_08166_));
 sg13g2_and2_1 _13815_ (.A(_08153_),
    .B(_08166_),
    .X(_08167_));
 sg13g2_nand3b_1 _13816_ (.B(_08152_),
    .C(_08167_),
    .Y(_08168_),
    .A_N(_08077_));
 sg13g2_buf_1 _13817_ (.A(\top_ihp.oisc.op_a[21] ),
    .X(_08169_));
 sg13g2_nor2b_1 _13818_ (.A(net1060),
    .B_N(_08166_),
    .Y(_08170_));
 sg13g2_nand3b_1 _13819_ (.B(_08152_),
    .C(_08170_),
    .Y(_08171_),
    .A_N(_08077_));
 sg13g2_nor2b_1 _13820_ (.A(_08154_),
    .B_N(_08155_),
    .Y(_08172_));
 sg13g2_nand2_1 _13821_ (.Y(_08173_),
    .A(_08158_),
    .B(_08172_));
 sg13g2_inv_1 _13822_ (.Y(_08174_),
    .A(_08157_));
 sg13g2_o21ai_1 _13823_ (.B1(_08174_),
    .Y(_08175_),
    .A1(_08158_),
    .A2(_08172_));
 sg13g2_nand2_1 _13824_ (.Y(_08176_),
    .A(_08173_),
    .B(_08175_));
 sg13g2_nor2b_1 _13825_ (.A(_08160_),
    .B_N(_08161_),
    .Y(_08177_));
 sg13g2_inv_1 _13826_ (.Y(_08178_),
    .A(net1061));
 sg13g2_a21oi_1 _13827_ (.A1(_08164_),
    .A2(_08177_),
    .Y(_08179_),
    .B1(_08178_));
 sg13g2_inv_1 _13828_ (.Y(_08180_),
    .A(_08160_));
 sg13g2_a21oi_1 _13829_ (.A1(_08180_),
    .A2(_08161_),
    .Y(_08181_),
    .B1(_08164_));
 sg13g2_nor4_1 _13830_ (.A(_08179_),
    .B(_08156_),
    .C(_08159_),
    .D(_08181_),
    .Y(_08182_));
 sg13g2_nor2b_1 _13831_ (.A(net1060),
    .B_N(_08153_),
    .Y(_08183_));
 sg13g2_buf_1 _13832_ (.A(_08183_),
    .X(_08184_));
 sg13g2_and2_1 _13833_ (.A(_08166_),
    .B(_08184_),
    .X(_08185_));
 sg13g2_nor3_1 _13834_ (.A(_08176_),
    .B(_08182_),
    .C(_08185_),
    .Y(_08186_));
 sg13g2_nand3_1 _13835_ (.B(_08171_),
    .C(_08186_),
    .A(_08168_),
    .Y(_08187_));
 sg13g2_buf_1 _13836_ (.A(_08187_),
    .X(_08188_));
 sg13g2_xnor2_1 _13837_ (.Y(_08189_),
    .A(_07989_),
    .B(_08188_));
 sg13g2_nor2_1 _13838_ (.A(net939),
    .B(_08189_),
    .Y(_08190_));
 sg13g2_xnor2_1 _13839_ (.Y(_08191_),
    .A(net974),
    .B(_08190_));
 sg13g2_buf_1 _13840_ (.A(\top_ihp.wb_spi.state ),
    .X(_08192_));
 sg13g2_buf_2 _13841_ (.A(_08192_),
    .X(_08193_));
 sg13g2_buf_1 _13842_ (.A(_08193_),
    .X(_08194_));
 sg13g2_buf_1 _13843_ (.A(_08194_),
    .X(_08195_));
 sg13g2_a21oi_1 _13844_ (.A1(net837),
    .A2(_08191_),
    .Y(_08196_),
    .B1(net972));
 sg13g2_buf_1 _13845_ (.A(\top_ihp.wb_spi.bits_left[0] ),
    .X(_08197_));
 sg13g2_buf_1 _13846_ (.A(\top_ihp.wb_spi.bits_left[1] ),
    .X(_08198_));
 sg13g2_or2_1 _13847_ (.X(_08199_),
    .B(\top_ihp.wb_spi.bits_left[2] ),
    .A(_08198_));
 sg13g2_buf_1 _13848_ (.A(_08199_),
    .X(_08200_));
 sg13g2_or3_1 _13849_ (.A(\top_ihp.wb_spi.bits_left[3] ),
    .B(\top_ihp.wb_spi.bits_left[4] ),
    .C(_08200_),
    .X(_08201_));
 sg13g2_nor2_1 _13850_ (.A(\top_ihp.wb_spi.bits_left[5] ),
    .B(_08201_),
    .Y(_08202_));
 sg13g2_nor2b_1 _13851_ (.A(\top_ihp.wb_spi.spi_clk_cnt[0] ),
    .B_N(\top_ihp.spi_clk_o ),
    .Y(_08203_));
 sg13g2_and4_1 _13852_ (.A(net1059),
    .B(_08192_),
    .C(_08202_),
    .D(_08203_),
    .X(_08204_));
 sg13g2_buf_1 _13853_ (.A(_08204_),
    .X(_08205_));
 sg13g2_nor2_1 _13854_ (.A(_08196_),
    .B(_08205_),
    .Y(_13605_));
 sg13g2_nand2_1 _13855_ (.Y(_08206_),
    .A(_07958_),
    .B(_07974_));
 sg13g2_buf_1 _13856_ (.A(_08206_),
    .X(_08207_));
 sg13g2_buf_1 _13857_ (.A(\top_ihp.oisc.decoder.decoded[11] ),
    .X(_08208_));
 sg13g2_o21ai_1 _13858_ (.B1(_07974_),
    .Y(_08209_),
    .A1(_07958_),
    .A2(net1058));
 sg13g2_buf_2 _13859_ (.A(_08209_),
    .X(_08210_));
 sg13g2_nor2_1 _13860_ (.A(net1047),
    .B(_08210_),
    .Y(_08211_));
 sg13g2_buf_2 _13861_ (.A(_08211_),
    .X(_08212_));
 sg13g2_buf_1 _13862_ (.A(_08212_),
    .X(_08213_));
 sg13g2_buf_1 _13863_ (.A(net809),
    .X(_08214_));
 sg13g2_nand2b_1 _13864_ (.Y(_08215_),
    .B(net790),
    .A_N(_08189_));
 sg13g2_nand2_1 _13865_ (.Y(_08216_),
    .A(_08189_),
    .B(net790));
 sg13g2_nor2_1 _13866_ (.A(net1019),
    .B(net974),
    .Y(_08217_));
 sg13g2_a221oi_1 _13867_ (.B2(_08217_),
    .C1(_08192_),
    .B1(_08216_),
    .A1(net974),
    .Y(_08218_),
    .A2(_08215_));
 sg13g2_a21o_1 _13868_ (.A2(_08218_),
    .A1(net883),
    .B1(_08205_),
    .X(_13604_));
 sg13g2_buf_1 _13869_ (.A(_00089_),
    .X(_08219_));
 sg13g2_inv_1 _13870_ (.Y(_08220_),
    .A(_07983_));
 sg13g2_buf_1 _13871_ (.A(_08220_),
    .X(_08221_));
 sg13g2_nand2b_1 _13872_ (.Y(_08222_),
    .B(net1017),
    .A_N(_08210_));
 sg13g2_buf_2 _13873_ (.A(_08222_),
    .X(_08223_));
 sg13g2_buf_1 _13874_ (.A(_08223_),
    .X(_08224_));
 sg13g2_nand2_1 _13875_ (.Y(_08225_),
    .A(_08045_),
    .B(_08048_));
 sg13g2_nor2_2 _13876_ (.A(_08225_),
    .B(_08063_),
    .Y(_08226_));
 sg13g2_nand2_1 _13877_ (.Y(_08227_),
    .A(_08042_),
    .B(_08043_));
 sg13g2_o21ai_1 _13878_ (.B1(_08039_),
    .Y(_08228_),
    .A1(_08028_),
    .A2(_08031_));
 sg13g2_o21ai_1 _13879_ (.B1(_08228_),
    .Y(_08229_),
    .A1(_08227_),
    .A2(_08145_));
 sg13g2_buf_2 _13880_ (.A(_08229_),
    .X(_08230_));
 sg13g2_inv_1 _13881_ (.Y(_08231_),
    .A(\top_ihp.oisc.op_b[14] ));
 sg13g2_nor2_1 _13882_ (.A(net1067),
    .B(_08231_),
    .Y(_08232_));
 sg13g2_nand2_1 _13883_ (.Y(_08233_),
    .A(net1046),
    .B(_08051_));
 sg13g2_inv_2 _13884_ (.Y(_08234_),
    .A(_08046_));
 sg13g2_o21ai_1 _13885_ (.B1(_08234_),
    .Y(_08235_),
    .A1(net1046),
    .A2(_08051_));
 sg13g2_a22oi_1 _13886_ (.Y(_08236_),
    .B1(_08233_),
    .B2(_08235_),
    .A2(_08231_),
    .A1(net1067));
 sg13g2_nor3_1 _13887_ (.A(_08009_),
    .B(_08232_),
    .C(_08236_),
    .Y(_08237_));
 sg13g2_o21ai_1 _13888_ (.B1(_08009_),
    .Y(_08238_),
    .A1(_08232_),
    .A2(_08236_));
 sg13g2_o21ai_1 _13889_ (.B1(_08238_),
    .Y(_08239_),
    .A1(net1068),
    .A2(_08237_));
 sg13g2_a21o_1 _13890_ (.A2(_08230_),
    .A1(_08226_),
    .B1(_08239_),
    .X(_08240_));
 sg13g2_nor2b_1 _13891_ (.A(_07999_),
    .B_N(net1071),
    .Y(_08241_));
 sg13g2_nor2_1 _13892_ (.A(_08000_),
    .B(net1071),
    .Y(_08242_));
 sg13g2_nand2b_1 _13893_ (.Y(_08243_),
    .B(_07996_),
    .A_N(net1070));
 sg13g2_nand2_1 _13894_ (.Y(_08244_),
    .A(_08071_),
    .B(_08243_));
 sg13g2_nor3_1 _13895_ (.A(_08241_),
    .B(_08242_),
    .C(_08244_),
    .Y(_08245_));
 sg13g2_nand2_1 _13896_ (.Y(_08246_),
    .A(_08067_),
    .B(_08245_));
 sg13g2_nor2b_1 _13897_ (.A(_08153_),
    .B_N(net1060),
    .Y(_08247_));
 sg13g2_buf_1 _13898_ (.A(_08247_),
    .X(_08248_));
 sg13g2_or4_1 _13899_ (.A(_08162_),
    .B(_08165_),
    .C(_08248_),
    .D(_08184_),
    .X(_08249_));
 sg13g2_nor4_1 _13900_ (.A(_07993_),
    .B(_08003_),
    .C(_08246_),
    .D(_08249_),
    .Y(_08250_));
 sg13g2_nor2b_1 _13901_ (.A(net1061),
    .B_N(_08164_),
    .Y(_08251_));
 sg13g2_buf_1 _13902_ (.A(_08251_),
    .X(_08252_));
 sg13g2_a21oi_1 _13903_ (.A1(_08240_),
    .A2(_08250_),
    .Y(_08253_),
    .B1(_08252_));
 sg13g2_nand2b_1 _13904_ (.Y(_08254_),
    .B(_07999_),
    .A_N(net1071));
 sg13g2_nand2_1 _13905_ (.Y(_08255_),
    .A(_08006_),
    .B(_08066_));
 sg13g2_inv_1 _13906_ (.Y(_08256_),
    .A(_08005_));
 sg13g2_o21ai_1 _13907_ (.B1(_08256_),
    .Y(_08257_),
    .A1(_08006_),
    .A2(_08066_));
 sg13g2_inv_1 _13908_ (.Y(_08258_),
    .A(_07996_));
 sg13g2_a21oi_1 _13909_ (.A1(_08255_),
    .A2(_08257_),
    .Y(_08259_),
    .B1(_08258_));
 sg13g2_nand3_1 _13910_ (.B(_08255_),
    .C(_08257_),
    .A(_08258_),
    .Y(_08260_));
 sg13g2_nor2_1 _13911_ (.A(net1070),
    .B(_08242_),
    .Y(_08261_));
 sg13g2_a221oi_1 _13912_ (.B2(_08261_),
    .C1(_08241_),
    .B1(_08260_),
    .A1(_08254_),
    .Y(_08262_),
    .A2(_08259_));
 sg13g2_buf_1 _13913_ (.A(_08262_),
    .X(_08263_));
 sg13g2_o21ai_1 _13914_ (.B1(_07990_),
    .Y(_08264_),
    .A1(_07991_),
    .A2(_08263_));
 sg13g2_a21oi_1 _13915_ (.A1(_07991_),
    .A2(_08263_),
    .Y(_08265_),
    .B1(_08248_));
 sg13g2_nand2b_1 _13916_ (.Y(_08266_),
    .B(_08153_),
    .A_N(net1060));
 sg13g2_nand2_1 _13917_ (.Y(_08267_),
    .A(_08160_),
    .B(_08266_));
 sg13g2_a21o_1 _13918_ (.A2(_08265_),
    .A1(_08264_),
    .B1(_08267_),
    .X(_08268_));
 sg13g2_nand2b_1 _13919_ (.Y(_08269_),
    .B(net1061),
    .A_N(_08164_));
 sg13g2_and2_1 _13920_ (.A(_08161_),
    .B(_08269_),
    .X(_08270_));
 sg13g2_nand2_1 _13921_ (.Y(_08271_),
    .A(_07991_),
    .B(_08263_));
 sg13g2_a21o_1 _13922_ (.A2(_08271_),
    .A1(_08264_),
    .B1(_08184_),
    .X(_08272_));
 sg13g2_nor2_1 _13923_ (.A(_08160_),
    .B(_08248_),
    .Y(_08273_));
 sg13g2_and2_1 _13924_ (.A(_08269_),
    .B(_08273_),
    .X(_08274_));
 sg13g2_a22oi_1 _13925_ (.Y(_08275_),
    .B1(_08272_),
    .B2(_08274_),
    .A2(_08270_),
    .A1(_08268_));
 sg13g2_buf_1 _13926_ (.A(\top_ihp.oisc.op_a[28] ),
    .X(_08276_));
 sg13g2_buf_1 _13927_ (.A(\top_ihp.oisc.op_b[28] ),
    .X(_08277_));
 sg13g2_xor2_1 _13928_ (.B(_08277_),
    .A(net1057),
    .X(_08278_));
 sg13g2_buf_1 _13929_ (.A(_08278_),
    .X(_08279_));
 sg13g2_xnor2_1 _13930_ (.Y(_08280_),
    .A(_08154_),
    .B(_08155_));
 sg13g2_xnor2_1 _13931_ (.Y(_08281_),
    .A(_08157_),
    .B(_08158_));
 sg13g2_xnor2_1 _13932_ (.Y(_08282_),
    .A(_07988_),
    .B(_07979_));
 sg13g2_buf_1 _13933_ (.A(\top_ihp.oisc.op_a[27] ),
    .X(_08283_));
 sg13g2_buf_2 _13934_ (.A(\top_ihp.oisc.op_b[27] ),
    .X(_08284_));
 sg13g2_xnor2_1 _13935_ (.Y(_08285_),
    .A(_08283_),
    .B(_08284_));
 sg13g2_and4_1 _13936_ (.A(_08280_),
    .B(_08281_),
    .C(_08282_),
    .D(_08285_),
    .X(_08286_));
 sg13g2_buf_1 _13937_ (.A(_08286_),
    .X(_08287_));
 sg13g2_nand2_1 _13938_ (.Y(_08288_),
    .A(_08279_),
    .B(_08287_));
 sg13g2_a21oi_1 _13939_ (.A1(_08253_),
    .A2(_08275_),
    .Y(_08289_),
    .B1(_08288_));
 sg13g2_buf_2 _13940_ (.A(_08283_),
    .X(_08290_));
 sg13g2_nand2b_1 _13941_ (.Y(_08291_),
    .B(_08284_),
    .A_N(net1044));
 sg13g2_nor2b_1 _13942_ (.A(_08284_),
    .B_N(net1044),
    .Y(_08292_));
 sg13g2_nor2_1 _13943_ (.A(_07982_),
    .B(_08176_),
    .Y(_08293_));
 sg13g2_a21oi_1 _13944_ (.A1(_07982_),
    .A2(_08176_),
    .Y(_08294_),
    .B1(_07988_));
 sg13g2_or3_1 _13945_ (.A(_08292_),
    .B(_08293_),
    .C(_08294_),
    .X(_08295_));
 sg13g2_nand2_1 _13946_ (.Y(_08296_),
    .A(_08291_),
    .B(_08295_));
 sg13g2_nor2_1 _13947_ (.A(_08279_),
    .B(_08296_),
    .Y(_08297_));
 sg13g2_and3_1 _13948_ (.X(_08298_),
    .A(_08253_),
    .B(_08275_),
    .C(_08297_));
 sg13g2_and2_1 _13949_ (.A(_08279_),
    .B(_08296_),
    .X(_08299_));
 sg13g2_nor3_1 _13950_ (.A(_08279_),
    .B(_08296_),
    .C(_08287_),
    .Y(_08300_));
 sg13g2_nor4_2 _13951_ (.A(_08289_),
    .B(_08298_),
    .C(_08299_),
    .Y(_08301_),
    .D(_08300_));
 sg13g2_nand2_1 _13952_ (.Y(_08302_),
    .A(net1019),
    .B(net1057));
 sg13g2_o21ai_1 _13953_ (.B1(_08302_),
    .Y(_08303_),
    .A1(net808),
    .A2(_08301_));
 sg13g2_and2_1 _13954_ (.A(_08219_),
    .B(_08303_),
    .X(_00004_));
 sg13g2_buf_2 _13955_ (.A(\top_ihp.wb_imem.state[0] ),
    .X(_08304_));
 sg13g2_inv_1 _13956_ (.Y(_08305_),
    .A(_08304_));
 sg13g2_buf_1 _13957_ (.A(\top_ihp.oisc.op_a[30] ),
    .X(_08306_));
 sg13g2_buf_1 _13958_ (.A(_08306_),
    .X(_08307_));
 sg13g2_nand2_1 _13959_ (.Y(_08308_),
    .A(net1019),
    .B(net1043));
 sg13g2_mux2_1 _13960_ (.A0(_08308_),
    .A1(_07958_),
    .S(_07974_),
    .X(_08309_));
 sg13g2_buf_1 _13961_ (.A(_08221_),
    .X(_08310_));
 sg13g2_inv_1 _13962_ (.Y(_08311_),
    .A(net1043));
 sg13g2_buf_2 _13963_ (.A(\top_ihp.oisc.op_b[30] ),
    .X(_08312_));
 sg13g2_nor2b_1 _13964_ (.A(_08312_),
    .B_N(net1058),
    .Y(_08313_));
 sg13g2_nand3_1 _13965_ (.B(_08311_),
    .C(_08313_),
    .A(net971),
    .Y(_08314_));
 sg13g2_inv_2 _13966_ (.Y(_08315_),
    .A(_08312_));
 sg13g2_nor2_1 _13967_ (.A(_08315_),
    .B(_08306_),
    .Y(_08316_));
 sg13g2_nand3_1 _13968_ (.B(net971),
    .C(_08316_),
    .A(net1058),
    .Y(_08317_));
 sg13g2_xnor2_1 _13969_ (.Y(_08318_),
    .A(_08160_),
    .B(_08161_));
 sg13g2_nor2b_1 _13970_ (.A(_08252_),
    .B_N(_08269_),
    .Y(_08319_));
 sg13g2_buf_2 _13971_ (.A(\top_ihp.oisc.op_a[29] ),
    .X(_08320_));
 sg13g2_buf_1 _13972_ (.A(\top_ihp.oisc.op_b[29] ),
    .X(_08321_));
 sg13g2_xor2_1 _13973_ (.B(_08321_),
    .A(_08320_),
    .X(_08322_));
 sg13g2_nor2_1 _13974_ (.A(_08279_),
    .B(_08322_),
    .Y(_08323_));
 sg13g2_and4_1 _13975_ (.A(_08318_),
    .B(_08319_),
    .C(_08287_),
    .D(_08323_),
    .X(_08324_));
 sg13g2_nor2b_1 _13976_ (.A(_08248_),
    .B_N(_08324_),
    .Y(_08325_));
 sg13g2_nand3b_1 _13977_ (.B(_08152_),
    .C(_08325_),
    .Y(_08326_),
    .A_N(_08077_));
 sg13g2_nor2_1 _13978_ (.A(_08176_),
    .B(_08182_),
    .Y(_08327_));
 sg13g2_inv_1 _13979_ (.Y(_08328_),
    .A(_08284_));
 sg13g2_nor2_1 _13980_ (.A(net1044),
    .B(_08328_),
    .Y(_08329_));
 sg13g2_a21oi_1 _13981_ (.A1(_07988_),
    .A2(_07981_),
    .Y(_08330_),
    .B1(_08329_));
 sg13g2_nand2b_1 _13982_ (.Y(_08331_),
    .B(net1057),
    .A_N(_08277_));
 sg13g2_inv_1 _13983_ (.Y(_08332_),
    .A(_08320_));
 sg13g2_a21o_1 _13984_ (.A2(_08331_),
    .A1(_08321_),
    .B1(_08332_),
    .X(_08333_));
 sg13g2_buf_1 _13985_ (.A(_08333_),
    .X(_08334_));
 sg13g2_nand2_1 _13986_ (.Y(_08335_),
    .A(_08277_),
    .B(_08334_));
 sg13g2_nand2b_1 _13987_ (.Y(_08336_),
    .B(_08334_),
    .A_N(net1057));
 sg13g2_nand2_1 _13988_ (.Y(_08337_),
    .A(_07989_),
    .B(net1048));
 sg13g2_nand2_1 _13989_ (.Y(_08338_),
    .A(net1044),
    .B(_08328_));
 sg13g2_o21ai_1 _13990_ (.B1(_08338_),
    .Y(_08339_),
    .A1(_08329_),
    .A2(_08337_));
 sg13g2_a221oi_1 _13991_ (.B2(_08336_),
    .C1(_08339_),
    .B1(_08335_),
    .A1(_08327_),
    .Y(_08340_),
    .A2(_08330_));
 sg13g2_nand2_1 _13992_ (.Y(_08341_),
    .A(_08338_),
    .B(_08337_));
 sg13g2_nand2_1 _13993_ (.Y(_08342_),
    .A(_08321_),
    .B(_08334_));
 sg13g2_a221oi_1 _13994_ (.B2(_08291_),
    .C1(_08342_),
    .B1(_08341_),
    .A1(_08327_),
    .Y(_08343_),
    .A2(_08330_));
 sg13g2_inv_1 _13995_ (.Y(_08344_),
    .A(_08321_));
 sg13g2_nand2b_1 _13996_ (.Y(_08345_),
    .B(_08277_),
    .A_N(net1057));
 sg13g2_nand2b_1 _13997_ (.Y(_08346_),
    .B(_08334_),
    .A_N(_08345_));
 sg13g2_o21ai_1 _13998_ (.B1(_08346_),
    .Y(_08347_),
    .A1(_08320_),
    .A2(_08344_));
 sg13g2_nor3_1 _13999_ (.A(_08340_),
    .B(_08343_),
    .C(_08347_),
    .Y(_08348_));
 sg13g2_nand2_1 _14000_ (.Y(_08349_),
    .A(_08184_),
    .B(_08324_));
 sg13g2_nand3_1 _14001_ (.B(_08348_),
    .C(_08349_),
    .A(_08326_),
    .Y(_08350_));
 sg13g2_buf_2 _14002_ (.A(_08350_),
    .X(_08351_));
 sg13g2_mux2_1 _14003_ (.A0(_08314_),
    .A1(_08317_),
    .S(_08351_),
    .X(_08352_));
 sg13g2_nand3_1 _14004_ (.B(_08312_),
    .C(net1043),
    .A(_08208_),
    .Y(_08353_));
 sg13g2_nand2_1 _14005_ (.Y(_08354_),
    .A(_08307_),
    .B(_08313_));
 sg13g2_mux2_1 _14006_ (.A0(_08353_),
    .A1(_08354_),
    .S(_08351_),
    .X(_08355_));
 sg13g2_and3_1 _14007_ (.X(_08356_),
    .A(_08308_),
    .B(_08352_),
    .C(_08355_));
 sg13g2_buf_1 _14008_ (.A(_08356_),
    .X(_08357_));
 sg13g2_or2_1 _14009_ (.X(_08358_),
    .B(_08357_),
    .A(_08309_));
 sg13g2_buf_2 _14010_ (.A(_08358_),
    .X(_08359_));
 sg13g2_buf_1 _14011_ (.A(\top_ihp.wb_imem.bits_left[0] ),
    .X(_08360_));
 sg13g2_inv_1 _14012_ (.Y(_08361_),
    .A(\top_ihp.wb_imem.bits_left[1] ));
 sg13g2_buf_8 _14013_ (.A(\top_ihp.wb_imem.bits_left[2] ),
    .X(_08362_));
 sg13g2_nor4_2 _14014_ (.A(_08362_),
    .B(\top_ihp.wb_imem.bits_left[3] ),
    .C(\top_ihp.wb_imem.bits_left[5] ),
    .Y(_08363_),
    .D(\top_ihp.wb_imem.bits_left[4] ));
 sg13g2_and3_1 _14015_ (.X(_08364_),
    .A(_08360_),
    .B(_08361_),
    .C(_08363_));
 sg13g2_buf_1 _14016_ (.A(_08364_),
    .X(_08365_));
 sg13g2_buf_1 _14017_ (.A(\top_ihp.wb_imem.state[2] ),
    .X(_08366_));
 sg13g2_nand2b_1 _14018_ (.Y(_08367_),
    .B(_08366_),
    .A_N(_08365_));
 sg13g2_o21ai_1 _14019_ (.B1(_08367_),
    .Y(_00001_),
    .A1(_08305_),
    .A2(_08359_));
 sg13g2_buf_1 _14020_ (.A(_00090_),
    .X(_08368_));
 sg13g2_nor2_2 _14021_ (.A(_08360_),
    .B(\top_ihp.wb_imem.bits_left[1] ),
    .Y(_08369_));
 sg13g2_and2_1 _14022_ (.A(_08363_),
    .B(_08369_),
    .X(_08370_));
 sg13g2_buf_2 _14023_ (.A(_08370_),
    .X(_08371_));
 sg13g2_buf_8 _14024_ (.A(_08371_),
    .X(_08372_));
 sg13g2_nand2_1 _14025_ (.Y(_08373_),
    .A(_08366_),
    .B(_08365_));
 sg13g2_o21ai_1 _14026_ (.B1(_08373_),
    .Y(_00000_),
    .A1(_08368_),
    .A2(_08372_));
 sg13g2_buf_2 _14027_ (.A(\top_ihp.wb_ack_coproc ),
    .X(_08374_));
 sg13g2_nor2b_1 _14028_ (.A(_08374_),
    .B_N(net1044),
    .Y(_08375_));
 sg13g2_nand3_1 _14029_ (.B(net809),
    .C(_08375_),
    .A(_08328_),
    .Y(_08376_));
 sg13g2_nor2_1 _14030_ (.A(_08374_),
    .B(net1044),
    .Y(_08377_));
 sg13g2_nand3_1 _14031_ (.B(_08212_),
    .C(_08377_),
    .A(_08284_),
    .Y(_08378_));
 sg13g2_nor2_1 _14032_ (.A(_08156_),
    .B(_08165_),
    .Y(_08379_));
 sg13g2_and3_1 _14033_ (.X(_08380_),
    .A(_08281_),
    .B(_08282_),
    .C(_08379_));
 sg13g2_buf_1 _14034_ (.A(_08380_),
    .X(_08381_));
 sg13g2_nor2b_1 _14035_ (.A(net1063),
    .B_N(_08028_),
    .Y(_08382_));
 sg13g2_nor2_1 _14036_ (.A(_08032_),
    .B(_08382_),
    .Y(_08383_));
 sg13g2_nand2_1 _14037_ (.Y(_08384_),
    .A(_08032_),
    .B(_08382_));
 sg13g2_o21ai_1 _14038_ (.B1(_08384_),
    .Y(_08385_),
    .A1(net1064),
    .A2(_08383_));
 sg13g2_nor2_1 _14039_ (.A(net1046),
    .B(_08385_),
    .Y(_08386_));
 sg13g2_a21oi_1 _14040_ (.A1(_08050_),
    .A2(_08385_),
    .Y(_08387_),
    .B1(_08234_));
 sg13g2_o21ai_1 _14041_ (.B1(_08016_),
    .Y(_08388_),
    .A1(_08386_),
    .A2(_08387_));
 sg13g2_nand2_1 _14042_ (.Y(_08389_),
    .A(_08061_),
    .B(_08388_));
 sg13g2_nor3_1 _14043_ (.A(_07993_),
    .B(_08003_),
    .C(_08246_),
    .Y(_08390_));
 sg13g2_nor3_2 _14044_ (.A(_08162_),
    .B(_08248_),
    .C(_08184_),
    .Y(_08391_));
 sg13g2_nand3_1 _14045_ (.B(_08390_),
    .C(_08391_),
    .A(_08060_),
    .Y(_08392_));
 sg13g2_inv_1 _14046_ (.Y(_08393_),
    .A(_08161_));
 sg13g2_a21oi_1 _14047_ (.A1(_08161_),
    .A2(_08184_),
    .Y(_08394_),
    .B1(_08180_));
 sg13g2_a21oi_1 _14048_ (.A1(_08393_),
    .A2(_08266_),
    .Y(_08395_),
    .B1(_08394_));
 sg13g2_inv_1 _14049_ (.Y(_08396_),
    .A(_08395_));
 sg13g2_o21ai_1 _14050_ (.B1(_08396_),
    .Y(_08397_),
    .A1(_08389_),
    .A2(_08392_));
 sg13g2_nand2_1 _14051_ (.Y(_08398_),
    .A(_08226_),
    .B(_08390_));
 sg13g2_inv_1 _14052_ (.Y(_08399_),
    .A(net1062));
 sg13g2_o21ai_1 _14053_ (.B1(net1045),
    .Y(_08400_),
    .A1(_08399_),
    .A2(_08129_));
 sg13g2_nand2_1 _14054_ (.Y(_08401_),
    .A(_08399_),
    .B(_08129_));
 sg13g2_a21oi_1 _14055_ (.A1(_08101_),
    .A2(_08119_),
    .Y(_08402_),
    .B1(_08112_));
 sg13g2_o21ai_1 _14056_ (.B1(_08402_),
    .Y(_08403_),
    .A1(_08100_),
    .A2(_08135_));
 sg13g2_a21oi_1 _14057_ (.A1(_08400_),
    .A2(_08401_),
    .Y(_08404_),
    .B1(_08403_));
 sg13g2_nand2_1 _14058_ (.Y(_08405_),
    .A(_08099_),
    .B(_08113_));
 sg13g2_inv_1 _14059_ (.Y(_08406_),
    .A(_08115_));
 sg13g2_inv_1 _14060_ (.Y(_08407_),
    .A(_08130_));
 sg13g2_a21oi_1 _14061_ (.A1(_08123_),
    .A2(_08130_),
    .Y(_08408_),
    .B1(_08139_));
 sg13g2_a221oi_1 _14062_ (.B2(_08407_),
    .C1(_08408_),
    .B1(_08399_),
    .A1(_08116_),
    .Y(_08409_),
    .A2(_08406_));
 sg13g2_o21ai_1 _14063_ (.B1(_08101_),
    .Y(_08410_),
    .A1(_08119_),
    .A2(_08409_));
 sg13g2_nor3_1 _14064_ (.A(_08101_),
    .B(_08119_),
    .C(_08409_),
    .Y(_08411_));
 sg13g2_a221oi_1 _14065_ (.B2(_08100_),
    .C1(_08411_),
    .B1(_08410_),
    .A1(_08404_),
    .Y(_08412_),
    .A2(_08405_));
 sg13g2_buf_1 _14066_ (.A(_08412_),
    .X(_08413_));
 sg13g2_inv_1 _14067_ (.Y(_08414_),
    .A(_08030_));
 sg13g2_nand2_1 _14068_ (.Y(_08415_),
    .A(net1065),
    .B(_08414_));
 sg13g2_and3_1 _14069_ (.X(_08416_),
    .A(_08042_),
    .B(_08415_),
    .C(_08105_));
 sg13g2_a21oi_1 _14070_ (.A1(_08414_),
    .A2(_08107_),
    .Y(_08417_),
    .B1(net1065));
 sg13g2_nor2_1 _14071_ (.A(_08414_),
    .B(_08107_),
    .Y(_08418_));
 sg13g2_nor2_1 _14072_ (.A(_08417_),
    .B(_08418_),
    .Y(_08419_));
 sg13g2_nor2b_1 _14073_ (.A(_08419_),
    .B_N(_08042_),
    .Y(_08420_));
 sg13g2_a21oi_1 _14074_ (.A1(_08413_),
    .A2(_08416_),
    .Y(_08421_),
    .B1(_08420_));
 sg13g2_nor2_1 _14075_ (.A(_07996_),
    .B(_08007_),
    .Y(_08422_));
 sg13g2_inv_1 _14076_ (.Y(_08423_),
    .A(net1070));
 sg13g2_a21oi_1 _14077_ (.A1(_07996_),
    .A2(_08007_),
    .Y(_08424_),
    .B1(_08423_));
 sg13g2_nor2_1 _14078_ (.A(_08422_),
    .B(_08424_),
    .Y(_08425_));
 sg13g2_nor2b_1 _14079_ (.A(net1068),
    .B_N(_08009_),
    .Y(_08426_));
 sg13g2_nor2_1 _14080_ (.A(net1066),
    .B(_08426_),
    .Y(_08427_));
 sg13g2_inv_1 _14081_ (.Y(_08428_),
    .A(_08010_));
 sg13g2_a21oi_1 _14082_ (.A1(net1066),
    .A2(_08426_),
    .Y(_08429_),
    .B1(_08428_));
 sg13g2_nor4_1 _14083_ (.A(_08064_),
    .B(_08244_),
    .C(_08427_),
    .D(_08429_),
    .Y(_08430_));
 sg13g2_o21ai_1 _14084_ (.B1(_07994_),
    .Y(_08431_),
    .A1(_08425_),
    .A2(_08430_));
 sg13g2_nor3_1 _14085_ (.A(_07994_),
    .B(_08425_),
    .C(_08430_),
    .Y(_08432_));
 sg13g2_a221oi_1 _14086_ (.B2(_08431_),
    .C1(_08432_),
    .B1(_07999_),
    .A1(_07990_),
    .Y(_08433_),
    .A2(_07991_));
 sg13g2_nor2_1 _14087_ (.A(_07993_),
    .B(_08433_),
    .Y(_08434_));
 sg13g2_o21ai_1 _14088_ (.B1(_08434_),
    .Y(_08435_),
    .A1(_08398_),
    .A2(_08421_));
 sg13g2_and2_1 _14089_ (.A(_08381_),
    .B(_08391_),
    .X(_08436_));
 sg13g2_inv_1 _14090_ (.Y(_08437_),
    .A(_08158_));
 sg13g2_nand2_1 _14091_ (.Y(_08438_),
    .A(_08155_),
    .B(_08252_));
 sg13g2_inv_1 _14092_ (.Y(_08439_),
    .A(_08154_));
 sg13g2_o21ai_1 _14093_ (.B1(_08439_),
    .Y(_08440_),
    .A1(_08155_),
    .A2(_08252_));
 sg13g2_a22oi_1 _14094_ (.Y(_08441_),
    .B1(_08438_),
    .B2(_08440_),
    .A2(_08437_),
    .A1(_08157_));
 sg13g2_a21oi_1 _14095_ (.A1(_08174_),
    .A2(_08158_),
    .Y(_08442_),
    .B1(_08441_));
 sg13g2_a21o_1 _14096_ (.A2(_08442_),
    .A1(net1048),
    .B1(_07989_),
    .X(_08443_));
 sg13g2_o21ai_1 _14097_ (.B1(_08443_),
    .Y(_08444_),
    .A1(net1048),
    .A2(_08442_));
 sg13g2_a221oi_1 _14098_ (.B2(_08436_),
    .C1(_08444_),
    .B1(_08435_),
    .A1(_08381_),
    .Y(_08445_),
    .A2(_08397_));
 sg13g2_buf_1 _14099_ (.A(_08445_),
    .X(_08446_));
 sg13g2_a21o_1 _14100_ (.A2(_08378_),
    .A1(_08376_),
    .B1(_08446_),
    .X(_08447_));
 sg13g2_nand4_1 _14101_ (.B(net809),
    .C(_08446_),
    .A(_08328_),
    .Y(_08448_),
    .D(_08377_));
 sg13g2_nand4_1 _14102_ (.B(net809),
    .C(_08446_),
    .A(_08284_),
    .Y(_08449_),
    .D(_08375_));
 sg13g2_nand3b_1 _14103_ (.B(net1044),
    .C(net1019),
    .Y(_08450_),
    .A_N(_08374_));
 sg13g2_nand4_1 _14104_ (.B(_08448_),
    .C(_08449_),
    .A(_08447_),
    .Y(_08451_),
    .D(_08450_));
 sg13g2_buf_1 _14105_ (.A(_08451_),
    .X(_00003_));
 sg13g2_inv_1 _14106_ (.Y(_08452_),
    .A(_08080_));
 sg13g2_xnor2_1 _14107_ (.Y(_08453_),
    .A(_08452_),
    .B(_08084_));
 sg13g2_a21o_1 _14108_ (.A2(_08453_),
    .A1(net809),
    .B1(net1019),
    .X(_08454_));
 sg13g2_nor2_1 _14109_ (.A(_08078_),
    .B(_08453_),
    .Y(_08455_));
 sg13g2_a22oi_1 _14110_ (.Y(_08456_),
    .B1(_08455_),
    .B2(_08213_),
    .A2(_08454_),
    .A1(_08078_));
 sg13g2_buf_2 _14111_ (.A(_08456_),
    .X(_08457_));
 sg13g2_inv_1 _14112_ (.Y(\top_ihp.oisc.wb_adr_o[1] ),
    .A(_08457_));
 sg13g2_o21ai_1 _14113_ (.B1(net971),
    .Y(_08458_),
    .A1(_08081_),
    .A2(_08210_));
 sg13g2_inv_1 _14114_ (.Y(_08459_),
    .A(_08081_));
 sg13g2_nor3_1 _14115_ (.A(_08459_),
    .B(_08082_),
    .C(_08223_),
    .Y(_08460_));
 sg13g2_a21o_1 _14116_ (.A2(_08458_),
    .A1(_08082_),
    .B1(_08460_),
    .X(_08461_));
 sg13g2_buf_2 _14117_ (.A(_08461_),
    .X(\top_ihp.oisc.wb_adr_o[0] ));
 sg13g2_buf_1 _14118_ (.A(_00093_),
    .X(_08462_));
 sg13g2_nand2b_1 _14119_ (.Y(_08463_),
    .B(_08152_),
    .A_N(_08077_));
 sg13g2_buf_2 _14120_ (.A(_08463_),
    .X(_08464_));
 sg13g2_nand2_1 _14121_ (.Y(_08465_),
    .A(_08291_),
    .B(_08338_));
 sg13g2_nor2_1 _14122_ (.A(_08279_),
    .B(_08465_),
    .Y(_08466_));
 sg13g2_nand3_1 _14123_ (.B(_08391_),
    .C(_08466_),
    .A(_08381_),
    .Y(_08467_));
 sg13g2_o21ai_1 _14124_ (.B1(_08345_),
    .Y(_08468_),
    .A1(_08292_),
    .A2(_08330_));
 sg13g2_nor2_1 _14125_ (.A(_07988_),
    .B(_07981_),
    .Y(_08469_));
 sg13g2_nor4_1 _14126_ (.A(_08186_),
    .B(_08279_),
    .C(_08469_),
    .D(_08465_),
    .Y(_08470_));
 sg13g2_a21oi_1 _14127_ (.A1(_08331_),
    .A2(_08468_),
    .Y(_08471_),
    .B1(_08470_));
 sg13g2_o21ai_1 _14128_ (.B1(_08471_),
    .Y(_08472_),
    .A1(_08464_),
    .A2(_08467_));
 sg13g2_xor2_1 _14129_ (.B(_08472_),
    .A(_08322_),
    .X(_08473_));
 sg13g2_buf_2 _14130_ (.A(\top_ihp.oisc.decoder.instruction[13] ),
    .X(_08474_));
 sg13g2_buf_1 _14131_ (.A(_08474_),
    .X(_08475_));
 sg13g2_buf_1 _14132_ (.A(_00074_),
    .X(_08476_));
 sg13g2_nor2b_1 _14133_ (.A(net1042),
    .B_N(_08476_),
    .Y(_08477_));
 sg13g2_buf_1 _14134_ (.A(_08477_),
    .X(_08478_));
 sg13g2_buf_8 _14135_ (.A(\top_ihp.oisc.decoder.instruction[12] ),
    .X(_08479_));
 sg13g2_nand2_1 _14136_ (.Y(_08480_),
    .A(_08474_),
    .B(_08476_));
 sg13g2_nand2_1 _14137_ (.Y(_08481_),
    .A(net1017),
    .B(_08210_));
 sg13g2_o21ai_1 _14138_ (.B1(_08481_),
    .Y(_08482_),
    .A1(net1056),
    .A2(_08480_));
 sg13g2_buf_2 _14139_ (.A(_08482_),
    .X(_08483_));
 sg13g2_o21ai_1 _14140_ (.B1(_08212_),
    .Y(_08484_),
    .A1(_08478_),
    .A2(_08483_));
 sg13g2_nand2_1 _14141_ (.Y(_08485_),
    .A(net1056),
    .B(net1042));
 sg13g2_nand4_1 _14142_ (.B(_08476_),
    .C(_08320_),
    .A(net1047),
    .Y(_08486_),
    .D(_08485_));
 sg13g2_o21ai_1 _14143_ (.B1(_08486_),
    .Y(_08487_),
    .A1(_08473_),
    .A2(_08484_));
 sg13g2_buf_2 _14144_ (.A(_08487_),
    .X(_08488_));
 sg13g2_buf_1 _14145_ (.A(\top_ihp.wb_uart.uart_rx.state[1] ),
    .X(_08489_));
 sg13g2_buf_1 _14146_ (.A(\top_ihp.wb_uart.uart_rx.state[0] ),
    .X(_08490_));
 sg13g2_nor2_1 _14147_ (.A(net1055),
    .B(_08490_),
    .Y(_08491_));
 sg13g2_nand4_1 _14148_ (.B(net883),
    .C(_08488_),
    .A(_08462_),
    .Y(_08492_),
    .D(_08491_));
 sg13g2_buf_1 _14149_ (.A(net2),
    .X(_08493_));
 sg13g2_buf_1 _14150_ (.A(\top_ihp.wb_uart.uart_rx.state[2] ),
    .X(_08494_));
 sg13g2_nand2b_1 _14151_ (.Y(_08495_),
    .B(_08490_),
    .A_N(_08494_));
 sg13g2_nor2_1 _14152_ (.A(_08489_),
    .B(_08495_),
    .Y(_08496_));
 sg13g2_buf_1 _14153_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[14] ),
    .X(_08497_));
 sg13g2_buf_1 _14154_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[13] ),
    .X(_08498_));
 sg13g2_nor4_1 _14155_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[15] ),
    .B(_08497_),
    .C(_08498_),
    .D(\top_ihp.wb_uart.uart_rx.cycle_cnt[16] ),
    .Y(_08499_));
 sg13g2_buf_1 _14156_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[18] ),
    .X(_08500_));
 sg13g2_nor4_1 _14157_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[21] ),
    .B(\top_ihp.wb_uart.uart_rx.cycle_cnt[19] ),
    .C(_08500_),
    .D(\top_ihp.wb_uart.uart_rx.cycle_cnt[17] ),
    .Y(_08501_));
 sg13g2_buf_1 _14158_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[27] ),
    .X(_08502_));
 sg13g2_buf_1 _14159_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[23] ),
    .X(_08503_));
 sg13g2_buf_2 _14160_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[20] ),
    .X(_08504_));
 sg13g2_nor4_1 _14161_ (.A(_08502_),
    .B(_08503_),
    .C(\top_ihp.wb_uart.uart_rx.cycle_cnt[22] ),
    .D(_08504_),
    .Y(_08505_));
 sg13g2_buf_1 _14162_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[26] ),
    .X(_08506_));
 sg13g2_buf_1 _14163_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[25] ),
    .X(_08507_));
 sg13g2_buf_1 _14164_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[24] ),
    .X(_08508_));
 sg13g2_nor3_1 _14165_ (.A(_08506_),
    .B(_08507_),
    .C(_08508_),
    .Y(_08509_));
 sg13g2_nand4_1 _14166_ (.B(_08501_),
    .C(_08505_),
    .A(_08499_),
    .Y(_08510_),
    .D(_08509_));
 sg13g2_buf_1 _14167_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[10] ),
    .X(_08511_));
 sg13g2_buf_1 _14168_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[29] ),
    .X(_08512_));
 sg13g2_nor4_1 _14169_ (.A(_08511_),
    .B(\top_ihp.wb_uart.uart_rx.cycle_cnt[31] ),
    .C(\top_ihp.wb_uart.uart_rx.cycle_cnt[30] ),
    .D(_08512_),
    .Y(_08513_));
 sg13g2_buf_1 _14170_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[11] ),
    .X(_08514_));
 sg13g2_nor4_1 _14171_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[12] ),
    .B(_08514_),
    .C(\top_ihp.wb_uart.uart_rx.cycle_cnt[9] ),
    .D(\top_ihp.wb_uart.uart_rx.cycle_cnt[28] ),
    .Y(_08515_));
 sg13g2_nand2_1 _14172_ (.Y(_08516_),
    .A(_08513_),
    .B(_08515_));
 sg13g2_buf_8 _14173_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[0] ),
    .X(_08517_));
 sg13g2_inv_1 _14174_ (.Y(_08518_),
    .A(_08517_));
 sg13g2_buf_1 _14175_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[6] ),
    .X(_08519_));
 sg13g2_buf_1 _14176_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[7] ),
    .X(_08520_));
 sg13g2_buf_2 _14177_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[4] ),
    .X(_08521_));
 sg13g2_inv_1 _14178_ (.Y(_08522_),
    .A(_08521_));
 sg13g2_buf_1 _14179_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[5] ),
    .X(_08523_));
 sg13g2_inv_1 _14180_ (.Y(_08524_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[8] ));
 sg13g2_nor4_1 _14181_ (.A(_08520_),
    .B(_08522_),
    .C(_08523_),
    .D(_08524_),
    .Y(_08525_));
 sg13g2_nand3_1 _14182_ (.B(_08519_),
    .C(_08525_),
    .A(_08518_),
    .Y(_08526_));
 sg13g2_buf_8 _14183_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[2] ),
    .X(_08527_));
 sg13g2_buf_8 _14184_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[3] ),
    .X(_08528_));
 sg13g2_buf_8 _14185_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[1] ),
    .X(_08529_));
 sg13g2_nand3b_1 _14186_ (.B(_08528_),
    .C(_08529_),
    .Y(_08530_),
    .A_N(_08527_));
 sg13g2_nor4_1 _14187_ (.A(_08510_),
    .B(_08516_),
    .C(_08526_),
    .D(_08530_),
    .Y(_08531_));
 sg13g2_buf_1 _14188_ (.A(_08531_),
    .X(_08532_));
 sg13g2_or2_1 _14189_ (.X(_08533_),
    .B(_08532_),
    .A(_08490_));
 sg13g2_buf_1 _14190_ (.A(_08533_),
    .X(_08534_));
 sg13g2_inv_1 _14191_ (.Y(_08535_),
    .A(_08490_));
 sg13g2_buf_2 _14192_ (.A(\top_ihp.wb_uart.uart_rx.bit_cnt[0] ),
    .X(_08536_));
 sg13g2_nand2_1 _14193_ (.Y(_08537_),
    .A(_08536_),
    .B(_08532_));
 sg13g2_buf_1 _14194_ (.A(\top_ihp.wb_uart.uart_rx.bit_cnt[1] ),
    .X(_08538_));
 sg13g2_buf_2 _14195_ (.A(\top_ihp.wb_uart.uart_rx.bit_cnt[2] ),
    .X(_08539_));
 sg13g2_nand2_1 _14196_ (.Y(_08540_),
    .A(_08538_),
    .B(_08539_));
 sg13g2_nor4_1 _14197_ (.A(_08535_),
    .B(\top_ihp.wb_uart.uart_rx.bit_cnt[3] ),
    .C(_08537_),
    .D(_08540_),
    .Y(_08541_));
 sg13g2_nand2_1 _14198_ (.Y(_08542_),
    .A(net1055),
    .B(_08462_));
 sg13g2_nor2_1 _14199_ (.A(_08541_),
    .B(_08542_),
    .Y(_08543_));
 sg13g2_a22oi_1 _14200_ (.Y(_08544_),
    .B1(_08534_),
    .B2(_08543_),
    .A2(_08496_),
    .A1(net1072));
 sg13g2_nand2_1 _14201_ (.Y(\top_ihp.wb_uart.uart_rx.next_state[0] ),
    .A(_08492_),
    .B(_08544_));
 sg13g2_nor3_1 _14202_ (.A(net1055),
    .B(net1072),
    .C(_08495_),
    .Y(_08545_));
 sg13g2_or2_1 _14203_ (.X(\top_ihp.wb_uart.uart_rx.next_state[1] ),
    .B(_08545_),
    .A(_08543_));
 sg13g2_nand2b_1 _14204_ (.Y(_08546_),
    .B(_08494_),
    .A_N(net1055));
 sg13g2_nand3_1 _14205_ (.B(_08462_),
    .C(_08541_),
    .A(net1055),
    .Y(_08547_));
 sg13g2_o21ai_1 _14206_ (.B1(_08547_),
    .Y(\top_ihp.wb_uart.uart_rx.next_state[2] ),
    .A1(_08534_),
    .A2(_08546_));
 sg13g2_a21o_1 _14207_ (.A2(_08532_),
    .A1(_08462_),
    .B1(_08494_),
    .X(_08548_));
 sg13g2_a22oi_1 _14208_ (.Y(_08549_),
    .B1(_08548_),
    .B2(net1055),
    .A2(_08534_),
    .A1(_08494_));
 sg13g2_nor2_1 _14209_ (.A(net2),
    .B(_08495_),
    .Y(_08550_));
 sg13g2_inv_1 _14210_ (.Y(_08551_),
    .A(_08543_));
 sg13g2_o21ai_1 _14211_ (.B1(_08551_),
    .Y(_08552_),
    .A1(net1055),
    .A2(_08550_));
 sg13g2_nand3_1 _14212_ (.B(_08549_),
    .C(_08552_),
    .A(_08492_),
    .Y(_08553_));
 sg13g2_buf_2 _14213_ (.A(_08553_),
    .X(_08554_));
 sg13g2_buf_8 _14214_ (.A(_08554_),
    .X(_08555_));
 sg13g2_nor2_1 _14215_ (.A(_08517_),
    .B(net159),
    .Y(_00005_));
 sg13g2_xnor2_1 _14216_ (.Y(_08556_),
    .A(_08517_),
    .B(_08529_));
 sg13g2_nor2_1 _14217_ (.A(net159),
    .B(_08556_),
    .Y(_00016_));
 sg13g2_nand2_1 _14218_ (.Y(_08557_),
    .A(_08517_),
    .B(_08529_));
 sg13g2_xor2_1 _14219_ (.B(_08557_),
    .A(_08527_),
    .X(_08558_));
 sg13g2_nor2_1 _14220_ (.A(net159),
    .B(_08558_),
    .Y(_00027_));
 sg13g2_nand3_1 _14221_ (.B(_08529_),
    .C(_08527_),
    .A(_08517_),
    .Y(_08559_));
 sg13g2_xor2_1 _14222_ (.B(_08559_),
    .A(_08528_),
    .X(_08560_));
 sg13g2_nor2_1 _14223_ (.A(net159),
    .B(_08560_),
    .Y(_00030_));
 sg13g2_and4_1 _14224_ (.A(_08517_),
    .B(_08529_),
    .C(_08528_),
    .D(_08527_),
    .X(_08561_));
 sg13g2_buf_1 _14225_ (.A(_08561_),
    .X(_08562_));
 sg13g2_xnor2_1 _14226_ (.Y(_08563_),
    .A(_08521_),
    .B(_08562_));
 sg13g2_nor2_1 _14227_ (.A(net159),
    .B(_08563_),
    .Y(_00031_));
 sg13g2_and2_1 _14228_ (.A(_08521_),
    .B(_08562_),
    .X(_08564_));
 sg13g2_xor2_1 _14229_ (.B(_08564_),
    .A(_00092_),
    .X(_08565_));
 sg13g2_nor2_1 _14230_ (.A(_08555_),
    .B(_08565_),
    .Y(_00032_));
 sg13g2_and2_1 _14231_ (.A(_08523_),
    .B(_08564_),
    .X(_08566_));
 sg13g2_buf_1 _14232_ (.A(_08566_),
    .X(_08567_));
 sg13g2_xnor2_1 _14233_ (.Y(_08568_),
    .A(_08519_),
    .B(_08567_));
 sg13g2_nor2_1 _14234_ (.A(net159),
    .B(_08568_),
    .Y(_00033_));
 sg13g2_inv_1 _14235_ (.Y(_08569_),
    .A(_08520_));
 sg13g2_nand2_1 _14236_ (.Y(_08570_),
    .A(_08519_),
    .B(_08567_));
 sg13g2_xnor2_1 _14237_ (.Y(_08571_),
    .A(_08569_),
    .B(_08570_));
 sg13g2_nor2_1 _14238_ (.A(net159),
    .B(_08571_),
    .Y(_00034_));
 sg13g2_and2_1 _14239_ (.A(_08519_),
    .B(_08520_),
    .X(_08572_));
 sg13g2_nand4_1 _14240_ (.B(_08523_),
    .C(_08562_),
    .A(_08521_),
    .Y(_08573_),
    .D(_08572_));
 sg13g2_buf_1 _14241_ (.A(_08573_),
    .X(_08574_));
 sg13g2_xnor2_1 _14242_ (.Y(_08575_),
    .A(_08524_),
    .B(_08574_));
 sg13g2_nor2_1 _14243_ (.A(_08555_),
    .B(_08575_),
    .Y(_00035_));
 sg13g2_o21ai_1 _14244_ (.B1(\top_ihp.wb_uart.uart_rx.cycle_cnt[9] ),
    .Y(_08576_),
    .A1(_08524_),
    .A2(_08574_));
 sg13g2_inv_1 _14245_ (.Y(_08577_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[9] ));
 sg13g2_nand4_1 _14246_ (.B(_08577_),
    .C(_08567_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[8] ),
    .Y(_08578_),
    .D(_08572_));
 sg13g2_a21oi_1 _14247_ (.A1(_08576_),
    .A2(_08578_),
    .Y(_00036_),
    .B1(_08554_));
 sg13g2_nor3_2 _14248_ (.A(_08524_),
    .B(_08577_),
    .C(_08574_),
    .Y(_08579_));
 sg13g2_xnor2_1 _14249_ (.Y(_08580_),
    .A(_08511_),
    .B(_08579_));
 sg13g2_nor2_1 _14250_ (.A(net159),
    .B(_08580_),
    .Y(_00006_));
 sg13g2_buf_8 _14251_ (.A(_08554_),
    .X(_08581_));
 sg13g2_nand2_1 _14252_ (.Y(_08582_),
    .A(_08511_),
    .B(_08579_));
 sg13g2_xor2_1 _14253_ (.B(_08582_),
    .A(_08514_),
    .X(_08583_));
 sg13g2_nor2_1 _14254_ (.A(net158),
    .B(_08583_),
    .Y(_00007_));
 sg13g2_nand3_1 _14255_ (.B(_08511_),
    .C(_08579_),
    .A(_08514_),
    .Y(_08584_));
 sg13g2_xor2_1 _14256_ (.B(_08584_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[12] ),
    .X(_08585_));
 sg13g2_nor2_1 _14257_ (.A(net158),
    .B(_08585_),
    .Y(_00008_));
 sg13g2_and4_1 _14258_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[12] ),
    .B(_08514_),
    .C(_08511_),
    .D(_08579_),
    .X(_08586_));
 sg13g2_buf_8 _14259_ (.A(_08586_),
    .X(_08587_));
 sg13g2_xnor2_1 _14260_ (.Y(_08588_),
    .A(_08498_),
    .B(_08587_));
 sg13g2_nor2_1 _14261_ (.A(net158),
    .B(_08588_),
    .Y(_00009_));
 sg13g2_nand2_1 _14262_ (.Y(_08589_),
    .A(_08498_),
    .B(_08587_));
 sg13g2_xor2_1 _14263_ (.B(_08589_),
    .A(_08497_),
    .X(_08590_));
 sg13g2_nor2_1 _14264_ (.A(net158),
    .B(_08590_),
    .Y(_00010_));
 sg13g2_nand3_1 _14265_ (.B(_08498_),
    .C(_08587_),
    .A(_08497_),
    .Y(_08591_));
 sg13g2_xor2_1 _14266_ (.B(_08591_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[15] ),
    .X(_08592_));
 sg13g2_nor2_1 _14267_ (.A(net158),
    .B(_08592_),
    .Y(_00011_));
 sg13g2_inv_1 _14268_ (.Y(_08593_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[16] ));
 sg13g2_nand4_1 _14269_ (.B(_08497_),
    .C(_08498_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[15] ),
    .Y(_08594_),
    .D(_08587_));
 sg13g2_xnor2_1 _14270_ (.Y(_08595_),
    .A(_08593_),
    .B(_08594_));
 sg13g2_nor2_1 _14271_ (.A(net158),
    .B(_08595_),
    .Y(_00012_));
 sg13g2_nor2_1 _14272_ (.A(_08593_),
    .B(_08594_),
    .Y(_08596_));
 sg13g2_xnor2_1 _14273_ (.Y(_08597_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[17] ),
    .B(_08596_));
 sg13g2_nor2_1 _14274_ (.A(_08581_),
    .B(_08597_),
    .Y(_00013_));
 sg13g2_and2_1 _14275_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[17] ),
    .B(_08596_),
    .X(_08598_));
 sg13g2_buf_8 _14276_ (.A(_08598_),
    .X(_08599_));
 sg13g2_xnor2_1 _14277_ (.Y(_08600_),
    .A(_08500_),
    .B(_08599_));
 sg13g2_nor2_1 _14278_ (.A(net158),
    .B(_08600_),
    .Y(_00014_));
 sg13g2_nand2_1 _14279_ (.Y(_08601_),
    .A(_08500_),
    .B(_08599_));
 sg13g2_xor2_1 _14280_ (.B(_08601_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[19] ),
    .X(_08602_));
 sg13g2_nor2_1 _14281_ (.A(net158),
    .B(_08602_),
    .Y(_00015_));
 sg13g2_and2_1 _14282_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[19] ),
    .B(_08500_),
    .X(_08603_));
 sg13g2_buf_1 _14283_ (.A(_08603_),
    .X(_08604_));
 sg13g2_nand2_1 _14284_ (.Y(_08605_),
    .A(_08599_),
    .B(_08604_));
 sg13g2_xor2_1 _14285_ (.B(_08605_),
    .A(_08504_),
    .X(_08606_));
 sg13g2_nor2_1 _14286_ (.A(_08581_),
    .B(_08606_),
    .Y(_00017_));
 sg13g2_buf_8 _14287_ (.A(_08554_),
    .X(_08607_));
 sg13g2_nand3_1 _14288_ (.B(_08599_),
    .C(_08604_),
    .A(_08504_),
    .Y(_08608_));
 sg13g2_xor2_1 _14289_ (.B(_08608_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[21] ),
    .X(_08609_));
 sg13g2_nor2_1 _14290_ (.A(_08607_),
    .B(_08609_),
    .Y(_00018_));
 sg13g2_inv_1 _14291_ (.Y(_08610_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[22] ));
 sg13g2_nand4_1 _14292_ (.B(_08504_),
    .C(_08599_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[21] ),
    .Y(_08611_),
    .D(_08604_));
 sg13g2_buf_1 _14293_ (.A(_08611_),
    .X(_08612_));
 sg13g2_xnor2_1 _14294_ (.Y(_08613_),
    .A(_08610_),
    .B(_08612_));
 sg13g2_nor2_1 _14295_ (.A(net157),
    .B(_08613_),
    .Y(_00019_));
 sg13g2_nor2_1 _14296_ (.A(_08610_),
    .B(_08612_),
    .Y(_08614_));
 sg13g2_buf_8 _14297_ (.A(_08614_),
    .X(_08615_));
 sg13g2_xnor2_1 _14298_ (.Y(_08616_),
    .A(_08503_),
    .B(_08615_));
 sg13g2_nor2_1 _14299_ (.A(net157),
    .B(_08616_),
    .Y(_00020_));
 sg13g2_nand2_1 _14300_ (.Y(_08617_),
    .A(_08503_),
    .B(_08615_));
 sg13g2_xor2_1 _14301_ (.B(_08617_),
    .A(_08508_),
    .X(_08618_));
 sg13g2_nor2_1 _14302_ (.A(net157),
    .B(_08618_),
    .Y(_00021_));
 sg13g2_nand3_1 _14303_ (.B(_08503_),
    .C(_08615_),
    .A(_08508_),
    .Y(_08619_));
 sg13g2_xor2_1 _14304_ (.B(_08619_),
    .A(_08507_),
    .X(_08620_));
 sg13g2_nor2_1 _14305_ (.A(_08607_),
    .B(_08620_),
    .Y(_00022_));
 sg13g2_and3_1 _14306_ (.X(_08621_),
    .A(_08507_),
    .B(_08508_),
    .C(_08503_));
 sg13g2_buf_1 _14307_ (.A(_08621_),
    .X(_08622_));
 sg13g2_nand2_1 _14308_ (.Y(_08623_),
    .A(_08615_),
    .B(_08622_));
 sg13g2_xor2_1 _14309_ (.B(_08623_),
    .A(_08506_),
    .X(_08624_));
 sg13g2_nor2_1 _14310_ (.A(net157),
    .B(_08624_),
    .Y(_00023_));
 sg13g2_nand3_1 _14311_ (.B(_08615_),
    .C(_08622_),
    .A(_08506_),
    .Y(_08625_));
 sg13g2_xor2_1 _14312_ (.B(_08625_),
    .A(_08502_),
    .X(_08626_));
 sg13g2_nor2_1 _14313_ (.A(net157),
    .B(_08626_),
    .Y(_00024_));
 sg13g2_nand4_1 _14314_ (.B(_08506_),
    .C(_08615_),
    .A(_08502_),
    .Y(_08627_),
    .D(_08622_));
 sg13g2_xor2_1 _14315_ (.B(_08627_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[28] ),
    .X(_08628_));
 sg13g2_nor2_1 _14316_ (.A(net157),
    .B(_08628_),
    .Y(_00025_));
 sg13g2_nand3_1 _14317_ (.B(_08508_),
    .C(_08503_),
    .A(_08507_),
    .Y(_08629_));
 sg13g2_nand4_1 _14318_ (.B(_08502_),
    .C(_08506_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[28] ),
    .Y(_08630_),
    .D(\top_ihp.wb_uart.uart_rx.cycle_cnt[22] ));
 sg13g2_nor3_2 _14319_ (.A(_08612_),
    .B(_08629_),
    .C(_08630_),
    .Y(_08631_));
 sg13g2_xnor2_1 _14320_ (.Y(_08632_),
    .A(_08512_),
    .B(_08631_));
 sg13g2_nor2_1 _14321_ (.A(net157),
    .B(_08632_),
    .Y(_00026_));
 sg13g2_nand2_1 _14322_ (.Y(_08633_),
    .A(_08512_),
    .B(_08631_));
 sg13g2_xor2_1 _14323_ (.B(_08633_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[30] ),
    .X(_08634_));
 sg13g2_nor2_1 _14324_ (.A(net157),
    .B(_08634_),
    .Y(_00028_));
 sg13g2_nand3_1 _14325_ (.B(_08512_),
    .C(_08631_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[30] ),
    .Y(_08635_));
 sg13g2_xor2_1 _14326_ (.B(_08635_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[31] ),
    .X(_08636_));
 sg13g2_nor2_1 _14327_ (.A(_08554_),
    .B(_08636_),
    .Y(_00029_));
 sg13g2_buf_1 _14328_ (.A(\top_ihp.wb_uart.uart_tx.state[0] ),
    .X(_08637_));
 sg13g2_inv_1 _14329_ (.Y(_08638_),
    .A(_08637_));
 sg13g2_buf_2 _14330_ (.A(\top_ihp.wb_uart.uart_tx.state[1] ),
    .X(_08639_));
 sg13g2_buf_1 _14331_ (.A(net857),
    .X(_08640_));
 sg13g2_and2_1 _14332_ (.A(net836),
    .B(_08488_),
    .X(_08641_));
 sg13g2_buf_2 _14333_ (.A(\top_ihp.wb_uart.uart_tx.bit_cnt[0] ),
    .X(_08642_));
 sg13g2_buf_2 _14334_ (.A(\top_ihp.wb_uart.uart_tx.bit_cnt[1] ),
    .X(_08643_));
 sg13g2_buf_1 _14335_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[25] ),
    .X(_08644_));
 sg13g2_buf_2 _14336_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[27] ),
    .X(_08645_));
 sg13g2_nor4_1 _14337_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[19] ),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[22] ),
    .C(_08644_),
    .D(_08645_),
    .Y(_08646_));
 sg13g2_buf_1 _14338_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[21] ),
    .X(_08647_));
 sg13g2_buf_1 _14339_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[23] ),
    .X(_08648_));
 sg13g2_nor4_1 _14340_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[18] ),
    .B(_08647_),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[20] ),
    .D(_08648_),
    .Y(_08649_));
 sg13g2_buf_1 _14341_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[29] ),
    .X(_08650_));
 sg13g2_buf_1 _14342_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[28] ),
    .X(_08651_));
 sg13g2_nor4_1 _14343_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[26] ),
    .B(_08650_),
    .C(_08651_),
    .D(\top_ihp.wb_uart.uart_tx.cycle_cnt[31] ),
    .Y(_08652_));
 sg13g2_buf_8 _14344_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[0] ),
    .X(_08653_));
 sg13g2_buf_8 _14345_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[1] ),
    .X(_08654_));
 sg13g2_inv_1 _14346_ (.Y(_08655_),
    .A(_08654_));
 sg13g2_buf_1 _14347_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[24] ),
    .X(_08656_));
 sg13g2_nor4_1 _14348_ (.A(_08653_),
    .B(_08655_),
    .C(_08656_),
    .D(\top_ihp.wb_uart.uart_tx.cycle_cnt[30] ),
    .Y(_08657_));
 sg13g2_nand4_1 _14349_ (.B(_08649_),
    .C(_08652_),
    .A(_08646_),
    .Y(_08658_),
    .D(_08657_));
 sg13g2_buf_1 _14350_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[9] ),
    .X(_08659_));
 sg13g2_inv_1 _14351_ (.Y(_08660_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[8] ));
 sg13g2_buf_1 _14352_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[16] ),
    .X(_08661_));
 sg13g2_nor4_1 _14353_ (.A(_08659_),
    .B(_08660_),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[10] ),
    .D(_08661_),
    .Y(_08662_));
 sg13g2_buf_8 _14354_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[2] ),
    .X(_08663_));
 sg13g2_buf_1 _14355_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[6] ),
    .X(_08664_));
 sg13g2_inv_1 _14356_ (.Y(_08665_),
    .A(_08664_));
 sg13g2_nor4_1 _14357_ (.A(_08663_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[5] ),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[7] ),
    .D(_08665_),
    .Y(_08666_));
 sg13g2_buf_1 _14358_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[14] ),
    .X(_08667_));
 sg13g2_nor4_1 _14359_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[13] ),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[12] ),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[15] ),
    .D(_08667_),
    .Y(_08668_));
 sg13g2_buf_1 _14360_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[11] ),
    .X(_08669_));
 sg13g2_buf_1 _14361_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[17] ),
    .X(_08670_));
 sg13g2_buf_8 _14362_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[3] ),
    .X(_08671_));
 sg13g2_nand2_1 _14363_ (.Y(_08672_),
    .A(_08671_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[4] ));
 sg13g2_nor3_1 _14364_ (.A(_08669_),
    .B(_08670_),
    .C(_08672_),
    .Y(_08673_));
 sg13g2_nand4_1 _14365_ (.B(_08666_),
    .C(_08668_),
    .A(_08662_),
    .Y(_08674_),
    .D(_08673_));
 sg13g2_nor2_1 _14366_ (.A(_08658_),
    .B(_08674_),
    .Y(_08675_));
 sg13g2_buf_1 _14367_ (.A(_08675_),
    .X(_08676_));
 sg13g2_nand4_1 _14368_ (.B(_08643_),
    .C(\top_ihp.wb_uart.uart_tx.bit_cnt[2] ),
    .A(_08642_),
    .Y(_08677_),
    .D(_08676_));
 sg13g2_o21ai_1 _14369_ (.B1(_08639_),
    .Y(_08678_),
    .A1(\top_ihp.wb_uart.uart_tx.bit_cnt[3] ),
    .A2(_08677_));
 sg13g2_o21ai_1 _14370_ (.B1(_08678_),
    .Y(_08679_),
    .A1(_08639_),
    .A2(_08641_));
 sg13g2_nand2_1 _14371_ (.Y(_08680_),
    .A(_08637_),
    .B(_08676_));
 sg13g2_inv_1 _14372_ (.Y(_08681_),
    .A(_08680_));
 sg13g2_a21oi_1 _14373_ (.A1(_08638_),
    .A2(_08679_),
    .Y(\top_ihp.wb_uart.uart_tx.next_state[0] ),
    .B1(_08681_));
 sg13g2_xnor2_1 _14374_ (.Y(\top_ihp.wb_uart.uart_tx.next_state[1] ),
    .A(_08639_),
    .B(_08680_));
 sg13g2_nor2_1 _14375_ (.A(_08639_),
    .B(_08637_),
    .Y(_08682_));
 sg13g2_nand2b_1 _14376_ (.Y(_08683_),
    .B(_08676_),
    .A_N(_08682_));
 sg13g2_nand3_1 _14377_ (.B(_08488_),
    .C(_08682_),
    .A(net857),
    .Y(_08684_));
 sg13g2_buf_2 _14378_ (.A(_08684_),
    .X(_08685_));
 sg13g2_nand2_1 _14379_ (.Y(_08686_),
    .A(_08683_),
    .B(net532));
 sg13g2_buf_8 _14380_ (.A(_08686_),
    .X(_08687_));
 sg13g2_buf_8 _14381_ (.A(_08687_),
    .X(_08688_));
 sg13g2_nor2_1 _14382_ (.A(_08653_),
    .B(net56),
    .Y(_00037_));
 sg13g2_xnor2_1 _14383_ (.Y(_08689_),
    .A(_08653_),
    .B(_08654_));
 sg13g2_nor2_1 _14384_ (.A(net56),
    .B(_08689_),
    .Y(_00048_));
 sg13g2_nand2_1 _14385_ (.Y(_08690_),
    .A(_08653_),
    .B(_08654_));
 sg13g2_xor2_1 _14386_ (.B(_08690_),
    .A(_08663_),
    .X(_08691_));
 sg13g2_nor2_1 _14387_ (.A(net56),
    .B(_08691_),
    .Y(_00059_));
 sg13g2_nand3_1 _14388_ (.B(_08654_),
    .C(_08663_),
    .A(_08653_),
    .Y(_08692_));
 sg13g2_buf_2 _14389_ (.A(_08692_),
    .X(_08693_));
 sg13g2_xor2_1 _14390_ (.B(_08693_),
    .A(_08671_),
    .X(_08694_));
 sg13g2_nor2_1 _14391_ (.A(net56),
    .B(_08694_),
    .Y(_00062_));
 sg13g2_nand4_1 _14392_ (.B(_08654_),
    .C(_08663_),
    .A(_08653_),
    .Y(_08695_),
    .D(_08671_));
 sg13g2_xor2_1 _14393_ (.B(_08695_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[4] ),
    .X(_08696_));
 sg13g2_nor2_1 _14394_ (.A(net56),
    .B(_08696_),
    .Y(_00063_));
 sg13g2_nor2_1 _14395_ (.A(_08672_),
    .B(_08693_),
    .Y(_08697_));
 sg13g2_xnor2_1 _14396_ (.Y(_08698_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[5] ),
    .B(_08697_));
 sg13g2_nor2_1 _14397_ (.A(net56),
    .B(_08698_),
    .Y(_00064_));
 sg13g2_nand3_1 _14398_ (.B(\top_ihp.wb_uart.uart_tx.cycle_cnt[5] ),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[4] ),
    .A(_08671_),
    .Y(_08699_));
 sg13g2_buf_1 _14399_ (.A(_08699_),
    .X(_08700_));
 sg13g2_nor2_1 _14400_ (.A(_08693_),
    .B(_08700_),
    .Y(_08701_));
 sg13g2_xnor2_1 _14401_ (.Y(_08702_),
    .A(_08664_),
    .B(_08701_));
 sg13g2_nor2_1 _14402_ (.A(_08688_),
    .B(_08702_),
    .Y(_00065_));
 sg13g2_nand2_1 _14403_ (.Y(_08703_),
    .A(_08664_),
    .B(_08701_));
 sg13g2_xor2_1 _14404_ (.B(_08703_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[7] ),
    .X(_08704_));
 sg13g2_nor2_1 _14405_ (.A(net56),
    .B(_08704_),
    .Y(_00066_));
 sg13g2_nand2_1 _14406_ (.Y(_08705_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[7] ),
    .B(_08664_));
 sg13g2_nor3_1 _14407_ (.A(_08693_),
    .B(_08700_),
    .C(_08705_),
    .Y(_08706_));
 sg13g2_xnor2_1 _14408_ (.Y(_08707_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[8] ),
    .B(_08706_));
 sg13g2_nor2_1 _14409_ (.A(_08688_),
    .B(_08707_),
    .Y(_00067_));
 sg13g2_nor4_2 _14410_ (.A(_08660_),
    .B(_08693_),
    .C(_08700_),
    .Y(_08708_),
    .D(_08705_));
 sg13g2_buf_8 _14411_ (.A(_08708_),
    .X(_08709_));
 sg13g2_xnor2_1 _14412_ (.Y(_08710_),
    .A(_08659_),
    .B(_08709_));
 sg13g2_nor2_1 _14413_ (.A(net56),
    .B(_08710_),
    .Y(_00068_));
 sg13g2_buf_8 _14414_ (.A(_08687_),
    .X(_08711_));
 sg13g2_nand2_1 _14415_ (.Y(_08712_),
    .A(_08659_),
    .B(_08709_));
 sg13g2_xor2_1 _14416_ (.B(_08712_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[10] ),
    .X(_08713_));
 sg13g2_nor2_1 _14417_ (.A(net55),
    .B(_08713_),
    .Y(_00038_));
 sg13g2_and2_1 _14418_ (.A(_08659_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[10] ),
    .X(_08714_));
 sg13g2_buf_1 _14419_ (.A(_08714_),
    .X(_08715_));
 sg13g2_nand2_1 _14420_ (.Y(_08716_),
    .A(_08709_),
    .B(_08715_));
 sg13g2_xor2_1 _14421_ (.B(_08716_),
    .A(_08669_),
    .X(_08717_));
 sg13g2_nor2_1 _14422_ (.A(net55),
    .B(_08717_),
    .Y(_00039_));
 sg13g2_nand3_1 _14423_ (.B(_08709_),
    .C(_08715_),
    .A(_08669_),
    .Y(_08718_));
 sg13g2_xor2_1 _14424_ (.B(_08718_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[12] ),
    .X(_08719_));
 sg13g2_nor2_1 _14425_ (.A(net55),
    .B(_08719_),
    .Y(_00040_));
 sg13g2_inv_1 _14426_ (.Y(_08720_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[13] ));
 sg13g2_nand4_1 _14427_ (.B(\top_ihp.wb_uart.uart_tx.cycle_cnt[12] ),
    .C(_08709_),
    .A(_08669_),
    .Y(_08721_),
    .D(_08715_));
 sg13g2_xnor2_1 _14428_ (.Y(_08722_),
    .A(_08720_),
    .B(_08721_));
 sg13g2_nor2_1 _14429_ (.A(net55),
    .B(_08722_),
    .Y(_00041_));
 sg13g2_nor2_1 _14430_ (.A(_08720_),
    .B(_08721_),
    .Y(_08723_));
 sg13g2_xnor2_1 _14431_ (.Y(_08724_),
    .A(_08667_),
    .B(_08723_));
 sg13g2_nor2_1 _14432_ (.A(_08711_),
    .B(_08724_),
    .Y(_00042_));
 sg13g2_nand2_1 _14433_ (.Y(_08725_),
    .A(_08667_),
    .B(_08723_));
 sg13g2_xor2_1 _14434_ (.B(_08725_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[15] ),
    .X(_08726_));
 sg13g2_nor2_1 _14435_ (.A(net55),
    .B(_08726_),
    .Y(_00043_));
 sg13g2_and3_1 _14436_ (.X(_08727_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[15] ),
    .B(_08667_),
    .C(_08723_));
 sg13g2_buf_8 _14437_ (.A(_08727_),
    .X(_08728_));
 sg13g2_xnor2_1 _14438_ (.Y(_08729_),
    .A(_08661_),
    .B(_08728_));
 sg13g2_nor2_1 _14439_ (.A(net55),
    .B(_08729_),
    .Y(_00044_));
 sg13g2_nand2_1 _14440_ (.Y(_08730_),
    .A(_08661_),
    .B(_08728_));
 sg13g2_xor2_1 _14441_ (.B(_08730_),
    .A(_08670_),
    .X(_08731_));
 sg13g2_nor2_1 _14442_ (.A(net55),
    .B(_08731_),
    .Y(_00045_));
 sg13g2_nand3_1 _14443_ (.B(_08661_),
    .C(_08728_),
    .A(_08670_),
    .Y(_08732_));
 sg13g2_xor2_1 _14444_ (.B(_08732_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[18] ),
    .X(_08733_));
 sg13g2_nor2_1 _14445_ (.A(net55),
    .B(_08733_),
    .Y(_00046_));
 sg13g2_inv_1 _14446_ (.Y(_08734_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[19] ));
 sg13g2_nand4_1 _14447_ (.B(_08661_),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[18] ),
    .A(_08670_),
    .Y(_08735_),
    .D(_08728_));
 sg13g2_buf_1 _14448_ (.A(_08735_),
    .X(_08736_));
 sg13g2_xnor2_1 _14449_ (.Y(_08737_),
    .A(_08734_),
    .B(_08736_));
 sg13g2_nor2_1 _14450_ (.A(_08711_),
    .B(_08737_),
    .Y(_00047_));
 sg13g2_buf_8 _14451_ (.A(_08687_),
    .X(_08738_));
 sg13g2_nor2_1 _14452_ (.A(_08734_),
    .B(_08736_),
    .Y(_08739_));
 sg13g2_xnor2_1 _14453_ (.Y(_08740_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[20] ),
    .B(_08739_));
 sg13g2_nor2_1 _14454_ (.A(net54),
    .B(_08740_),
    .Y(_00049_));
 sg13g2_inv_1 _14455_ (.Y(_08741_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[20] ));
 sg13g2_nor3_2 _14456_ (.A(_08734_),
    .B(_08741_),
    .C(_08736_),
    .Y(_08742_));
 sg13g2_xnor2_1 _14457_ (.Y(_08743_),
    .A(_08647_),
    .B(_08742_));
 sg13g2_nor2_1 _14458_ (.A(net54),
    .B(_08743_),
    .Y(_00050_));
 sg13g2_nand2_1 _14459_ (.Y(_08744_),
    .A(_08647_),
    .B(_08742_));
 sg13g2_xor2_1 _14460_ (.B(_08744_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[22] ),
    .X(_08745_));
 sg13g2_nor2_1 _14461_ (.A(net54),
    .B(_08745_),
    .Y(_00051_));
 sg13g2_and3_1 _14462_ (.X(_08746_),
    .A(_08647_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[22] ),
    .C(_08742_));
 sg13g2_buf_8 _14463_ (.A(_08746_),
    .X(_08747_));
 sg13g2_xnor2_1 _14464_ (.Y(_08748_),
    .A(_08648_),
    .B(_08747_));
 sg13g2_nor2_1 _14465_ (.A(net54),
    .B(_08748_),
    .Y(_00052_));
 sg13g2_nand2_1 _14466_ (.Y(_08749_),
    .A(_08648_),
    .B(_08747_));
 sg13g2_xor2_1 _14467_ (.B(_08749_),
    .A(_08656_),
    .X(_08750_));
 sg13g2_nor2_1 _14468_ (.A(net54),
    .B(_08750_),
    .Y(_00053_));
 sg13g2_nand3_1 _14469_ (.B(_08656_),
    .C(_08747_),
    .A(_08648_),
    .Y(_08751_));
 sg13g2_xor2_1 _14470_ (.B(_08751_),
    .A(_08644_),
    .X(_08752_));
 sg13g2_nor2_1 _14471_ (.A(net54),
    .B(_08752_),
    .Y(_00054_));
 sg13g2_nand4_1 _14472_ (.B(_08644_),
    .C(_08656_),
    .A(_08648_),
    .Y(_08753_),
    .D(_08747_));
 sg13g2_xor2_1 _14473_ (.B(_08753_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[26] ),
    .X(_08754_));
 sg13g2_nor2_1 _14474_ (.A(_08738_),
    .B(_08754_),
    .Y(_00055_));
 sg13g2_and4_1 _14475_ (.A(_08648_),
    .B(_08644_),
    .C(_08656_),
    .D(\top_ihp.wb_uart.uart_tx.cycle_cnt[26] ),
    .X(_08755_));
 sg13g2_and2_1 _14476_ (.A(_08747_),
    .B(_08755_),
    .X(_08756_));
 sg13g2_buf_8 _14477_ (.A(_08756_),
    .X(_08757_));
 sg13g2_xnor2_1 _14478_ (.Y(_08758_),
    .A(_08645_),
    .B(_08757_));
 sg13g2_nor2_1 _14479_ (.A(net54),
    .B(_08758_),
    .Y(_00056_));
 sg13g2_nand2_1 _14480_ (.Y(_08759_),
    .A(_08645_),
    .B(_08757_));
 sg13g2_xor2_1 _14481_ (.B(_08759_),
    .A(_08651_),
    .X(_08760_));
 sg13g2_nor2_1 _14482_ (.A(net54),
    .B(_08760_),
    .Y(_00057_));
 sg13g2_nand3_1 _14483_ (.B(_08651_),
    .C(_08757_),
    .A(_08645_),
    .Y(_08761_));
 sg13g2_xor2_1 _14484_ (.B(_08761_),
    .A(_08650_),
    .X(_08762_));
 sg13g2_nor2_1 _14485_ (.A(_08738_),
    .B(_08762_),
    .Y(_00058_));
 sg13g2_nand4_1 _14486_ (.B(_08650_),
    .C(_08651_),
    .A(_08645_),
    .Y(_08763_),
    .D(_08757_));
 sg13g2_xor2_1 _14487_ (.B(_08763_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[30] ),
    .X(_08764_));
 sg13g2_nor2_1 _14488_ (.A(_08687_),
    .B(_08764_),
    .Y(_00060_));
 sg13g2_and4_1 _14489_ (.A(_08645_),
    .B(_08650_),
    .C(_08651_),
    .D(\top_ihp.wb_uart.uart_tx.cycle_cnt[30] ),
    .X(_08765_));
 sg13g2_and2_1 _14490_ (.A(_08757_),
    .B(_08765_),
    .X(_08766_));
 sg13g2_xnor2_1 _14491_ (.Y(_08767_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[31] ),
    .B(_08766_));
 sg13g2_nor2_1 _14492_ (.A(_08687_),
    .B(_08767_),
    .Y(_00061_));
 sg13g2_nand3_1 _14493_ (.B(_08363_),
    .C(_08369_),
    .A(\top_ihp.wb_imem.state[1] ),
    .Y(_08768_));
 sg13g2_buf_1 _14494_ (.A(_08768_),
    .X(_08769_));
 sg13g2_buf_8 _14495_ (.A(_08769_),
    .X(_08770_));
 sg13g2_nor2_1 _14496_ (.A(_00112_),
    .B(net904),
    .Y(_08771_));
 sg13g2_buf_8 _14497_ (.A(\top_ihp.wb_imem.state[1] ),
    .X(_08772_));
 sg13g2_buf_1 _14498_ (.A(\top_ihp.wb_emem.last_bit ),
    .X(_08773_));
 sg13g2_buf_1 _14499_ (.A(\top_ihp.wb_emem.state[2] ),
    .X(_08774_));
 sg13g2_buf_1 _14500_ (.A(\top_ihp.wb_emem.state[3] ),
    .X(_08775_));
 sg13g2_nor2_1 _14501_ (.A(_08774_),
    .B(_08775_),
    .Y(_08776_));
 sg13g2_buf_1 _14502_ (.A(_08776_),
    .X(_08777_));
 sg13g2_buf_8 _14503_ (.A(\top_ihp.wb_emem.state[0] ),
    .X(_08778_));
 sg13g2_buf_8 _14504_ (.A(\top_ihp.wb_emem.state[1] ),
    .X(_08779_));
 sg13g2_and2_1 _14505_ (.A(_08778_),
    .B(_08779_),
    .X(_08780_));
 sg13g2_buf_8 _14506_ (.A(_08780_),
    .X(_08781_));
 sg13g2_nand3_1 _14507_ (.B(net970),
    .C(_08781_),
    .A(_08773_),
    .Y(_08782_));
 sg13g2_buf_1 _14508_ (.A(_08782_),
    .X(_08783_));
 sg13g2_buf_8 _14509_ (.A(_08783_),
    .X(_08784_));
 sg13g2_buf_8 _14510_ (.A(\top_ihp.wb_ack_spi ),
    .X(_08785_));
 sg13g2_inv_1 _14511_ (.Y(_08786_),
    .A(_00114_));
 sg13g2_nor2b_1 _14512_ (.A(_08785_),
    .B_N(_08374_),
    .Y(_08787_));
 sg13g2_buf_2 _14513_ (.A(_08787_),
    .X(_08788_));
 sg13g2_a22oi_1 _14514_ (.Y(_08789_),
    .B1(_08788_),
    .B2(\top_ihp.wb_coproc.dat_o[15] ),
    .A2(_08786_),
    .A1(_08785_));
 sg13g2_and4_1 _14515_ (.A(_08773_),
    .B(_00113_),
    .C(net970),
    .D(_08781_),
    .X(_08790_));
 sg13g2_a221oi_1 _14516_ (.B2(_08789_),
    .C1(_08790_),
    .B1(net891),
    .A1(net1041),
    .Y(_08791_),
    .A2(_08371_));
 sg13g2_buf_1 _14517_ (.A(\top_ihp.wb_ack_gpio ),
    .X(_08792_));
 sg13g2_nor2b_1 _14518_ (.A(_08792_),
    .B_N(_00075_),
    .Y(_08793_));
 sg13g2_buf_8 _14519_ (.A(_08793_),
    .X(_08794_));
 sg13g2_o21ai_1 _14520_ (.B1(_08794_),
    .Y(_08795_),
    .A1(_08771_),
    .A2(_08791_));
 sg13g2_buf_2 _14521_ (.A(_08795_),
    .X(_08796_));
 sg13g2_buf_1 _14522_ (.A(\top_ihp.wb_ack_uart ),
    .X(_08797_));
 sg13g2_nor2_1 _14523_ (.A(_08792_),
    .B(_08797_),
    .Y(_08798_));
 sg13g2_buf_2 _14524_ (.A(_08798_),
    .X(_08799_));
 sg13g2_nor2_1 _14525_ (.A(_08374_),
    .B(_08785_),
    .Y(_08800_));
 sg13g2_nand4_1 _14526_ (.B(_08783_),
    .C(_08799_),
    .A(_08769_),
    .Y(_08801_),
    .D(_08800_));
 sg13g2_buf_8 _14527_ (.A(_08801_),
    .X(_08802_));
 sg13g2_nand2_1 _14528_ (.Y(_08803_),
    .A(_07983_),
    .B(_08802_));
 sg13g2_buf_2 _14529_ (.A(_08803_),
    .X(_08804_));
 sg13g2_buf_8 _14530_ (.A(_08804_),
    .X(_08805_));
 sg13g2_buf_1 _14531_ (.A(net807),
    .X(_08806_));
 sg13g2_buf_1 _14532_ (.A(net789),
    .X(_08807_));
 sg13g2_buf_1 _14533_ (.A(net789),
    .X(_08808_));
 sg13g2_nand2_1 _14534_ (.Y(_08809_),
    .A(\top_ihp.oisc.decoder.instruction[15] ),
    .B(net768));
 sg13g2_o21ai_1 _14535_ (.B1(_08809_),
    .Y(_00204_),
    .A1(_08796_),
    .A2(net769));
 sg13g2_buf_1 _14536_ (.A(\top_ihp.oisc.micro_op[9] ),
    .X(_08810_));
 sg13g2_and2_1 _14537_ (.A(\top_ihp.oisc.micro_state[1] ),
    .B(_07959_),
    .X(_08811_));
 sg13g2_buf_1 _14538_ (.A(_08811_),
    .X(_08812_));
 sg13g2_nand2_1 _14539_ (.Y(_08813_),
    .A(_08810_),
    .B(net1016));
 sg13g2_inv_1 _14540_ (.Y(\top_ihp.oisc.reg_rb[1] ),
    .A(_08813_));
 sg13g2_buf_1 _14541_ (.A(\top_ihp.oisc.micro_op[8] ),
    .X(_08814_));
 sg13g2_nand2_1 _14542_ (.Y(_08815_),
    .A(_08814_),
    .B(net1016));
 sg13g2_inv_1 _14543_ (.Y(\top_ihp.oisc.reg_rb[0] ),
    .A(_08815_));
 sg13g2_nand2_1 _14544_ (.Y(_08816_),
    .A(\top_ihp.oisc.micro_op[11] ),
    .B(_08812_));
 sg13g2_buf_2 _14545_ (.A(_08816_),
    .X(_08817_));
 sg13g2_inv_1 _14546_ (.Y(\top_ihp.oisc.reg_rb[3] ),
    .A(_08817_));
 sg13g2_buf_2 _14547_ (.A(\top_ihp.oisc.micro_op[10] ),
    .X(_08818_));
 sg13g2_nand2_1 _14548_ (.Y(_08819_),
    .A(_08818_),
    .B(net1016));
 sg13g2_o21ai_1 _14549_ (.B1(_08819_),
    .Y(_08820_),
    .A1(_07973_),
    .A2(net1016));
 sg13g2_buf_2 _14550_ (.A(_08820_),
    .X(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_nand2_2 _14551_ (.Y(_08821_),
    .A(_07960_),
    .B(_07973_));
 sg13g2_inv_1 _14552_ (.Y(_08822_),
    .A(_00088_));
 sg13g2_buf_2 _14553_ (.A(\top_ihp.oisc.state[6] ),
    .X(_08823_));
 sg13g2_and4_1 _14554_ (.A(net904),
    .B(net891),
    .C(_08799_),
    .D(_08800_),
    .X(_08824_));
 sg13g2_buf_8 _14555_ (.A(_08824_),
    .X(_08825_));
 sg13g2_o21ai_1 _14556_ (.B1(net856),
    .Y(_08826_),
    .A1(_07985_),
    .A2(_08823_));
 sg13g2_buf_1 _14557_ (.A(_08826_),
    .X(_08827_));
 sg13g2_nand3_1 _14558_ (.B(_08822_),
    .C(net806),
    .A(_07961_),
    .Y(_08828_));
 sg13g2_nand2_1 _14559_ (.Y(_00002_),
    .A(_08821_),
    .B(_08828_));
 sg13g2_xor2_1 _14560_ (.B(\top_ihp.wb_spi.spi_clk_cnt[0] ),
    .A(\top_ihp.spi_clk_o ),
    .X(_00234_));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_nand2_2 _14562_ (.Y(_08829_),
    .A(net1049),
    .B(\top_ihp.oisc.micro_state[0] ));
 sg13g2_and2_1 _14563_ (.A(_07973_),
    .B(_08829_),
    .X(_08830_));
 sg13g2_buf_1 _14564_ (.A(_08830_),
    .X(_08831_));
 sg13g2_buf_1 _14565_ (.A(_08831_),
    .X(_08832_));
 sg13g2_buf_2 _14566_ (.A(\top_ihp.oisc.micro_pc[7] ),
    .X(_08833_));
 sg13g2_buf_1 _14567_ (.A(_08833_),
    .X(_08834_));
 sg13g2_buf_2 _14568_ (.A(\top_ihp.oisc.micro_pc[5] ),
    .X(_08835_));
 sg13g2_inv_2 _14569_ (.Y(_08836_),
    .A(_08835_));
 sg13g2_buf_1 _14570_ (.A(_08836_),
    .X(_08837_));
 sg13g2_buf_1 _14571_ (.A(net1015),
    .X(_08838_));
 sg13g2_buf_2 _14572_ (.A(\top_ihp.oisc.micro_pc[6] ),
    .X(_08839_));
 sg13g2_buf_1 _14573_ (.A(_08839_),
    .X(_08840_));
 sg13g2_buf_1 _14574_ (.A(net1039),
    .X(_08841_));
 sg13g2_buf_1 _14575_ (.A(\top_ihp.oisc.micro_pc[0] ),
    .X(_08842_));
 sg13g2_buf_1 _14576_ (.A(_08842_),
    .X(_08843_));
 sg13g2_inv_2 _14577_ (.Y(_08844_),
    .A(net1038));
 sg13g2_buf_1 _14578_ (.A(_08844_),
    .X(_08845_));
 sg13g2_buf_1 _14579_ (.A(_08845_),
    .X(_08846_));
 sg13g2_buf_2 _14580_ (.A(_00180_),
    .X(_08847_));
 sg13g2_inv_1 _14581_ (.Y(_08848_),
    .A(_08847_));
 sg13g2_buf_1 _14582_ (.A(_08848_),
    .X(_08849_));
 sg13g2_nor2_1 _14583_ (.A(net938),
    .B(net1013),
    .Y(_08850_));
 sg13g2_buf_1 _14584_ (.A(\top_ihp.oisc.micro_pc[1] ),
    .X(_08851_));
 sg13g2_inv_1 _14585_ (.Y(_08852_),
    .A(_08851_));
 sg13g2_buf_1 _14586_ (.A(_08852_),
    .X(_08853_));
 sg13g2_buf_1 _14587_ (.A(net1012),
    .X(_08854_));
 sg13g2_buf_1 _14588_ (.A(\top_ihp.oisc.micro_pc[3] ),
    .X(_08855_));
 sg13g2_buf_1 _14589_ (.A(\top_ihp.oisc.micro_pc[4] ),
    .X(_08856_));
 sg13g2_inv_1 _14590_ (.Y(_08857_),
    .A(net1053));
 sg13g2_buf_1 _14591_ (.A(_08857_),
    .X(_08858_));
 sg13g2_nand2_1 _14592_ (.Y(_08859_),
    .A(net1054),
    .B(net1011));
 sg13g2_buf_1 _14593_ (.A(_08859_),
    .X(_08860_));
 sg13g2_buf_1 _14594_ (.A(net1053),
    .X(_08861_));
 sg13g2_nand2_1 _14595_ (.Y(_08862_),
    .A(net1012),
    .B(net1037));
 sg13g2_buf_2 _14596_ (.A(_08862_),
    .X(_08863_));
 sg13g2_o21ai_1 _14597_ (.B1(_08863_),
    .Y(_08864_),
    .A1(_08854_),
    .A2(_08860_));
 sg13g2_buf_1 _14598_ (.A(net1038),
    .X(_08865_));
 sg13g2_buf_1 _14599_ (.A(\top_ihp.oisc.micro_pc[2] ),
    .X(_08866_));
 sg13g2_buf_1 _14600_ (.A(_08866_),
    .X(_08867_));
 sg13g2_inv_1 _14601_ (.Y(_08868_),
    .A(net1036));
 sg13g2_buf_2 _14602_ (.A(_08868_),
    .X(_08869_));
 sg13g2_nor2_1 _14603_ (.A(net1010),
    .B(_08869_),
    .Y(_08870_));
 sg13g2_buf_1 _14604_ (.A(_08870_),
    .X(_08871_));
 sg13g2_buf_1 _14605_ (.A(net1054),
    .X(_08872_));
 sg13g2_buf_1 _14606_ (.A(net1035),
    .X(_08873_));
 sg13g2_nor2_1 _14607_ (.A(net1009),
    .B(net1053),
    .Y(_08874_));
 sg13g2_buf_1 _14608_ (.A(_08874_),
    .X(_08875_));
 sg13g2_a22oi_1 _14609_ (.Y(_08876_),
    .B1(_08871_),
    .B2(net936),
    .A2(_08864_),
    .A1(_08850_));
 sg13g2_buf_1 _14610_ (.A(_08851_),
    .X(_08877_));
 sg13g2_nor2_1 _14611_ (.A(net1038),
    .B(_08877_),
    .Y(_08878_));
 sg13g2_buf_2 _14612_ (.A(_08878_),
    .X(_08879_));
 sg13g2_buf_1 _14613_ (.A(_08879_),
    .X(_08880_));
 sg13g2_buf_1 _14614_ (.A(_08847_),
    .X(_08881_));
 sg13g2_inv_2 _14615_ (.Y(_08882_),
    .A(net1054));
 sg13g2_nor2_2 _14616_ (.A(net1033),
    .B(_08882_),
    .Y(_08883_));
 sg13g2_nand2_2 _14617_ (.Y(_08884_),
    .A(_08843_),
    .B(net1036));
 sg13g2_buf_1 _14618_ (.A(net1034),
    .X(_08885_));
 sg13g2_nand2_1 _14619_ (.Y(_08886_),
    .A(net1008),
    .B(net1053));
 sg13g2_buf_1 _14620_ (.A(_08886_),
    .X(_08887_));
 sg13g2_buf_1 _14621_ (.A(_08869_),
    .X(_08888_));
 sg13g2_buf_1 _14622_ (.A(_08861_),
    .X(_08889_));
 sg13g2_nor2_1 _14623_ (.A(_08888_),
    .B(net1007),
    .Y(_08890_));
 sg13g2_buf_1 _14624_ (.A(net1036),
    .X(_08891_));
 sg13g2_nor2_1 _14625_ (.A(net1006),
    .B(_08887_),
    .Y(_08892_));
 sg13g2_o21ai_1 _14626_ (.B1(net968),
    .Y(_08893_),
    .A1(_08890_),
    .A2(_08892_));
 sg13g2_o21ai_1 _14627_ (.B1(_08893_),
    .Y(_08894_),
    .A1(_08884_),
    .A2(_08887_));
 sg13g2_buf_1 _14628_ (.A(net1039),
    .X(_08895_));
 sg13g2_a221oi_1 _14629_ (.B2(_08882_),
    .C1(net1005),
    .B1(_08894_),
    .A1(net935),
    .Y(_08896_),
    .A2(_08883_));
 sg13g2_a21oi_1 _14630_ (.A1(net1014),
    .A2(_08876_),
    .Y(_08897_),
    .B1(_08896_));
 sg13g2_buf_1 _14631_ (.A(net1008),
    .X(_08898_));
 sg13g2_buf_1 _14632_ (.A(net966),
    .X(_08899_));
 sg13g2_buf_1 _14633_ (.A(net933),
    .X(_08900_));
 sg13g2_nor2_1 _14634_ (.A(net903),
    .B(_08840_),
    .Y(_08901_));
 sg13g2_buf_1 _14635_ (.A(net1010),
    .X(_08902_));
 sg13g2_buf_1 _14636_ (.A(net965),
    .X(_08903_));
 sg13g2_buf_1 _14637_ (.A(_08903_),
    .X(_08904_));
 sg13g2_nand2_2 _14638_ (.Y(_08905_),
    .A(net1013),
    .B(net1037));
 sg13g2_nor2_1 _14639_ (.A(_08848_),
    .B(net1009),
    .Y(_08906_));
 sg13g2_buf_1 _14640_ (.A(_08906_),
    .X(_08907_));
 sg13g2_buf_1 _14641_ (.A(_08861_),
    .X(_08908_));
 sg13g2_nor2_1 _14642_ (.A(net968),
    .B(_08908_),
    .Y(_08909_));
 sg13g2_nand2_1 _14643_ (.Y(_08910_),
    .A(_08907_),
    .B(_08909_));
 sg13g2_o21ai_1 _14644_ (.B1(_08910_),
    .Y(_08911_),
    .A1(net902),
    .A2(_08905_));
 sg13g2_buf_1 _14645_ (.A(net1009),
    .X(_08912_));
 sg13g2_buf_1 _14646_ (.A(net964),
    .X(_08913_));
 sg13g2_nor2_1 _14647_ (.A(net1038),
    .B(net1036),
    .Y(_08914_));
 sg13g2_buf_1 _14648_ (.A(_08914_),
    .X(_08915_));
 sg13g2_nor2_1 _14649_ (.A(net1012),
    .B(net1007),
    .Y(_08916_));
 sg13g2_nor2_1 _14650_ (.A(_08866_),
    .B(_08852_),
    .Y(_08917_));
 sg13g2_buf_2 _14651_ (.A(_08917_),
    .X(_08918_));
 sg13g2_nor2_2 _14652_ (.A(_08869_),
    .B(net1034),
    .Y(_08919_));
 sg13g2_o21ai_1 _14653_ (.B1(net1010),
    .Y(_08920_),
    .A1(_08918_),
    .A2(_08919_));
 sg13g2_nand2_1 _14654_ (.Y(_08921_),
    .A(_08869_),
    .B(_08879_));
 sg13g2_nand2_1 _14655_ (.Y(_08922_),
    .A(_08920_),
    .B(_08921_));
 sg13g2_buf_1 _14656_ (.A(net1007),
    .X(_08923_));
 sg13g2_a22oi_1 _14657_ (.Y(_08924_),
    .B1(_08922_),
    .B2(net962),
    .A2(_08916_),
    .A1(net963));
 sg13g2_nor2_1 _14658_ (.A(_08882_),
    .B(net1011),
    .Y(_08925_));
 sg13g2_buf_2 _14659_ (.A(_08925_),
    .X(_08926_));
 sg13g2_and2_1 _14660_ (.A(net966),
    .B(net963),
    .X(_08927_));
 sg13g2_buf_1 _14661_ (.A(_08927_),
    .X(_08928_));
 sg13g2_nand2_1 _14662_ (.Y(_08929_),
    .A(_08926_),
    .B(_08928_));
 sg13g2_o21ai_1 _14663_ (.B1(_08929_),
    .Y(_08930_),
    .A1(_08913_),
    .A2(_08924_));
 sg13g2_a22oi_1 _14664_ (.Y(_08931_),
    .B1(_08930_),
    .B2(net1005),
    .A2(_08911_),
    .A1(_08901_));
 sg13g2_nor2_1 _14665_ (.A(net969),
    .B(_08931_),
    .Y(_08932_));
 sg13g2_a21oi_1 _14666_ (.A1(net969),
    .A2(_08897_),
    .Y(_08933_),
    .B1(_08932_));
 sg13g2_inv_1 _14667_ (.Y(_08934_),
    .A(_08839_));
 sg13g2_buf_1 _14668_ (.A(_08934_),
    .X(_08935_));
 sg13g2_buf_1 _14669_ (.A(net1036),
    .X(_08936_));
 sg13g2_buf_1 _14670_ (.A(net1002),
    .X(_08937_));
 sg13g2_buf_1 _14671_ (.A(net961),
    .X(_08938_));
 sg13g2_buf_1 _14672_ (.A(net966),
    .X(_08939_));
 sg13g2_buf_1 _14673_ (.A(net1011),
    .X(_08940_));
 sg13g2_buf_2 _14674_ (.A(_00179_),
    .X(_08941_));
 sg13g2_nor2_2 _14675_ (.A(net960),
    .B(_08941_),
    .Y(_08942_));
 sg13g2_nor2_1 _14676_ (.A(_08882_),
    .B(net1053),
    .Y(_08943_));
 sg13g2_buf_1 _14677_ (.A(_08943_),
    .X(_08944_));
 sg13g2_a21oi_1 _14678_ (.A1(net1007),
    .A2(_08941_),
    .Y(_08945_),
    .B1(_08944_));
 sg13g2_buf_1 _14679_ (.A(net1010),
    .X(_08946_));
 sg13g2_buf_1 _14680_ (.A(net959),
    .X(_08947_));
 sg13g2_a22oi_1 _14681_ (.Y(_08948_),
    .B1(_08945_),
    .B2(_08947_),
    .A2(_08942_),
    .A1(net929));
 sg13g2_nor2_1 _14682_ (.A(net930),
    .B(_08948_),
    .Y(_08949_));
 sg13g2_nor2_1 _14683_ (.A(net937),
    .B(_08884_),
    .Y(_08950_));
 sg13g2_o21ai_1 _14684_ (.B1(net969),
    .Y(_08951_),
    .A1(_08949_),
    .A2(_08950_));
 sg13g2_buf_1 _14685_ (.A(_08835_),
    .X(_08952_));
 sg13g2_buf_1 _14686_ (.A(net1032),
    .X(_08953_));
 sg13g2_buf_1 _14687_ (.A(_08953_),
    .X(_08954_));
 sg13g2_nand2_1 _14688_ (.Y(_08955_),
    .A(net1038),
    .B(net1034));
 sg13g2_buf_1 _14689_ (.A(_08955_),
    .X(_08956_));
 sg13g2_nor2_1 _14690_ (.A(_08847_),
    .B(net1035),
    .Y(_08957_));
 sg13g2_buf_2 _14691_ (.A(_08957_),
    .X(_08958_));
 sg13g2_nand4_1 _14692_ (.B(_08863_),
    .C(net957),
    .A(net958),
    .Y(_08959_),
    .D(_08958_));
 sg13g2_nand3_1 _14693_ (.B(_08951_),
    .C(_08959_),
    .A(net1003),
    .Y(_08960_));
 sg13g2_buf_1 _14694_ (.A(_00177_),
    .X(_08961_));
 sg13g2_nand2_1 _14695_ (.Y(_08962_),
    .A(_08839_),
    .B(_08961_));
 sg13g2_nand3_1 _14696_ (.B(_08960_),
    .C(_08962_),
    .A(net1040),
    .Y(_08963_));
 sg13g2_o21ai_1 _14697_ (.B1(_08963_),
    .Y(_08964_),
    .A1(net1040),
    .A2(_08933_));
 sg13g2_buf_1 _14698_ (.A(_08831_),
    .X(_08965_));
 sg13g2_nand2_1 _14699_ (.Y(_08966_),
    .A(_07963_),
    .B(net881));
 sg13g2_o21ai_1 _14700_ (.B1(_08966_),
    .Y(_00363_),
    .A1(net882),
    .A2(_08964_));
 sg13g2_inv_1 _14701_ (.Y(_08967_),
    .A(_08833_));
 sg13g2_buf_1 _14702_ (.A(_08967_),
    .X(_08968_));
 sg13g2_buf_1 _14703_ (.A(net1005),
    .X(_08969_));
 sg13g2_nand2_2 _14704_ (.Y(_08970_),
    .A(_08844_),
    .B(_08853_));
 sg13g2_nor2_1 _14705_ (.A(net934),
    .B(_08970_),
    .Y(_08971_));
 sg13g2_nor2_1 _14706_ (.A(net1006),
    .B(net957),
    .Y(_08972_));
 sg13g2_o21ai_1 _14707_ (.B1(_08945_),
    .Y(_08973_),
    .A1(_08971_),
    .A2(_08972_));
 sg13g2_o21ai_1 _14708_ (.B1(_08973_),
    .Y(_08974_),
    .A1(net937),
    .A2(_08921_));
 sg13g2_buf_1 _14709_ (.A(_08944_),
    .X(_08975_));
 sg13g2_nor2_1 _14710_ (.A(_08844_),
    .B(_08936_),
    .Y(_08976_));
 sg13g2_buf_2 _14711_ (.A(_08976_),
    .X(_08977_));
 sg13g2_nor2_1 _14712_ (.A(net1054),
    .B(net1011),
    .Y(_08978_));
 sg13g2_buf_2 _14713_ (.A(_08978_),
    .X(_08979_));
 sg13g2_a22oi_1 _14714_ (.Y(_08980_),
    .B1(_08977_),
    .B2(_08979_),
    .A2(net927),
    .A1(net930));
 sg13g2_nor2_1 _14715_ (.A(net966),
    .B(_08835_),
    .Y(_08981_));
 sg13g2_nor2b_1 _14716_ (.A(_08980_),
    .B_N(_08981_),
    .Y(_08982_));
 sg13g2_a21oi_1 _14717_ (.A1(net958),
    .A2(_08974_),
    .Y(_08983_),
    .B1(_08982_));
 sg13g2_nor2_1 _14718_ (.A(net1037),
    .B(_08836_),
    .Y(_08984_));
 sg13g2_buf_1 _14719_ (.A(_08984_),
    .X(_08985_));
 sg13g2_nand2_1 _14720_ (.Y(_08986_),
    .A(_08848_),
    .B(_08882_));
 sg13g2_nor2_1 _14721_ (.A(net1034),
    .B(_08847_),
    .Y(_08987_));
 sg13g2_nor2b_1 _14722_ (.A(net1038),
    .B_N(_08855_),
    .Y(_08988_));
 sg13g2_o21ai_1 _14723_ (.B1(_08988_),
    .Y(_08989_),
    .A1(_08918_),
    .A2(_08987_));
 sg13g2_o21ai_1 _14724_ (.B1(_08989_),
    .Y(_08990_),
    .A1(net957),
    .A2(_08986_));
 sg13g2_nor2_1 _14725_ (.A(net1012),
    .B(net1011),
    .Y(_08991_));
 sg13g2_nor2_1 _14726_ (.A(_08847_),
    .B(net1053),
    .Y(_08992_));
 sg13g2_buf_2 _14727_ (.A(_08992_),
    .X(_08993_));
 sg13g2_nor2_2 _14728_ (.A(net1008),
    .B(_08858_),
    .Y(_08994_));
 sg13g2_a21o_1 _14729_ (.A2(_08993_),
    .A1(net966),
    .B1(_08994_),
    .X(_08995_));
 sg13g2_a22oi_1 _14730_ (.Y(_08996_),
    .B1(_08995_),
    .B2(net928),
    .A2(_08871_),
    .A1(_08991_));
 sg13g2_nand2_1 _14731_ (.Y(_08997_),
    .A(_08856_),
    .B(_08835_));
 sg13g2_buf_1 _14732_ (.A(_08997_),
    .X(_08998_));
 sg13g2_nor2_1 _14733_ (.A(net1033),
    .B(_08970_),
    .Y(_08999_));
 sg13g2_nand2b_1 _14734_ (.Y(_09000_),
    .B(_08999_),
    .A_N(net999));
 sg13g2_o21ai_1 _14735_ (.B1(_09000_),
    .Y(_09001_),
    .A1(net1001),
    .A2(_08996_));
 sg13g2_inv_1 _14736_ (.Y(_09002_),
    .A(_08941_));
 sg13g2_a221oi_1 _14737_ (.B2(_09002_),
    .C1(net1014),
    .B1(_09001_),
    .A1(_08985_),
    .Y(_09003_),
    .A2(_08990_));
 sg13g2_a21o_1 _14738_ (.A2(_08983_),
    .A1(net956),
    .B1(_09003_),
    .X(_09004_));
 sg13g2_nand2_1 _14739_ (.Y(_09005_),
    .A(_08848_),
    .B(net1035));
 sg13g2_nand2_1 _14740_ (.Y(_09006_),
    .A(net965),
    .B(net1012));
 sg13g2_nor3_1 _14741_ (.A(net962),
    .B(_09005_),
    .C(_09006_),
    .Y(_09007_));
 sg13g2_nor2_1 _14742_ (.A(net1001),
    .B(_09007_),
    .Y(_09008_));
 sg13g2_nor2_1 _14743_ (.A(_08891_),
    .B(net966),
    .Y(_09009_));
 sg13g2_nor2_1 _14744_ (.A(net968),
    .B(_08912_),
    .Y(_09010_));
 sg13g2_nor2_1 _14745_ (.A(net1008),
    .B(net1037),
    .Y(_09011_));
 sg13g2_nand2_1 _14746_ (.Y(_09012_),
    .A(net934),
    .B(_09011_));
 sg13g2_o21ai_1 _14747_ (.B1(_09012_),
    .Y(_09013_),
    .A1(net967),
    .A2(_08905_));
 sg13g2_a22oi_1 _14748_ (.Y(_09014_),
    .B1(_09010_),
    .B2(_09013_),
    .A2(_08926_),
    .A1(_09009_));
 sg13g2_buf_1 _14749_ (.A(net1033),
    .X(_09015_));
 sg13g2_xor2_1 _14750_ (.B(net1007),
    .A(net959),
    .X(_09016_));
 sg13g2_nor4_1 _14751_ (.A(net929),
    .B(net998),
    .C(net931),
    .D(_09016_),
    .Y(_09017_));
 sg13g2_nor2_1 _14752_ (.A(net1015),
    .B(_09017_),
    .Y(_09018_));
 sg13g2_o21ai_1 _14753_ (.B1(_08926_),
    .Y(_09019_),
    .A1(_08918_),
    .A2(_08971_));
 sg13g2_a221oi_1 _14754_ (.B2(_09019_),
    .C1(net1014),
    .B1(_09018_),
    .A1(_09008_),
    .Y(_09020_),
    .A2(_09014_));
 sg13g2_nand2_1 _14755_ (.Y(_09021_),
    .A(_09009_),
    .B(_08926_));
 sg13g2_nand2b_1 _14756_ (.Y(_09022_),
    .B(net1034),
    .A_N(net1054));
 sg13g2_buf_1 _14757_ (.A(_09022_),
    .X(_09023_));
 sg13g2_a21oi_1 _14758_ (.A1(_09021_),
    .A2(_09023_),
    .Y(_09024_),
    .B1(net902));
 sg13g2_buf_1 _14759_ (.A(net1009),
    .X(_09025_));
 sg13g2_buf_1 _14760_ (.A(_09025_),
    .X(_09026_));
 sg13g2_nand2_1 _14761_ (.Y(_09027_),
    .A(net1038),
    .B(_08869_));
 sg13g2_buf_2 _14762_ (.A(_09027_),
    .X(_09028_));
 sg13g2_nand2_1 _14763_ (.Y(_09029_),
    .A(net1008),
    .B(net1011));
 sg13g2_a21oi_1 _14764_ (.A1(net926),
    .A2(_09028_),
    .Y(_09030_),
    .B1(_09029_));
 sg13g2_o21ai_1 _14765_ (.B1(net969),
    .Y(_09031_),
    .A1(_09024_),
    .A2(_09030_));
 sg13g2_nor2_1 _14766_ (.A(net1003),
    .B(_09031_),
    .Y(_09032_));
 sg13g2_nor3_1 _14767_ (.A(_08967_),
    .B(_09020_),
    .C(_09032_),
    .Y(_09033_));
 sg13g2_a21oi_1 _14768_ (.A1(net1000),
    .A2(_09004_),
    .Y(_09034_),
    .B1(_09033_));
 sg13g2_mux2_1 _14769_ (.A0(_09034_),
    .A1(_08818_),
    .S(net882),
    .X(_00364_));
 sg13g2_a22oi_1 _14770_ (.Y(_09035_),
    .B1(_08993_),
    .B2(_08880_),
    .A2(_08977_),
    .A1(_08991_));
 sg13g2_inv_1 _14771_ (.Y(_09036_),
    .A(_00178_));
 sg13g2_nand3_1 _14772_ (.B(_09036_),
    .C(_08928_),
    .A(_08895_),
    .Y(_09037_));
 sg13g2_o21ai_1 _14773_ (.B1(_09037_),
    .Y(_09038_),
    .A1(_08841_),
    .A2(_09035_));
 sg13g2_nor2_1 _14774_ (.A(net1009),
    .B(_08835_),
    .Y(_09039_));
 sg13g2_buf_1 _14775_ (.A(_08940_),
    .X(_09040_));
 sg13g2_nand2_1 _14776_ (.Y(_09041_),
    .A(net1002),
    .B(net1008));
 sg13g2_nor2_1 _14777_ (.A(net965),
    .B(_09041_),
    .Y(_09042_));
 sg13g2_inv_1 _14778_ (.Y(_09043_),
    .A(_09042_));
 sg13g2_a21oi_1 _14779_ (.A1(_08920_),
    .A2(_09043_),
    .Y(_09044_),
    .B1(net931));
 sg13g2_nor2_1 _14780_ (.A(net998),
    .B(_09006_),
    .Y(_09045_));
 sg13g2_a22oi_1 _14781_ (.Y(_09046_),
    .B1(_09045_),
    .B2(_08942_),
    .A2(_09044_),
    .A1(net925));
 sg13g2_nor2b_1 _14782_ (.A(_08877_),
    .B_N(_08855_),
    .Y(_09047_));
 sg13g2_buf_1 _14783_ (.A(_09047_),
    .X(_09048_));
 sg13g2_nand4_1 _14784_ (.B(_00178_),
    .C(_08977_),
    .A(_08895_),
    .Y(_09049_),
    .D(_09048_));
 sg13g2_o21ai_1 _14785_ (.B1(_09049_),
    .Y(_09050_),
    .A1(net1014),
    .A2(_09046_));
 sg13g2_a221oi_1 _14786_ (.B2(_08954_),
    .C1(_08833_),
    .B1(_09050_),
    .A1(_09038_),
    .Y(_09051_),
    .A2(_09039_));
 sg13g2_nand2_1 _14787_ (.Y(_09052_),
    .A(_08852_),
    .B(net1054));
 sg13g2_buf_1 _14788_ (.A(_09052_),
    .X(_09053_));
 sg13g2_nand2_1 _14789_ (.Y(_09054_),
    .A(_09023_),
    .B(_09053_));
 sg13g2_nor3_1 _14790_ (.A(net938),
    .B(net1039),
    .C(_08998_),
    .Y(_09055_));
 sg13g2_nor3_1 _14791_ (.A(_08913_),
    .B(_09036_),
    .C(_08962_),
    .Y(_09056_));
 sg13g2_a22oi_1 _14792_ (.Y(_09057_),
    .B1(_09056_),
    .B2(net935),
    .A2(_09055_),
    .A1(_09054_));
 sg13g2_nor2_1 _14793_ (.A(net1039),
    .B(net999),
    .Y(_09058_));
 sg13g2_nor2_1 _14794_ (.A(net1034),
    .B(net1035),
    .Y(_09059_));
 sg13g2_buf_2 _14795_ (.A(_09059_),
    .X(_09060_));
 sg13g2_nand3_1 _14796_ (.B(_09058_),
    .C(_09060_),
    .A(_08871_),
    .Y(_09061_));
 sg13g2_o21ai_1 _14797_ (.B1(_09061_),
    .Y(_09062_),
    .A1(_08938_),
    .A2(_09057_));
 sg13g2_nor2_1 _14798_ (.A(net1000),
    .B(_09062_),
    .Y(_09063_));
 sg13g2_nor3_1 _14799_ (.A(net881),
    .B(_09051_),
    .C(_09063_),
    .Y(_09064_));
 sg13g2_a21o_1 _14800_ (.A2(net882),
    .A1(\top_ihp.oisc.micro_op[11] ),
    .B1(_09064_),
    .X(_00365_));
 sg13g2_buf_1 _14801_ (.A(\top_ihp.oisc.micro_op[12] ),
    .X(_09065_));
 sg13g2_inv_1 _14802_ (.Y(_09066_),
    .A(_09065_));
 sg13g2_and2_1 _14803_ (.A(_08840_),
    .B(_08961_),
    .X(_09067_));
 sg13g2_buf_1 _14804_ (.A(_09067_),
    .X(_09068_));
 sg13g2_o21ai_1 _14805_ (.B1(_08887_),
    .Y(_09069_),
    .A1(_08899_),
    .A2(net937));
 sg13g2_buf_1 _14806_ (.A(net934),
    .X(_09070_));
 sg13g2_nand2_1 _14807_ (.Y(_09071_),
    .A(net1036),
    .B(net1011));
 sg13g2_buf_1 _14808_ (.A(_09071_),
    .X(_09072_));
 sg13g2_a21oi_1 _14809_ (.A1(net931),
    .A2(_09072_),
    .Y(_09073_),
    .B1(net967));
 sg13g2_a221oi_1 _14810_ (.B2(net901),
    .C1(_09073_),
    .B1(_09069_),
    .A1(_08926_),
    .Y(_09074_),
    .A2(_08987_));
 sg13g2_and2_1 _14811_ (.A(net1034),
    .B(net1035),
    .X(_09075_));
 sg13g2_buf_1 _14812_ (.A(_09075_),
    .X(_09076_));
 sg13g2_or2_1 _14813_ (.X(_09077_),
    .B(net1035),
    .A(net1034));
 sg13g2_buf_1 _14814_ (.A(_09077_),
    .X(_09078_));
 sg13g2_o21ai_1 _14815_ (.B1(_09078_),
    .Y(_09079_),
    .A1(_09070_),
    .A2(_09076_));
 sg13g2_nand3_1 _14816_ (.B(net925),
    .C(_09079_),
    .A(net938),
    .Y(_09080_));
 sg13g2_o21ai_1 _14817_ (.B1(_09080_),
    .Y(_09081_),
    .A1(net938),
    .A2(_09074_));
 sg13g2_buf_1 _14818_ (.A(net1006),
    .X(_09082_));
 sg13g2_a22oi_1 _14819_ (.Y(_09083_),
    .B1(net936),
    .B2(_08977_),
    .A2(_09025_),
    .A1(net954));
 sg13g2_nand2_1 _14820_ (.Y(_09084_),
    .A(net1010),
    .B(net1009));
 sg13g2_o21ai_1 _14821_ (.B1(_09084_),
    .Y(_09085_),
    .A1(_08902_),
    .A2(_09078_));
 sg13g2_nand2_1 _14822_ (.Y(_09086_),
    .A(net964),
    .B(net1007));
 sg13g2_o21ai_1 _14823_ (.B1(_09086_),
    .Y(_09087_),
    .A1(_08899_),
    .A2(_08874_));
 sg13g2_a22oi_1 _14824_ (.Y(_09088_),
    .B1(_09087_),
    .B2(_08977_),
    .A2(_09085_),
    .A1(_08890_));
 sg13g2_o21ai_1 _14825_ (.B1(_09088_),
    .Y(_09089_),
    .A1(net967),
    .A2(_09083_));
 sg13g2_nor2_1 _14826_ (.A(net1012),
    .B(net1035),
    .Y(_09090_));
 sg13g2_buf_2 _14827_ (.A(_09090_),
    .X(_09091_));
 sg13g2_nor2_1 _14828_ (.A(_09091_),
    .B(_09048_),
    .Y(_09092_));
 sg13g2_buf_2 _14829_ (.A(_00181_),
    .X(_09093_));
 sg13g2_nand2_1 _14830_ (.Y(_09094_),
    .A(_08869_),
    .B(_09093_));
 sg13g2_o21ai_1 _14831_ (.B1(net960),
    .Y(_09095_),
    .A1(net964),
    .A2(_09094_));
 sg13g2_a21oi_1 _14832_ (.A1(_08871_),
    .A2(_09092_),
    .Y(_09096_),
    .B1(_09095_));
 sg13g2_nor2_1 _14833_ (.A(net934),
    .B(_09023_),
    .Y(_09097_));
 sg13g2_nor2_1 _14834_ (.A(net1006),
    .B(_09053_),
    .Y(_09098_));
 sg13g2_buf_1 _14835_ (.A(net959),
    .X(_09099_));
 sg13g2_o21ai_1 _14836_ (.B1(_09099_),
    .Y(_09100_),
    .A1(_09097_),
    .A2(_09098_));
 sg13g2_nor2_1 _14837_ (.A(net1008),
    .B(_08848_),
    .Y(_09101_));
 sg13g2_nand2_1 _14838_ (.Y(_09102_),
    .A(_08844_),
    .B(_09101_));
 sg13g2_nor2_1 _14839_ (.A(net1012),
    .B(net1013),
    .Y(_09103_));
 sg13g2_o21ai_1 _14840_ (.B1(_08902_),
    .Y(_09104_),
    .A1(_08919_),
    .A2(_09103_));
 sg13g2_a21oi_1 _14841_ (.A1(_09102_),
    .A2(_09104_),
    .Y(_09105_),
    .B1(net955));
 sg13g2_buf_1 _14842_ (.A(_00182_),
    .X(_09106_));
 sg13g2_nor2b_1 _14843_ (.A(_08867_),
    .B_N(_08872_),
    .Y(_09107_));
 sg13g2_buf_2 _14844_ (.A(_09107_),
    .X(_09108_));
 sg13g2_a21o_1 _14845_ (.A2(_09108_),
    .A1(_09106_),
    .B1(_08940_),
    .X(_09109_));
 sg13g2_nor3_1 _14846_ (.A(_09042_),
    .B(_09105_),
    .C(_09109_),
    .Y(_09110_));
 sg13g2_a21oi_1 _14847_ (.A1(_09096_),
    .A2(_09100_),
    .Y(_09111_),
    .B1(_09110_));
 sg13g2_mux2_1 _14848_ (.A0(_09089_),
    .A1(_09111_),
    .S(net1015),
    .X(_09112_));
 sg13g2_a22oi_1 _14849_ (.Y(_09113_),
    .B1(_09112_),
    .B2(net1003),
    .A2(_09081_),
    .A1(_09068_));
 sg13g2_a22oi_1 _14850_ (.Y(_09114_),
    .B1(_08879_),
    .B2(_08979_),
    .A2(net927),
    .A1(net932));
 sg13g2_nor2_1 _14851_ (.A(net954),
    .B(_09114_),
    .Y(_09115_));
 sg13g2_a21oi_1 _14852_ (.A1(net927),
    .A2(_08919_),
    .Y(_09116_),
    .B1(_09115_));
 sg13g2_nand2b_1 _14853_ (.Y(_09117_),
    .B(net1053),
    .A_N(net1054));
 sg13g2_buf_2 _14854_ (.A(_09117_),
    .X(_09118_));
 sg13g2_o21ai_1 _14855_ (.B1(_09118_),
    .Y(_09119_),
    .A1(net1004),
    .A2(_08941_));
 sg13g2_nor2_1 _14856_ (.A(_09042_),
    .B(_09119_),
    .Y(_09120_));
 sg13g2_nor2_2 _14857_ (.A(_08869_),
    .B(net1011),
    .Y(_09121_));
 sg13g2_o21ai_1 _14858_ (.B1(net928),
    .Y(_09122_),
    .A1(net967),
    .A2(_09121_));
 sg13g2_a21oi_1 _14859_ (.A1(_09120_),
    .A2(_09122_),
    .Y(_09123_),
    .B1(net1015));
 sg13g2_a21oi_1 _14860_ (.A1(net1015),
    .A2(_09116_),
    .Y(_09124_),
    .B1(_09123_));
 sg13g2_nor2_1 _14861_ (.A(net1036),
    .B(net1053),
    .Y(_09125_));
 sg13g2_nand3_1 _14862_ (.B(_08863_),
    .C(_09029_),
    .A(net961),
    .Y(_09126_));
 sg13g2_o21ai_1 _14863_ (.B1(_09126_),
    .Y(_09127_),
    .A1(net954),
    .A2(_08863_));
 sg13g2_a22oi_1 _14864_ (.Y(_09128_),
    .B1(_09127_),
    .B2(net902),
    .A2(_09125_),
    .A1(_09106_));
 sg13g2_o21ai_1 _14865_ (.B1(_09008_),
    .Y(_09129_),
    .A1(net926),
    .A2(_09128_));
 sg13g2_nand2_1 _14866_ (.Y(_09130_),
    .A(net1036),
    .B(net1054));
 sg13g2_buf_2 _14867_ (.A(_09130_),
    .X(_09131_));
 sg13g2_and2_1 _14868_ (.A(net1010),
    .B(_09131_),
    .X(_09132_));
 sg13g2_nor2_2 _14869_ (.A(_08936_),
    .B(_08873_),
    .Y(_09133_));
 sg13g2_o21ai_1 _14870_ (.B1(net1004),
    .Y(_09134_),
    .A1(_09132_),
    .A2(_09133_));
 sg13g2_o21ai_1 _14871_ (.B1(_09134_),
    .Y(_09135_),
    .A1(_09072_),
    .A2(_09010_));
 sg13g2_nor2_2 _14872_ (.A(net1008),
    .B(_08884_),
    .Y(_09136_));
 sg13g2_a221oi_1 _14873_ (.B2(net936),
    .C1(_08837_),
    .B1(_09136_),
    .A1(net903),
    .Y(_09137_),
    .A2(_09135_));
 sg13g2_nor2_1 _14874_ (.A(net1005),
    .B(_09137_),
    .Y(_09138_));
 sg13g2_a221oi_1 _14875_ (.B2(_09138_),
    .C1(_08833_),
    .B1(_09129_),
    .A1(net956),
    .Y(_09139_),
    .A2(_09124_));
 sg13g2_a21oi_1 _14876_ (.A1(net1040),
    .A2(_09113_),
    .Y(_09140_),
    .B1(_09139_));
 sg13g2_nor2_1 _14877_ (.A(net881),
    .B(_09140_),
    .Y(_09141_));
 sg13g2_a21oi_1 _14878_ (.A1(_09066_),
    .A2(net882),
    .Y(_00366_),
    .B1(_09141_));
 sg13g2_nand2_1 _14879_ (.Y(_09142_),
    .A(_08836_),
    .B(_08839_));
 sg13g2_nor2_1 _14880_ (.A(net928),
    .B(_09023_),
    .Y(_09143_));
 sg13g2_a21oi_1 _14881_ (.A1(net902),
    .A2(_09048_),
    .Y(_09144_),
    .B1(_09143_));
 sg13g2_nor2_1 _14882_ (.A(net966),
    .B(_09005_),
    .Y(_09145_));
 sg13g2_o21ai_1 _14883_ (.B1(_08845_),
    .Y(_09146_),
    .A1(_09097_),
    .A2(_09145_));
 sg13g2_o21ai_1 _14884_ (.B1(_09146_),
    .Y(_09147_),
    .A1(_09091_),
    .A2(_09028_));
 sg13g2_nand2_1 _14885_ (.Y(_09148_),
    .A(net925),
    .B(_09147_));
 sg13g2_o21ai_1 _14886_ (.B1(_09148_),
    .Y(_09149_),
    .A1(_08905_),
    .A2(_09144_));
 sg13g2_nor2b_1 _14887_ (.A(_08851_),
    .B_N(_08843_),
    .Y(_09150_));
 sg13g2_buf_1 _14888_ (.A(_09150_),
    .X(_09151_));
 sg13g2_a21oi_1 _14889_ (.A1(net961),
    .A2(_09048_),
    .Y(_09152_),
    .B1(_09091_));
 sg13g2_and2_1 _14890_ (.A(net934),
    .B(_09076_),
    .X(_09153_));
 sg13g2_nor3_1 _14891_ (.A(net932),
    .B(_09060_),
    .C(_09153_),
    .Y(_09154_));
 sg13g2_a21oi_1 _14892_ (.A1(net928),
    .A2(_09152_),
    .Y(_09155_),
    .B1(_09154_));
 sg13g2_a221oi_1 _14893_ (.B2(net925),
    .C1(net1005),
    .B1(_09155_),
    .A1(_08958_),
    .Y(_09156_),
    .A2(_09151_));
 sg13g2_nand2_2 _14894_ (.Y(_09157_),
    .A(net937),
    .B(_09118_));
 sg13g2_nor2_1 _14895_ (.A(_09151_),
    .B(_09157_),
    .Y(_09158_));
 sg13g2_a22oi_1 _14896_ (.Y(_09159_),
    .B1(_09158_),
    .B2(net998),
    .A2(_09157_),
    .A1(_09045_));
 sg13g2_nor3_1 _14897_ (.A(_08912_),
    .B(_08879_),
    .C(net999),
    .Y(_09160_));
 sg13g2_nor2_1 _14898_ (.A(_08839_),
    .B(_09160_),
    .Y(_09161_));
 sg13g2_o21ai_1 _14899_ (.B1(net1002),
    .Y(_09162_),
    .A1(net1010),
    .A2(_08847_));
 sg13g2_a22oi_1 _14900_ (.Y(_09163_),
    .B1(_09076_),
    .B2(_09162_),
    .A2(_09060_),
    .A1(net965));
 sg13g2_nand2b_1 _14901_ (.Y(_09164_),
    .B(_08985_),
    .A_N(_09163_));
 sg13g2_and2_1 _14902_ (.A(_09161_),
    .B(_09164_),
    .X(_09165_));
 sg13g2_a21o_1 _14903_ (.A2(_09159_),
    .A1(net1005),
    .B1(_09165_),
    .X(_09166_));
 sg13g2_o21ai_1 _14904_ (.B1(_09166_),
    .Y(_09167_),
    .A1(net958),
    .A2(_09156_));
 sg13g2_o21ai_1 _14905_ (.B1(_09167_),
    .Y(_09168_),
    .A1(_09142_),
    .A2(_09149_));
 sg13g2_buf_1 _14906_ (.A(net962),
    .X(_09169_));
 sg13g2_nor2b_1 _14907_ (.A(_08999_),
    .B_N(net926),
    .Y(_09170_));
 sg13g2_nor4_1 _14908_ (.A(_09169_),
    .B(_08962_),
    .C(_09044_),
    .D(_09170_),
    .Y(_09171_));
 sg13g2_nor3_1 _14909_ (.A(net1033),
    .B(net964),
    .C(_08970_),
    .Y(_09172_));
 sg13g2_a21oi_1 _14910_ (.A1(net955),
    .A2(_09106_),
    .Y(_09173_),
    .B1(_09172_));
 sg13g2_nand2_1 _14911_ (.Y(_09174_),
    .A(net959),
    .B(_09133_));
 sg13g2_a21o_1 _14912_ (.A2(_09174_),
    .A1(_09131_),
    .B1(_08887_),
    .X(_09175_));
 sg13g2_o21ai_1 _14913_ (.B1(_09175_),
    .Y(_09176_),
    .A1(net923),
    .A2(_09173_));
 sg13g2_a22oi_1 _14914_ (.Y(_09177_),
    .B1(_08991_),
    .B2(_08946_),
    .A2(net960),
    .A1(net1033));
 sg13g2_nor2b_1 _14915_ (.A(_09177_),
    .B_N(net955),
    .Y(_09178_));
 sg13g2_nor2b_1 _14916_ (.A(_08842_),
    .B_N(_08851_),
    .Y(_09179_));
 sg13g2_buf_1 _14917_ (.A(_09179_),
    .X(_09180_));
 sg13g2_o21ai_1 _14918_ (.B1(net961),
    .Y(_09181_),
    .A1(net1007),
    .A2(net997));
 sg13g2_nor2_1 _14919_ (.A(net931),
    .B(_09181_),
    .Y(_09182_));
 sg13g2_nand3_1 _14920_ (.B(_08863_),
    .C(_09029_),
    .A(net934),
    .Y(_09183_));
 sg13g2_a21oi_1 _14921_ (.A1(_09053_),
    .A2(_09183_),
    .Y(_09184_),
    .B1(net924));
 sg13g2_nor4_1 _14922_ (.A(net1001),
    .B(_09178_),
    .C(_09182_),
    .D(_09184_),
    .Y(_09185_));
 sg13g2_a21oi_1 _14923_ (.A1(net958),
    .A2(_09176_),
    .Y(_09186_),
    .B1(_09185_));
 sg13g2_nor2_1 _14924_ (.A(net956),
    .B(_09186_),
    .Y(_09187_));
 sg13g2_o21ai_1 _14925_ (.B1(net1040),
    .Y(_09188_),
    .A1(_09171_),
    .A2(_09187_));
 sg13g2_o21ai_1 _14926_ (.B1(_09188_),
    .Y(_09189_),
    .A1(net1040),
    .A2(_09168_));
 sg13g2_mux2_1 _14927_ (.A0(_09189_),
    .A1(\top_ihp.oisc.micro_op[13] ),
    .S(_08965_),
    .X(_00367_));
 sg13g2_nor2_1 _14928_ (.A(_08848_),
    .B(_08858_),
    .Y(_09190_));
 sg13g2_nand2_1 _14929_ (.Y(_09191_),
    .A(net966),
    .B(_09190_));
 sg13g2_nand2_1 _14930_ (.Y(_09192_),
    .A(_09012_),
    .B(_09191_));
 sg13g2_a22oi_1 _14931_ (.Y(_09193_),
    .B1(_09192_),
    .B2(net928),
    .A2(_09190_),
    .A1(net935));
 sg13g2_a21oi_1 _14932_ (.A1(_08946_),
    .A2(_08994_),
    .Y(_09194_),
    .B1(net997));
 sg13g2_nor2_1 _14933_ (.A(net901),
    .B(_09194_),
    .Y(_09195_));
 sg13g2_a21oi_1 _14934_ (.A1(_08887_),
    .A2(_09012_),
    .Y(_09196_),
    .B1(net924));
 sg13g2_nor3_1 _14935_ (.A(net931),
    .B(_09195_),
    .C(_09196_),
    .Y(_09197_));
 sg13g2_a21oi_1 _14936_ (.A1(net926),
    .A2(_09193_),
    .Y(_09198_),
    .B1(_09197_));
 sg13g2_a21o_1 _14937_ (.A2(_09041_),
    .A1(net932),
    .B1(_09098_),
    .X(_09199_));
 sg13g2_o21ai_1 _14938_ (.B1(_09028_),
    .Y(_09200_),
    .A1(net924),
    .A2(_09072_));
 sg13g2_a22oi_1 _14939_ (.Y(_09201_),
    .B1(_09200_),
    .B2(_09091_),
    .A2(_09199_),
    .A1(net923));
 sg13g2_nor2_1 _14940_ (.A(_08837_),
    .B(_09201_),
    .Y(_09202_));
 sg13g2_a21oi_1 _14941_ (.A1(net969),
    .A2(_09198_),
    .Y(_09203_),
    .B1(_09202_));
 sg13g2_nand2_1 _14942_ (.Y(_09204_),
    .A(_08891_),
    .B(_08860_));
 sg13g2_nand2_1 _14943_ (.Y(_09205_),
    .A(_08882_),
    .B(net960));
 sg13g2_nor2_1 _14944_ (.A(net961),
    .B(_09205_),
    .Y(_09206_));
 sg13g2_a21o_1 _14945_ (.A2(_09204_),
    .A1(net928),
    .B1(_09206_),
    .X(_09207_));
 sg13g2_nand3_1 _14946_ (.B(net1013),
    .C(_08875_),
    .A(net933),
    .Y(_09208_));
 sg13g2_a21oi_1 _14947_ (.A1(_09021_),
    .A2(_09208_),
    .Y(_09209_),
    .B1(net902));
 sg13g2_a221oi_1 _14948_ (.B2(net903),
    .C1(_09209_),
    .B1(_09207_),
    .A1(_08926_),
    .Y(_09210_),
    .A2(_09136_));
 sg13g2_nand2b_1 _14949_ (.Y(_09211_),
    .B(_09068_),
    .A_N(_09210_));
 sg13g2_o21ai_1 _14950_ (.B1(_09211_),
    .Y(_09212_),
    .A1(net956),
    .A2(_09203_));
 sg13g2_and2_1 _14951_ (.A(_08842_),
    .B(_08851_),
    .X(_09213_));
 sg13g2_buf_2 _14952_ (.A(_09213_),
    .X(_09214_));
 sg13g2_xnor2_1 _14953_ (.Y(_09215_),
    .A(net1002),
    .B(net1037));
 sg13g2_nand2b_1 _14954_ (.Y(_09216_),
    .B(net955),
    .A_N(_09215_));
 sg13g2_o21ai_1 _14955_ (.B1(_09216_),
    .Y(_09217_),
    .A1(net998),
    .A2(_09205_));
 sg13g2_o21ai_1 _14956_ (.B1(_09131_),
    .Y(_09218_),
    .A1(net930),
    .A2(_09118_));
 sg13g2_a22oi_1 _14957_ (.Y(_09219_),
    .B1(_09218_),
    .B2(net935),
    .A2(_09217_),
    .A1(_09214_));
 sg13g2_xnor2_1 _14958_ (.Y(_09220_),
    .A(net1006),
    .B(net964));
 sg13g2_nand2_1 _14959_ (.Y(_09221_),
    .A(_08937_),
    .B(_09214_));
 sg13g2_o21ai_1 _14960_ (.B1(_09221_),
    .Y(_09222_),
    .A1(_08970_),
    .A2(_09220_));
 sg13g2_a22oi_1 _14961_ (.Y(_09223_),
    .B1(_09222_),
    .B2(_09040_),
    .A2(_08999_),
    .A1(_08942_));
 sg13g2_a22oi_1 _14962_ (.Y(_09224_),
    .B1(_09220_),
    .B2(net924),
    .A2(_09076_),
    .A1(_08915_));
 sg13g2_inv_1 _14963_ (.Y(_09225_),
    .A(_09224_));
 sg13g2_a22oi_1 _14964_ (.Y(_09226_),
    .B1(_09225_),
    .B2(net923),
    .A2(_09060_),
    .A1(_08977_));
 sg13g2_nor2_1 _14965_ (.A(net961),
    .B(_09023_),
    .Y(_09227_));
 sg13g2_o21ai_1 _14966_ (.B1(_08909_),
    .Y(_09228_),
    .A1(_09145_),
    .A2(_09227_));
 sg13g2_o21ai_1 _14967_ (.B1(_08994_),
    .Y(_09229_),
    .A1(_08988_),
    .A2(_09133_));
 sg13g2_and2_1 _14968_ (.A(_09228_),
    .B(_09229_),
    .X(_09230_));
 sg13g2_mux4_1 _14969_ (.S0(net1005),
    .A0(_09219_),
    .A1(_09223_),
    .A2(_09226_),
    .A3(_09230_),
    .S1(net969),
    .X(_09231_));
 sg13g2_nor2_1 _14970_ (.A(net1040),
    .B(_09231_),
    .Y(_09232_));
 sg13g2_a21oi_1 _14971_ (.A1(net1040),
    .A2(_09212_),
    .Y(_09233_),
    .B1(_09232_));
 sg13g2_nand2_1 _14972_ (.Y(_09234_),
    .A(\top_ihp.oisc.micro_op[14] ),
    .B(net881));
 sg13g2_o21ai_1 _14973_ (.B1(_09234_),
    .Y(_00368_),
    .A1(net882),
    .A2(_09233_));
 sg13g2_nand2_1 _14974_ (.Y(_09235_),
    .A(net933),
    .B(_08907_));
 sg13g2_a21o_1 _14975_ (.A2(_09235_),
    .A1(_09053_),
    .B1(net968),
    .X(_09236_));
 sg13g2_nor2_1 _14976_ (.A(_08903_),
    .B(_09054_),
    .Y(_09237_));
 sg13g2_nor2_1 _14977_ (.A(_09108_),
    .B(_09237_),
    .Y(_09238_));
 sg13g2_a21oi_1 _14978_ (.A1(_09236_),
    .A2(_09238_),
    .Y(_09239_),
    .B1(_09109_));
 sg13g2_nor3_1 _14979_ (.A(net928),
    .B(_08958_),
    .C(_09108_),
    .Y(_09240_));
 sg13g2_nor3_1 _14980_ (.A(_09029_),
    .B(_09132_),
    .C(_09240_),
    .Y(_09241_));
 sg13g2_o21ai_1 _14981_ (.B1(_08961_),
    .Y(_09242_),
    .A1(_09239_),
    .A2(_09241_));
 sg13g2_a21o_1 _14982_ (.A2(_08970_),
    .A1(_08907_),
    .B1(_09082_),
    .X(_09243_));
 sg13g2_a22oi_1 _14983_ (.Y(_09244_),
    .B1(_09243_),
    .B2(net957),
    .A2(_09108_),
    .A1(_09093_));
 sg13g2_nor3_1 _14984_ (.A(_09082_),
    .B(_08923_),
    .C(net1001),
    .Y(_09245_));
 sg13g2_nor2_1 _14985_ (.A(net1032),
    .B(_09002_),
    .Y(_09246_));
 sg13g2_a22oi_1 _14986_ (.Y(_09247_),
    .B1(_09246_),
    .B2(_09121_),
    .A2(_09133_),
    .A1(_08985_));
 sg13g2_nor2_1 _14987_ (.A(net938),
    .B(_09247_),
    .Y(_09248_));
 sg13g2_a21oi_1 _14988_ (.A1(_09085_),
    .A2(_09245_),
    .Y(_09249_),
    .B1(_09248_));
 sg13g2_o21ai_1 _14989_ (.B1(_09249_),
    .Y(_09250_),
    .A1(net999),
    .A2(_09244_));
 sg13g2_nor2_1 _14990_ (.A(net956),
    .B(_09250_),
    .Y(_09251_));
 sg13g2_a21oi_1 _14991_ (.A1(net956),
    .A2(_09242_),
    .Y(_09252_),
    .B1(_09251_));
 sg13g2_nand2_1 _14992_ (.Y(_09253_),
    .A(_09093_),
    .B(_09108_));
 sg13g2_o21ai_1 _14993_ (.B1(_09253_),
    .Y(_09254_),
    .A1(net957),
    .A2(_09108_));
 sg13g2_nand3_1 _14994_ (.B(_08986_),
    .C(_09131_),
    .A(_08865_),
    .Y(_09255_));
 sg13g2_o21ai_1 _14995_ (.B1(_09255_),
    .Y(_09256_),
    .A1(net965),
    .A2(_09131_));
 sg13g2_a22oi_1 _14996_ (.Y(_09257_),
    .B1(_09256_),
    .B2(net933),
    .A2(net935),
    .A1(_08907_));
 sg13g2_nor2_1 _14997_ (.A(net960),
    .B(_09257_),
    .Y(_09258_));
 sg13g2_a21oi_1 _14998_ (.A1(net925),
    .A2(_09254_),
    .Y(_09259_),
    .B1(_09258_));
 sg13g2_nand2_1 _14999_ (.Y(_09260_),
    .A(_08863_),
    .B(_09072_));
 sg13g2_a22oi_1 _15000_ (.Y(_09261_),
    .B1(_09260_),
    .B2(net968),
    .A2(_09011_),
    .A1(net954));
 sg13g2_nor2_1 _15001_ (.A(net965),
    .B(_09125_),
    .Y(_09262_));
 sg13g2_a21oi_1 _15002_ (.A1(net932),
    .A2(_09215_),
    .Y(_09263_),
    .B1(_09262_));
 sg13g2_a22oi_1 _15003_ (.Y(_09264_),
    .B1(_09263_),
    .B2(net929),
    .A2(_09121_),
    .A1(_09093_));
 sg13g2_mux2_1 _15004_ (.A0(_09261_),
    .A1(_09264_),
    .S(net931),
    .X(_09265_));
 sg13g2_a21oi_1 _15005_ (.A1(_08863_),
    .A2(net957),
    .Y(_09266_),
    .B1(net961));
 sg13g2_a21o_1 _15006_ (.A2(_09011_),
    .A1(_08871_),
    .B1(_09266_),
    .X(_09267_));
 sg13g2_o21ai_1 _15007_ (.B1(_08879_),
    .Y(_09268_),
    .A1(_08993_),
    .A2(_09121_));
 sg13g2_nand3_1 _15008_ (.B(_08908_),
    .C(_09106_),
    .A(net901),
    .Y(_09269_));
 sg13g2_nand3_1 _15009_ (.B(_09268_),
    .C(_09269_),
    .A(net931),
    .Y(_09270_));
 sg13g2_o21ai_1 _15010_ (.B1(_09270_),
    .Y(_09271_),
    .A1(net926),
    .A2(_09267_));
 sg13g2_nor3_1 _15011_ (.A(net929),
    .B(_09005_),
    .C(_09016_),
    .Y(_09272_));
 sg13g2_nand2b_1 _15012_ (.Y(_09273_),
    .B(net1038),
    .A_N(net1009));
 sg13g2_buf_1 _15013_ (.A(_09273_),
    .X(_09274_));
 sg13g2_a21oi_1 _15014_ (.A1(net930),
    .A2(_08887_),
    .Y(_09275_),
    .B1(_09274_));
 sg13g2_nor2_1 _15015_ (.A(_09272_),
    .B(_09275_),
    .Y(_09276_));
 sg13g2_mux4_1 _15016_ (.S0(net1003),
    .A0(_09259_),
    .A1(_09265_),
    .A2(_09271_),
    .A3(_09276_),
    .S1(net969),
    .X(_09277_));
 sg13g2_nand2_1 _15017_ (.Y(_09278_),
    .A(net1000),
    .B(_09277_));
 sg13g2_o21ai_1 _15018_ (.B1(_09278_),
    .Y(_09279_),
    .A1(net1000),
    .A2(_09252_));
 sg13g2_buf_1 _15019_ (.A(\top_ihp.oisc.micro_op[15] ),
    .X(_09280_));
 sg13g2_nand2_1 _15020_ (.Y(_09281_),
    .A(_09280_),
    .B(net881));
 sg13g2_o21ai_1 _15021_ (.B1(_09281_),
    .Y(_00369_),
    .A1(net882),
    .A2(_09279_));
 sg13g2_a22oi_1 _15022_ (.Y(_09282_),
    .B1(_08993_),
    .B2(_09237_),
    .A2(_09151_),
    .A1(_08942_));
 sg13g2_o21ai_1 _15023_ (.B1(_09072_),
    .Y(_09283_),
    .A1(_08881_),
    .A2(_09118_));
 sg13g2_a22oi_1 _15024_ (.Y(_09284_),
    .B1(_09283_),
    .B2(net924),
    .A2(net963),
    .A1(net927));
 sg13g2_inv_1 _15025_ (.Y(_09285_),
    .A(_09284_));
 sg13g2_a221oi_1 _15026_ (.B2(net903),
    .C1(net1005),
    .B1(_09285_),
    .A1(net936),
    .Y(_09286_),
    .A2(net935));
 sg13g2_a21oi_1 _15027_ (.A1(net1014),
    .A2(_09282_),
    .Y(_09287_),
    .B1(_09286_));
 sg13g2_o21ai_1 _15028_ (.B1(net967),
    .Y(_09288_),
    .A1(_08941_),
    .A2(net999));
 sg13g2_a21oi_1 _15029_ (.A1(_08871_),
    .A2(_09288_),
    .Y(_09289_),
    .B1(_08977_));
 sg13g2_a221oi_1 _15030_ (.B2(net929),
    .C1(_09289_),
    .B1(net937),
    .A1(net962),
    .Y(_09290_),
    .A2(_08941_));
 sg13g2_nor2_1 _15031_ (.A(_08881_),
    .B(_09157_),
    .Y(_09291_));
 sg13g2_a22oi_1 _15032_ (.Y(_09292_),
    .B1(_09291_),
    .B2(net928),
    .A2(_09157_),
    .A1(net963));
 sg13g2_nor3_1 _15033_ (.A(net903),
    .B(net1003),
    .C(_09292_),
    .Y(_09293_));
 sg13g2_a21oi_1 _15034_ (.A1(net1003),
    .A2(_09290_),
    .Y(_09294_),
    .B1(_09293_));
 sg13g2_nor2_1 _15035_ (.A(net969),
    .B(_09294_),
    .Y(_09295_));
 sg13g2_a21oi_1 _15036_ (.A1(_08838_),
    .A2(_09287_),
    .Y(_09296_),
    .B1(_09295_));
 sg13g2_a21oi_1 _15037_ (.A1(_08849_),
    .A2(_09180_),
    .Y(_09297_),
    .B1(_08889_));
 sg13g2_nand2_1 _15038_ (.Y(_09298_),
    .A(net1037),
    .B(_08989_));
 sg13g2_a21oi_1 _15039_ (.A1(net963),
    .A2(_09091_),
    .Y(_09299_),
    .B1(_09298_));
 sg13g2_nor3_1 _15040_ (.A(_09142_),
    .B(_09297_),
    .C(_09299_),
    .Y(_09300_));
 sg13g2_o21ai_1 _15041_ (.B1(net1002),
    .Y(_09301_),
    .A1(_08853_),
    .A2(_08847_));
 sg13g2_a21oi_1 _15042_ (.A1(_09102_),
    .A2(_09301_),
    .Y(_09302_),
    .B1(net955));
 sg13g2_a21oi_1 _15043_ (.A1(_08986_),
    .A2(_08972_),
    .Y(_09303_),
    .B1(_09302_));
 sg13g2_nand2_1 _15044_ (.Y(_09304_),
    .A(net934),
    .B(net960));
 sg13g2_nand3_1 _15045_ (.B(_09304_),
    .C(net997),
    .A(_08958_),
    .Y(_09305_));
 sg13g2_o21ai_1 _15046_ (.B1(_09305_),
    .Y(_09306_),
    .A1(net923),
    .A2(_09303_));
 sg13g2_nor2_2 _15047_ (.A(_09151_),
    .B(net997),
    .Y(_09307_));
 sg13g2_nand2_1 _15048_ (.Y(_09308_),
    .A(net1002),
    .B(_09307_));
 sg13g2_o21ai_1 _15049_ (.B1(_09308_),
    .Y(_09309_),
    .A1(net1006),
    .A2(_09093_));
 sg13g2_nor2_1 _15050_ (.A(net955),
    .B(_09309_),
    .Y(_09310_));
 sg13g2_nor3_1 _15051_ (.A(net960),
    .B(_09153_),
    .C(_09310_),
    .Y(_09311_));
 sg13g2_xnor2_1 _15052_ (.Y(_09312_),
    .A(_08898_),
    .B(net1033));
 sg13g2_nor2_1 _15053_ (.A(_09084_),
    .B(_09312_),
    .Y(_09313_));
 sg13g2_nand2_1 _15054_ (.Y(_09314_),
    .A(_08885_),
    .B(_08847_));
 sg13g2_a21oi_1 _15055_ (.A1(net964),
    .A2(_09314_),
    .Y(_09315_),
    .B1(net932));
 sg13g2_nor4_1 _15056_ (.A(net962),
    .B(_09133_),
    .C(_09313_),
    .D(_09315_),
    .Y(_09316_));
 sg13g2_nor3_1 _15057_ (.A(net1001),
    .B(_09311_),
    .C(_09316_),
    .Y(_09317_));
 sg13g2_a21oi_1 _15058_ (.A1(net958),
    .A2(_09306_),
    .Y(_09318_),
    .B1(_09317_));
 sg13g2_nor2_1 _15059_ (.A(_08841_),
    .B(_09318_),
    .Y(_09319_));
 sg13g2_o21ai_1 _15060_ (.B1(_08834_),
    .Y(_09320_),
    .A1(_09300_),
    .A2(_09319_));
 sg13g2_o21ai_1 _15061_ (.B1(_09320_),
    .Y(_09321_),
    .A1(_08834_),
    .A2(_09296_));
 sg13g2_mux2_1 _15062_ (.A0(_09321_),
    .A1(_07962_),
    .S(net881),
    .X(_00370_));
 sg13g2_a22oi_1 _15063_ (.Y(_09322_),
    .B1(_08979_),
    .B2(net929),
    .A2(net935),
    .A1(net927));
 sg13g2_o21ai_1 _15064_ (.B1(net937),
    .Y(_09323_),
    .A1(_08928_),
    .A2(_09136_));
 sg13g2_o21ai_1 _15065_ (.B1(_09323_),
    .Y(_09324_),
    .A1(net930),
    .A2(_09322_));
 sg13g2_o21ai_1 _15066_ (.B1(_09070_),
    .Y(_09325_),
    .A1(_08942_),
    .A2(_08975_));
 sg13g2_or4_1 _15067_ (.A(net924),
    .B(_08923_),
    .C(_08907_),
    .D(_09108_),
    .X(_09326_));
 sg13g2_o21ai_1 _15068_ (.B1(_09326_),
    .Y(_09327_),
    .A1(net938),
    .A2(_09325_));
 sg13g2_nor2_2 _15069_ (.A(net1012),
    .B(_08835_),
    .Y(_09328_));
 sg13g2_a22oi_1 _15070_ (.Y(_09329_),
    .B1(_09327_),
    .B2(_09328_),
    .A2(_09324_),
    .A1(net958));
 sg13g2_a22oi_1 _15071_ (.Y(_09330_),
    .B1(_09328_),
    .B2(_08958_),
    .A2(_09098_),
    .A1(net1032));
 sg13g2_nand2b_1 _15072_ (.Y(_09331_),
    .B(net902),
    .A_N(_09330_));
 sg13g2_nor2_1 _15073_ (.A(_08835_),
    .B(_09005_),
    .Y(_09332_));
 sg13g2_nor2_1 _15074_ (.A(_08873_),
    .B(_08836_),
    .Y(_09333_));
 sg13g2_o21ai_1 _15075_ (.B1(net935),
    .Y(_09334_),
    .A1(_09332_),
    .A2(_09333_));
 sg13g2_nand3_1 _15076_ (.B(_09331_),
    .C(_09334_),
    .A(net923),
    .Y(_09335_));
 sg13g2_a22oi_1 _15077_ (.Y(_09336_),
    .B1(net997),
    .B2(_08883_),
    .A2(_09060_),
    .A1(_08977_));
 sg13g2_o21ai_1 _15078_ (.B1(_09308_),
    .Y(_09337_),
    .A1(net1013),
    .A2(_09307_));
 sg13g2_nand2_1 _15079_ (.Y(_09338_),
    .A(_09026_),
    .B(_09337_));
 sg13g2_nor4_1 _15080_ (.A(net932),
    .B(net955),
    .C(_08918_),
    .D(_08919_),
    .Y(_09339_));
 sg13g2_nor2_1 _15081_ (.A(net1004),
    .B(net1032),
    .Y(_09340_));
 sg13g2_nor2b_1 _15082_ (.A(_09339_),
    .B_N(_09340_),
    .Y(_09341_));
 sg13g2_a22oi_1 _15083_ (.Y(_09342_),
    .B1(_09338_),
    .B2(_09341_),
    .A2(_09336_),
    .A1(_08985_));
 sg13g2_a21oi_1 _15084_ (.A1(_09335_),
    .A2(_09342_),
    .Y(_09343_),
    .B1(net956));
 sg13g2_a21oi_1 _15085_ (.A1(_08969_),
    .A2(_09329_),
    .Y(_09344_),
    .B1(_09343_));
 sg13g2_o21ai_1 _15086_ (.B1(net937),
    .Y(_09345_),
    .A1(net901),
    .A2(_09118_));
 sg13g2_a22oi_1 _15087_ (.Y(_09346_),
    .B1(_09345_),
    .B2(net903),
    .A2(_09009_),
    .A1(net936));
 sg13g2_a21oi_1 _15088_ (.A1(_08938_),
    .A2(_08926_),
    .Y(_09347_),
    .B1(_09206_));
 sg13g2_nand2_1 _15089_ (.Y(_09348_),
    .A(_09151_),
    .B(_09347_));
 sg13g2_o21ai_1 _15090_ (.B1(_09348_),
    .Y(_09349_),
    .A1(net902),
    .A2(_09346_));
 sg13g2_nor2_1 _15091_ (.A(_08952_),
    .B(_08839_),
    .Y(_09350_));
 sg13g2_nor2_1 _15092_ (.A(net1010),
    .B(_08941_),
    .Y(_09351_));
 sg13g2_a22oi_1 _15093_ (.Y(_09352_),
    .B1(_09351_),
    .B2(_08994_),
    .A2(_09214_),
    .A1(_08944_));
 sg13g2_nand3_1 _15094_ (.B(_08874_),
    .C(_09307_),
    .A(net1033),
    .Y(_09353_));
 sg13g2_o21ai_1 _15095_ (.B1(_09353_),
    .Y(_09354_),
    .A1(net1006),
    .A2(_09352_));
 sg13g2_nand3_1 _15096_ (.B(_08934_),
    .C(_09354_),
    .A(_08952_),
    .Y(_09355_));
 sg13g2_nand2b_1 _15097_ (.Y(_09356_),
    .B(_09355_),
    .A_N(_09300_));
 sg13g2_a21oi_1 _15098_ (.A1(_09349_),
    .A2(_09350_),
    .Y(_09357_),
    .B1(_09356_));
 sg13g2_nor2_1 _15099_ (.A(_08968_),
    .B(_09357_),
    .Y(_09358_));
 sg13g2_a21oi_1 _15100_ (.A1(net1000),
    .A2(_09344_),
    .Y(_09359_),
    .B1(_09358_));
 sg13g2_nand2_1 _15101_ (.Y(_09360_),
    .A(_07967_),
    .B(_08965_));
 sg13g2_o21ai_1 _15102_ (.B1(_09360_),
    .Y(_00371_),
    .A1(_08832_),
    .A2(_09359_));
 sg13g2_inv_1 _15103_ (.Y(_09361_),
    .A(_07964_));
 sg13g2_nand3_1 _15104_ (.B(net963),
    .C(_09060_),
    .A(net1032),
    .Y(_09362_));
 sg13g2_and3_1 _15105_ (.X(_09363_),
    .A(_09002_),
    .B(_08993_),
    .C(net997));
 sg13g2_inv_1 _15106_ (.Y(_09364_),
    .A(_09363_));
 sg13g2_a221oi_1 _15107_ (.B2(net963),
    .C1(net1032),
    .B1(_09060_),
    .A1(_09214_),
    .Y(_09365_),
    .A2(_08883_));
 sg13g2_a221oi_1 _15108_ (.B2(_08985_),
    .C1(_09365_),
    .B1(_09364_),
    .A1(net962),
    .Y(_09366_),
    .A2(_09362_));
 sg13g2_nor3_1 _15109_ (.A(_09028_),
    .B(net999),
    .C(_09053_),
    .Y(_09367_));
 sg13g2_o21ai_1 _15110_ (.B1(_08935_),
    .Y(_09368_),
    .A1(_09366_),
    .A2(_09367_));
 sg13g2_nor2_1 _15111_ (.A(net1001),
    .B(_09364_),
    .Y(_09369_));
 sg13g2_and3_1 _15112_ (.X(_09370_),
    .A(net1001),
    .B(_08945_),
    .C(_09045_));
 sg13g2_o21ai_1 _15113_ (.B1(net1014),
    .Y(_09371_),
    .A1(_09369_),
    .A2(_09370_));
 sg13g2_nand4_1 _15114_ (.B(_08915_),
    .C(_08985_),
    .A(net1014),
    .Y(_09372_),
    .D(_09048_));
 sg13g2_nand3_1 _15115_ (.B(_09371_),
    .C(_09372_),
    .A(_09368_),
    .Y(_09373_));
 sg13g2_a22oi_1 _15116_ (.Y(_09374_),
    .B1(_08979_),
    .B2(net954),
    .A2(_08975_),
    .A1(_09015_));
 sg13g2_nand3_1 _15117_ (.B(_08875_),
    .C(_08880_),
    .A(net901),
    .Y(_09375_));
 sg13g2_o21ai_1 _15118_ (.B1(_09375_),
    .Y(_09376_),
    .A1(_09307_),
    .A2(_09374_));
 sg13g2_a21o_1 _15119_ (.A2(_09376_),
    .A1(_09350_),
    .B1(_09356_),
    .X(_09377_));
 sg13g2_a21o_1 _15120_ (.A2(_09377_),
    .A1(_08833_),
    .B1(_08831_),
    .X(_09378_));
 sg13g2_a21oi_1 _15121_ (.A1(net1000),
    .A2(_09373_),
    .Y(_09379_),
    .B1(_09378_));
 sg13g2_a21oi_1 _15122_ (.A1(_09361_),
    .A2(_08829_),
    .Y(_00372_),
    .B1(_09379_));
 sg13g2_inv_1 _15123_ (.Y(_09380_),
    .A(_07968_));
 sg13g2_and2_1 _15124_ (.A(net1009),
    .B(_08835_),
    .X(_09381_));
 sg13g2_buf_1 _15125_ (.A(_09381_),
    .X(_09382_));
 sg13g2_nor2_1 _15126_ (.A(_08898_),
    .B(_09028_),
    .Y(_09383_));
 sg13g2_a22oi_1 _15127_ (.Y(_09384_),
    .B1(_09382_),
    .B2(_08919_),
    .A2(_09039_),
    .A1(_08918_));
 sg13g2_nor2_1 _15128_ (.A(net924),
    .B(_09384_),
    .Y(_09385_));
 sg13g2_a21oi_1 _15129_ (.A1(_09382_),
    .A2(_09383_),
    .Y(_09386_),
    .B1(_09385_));
 sg13g2_nor2_1 _15130_ (.A(net925),
    .B(_09386_),
    .Y(_09387_));
 sg13g2_o21ai_1 _15131_ (.B1(_08935_),
    .Y(_09388_),
    .A1(_09366_),
    .A2(_09387_));
 sg13g2_or4_1 _15132_ (.A(net925),
    .B(_09028_),
    .C(_09078_),
    .D(_09142_),
    .X(_09389_));
 sg13g2_nand3_1 _15133_ (.B(_09388_),
    .C(_09389_),
    .A(_09371_),
    .Y(_09390_));
 sg13g2_a21oi_1 _15134_ (.A1(net1000),
    .A2(_09390_),
    .Y(_09391_),
    .B1(_09378_));
 sg13g2_a21oi_1 _15135_ (.A1(_09380_),
    .A2(_08832_),
    .Y(_00373_),
    .B1(_09391_));
 sg13g2_inv_1 _15136_ (.Y(_09392_),
    .A(_07969_));
 sg13g2_nand2b_1 _15137_ (.Y(_09393_),
    .B(net1000),
    .A_N(_09372_));
 sg13g2_a22oi_1 _15138_ (.Y(_00374_),
    .B1(_09391_),
    .B2(_09393_),
    .A2(_08829_),
    .A1(_09392_));
 sg13g2_nor2_1 _15139_ (.A(net1002),
    .B(_09190_),
    .Y(_09394_));
 sg13g2_a21oi_1 _15140_ (.A1(_08865_),
    .A2(_09125_),
    .Y(_09395_),
    .B1(_09121_));
 sg13g2_o21ai_1 _15141_ (.B1(_09395_),
    .Y(_09396_),
    .A1(net965),
    .A2(_09394_));
 sg13g2_a22oi_1 _15142_ (.Y(_09397_),
    .B1(_09396_),
    .B2(net933),
    .A2(_09136_),
    .A1(_08905_));
 sg13g2_a22oi_1 _15143_ (.Y(_09398_),
    .B1(_08993_),
    .B2(_08885_),
    .A2(net1037),
    .A1(_08869_));
 sg13g2_nand3_1 _15144_ (.B(net1037),
    .C(_08879_),
    .A(net1013),
    .Y(_09399_));
 sg13g2_o21ai_1 _15145_ (.B1(_09399_),
    .Y(_09400_),
    .A1(_08844_),
    .A2(_09398_));
 sg13g2_a22oi_1 _15146_ (.Y(_09401_),
    .B1(_09400_),
    .B2(net955),
    .A2(_09383_),
    .A1(_09190_));
 sg13g2_o21ai_1 _15147_ (.B1(_09401_),
    .Y(_09402_),
    .A1(net931),
    .A2(_09397_));
 sg13g2_nor2_1 _15148_ (.A(_08944_),
    .B(_08979_),
    .Y(_09403_));
 sg13g2_nand2_1 _15149_ (.Y(_09404_),
    .A(_08986_),
    .B(_09072_));
 sg13g2_a221oi_1 _15150_ (.B2(net959),
    .C1(net967),
    .B1(_09404_),
    .A1(net934),
    .Y(_09405_),
    .A2(_09403_));
 sg13g2_a221oi_1 _15151_ (.B2(net1006),
    .C1(net933),
    .B1(_09403_),
    .A1(_08944_),
    .Y(_09406_),
    .A2(net963));
 sg13g2_o21ai_1 _15152_ (.B1(net1039),
    .Y(_09407_),
    .A1(_09405_),
    .A2(_09406_));
 sg13g2_o21ai_1 _15153_ (.B1(_09407_),
    .Y(_09408_),
    .A1(net1039),
    .A2(_09402_));
 sg13g2_o21ai_1 _15154_ (.B1(net930),
    .Y(_09409_),
    .A1(_08939_),
    .A2(net962));
 sg13g2_a21oi_1 _15155_ (.A1(_09010_),
    .A2(_09409_),
    .Y(_09410_),
    .B1(net1039));
 sg13g2_o21ai_1 _15156_ (.B1(_08937_),
    .Y(_09411_),
    .A1(net1004),
    .A2(_08956_));
 sg13g2_nor2_1 _15157_ (.A(_08879_),
    .B(_08890_),
    .Y(_09412_));
 sg13g2_a22oi_1 _15158_ (.Y(_09413_),
    .B1(_09412_),
    .B2(_09221_),
    .A2(_09411_),
    .A1(_08849_));
 sg13g2_nor3_1 _15159_ (.A(net1004),
    .B(net957),
    .C(_08883_),
    .Y(_09414_));
 sg13g2_a21o_1 _15160_ (.A2(_09084_),
    .A1(_08994_),
    .B1(_09414_),
    .X(_09415_));
 sg13g2_a221oi_1 _15161_ (.B2(net901),
    .C1(_09142_),
    .B1(_09415_),
    .A1(net926),
    .Y(_09416_),
    .A2(_09413_));
 sg13g2_a221oi_1 _15162_ (.B2(_09008_),
    .C1(_09416_),
    .B1(_09410_),
    .A1(net958),
    .Y(_09417_),
    .A2(_09408_));
 sg13g2_nor2_1 _15163_ (.A(_08833_),
    .B(_09417_),
    .Y(_09418_));
 sg13g2_o21ai_1 _15164_ (.B1(_09304_),
    .Y(_09419_),
    .A1(net998),
    .A2(_09086_));
 sg13g2_nor3_1 _15165_ (.A(net924),
    .B(net962),
    .C(_08907_),
    .Y(_09420_));
 sg13g2_a21oi_1 _15166_ (.A1(net902),
    .A2(_09419_),
    .Y(_09421_),
    .B1(_09420_));
 sg13g2_nand2_1 _15167_ (.Y(_09422_),
    .A(net901),
    .B(net927));
 sg13g2_nand3_1 _15168_ (.B(_09204_),
    .C(_09422_),
    .A(_09214_),
    .Y(_09423_));
 sg13g2_o21ai_1 _15169_ (.B1(_09423_),
    .Y(_09424_),
    .A1(net903),
    .A2(_09421_));
 sg13g2_a21oi_1 _15170_ (.A1(_09078_),
    .A2(_09314_),
    .Y(_09425_),
    .B1(net959));
 sg13g2_a21oi_1 _15171_ (.A1(_09274_),
    .A2(_09131_),
    .Y(_09426_),
    .B1(net967));
 sg13g2_a21oi_1 _15172_ (.A1(net964),
    .A2(_09101_),
    .Y(_09427_),
    .B1(_08958_));
 sg13g2_nor2_1 _15173_ (.A(net968),
    .B(_09427_),
    .Y(_09428_));
 sg13g2_nor3_1 _15174_ (.A(_09425_),
    .B(_09426_),
    .C(_09428_),
    .Y(_09429_));
 sg13g2_a21o_1 _15175_ (.A2(_09093_),
    .A1(net964),
    .B1(_09091_),
    .X(_09430_));
 sg13g2_nand3_1 _15176_ (.B(_08921_),
    .C(_09274_),
    .A(net1004),
    .Y(_09431_));
 sg13g2_a21oi_1 _15177_ (.A1(net954),
    .A2(_09430_),
    .Y(_09432_),
    .B1(_09431_));
 sg13g2_a21oi_1 _15178_ (.A1(net960),
    .A2(_09429_),
    .Y(_09433_),
    .B1(_09432_));
 sg13g2_nor2_1 _15179_ (.A(net961),
    .B(_09086_),
    .Y(_09434_));
 sg13g2_a221oi_1 _15180_ (.B2(net1033),
    .C1(net965),
    .B1(_08979_),
    .A1(net1002),
    .Y(_09435_),
    .A2(_08944_));
 sg13g2_a21oi_1 _15181_ (.A1(net959),
    .A2(_09157_),
    .Y(_09436_),
    .B1(_09435_));
 sg13g2_nor3_1 _15182_ (.A(net967),
    .B(_09434_),
    .C(_09436_),
    .Y(_09437_));
 sg13g2_o21ai_1 _15183_ (.B1(net937),
    .Y(_09438_),
    .A1(net1013),
    .A2(_09118_));
 sg13g2_nor2_1 _15184_ (.A(net959),
    .B(net1013),
    .Y(_09439_));
 sg13g2_a221oi_1 _15185_ (.B2(net936),
    .C1(net929),
    .B1(_09439_),
    .A1(net932),
    .Y(_09440_),
    .A2(_09438_));
 sg13g2_nor3_1 _15186_ (.A(net1015),
    .B(_09437_),
    .C(_09440_),
    .Y(_09441_));
 sg13g2_a21o_1 _15187_ (.A2(_09433_),
    .A1(net1015),
    .B1(_09441_),
    .X(_09442_));
 sg13g2_a221oi_1 _15188_ (.B2(net1003),
    .C1(_08967_),
    .B1(_09442_),
    .A1(_09068_),
    .Y(_09443_),
    .A2(_09424_));
 sg13g2_or2_1 _15189_ (.X(_09444_),
    .B(_09443_),
    .A(_09418_));
 sg13g2_nand2_1 _15190_ (.Y(_09445_),
    .A(_08814_),
    .B(net881));
 sg13g2_o21ai_1 _15191_ (.B1(_09445_),
    .Y(_00375_),
    .A1(net882),
    .A2(_09444_));
 sg13g2_nand2_1 _15192_ (.Y(_09446_),
    .A(_08844_),
    .B(_09048_));
 sg13g2_o21ai_1 _15193_ (.B1(_09446_),
    .Y(_09447_),
    .A1(net968),
    .A2(_09054_));
 sg13g2_a22oi_1 _15194_ (.Y(_09448_),
    .B1(_09447_),
    .B2(net1004),
    .A2(net936),
    .A1(net933));
 sg13g2_a221oi_1 _15195_ (.B2(net997),
    .C1(net954),
    .B1(_08979_),
    .A1(net932),
    .Y(_09449_),
    .A2(net927));
 sg13g2_a21oi_1 _15196_ (.A1(net930),
    .A2(_09448_),
    .Y(_09450_),
    .B1(_09449_));
 sg13g2_a21oi_1 _15197_ (.A1(net927),
    .A2(_08999_),
    .Y(_09451_),
    .B1(_09450_));
 sg13g2_a21oi_1 _15198_ (.A1(net1004),
    .A2(_09093_),
    .Y(_09452_),
    .B1(_08916_));
 sg13g2_a21o_1 _15199_ (.A2(_09078_),
    .A1(net957),
    .B1(_09215_),
    .X(_09453_));
 sg13g2_o21ai_1 _15200_ (.B1(_09453_),
    .Y(_09454_),
    .A1(_09131_),
    .A2(_09452_));
 sg13g2_a21oi_1 _15201_ (.A1(net936),
    .A2(_08918_),
    .Y(_09455_),
    .B1(_09454_));
 sg13g2_mux2_1 _15202_ (.A0(_09451_),
    .A1(_09455_),
    .S(net1015),
    .X(_09456_));
 sg13g2_a21oi_1 _15203_ (.A1(_09131_),
    .A2(_09235_),
    .Y(_09457_),
    .B1(_08947_));
 sg13g2_nand2_1 _15204_ (.Y(_09458_),
    .A(net968),
    .B(_08958_));
 sg13g2_a21oi_1 _15205_ (.A1(_09255_),
    .A2(_09458_),
    .Y(_09459_),
    .B1(_08939_));
 sg13g2_or3_1 _15206_ (.A(net923),
    .B(_09457_),
    .C(_09459_),
    .X(_09460_));
 sg13g2_nand3_1 _15207_ (.B(_09298_),
    .C(_09460_),
    .A(_09068_),
    .Y(_09461_));
 sg13g2_o21ai_1 _15208_ (.B1(_09461_),
    .Y(_09462_),
    .A1(net956),
    .A2(_09456_));
 sg13g2_a21oi_1 _15209_ (.A1(net1032),
    .A2(_08918_),
    .Y(_09463_),
    .B1(_08981_));
 sg13g2_nand2b_1 _15210_ (.Y(_09464_),
    .B(_09328_),
    .A_N(_08884_));
 sg13g2_o21ai_1 _15211_ (.B1(_09464_),
    .Y(_09465_),
    .A1(_09099_),
    .A2(_09463_));
 sg13g2_nor2_1 _15212_ (.A(net933),
    .B(_08836_),
    .Y(_09466_));
 sg13g2_nor4_1 _15213_ (.A(_09015_),
    .B(_09274_),
    .C(_09328_),
    .D(_09466_),
    .Y(_09467_));
 sg13g2_a21o_1 _15214_ (.A2(_09465_),
    .A1(net926),
    .B1(_09467_),
    .X(_09468_));
 sg13g2_a22oi_1 _15215_ (.Y(_09469_),
    .B1(_09382_),
    .B2(net954),
    .A2(_08836_),
    .A1(net998));
 sg13g2_nand2b_1 _15216_ (.Y(_09470_),
    .B(_09307_),
    .A_N(_09469_));
 sg13g2_a21oi_1 _15217_ (.A1(_08888_),
    .A2(_09333_),
    .Y(_09471_),
    .B1(_09332_));
 sg13g2_nor2b_1 _15218_ (.A(_09471_),
    .B_N(net997),
    .Y(_09472_));
 sg13g2_a21oi_1 _15219_ (.A1(_09136_),
    .A2(_09333_),
    .Y(_09473_),
    .B1(_09472_));
 sg13g2_a21oi_1 _15220_ (.A1(_09470_),
    .A2(_09473_),
    .Y(_09474_),
    .B1(net923));
 sg13g2_a21oi_1 _15221_ (.A1(net923),
    .A2(_09468_),
    .Y(_09475_),
    .B1(_09474_));
 sg13g2_a21oi_1 _15222_ (.A1(net938),
    .A2(_08979_),
    .Y(_09476_),
    .B1(_08909_));
 sg13g2_nor4_1 _15223_ (.A(net903),
    .B(net998),
    .C(net958),
    .D(_09476_),
    .Y(_09477_));
 sg13g2_a21oi_1 _15224_ (.A1(_08954_),
    .A2(_09363_),
    .Y(_09478_),
    .B1(_09477_));
 sg13g2_nor2_1 _15225_ (.A(net929),
    .B(net999),
    .Y(_09479_));
 sg13g2_a21oi_1 _15226_ (.A1(_09091_),
    .A2(_09340_),
    .Y(_09480_),
    .B1(_09479_));
 sg13g2_nor2_1 _15227_ (.A(_09028_),
    .B(_09480_),
    .Y(_09481_));
 sg13g2_nor2b_1 _15228_ (.A(_09481_),
    .B_N(_09161_),
    .Y(_09482_));
 sg13g2_a221oi_1 _15229_ (.B2(_09482_),
    .C1(_08833_),
    .B1(_09478_),
    .A1(_08969_),
    .Y(_09483_),
    .A2(_09475_));
 sg13g2_a21oi_1 _15230_ (.A1(net1040),
    .A2(_09462_),
    .Y(_09484_),
    .B1(_09483_));
 sg13g2_nand2_1 _15231_ (.Y(_09485_),
    .A(_08810_),
    .B(net881));
 sg13g2_o21ai_1 _15232_ (.B1(_09485_),
    .Y(_00376_),
    .A1(net882),
    .A2(_09484_));
 sg13g2_and2_1 _15233_ (.A(_07966_),
    .B(_07971_),
    .X(_09486_));
 sg13g2_buf_8 _15234_ (.A(_09486_),
    .X(_09487_));
 sg13g2_nand2_2 _15235_ (.Y(_09488_),
    .A(_07959_),
    .B(\top_ihp.oisc.micro_state[2] ));
 sg13g2_nand2_1 _15236_ (.Y(_09489_),
    .A(_00086_),
    .B(_09488_));
 sg13g2_buf_1 _15237_ (.A(net1108),
    .X(_09490_));
 sg13g2_o21ai_1 _15238_ (.B1(_09490_),
    .Y(_09491_),
    .A1(_09487_),
    .A2(_09489_));
 sg13g2_buf_2 _15239_ (.A(_09491_),
    .X(_09492_));
 sg13g2_buf_1 _15240_ (.A(_09492_),
    .X(_09493_));
 sg13g2_buf_2 _15241_ (.A(\top_ihp.oisc.state[3] ),
    .X(_09494_));
 sg13g2_buf_1 _15242_ (.A(_09494_),
    .X(_09495_));
 sg13g2_inv_1 _15243_ (.Y(_09496_),
    .A(_07963_));
 sg13g2_buf_8 _15244_ (.A(\top_ihp.oisc.op_a[31] ),
    .X(_09497_));
 sg13g2_buf_2 _15245_ (.A(\top_ihp.oisc.op_b[31] ),
    .X(_09498_));
 sg13g2_nand2b_1 _15246_ (.Y(_09499_),
    .B(_09498_),
    .A_N(_09497_));
 sg13g2_nand2b_1 _15247_ (.Y(_09500_),
    .B(_08226_),
    .A_N(_08227_));
 sg13g2_nand2b_1 _15248_ (.Y(_09501_),
    .B(_08095_),
    .A_N(_08092_));
 sg13g2_xor2_1 _15249_ (.B(_08087_),
    .A(_08086_),
    .X(_09502_));
 sg13g2_xor2_1 _15250_ (.B(_09497_),
    .A(_09498_),
    .X(_09503_));
 sg13g2_xor2_1 _15251_ (.B(_08306_),
    .A(_08312_),
    .X(_09504_));
 sg13g2_nor4_1 _15252_ (.A(_09501_),
    .B(_09502_),
    .C(_09503_),
    .D(_09504_),
    .Y(_09505_));
 sg13g2_nor2_1 _15253_ (.A(_08079_),
    .B(_08080_),
    .Y(_09506_));
 sg13g2_xor2_1 _15254_ (.B(_08082_),
    .A(_08081_),
    .X(_09507_));
 sg13g2_nor3_1 _15255_ (.A(_09506_),
    .B(_08089_),
    .C(_09507_),
    .Y(_09508_));
 sg13g2_nand3_1 _15256_ (.B(_09505_),
    .C(_09508_),
    .A(_08323_),
    .Y(_09509_));
 sg13g2_nor2_1 _15257_ (.A(_09500_),
    .B(_09509_),
    .Y(_09510_));
 sg13g2_nand4_1 _15258_ (.B(_08250_),
    .C(_08287_),
    .A(_08132_),
    .Y(_09511_),
    .D(_09510_));
 sg13g2_and3_1 _15259_ (.X(_09512_),
    .A(_08311_),
    .B(_09499_),
    .C(_09511_));
 sg13g2_and3_1 _15260_ (.X(_09513_),
    .A(_08312_),
    .B(_09499_),
    .C(_09511_));
 sg13g2_o21ai_1 _15261_ (.B1(_08351_),
    .Y(_09514_),
    .A1(_09512_),
    .A2(_09513_));
 sg13g2_nor2b_1 _15262_ (.A(_09498_),
    .B_N(_09497_),
    .Y(_09515_));
 sg13g2_a21oi_1 _15263_ (.A1(_08316_),
    .A2(_09499_),
    .Y(_09516_),
    .B1(_09515_));
 sg13g2_nand3_1 _15264_ (.B(_09514_),
    .C(_09516_),
    .A(_09496_),
    .Y(_09517_));
 sg13g2_nor3_1 _15265_ (.A(_09494_),
    .B(net922),
    .C(_09488_),
    .Y(_09518_));
 sg13g2_buf_1 _15266_ (.A(_09518_),
    .X(_09519_));
 sg13g2_and2_1 _15267_ (.A(net938),
    .B(_09519_),
    .X(_09520_));
 sg13g2_a22oi_1 _15268_ (.Y(_09521_),
    .B1(_09517_),
    .B2(_09520_),
    .A2(\top_ihp.oisc.decoder.decoded[0] ),
    .A1(net1031));
 sg13g2_nor2b_1 _15269_ (.A(_09517_),
    .B_N(_09519_),
    .Y(_09522_));
 sg13g2_o21ai_1 _15270_ (.B1(_08904_),
    .Y(_09523_),
    .A1(_09492_),
    .A2(_09522_));
 sg13g2_o21ai_1 _15271_ (.B1(_09523_),
    .Y(_00377_),
    .A1(_09493_),
    .A2(_09521_));
 sg13g2_nand3b_1 _15272_ (.B(_07963_),
    .C(_08904_),
    .Y(_09524_),
    .A_N(_07962_));
 sg13g2_o21ai_1 _15273_ (.B1(_07962_),
    .Y(_09525_),
    .A1(_09496_),
    .A2(_08846_));
 sg13g2_nand2_1 _15274_ (.Y(_09526_),
    .A(_09514_),
    .B(_09516_));
 sg13g2_buf_2 _15275_ (.A(_09526_),
    .X(_09527_));
 sg13g2_mux2_1 _15276_ (.A0(_09525_),
    .A1(_08846_),
    .S(_09527_),
    .X(_09528_));
 sg13g2_nand3b_1 _15277_ (.B(net890),
    .C(_08854_),
    .Y(_09529_),
    .A_N(_09492_));
 sg13g2_a21oi_1 _15278_ (.A1(_09524_),
    .A2(_09528_),
    .Y(_09530_),
    .B1(_09529_));
 sg13g2_nand4_1 _15279_ (.B(net890),
    .C(_09524_),
    .A(_08900_),
    .Y(_09531_),
    .D(_09528_));
 sg13g2_inv_2 _15280_ (.Y(_09532_),
    .A(_09494_));
 sg13g2_inv_1 _15281_ (.Y(_09533_),
    .A(\top_ihp.oisc.decoder.decoded[1] ));
 sg13g2_nor3_1 _15282_ (.A(_09532_),
    .B(_09533_),
    .C(_09492_),
    .Y(_09534_));
 sg13g2_a21oi_1 _15283_ (.A1(_08900_),
    .A2(_09492_),
    .Y(_09535_),
    .B1(_09534_));
 sg13g2_nand3b_1 _15284_ (.B(_09531_),
    .C(_09535_),
    .Y(_00378_),
    .A_N(_09530_));
 sg13g2_a21o_1 _15285_ (.A2(_08842_),
    .A1(_07963_),
    .B1(_08851_),
    .X(_09536_));
 sg13g2_a22oi_1 _15286_ (.Y(_09537_),
    .B1(_09536_),
    .B2(_07962_),
    .A2(_09214_),
    .A1(_07963_));
 sg13g2_xor2_1 _15287_ (.B(net930),
    .A(_07967_),
    .X(_09538_));
 sg13g2_xnor2_1 _15288_ (.Y(_09539_),
    .A(_09537_),
    .B(_09538_));
 sg13g2_xnor2_1 _15289_ (.Y(_09540_),
    .A(net998),
    .B(_09214_));
 sg13g2_mux2_1 _15290_ (.A0(_09539_),
    .A1(_09540_),
    .S(_09527_),
    .X(_09541_));
 sg13g2_a221oi_1 _15291_ (.B2(_09541_),
    .C1(net880),
    .B1(net890),
    .A1(net1031),
    .Y(_09542_),
    .A2(\top_ihp.oisc.decoder.decoded[2] ));
 sg13g2_a21oi_1 _15292_ (.A1(net901),
    .A2(net880),
    .Y(_00379_),
    .B1(_09542_));
 sg13g2_nand2_1 _15293_ (.Y(_09543_),
    .A(_07967_),
    .B(_08866_));
 sg13g2_nor2_1 _15294_ (.A(_07967_),
    .B(_08867_),
    .Y(_09544_));
 sg13g2_a21oi_1 _15295_ (.A1(_09537_),
    .A2(_09543_),
    .Y(_09545_),
    .B1(_09544_));
 sg13g2_xnor2_1 _15296_ (.Y(_09546_),
    .A(_07964_),
    .B(_09026_));
 sg13g2_xnor2_1 _15297_ (.Y(_09547_),
    .A(_09545_),
    .B(_09546_));
 sg13g2_nor2_1 _15298_ (.A(_09093_),
    .B(_09041_),
    .Y(_09548_));
 sg13g2_xnor2_1 _15299_ (.Y(_09549_),
    .A(_08941_),
    .B(_09548_));
 sg13g2_mux2_1 _15300_ (.A0(_09547_),
    .A1(_09549_),
    .S(_09527_),
    .X(_09550_));
 sg13g2_a22oi_1 _15301_ (.Y(_09551_),
    .B1(net890),
    .B2(_09550_),
    .A2(\top_ihp.oisc.decoder.decoded[3] ),
    .A1(net1031));
 sg13g2_nand2_1 _15302_ (.Y(_09552_),
    .A(net926),
    .B(net880));
 sg13g2_o21ai_1 _15303_ (.B1(_09552_),
    .Y(_00380_),
    .A1(net880),
    .A2(_09551_));
 sg13g2_nor2_1 _15304_ (.A(net1035),
    .B(_09545_),
    .Y(_09553_));
 sg13g2_a21oi_1 _15305_ (.A1(_08872_),
    .A2(_09545_),
    .Y(_09554_),
    .B1(_07964_));
 sg13g2_nor2_1 _15306_ (.A(_09553_),
    .B(_09554_),
    .Y(_09555_));
 sg13g2_xnor2_1 _15307_ (.Y(_09556_),
    .A(_07968_),
    .B(_09169_));
 sg13g2_xnor2_1 _15308_ (.Y(_09557_),
    .A(_09555_),
    .B(_09556_));
 sg13g2_nand2b_1 _15309_ (.Y(_09558_),
    .B(_09076_),
    .A_N(_08884_));
 sg13g2_xnor2_1 _15310_ (.Y(_09559_),
    .A(_09036_),
    .B(_09558_));
 sg13g2_mux2_1 _15311_ (.A0(_09557_),
    .A1(_09559_),
    .S(_09527_),
    .X(_09560_));
 sg13g2_a221oi_1 _15312_ (.B2(_09560_),
    .C1(net880),
    .B1(net890),
    .A1(net1031),
    .Y(_09561_),
    .A2(\top_ihp.oisc.decoder.decoded[4] ));
 sg13g2_a21oi_1 _15313_ (.A1(net925),
    .A2(net880),
    .Y(_00381_),
    .B1(_09561_));
 sg13g2_nor2_1 _15314_ (.A(_08889_),
    .B(_09555_),
    .Y(_09562_));
 sg13g2_a21oi_1 _15315_ (.A1(net1007),
    .A2(_09555_),
    .Y(_09563_),
    .B1(_07968_));
 sg13g2_nor2_2 _15316_ (.A(_09562_),
    .B(_09563_),
    .Y(_09564_));
 sg13g2_nand2_1 _15317_ (.Y(_09565_),
    .A(_07969_),
    .B(_08836_));
 sg13g2_nand2_1 _15318_ (.Y(_09566_),
    .A(_09392_),
    .B(net1032));
 sg13g2_and2_1 _15319_ (.A(_09565_),
    .B(_09566_),
    .X(_09567_));
 sg13g2_xnor2_1 _15320_ (.Y(_09568_),
    .A(_09564_),
    .B(_09567_));
 sg13g2_nor2_1 _15321_ (.A(_09040_),
    .B(_09558_),
    .Y(_09569_));
 sg13g2_xnor2_1 _15322_ (.Y(_09570_),
    .A(_08961_),
    .B(_09569_));
 sg13g2_mux2_1 _15323_ (.A0(_09568_),
    .A1(_09570_),
    .S(_09527_),
    .X(_09571_));
 sg13g2_a221oi_1 _15324_ (.B2(_09571_),
    .C1(_09492_),
    .B1(net890),
    .A1(net1031),
    .Y(_09572_),
    .A2(\top_ihp.oisc.decoder.decoded[5] ));
 sg13g2_a21oi_1 _15325_ (.A1(_08838_),
    .A2(net880),
    .Y(_00382_),
    .B1(_09572_));
 sg13g2_mux2_1 _15326_ (.A0(_09565_),
    .A1(_09566_),
    .S(_09564_),
    .X(_09573_));
 sg13g2_xnor2_1 _15327_ (.Y(_09574_),
    .A(net1014),
    .B(_09573_));
 sg13g2_nor2_1 _15328_ (.A(net999),
    .B(_09558_),
    .Y(_09575_));
 sg13g2_xnor2_1 _15329_ (.Y(_09576_),
    .A(_00176_),
    .B(_09575_));
 sg13g2_mux2_1 _15330_ (.A0(_09574_),
    .A1(_09576_),
    .S(_09527_),
    .X(_09577_));
 sg13g2_a221oi_1 _15331_ (.B2(_09577_),
    .C1(_09492_),
    .B1(net890),
    .A1(net1031),
    .Y(_09578_),
    .A2(\top_ihp.oisc.decoder.decoded[6] ));
 sg13g2_a21oi_1 _15332_ (.A1(net1003),
    .A2(net880),
    .Y(_00383_),
    .B1(_09578_));
 sg13g2_nand2_1 _15333_ (.Y(_09579_),
    .A(_07969_),
    .B(_09350_));
 sg13g2_nand3_1 _15334_ (.B(_08953_),
    .C(_08839_),
    .A(_09392_),
    .Y(_09580_));
 sg13g2_mux2_1 _15335_ (.A0(_09579_),
    .A1(_09580_),
    .S(_09564_),
    .X(_09581_));
 sg13g2_xnor2_1 _15336_ (.Y(_09582_),
    .A(_08833_),
    .B(_09581_));
 sg13g2_nand4_1 _15337_ (.B(net1039),
    .C(_08926_),
    .A(net1001),
    .Y(_09583_),
    .D(_09548_));
 sg13g2_xor2_1 _15338_ (.B(_09583_),
    .A(_00175_),
    .X(_09584_));
 sg13g2_mux2_1 _15339_ (.A0(_09582_),
    .A1(_09584_),
    .S(_09527_),
    .X(_09585_));
 sg13g2_a221oi_1 _15340_ (.B2(_09585_),
    .C1(_09492_),
    .B1(net890),
    .A1(net1031),
    .Y(_09586_),
    .A2(\top_ihp.oisc.decoder.decoded[7] ));
 sg13g2_a21oi_1 _15341_ (.A1(_08968_),
    .A2(_09493_),
    .Y(_00384_),
    .B1(_09586_));
 sg13g2_inv_1 _15342_ (.Y(_09587_),
    .A(\top_ihp.oisc.micro_state[2] ));
 sg13g2_mux2_1 _15343_ (.A0(_09587_),
    .A1(_13599_),
    .S(_07961_),
    .X(_00385_));
 sg13g2_nand2_1 _15344_ (.Y(_09588_),
    .A(\top_ihp.oisc.micro_state[1] ),
    .B(_07961_));
 sg13g2_o21ai_1 _15345_ (.B1(_09588_),
    .Y(_00386_),
    .A1(net922),
    .A2(_08829_));
 sg13g2_nand2_1 _15346_ (.Y(_09589_),
    .A(_07973_),
    .B(net1016));
 sg13g2_o21ai_1 _15347_ (.B1(_09589_),
    .Y(_00387_),
    .A1(net1049),
    .A2(_09587_));
 sg13g2_buf_1 _15348_ (.A(\top_ihp.oisc.state[2] ),
    .X(_09590_));
 sg13g2_nor2_1 _15349_ (.A(net1052),
    .B(_09494_),
    .Y(_09591_));
 sg13g2_buf_1 _15350_ (.A(_09591_),
    .X(_09592_));
 sg13g2_buf_8 _15351_ (.A(_09592_),
    .X(_09593_));
 sg13g2_buf_1 _15352_ (.A(\top_ihp.oisc.state[4] ),
    .X(_09594_));
 sg13g2_inv_2 _15353_ (.Y(_09595_),
    .A(net1051));
 sg13g2_buf_1 _15354_ (.A(_09595_),
    .X(_09596_));
 sg13g2_and2_1 _15355_ (.A(net1058),
    .B(_08823_),
    .X(_09597_));
 sg13g2_buf_1 _15356_ (.A(_09597_),
    .X(_09598_));
 sg13g2_buf_1 _15357_ (.A(_09598_),
    .X(_09599_));
 sg13g2_buf_1 _15358_ (.A(net952),
    .X(_09600_));
 sg13g2_buf_8 _15359_ (.A(\top_ihp.oisc.mem_addr_lowbits[1] ),
    .X(_09601_));
 sg13g2_buf_1 _15360_ (.A(_09601_),
    .X(_09602_));
 sg13g2_and3_1 _15361_ (.X(_09603_),
    .A(_08772_),
    .B(_08363_),
    .C(_08369_));
 sg13g2_buf_8 _15362_ (.A(_09603_),
    .X(_09604_));
 sg13g2_buf_1 _15363_ (.A(_09604_),
    .X(_09605_));
 sg13g2_nand2b_1 _15364_ (.Y(_09606_),
    .B(net900),
    .A_N(_00154_));
 sg13g2_buf_8 _15365_ (.A(_08770_),
    .X(_09607_));
 sg13g2_buf_1 _15366_ (.A(net889),
    .X(_09608_));
 sg13g2_buf_8 _15367_ (.A(_09608_),
    .X(_09609_));
 sg13g2_and3_1 _15368_ (.X(_09610_),
    .A(_08773_),
    .B(net970),
    .C(_08781_));
 sg13g2_buf_2 _15369_ (.A(_09610_),
    .X(_09611_));
 sg13g2_buf_1 _15370_ (.A(_09611_),
    .X(_09612_));
 sg13g2_nand2_1 _15371_ (.Y(_09613_),
    .A(_00155_),
    .B(net888));
 sg13g2_buf_8 _15372_ (.A(net891),
    .X(_09614_));
 sg13g2_buf_1 _15373_ (.A(net878),
    .X(_09615_));
 sg13g2_buf_1 _15374_ (.A(_08785_),
    .X(_09616_));
 sg13g2_buf_1 _15375_ (.A(net1029),
    .X(_09617_));
 sg13g2_buf_1 _15376_ (.A(_09617_),
    .X(_09618_));
 sg13g2_inv_1 _15377_ (.Y(_09619_),
    .A(_00156_));
 sg13g2_buf_8 _15378_ (.A(_08788_),
    .X(_09620_));
 sg13g2_buf_1 _15379_ (.A(net950),
    .X(_09621_));
 sg13g2_buf_8 _15380_ (.A(net919),
    .X(_09622_));
 sg13g2_a22oi_1 _15381_ (.Y(_09623_),
    .B1(net899),
    .B2(\top_ihp.wb_coproc.dat_o[24] ),
    .A2(_09619_),
    .A1(net951));
 sg13g2_nand2_1 _15382_ (.Y(_09624_),
    .A(_09615_),
    .B(_09623_));
 sg13g2_nand3_1 _15383_ (.B(_09613_),
    .C(_09624_),
    .A(net855),
    .Y(_09625_));
 sg13g2_nand2b_1 _15384_ (.Y(_09626_),
    .B(_00075_),
    .A_N(_08792_));
 sg13g2_buf_1 _15385_ (.A(_09626_),
    .X(_09627_));
 sg13g2_a21oi_2 _15386_ (.B1(net993),
    .Y(_09628_),
    .A2(_09625_),
    .A1(_09606_));
 sg13g2_and2_1 _15387_ (.A(net1030),
    .B(_09628_),
    .X(_09629_));
 sg13g2_nor2_1 _15388_ (.A(_00130_),
    .B(net879),
    .Y(_09630_));
 sg13g2_buf_1 _15389_ (.A(_08772_),
    .X(_09631_));
 sg13g2_buf_8 _15390_ (.A(net888),
    .X(_09632_));
 sg13g2_inv_1 _15391_ (.Y(_09633_),
    .A(_00132_));
 sg13g2_a221oi_1 _15392_ (.B2(\top_ihp.wb_coproc.dat_o[8] ),
    .C1(net888),
    .B1(net899),
    .A1(net951),
    .Y(_09634_),
    .A2(_09633_));
 sg13g2_a221oi_1 _15393_ (.B2(_00131_),
    .C1(_09634_),
    .B1(net877),
    .A1(net992),
    .Y(_09635_),
    .A2(net905));
 sg13g2_o21ai_1 _15394_ (.B1(_08794_),
    .Y(_09636_),
    .A1(_09630_),
    .A2(_09635_));
 sg13g2_nor2_1 _15395_ (.A(net1030),
    .B(_09636_),
    .Y(_09637_));
 sg13g2_buf_8 _15396_ (.A(\top_ihp.oisc.mem_addr_lowbits[0] ),
    .X(_09638_));
 sg13g2_nor2_1 _15397_ (.A(net1056),
    .B(_08474_),
    .Y(_09639_));
 sg13g2_and2_1 _15398_ (.A(_09638_),
    .B(_09639_),
    .X(_09640_));
 sg13g2_buf_1 _15399_ (.A(_09640_),
    .X(_09641_));
 sg13g2_o21ai_1 _15400_ (.B1(_09641_),
    .Y(_09642_),
    .A1(_09629_),
    .A2(_09637_));
 sg13g2_nand2b_1 _15401_ (.Y(_09643_),
    .B(_09638_),
    .A_N(_08479_));
 sg13g2_buf_1 _15402_ (.A(_09643_),
    .X(_09644_));
 sg13g2_nand2_1 _15403_ (.Y(_09645_),
    .A(_00115_),
    .B(net920));
 sg13g2_nand3_1 _15404_ (.B(net904),
    .C(_09611_),
    .A(_00116_),
    .Y(_09646_));
 sg13g2_inv_1 _15405_ (.Y(_09647_),
    .A(_00117_));
 sg13g2_a22oi_1 _15406_ (.Y(_09648_),
    .B1(net950),
    .B2(\top_ihp.wb_coproc.dat_o[16] ),
    .A2(_09647_),
    .A1(_08785_));
 sg13g2_nand3_1 _15407_ (.B(net891),
    .C(_09648_),
    .A(net904),
    .Y(_09649_));
 sg13g2_and4_1 _15408_ (.A(_08799_),
    .B(_09645_),
    .C(_09646_),
    .D(_09649_),
    .X(_09650_));
 sg13g2_buf_1 _15409_ (.A(_09650_),
    .X(_09651_));
 sg13g2_inv_1 _15410_ (.Y(_09652_),
    .A(_09601_));
 sg13g2_buf_1 _15411_ (.A(_09652_),
    .X(_09653_));
 sg13g2_nor2_1 _15412_ (.A(net1042),
    .B(net991),
    .Y(_09654_));
 sg13g2_buf_1 _15413_ (.A(_09654_),
    .X(_09655_));
 sg13g2_nand3_1 _15414_ (.B(_09651_),
    .C(net918),
    .A(_09644_),
    .Y(_09656_));
 sg13g2_buf_8 _15415_ (.A(net1042),
    .X(_09657_));
 sg13g2_nor2b_1 _15416_ (.A(net1056),
    .B_N(_09638_),
    .Y(_09658_));
 sg13g2_buf_1 _15417_ (.A(_09658_),
    .X(_09659_));
 sg13g2_nor2_1 _15418_ (.A(net1030),
    .B(_09659_),
    .Y(_09660_));
 sg13g2_buf_1 _15419_ (.A(_08797_),
    .X(_09661_));
 sg13g2_inv_1 _15420_ (.Y(_09662_),
    .A(\top_ihp.wb_dati_ram[0] ));
 sg13g2_a22oi_1 _15421_ (.Y(_09663_),
    .B1(\top_ihp.wb_coproc.dat_o[0] ),
    .B2(net899),
    .A2(\top_ihp.wb_dati_spi[0] ),
    .A1(net951));
 sg13g2_mux2_1 _15422_ (.A0(_09662_),
    .A1(_09663_),
    .S(net854),
    .X(_09664_));
 sg13g2_nand2_1 _15423_ (.Y(_09665_),
    .A(\top_ihp.wb_dati_rom[0] ),
    .B(net920));
 sg13g2_o21ai_1 _15424_ (.B1(_09665_),
    .Y(_09666_),
    .A1(net900),
    .A2(_09664_));
 sg13g2_nand2b_1 _15425_ (.Y(_09667_),
    .B(_08792_),
    .A_N(\top_ihp.wb_dati_gpio[0] ));
 sg13g2_o21ai_1 _15426_ (.B1(_09667_),
    .Y(_09668_),
    .A1(_08792_),
    .A2(_09666_));
 sg13g2_nand2_1 _15427_ (.Y(_09669_),
    .A(net1028),
    .B(\top_ihp.wb_dati_uart[0] ));
 sg13g2_o21ai_1 _15428_ (.B1(_09669_),
    .Y(_09670_),
    .A1(_09661_),
    .A2(_09668_));
 sg13g2_o21ai_1 _15429_ (.B1(_09670_),
    .Y(_09671_),
    .A1(net990),
    .A2(_09660_));
 sg13g2_nand4_1 _15430_ (.B(_09656_),
    .C(_09671_),
    .A(_09642_),
    .Y(_09672_),
    .D(net952));
 sg13g2_o21ai_1 _15431_ (.B1(_09672_),
    .Y(_09673_),
    .A1(_09507_),
    .A2(net921));
 sg13g2_buf_1 _15432_ (.A(\top_ihp.oisc.decoder.decoded[13] ),
    .X(_09674_));
 sg13g2_buf_1 _15433_ (.A(_09674_),
    .X(_09675_));
 sg13g2_buf_1 _15434_ (.A(net1027),
    .X(_09676_));
 sg13g2_buf_2 _15435_ (.A(_00085_),
    .X(_09677_));
 sg13g2_buf_1 _15436_ (.A(_09677_),
    .X(_09678_));
 sg13g2_buf_1 _15437_ (.A(\top_ihp.oisc.decoder.instruction[7] ),
    .X(_09679_));
 sg13g2_nand3_1 _15438_ (.B(net1026),
    .C(_09679_),
    .A(_09676_),
    .Y(_09680_));
 sg13g2_buf_2 _15439_ (.A(\top_ihp.oisc.decoder.instruction[20] ),
    .X(_09681_));
 sg13g2_buf_1 _15440_ (.A(\top_ihp.oisc.decoder.decoded[15] ),
    .X(_09682_));
 sg13g2_nand2_1 _15441_ (.Y(_09683_),
    .A(net1027),
    .B(_09682_));
 sg13g2_inv_1 _15442_ (.Y(_09684_),
    .A(_09675_));
 sg13g2_nand2_1 _15443_ (.Y(_09685_),
    .A(_09684_),
    .B(_09677_));
 sg13g2_o21ai_1 _15444_ (.B1(_09685_),
    .Y(_09686_),
    .A1(_09678_),
    .A2(_09683_));
 sg13g2_nand2_1 _15445_ (.Y(_09687_),
    .A(_09681_),
    .B(_09686_));
 sg13g2_buf_2 _15446_ (.A(\top_ihp.oisc.decoder.decoded[14] ),
    .X(_09688_));
 sg13g2_buf_1 _15447_ (.A(_09688_),
    .X(_09689_));
 sg13g2_a21oi_1 _15448_ (.A1(_09680_),
    .A2(_09687_),
    .Y(_09690_),
    .B1(net1025));
 sg13g2_nor2_1 _15449_ (.A(net995),
    .B(_09690_),
    .Y(_09691_));
 sg13g2_a21oi_1 _15450_ (.A1(net995),
    .A2(_09673_),
    .Y(_09692_),
    .B1(_09691_));
 sg13g2_buf_1 _15451_ (.A(net996),
    .X(_09693_));
 sg13g2_nor2b_1 _15452_ (.A(net949),
    .B_N(_08082_),
    .Y(_09694_));
 sg13g2_a21oi_1 _15453_ (.A1(net953),
    .A2(_09692_),
    .Y(_09695_),
    .B1(_09694_));
 sg13g2_buf_2 _15454_ (.A(_09695_),
    .X(_09696_));
 sg13g2_buf_8 _15455_ (.A(_09696_),
    .X(_09697_));
 sg13g2_buf_8 _15456_ (.A(net156),
    .X(_09698_));
 sg13g2_inv_1 _15457_ (.Y(_09699_),
    .A(_09682_));
 sg13g2_nor2_2 _15458_ (.A(_09674_),
    .B(_09699_),
    .Y(_09700_));
 sg13g2_nand2_1 _15459_ (.Y(_09701_),
    .A(_09688_),
    .B(_09700_));
 sg13g2_inv_1 _15460_ (.Y(_09702_),
    .A(_09701_));
 sg13g2_buf_1 _15461_ (.A(\top_ihp.oisc.decoder.decoded[12] ),
    .X(_09703_));
 sg13g2_a221oi_1 _15462_ (.B2(_09703_),
    .C1(_09488_),
    .B1(_09487_),
    .A1(net1058),
    .Y(_09704_),
    .A2(_08823_));
 sg13g2_buf_1 _15463_ (.A(_09704_),
    .X(_09705_));
 sg13g2_nand2_1 _15464_ (.Y(_09706_),
    .A(net1058),
    .B(_08823_));
 sg13g2_buf_8 _15465_ (.A(_09706_),
    .X(_09707_));
 sg13g2_nand4_1 _15466_ (.B(_09703_),
    .C(_07966_),
    .A(_07959_),
    .Y(_09708_),
    .D(_07971_));
 sg13g2_xor2_1 _15467_ (.B(_09674_),
    .A(_09688_),
    .X(_09709_));
 sg13g2_a22oi_1 _15468_ (.Y(_09710_),
    .B1(_09709_),
    .B2(_09677_),
    .A2(_09708_),
    .A1(_09707_));
 sg13g2_buf_2 _15469_ (.A(_09710_),
    .X(_09711_));
 sg13g2_buf_1 _15470_ (.A(\top_ihp.oisc.decoder.instruction[10] ),
    .X(_09712_));
 sg13g2_a221oi_1 _15471_ (.B2(_09712_),
    .C1(_09594_),
    .B1(_09711_),
    .A1(\top_ihp.oisc.micro_res_addr[3] ),
    .Y(_09713_),
    .A2(_09705_));
 sg13g2_a21oi_2 _15472_ (.B1(_09713_),
    .Y(_09714_),
    .A2(_09702_),
    .A1(net1051));
 sg13g2_buf_1 _15473_ (.A(\top_ihp.oisc.decoder.instruction[9] ),
    .X(_09715_));
 sg13g2_inv_1 _15474_ (.Y(_09716_),
    .A(\top_ihp.oisc.micro_res_addr[2] ));
 sg13g2_nor3_1 _15475_ (.A(_09716_),
    .B(_09488_),
    .C(_09598_),
    .Y(_09717_));
 sg13g2_nand2_1 _15476_ (.Y(_09718_),
    .A(_09703_),
    .B(net922));
 sg13g2_a221oi_1 _15477_ (.B2(_09718_),
    .C1(net1051),
    .B1(_09717_),
    .A1(_09715_),
    .Y(_09719_),
    .A2(_09711_));
 sg13g2_a21oi_1 _15478_ (.A1(net1051),
    .A2(_09701_),
    .Y(_09720_),
    .B1(_09719_));
 sg13g2_or2_1 _15479_ (.X(_09721_),
    .B(_09720_),
    .A(_09494_));
 sg13g2_buf_1 _15480_ (.A(_09721_),
    .X(_09722_));
 sg13g2_buf_2 _15481_ (.A(_00087_),
    .X(_09723_));
 sg13g2_o21ai_1 _15482_ (.B1(_09723_),
    .Y(_09724_),
    .A1(_09714_),
    .A2(_09722_));
 sg13g2_buf_1 _15483_ (.A(_09724_),
    .X(_09725_));
 sg13g2_buf_1 _15484_ (.A(_09725_),
    .X(_09726_));
 sg13g2_nand2_1 _15485_ (.Y(_09727_),
    .A(_09532_),
    .B(_09723_));
 sg13g2_nor2_1 _15486_ (.A(net1051),
    .B(_09727_),
    .Y(_09728_));
 sg13g2_nand2b_1 _15487_ (.Y(_09729_),
    .B(_09728_),
    .A_N(_09705_));
 sg13g2_buf_1 _15488_ (.A(\top_ihp.oisc.decoder.instruction[11] ),
    .X(_09730_));
 sg13g2_nand3_1 _15489_ (.B(_09711_),
    .C(_09728_),
    .A(_09730_),
    .Y(_09731_));
 sg13g2_inv_1 _15490_ (.Y(_09732_),
    .A(net1052));
 sg13g2_nand2_1 _15491_ (.Y(_09733_),
    .A(_09732_),
    .B(_09532_));
 sg13g2_nor2_1 _15492_ (.A(net1051),
    .B(_09733_),
    .Y(_09734_));
 sg13g2_buf_2 _15493_ (.A(\top_ihp.oisc.state[0] ),
    .X(_09735_));
 sg13g2_a21oi_1 _15494_ (.A1(_09703_),
    .A2(_08823_),
    .Y(_09736_),
    .B1(_09735_));
 sg13g2_nand3_1 _15495_ (.B(_09734_),
    .C(_09736_),
    .A(_09488_),
    .Y(_09737_));
 sg13g2_and2_1 _15496_ (.A(_09731_),
    .B(_09737_),
    .X(_09738_));
 sg13g2_nand2_2 _15497_ (.Y(_09739_),
    .A(_09729_),
    .B(_09738_));
 sg13g2_buf_1 _15498_ (.A(\top_ihp.oisc.decoder.instruction[8] ),
    .X(_09740_));
 sg13g2_a22oi_1 _15499_ (.Y(_09741_),
    .B1(_09711_),
    .B2(_09740_),
    .A2(_09705_),
    .A1(\top_ihp.oisc.micro_res_addr[1] ));
 sg13g2_nand2b_1 _15500_ (.Y(_09742_),
    .B(_00086_),
    .A_N(_09741_));
 sg13g2_buf_2 _15501_ (.A(_09742_),
    .X(_09743_));
 sg13g2_o21ai_1 _15502_ (.B1(_09732_),
    .Y(_09744_),
    .A1(net1051),
    .A2(_09743_));
 sg13g2_nand2_1 _15503_ (.Y(_09745_),
    .A(_09679_),
    .B(_09711_));
 sg13g2_nand2_1 _15504_ (.Y(_09746_),
    .A(\top_ihp.oisc.micro_res_addr[0] ),
    .B(_09705_));
 sg13g2_nand2_1 _15505_ (.Y(_09747_),
    .A(_09595_),
    .B(net996));
 sg13g2_buf_1 _15506_ (.A(_09747_),
    .X(_09748_));
 sg13g2_a21o_1 _15507_ (.A2(_09746_),
    .A1(_09745_),
    .B1(net917),
    .X(_09749_));
 sg13g2_buf_2 _15508_ (.A(_09749_),
    .X(_09750_));
 sg13g2_nor2b_1 _15509_ (.A(_09744_),
    .B_N(_09750_),
    .Y(_09751_));
 sg13g2_buf_8 _15510_ (.A(_09751_),
    .X(_09752_));
 sg13g2_nor2b_1 _15511_ (.A(_09739_),
    .B_N(net766),
    .Y(_09753_));
 sg13g2_buf_1 _15512_ (.A(_09753_),
    .X(_09754_));
 sg13g2_nand2_1 _15513_ (.Y(_09755_),
    .A(net767),
    .B(_09754_));
 sg13g2_buf_1 _15514_ (.A(_09755_),
    .X(_09756_));
 sg13g2_buf_1 _15515_ (.A(net661),
    .X(_09757_));
 sg13g2_buf_1 _15516_ (.A(_09755_),
    .X(_09758_));
 sg13g2_nand2_1 _15517_ (.Y(_09759_),
    .A(\top_ihp.oisc.regs[0][0] ),
    .B(net660));
 sg13g2_o21ai_1 _15518_ (.B1(_09759_),
    .Y(_00452_),
    .A1(net53),
    .A2(_09757_));
 sg13g2_inv_1 _15519_ (.Y(_09760_),
    .A(net1065));
 sg13g2_inv_1 _15520_ (.Y(_09761_),
    .A(_09688_));
 sg13g2_o21ai_1 _15521_ (.B1(_09761_),
    .Y(_09762_),
    .A1(_09677_),
    .A2(_09700_));
 sg13g2_a21oi_1 _15522_ (.A1(_09685_),
    .A2(_09762_),
    .Y(_09763_),
    .B1(_09595_));
 sg13g2_buf_2 _15523_ (.A(_09763_),
    .X(_09764_));
 sg13g2_a21o_1 _15524_ (.A2(_08789_),
    .A1(net891),
    .B1(_08790_),
    .X(_09765_));
 sg13g2_inv_1 _15525_ (.Y(_09766_),
    .A(_00174_));
 sg13g2_a22oi_1 _15526_ (.Y(_09767_),
    .B1(net950),
    .B2(\top_ihp.wb_coproc.dat_o[31] ),
    .A2(_09766_),
    .A1(net1029));
 sg13g2_mux2_1 _15527_ (.A0(_00173_),
    .A1(_09767_),
    .S(net891),
    .X(_09768_));
 sg13g2_mux4_1 _15528_ (.S0(_09601_),
    .A0(_00112_),
    .A1(_00172_),
    .A2(_09765_),
    .A3(_09768_),
    .S1(net889),
    .X(_09769_));
 sg13g2_nor2_2 _15529_ (.A(net993),
    .B(_09769_),
    .Y(_09770_));
 sg13g2_and2_1 _15530_ (.A(_09638_),
    .B(_09770_),
    .X(_09771_));
 sg13g2_nor2_1 _15531_ (.A(_00151_),
    .B(net904),
    .Y(_09772_));
 sg13g2_inv_1 _15532_ (.Y(_09773_),
    .A(_00153_));
 sg13g2_a22oi_1 _15533_ (.Y(_09774_),
    .B1(_08788_),
    .B2(\top_ihp.wb_coproc.dat_o[23] ),
    .A2(_09773_),
    .A1(_08785_));
 sg13g2_and4_1 _15534_ (.A(_08773_),
    .B(_00152_),
    .C(net970),
    .D(_08781_),
    .X(_09775_));
 sg13g2_a221oi_1 _15535_ (.B2(_09774_),
    .C1(_09775_),
    .B1(_08784_),
    .A1(net1041),
    .Y(_09776_),
    .A2(_08371_));
 sg13g2_o21ai_1 _15536_ (.B1(_08794_),
    .Y(_09777_),
    .A1(_09772_),
    .A2(_09776_));
 sg13g2_and2_1 _15537_ (.A(_09601_),
    .B(_09777_),
    .X(_09778_));
 sg13g2_buf_1 _15538_ (.A(_09778_),
    .X(_09779_));
 sg13g2_nand2_1 _15539_ (.Y(_09780_),
    .A(net1028),
    .B(\top_ihp.wb_dati_uart[7] ));
 sg13g2_nor2_1 _15540_ (.A(_00127_),
    .B(_08770_),
    .Y(_09781_));
 sg13g2_inv_1 _15541_ (.Y(_09782_),
    .A(_00129_));
 sg13g2_a22oi_1 _15542_ (.Y(_09783_),
    .B1(net950),
    .B2(\top_ihp.wb_coproc.dat_o[7] ),
    .A2(_09782_),
    .A1(_08785_));
 sg13g2_buf_1 _15543_ (.A(_08773_),
    .X(_09784_));
 sg13g2_and4_1 _15544_ (.A(net1024),
    .B(_00128_),
    .C(net970),
    .D(_08781_),
    .X(_09785_));
 sg13g2_a221oi_1 _15545_ (.B2(_09783_),
    .C1(_09785_),
    .B1(net891),
    .A1(net1041),
    .Y(_09786_),
    .A2(_08371_));
 sg13g2_nor2b_1 _15546_ (.A(_08797_),
    .B_N(_08219_),
    .Y(_09787_));
 sg13g2_buf_1 _15547_ (.A(_09787_),
    .X(_09788_));
 sg13g2_o21ai_1 _15548_ (.B1(net987),
    .Y(_09789_),
    .A1(_09781_),
    .A2(_09786_));
 sg13g2_and3_1 _15549_ (.X(_09790_),
    .A(net991),
    .B(_09780_),
    .C(_09789_));
 sg13g2_buf_1 _15550_ (.A(_09790_),
    .X(_09791_));
 sg13g2_nor3_1 _15551_ (.A(_09638_),
    .B(_09779_),
    .C(_09791_),
    .Y(_09792_));
 sg13g2_buf_1 _15552_ (.A(\top_ihp.oisc.decoder.instruction[14] ),
    .X(_09793_));
 sg13g2_nor3_1 _15553_ (.A(net1056),
    .B(_08475_),
    .C(_09793_),
    .Y(_09794_));
 sg13g2_o21ai_1 _15554_ (.B1(_09794_),
    .Y(_09795_),
    .A1(_09771_),
    .A2(_09792_));
 sg13g2_and2_1 _15555_ (.A(_09598_),
    .B(_09795_),
    .X(_09796_));
 sg13g2_buf_8 _15556_ (.A(_09796_),
    .X(_09797_));
 sg13g2_buf_1 _15557_ (.A(_08475_),
    .X(_09798_));
 sg13g2_nand2b_1 _15558_ (.Y(_09799_),
    .B(net920),
    .A_N(_00136_));
 sg13g2_nand2_1 _15559_ (.Y(_09800_),
    .A(_00137_),
    .B(net888));
 sg13g2_inv_1 _15560_ (.Y(_09801_),
    .A(_00138_));
 sg13g2_a22oi_1 _15561_ (.Y(_09802_),
    .B1(net919),
    .B2(\top_ihp.wb_coproc.dat_o[10] ),
    .A2(_09801_),
    .A1(net994));
 sg13g2_nand2_1 _15562_ (.Y(_09803_),
    .A(net854),
    .B(_09802_));
 sg13g2_nand3_1 _15563_ (.B(_09800_),
    .C(_09803_),
    .A(net879),
    .Y(_09804_));
 sg13g2_a21oi_2 _15564_ (.B1(net993),
    .Y(_09805_),
    .A2(_09804_),
    .A1(_09799_));
 sg13g2_nand2b_1 _15565_ (.Y(_09806_),
    .B(net920),
    .A_N(_00160_));
 sg13g2_nand2_1 _15566_ (.Y(_09807_),
    .A(_00161_),
    .B(_09612_));
 sg13g2_inv_1 _15567_ (.Y(_09808_),
    .A(_00162_));
 sg13g2_a22oi_1 _15568_ (.Y(_09809_),
    .B1(net919),
    .B2(\top_ihp.wb_coproc.dat_o[26] ),
    .A2(_09808_),
    .A1(net994));
 sg13g2_nand2_1 _15569_ (.Y(_09810_),
    .A(net854),
    .B(_09809_));
 sg13g2_nand3_1 _15570_ (.B(_09807_),
    .C(_09810_),
    .A(net879),
    .Y(_09811_));
 sg13g2_a21oi_2 _15571_ (.B1(net993),
    .Y(_09812_),
    .A2(_09811_),
    .A1(_09806_));
 sg13g2_a22oi_1 _15572_ (.Y(_09813_),
    .B1(_09812_),
    .B2(net918),
    .A2(_09805_),
    .A1(net991));
 sg13g2_inv_1 _15573_ (.Y(_09814_),
    .A(_09813_));
 sg13g2_buf_1 _15574_ (.A(net1056),
    .X(_09815_));
 sg13g2_a22oi_1 _15575_ (.Y(_09816_),
    .B1(_09814_),
    .B2(net1023),
    .A2(_09805_),
    .A1(net986));
 sg13g2_xnor2_1 _15576_ (.Y(_09817_),
    .A(_08030_),
    .B(_08145_));
 sg13g2_xnor2_1 _15577_ (.Y(_09818_),
    .A(_09760_),
    .B(_09817_));
 sg13g2_buf_1 _15578_ (.A(net988),
    .X(_09819_));
 sg13g2_buf_8 _15579_ (.A(net1051),
    .X(_09820_));
 sg13g2_a221oi_1 _15580_ (.B2(net948),
    .C1(net1022),
    .B1(_09818_),
    .A1(_09797_),
    .Y(_09821_),
    .A2(_09816_));
 sg13g2_a21oi_1 _15581_ (.A1(\top_ihp.oisc.decoder.instruction[30] ),
    .A2(_09764_),
    .Y(_09822_),
    .B1(_09821_));
 sg13g2_mux2_1 _15582_ (.A0(_09760_),
    .A1(_09822_),
    .S(net949),
    .X(_09823_));
 sg13g2_buf_2 _15583_ (.A(_09823_),
    .X(_09824_));
 sg13g2_buf_2 _15584_ (.A(_09824_),
    .X(_09825_));
 sg13g2_nand2_1 _15585_ (.Y(_09826_),
    .A(\top_ihp.oisc.regs[0][10] ),
    .B(net660));
 sg13g2_o21ai_1 _15586_ (.B1(_09826_),
    .Y(_00453_),
    .A1(net531),
    .A2(net155));
 sg13g2_nand2b_1 _15587_ (.Y(_09827_),
    .B(net920),
    .A_N(_00139_));
 sg13g2_nand2_1 _15588_ (.Y(_09828_),
    .A(_00140_),
    .B(_09612_));
 sg13g2_inv_1 _15589_ (.Y(_09829_),
    .A(_00141_));
 sg13g2_a22oi_1 _15590_ (.Y(_09830_),
    .B1(net919),
    .B2(\top_ihp.wb_coproc.dat_o[11] ),
    .A2(_09829_),
    .A1(net994));
 sg13g2_nand2_1 _15591_ (.Y(_09831_),
    .A(net854),
    .B(_09830_));
 sg13g2_nand3_1 _15592_ (.B(_09828_),
    .C(_09831_),
    .A(net879),
    .Y(_09832_));
 sg13g2_a21oi_1 _15593_ (.A1(_09827_),
    .A2(_09832_),
    .Y(_09833_),
    .B1(net993));
 sg13g2_inv_1 _15594_ (.Y(_09834_),
    .A(net1042));
 sg13g2_nand2_1 _15595_ (.Y(_09835_),
    .A(_09834_),
    .B(_09601_));
 sg13g2_nor2_1 _15596_ (.A(_00163_),
    .B(net879),
    .Y(_09836_));
 sg13g2_inv_1 _15597_ (.Y(_09837_),
    .A(_00165_));
 sg13g2_a221oi_1 _15598_ (.B2(\top_ihp.wb_coproc.dat_o[27] ),
    .C1(_09611_),
    .B1(_09621_),
    .A1(_09617_),
    .Y(_09838_),
    .A2(_09837_));
 sg13g2_a221oi_1 _15599_ (.B2(_00164_),
    .C1(_09838_),
    .B1(net888),
    .A1(net992),
    .Y(_09839_),
    .A2(net905));
 sg13g2_o21ai_1 _15600_ (.B1(_08794_),
    .Y(_09840_),
    .A1(_09836_),
    .A2(_09839_));
 sg13g2_buf_1 _15601_ (.A(_09840_),
    .X(_09841_));
 sg13g2_nand2_1 _15602_ (.Y(_09842_),
    .A(net991),
    .B(_09833_));
 sg13g2_o21ai_1 _15603_ (.B1(_09842_),
    .Y(_09843_),
    .A1(_09835_),
    .A2(_09841_));
 sg13g2_a22oi_1 _15604_ (.Y(_09844_),
    .B1(_09843_),
    .B2(net1023),
    .A2(_09833_),
    .A1(net986));
 sg13g2_a21oi_1 _15605_ (.A1(_08029_),
    .A2(_08414_),
    .Y(_09845_),
    .B1(_08145_));
 sg13g2_or2_1 _15606_ (.X(_09846_),
    .B(_09845_),
    .A(_08031_));
 sg13g2_o21ai_1 _15607_ (.B1(_08421_),
    .Y(_09847_),
    .A1(_08042_),
    .A2(_09846_));
 sg13g2_buf_1 _15608_ (.A(net988),
    .X(_09848_));
 sg13g2_buf_1 _15609_ (.A(net1022),
    .X(_09849_));
 sg13g2_a221oi_1 _15610_ (.B2(net947),
    .C1(net985),
    .B1(_09847_),
    .A1(_09797_),
    .Y(_09850_),
    .A2(_09844_));
 sg13g2_buf_2 _15611_ (.A(\top_ihp.oisc.decoder.instruction[31] ),
    .X(_09851_));
 sg13g2_nor2b_1 _15612_ (.A(net1026),
    .B_N(_09681_),
    .Y(_09852_));
 sg13g2_a22oi_1 _15613_ (.Y(_09853_),
    .B1(_09700_),
    .B2(_09852_),
    .A2(_09851_),
    .A1(net1026));
 sg13g2_nand4_1 _15614_ (.B(_09684_),
    .C(net1026),
    .A(net1025),
    .Y(_09854_),
    .D(_09679_));
 sg13g2_o21ai_1 _15615_ (.B1(_09854_),
    .Y(_09855_),
    .A1(net1025),
    .A2(_09853_));
 sg13g2_buf_8 _15616_ (.A(_09733_),
    .X(_09856_));
 sg13g2_a21oi_1 _15617_ (.A1(net985),
    .A2(_09855_),
    .Y(_09857_),
    .B1(_09856_));
 sg13g2_nand2b_1 _15618_ (.Y(_09858_),
    .B(_09857_),
    .A_N(_09850_));
 sg13g2_o21ai_1 _15619_ (.B1(_09858_),
    .Y(_09859_),
    .A1(net1063),
    .A2(net953));
 sg13g2_buf_2 _15620_ (.A(_09859_),
    .X(_09860_));
 sg13g2_buf_2 _15621_ (.A(_09860_),
    .X(_09861_));
 sg13g2_nand2_1 _15622_ (.Y(_09862_),
    .A(\top_ihp.oisc.regs[0][11] ),
    .B(net660));
 sg13g2_o21ai_1 _15623_ (.B1(_09862_),
    .Y(_00454_),
    .A1(net531),
    .A2(net154));
 sg13g2_buf_1 _15624_ (.A(net946),
    .X(_09863_));
 sg13g2_buf_1 _15625_ (.A(net916),
    .X(_09864_));
 sg13g2_buf_1 _15626_ (.A(net946),
    .X(_09865_));
 sg13g2_nor2_1 _15627_ (.A(_00076_),
    .B(net889),
    .Y(_09866_));
 sg13g2_a21oi_1 _15628_ (.A1(\top_ihp.wb_coproc.dat_o[12] ),
    .A2(_08374_),
    .Y(_09867_),
    .B1(net1029));
 sg13g2_a21o_1 _15629_ (.A2(net1029),
    .A1(_00078_),
    .B1(_09867_),
    .X(_09868_));
 sg13g2_buf_1 _15630_ (.A(net970),
    .X(_09869_));
 sg13g2_buf_1 _15631_ (.A(_08781_),
    .X(_09870_));
 sg13g2_and4_1 _15632_ (.A(_09784_),
    .B(_00077_),
    .C(net914),
    .D(net913),
    .X(_09871_));
 sg13g2_a221oi_1 _15633_ (.B2(_09868_),
    .C1(_09871_),
    .B1(net878),
    .A1(net1041),
    .Y(_09872_),
    .A2(net905));
 sg13g2_nor2_1 _15634_ (.A(_09866_),
    .B(_09872_),
    .Y(_09873_));
 sg13g2_nor2_1 _15635_ (.A(_09627_),
    .B(_09873_),
    .Y(_09874_));
 sg13g2_buf_1 _15636_ (.A(_09874_),
    .X(_09875_));
 sg13g2_nand2b_1 _15637_ (.Y(_09876_),
    .B(net900),
    .A_N(_00166_));
 sg13g2_nand2_1 _15638_ (.Y(_09877_),
    .A(_00167_),
    .B(net888));
 sg13g2_inv_1 _15639_ (.Y(_09878_),
    .A(_00168_));
 sg13g2_a22oi_1 _15640_ (.Y(_09879_),
    .B1(net899),
    .B2(\top_ihp.wb_coproc.dat_o[28] ),
    .A2(_09878_),
    .A1(net951));
 sg13g2_nand2_1 _15641_ (.Y(_09880_),
    .A(net854),
    .B(_09879_));
 sg13g2_nand3_1 _15642_ (.B(_09877_),
    .C(_09880_),
    .A(net879),
    .Y(_09881_));
 sg13g2_a21oi_2 _15643_ (.B1(net993),
    .Y(_09882_),
    .A2(_09881_),
    .A1(_09876_));
 sg13g2_o21ai_1 _15644_ (.B1(_08794_),
    .Y(_09883_),
    .A1(_09866_),
    .A2(_09872_));
 sg13g2_buf_1 _15645_ (.A(_09883_),
    .X(_09884_));
 sg13g2_nor2_1 _15646_ (.A(_09601_),
    .B(_09884_),
    .Y(_09885_));
 sg13g2_a21o_1 _15647_ (.A2(_09882_),
    .A1(_09655_),
    .B1(_09885_),
    .X(_09886_));
 sg13g2_a22oi_1 _15648_ (.Y(_09887_),
    .B1(_09886_),
    .B2(net1023),
    .A2(net788),
    .A1(_09798_));
 sg13g2_nand3_1 _15649_ (.B(_09795_),
    .C(_09887_),
    .A(_09599_),
    .Y(_09888_));
 sg13g2_xnor2_1 _15650_ (.Y(_09889_),
    .A(_08045_),
    .B(_08230_));
 sg13g2_nand2_1 _15651_ (.Y(_09890_),
    .A(net948),
    .B(_09889_));
 sg13g2_a21oi_1 _15652_ (.A1(_09888_),
    .A2(_09890_),
    .Y(_09891_),
    .B1(net985));
 sg13g2_and3_1 _15653_ (.X(_09892_),
    .A(net1025),
    .B(net1027),
    .C(_09677_));
 sg13g2_buf_2 _15654_ (.A(_09892_),
    .X(_09893_));
 sg13g2_nor2_1 _15655_ (.A(_09688_),
    .B(_09677_),
    .Y(_09894_));
 sg13g2_nand2_1 _15656_ (.Y(_09895_),
    .A(_09700_),
    .B(_09894_));
 sg13g2_buf_1 _15657_ (.A(_09895_),
    .X(_09896_));
 sg13g2_nand2b_1 _15658_ (.Y(_09897_),
    .B(_09896_),
    .A_N(_09893_));
 sg13g2_nand2_1 _15659_ (.Y(_09898_),
    .A(net1025),
    .B(net1027));
 sg13g2_nand3_1 _15660_ (.B(_09851_),
    .C(_09898_),
    .A(_09677_),
    .Y(_09899_));
 sg13g2_nand2_1 _15661_ (.Y(_09900_),
    .A(net1022),
    .B(_09899_));
 sg13g2_buf_2 _15662_ (.A(_09900_),
    .X(_09901_));
 sg13g2_a21oi_1 _15663_ (.A1(net1023),
    .A2(_09897_),
    .Y(_09902_),
    .B1(_09901_));
 sg13g2_nor3_2 _15664_ (.A(net915),
    .B(_09891_),
    .C(_09902_),
    .Y(_09903_));
 sg13g2_a21oi_1 _15665_ (.A1(net1064),
    .A2(net898),
    .Y(_09904_),
    .B1(_09903_));
 sg13g2_buf_2 _15666_ (.A(_09904_),
    .X(_09905_));
 sg13g2_buf_8 _15667_ (.A(net332),
    .X(_09906_));
 sg13g2_nand2_1 _15668_ (.Y(_09907_),
    .A(\top_ihp.oisc.regs[0][12] ),
    .B(net660));
 sg13g2_o21ai_1 _15669_ (.B1(_09907_),
    .Y(_00455_),
    .A1(net531),
    .A2(_09906_));
 sg13g2_buf_1 _15670_ (.A(net990),
    .X(_09908_));
 sg13g2_buf_1 _15671_ (.A(net993),
    .X(_09909_));
 sg13g2_nor2_1 _15672_ (.A(_00082_),
    .B(net889),
    .Y(_09910_));
 sg13g2_inv_1 _15673_ (.Y(_09911_),
    .A(_00084_));
 sg13g2_a22oi_1 _15674_ (.Y(_09912_),
    .B1(net950),
    .B2(\top_ihp.wb_coproc.dat_o[13] ),
    .A2(_09911_),
    .A1(net1029));
 sg13g2_and4_1 _15675_ (.A(net1024),
    .B(_00083_),
    .C(net970),
    .D(net913),
    .X(_09913_));
 sg13g2_a221oi_1 _15676_ (.B2(_09912_),
    .C1(_09913_),
    .B1(_09614_),
    .A1(net1041),
    .Y(_09914_),
    .A2(_08371_));
 sg13g2_nor2_1 _15677_ (.A(_09910_),
    .B(_09914_),
    .Y(_09915_));
 sg13g2_nor2_1 _15678_ (.A(net944),
    .B(_09915_),
    .Y(_09916_));
 sg13g2_buf_1 _15679_ (.A(_09916_),
    .X(_09917_));
 sg13g2_nand2b_1 _15680_ (.Y(_09918_),
    .B(net900),
    .A_N(_00169_));
 sg13g2_inv_1 _15681_ (.Y(_09919_),
    .A(_00171_));
 sg13g2_a221oi_1 _15682_ (.B2(\top_ihp.wb_coproc.dat_o[29] ),
    .C1(net877),
    .B1(net899),
    .A1(_09618_),
    .Y(_09920_),
    .A2(_09919_));
 sg13g2_a21oi_1 _15683_ (.A1(_00170_),
    .A2(net877),
    .Y(_09921_),
    .B1(_09920_));
 sg13g2_nand2_1 _15684_ (.Y(_09922_),
    .A(net855),
    .B(_09921_));
 sg13g2_a21oi_2 _15685_ (.B1(net944),
    .Y(_09923_),
    .A2(_09922_),
    .A1(_09918_));
 sg13g2_o21ai_1 _15686_ (.B1(_08794_),
    .Y(_09924_),
    .A1(_09910_),
    .A2(_09914_));
 sg13g2_buf_1 _15687_ (.A(_09924_),
    .X(_09925_));
 sg13g2_nor2_1 _15688_ (.A(_09602_),
    .B(net805),
    .Y(_09926_));
 sg13g2_a21o_1 _15689_ (.A2(_09923_),
    .A1(net918),
    .B1(_09926_),
    .X(_09927_));
 sg13g2_a22oi_1 _15690_ (.Y(_09928_),
    .B1(_09927_),
    .B2(_09815_),
    .A2(_09917_),
    .A1(net945));
 sg13g2_and4_1 _15691_ (.A(_08042_),
    .B(_08415_),
    .C(_08045_),
    .D(_08105_),
    .X(_09929_));
 sg13g2_nand2_1 _15692_ (.Y(_09930_),
    .A(_08042_),
    .B(_08045_));
 sg13g2_inv_1 _15693_ (.Y(_09931_),
    .A(_08385_));
 sg13g2_o21ai_1 _15694_ (.B1(_09931_),
    .Y(_09932_),
    .A1(_08419_),
    .A2(_09930_));
 sg13g2_a21oi_1 _15695_ (.A1(_08413_),
    .A2(_09929_),
    .Y(_09933_),
    .B1(_09932_));
 sg13g2_xnor2_1 _15696_ (.Y(_09934_),
    .A(net1046),
    .B(_09933_));
 sg13g2_xnor2_1 _15697_ (.Y(_09935_),
    .A(_08234_),
    .B(_09934_));
 sg13g2_a22oi_1 _15698_ (.Y(_09936_),
    .B1(_09935_),
    .B2(net947),
    .A2(_09928_),
    .A1(_09797_));
 sg13g2_a21oi_1 _15699_ (.A1(net945),
    .A2(_09897_),
    .Y(_09937_),
    .B1(_09901_));
 sg13g2_nor2_1 _15700_ (.A(_08046_),
    .B(net996),
    .Y(_09938_));
 sg13g2_a21oi_1 _15701_ (.A1(net949),
    .A2(_09937_),
    .Y(_09939_),
    .B1(_09938_));
 sg13g2_o21ai_1 _15702_ (.B1(_09939_),
    .Y(_09940_),
    .A1(net917),
    .A2(_09936_));
 sg13g2_buf_1 _15703_ (.A(_09940_),
    .X(_09941_));
 sg13g2_buf_2 _15704_ (.A(_09941_),
    .X(_09942_));
 sg13g2_nand2_1 _15705_ (.Y(_09943_),
    .A(\top_ihp.oisc.regs[0][13] ),
    .B(net660));
 sg13g2_o21ai_1 _15706_ (.B1(_09943_),
    .Y(_00456_),
    .A1(net531),
    .A2(net331));
 sg13g2_inv_1 _15707_ (.Y(_09944_),
    .A(_00081_));
 sg13g2_a22oi_1 _15708_ (.Y(_09945_),
    .B1(net950),
    .B2(\top_ihp.wb_coproc.dat_o[14] ),
    .A2(_09944_),
    .A1(net1029));
 sg13g2_mux2_1 _15709_ (.A0(_00080_),
    .A1(_09945_),
    .S(net878),
    .X(_09946_));
 sg13g2_mux2_1 _15710_ (.A0(_00079_),
    .A1(_09946_),
    .S(net889),
    .X(_09947_));
 sg13g2_nor2_1 _15711_ (.A(net944),
    .B(_09947_),
    .Y(_09948_));
 sg13g2_buf_1 _15712_ (.A(_09948_),
    .X(_09949_));
 sg13g2_nand2b_1 _15713_ (.Y(_09950_),
    .B(_09605_),
    .A_N(_00109_));
 sg13g2_nand2_1 _15714_ (.Y(_09951_),
    .A(_00110_),
    .B(net877));
 sg13g2_inv_1 _15715_ (.Y(_09952_),
    .A(_00111_));
 sg13g2_a22oi_1 _15716_ (.Y(_09953_),
    .B1(net899),
    .B2(\top_ihp.wb_coproc.dat_o[30] ),
    .A2(_09952_),
    .A1(net951));
 sg13g2_nand2_1 _15717_ (.Y(_09954_),
    .A(net854),
    .B(_09953_));
 sg13g2_nand3_1 _15718_ (.B(_09951_),
    .C(_09954_),
    .A(net855),
    .Y(_09955_));
 sg13g2_a21oi_1 _15719_ (.A1(_09950_),
    .A2(_09955_),
    .Y(_09956_),
    .B1(_09909_));
 sg13g2_nand2b_1 _15720_ (.Y(_09957_),
    .B(_08794_),
    .A_N(_09947_));
 sg13g2_buf_2 _15721_ (.A(_09957_),
    .X(_09958_));
 sg13g2_nor2_1 _15722_ (.A(_09601_),
    .B(_09958_),
    .Y(_09959_));
 sg13g2_a21o_1 _15723_ (.A2(_09956_),
    .A1(_09655_),
    .B1(_09959_),
    .X(_09960_));
 sg13g2_a221oi_1 _15724_ (.B2(_08479_),
    .C1(_09820_),
    .B1(_09960_),
    .A1(net986),
    .Y(_09961_),
    .A2(net786));
 sg13g2_nand2_1 _15725_ (.Y(_09962_),
    .A(_09793_),
    .B(_09893_));
 sg13g2_o21ai_1 _15726_ (.B1(_09962_),
    .Y(_09963_),
    .A1(_08476_),
    .A2(_09896_));
 sg13g2_o21ai_1 _15727_ (.B1(net996),
    .Y(_09964_),
    .A1(_09901_),
    .A2(_09963_));
 sg13g2_a21o_1 _15728_ (.A2(_09961_),
    .A1(_09797_),
    .B1(_09964_),
    .X(_09965_));
 sg13g2_nor2_1 _15729_ (.A(_08234_),
    .B(net1046),
    .Y(_09966_));
 sg13g2_nand2_1 _15730_ (.Y(_09967_),
    .A(_08234_),
    .B(net1046));
 sg13g2_o21ai_1 _15731_ (.B1(_09967_),
    .Y(_09968_),
    .A1(_09966_),
    .A2(_09933_));
 sg13g2_xnor2_1 _15732_ (.Y(_09969_),
    .A(_08231_),
    .B(_09968_));
 sg13g2_inv_1 _15733_ (.Y(_09970_),
    .A(_09969_));
 sg13g2_o21ai_1 _15734_ (.B1(net953),
    .Y(_09971_),
    .A1(_09965_),
    .A2(_09970_));
 sg13g2_nor2_1 _15735_ (.A(net1022),
    .B(_09598_),
    .Y(_09972_));
 sg13g2_buf_2 _15736_ (.A(_09972_),
    .X(_09973_));
 sg13g2_o21ai_1 _15737_ (.B1(_09973_),
    .Y(_09974_),
    .A1(net1067),
    .A2(_09969_));
 sg13g2_nor2b_1 _15738_ (.A(_09965_),
    .B_N(_09974_),
    .Y(_09975_));
 sg13g2_a21oi_2 _15739_ (.B1(_09975_),
    .Y(_09976_),
    .A2(_09971_),
    .A1(net1067));
 sg13g2_buf_8 _15740_ (.A(_09976_),
    .X(_09977_));
 sg13g2_buf_8 _15741_ (.A(net330),
    .X(_09978_));
 sg13g2_nand2_1 _15742_ (.Y(_09979_),
    .A(\top_ihp.oisc.regs[0][14] ),
    .B(net660));
 sg13g2_o21ai_1 _15743_ (.B1(_09979_),
    .Y(_00457_),
    .A1(net531),
    .A2(net152));
 sg13g2_nand4_1 _15744_ (.B(_08045_),
    .C(_08048_),
    .A(_08016_),
    .Y(_09980_),
    .D(_08061_));
 sg13g2_o21ai_1 _15745_ (.B1(_08389_),
    .Y(_09981_),
    .A1(_08421_),
    .A2(_09980_));
 sg13g2_xor2_1 _15746_ (.B(_09981_),
    .A(_08060_),
    .X(_09982_));
 sg13g2_a21oi_1 _15747_ (.A1(net1056),
    .A2(_09770_),
    .Y(_09983_),
    .B1(net1042));
 sg13g2_a21o_1 _15748_ (.A2(_08796_),
    .A1(net986),
    .B1(_09983_),
    .X(_09984_));
 sg13g2_nand3_1 _15749_ (.B(_09795_),
    .C(_09984_),
    .A(net952),
    .Y(_09985_));
 sg13g2_o21ai_1 _15750_ (.B1(_09985_),
    .Y(_09986_),
    .A1(net921),
    .A2(_09982_));
 sg13g2_nand2_1 _15751_ (.Y(_09987_),
    .A(net995),
    .B(_09986_));
 sg13g2_a21oi_1 _15752_ (.A1(\top_ihp.oisc.decoder.instruction[15] ),
    .A2(_09897_),
    .Y(_09988_),
    .B1(_09901_));
 sg13g2_nor2_1 _15753_ (.A(net915),
    .B(_09988_),
    .Y(_09989_));
 sg13g2_a22oi_1 _15754_ (.Y(_09990_),
    .B1(_09987_),
    .B2(_09989_),
    .A2(net898),
    .A1(_08012_));
 sg13g2_buf_1 _15755_ (.A(_09990_),
    .X(_09991_));
 sg13g2_buf_2 _15756_ (.A(_09991_),
    .X(_09992_));
 sg13g2_buf_8 _15757_ (.A(_09992_),
    .X(_09993_));
 sg13g2_nand2_1 _15758_ (.Y(_09994_),
    .A(\top_ihp.oisc.regs[0][15] ),
    .B(net660));
 sg13g2_o21ai_1 _15759_ (.B1(_09994_),
    .Y(_00458_),
    .A1(net531),
    .A2(net151));
 sg13g2_nor2_1 _15760_ (.A(_09779_),
    .B(_09791_),
    .Y(_09995_));
 sg13g2_nor4_2 _15761_ (.A(net1056),
    .B(_08474_),
    .C(_09638_),
    .Y(_09996_),
    .D(_09793_));
 sg13g2_nor3_1 _15762_ (.A(\top_ihp.oisc.decoder.instruction[12] ),
    .B(_08474_),
    .C(_09638_),
    .Y(_09997_));
 sg13g2_nor3_1 _15763_ (.A(_08474_),
    .B(_09793_),
    .C(_09997_),
    .Y(_09998_));
 sg13g2_and2_1 _15764_ (.A(_09770_),
    .B(_09998_),
    .X(_09999_));
 sg13g2_a21o_1 _15765_ (.A2(_09996_),
    .A1(_09995_),
    .B1(_09999_),
    .X(_10000_));
 sg13g2_buf_8 _15766_ (.A(_10000_),
    .X(_10001_));
 sg13g2_a21oi_1 _15767_ (.A1(_09657_),
    .A2(_09651_),
    .Y(_10002_),
    .B1(_10001_));
 sg13g2_o21ai_1 _15768_ (.B1(_09734_),
    .Y(_10003_),
    .A1(net948),
    .A2(_10002_));
 sg13g2_a21oi_1 _15769_ (.A1(_08226_),
    .A2(_08230_),
    .Y(_10004_),
    .B1(_08239_));
 sg13g2_xnor2_1 _15770_ (.Y(_10005_),
    .A(_08022_),
    .B(_10004_));
 sg13g2_o21ai_1 _15771_ (.B1(net949),
    .Y(_10006_),
    .A1(_10003_),
    .A2(_10005_));
 sg13g2_a21oi_1 _15772_ (.A1(net1069),
    .A2(_10005_),
    .Y(_10007_),
    .B1(net921));
 sg13g2_or2_1 _15773_ (.X(_10008_),
    .B(_09896_),
    .A(_00200_));
 sg13g2_buf_1 _15774_ (.A(_09893_),
    .X(_10009_));
 sg13g2_a21oi_1 _15775_ (.A1(\top_ihp.oisc.decoder.instruction[16] ),
    .A2(net912),
    .Y(_10010_),
    .B1(_09901_));
 sg13g2_nand3_1 _15776_ (.B(_10008_),
    .C(_10010_),
    .A(net996),
    .Y(_10011_));
 sg13g2_o21ai_1 _15777_ (.B1(_10011_),
    .Y(_10012_),
    .A1(_10003_),
    .A2(_10007_));
 sg13g2_a21o_1 _15778_ (.A2(_10006_),
    .A1(_08428_),
    .B1(_10012_),
    .X(_10013_));
 sg13g2_buf_2 _15779_ (.A(_10013_),
    .X(_10014_));
 sg13g2_buf_1 _15780_ (.A(_10014_),
    .X(_10015_));
 sg13g2_nand2_1 _15781_ (.Y(_10016_),
    .A(\top_ihp.oisc.regs[0][16] ),
    .B(net660));
 sg13g2_o21ai_1 _15782_ (.B1(_10016_),
    .Y(_00459_),
    .A1(net531),
    .A2(net150));
 sg13g2_o21ai_1 _15783_ (.B1(_08239_),
    .Y(_10017_),
    .A1(_08428_),
    .A2(net1066));
 sg13g2_nand3_1 _15784_ (.B(_08226_),
    .C(_08230_),
    .A(net1066),
    .Y(_10018_));
 sg13g2_nor3_1 _15785_ (.A(net1069),
    .B(_08225_),
    .C(_08063_),
    .Y(_10019_));
 sg13g2_a21oi_1 _15786_ (.A1(_08230_),
    .A2(_10019_),
    .Y(_10020_),
    .B1(_08066_));
 sg13g2_nand3_1 _15787_ (.B(_10018_),
    .C(_10020_),
    .A(_10017_),
    .Y(_10021_));
 sg13g2_xor2_1 _15788_ (.B(_10021_),
    .A(_08064_),
    .X(_10022_));
 sg13g2_nand2_1 _15789_ (.Y(_10023_),
    .A(_00118_),
    .B(net920));
 sg13g2_nand3_1 _15790_ (.B(net904),
    .C(_09611_),
    .A(_00119_),
    .Y(_10024_));
 sg13g2_inv_1 _15791_ (.Y(_10025_),
    .A(_00120_));
 sg13g2_a22oi_1 _15792_ (.Y(_10026_),
    .B1(net950),
    .B2(\top_ihp.wb_coproc.dat_o[17] ),
    .A2(_10025_),
    .A1(net1029));
 sg13g2_nand3_1 _15793_ (.B(net891),
    .C(_10026_),
    .A(net904),
    .Y(_10027_));
 sg13g2_nand4_1 _15794_ (.B(_10023_),
    .C(_10024_),
    .A(_08799_),
    .Y(_10028_),
    .D(_10027_));
 sg13g2_buf_1 _15795_ (.A(_10028_),
    .X(_10029_));
 sg13g2_nor2_1 _15796_ (.A(_09834_),
    .B(_10029_),
    .Y(_10030_));
 sg13g2_nor3_1 _15797_ (.A(net947),
    .B(_10001_),
    .C(_10030_),
    .Y(_10031_));
 sg13g2_a21oi_1 _15798_ (.A1(net947),
    .A2(_10022_),
    .Y(_10032_),
    .B1(_10031_));
 sg13g2_nand2_1 _15799_ (.Y(_10033_),
    .A(\top_ihp.oisc.decoder.instruction[17] ),
    .B(_09893_));
 sg13g2_o21ai_1 _15800_ (.B1(_10033_),
    .Y(_10034_),
    .A1(_00201_),
    .A2(_09896_));
 sg13g2_o21ai_1 _15801_ (.B1(net996),
    .Y(_10035_),
    .A1(_09901_),
    .A2(_10034_));
 sg13g2_o21ai_1 _15802_ (.B1(_10035_),
    .Y(_10036_),
    .A1(_08256_),
    .A2(net949));
 sg13g2_o21ai_1 _15803_ (.B1(_10036_),
    .Y(_10037_),
    .A1(net917),
    .A2(_10032_));
 sg13g2_buf_1 _15804_ (.A(_10037_),
    .X(_10038_));
 sg13g2_buf_2 _15805_ (.A(_10038_),
    .X(_10039_));
 sg13g2_buf_1 _15806_ (.A(net661),
    .X(_10040_));
 sg13g2_nand2_1 _15807_ (.Y(_10041_),
    .A(\top_ihp.oisc.regs[0][17] ),
    .B(net530));
 sg13g2_o21ai_1 _15808_ (.B1(_10041_),
    .Y(_00460_),
    .A1(net531),
    .A2(net328));
 sg13g2_nand2_1 _15809_ (.Y(_10042_),
    .A(_00121_),
    .B(net920));
 sg13g2_nand3_1 _15810_ (.B(net889),
    .C(_09611_),
    .A(_00122_),
    .Y(_10043_));
 sg13g2_inv_1 _15811_ (.Y(_10044_),
    .A(_00123_));
 sg13g2_a22oi_1 _15812_ (.Y(_10045_),
    .B1(net950),
    .B2(\top_ihp.wb_coproc.dat_o[18] ),
    .A2(_10044_),
    .A1(net1029));
 sg13g2_nand3_1 _15813_ (.B(_09614_),
    .C(_10045_),
    .A(net889),
    .Y(_10046_));
 sg13g2_and4_1 _15814_ (.A(_08799_),
    .B(_10042_),
    .C(_10043_),
    .D(_10046_),
    .X(_10047_));
 sg13g2_buf_8 _15815_ (.A(_10047_),
    .X(_10048_));
 sg13g2_a21oi_1 _15816_ (.A1(net945),
    .A2(_10048_),
    .Y(_10049_),
    .B1(_10001_));
 sg13g2_o21ai_1 _15817_ (.B1(_08150_),
    .Y(_10050_),
    .A1(_08145_),
    .A2(_09500_));
 sg13g2_a221oi_1 _15818_ (.B2(_10050_),
    .C1(_08026_),
    .B1(_08067_),
    .A1(_08256_),
    .Y(_10051_),
    .A2(_08006_));
 sg13g2_xor2_1 _15819_ (.B(_10051_),
    .A(_08244_),
    .X(_10052_));
 sg13g2_nor2_1 _15820_ (.A(net921),
    .B(_10052_),
    .Y(_10053_));
 sg13g2_a21oi_1 _15821_ (.A1(net921),
    .A2(_10049_),
    .Y(_10054_),
    .B1(_10053_));
 sg13g2_a21oi_1 _15822_ (.A1(\top_ihp.oisc.decoder.instruction[18] ),
    .A2(_09893_),
    .Y(_10055_),
    .B1(_09901_));
 sg13g2_o21ai_1 _15823_ (.B1(_10055_),
    .Y(_10056_),
    .A1(_00202_),
    .A2(_09896_));
 sg13g2_mux2_1 _15824_ (.A0(net1070),
    .A1(_10056_),
    .S(net996),
    .X(_10057_));
 sg13g2_o21ai_1 _15825_ (.B1(_10057_),
    .Y(_10058_),
    .A1(net917),
    .A2(_10054_));
 sg13g2_buf_1 _15826_ (.A(_10058_),
    .X(_10059_));
 sg13g2_buf_2 _15827_ (.A(_10059_),
    .X(_10060_));
 sg13g2_nand2_1 _15828_ (.Y(_10061_),
    .A(\top_ihp.oisc.regs[0][18] ),
    .B(net530));
 sg13g2_o21ai_1 _15829_ (.B1(_10061_),
    .Y(_00461_),
    .A1(_09757_),
    .A2(net327));
 sg13g2_buf_1 _15830_ (.A(net661),
    .X(_10062_));
 sg13g2_inv_1 _15831_ (.Y(_10063_),
    .A(_08071_));
 sg13g2_o21ai_1 _15832_ (.B1(_08243_),
    .Y(_10064_),
    .A1(_10063_),
    .A2(_10051_));
 sg13g2_xnor2_1 _15833_ (.Y(_10065_),
    .A(net1071),
    .B(_10064_));
 sg13g2_nand3_1 _15834_ (.B(_09973_),
    .C(_10065_),
    .A(_07999_),
    .Y(_10066_));
 sg13g2_a21oi_1 _15835_ (.A1(\top_ihp.oisc.decoder.instruction[19] ),
    .A2(_09893_),
    .Y(_10067_),
    .B1(_09901_));
 sg13g2_o21ai_1 _15836_ (.B1(_10067_),
    .Y(_10068_),
    .A1(_00203_),
    .A2(_09896_));
 sg13g2_nor2_1 _15837_ (.A(_00124_),
    .B(net904),
    .Y(_10069_));
 sg13g2_inv_1 _15838_ (.Y(_10070_),
    .A(_00126_));
 sg13g2_a22oi_1 _15839_ (.Y(_10071_),
    .B1(_08788_),
    .B2(\top_ihp.wb_coproc.dat_o[19] ),
    .A2(_10070_),
    .A1(_08785_));
 sg13g2_and4_1 _15840_ (.A(net1024),
    .B(_00125_),
    .C(_08777_),
    .D(_08781_),
    .X(_10072_));
 sg13g2_a221oi_1 _15841_ (.B2(_10071_),
    .C1(_10072_),
    .B1(_08784_),
    .A1(net1041),
    .Y(_10073_),
    .A2(_08371_));
 sg13g2_o21ai_1 _15842_ (.B1(_08799_),
    .Y(_10074_),
    .A1(_10069_),
    .A2(_10073_));
 sg13g2_buf_2 _15843_ (.A(_10074_),
    .X(_10075_));
 sg13g2_nand2_1 _15844_ (.Y(_10076_),
    .A(_09595_),
    .B(_09598_));
 sg13g2_a221oi_1 _15845_ (.B2(_09995_),
    .C1(_10076_),
    .B1(_09996_),
    .A1(_09770_),
    .Y(_10077_),
    .A2(_09998_));
 sg13g2_buf_1 _15846_ (.A(_10077_),
    .X(_10078_));
 sg13g2_o21ai_1 _15847_ (.B1(_10078_),
    .Y(_10079_),
    .A1(_09834_),
    .A2(_10075_));
 sg13g2_nand3_1 _15848_ (.B(_10068_),
    .C(_10079_),
    .A(_10066_),
    .Y(_10080_));
 sg13g2_nand3b_1 _15849_ (.B(net947),
    .C(_09595_),
    .Y(_10081_),
    .A_N(_10065_));
 sg13g2_a21oi_1 _15850_ (.A1(net949),
    .A2(_10081_),
    .Y(_10082_),
    .B1(_07999_));
 sg13g2_a21o_1 _15851_ (.A2(_10080_),
    .A1(net953),
    .B1(_10082_),
    .X(_10083_));
 sg13g2_buf_1 _15852_ (.A(_10083_),
    .X(_10084_));
 sg13g2_buf_2 _15853_ (.A(_10084_),
    .X(_10085_));
 sg13g2_nand2_1 _15854_ (.Y(_10086_),
    .A(\top_ihp.oisc.regs[0][19] ),
    .B(net530));
 sg13g2_o21ai_1 _15855_ (.B1(_10086_),
    .Y(_00462_),
    .A1(net529),
    .A2(net326));
 sg13g2_buf_1 _15856_ (.A(\top_ihp.oisc.decoder.instruction[21] ),
    .X(_10087_));
 sg13g2_and2_1 _15857_ (.A(net1027),
    .B(_09740_),
    .X(_10088_));
 sg13g2_a21oi_1 _15858_ (.A1(_09684_),
    .A2(_10087_),
    .Y(_10089_),
    .B1(_10088_));
 sg13g2_nor2_1 _15859_ (.A(_09761_),
    .B(_09675_),
    .Y(_10090_));
 sg13g2_nand2_1 _15860_ (.Y(_10091_),
    .A(_09740_),
    .B(_10090_));
 sg13g2_o21ai_1 _15861_ (.B1(_10091_),
    .Y(_10092_),
    .A1(net1025),
    .A2(_10089_));
 sg13g2_and2_1 _15862_ (.A(_09682_),
    .B(_09894_),
    .X(_10093_));
 sg13g2_buf_1 _15863_ (.A(_10093_),
    .X(_10094_));
 sg13g2_nand2_1 _15864_ (.Y(_10095_),
    .A(net989),
    .B(_10087_));
 sg13g2_o21ai_1 _15865_ (.B1(_10095_),
    .Y(_10096_),
    .A1(net989),
    .A2(_00196_));
 sg13g2_a221oi_1 _15866_ (.B2(_10096_),
    .C1(_09596_),
    .B1(_10094_),
    .A1(net1026),
    .Y(_10097_),
    .A2(_10092_));
 sg13g2_inv_1 _15867_ (.Y(_10098_),
    .A(_00159_));
 sg13g2_a22oi_1 _15868_ (.Y(_10099_),
    .B1(net919),
    .B2(\top_ihp.wb_coproc.dat_o[25] ),
    .A2(_10098_),
    .A1(net994));
 sg13g2_mux2_1 _15869_ (.A0(_00158_),
    .A1(_10099_),
    .S(net878),
    .X(_10100_));
 sg13g2_mux2_1 _15870_ (.A0(_00157_),
    .A1(_10100_),
    .S(net879),
    .X(_10101_));
 sg13g2_nor3_1 _15871_ (.A(net993),
    .B(_09644_),
    .C(_10101_),
    .Y(_10102_));
 sg13g2_and4_1 _15872_ (.A(_08799_),
    .B(_10023_),
    .C(_10024_),
    .D(_10027_),
    .X(_10103_));
 sg13g2_nand2_1 _15873_ (.Y(_10104_),
    .A(_09644_),
    .B(_10103_));
 sg13g2_nand3b_1 _15874_ (.B(_10104_),
    .C(net1030),
    .Y(_10105_),
    .A_N(_10102_));
 sg13g2_nor2_1 _15875_ (.A(_00133_),
    .B(_09608_),
    .Y(_10106_));
 sg13g2_inv_1 _15876_ (.Y(_10107_),
    .A(_00135_));
 sg13g2_a221oi_1 _15877_ (.B2(\top_ihp.wb_coproc.dat_o[9] ),
    .C1(net888),
    .B1(_09621_),
    .A1(net994),
    .Y(_10108_),
    .A2(_10107_));
 sg13g2_a221oi_1 _15878_ (.B2(_00134_),
    .C1(_10108_),
    .B1(net888),
    .A1(net992),
    .Y(_10109_),
    .A2(net905));
 sg13g2_o21ai_1 _15879_ (.B1(_08794_),
    .Y(_10110_),
    .A1(_10106_),
    .A2(_10109_));
 sg13g2_nand3_1 _15880_ (.B(_09659_),
    .C(_10110_),
    .A(net991),
    .Y(_10111_));
 sg13g2_a21o_1 _15881_ (.A2(_10111_),
    .A1(_10105_),
    .B1(net990),
    .X(_10112_));
 sg13g2_nand2_1 _15882_ (.Y(_10113_),
    .A(_00194_),
    .B(net877));
 sg13g2_inv_1 _15883_ (.Y(_10114_),
    .A(_00195_));
 sg13g2_a22oi_1 _15884_ (.Y(_10115_),
    .B1(net899),
    .B2(\top_ihp.wb_coproc.dat_o[1] ),
    .A2(_10114_),
    .A1(net951));
 sg13g2_nand2_1 _15885_ (.Y(_10116_),
    .A(net854),
    .B(_10115_));
 sg13g2_nand3_1 _15886_ (.B(_10113_),
    .C(_10116_),
    .A(net855),
    .Y(_10117_));
 sg13g2_o21ai_1 _15887_ (.B1(_10117_),
    .Y(_10118_),
    .A1(_00193_),
    .A2(net855));
 sg13g2_a22oi_1 _15888_ (.Y(_10119_),
    .B1(net987),
    .B2(_10118_),
    .A2(\top_ihp.wb_dati_uart[1] ),
    .A1(net1028));
 sg13g2_o21ai_1 _15889_ (.B1(_10119_),
    .Y(_10120_),
    .A1(net990),
    .A2(_09660_));
 sg13g2_and3_1 _15890_ (.X(_10121_),
    .A(net952),
    .B(_10112_),
    .C(_10120_));
 sg13g2_xnor2_1 _15891_ (.Y(_10122_),
    .A(_08079_),
    .B(_08453_));
 sg13g2_nor2_1 _15892_ (.A(net921),
    .B(_10122_),
    .Y(_10123_));
 sg13g2_nor3_1 _15893_ (.A(net985),
    .B(_10121_),
    .C(_10123_),
    .Y(_10124_));
 sg13g2_nor3_2 _15894_ (.A(net915),
    .B(_10097_),
    .C(_10124_),
    .Y(_10125_));
 sg13g2_a21oi_1 _15895_ (.A1(_08078_),
    .A2(net898),
    .Y(_10126_),
    .B1(_10125_));
 sg13g2_buf_2 _15896_ (.A(_10126_),
    .X(_10127_));
 sg13g2_buf_1 _15897_ (.A(net325),
    .X(_10128_));
 sg13g2_nand2_1 _15898_ (.Y(_10129_),
    .A(\top_ihp.oisc.regs[0][1] ),
    .B(net530));
 sg13g2_o21ai_1 _15899_ (.B1(_10129_),
    .Y(_00463_),
    .A1(net529),
    .A2(net149));
 sg13g2_a21oi_2 _15900_ (.B1(_09999_),
    .Y(_10130_),
    .A2(_09996_),
    .A1(_09995_));
 sg13g2_nand2b_1 _15901_ (.Y(_10131_),
    .B(net900),
    .A_N(_00142_));
 sg13g2_inv_1 _15902_ (.Y(_10132_),
    .A(_00144_));
 sg13g2_a221oi_1 _15903_ (.B2(\top_ihp.wb_coproc.dat_o[20] ),
    .C1(net877),
    .B1(net899),
    .A1(net951),
    .Y(_10133_),
    .A2(_10132_));
 sg13g2_a21oi_1 _15904_ (.A1(_00143_),
    .A2(net877),
    .Y(_10134_),
    .B1(_10133_));
 sg13g2_nand2_1 _15905_ (.Y(_10135_),
    .A(net855),
    .B(_10134_));
 sg13g2_a21oi_1 _15906_ (.A1(_10131_),
    .A2(_10135_),
    .Y(_10136_),
    .B1(net944));
 sg13g2_nand2_1 _15907_ (.Y(_10137_),
    .A(net986),
    .B(_10136_));
 sg13g2_a21oi_1 _15908_ (.A1(_10130_),
    .A2(_10137_),
    .Y(_10138_),
    .B1(net948));
 sg13g2_nor2_1 _15909_ (.A(_07993_),
    .B(_08003_),
    .Y(_10139_));
 sg13g2_o21ai_1 _15910_ (.B1(_08263_),
    .Y(_10140_),
    .A1(_10004_),
    .A2(_08246_));
 sg13g2_xnor2_1 _15911_ (.Y(_10141_),
    .A(_10139_),
    .B(_10140_));
 sg13g2_nor2_1 _15912_ (.A(net952),
    .B(_10141_),
    .Y(_10142_));
 sg13g2_nor3_1 _15913_ (.A(net917),
    .B(_10138_),
    .C(_10142_),
    .Y(_10143_));
 sg13g2_buf_2 _15914_ (.A(_10143_),
    .X(_10144_));
 sg13g2_nand2_1 _15915_ (.Y(_10145_),
    .A(_09685_),
    .B(_09762_));
 sg13g2_a21oi_1 _15916_ (.A1(_09851_),
    .A2(_10145_),
    .Y(_10146_),
    .B1(_09595_));
 sg13g2_buf_2 _15917_ (.A(_10146_),
    .X(_10147_));
 sg13g2_nand2_1 _15918_ (.Y(_10148_),
    .A(_09681_),
    .B(_10009_));
 sg13g2_a21oi_1 _15919_ (.A1(_10147_),
    .A2(_10148_),
    .Y(_10149_),
    .B1(_09863_));
 sg13g2_a21oi_1 _15920_ (.A1(_07990_),
    .A2(net898),
    .Y(_10150_),
    .B1(_10149_));
 sg13g2_or2_1 _15921_ (.X(_10151_),
    .B(_10150_),
    .A(_10144_));
 sg13g2_buf_2 _15922_ (.A(_10151_),
    .X(_10152_));
 sg13g2_buf_8 _15923_ (.A(_10152_),
    .X(_10153_));
 sg13g2_nand2_1 _15924_ (.Y(_10154_),
    .A(\top_ihp.oisc.regs[0][20] ),
    .B(net530));
 sg13g2_o21ai_1 _15925_ (.B1(_10154_),
    .Y(_00464_),
    .A1(net529),
    .A2(net324));
 sg13g2_nand2_1 _15926_ (.Y(_10155_),
    .A(_10087_),
    .B(_09893_));
 sg13g2_nand2b_1 _15927_ (.Y(_10156_),
    .B(net900),
    .A_N(_00145_));
 sg13g2_inv_1 _15928_ (.Y(_10157_),
    .A(_00147_));
 sg13g2_a221oi_1 _15929_ (.B2(\top_ihp.wb_coproc.dat_o[21] ),
    .C1(net877),
    .B1(_09622_),
    .A1(net951),
    .Y(_10158_),
    .A2(_10157_));
 sg13g2_a21oi_1 _15930_ (.A1(_00146_),
    .A2(_09632_),
    .Y(_10159_),
    .B1(_10158_));
 sg13g2_nand2_1 _15931_ (.Y(_10160_),
    .A(net855),
    .B(_10159_));
 sg13g2_a21oi_2 _15932_ (.B1(net944),
    .Y(_10161_),
    .A2(_10160_),
    .A1(_10156_));
 sg13g2_nand2_1 _15933_ (.Y(_10162_),
    .A(net986),
    .B(_10161_));
 sg13g2_a221oi_1 _15934_ (.B2(_10078_),
    .C1(net946),
    .B1(_10162_),
    .A1(_10147_),
    .Y(_10163_),
    .A2(_10155_));
 sg13g2_xnor2_1 _15935_ (.Y(_10164_),
    .A(_08153_),
    .B(_08464_));
 sg13g2_o21ai_1 _15936_ (.B1(_09973_),
    .Y(_10165_),
    .A1(net1060),
    .A2(_10164_));
 sg13g2_a21o_1 _15937_ (.A2(_10164_),
    .A1(_10163_),
    .B1(net916),
    .X(_10166_));
 sg13g2_a22oi_1 _15938_ (.Y(_10167_),
    .B1(_10166_),
    .B2(net1060),
    .A2(_10165_),
    .A1(_10163_));
 sg13g2_buf_1 _15939_ (.A(_10167_),
    .X(_10168_));
 sg13g2_buf_2 _15940_ (.A(_10168_),
    .X(_10169_));
 sg13g2_nand2_1 _15941_ (.Y(_10170_),
    .A(\top_ihp.oisc.regs[0][21] ),
    .B(net530));
 sg13g2_o21ai_1 _15942_ (.B1(_10170_),
    .Y(_00465_),
    .A1(net529),
    .A2(net323));
 sg13g2_a21o_1 _15943_ (.A2(_08266_),
    .A1(_08464_),
    .B1(_08248_),
    .X(_10171_));
 sg13g2_xnor2_1 _15944_ (.Y(_10172_),
    .A(_08318_),
    .B(_10171_));
 sg13g2_nand2b_1 _15945_ (.Y(_10173_),
    .B(net900),
    .A_N(_00148_));
 sg13g2_nand2_1 _15946_ (.Y(_10174_),
    .A(_00149_),
    .B(_09632_));
 sg13g2_inv_1 _15947_ (.Y(_10175_),
    .A(_00150_));
 sg13g2_a22oi_1 _15948_ (.Y(_10176_),
    .B1(_09622_),
    .B2(\top_ihp.wb_coproc.dat_o[22] ),
    .A2(_10175_),
    .A1(_09618_));
 sg13g2_nand2_1 _15949_ (.Y(_10177_),
    .A(_09615_),
    .B(_10176_));
 sg13g2_nand3_1 _15950_ (.B(_10174_),
    .C(_10177_),
    .A(net855),
    .Y(_10178_));
 sg13g2_a21oi_1 _15951_ (.A1(_10173_),
    .A2(_10178_),
    .Y(_10179_),
    .B1(net944));
 sg13g2_nand2_1 _15952_ (.Y(_10180_),
    .A(net1042),
    .B(_10179_));
 sg13g2_a21oi_1 _15953_ (.A1(_10130_),
    .A2(_10180_),
    .Y(_10181_),
    .B1(net988));
 sg13g2_a21oi_1 _15954_ (.A1(net948),
    .A2(_10172_),
    .Y(_10182_),
    .B1(_10181_));
 sg13g2_buf_1 _15955_ (.A(\top_ihp.oisc.decoder.instruction[22] ),
    .X(_10183_));
 sg13g2_nand2_1 _15956_ (.Y(_10184_),
    .A(_10183_),
    .B(net912));
 sg13g2_a221oi_1 _15957_ (.B2(_10147_),
    .C1(net916),
    .B1(_10184_),
    .A1(net995),
    .Y(_10185_),
    .A2(_10182_));
 sg13g2_buf_2 _15958_ (.A(_10185_),
    .X(_10186_));
 sg13g2_a21oi_1 _15959_ (.A1(_08160_),
    .A2(net898),
    .Y(_10187_),
    .B1(_10186_));
 sg13g2_buf_2 _15960_ (.A(_10187_),
    .X(_10188_));
 sg13g2_buf_8 _15961_ (.A(net322),
    .X(_10189_));
 sg13g2_nand2_1 _15962_ (.Y(_10190_),
    .A(\top_ihp.oisc.regs[0][22] ),
    .B(net530));
 sg13g2_o21ai_1 _15963_ (.B1(_10190_),
    .Y(_00466_),
    .A1(net529),
    .A2(net148));
 sg13g2_a21oi_1 _15964_ (.A1(_08391_),
    .A2(_08435_),
    .Y(_10191_),
    .B1(_08397_));
 sg13g2_xnor2_1 _15965_ (.Y(_10192_),
    .A(_08319_),
    .B(_10191_));
 sg13g2_o21ai_1 _15966_ (.B1(_10130_),
    .Y(_10193_),
    .A1(_09834_),
    .A2(_09777_));
 sg13g2_mux2_1 _15967_ (.A0(_10192_),
    .A1(_10193_),
    .S(net921),
    .X(_10194_));
 sg13g2_buf_1 _15968_ (.A(_10194_),
    .X(_10195_));
 sg13g2_buf_1 _15969_ (.A(\top_ihp.oisc.decoder.instruction[23] ),
    .X(_10196_));
 sg13g2_a21o_1 _15970_ (.A2(_10145_),
    .A1(_09851_),
    .B1(_09595_),
    .X(_10197_));
 sg13g2_buf_1 _15971_ (.A(_10197_),
    .X(_10198_));
 sg13g2_a21oi_1 _15972_ (.A1(_10196_),
    .A2(net912),
    .Y(_10199_),
    .B1(_10198_));
 sg13g2_nor2_1 _15973_ (.A(net1061),
    .B(net949),
    .Y(_10200_));
 sg13g2_a21oi_1 _15974_ (.A1(net953),
    .A2(_10199_),
    .Y(_10201_),
    .B1(_10200_));
 sg13g2_o21ai_1 _15975_ (.B1(_10201_),
    .Y(_10202_),
    .A1(net917),
    .A2(_10195_));
 sg13g2_buf_1 _15976_ (.A(_10202_),
    .X(_10203_));
 sg13g2_buf_8 _15977_ (.A(net528),
    .X(_10204_));
 sg13g2_nand2_1 _15978_ (.Y(_10205_),
    .A(\top_ihp.oisc.regs[0][23] ),
    .B(_10040_));
 sg13g2_o21ai_1 _15979_ (.B1(_10205_),
    .Y(_00467_),
    .A1(_10062_),
    .A2(net321));
 sg13g2_nand2_1 _15980_ (.Y(_10206_),
    .A(net945),
    .B(_09628_));
 sg13g2_nor2_1 _15981_ (.A(net988),
    .B(_10001_),
    .Y(_10207_));
 sg13g2_nand2_1 _15982_ (.Y(_10208_),
    .A(_08253_),
    .B(_08275_));
 sg13g2_xnor2_1 _15983_ (.Y(_10209_),
    .A(_08280_),
    .B(_10208_));
 sg13g2_a22oi_1 _15984_ (.Y(_10210_),
    .B1(_10209_),
    .B2(net947),
    .A2(_10207_),
    .A1(_10206_));
 sg13g2_buf_1 _15985_ (.A(\top_ihp.oisc.decoder.instruction[24] ),
    .X(_10211_));
 sg13g2_a21oi_1 _15986_ (.A1(_10211_),
    .A2(net912),
    .Y(_10212_),
    .B1(_10198_));
 sg13g2_nand2_1 _15987_ (.Y(_10213_),
    .A(_08154_),
    .B(net946));
 sg13g2_o21ai_1 _15988_ (.B1(_10213_),
    .Y(_10214_),
    .A1(_09865_),
    .A2(_10212_));
 sg13g2_o21ai_1 _15989_ (.B1(_10214_),
    .Y(_10215_),
    .A1(net917),
    .A2(_10210_));
 sg13g2_buf_2 _15990_ (.A(_10215_),
    .X(_10216_));
 sg13g2_buf_1 _15991_ (.A(_10216_),
    .X(_10217_));
 sg13g2_nand2_1 _15992_ (.Y(_10218_),
    .A(\top_ihp.oisc.regs[0][24] ),
    .B(_10040_));
 sg13g2_o21ai_1 _15993_ (.B1(_10218_),
    .Y(_00468_),
    .A1(_10062_),
    .A2(net320));
 sg13g2_nand2_1 _15994_ (.Y(_10219_),
    .A(_08379_),
    .B(_08391_));
 sg13g2_inv_1 _15995_ (.Y(_10220_),
    .A(_08164_));
 sg13g2_o21ai_1 _15996_ (.B1(_08178_),
    .Y(_10221_),
    .A1(_08164_),
    .A2(_08395_));
 sg13g2_o21ai_1 _15997_ (.B1(_10221_),
    .Y(_10222_),
    .A1(_10220_),
    .A2(_08396_));
 sg13g2_nand2b_1 _15998_ (.Y(_10223_),
    .B(_08154_),
    .A_N(_08155_));
 sg13g2_o21ai_1 _15999_ (.B1(_10223_),
    .Y(_10224_),
    .A1(_08172_),
    .A2(_10222_));
 sg13g2_o21ai_1 _16000_ (.B1(_10224_),
    .Y(_10225_),
    .A1(_08464_),
    .A2(_10219_));
 sg13g2_xnor2_1 _16001_ (.Y(_10226_),
    .A(_08159_),
    .B(_10225_));
 sg13g2_nor2_1 _16002_ (.A(_09627_),
    .B(_10101_),
    .Y(_10227_));
 sg13g2_nand2_1 _16003_ (.Y(_10228_),
    .A(net990),
    .B(_10227_));
 sg13g2_a21oi_1 _16004_ (.A1(_10130_),
    .A2(_10228_),
    .Y(_10229_),
    .B1(net988));
 sg13g2_a21oi_1 _16005_ (.A1(net948),
    .A2(_10226_),
    .Y(_10230_),
    .B1(_10229_));
 sg13g2_buf_1 _16006_ (.A(\top_ihp.oisc.decoder.instruction[25] ),
    .X(_10231_));
 sg13g2_nand2_1 _16007_ (.Y(_10232_),
    .A(_10231_),
    .B(net912));
 sg13g2_a221oi_1 _16008_ (.B2(_10147_),
    .C1(net916),
    .B1(_10232_),
    .A1(net995),
    .Y(_10233_),
    .A2(_10230_));
 sg13g2_buf_1 _16009_ (.A(_10233_),
    .X(_10234_));
 sg13g2_a21oi_1 _16010_ (.A1(_08157_),
    .A2(net898),
    .Y(_10235_),
    .B1(_10234_));
 sg13g2_buf_2 _16011_ (.A(_10235_),
    .X(_10236_));
 sg13g2_buf_1 _16012_ (.A(net319),
    .X(_10237_));
 sg13g2_nand2_1 _16013_ (.Y(_10238_),
    .A(\top_ihp.oisc.regs[0][25] ),
    .B(net530));
 sg13g2_o21ai_1 _16014_ (.B1(_10238_),
    .Y(_00469_),
    .A1(net529),
    .A2(net147));
 sg13g2_a21oi_1 _16015_ (.A1(net945),
    .A2(_09812_),
    .Y(_10239_),
    .B1(_10001_));
 sg13g2_xnor2_1 _16016_ (.Y(_10240_),
    .A(_08188_),
    .B(_08282_));
 sg13g2_mux2_1 _16017_ (.A0(_10239_),
    .A1(_10240_),
    .S(net948),
    .X(_10241_));
 sg13g2_nand2_1 _16018_ (.Y(_10242_),
    .A(net995),
    .B(_10241_));
 sg13g2_buf_1 _16019_ (.A(\top_ihp.oisc.decoder.instruction[26] ),
    .X(_10243_));
 sg13g2_nand2_1 _16020_ (.Y(_10244_),
    .A(_10243_),
    .B(net912));
 sg13g2_a21oi_1 _16021_ (.A1(_10147_),
    .A2(_10244_),
    .Y(_10245_),
    .B1(net915));
 sg13g2_a22oi_1 _16022_ (.Y(_10246_),
    .B1(_10242_),
    .B2(_10245_),
    .A2(_09864_),
    .A1(net1048));
 sg13g2_buf_1 _16023_ (.A(_10246_),
    .X(_10247_));
 sg13g2_buf_2 _16024_ (.A(_10247_),
    .X(_10248_));
 sg13g2_buf_8 _16025_ (.A(net661),
    .X(_10249_));
 sg13g2_nand2_1 _16026_ (.Y(_10250_),
    .A(\top_ihp.oisc.regs[0][26] ),
    .B(net527));
 sg13g2_o21ai_1 _16027_ (.B1(_10250_),
    .Y(_00470_),
    .A1(net529),
    .A2(net146));
 sg13g2_xnor2_1 _16028_ (.Y(_10251_),
    .A(_08465_),
    .B(_08446_));
 sg13g2_nor2_1 _16029_ (.A(_09834_),
    .B(_09841_),
    .Y(_10252_));
 sg13g2_nor3_1 _16030_ (.A(_09848_),
    .B(_10001_),
    .C(_10252_),
    .Y(_10253_));
 sg13g2_a21oi_1 _16031_ (.A1(net947),
    .A2(_10251_),
    .Y(_10254_),
    .B1(_10253_));
 sg13g2_a21oi_1 _16032_ (.A1(\top_ihp.oisc.decoder.instruction[27] ),
    .A2(net912),
    .Y(_10255_),
    .B1(_10198_));
 sg13g2_nand2_1 _16033_ (.Y(_10256_),
    .A(net1044),
    .B(net946));
 sg13g2_o21ai_1 _16034_ (.B1(_10256_),
    .Y(_10257_),
    .A1(net916),
    .A2(_10255_));
 sg13g2_o21ai_1 _16035_ (.B1(_10257_),
    .Y(_10258_),
    .A1(net917),
    .A2(_10254_));
 sg13g2_buf_1 _16036_ (.A(_10258_),
    .X(_10259_));
 sg13g2_buf_2 _16037_ (.A(_10259_),
    .X(_10260_));
 sg13g2_nand2_1 _16038_ (.Y(_10261_),
    .A(\top_ihp.oisc.regs[0][27] ),
    .B(net527));
 sg13g2_o21ai_1 _16039_ (.B1(_10261_),
    .Y(_00471_),
    .A1(net529),
    .A2(net318));
 sg13g2_buf_1 _16040_ (.A(net661),
    .X(_10262_));
 sg13g2_nand2_1 _16041_ (.Y(_10263_),
    .A(_08301_),
    .B(_09973_));
 sg13g2_nand2_1 _16042_ (.Y(_10264_),
    .A(\top_ihp.oisc.decoder.instruction[28] ),
    .B(_10009_));
 sg13g2_nand2_1 _16043_ (.Y(_10265_),
    .A(net945),
    .B(_09882_));
 sg13g2_a221oi_1 _16044_ (.B2(_10078_),
    .C1(net915),
    .B1(_10265_),
    .A1(_10147_),
    .Y(_10266_),
    .A2(_10264_));
 sg13g2_a22oi_1 _16045_ (.Y(_10267_),
    .B1(_10263_),
    .B2(_10266_),
    .A2(net898),
    .A1(net1057));
 sg13g2_buf_1 _16046_ (.A(_10267_),
    .X(_10268_));
 sg13g2_buf_2 _16047_ (.A(_10268_),
    .X(_10269_));
 sg13g2_nand2_1 _16048_ (.Y(_10270_),
    .A(\top_ihp.oisc.regs[0][28] ),
    .B(net527));
 sg13g2_o21ai_1 _16049_ (.B1(_10270_),
    .Y(_00472_),
    .A1(net526),
    .A2(net525));
 sg13g2_xnor2_1 _16050_ (.Y(_10271_),
    .A(_08321_),
    .B(_08472_));
 sg13g2_nor3_1 _16051_ (.A(_09820_),
    .B(_09600_),
    .C(_10271_),
    .Y(_10272_));
 sg13g2_nor2_1 _16052_ (.A(net915),
    .B(_10272_),
    .Y(_10273_));
 sg13g2_nand2_1 _16053_ (.Y(_10274_),
    .A(net945),
    .B(_09923_));
 sg13g2_nand2_1 _16054_ (.Y(_10275_),
    .A(\top_ihp.oisc.decoder.instruction[29] ),
    .B(net912));
 sg13g2_a22oi_1 _16055_ (.Y(_10276_),
    .B1(_10275_),
    .B2(_10147_),
    .A2(_10274_),
    .A1(_10078_));
 sg13g2_nand3_1 _16056_ (.B(_09973_),
    .C(_10271_),
    .A(_08320_),
    .Y(_10277_));
 sg13g2_a21o_1 _16057_ (.A2(_10277_),
    .A1(_10276_),
    .B1(net916),
    .X(_10278_));
 sg13g2_o21ai_1 _16058_ (.B1(_10278_),
    .Y(_10279_),
    .A1(_08320_),
    .A2(_10273_));
 sg13g2_buf_2 _16059_ (.A(_10279_),
    .X(_10280_));
 sg13g2_buf_1 _16060_ (.A(_10280_),
    .X(_10281_));
 sg13g2_nand2_1 _16061_ (.Y(_10282_),
    .A(\top_ihp.oisc.regs[0][29] ),
    .B(_10249_));
 sg13g2_o21ai_1 _16062_ (.B1(_10282_),
    .Y(_00473_),
    .A1(_10262_),
    .A2(net317));
 sg13g2_inv_1 _16063_ (.Y(_10283_),
    .A(_00096_));
 sg13g2_a22oi_1 _16064_ (.Y(_10284_),
    .B1(_09620_),
    .B2(\top_ihp.wb_coproc.dat_o[2] ),
    .A2(_10283_),
    .A1(_09616_));
 sg13g2_mux2_1 _16065_ (.A0(_00095_),
    .A1(_10284_),
    .S(net878),
    .X(_10285_));
 sg13g2_nand2b_1 _16066_ (.Y(_10286_),
    .B(net920),
    .A_N(_00094_));
 sg13g2_o21ai_1 _16067_ (.B1(_10286_),
    .Y(_10287_),
    .A1(_09604_),
    .A2(_10285_));
 sg13g2_and2_1 _16068_ (.A(net1028),
    .B(\top_ihp.wb_dati_uart[2] ),
    .X(_10288_));
 sg13g2_buf_1 _16069_ (.A(_10288_),
    .X(_10289_));
 sg13g2_a21oi_1 _16070_ (.A1(net987),
    .A2(_10287_),
    .Y(_10290_),
    .B1(_10289_));
 sg13g2_buf_2 _16071_ (.A(_10290_),
    .X(_10291_));
 sg13g2_nand2_1 _16072_ (.Y(_10292_),
    .A(_09654_),
    .B(_10048_));
 sg13g2_o21ai_1 _16073_ (.B1(_10292_),
    .Y(_10293_),
    .A1(net1030),
    .A2(_10291_));
 sg13g2_mux2_1 _16074_ (.A0(_09805_),
    .A1(_09812_),
    .S(_09601_),
    .X(_10294_));
 sg13g2_nor2_1 _16075_ (.A(_09834_),
    .B(_10291_),
    .Y(_10295_));
 sg13g2_a221oi_1 _16076_ (.B2(_09641_),
    .C1(_10295_),
    .B1(_10294_),
    .A1(_09644_),
    .Y(_10296_),
    .A2(_10293_));
 sg13g2_nand2_1 _16077_ (.Y(_10297_),
    .A(_08080_),
    .B(_08084_));
 sg13g2_o21ai_1 _16078_ (.B1(_08079_),
    .Y(_10298_),
    .A1(_08080_),
    .A2(_08084_));
 sg13g2_nand2_1 _16079_ (.Y(_10299_),
    .A(_10297_),
    .B(_10298_));
 sg13g2_xnor2_1 _16080_ (.Y(_10300_),
    .A(_09501_),
    .B(_10299_));
 sg13g2_nor2_1 _16081_ (.A(net952),
    .B(_10300_),
    .Y(_10301_));
 sg13g2_a21oi_1 _16082_ (.A1(net952),
    .A2(_10296_),
    .Y(_10302_),
    .B1(_10301_));
 sg13g2_and2_1 _16083_ (.A(net1027),
    .B(_09715_),
    .X(_10303_));
 sg13g2_a21oi_1 _16084_ (.A1(_09684_),
    .A2(_10183_),
    .Y(_10304_),
    .B1(_10303_));
 sg13g2_nand2_1 _16085_ (.Y(_10305_),
    .A(_09715_),
    .B(_10090_));
 sg13g2_o21ai_1 _16086_ (.B1(_10305_),
    .Y(_10306_),
    .A1(net1025),
    .A2(_10304_));
 sg13g2_nand2_1 _16087_ (.Y(_10307_),
    .A(net989),
    .B(_10183_));
 sg13g2_o21ai_1 _16088_ (.B1(_10307_),
    .Y(_10308_),
    .A1(net989),
    .A2(_00197_));
 sg13g2_a22oi_1 _16089_ (.Y(_10309_),
    .B1(_10308_),
    .B2(_10094_),
    .A2(_10306_),
    .A1(net1026));
 sg13g2_nand2_1 _16090_ (.Y(_10310_),
    .A(net1022),
    .B(_10309_));
 sg13g2_o21ai_1 _16091_ (.B1(_10310_),
    .Y(_10311_),
    .A1(_09849_),
    .A2(_10302_));
 sg13g2_nor2_1 _16092_ (.A(net915),
    .B(_10311_),
    .Y(_10312_));
 sg13g2_a21oi_1 _16093_ (.A1(_08090_),
    .A2(_09864_),
    .Y(_10313_),
    .B1(_10312_));
 sg13g2_buf_2 _16094_ (.A(_10313_),
    .X(_10314_));
 sg13g2_buf_2 _16095_ (.A(_10314_),
    .X(_10315_));
 sg13g2_nand2_1 _16096_ (.Y(_10316_),
    .A(\top_ihp.oisc.regs[0][2] ),
    .B(_10249_));
 sg13g2_o21ai_1 _16097_ (.B1(_10316_),
    .Y(_00474_),
    .A1(net526),
    .A2(net145));
 sg13g2_xnor2_1 _16098_ (.Y(_10317_),
    .A(_08315_),
    .B(_08351_));
 sg13g2_a21oi_1 _16099_ (.A1(_10317_),
    .A2(_09973_),
    .Y(_10318_),
    .B1(net916));
 sg13g2_nand2_1 _16100_ (.Y(_10319_),
    .A(net1043),
    .B(_09973_));
 sg13g2_nand2_1 _16101_ (.Y(_10320_),
    .A(net986),
    .B(_09956_));
 sg13g2_nand2_1 _16102_ (.Y(_10321_),
    .A(\top_ihp.oisc.decoder.instruction[30] ),
    .B(_09893_));
 sg13g2_a22oi_1 _16103_ (.Y(_10322_),
    .B1(_10321_),
    .B2(_10147_),
    .A2(_10320_),
    .A1(_10078_));
 sg13g2_o21ai_1 _16104_ (.B1(_10322_),
    .Y(_10323_),
    .A1(_10317_),
    .A2(_10319_));
 sg13g2_nand2_1 _16105_ (.Y(_10324_),
    .A(_09693_),
    .B(_10323_));
 sg13g2_o21ai_1 _16106_ (.B1(_10324_),
    .Y(_10325_),
    .A1(net1043),
    .A2(_10318_));
 sg13g2_buf_2 _16107_ (.A(_10325_),
    .X(_10326_));
 sg13g2_buf_2 _16108_ (.A(_10326_),
    .X(_10327_));
 sg13g2_nand2_1 _16109_ (.Y(_10328_),
    .A(\top_ihp.oisc.regs[0][30] ),
    .B(net527));
 sg13g2_o21ai_1 _16110_ (.B1(_10328_),
    .Y(_00475_),
    .A1(net526),
    .A2(net144));
 sg13g2_xnor2_1 _16111_ (.Y(_10329_),
    .A(_09498_),
    .B(_09497_));
 sg13g2_buf_1 _16112_ (.A(_10329_),
    .X(_10330_));
 sg13g2_nand2_1 _16113_ (.Y(_10331_),
    .A(_10330_),
    .B(_09707_));
 sg13g2_nand2_1 _16114_ (.Y(_10332_),
    .A(_09503_),
    .B(net988));
 sg13g2_nand2_1 _16115_ (.Y(_10333_),
    .A(_08306_),
    .B(_08349_));
 sg13g2_nor4_1 _16116_ (.A(_08340_),
    .B(_08343_),
    .C(_08347_),
    .D(_10333_),
    .Y(_10334_));
 sg13g2_a21oi_1 _16117_ (.A1(_08326_),
    .A2(_10334_),
    .Y(_10335_),
    .B1(_08315_));
 sg13g2_a21oi_1 _16118_ (.A1(_08311_),
    .A2(_08351_),
    .Y(_10336_),
    .B1(_10335_));
 sg13g2_mux2_1 _16119_ (.A0(_10331_),
    .A1(_10332_),
    .S(_10336_),
    .X(_10337_));
 sg13g2_mux2_1 _16120_ (.A0(_00172_),
    .A1(_09768_),
    .S(_09609_),
    .X(_10338_));
 sg13g2_nor2_1 _16121_ (.A(_09909_),
    .B(_10338_),
    .Y(_10339_));
 sg13g2_nand2_1 _16122_ (.Y(_10340_),
    .A(_09657_),
    .B(_10339_));
 sg13g2_a21oi_1 _16123_ (.A1(_10207_),
    .A2(_10340_),
    .Y(_10341_),
    .B1(net1022));
 sg13g2_a21oi_1 _16124_ (.A1(_09761_),
    .A2(_09700_),
    .Y(_10342_),
    .B1(_09678_));
 sg13g2_nor2b_1 _16125_ (.A(_10342_),
    .B_N(_09851_),
    .Y(_10343_));
 sg13g2_a221oi_1 _16126_ (.B2(net1022),
    .C1(_09856_),
    .B1(_10343_),
    .A1(_10337_),
    .Y(_10344_),
    .A2(_10341_));
 sg13g2_buf_2 _16127_ (.A(_10344_),
    .X(_10345_));
 sg13g2_nor2_1 _16128_ (.A(_09497_),
    .B(_09593_),
    .Y(_10346_));
 sg13g2_or2_1 _16129_ (.X(_10347_),
    .B(_10346_),
    .A(_10345_));
 sg13g2_buf_8 _16130_ (.A(_10347_),
    .X(_10348_));
 sg13g2_buf_8 _16131_ (.A(_10348_),
    .X(_10349_));
 sg13g2_nand2_1 _16132_ (.Y(_10350_),
    .A(\top_ihp.oisc.regs[0][31] ),
    .B(net527));
 sg13g2_o21ai_1 _16133_ (.B1(_10350_),
    .Y(_00476_),
    .A1(net526),
    .A2(net52));
 sg13g2_nand2_1 _16134_ (.Y(_10351_),
    .A(net1028),
    .B(\top_ihp.wb_dati_uart[3] ));
 sg13g2_nor2_1 _16135_ (.A(_00100_),
    .B(net889),
    .Y(_10352_));
 sg13g2_inv_1 _16136_ (.Y(_10353_),
    .A(_00102_));
 sg13g2_a22oi_1 _16137_ (.Y(_10354_),
    .B1(net919),
    .B2(\top_ihp.wb_coproc.dat_o[3] ),
    .A2(_10353_),
    .A1(net994));
 sg13g2_and4_1 _16138_ (.A(net1024),
    .B(_00101_),
    .C(net914),
    .D(net913),
    .X(_10355_));
 sg13g2_a221oi_1 _16139_ (.B2(_10354_),
    .C1(_10355_),
    .B1(net878),
    .A1(net1041),
    .Y(_10356_),
    .A2(net905));
 sg13g2_o21ai_1 _16140_ (.B1(net987),
    .Y(_10357_),
    .A1(_10352_),
    .A2(_10356_));
 sg13g2_nand2_1 _16141_ (.Y(_10358_),
    .A(_10351_),
    .B(_10357_));
 sg13g2_buf_2 _16142_ (.A(_10358_),
    .X(_10359_));
 sg13g2_nand2_1 _16143_ (.Y(_10360_),
    .A(_09653_),
    .B(_10359_));
 sg13g2_o21ai_1 _16144_ (.B1(_10360_),
    .Y(_10361_),
    .A1(_09835_),
    .A2(_10075_));
 sg13g2_or2_1 _16145_ (.X(_10362_),
    .B(_09841_),
    .A(_09653_));
 sg13g2_nand2_1 _16146_ (.Y(_10363_),
    .A(_09638_),
    .B(_09639_));
 sg13g2_a21oi_1 _16147_ (.A1(_09842_),
    .A2(_10362_),
    .Y(_10364_),
    .B1(_10363_));
 sg13g2_a221oi_1 _16148_ (.B2(_09644_),
    .C1(_10364_),
    .B1(_10361_),
    .A1(_09798_),
    .Y(_10365_),
    .A2(_10359_));
 sg13g2_o21ai_1 _16149_ (.B1(_08095_),
    .Y(_10366_),
    .A1(_08092_),
    .A2(_10299_));
 sg13g2_xnor2_1 _16150_ (.Y(_10367_),
    .A(_09502_),
    .B(_10366_));
 sg13g2_mux2_1 _16151_ (.A0(_10365_),
    .A1(_10367_),
    .S(net948),
    .X(_10368_));
 sg13g2_and2_1 _16152_ (.A(net1027),
    .B(_09712_),
    .X(_10369_));
 sg13g2_a21oi_1 _16153_ (.A1(_09684_),
    .A2(_10196_),
    .Y(_10370_),
    .B1(_10369_));
 sg13g2_nand2_1 _16154_ (.Y(_10371_),
    .A(_09712_),
    .B(_10090_));
 sg13g2_o21ai_1 _16155_ (.B1(_10371_),
    .Y(_10372_),
    .A1(net1025),
    .A2(_10370_));
 sg13g2_nand2_1 _16156_ (.Y(_10373_),
    .A(net989),
    .B(_10196_));
 sg13g2_o21ai_1 _16157_ (.B1(_10373_),
    .Y(_10374_),
    .A1(net989),
    .A2(_00198_));
 sg13g2_a22oi_1 _16158_ (.Y(_10375_),
    .B1(_10374_),
    .B2(_10094_),
    .A2(_10372_),
    .A1(net1026));
 sg13g2_nand2b_1 _16159_ (.Y(_10376_),
    .B(net985),
    .A_N(_10375_));
 sg13g2_o21ai_1 _16160_ (.B1(_10376_),
    .Y(_10377_),
    .A1(net985),
    .A2(_10368_));
 sg13g2_nor2b_1 _16161_ (.A(net949),
    .B_N(_08086_),
    .Y(_10378_));
 sg13g2_a21oi_1 _16162_ (.A1(net953),
    .A2(_10377_),
    .Y(_10379_),
    .B1(_10378_));
 sg13g2_buf_1 _16163_ (.A(_10379_),
    .X(_10380_));
 sg13g2_buf_2 _16164_ (.A(_10380_),
    .X(_10381_));
 sg13g2_nand2_1 _16165_ (.Y(_10382_),
    .A(\top_ihp.oisc.regs[0][3] ),
    .B(net527));
 sg13g2_o21ai_1 _16166_ (.B1(_10382_),
    .Y(_00477_),
    .A1(net526),
    .A2(net143));
 sg13g2_nand2_1 _16167_ (.Y(_10383_),
    .A(net1028),
    .B(\top_ihp.wb_dati_uart[4] ));
 sg13g2_nor2_1 _16168_ (.A(_00097_),
    .B(_09607_),
    .Y(_10384_));
 sg13g2_inv_1 _16169_ (.Y(_10385_),
    .A(_00099_));
 sg13g2_a22oi_1 _16170_ (.Y(_10386_),
    .B1(_09620_),
    .B2(\top_ihp.wb_coproc.dat_o[4] ),
    .A2(_10385_),
    .A1(_09616_));
 sg13g2_and4_1 _16171_ (.A(net1024),
    .B(_00098_),
    .C(net970),
    .D(net913),
    .X(_10387_));
 sg13g2_a221oi_1 _16172_ (.B2(_10386_),
    .C1(_10387_),
    .B1(net878),
    .A1(net1041),
    .Y(_10388_),
    .A2(net905));
 sg13g2_o21ai_1 _16173_ (.B1(net987),
    .Y(_10389_),
    .A1(_10384_),
    .A2(_10388_));
 sg13g2_buf_1 _16174_ (.A(_10389_),
    .X(_10390_));
 sg13g2_nand2_1 _16175_ (.Y(_10391_),
    .A(_10383_),
    .B(_10390_));
 sg13g2_buf_1 _16176_ (.A(_10391_),
    .X(_10392_));
 sg13g2_a22oi_1 _16177_ (.Y(_10393_),
    .B1(net765),
    .B2(net991),
    .A2(_10136_),
    .A1(net918));
 sg13g2_a21o_1 _16178_ (.A2(_09882_),
    .A1(_09602_),
    .B1(_09885_),
    .X(_10394_));
 sg13g2_a22oi_1 _16179_ (.Y(_10395_),
    .B1(_10394_),
    .B2(_09641_),
    .A2(net765),
    .A1(net990));
 sg13g2_o21ai_1 _16180_ (.B1(_10395_),
    .Y(_10396_),
    .A1(_09659_),
    .A2(_10393_));
 sg13g2_xnor2_1 _16181_ (.Y(_10397_),
    .A(_08110_),
    .B(_08099_));
 sg13g2_xnor2_1 _16182_ (.Y(_10398_),
    .A(_08109_),
    .B(_10397_));
 sg13g2_nor2_1 _16183_ (.A(_09599_),
    .B(_10398_),
    .Y(_10399_));
 sg13g2_a21oi_1 _16184_ (.A1(net921),
    .A2(_10396_),
    .Y(_10400_),
    .B1(_10399_));
 sg13g2_and2_1 _16185_ (.A(net1027),
    .B(_09730_),
    .X(_10401_));
 sg13g2_a21oi_1 _16186_ (.A1(_09684_),
    .A2(_10211_),
    .Y(_10402_),
    .B1(_10401_));
 sg13g2_nand2_1 _16187_ (.Y(_10403_),
    .A(_09730_),
    .B(_10090_));
 sg13g2_o21ai_1 _16188_ (.B1(_10403_),
    .Y(_10404_),
    .A1(_09689_),
    .A2(_10402_));
 sg13g2_nand2_1 _16189_ (.Y(_10405_),
    .A(net989),
    .B(_10211_));
 sg13g2_o21ai_1 _16190_ (.B1(_10405_),
    .Y(_10406_),
    .A1(net989),
    .A2(_00199_));
 sg13g2_a22oi_1 _16191_ (.Y(_10407_),
    .B1(_10406_),
    .B2(_10094_),
    .A2(_10404_),
    .A1(net1026));
 sg13g2_nand2b_1 _16192_ (.Y(_10408_),
    .B(net985),
    .A_N(_10407_));
 sg13g2_o21ai_1 _16193_ (.B1(_10408_),
    .Y(_10409_),
    .A1(net985),
    .A2(_10400_));
 sg13g2_nor2b_1 _16194_ (.A(_09693_),
    .B_N(_08109_),
    .Y(_10410_));
 sg13g2_a21oi_1 _16195_ (.A1(_09593_),
    .A2(_10409_),
    .Y(_10411_),
    .B1(_10410_));
 sg13g2_buf_1 _16196_ (.A(_10411_),
    .X(_10412_));
 sg13g2_buf_2 _16197_ (.A(_10412_),
    .X(_10413_));
 sg13g2_nand2_1 _16198_ (.Y(_10414_),
    .A(\top_ihp.oisc.regs[0][4] ),
    .B(net527));
 sg13g2_o21ai_1 _16199_ (.B1(_10414_),
    .Y(_00478_),
    .A1(net526),
    .A2(net142));
 sg13g2_o21ai_1 _16200_ (.B1(_08113_),
    .Y(_10415_),
    .A1(_08112_),
    .A2(_08099_));
 sg13g2_xnor2_1 _16201_ (.Y(_10416_),
    .A(_08127_),
    .B(_10415_));
 sg13g2_a21oi_1 _16202_ (.A1(_10231_),
    .A2(_09764_),
    .Y(_10417_),
    .B1(_09600_));
 sg13g2_a21oi_1 _16203_ (.A1(_10416_),
    .A2(_10417_),
    .Y(_10418_),
    .B1(net916));
 sg13g2_nand2_1 _16204_ (.Y(_10419_),
    .A(_08126_),
    .B(_09819_));
 sg13g2_o21ai_1 _16205_ (.B1(net995),
    .Y(_10420_),
    .A1(_10416_),
    .A2(_10419_));
 sg13g2_nand2_1 _16206_ (.Y(_10421_),
    .A(_09661_),
    .B(\top_ihp.wb_dati_uart[5] ));
 sg13g2_nor2_1 _16207_ (.A(_00103_),
    .B(net879),
    .Y(_10422_));
 sg13g2_inv_1 _16208_ (.Y(_10423_),
    .A(_00105_));
 sg13g2_a22oi_1 _16209_ (.Y(_10424_),
    .B1(net919),
    .B2(\top_ihp.wb_coproc.dat_o[5] ),
    .A2(_10423_),
    .A1(net994));
 sg13g2_and4_1 _16210_ (.A(net1024),
    .B(_00104_),
    .C(net914),
    .D(_09870_),
    .X(_10425_));
 sg13g2_a221oi_1 _16211_ (.B2(_10424_),
    .C1(_10425_),
    .B1(net854),
    .A1(net992),
    .Y(_10426_),
    .A2(net905));
 sg13g2_o21ai_1 _16212_ (.B1(net987),
    .Y(_10427_),
    .A1(_10422_),
    .A2(_10426_));
 sg13g2_nand2_1 _16213_ (.Y(_10428_),
    .A(_10421_),
    .B(_10427_));
 sg13g2_buf_2 _16214_ (.A(_10428_),
    .X(_10429_));
 sg13g2_buf_8 _16215_ (.A(_10429_),
    .X(_10430_));
 sg13g2_a22oi_1 _16216_ (.Y(_10431_),
    .B1(_10429_),
    .B2(net991),
    .A2(_10161_),
    .A1(net918));
 sg13g2_inv_1 _16217_ (.Y(_10432_),
    .A(_10431_));
 sg13g2_a21oi_1 _16218_ (.A1(net1030),
    .A2(_09923_),
    .Y(_10433_),
    .B1(_09926_));
 sg13g2_o21ai_1 _16219_ (.B1(net952),
    .Y(_10434_),
    .A1(_10363_),
    .A2(_10433_));
 sg13g2_a221oi_1 _16220_ (.B2(_09644_),
    .C1(_10434_),
    .B1(_10432_),
    .A1(_09908_),
    .Y(_10435_),
    .A2(_10430_));
 sg13g2_a21oi_1 _16221_ (.A1(_10231_),
    .A2(_09764_),
    .Y(_10436_),
    .B1(net946));
 sg13g2_o21ai_1 _16222_ (.B1(_10436_),
    .Y(_10437_),
    .A1(_10420_),
    .A2(_10435_));
 sg13g2_o21ai_1 _16223_ (.B1(_10437_),
    .Y(_10438_),
    .A1(_08126_),
    .A2(_10418_));
 sg13g2_buf_1 _16224_ (.A(_10438_),
    .X(_10439_));
 sg13g2_buf_2 _16225_ (.A(_10439_),
    .X(_10440_));
 sg13g2_nand2_1 _16226_ (.Y(_10441_),
    .A(\top_ihp.oisc.regs[0][5] ),
    .B(net527));
 sg13g2_o21ai_1 _16227_ (.B1(_10441_),
    .Y(_00479_),
    .A1(net526),
    .A2(net141));
 sg13g2_o21ai_1 _16228_ (.B1(_08129_),
    .Y(_10442_),
    .A1(_08407_),
    .A2(_10415_));
 sg13g2_nor2_1 _16229_ (.A(net1062),
    .B(_10442_),
    .Y(_10443_));
 sg13g2_nand2_1 _16230_ (.Y(_10444_),
    .A(net1062),
    .B(_10442_));
 sg13g2_nand2b_1 _16231_ (.Y(_10445_),
    .B(_10444_),
    .A_N(_10443_));
 sg13g2_buf_1 _16232_ (.A(_10445_),
    .X(_10446_));
 sg13g2_a221oi_1 _16233_ (.B2(_09764_),
    .C1(_10446_),
    .B1(_10243_),
    .A1(net1058),
    .Y(_10447_),
    .A2(_08823_));
 sg13g2_o21ai_1 _16234_ (.B1(_08139_),
    .Y(_10448_),
    .A1(_09865_),
    .A2(_10447_));
 sg13g2_nand2_1 _16235_ (.Y(_10449_),
    .A(net1028),
    .B(\top_ihp.wb_dati_uart[6] ));
 sg13g2_nor2_1 _16236_ (.A(_00106_),
    .B(_09607_),
    .Y(_10450_));
 sg13g2_inv_1 _16237_ (.Y(_10451_),
    .A(_00108_));
 sg13g2_a22oi_1 _16238_ (.Y(_10452_),
    .B1(net919),
    .B2(\top_ihp.wb_coproc.dat_o[6] ),
    .A2(_10451_),
    .A1(net994));
 sg13g2_and4_1 _16239_ (.A(_09784_),
    .B(_00107_),
    .C(_09869_),
    .D(_09870_),
    .X(_10453_));
 sg13g2_a221oi_1 _16240_ (.B2(_10452_),
    .C1(_10453_),
    .B1(net878),
    .A1(net992),
    .Y(_10454_),
    .A2(net905));
 sg13g2_o21ai_1 _16241_ (.B1(net987),
    .Y(_10455_),
    .A1(_10450_),
    .A2(_10454_));
 sg13g2_nand2_1 _16242_ (.Y(_10456_),
    .A(_10449_),
    .B(_10455_));
 sg13g2_buf_2 _16243_ (.A(_10456_),
    .X(_10457_));
 sg13g2_a22oi_1 _16244_ (.Y(_10458_),
    .B1(_10457_),
    .B2(net991),
    .A2(_10179_),
    .A1(net918));
 sg13g2_nor2_1 _16245_ (.A(_09659_),
    .B(_10458_),
    .Y(_10459_));
 sg13g2_a21oi_1 _16246_ (.A1(net1030),
    .A2(_09956_),
    .Y(_10460_),
    .B1(_09959_));
 sg13g2_a21oi_1 _16247_ (.A1(net990),
    .A2(_10457_),
    .Y(_10461_),
    .B1(net988));
 sg13g2_o21ai_1 _16248_ (.B1(_10461_),
    .Y(_10462_),
    .A1(_10363_),
    .A2(_10460_));
 sg13g2_nand3_1 _16249_ (.B(_09819_),
    .C(_10446_),
    .A(net1045),
    .Y(_10463_));
 sg13g2_o21ai_1 _16250_ (.B1(_10463_),
    .Y(_10464_),
    .A1(_10459_),
    .A2(_10462_));
 sg13g2_a21oi_1 _16251_ (.A1(_10243_),
    .A2(_09764_),
    .Y(_10465_),
    .B1(_09863_));
 sg13g2_o21ai_1 _16252_ (.B1(_10465_),
    .Y(_10466_),
    .A1(_09849_),
    .A2(_10464_));
 sg13g2_nand2_1 _16253_ (.Y(_10467_),
    .A(_10448_),
    .B(_10466_));
 sg13g2_buf_2 _16254_ (.A(_10467_),
    .X(_10468_));
 sg13g2_buf_1 _16255_ (.A(_10468_),
    .X(_10469_));
 sg13g2_nand2_1 _16256_ (.Y(_10470_),
    .A(\top_ihp.oisc.regs[0][6] ),
    .B(net661));
 sg13g2_o21ai_1 _16257_ (.B1(_10470_),
    .Y(_00480_),
    .A1(net526),
    .A2(net140));
 sg13g2_nor3_1 _16258_ (.A(_09659_),
    .B(_09779_),
    .C(_09791_),
    .Y(_10471_));
 sg13g2_a21oi_1 _16259_ (.A1(_09659_),
    .A2(_09770_),
    .Y(_10472_),
    .B1(_10471_));
 sg13g2_nand2_1 _16260_ (.Y(_10473_),
    .A(_09780_),
    .B(_09789_));
 sg13g2_nand2_1 _16261_ (.Y(_10474_),
    .A(net1042),
    .B(_10473_));
 sg13g2_o21ai_1 _16262_ (.B1(_10474_),
    .Y(_10475_),
    .A1(net990),
    .A2(_10472_));
 sg13g2_o21ai_1 _16263_ (.B1(_10444_),
    .Y(_10476_),
    .A1(net1045),
    .A2(_10443_));
 sg13g2_xnor2_1 _16264_ (.Y(_10477_),
    .A(_08120_),
    .B(_10476_));
 sg13g2_mux2_1 _16265_ (.A0(_10475_),
    .A1(_10477_),
    .S(net988),
    .X(_10478_));
 sg13g2_a221oi_1 _16266_ (.B2(_09595_),
    .C1(net946),
    .B1(_10478_),
    .A1(\top_ihp.oisc.decoder.instruction[27] ),
    .Y(_10479_),
    .A2(_09764_));
 sg13g2_buf_2 _16267_ (.A(_10479_),
    .X(_10480_));
 sg13g2_nor2_1 _16268_ (.A(_08116_),
    .B(net953),
    .Y(_10481_));
 sg13g2_or2_1 _16269_ (.X(_10482_),
    .B(_10481_),
    .A(_10480_));
 sg13g2_buf_2 _16270_ (.A(_10482_),
    .X(_10483_));
 sg13g2_buf_1 _16271_ (.A(_10483_),
    .X(_10484_));
 sg13g2_nand2_1 _16272_ (.Y(_10485_),
    .A(\top_ihp.oisc.regs[0][7] ),
    .B(net661));
 sg13g2_o21ai_1 _16273_ (.B1(_10485_),
    .Y(_00481_),
    .A1(_10262_),
    .A2(net139));
 sg13g2_and2_1 _16274_ (.A(\top_ihp.oisc.decoder.instruction[28] ),
    .B(net996),
    .X(_10486_));
 sg13g2_inv_1 _16275_ (.Y(_10487_),
    .A(_08116_));
 sg13g2_a221oi_1 _16276_ (.B2(net1062),
    .C1(_10442_),
    .B1(_08139_),
    .A1(_10487_),
    .Y(_10488_),
    .A2(_08115_));
 sg13g2_nor2_1 _16277_ (.A(_08125_),
    .B(_08119_),
    .Y(_10489_));
 sg13g2_nor3_1 _16278_ (.A(_08117_),
    .B(_10488_),
    .C(_10489_),
    .Y(_10490_));
 sg13g2_xor2_1 _16279_ (.B(_10490_),
    .A(_08101_),
    .X(_10491_));
 sg13g2_xnor2_1 _16280_ (.Y(_10492_),
    .A(_08133_),
    .B(_10491_));
 sg13g2_inv_1 _16281_ (.Y(_10493_),
    .A(_09636_));
 sg13g2_a21o_1 _16282_ (.A2(net918),
    .A1(_09628_),
    .B1(_09637_),
    .X(_10494_));
 sg13g2_a22oi_1 _16283_ (.Y(_10495_),
    .B1(_10494_),
    .B2(_09815_),
    .A2(_10493_),
    .A1(_09908_));
 sg13g2_a221oi_1 _16284_ (.B2(_09797_),
    .C1(_09748_),
    .B1(_10495_),
    .A1(net947),
    .Y(_10496_),
    .A2(_10492_));
 sg13g2_a221oi_1 _16285_ (.B2(_10486_),
    .C1(_10496_),
    .B1(_09764_),
    .A1(_08100_),
    .Y(_10497_),
    .A2(net915));
 sg13g2_buf_2 _16286_ (.A(_10497_),
    .X(_10498_));
 sg13g2_buf_8 _16287_ (.A(_10498_),
    .X(_10499_));
 sg13g2_nand2_1 _16288_ (.Y(_10500_),
    .A(\top_ihp.oisc.regs[0][8] ),
    .B(_09756_));
 sg13g2_o21ai_1 _16289_ (.B1(_10500_),
    .Y(_00482_),
    .A1(_09758_),
    .A2(net316));
 sg13g2_nor2_1 _16290_ (.A(_10106_),
    .B(_10109_),
    .Y(_10501_));
 sg13g2_nor2_1 _16291_ (.A(net944),
    .B(_10501_),
    .Y(_10502_));
 sg13g2_nand2_1 _16292_ (.Y(_10503_),
    .A(net918),
    .B(_10227_));
 sg13g2_o21ai_1 _16293_ (.B1(_10503_),
    .Y(_10504_),
    .A1(net1030),
    .A2(_10110_));
 sg13g2_a22oi_1 _16294_ (.Y(_10505_),
    .B1(_10504_),
    .B2(net1023),
    .A2(_10502_),
    .A1(net986));
 sg13g2_inv_1 _16295_ (.Y(_10506_),
    .A(\top_ihp.oisc.op_b[9] ));
 sg13g2_xnor2_1 _16296_ (.Y(_10507_),
    .A(_10506_),
    .B(_08413_));
 sg13g2_xor2_1 _16297_ (.B(_10507_),
    .A(_08103_),
    .X(_10508_));
 sg13g2_a221oi_1 _16298_ (.B2(_09848_),
    .C1(net1022),
    .B1(_10508_),
    .A1(_09797_),
    .Y(_10509_),
    .A2(_10505_));
 sg13g2_a21oi_1 _16299_ (.A1(\top_ihp.oisc.decoder.instruction[29] ),
    .A2(_09764_),
    .Y(_10510_),
    .B1(net946));
 sg13g2_nand2b_1 _16300_ (.Y(_10511_),
    .B(_10510_),
    .A_N(_10509_));
 sg13g2_o21ai_1 _16301_ (.B1(_10511_),
    .Y(_10512_),
    .A1(_08103_),
    .A2(net953));
 sg13g2_buf_2 _16302_ (.A(_10512_),
    .X(_10513_));
 sg13g2_buf_1 _16303_ (.A(_10513_),
    .X(_10514_));
 sg13g2_nand2_1 _16304_ (.Y(_10515_),
    .A(\top_ihp.oisc.regs[0][9] ),
    .B(net661));
 sg13g2_o21ai_1 _16305_ (.B1(_10515_),
    .Y(_00483_),
    .A1(_09758_),
    .A2(_10514_));
 sg13g2_nor2_1 _16306_ (.A(_09494_),
    .B(_09720_),
    .Y(_10516_));
 sg13g2_a22oi_1 _16307_ (.Y(_10517_),
    .B1(_09714_),
    .B2(_10516_),
    .A2(_09702_),
    .A1(_09494_));
 sg13g2_nor2b_1 _16308_ (.A(_10517_),
    .B_N(_09723_),
    .Y(_10518_));
 sg13g2_buf_2 _16309_ (.A(_10518_),
    .X(_10519_));
 sg13g2_buf_8 _16310_ (.A(_10519_),
    .X(_10520_));
 sg13g2_and2_1 _16311_ (.A(_09750_),
    .B(_09744_),
    .X(_10521_));
 sg13g2_buf_1 _16312_ (.A(_10521_),
    .X(_10522_));
 sg13g2_nor2b_1 _16313_ (.A(_09739_),
    .B_N(_10522_),
    .Y(_10523_));
 sg13g2_buf_1 _16314_ (.A(_10523_),
    .X(_10524_));
 sg13g2_nand2_1 _16315_ (.Y(_10525_),
    .A(net764),
    .B(_10524_));
 sg13g2_buf_1 _16316_ (.A(_10525_),
    .X(_10526_));
 sg13g2_buf_1 _16317_ (.A(net659),
    .X(_10527_));
 sg13g2_mux2_1 _16318_ (.A0(net156),
    .A1(_00235_),
    .S(net524),
    .X(_00484_));
 sg13g2_buf_1 _16319_ (.A(net659),
    .X(_10528_));
 sg13g2_nand2_1 _16320_ (.Y(_10529_),
    .A(\top_ihp.oisc.regs[10][10] ),
    .B(net524));
 sg13g2_o21ai_1 _16321_ (.B1(_10529_),
    .Y(_00485_),
    .A1(net155),
    .A2(net523));
 sg13g2_nand2_1 _16322_ (.Y(_10530_),
    .A(\top_ihp.oisc.regs[10][11] ),
    .B(net524));
 sg13g2_o21ai_1 _16323_ (.B1(_10530_),
    .Y(_00486_),
    .A1(net154),
    .A2(net523));
 sg13g2_buf_8 _16324_ (.A(_09905_),
    .X(_10531_));
 sg13g2_nand2_1 _16325_ (.Y(_10532_),
    .A(\top_ihp.oisc.regs[10][12] ),
    .B(net524));
 sg13g2_o21ai_1 _16326_ (.B1(_10532_),
    .Y(_00487_),
    .A1(net137),
    .A2(_10528_));
 sg13g2_nand2_1 _16327_ (.Y(_10533_),
    .A(\top_ihp.oisc.regs[10][13] ),
    .B(net524));
 sg13g2_o21ai_1 _16328_ (.B1(_10533_),
    .Y(_00488_),
    .A1(net331),
    .A2(net523));
 sg13g2_buf_8 _16329_ (.A(_09977_),
    .X(_10534_));
 sg13g2_nand2_1 _16330_ (.Y(_10535_),
    .A(\top_ihp.oisc.regs[10][14] ),
    .B(net524));
 sg13g2_o21ai_1 _16331_ (.B1(_10535_),
    .Y(_00489_),
    .A1(net136),
    .A2(net523));
 sg13g2_buf_8 _16332_ (.A(_09992_),
    .X(_10536_));
 sg13g2_nand2_1 _16333_ (.Y(_10537_),
    .A(\top_ihp.oisc.regs[10][15] ),
    .B(net524));
 sg13g2_o21ai_1 _16334_ (.B1(_10537_),
    .Y(_00490_),
    .A1(net135),
    .A2(net523));
 sg13g2_nand2_1 _16335_ (.Y(_10538_),
    .A(\top_ihp.oisc.regs[10][16] ),
    .B(net524));
 sg13g2_o21ai_1 _16336_ (.B1(_10538_),
    .Y(_00491_),
    .A1(net150),
    .A2(net523));
 sg13g2_nand2_1 _16337_ (.Y(_10539_),
    .A(\top_ihp.oisc.regs[10][17] ),
    .B(_10527_));
 sg13g2_o21ai_1 _16338_ (.B1(_10539_),
    .Y(_00492_),
    .A1(net328),
    .A2(_10528_));
 sg13g2_buf_1 _16339_ (.A(net659),
    .X(_10540_));
 sg13g2_nand2_1 _16340_ (.Y(_10541_),
    .A(\top_ihp.oisc.regs[10][18] ),
    .B(net522));
 sg13g2_o21ai_1 _16341_ (.B1(_10541_),
    .Y(_00493_),
    .A1(net327),
    .A2(net523));
 sg13g2_nand2_1 _16342_ (.Y(_10542_),
    .A(\top_ihp.oisc.regs[10][19] ),
    .B(net522));
 sg13g2_o21ai_1 _16343_ (.B1(_10542_),
    .Y(_00494_),
    .A1(net326),
    .A2(net523));
 sg13g2_buf_1 _16344_ (.A(net325),
    .X(_10543_));
 sg13g2_buf_1 _16345_ (.A(_10526_),
    .X(_10544_));
 sg13g2_nand2_1 _16346_ (.Y(_10545_),
    .A(\top_ihp.oisc.regs[10][1] ),
    .B(_10540_));
 sg13g2_o21ai_1 _16347_ (.B1(_10545_),
    .Y(_00495_),
    .A1(net134),
    .A2(net521));
 sg13g2_nand2_1 _16348_ (.Y(_10546_),
    .A(\top_ihp.oisc.regs[10][20] ),
    .B(net522));
 sg13g2_o21ai_1 _16349_ (.B1(_10546_),
    .Y(_00496_),
    .A1(net324),
    .A2(net521));
 sg13g2_nand2_1 _16350_ (.Y(_10547_),
    .A(\top_ihp.oisc.regs[10][21] ),
    .B(net522));
 sg13g2_o21ai_1 _16351_ (.B1(_10547_),
    .Y(_00497_),
    .A1(net323),
    .A2(net521));
 sg13g2_buf_8 _16352_ (.A(_10188_),
    .X(_10548_));
 sg13g2_nand2_1 _16353_ (.Y(_10549_),
    .A(\top_ihp.oisc.regs[10][22] ),
    .B(_10540_));
 sg13g2_o21ai_1 _16354_ (.B1(_10549_),
    .Y(_00498_),
    .A1(net133),
    .A2(net521));
 sg13g2_nand2_1 _16355_ (.Y(_10550_),
    .A(\top_ihp.oisc.regs[10][23] ),
    .B(net522));
 sg13g2_o21ai_1 _16356_ (.B1(_10550_),
    .Y(_00499_),
    .A1(net321),
    .A2(net521));
 sg13g2_nand2_1 _16357_ (.Y(_10551_),
    .A(\top_ihp.oisc.regs[10][24] ),
    .B(net522));
 sg13g2_o21ai_1 _16358_ (.B1(_10551_),
    .Y(_00500_),
    .A1(net320),
    .A2(_10544_));
 sg13g2_nand2_1 _16359_ (.Y(_10552_),
    .A(\top_ihp.oisc.regs[10][25] ),
    .B(net522));
 sg13g2_o21ai_1 _16360_ (.B1(_10552_),
    .Y(_00501_),
    .A1(net147),
    .A2(net521));
 sg13g2_nand2_1 _16361_ (.Y(_10553_),
    .A(\top_ihp.oisc.regs[10][26] ),
    .B(net522));
 sg13g2_o21ai_1 _16362_ (.B1(_10553_),
    .Y(_00502_),
    .A1(net146),
    .A2(net521));
 sg13g2_buf_8 _16363_ (.A(net659),
    .X(_10554_));
 sg13g2_nand2_1 _16364_ (.Y(_10555_),
    .A(\top_ihp.oisc.regs[10][27] ),
    .B(net520));
 sg13g2_o21ai_1 _16365_ (.B1(_10555_),
    .Y(_00503_),
    .A1(net318),
    .A2(net521));
 sg13g2_nand2_1 _16366_ (.Y(_10556_),
    .A(\top_ihp.oisc.regs[10][28] ),
    .B(_10554_));
 sg13g2_o21ai_1 _16367_ (.B1(_10556_),
    .Y(_00504_),
    .A1(net525),
    .A2(_10544_));
 sg13g2_buf_8 _16368_ (.A(net659),
    .X(_10557_));
 sg13g2_nand2_1 _16369_ (.Y(_10558_),
    .A(\top_ihp.oisc.regs[10][29] ),
    .B(net520));
 sg13g2_o21ai_1 _16370_ (.B1(_10558_),
    .Y(_00505_),
    .A1(net317),
    .A2(net519));
 sg13g2_nand2_1 _16371_ (.Y(_10559_),
    .A(\top_ihp.oisc.regs[10][2] ),
    .B(net520));
 sg13g2_o21ai_1 _16372_ (.B1(_10559_),
    .Y(_00506_),
    .A1(net145),
    .A2(net519));
 sg13g2_nand2_1 _16373_ (.Y(_10560_),
    .A(\top_ihp.oisc.regs[10][30] ),
    .B(net520));
 sg13g2_o21ai_1 _16374_ (.B1(_10560_),
    .Y(_00507_),
    .A1(net144),
    .A2(net519));
 sg13g2_nand2_1 _16375_ (.Y(_10561_),
    .A(\top_ihp.oisc.regs[10][31] ),
    .B(net520));
 sg13g2_o21ai_1 _16376_ (.B1(_10561_),
    .Y(_00508_),
    .A1(net52),
    .A2(net519));
 sg13g2_nand2_1 _16377_ (.Y(_10562_),
    .A(\top_ihp.oisc.regs[10][3] ),
    .B(net520));
 sg13g2_o21ai_1 _16378_ (.B1(_10562_),
    .Y(_00509_),
    .A1(net143),
    .A2(net519));
 sg13g2_nand2_1 _16379_ (.Y(_10563_),
    .A(\top_ihp.oisc.regs[10][4] ),
    .B(net520));
 sg13g2_o21ai_1 _16380_ (.B1(_10563_),
    .Y(_00510_),
    .A1(net142),
    .A2(net519));
 sg13g2_nand2_1 _16381_ (.Y(_10564_),
    .A(\top_ihp.oisc.regs[10][5] ),
    .B(net520));
 sg13g2_o21ai_1 _16382_ (.B1(_10564_),
    .Y(_00511_),
    .A1(net141),
    .A2(net519));
 sg13g2_nand2_1 _16383_ (.Y(_10565_),
    .A(\top_ihp.oisc.regs[10][6] ),
    .B(_10554_));
 sg13g2_o21ai_1 _16384_ (.B1(_10565_),
    .Y(_00512_),
    .A1(net140),
    .A2(_10557_));
 sg13g2_nand2_1 _16385_ (.Y(_10566_),
    .A(\top_ihp.oisc.regs[10][7] ),
    .B(net659));
 sg13g2_o21ai_1 _16386_ (.B1(_10566_),
    .Y(_00513_),
    .A1(net139),
    .A2(_10557_));
 sg13g2_nand2_1 _16387_ (.Y(_10567_),
    .A(\top_ihp.oisc.regs[10][8] ),
    .B(net659));
 sg13g2_o21ai_1 _16388_ (.B1(_10567_),
    .Y(_00514_),
    .A1(net316),
    .A2(net519));
 sg13g2_nand2_1 _16389_ (.Y(_10568_),
    .A(\top_ihp.oisc.regs[10][9] ),
    .B(net659));
 sg13g2_o21ai_1 _16390_ (.B1(_10568_),
    .Y(_00515_),
    .A1(net138),
    .A2(_10527_));
 sg13g2_nor2_1 _16391_ (.A(_09750_),
    .B(_09743_),
    .Y(_10569_));
 sg13g2_buf_1 _16392_ (.A(_10569_),
    .X(_10570_));
 sg13g2_nor2b_1 _16393_ (.A(_09739_),
    .B_N(net785),
    .Y(_10571_));
 sg13g2_buf_1 _16394_ (.A(_10571_),
    .X(_10572_));
 sg13g2_nand2_1 _16395_ (.Y(_10573_),
    .A(net764),
    .B(_10572_));
 sg13g2_buf_2 _16396_ (.A(_10573_),
    .X(_10574_));
 sg13g2_buf_1 _16397_ (.A(_10574_),
    .X(_10575_));
 sg13g2_mux2_1 _16398_ (.A0(net156),
    .A1(_00236_),
    .S(_10575_),
    .X(_00516_));
 sg13g2_buf_1 _16399_ (.A(_10574_),
    .X(_10576_));
 sg13g2_buf_1 _16400_ (.A(_10574_),
    .X(_10577_));
 sg13g2_nand2_1 _16401_ (.Y(_10578_),
    .A(\top_ihp.oisc.regs[11][10] ),
    .B(net656));
 sg13g2_o21ai_1 _16402_ (.B1(_10578_),
    .Y(_00517_),
    .A1(net155),
    .A2(net657));
 sg13g2_nand2_1 _16403_ (.Y(_10579_),
    .A(\top_ihp.oisc.regs[11][11] ),
    .B(net656));
 sg13g2_o21ai_1 _16404_ (.B1(_10579_),
    .Y(_00518_),
    .A1(net154),
    .A2(net657));
 sg13g2_nand2_1 _16405_ (.Y(_10580_),
    .A(\top_ihp.oisc.regs[11][12] ),
    .B(net656));
 sg13g2_o21ai_1 _16406_ (.B1(_10580_),
    .Y(_00519_),
    .A1(net137),
    .A2(_10576_));
 sg13g2_nand2_1 _16407_ (.Y(_10581_),
    .A(\top_ihp.oisc.regs[11][13] ),
    .B(net656));
 sg13g2_o21ai_1 _16408_ (.B1(_10581_),
    .Y(_00520_),
    .A1(net331),
    .A2(net657));
 sg13g2_nand2_1 _16409_ (.Y(_10582_),
    .A(\top_ihp.oisc.regs[11][14] ),
    .B(net656));
 sg13g2_o21ai_1 _16410_ (.B1(_10582_),
    .Y(_00521_),
    .A1(net136),
    .A2(net657));
 sg13g2_nand2_1 _16411_ (.Y(_10583_),
    .A(\top_ihp.oisc.regs[11][15] ),
    .B(_10577_));
 sg13g2_o21ai_1 _16412_ (.B1(_10583_),
    .Y(_00522_),
    .A1(net135),
    .A2(net657));
 sg13g2_nand2_1 _16413_ (.Y(_10584_),
    .A(\top_ihp.oisc.regs[11][16] ),
    .B(_10577_));
 sg13g2_o21ai_1 _16414_ (.B1(_10584_),
    .Y(_00523_),
    .A1(net150),
    .A2(net657));
 sg13g2_nand2_1 _16415_ (.Y(_10585_),
    .A(\top_ihp.oisc.regs[11][17] ),
    .B(net656));
 sg13g2_o21ai_1 _16416_ (.B1(_10585_),
    .Y(_00524_),
    .A1(net328),
    .A2(net657));
 sg13g2_buf_1 _16417_ (.A(_10574_),
    .X(_10586_));
 sg13g2_nand2_1 _16418_ (.Y(_10587_),
    .A(\top_ihp.oisc.regs[11][18] ),
    .B(net655));
 sg13g2_o21ai_1 _16419_ (.B1(_10587_),
    .Y(_00525_),
    .A1(net327),
    .A2(_10576_));
 sg13g2_nand2_1 _16420_ (.Y(_10588_),
    .A(\top_ihp.oisc.regs[11][19] ),
    .B(net655));
 sg13g2_o21ai_1 _16421_ (.B1(_10588_),
    .Y(_00526_),
    .A1(net326),
    .A2(net657));
 sg13g2_buf_1 _16422_ (.A(_10574_),
    .X(_10589_));
 sg13g2_nand2_1 _16423_ (.Y(_10590_),
    .A(_00237_),
    .B(_10586_));
 sg13g2_o21ai_1 _16424_ (.B1(_10590_),
    .Y(_00527_),
    .A1(_10125_),
    .A2(net654));
 sg13g2_buf_2 _16425_ (.A(_10144_),
    .X(_10591_));
 sg13g2_nand2_1 _16426_ (.Y(_10592_),
    .A(\top_ihp.oisc.regs[11][20] ),
    .B(_10586_));
 sg13g2_o21ai_1 _16427_ (.B1(_10592_),
    .Y(_00528_),
    .A1(net653),
    .A2(net654));
 sg13g2_nand2_1 _16428_ (.Y(_10593_),
    .A(\top_ihp.oisc.regs[11][21] ),
    .B(net655));
 sg13g2_o21ai_1 _16429_ (.B1(_10593_),
    .Y(_00529_),
    .A1(net323),
    .A2(net654));
 sg13g2_nand2_1 _16430_ (.Y(_10594_),
    .A(\top_ihp.oisc.regs[11][22] ),
    .B(net655));
 sg13g2_o21ai_1 _16431_ (.B1(_10594_),
    .Y(_00530_),
    .A1(net133),
    .A2(net654));
 sg13g2_nand2_1 _16432_ (.Y(_10595_),
    .A(\top_ihp.oisc.regs[11][23] ),
    .B(net655));
 sg13g2_o21ai_1 _16433_ (.B1(_10595_),
    .Y(_00531_),
    .A1(net321),
    .A2(net654));
 sg13g2_nand2_1 _16434_ (.Y(_10596_),
    .A(\top_ihp.oisc.regs[11][24] ),
    .B(net655));
 sg13g2_o21ai_1 _16435_ (.B1(_10596_),
    .Y(_00532_),
    .A1(net320),
    .A2(_10589_));
 sg13g2_buf_8 _16436_ (.A(_10236_),
    .X(_10597_));
 sg13g2_nand2_1 _16437_ (.Y(_10598_),
    .A(\top_ihp.oisc.regs[11][25] ),
    .B(net655));
 sg13g2_o21ai_1 _16438_ (.B1(_10598_),
    .Y(_00533_),
    .A1(net132),
    .A2(net654));
 sg13g2_nand2_1 _16439_ (.Y(_10599_),
    .A(\top_ihp.oisc.regs[11][26] ),
    .B(net655));
 sg13g2_o21ai_1 _16440_ (.B1(_10599_),
    .Y(_00534_),
    .A1(net146),
    .A2(_10589_));
 sg13g2_buf_1 _16441_ (.A(_10574_),
    .X(_10600_));
 sg13g2_nand2_1 _16442_ (.Y(_10601_),
    .A(\top_ihp.oisc.regs[11][27] ),
    .B(net652));
 sg13g2_o21ai_1 _16443_ (.B1(_10601_),
    .Y(_00535_),
    .A1(net318),
    .A2(net654));
 sg13g2_nand2_1 _16444_ (.Y(_10602_),
    .A(\top_ihp.oisc.regs[11][28] ),
    .B(net652));
 sg13g2_o21ai_1 _16445_ (.B1(_10602_),
    .Y(_00536_),
    .A1(net525),
    .A2(net654));
 sg13g2_nand2_1 _16446_ (.Y(_10603_),
    .A(\top_ihp.oisc.regs[11][29] ),
    .B(net652));
 sg13g2_o21ai_1 _16447_ (.B1(_10603_),
    .Y(_00537_),
    .A1(net317),
    .A2(net658));
 sg13g2_buf_8 _16448_ (.A(_10314_),
    .X(_10604_));
 sg13g2_mux2_1 _16449_ (.A0(net131),
    .A1(_00238_),
    .S(net658),
    .X(_00538_));
 sg13g2_nand2_1 _16450_ (.Y(_10605_),
    .A(\top_ihp.oisc.regs[11][30] ),
    .B(net652));
 sg13g2_o21ai_1 _16451_ (.B1(_10605_),
    .Y(_00539_),
    .A1(net144),
    .A2(net658));
 sg13g2_buf_8 _16452_ (.A(_10345_),
    .X(_10606_));
 sg13g2_nand2_1 _16453_ (.Y(_10607_),
    .A(\top_ihp.oisc.regs[11][31] ),
    .B(net652));
 sg13g2_o21ai_1 _16454_ (.B1(_10607_),
    .Y(_00540_),
    .A1(net315),
    .A2(net658));
 sg13g2_buf_1 _16455_ (.A(_10380_),
    .X(_10608_));
 sg13g2_mux2_1 _16456_ (.A0(net130),
    .A1(_00239_),
    .S(net656),
    .X(_00541_));
 sg13g2_buf_1 _16457_ (.A(_10412_),
    .X(_10609_));
 sg13g2_mux2_1 _16458_ (.A0(net129),
    .A1(_00240_),
    .S(net656),
    .X(_00542_));
 sg13g2_nand2_1 _16459_ (.Y(_10610_),
    .A(\top_ihp.oisc.regs[11][5] ),
    .B(net652));
 sg13g2_o21ai_1 _16460_ (.B1(_10610_),
    .Y(_00543_),
    .A1(net141),
    .A2(net658));
 sg13g2_nand2_1 _16461_ (.Y(_10611_),
    .A(\top_ihp.oisc.regs[11][6] ),
    .B(net652));
 sg13g2_o21ai_1 _16462_ (.B1(_10611_),
    .Y(_00544_),
    .A1(net140),
    .A2(net658));
 sg13g2_buf_2 _16463_ (.A(_10480_),
    .X(_10612_));
 sg13g2_nand2_1 _16464_ (.Y(_10613_),
    .A(\top_ihp.oisc.regs[11][7] ),
    .B(_10600_));
 sg13g2_o21ai_1 _16465_ (.B1(_10613_),
    .Y(_00545_),
    .A1(net518),
    .A2(net658));
 sg13g2_nand2_1 _16466_ (.Y(_10614_),
    .A(\top_ihp.oisc.regs[11][8] ),
    .B(net652));
 sg13g2_o21ai_1 _16467_ (.B1(_10614_),
    .Y(_00546_),
    .A1(net316),
    .A2(net658));
 sg13g2_nand2_1 _16468_ (.Y(_10615_),
    .A(\top_ihp.oisc.regs[11][9] ),
    .B(_10600_));
 sg13g2_o21ai_1 _16469_ (.B1(_10615_),
    .Y(_00547_),
    .A1(net138),
    .A2(_10575_));
 sg13g2_inv_1 _16470_ (.Y(_10616_),
    .A(_09714_));
 sg13g2_nor3_2 _16471_ (.A(_10616_),
    .B(_10516_),
    .C(_09727_),
    .Y(_10617_));
 sg13g2_buf_2 _16472_ (.A(_10617_),
    .X(_10618_));
 sg13g2_buf_1 _16473_ (.A(_10618_),
    .X(_10619_));
 sg13g2_nand2_1 _16474_ (.Y(_10620_),
    .A(_09754_),
    .B(net763));
 sg13g2_buf_1 _16475_ (.A(_10620_),
    .X(_10621_));
 sg13g2_buf_2 _16476_ (.A(net651),
    .X(_10622_));
 sg13g2_mux2_1 _16477_ (.A0(net156),
    .A1(_00241_),
    .S(net517),
    .X(_00548_));
 sg13g2_buf_8 _16478_ (.A(_09824_),
    .X(_10623_));
 sg13g2_mux2_1 _16479_ (.A0(net128),
    .A1(_00242_),
    .S(net517),
    .X(_00549_));
 sg13g2_buf_8 _16480_ (.A(_09860_),
    .X(_10624_));
 sg13g2_mux2_1 _16481_ (.A0(net127),
    .A1(_00243_),
    .S(net517),
    .X(_00550_));
 sg13g2_nand2_1 _16482_ (.Y(_10625_),
    .A(_00244_),
    .B(net651));
 sg13g2_o21ai_1 _16483_ (.B1(_10625_),
    .Y(_00551_),
    .A1(_09903_),
    .A2(net517));
 sg13g2_buf_8 _16484_ (.A(_09941_),
    .X(_10626_));
 sg13g2_mux2_1 _16485_ (.A0(net314),
    .A1(_00245_),
    .S(net517),
    .X(_00552_));
 sg13g2_mux2_1 _16486_ (.A0(net330),
    .A1(_00246_),
    .S(_10622_),
    .X(_00553_));
 sg13g2_buf_1 _16487_ (.A(net651),
    .X(_10627_));
 sg13g2_mux2_1 _16488_ (.A0(net329),
    .A1(_00247_),
    .S(_10627_),
    .X(_00554_));
 sg13g2_buf_8 _16489_ (.A(_10014_),
    .X(_10628_));
 sg13g2_mux2_1 _16490_ (.A0(net126),
    .A1(_00248_),
    .S(_10627_),
    .X(_00555_));
 sg13g2_buf_1 _16491_ (.A(_10038_),
    .X(_10629_));
 sg13g2_mux2_1 _16492_ (.A0(net313),
    .A1(_00249_),
    .S(net516),
    .X(_00556_));
 sg13g2_buf_1 _16493_ (.A(_10059_),
    .X(_10630_));
 sg13g2_mux2_1 _16494_ (.A0(net312),
    .A1(_00250_),
    .S(net516),
    .X(_00557_));
 sg13g2_buf_8 _16495_ (.A(_10084_),
    .X(_10631_));
 sg13g2_mux2_1 _16496_ (.A0(net311),
    .A1(_00251_),
    .S(net516),
    .X(_00558_));
 sg13g2_nand2_1 _16497_ (.Y(_10632_),
    .A(_00252_),
    .B(net651));
 sg13g2_o21ai_1 _16498_ (.B1(_10632_),
    .Y(_00559_),
    .A1(_10125_),
    .A2(net517));
 sg13g2_mux2_1 _16499_ (.A0(_10144_),
    .A1(_00253_),
    .S(net516),
    .X(_00560_));
 sg13g2_buf_8 _16500_ (.A(_10168_),
    .X(_10633_));
 sg13g2_mux2_1 _16501_ (.A0(net310),
    .A1(_00254_),
    .S(net516),
    .X(_00561_));
 sg13g2_nand2_1 _16502_ (.Y(_10634_),
    .A(_00255_),
    .B(_10621_));
 sg13g2_o21ai_1 _16503_ (.B1(_10634_),
    .Y(_00562_),
    .A1(_10186_),
    .A2(_10622_));
 sg13g2_nand2_1 _16504_ (.Y(_10635_),
    .A(_00256_),
    .B(net651));
 sg13g2_o21ai_1 _16505_ (.B1(_10635_),
    .Y(_00563_),
    .A1(_10195_),
    .A2(net517));
 sg13g2_buf_8 _16506_ (.A(_10216_),
    .X(_10636_));
 sg13g2_mux2_1 _16507_ (.A0(net309),
    .A1(_00257_),
    .S(net516),
    .X(_00564_));
 sg13g2_nand2_1 _16508_ (.Y(_10637_),
    .A(_00258_),
    .B(net651));
 sg13g2_o21ai_1 _16509_ (.B1(_10637_),
    .Y(_00565_),
    .A1(_10234_),
    .A2(net517));
 sg13g2_buf_1 _16510_ (.A(_10247_),
    .X(_10638_));
 sg13g2_mux2_1 _16511_ (.A0(net125),
    .A1(_00259_),
    .S(net516),
    .X(_00566_));
 sg13g2_buf_1 _16512_ (.A(_10259_),
    .X(_10639_));
 sg13g2_mux2_1 _16513_ (.A0(net308),
    .A1(_00260_),
    .S(net516),
    .X(_00567_));
 sg13g2_buf_8 _16514_ (.A(_10268_),
    .X(_10640_));
 sg13g2_buf_2 _16515_ (.A(net651),
    .X(_10641_));
 sg13g2_mux2_1 _16516_ (.A0(net515),
    .A1(_00261_),
    .S(_10641_),
    .X(_00568_));
 sg13g2_buf_8 _16517_ (.A(_10280_),
    .X(_10642_));
 sg13g2_mux2_1 _16518_ (.A0(net307),
    .A1(_00262_),
    .S(net514),
    .X(_00569_));
 sg13g2_mux2_1 _16519_ (.A0(net131),
    .A1(_00263_),
    .S(_10641_),
    .X(_00570_));
 sg13g2_buf_8 _16520_ (.A(_10326_),
    .X(_10643_));
 sg13g2_mux2_1 _16521_ (.A0(net124),
    .A1(_00264_),
    .S(net514),
    .X(_00571_));
 sg13g2_buf_8 _16522_ (.A(_10345_),
    .X(_10644_));
 sg13g2_mux2_1 _16523_ (.A0(net306),
    .A1(_00265_),
    .S(net514),
    .X(_00572_));
 sg13g2_mux2_1 _16524_ (.A0(net130),
    .A1(_00266_),
    .S(net514),
    .X(_00573_));
 sg13g2_mux2_1 _16525_ (.A0(net129),
    .A1(_00267_),
    .S(net514),
    .X(_00574_));
 sg13g2_buf_1 _16526_ (.A(_10439_),
    .X(_10645_));
 sg13g2_mux2_1 _16527_ (.A0(net123),
    .A1(_00268_),
    .S(net514),
    .X(_00575_));
 sg13g2_buf_2 _16528_ (.A(_10468_),
    .X(_10646_));
 sg13g2_mux2_1 _16529_ (.A0(net122),
    .A1(_00269_),
    .S(net514),
    .X(_00576_));
 sg13g2_mux2_1 _16530_ (.A0(_10480_),
    .A1(_00270_),
    .S(net514),
    .X(_00577_));
 sg13g2_buf_8 _16531_ (.A(_10498_),
    .X(_10647_));
 sg13g2_mux2_1 _16532_ (.A0(net305),
    .A1(_00271_),
    .S(net651),
    .X(_00578_));
 sg13g2_buf_8 _16533_ (.A(_10513_),
    .X(_10648_));
 sg13g2_mux2_1 _16534_ (.A0(net121),
    .A1(_00272_),
    .S(_10621_),
    .X(_00579_));
 sg13g2_nor2b_1 _16535_ (.A(_09750_),
    .B_N(_09743_),
    .Y(_10649_));
 sg13g2_nor2b_1 _16536_ (.A(_09739_),
    .B_N(_10649_),
    .Y(_10650_));
 sg13g2_buf_1 _16537_ (.A(_10650_),
    .X(_10651_));
 sg13g2_nand2_1 _16538_ (.Y(_10652_),
    .A(net763),
    .B(_10651_));
 sg13g2_buf_1 _16539_ (.A(_10652_),
    .X(_10653_));
 sg13g2_buf_1 _16540_ (.A(net736),
    .X(_10654_));
 sg13g2_nand2_1 _16541_ (.Y(_10655_),
    .A(\top_ihp.oisc.regs[13][0] ),
    .B(net736));
 sg13g2_o21ai_1 _16542_ (.B1(_10655_),
    .Y(_00580_),
    .A1(net53),
    .A2(net718));
 sg13g2_mux2_1 _16543_ (.A0(net128),
    .A1(_00273_),
    .S(net718),
    .X(_00581_));
 sg13g2_mux2_1 _16544_ (.A0(net127),
    .A1(_00274_),
    .S(_10654_),
    .X(_00582_));
 sg13g2_nand2_1 _16545_ (.Y(_10656_),
    .A(_00275_),
    .B(net736));
 sg13g2_o21ai_1 _16546_ (.B1(_10656_),
    .Y(_00583_),
    .A1(_09903_),
    .A2(net718));
 sg13g2_mux2_1 _16547_ (.A0(net314),
    .A1(_00276_),
    .S(net718),
    .X(_00584_));
 sg13g2_mux2_1 _16548_ (.A0(net330),
    .A1(_00277_),
    .S(_10654_),
    .X(_00585_));
 sg13g2_buf_2 _16549_ (.A(net736),
    .X(_10657_));
 sg13g2_mux2_1 _16550_ (.A0(net329),
    .A1(_00278_),
    .S(_10657_),
    .X(_00586_));
 sg13g2_mux2_1 _16551_ (.A0(net126),
    .A1(_00279_),
    .S(net717),
    .X(_00587_));
 sg13g2_mux2_1 _16552_ (.A0(net313),
    .A1(_00280_),
    .S(net717),
    .X(_00588_));
 sg13g2_mux2_1 _16553_ (.A0(net312),
    .A1(_00281_),
    .S(net717),
    .X(_00589_));
 sg13g2_mux2_1 _16554_ (.A0(net311),
    .A1(_00282_),
    .S(net717),
    .X(_00590_));
 sg13g2_nand2_1 _16555_ (.Y(_10658_),
    .A(\top_ihp.oisc.regs[13][1] ),
    .B(_10653_));
 sg13g2_o21ai_1 _16556_ (.B1(_10658_),
    .Y(_00591_),
    .A1(net134),
    .A2(net718));
 sg13g2_mux2_1 _16557_ (.A0(_10144_),
    .A1(_00283_),
    .S(net717),
    .X(_00592_));
 sg13g2_mux2_1 _16558_ (.A0(net310),
    .A1(_00284_),
    .S(net717),
    .X(_00593_));
 sg13g2_nand2_1 _16559_ (.Y(_10659_),
    .A(_00285_),
    .B(net736));
 sg13g2_o21ai_1 _16560_ (.B1(_10659_),
    .Y(_00594_),
    .A1(_10186_),
    .A2(net718));
 sg13g2_nand2_1 _16561_ (.Y(_10660_),
    .A(_00286_),
    .B(net736));
 sg13g2_o21ai_1 _16562_ (.B1(_10660_),
    .Y(_00595_),
    .A1(_10195_),
    .A2(net718));
 sg13g2_mux2_1 _16563_ (.A0(net309),
    .A1(_00287_),
    .S(_10657_),
    .X(_00596_));
 sg13g2_nand2_1 _16564_ (.Y(_10661_),
    .A(_00288_),
    .B(net736));
 sg13g2_o21ai_1 _16565_ (.B1(_10661_),
    .Y(_00597_),
    .A1(_10234_),
    .A2(net718));
 sg13g2_mux2_1 _16566_ (.A0(net125),
    .A1(_00289_),
    .S(net717),
    .X(_00598_));
 sg13g2_mux2_1 _16567_ (.A0(net308),
    .A1(_00290_),
    .S(net717),
    .X(_00599_));
 sg13g2_buf_2 _16568_ (.A(_10652_),
    .X(_10662_));
 sg13g2_mux2_1 _16569_ (.A0(net515),
    .A1(_00291_),
    .S(net735),
    .X(_00600_));
 sg13g2_mux2_1 _16570_ (.A0(_10642_),
    .A1(_00292_),
    .S(_10662_),
    .X(_00601_));
 sg13g2_mux2_1 _16571_ (.A0(_10604_),
    .A1(_00293_),
    .S(net735),
    .X(_00602_));
 sg13g2_mux2_1 _16572_ (.A0(net124),
    .A1(_00294_),
    .S(net735),
    .X(_00603_));
 sg13g2_mux2_1 _16573_ (.A0(_10345_),
    .A1(_00295_),
    .S(net735),
    .X(_00604_));
 sg13g2_mux2_1 _16574_ (.A0(net130),
    .A1(_00296_),
    .S(net735),
    .X(_00605_));
 sg13g2_mux2_1 _16575_ (.A0(net129),
    .A1(_00297_),
    .S(net735),
    .X(_00606_));
 sg13g2_mux2_1 _16576_ (.A0(net123),
    .A1(_00298_),
    .S(net735),
    .X(_00607_));
 sg13g2_mux2_1 _16577_ (.A0(_10646_),
    .A1(_00299_),
    .S(net735),
    .X(_00608_));
 sg13g2_mux2_1 _16578_ (.A0(_10480_),
    .A1(_00300_),
    .S(_10662_),
    .X(_00609_));
 sg13g2_mux2_1 _16579_ (.A0(net305),
    .A1(_00301_),
    .S(net736),
    .X(_00610_));
 sg13g2_mux2_1 _16580_ (.A0(_10648_),
    .A1(_00302_),
    .S(_10653_),
    .X(_00611_));
 sg13g2_nand2_1 _16581_ (.Y(_10663_),
    .A(_10524_),
    .B(net763));
 sg13g2_buf_1 _16582_ (.A(_10663_),
    .X(_10664_));
 sg13g2_buf_1 _16583_ (.A(net650),
    .X(_10665_));
 sg13g2_buf_1 _16584_ (.A(_10663_),
    .X(_10666_));
 sg13g2_nand2_1 _16585_ (.Y(_10667_),
    .A(\top_ihp.oisc.regs[14][0] ),
    .B(net649));
 sg13g2_o21ai_1 _16586_ (.B1(_10667_),
    .Y(_00612_),
    .A1(net53),
    .A2(net513));
 sg13g2_nand2_1 _16587_ (.Y(_10668_),
    .A(\top_ihp.oisc.regs[14][10] ),
    .B(net649));
 sg13g2_o21ai_1 _16588_ (.B1(_10668_),
    .Y(_00613_),
    .A1(net155),
    .A2(net513));
 sg13g2_nand2_1 _16589_ (.Y(_10669_),
    .A(\top_ihp.oisc.regs[14][11] ),
    .B(net649));
 sg13g2_o21ai_1 _16590_ (.B1(_10669_),
    .Y(_00614_),
    .A1(net154),
    .A2(net513));
 sg13g2_nand2_1 _16591_ (.Y(_10670_),
    .A(\top_ihp.oisc.regs[14][12] ),
    .B(_10666_));
 sg13g2_o21ai_1 _16592_ (.B1(_10670_),
    .Y(_00615_),
    .A1(net137),
    .A2(_10665_));
 sg13g2_nand2_1 _16593_ (.Y(_10671_),
    .A(\top_ihp.oisc.regs[14][13] ),
    .B(net649));
 sg13g2_o21ai_1 _16594_ (.B1(_10671_),
    .Y(_00616_),
    .A1(net331),
    .A2(net513));
 sg13g2_nand2_1 _16595_ (.Y(_10672_),
    .A(\top_ihp.oisc.regs[14][14] ),
    .B(net649));
 sg13g2_o21ai_1 _16596_ (.B1(_10672_),
    .Y(_00617_),
    .A1(net136),
    .A2(net513));
 sg13g2_nand2_1 _16597_ (.Y(_10673_),
    .A(\top_ihp.oisc.regs[14][15] ),
    .B(net649));
 sg13g2_o21ai_1 _16598_ (.B1(_10673_),
    .Y(_00618_),
    .A1(net135),
    .A2(net513));
 sg13g2_nand2_1 _16599_ (.Y(_10674_),
    .A(\top_ihp.oisc.regs[14][16] ),
    .B(_10666_));
 sg13g2_o21ai_1 _16600_ (.B1(_10674_),
    .Y(_00619_),
    .A1(net150),
    .A2(_10665_));
 sg13g2_buf_1 _16601_ (.A(net650),
    .X(_10675_));
 sg13g2_nand2_1 _16602_ (.Y(_10676_),
    .A(\top_ihp.oisc.regs[14][17] ),
    .B(net512));
 sg13g2_o21ai_1 _16603_ (.B1(_10676_),
    .Y(_00620_),
    .A1(net328),
    .A2(net513));
 sg13g2_nand2_1 _16604_ (.Y(_10677_),
    .A(\top_ihp.oisc.regs[14][18] ),
    .B(net512));
 sg13g2_o21ai_1 _16605_ (.B1(_10677_),
    .Y(_00621_),
    .A1(net327),
    .A2(net513));
 sg13g2_buf_1 _16606_ (.A(net650),
    .X(_10678_));
 sg13g2_nand2_1 _16607_ (.Y(_10679_),
    .A(\top_ihp.oisc.regs[14][19] ),
    .B(net512));
 sg13g2_o21ai_1 _16608_ (.B1(_10679_),
    .Y(_00622_),
    .A1(net326),
    .A2(net511));
 sg13g2_nand2_1 _16609_ (.Y(_10680_),
    .A(\top_ihp.oisc.regs[14][1] ),
    .B(_10675_));
 sg13g2_o21ai_1 _16610_ (.B1(_10680_),
    .Y(_00623_),
    .A1(net134),
    .A2(_10678_));
 sg13g2_nand2_1 _16611_ (.Y(_10681_),
    .A(\top_ihp.oisc.regs[14][20] ),
    .B(net512));
 sg13g2_o21ai_1 _16612_ (.B1(_10681_),
    .Y(_00624_),
    .A1(net324),
    .A2(net511));
 sg13g2_nand2_1 _16613_ (.Y(_10682_),
    .A(\top_ihp.oisc.regs[14][21] ),
    .B(net512));
 sg13g2_o21ai_1 _16614_ (.B1(_10682_),
    .Y(_00625_),
    .A1(net323),
    .A2(net511));
 sg13g2_nand2_1 _16615_ (.Y(_10683_),
    .A(\top_ihp.oisc.regs[14][22] ),
    .B(net512));
 sg13g2_o21ai_1 _16616_ (.B1(_10683_),
    .Y(_00626_),
    .A1(net133),
    .A2(net511));
 sg13g2_nand2_1 _16617_ (.Y(_10684_),
    .A(\top_ihp.oisc.regs[14][23] ),
    .B(net512));
 sg13g2_o21ai_1 _16618_ (.B1(_10684_),
    .Y(_00627_),
    .A1(net321),
    .A2(net511));
 sg13g2_nand2_1 _16619_ (.Y(_10685_),
    .A(\top_ihp.oisc.regs[14][24] ),
    .B(_10675_));
 sg13g2_o21ai_1 _16620_ (.B1(_10685_),
    .Y(_00628_),
    .A1(net320),
    .A2(_10678_));
 sg13g2_nand2_1 _16621_ (.Y(_10686_),
    .A(\top_ihp.oisc.regs[14][25] ),
    .B(net512));
 sg13g2_o21ai_1 _16622_ (.B1(_10686_),
    .Y(_00629_),
    .A1(net132),
    .A2(net511));
 sg13g2_buf_8 _16623_ (.A(net650),
    .X(_10687_));
 sg13g2_nand2_1 _16624_ (.Y(_10688_),
    .A(\top_ihp.oisc.regs[14][26] ),
    .B(_10687_));
 sg13g2_o21ai_1 _16625_ (.B1(_10688_),
    .Y(_00630_),
    .A1(net146),
    .A2(net511));
 sg13g2_nand2_1 _16626_ (.Y(_10689_),
    .A(\top_ihp.oisc.regs[14][27] ),
    .B(net510));
 sg13g2_o21ai_1 _16627_ (.B1(_10689_),
    .Y(_00631_),
    .A1(net318),
    .A2(net511));
 sg13g2_buf_8 _16628_ (.A(net650),
    .X(_10690_));
 sg13g2_nand2_1 _16629_ (.Y(_10691_),
    .A(\top_ihp.oisc.regs[14][28] ),
    .B(net510));
 sg13g2_o21ai_1 _16630_ (.B1(_10691_),
    .Y(_00632_),
    .A1(net525),
    .A2(net509));
 sg13g2_nand2_1 _16631_ (.Y(_10692_),
    .A(\top_ihp.oisc.regs[14][29] ),
    .B(net510));
 sg13g2_o21ai_1 _16632_ (.B1(_10692_),
    .Y(_00633_),
    .A1(net317),
    .A2(net509));
 sg13g2_nand2_1 _16633_ (.Y(_10693_),
    .A(\top_ihp.oisc.regs[14][2] ),
    .B(_10687_));
 sg13g2_o21ai_1 _16634_ (.B1(_10693_),
    .Y(_00634_),
    .A1(net145),
    .A2(_10690_));
 sg13g2_nand2_1 _16635_ (.Y(_10694_),
    .A(\top_ihp.oisc.regs[14][30] ),
    .B(net510));
 sg13g2_o21ai_1 _16636_ (.B1(_10694_),
    .Y(_00635_),
    .A1(net144),
    .A2(net509));
 sg13g2_nand2_1 _16637_ (.Y(_10695_),
    .A(\top_ihp.oisc.regs[14][31] ),
    .B(net510));
 sg13g2_o21ai_1 _16638_ (.B1(_10695_),
    .Y(_00636_),
    .A1(net52),
    .A2(net509));
 sg13g2_nand2_1 _16639_ (.Y(_10696_),
    .A(\top_ihp.oisc.regs[14][3] ),
    .B(net510));
 sg13g2_o21ai_1 _16640_ (.B1(_10696_),
    .Y(_00637_),
    .A1(net143),
    .A2(net509));
 sg13g2_nand2_1 _16641_ (.Y(_10697_),
    .A(\top_ihp.oisc.regs[14][4] ),
    .B(net510));
 sg13g2_o21ai_1 _16642_ (.B1(_10697_),
    .Y(_00638_),
    .A1(net142),
    .A2(net509));
 sg13g2_nand2_1 _16643_ (.Y(_10698_),
    .A(\top_ihp.oisc.regs[14][5] ),
    .B(net510));
 sg13g2_o21ai_1 _16644_ (.B1(_10698_),
    .Y(_00639_),
    .A1(net141),
    .A2(net509));
 sg13g2_nand2_1 _16645_ (.Y(_10699_),
    .A(\top_ihp.oisc.regs[14][6] ),
    .B(net650));
 sg13g2_o21ai_1 _16646_ (.B1(_10699_),
    .Y(_00640_),
    .A1(net140),
    .A2(_10690_));
 sg13g2_nand2_1 _16647_ (.Y(_10700_),
    .A(\top_ihp.oisc.regs[14][7] ),
    .B(net650));
 sg13g2_o21ai_1 _16648_ (.B1(_10700_),
    .Y(_00641_),
    .A1(net139),
    .A2(net509));
 sg13g2_nand2_1 _16649_ (.Y(_10701_),
    .A(\top_ihp.oisc.regs[14][8] ),
    .B(_10664_));
 sg13g2_o21ai_1 _16650_ (.B1(_10701_),
    .Y(_00642_),
    .A1(net316),
    .A2(net649));
 sg13g2_nand2_1 _16651_ (.Y(_10702_),
    .A(\top_ihp.oisc.regs[14][9] ),
    .B(net650));
 sg13g2_o21ai_1 _16652_ (.B1(_10702_),
    .Y(_00643_),
    .A1(net138),
    .A2(net649));
 sg13g2_nand2_1 _16653_ (.Y(_10703_),
    .A(_10572_),
    .B(net763));
 sg13g2_buf_1 _16654_ (.A(_10703_),
    .X(_10704_));
 sg13g2_buf_1 _16655_ (.A(net716),
    .X(_10705_));
 sg13g2_buf_1 _16656_ (.A(_10703_),
    .X(_10706_));
 sg13g2_nand2_1 _16657_ (.Y(_10707_),
    .A(\top_ihp.oisc.regs[15][0] ),
    .B(net715));
 sg13g2_o21ai_1 _16658_ (.B1(_10707_),
    .Y(_00644_),
    .A1(net53),
    .A2(net648));
 sg13g2_nand2_1 _16659_ (.Y(_10708_),
    .A(\top_ihp.oisc.regs[15][10] ),
    .B(net715));
 sg13g2_o21ai_1 _16660_ (.B1(_10708_),
    .Y(_00645_),
    .A1(net155),
    .A2(net648));
 sg13g2_nand2_1 _16661_ (.Y(_10709_),
    .A(\top_ihp.oisc.regs[15][11] ),
    .B(net715));
 sg13g2_o21ai_1 _16662_ (.B1(_10709_),
    .Y(_00646_),
    .A1(net154),
    .A2(net648));
 sg13g2_nand2_1 _16663_ (.Y(_10710_),
    .A(\top_ihp.oisc.regs[15][12] ),
    .B(net715));
 sg13g2_o21ai_1 _16664_ (.B1(_10710_),
    .Y(_00647_),
    .A1(net137),
    .A2(net648));
 sg13g2_nand2_1 _16665_ (.Y(_10711_),
    .A(\top_ihp.oisc.regs[15][13] ),
    .B(net715));
 sg13g2_o21ai_1 _16666_ (.B1(_10711_),
    .Y(_00648_),
    .A1(net331),
    .A2(net648));
 sg13g2_nand2_1 _16667_ (.Y(_10712_),
    .A(\top_ihp.oisc.regs[15][14] ),
    .B(net715));
 sg13g2_o21ai_1 _16668_ (.B1(_10712_),
    .Y(_00649_),
    .A1(net136),
    .A2(net648));
 sg13g2_nand2_1 _16669_ (.Y(_10713_),
    .A(\top_ihp.oisc.regs[15][15] ),
    .B(net715));
 sg13g2_o21ai_1 _16670_ (.B1(_10713_),
    .Y(_00650_),
    .A1(net135),
    .A2(_10705_));
 sg13g2_nand2_1 _16671_ (.Y(_10714_),
    .A(\top_ihp.oisc.regs[15][16] ),
    .B(net715));
 sg13g2_o21ai_1 _16672_ (.B1(_10714_),
    .Y(_00651_),
    .A1(net150),
    .A2(net648));
 sg13g2_buf_1 _16673_ (.A(net716),
    .X(_10715_));
 sg13g2_nand2_1 _16674_ (.Y(_10716_),
    .A(\top_ihp.oisc.regs[15][17] ),
    .B(_10715_));
 sg13g2_o21ai_1 _16675_ (.B1(_10716_),
    .Y(_00652_),
    .A1(net328),
    .A2(_10705_));
 sg13g2_nand2_1 _16676_ (.Y(_10717_),
    .A(\top_ihp.oisc.regs[15][18] ),
    .B(net647));
 sg13g2_o21ai_1 _16677_ (.B1(_10717_),
    .Y(_00653_),
    .A1(net327),
    .A2(net648));
 sg13g2_buf_1 _16678_ (.A(net716),
    .X(_10718_));
 sg13g2_nand2_1 _16679_ (.Y(_10719_),
    .A(\top_ihp.oisc.regs[15][19] ),
    .B(net647));
 sg13g2_o21ai_1 _16680_ (.B1(_10719_),
    .Y(_00654_),
    .A1(net326),
    .A2(net646));
 sg13g2_nand2_1 _16681_ (.Y(_10720_),
    .A(\top_ihp.oisc.regs[15][1] ),
    .B(_10715_));
 sg13g2_o21ai_1 _16682_ (.B1(_10720_),
    .Y(_00655_),
    .A1(net134),
    .A2(_10718_));
 sg13g2_nand2_1 _16683_ (.Y(_10721_),
    .A(\top_ihp.oisc.regs[15][20] ),
    .B(net647));
 sg13g2_o21ai_1 _16684_ (.B1(_10721_),
    .Y(_00656_),
    .A1(net653),
    .A2(_10718_));
 sg13g2_nand2_1 _16685_ (.Y(_10722_),
    .A(\top_ihp.oisc.regs[15][21] ),
    .B(net647));
 sg13g2_o21ai_1 _16686_ (.B1(_10722_),
    .Y(_00657_),
    .A1(net323),
    .A2(net646));
 sg13g2_nand2_1 _16687_ (.Y(_10723_),
    .A(\top_ihp.oisc.regs[15][22] ),
    .B(net647));
 sg13g2_o21ai_1 _16688_ (.B1(_10723_),
    .Y(_00658_),
    .A1(net133),
    .A2(net646));
 sg13g2_nand2_1 _16689_ (.Y(_10724_),
    .A(\top_ihp.oisc.regs[15][23] ),
    .B(net647));
 sg13g2_o21ai_1 _16690_ (.B1(_10724_),
    .Y(_00659_),
    .A1(net321),
    .A2(net646));
 sg13g2_nand2_1 _16691_ (.Y(_10725_),
    .A(\top_ihp.oisc.regs[15][24] ),
    .B(net647));
 sg13g2_o21ai_1 _16692_ (.B1(_10725_),
    .Y(_00660_),
    .A1(net320),
    .A2(net646));
 sg13g2_nand2_1 _16693_ (.Y(_10726_),
    .A(\top_ihp.oisc.regs[15][25] ),
    .B(net647));
 sg13g2_o21ai_1 _16694_ (.B1(_10726_),
    .Y(_00661_),
    .A1(net132),
    .A2(net646));
 sg13g2_buf_1 _16695_ (.A(net716),
    .X(_10727_));
 sg13g2_nand2_1 _16696_ (.Y(_10728_),
    .A(\top_ihp.oisc.regs[15][26] ),
    .B(net645));
 sg13g2_o21ai_1 _16697_ (.B1(_10728_),
    .Y(_00662_),
    .A1(net146),
    .A2(net646));
 sg13g2_nand2_1 _16698_ (.Y(_10729_),
    .A(\top_ihp.oisc.regs[15][27] ),
    .B(net645));
 sg13g2_o21ai_1 _16699_ (.B1(_10729_),
    .Y(_00663_),
    .A1(net318),
    .A2(net646));
 sg13g2_buf_1 _16700_ (.A(net716),
    .X(_10730_));
 sg13g2_nand2_1 _16701_ (.Y(_10731_),
    .A(\top_ihp.oisc.regs[15][28] ),
    .B(net645));
 sg13g2_o21ai_1 _16702_ (.B1(_10731_),
    .Y(_00664_),
    .A1(net525),
    .A2(net644));
 sg13g2_nand2_1 _16703_ (.Y(_10732_),
    .A(\top_ihp.oisc.regs[15][29] ),
    .B(_10727_));
 sg13g2_o21ai_1 _16704_ (.B1(_10732_),
    .Y(_00665_),
    .A1(net317),
    .A2(_10730_));
 sg13g2_nand2_1 _16705_ (.Y(_10733_),
    .A(\top_ihp.oisc.regs[15][2] ),
    .B(_10727_));
 sg13g2_o21ai_1 _16706_ (.B1(_10733_),
    .Y(_00666_),
    .A1(net145),
    .A2(net644));
 sg13g2_nand2_1 _16707_ (.Y(_10734_),
    .A(\top_ihp.oisc.regs[15][30] ),
    .B(net645));
 sg13g2_o21ai_1 _16708_ (.B1(_10734_),
    .Y(_00667_),
    .A1(net144),
    .A2(net644));
 sg13g2_nand2_1 _16709_ (.Y(_10735_),
    .A(\top_ihp.oisc.regs[15][31] ),
    .B(net645));
 sg13g2_o21ai_1 _16710_ (.B1(_10735_),
    .Y(_00668_),
    .A1(net315),
    .A2(net644));
 sg13g2_nand2_1 _16711_ (.Y(_10736_),
    .A(\top_ihp.oisc.regs[15][3] ),
    .B(net645));
 sg13g2_o21ai_1 _16712_ (.B1(_10736_),
    .Y(_00669_),
    .A1(net143),
    .A2(net644));
 sg13g2_nand2_1 _16713_ (.Y(_10737_),
    .A(\top_ihp.oisc.regs[15][4] ),
    .B(net645));
 sg13g2_o21ai_1 _16714_ (.B1(_10737_),
    .Y(_00670_),
    .A1(net142),
    .A2(net644));
 sg13g2_nand2_1 _16715_ (.Y(_10738_),
    .A(\top_ihp.oisc.regs[15][5] ),
    .B(net645));
 sg13g2_o21ai_1 _16716_ (.B1(_10738_),
    .Y(_00671_),
    .A1(net141),
    .A2(net644));
 sg13g2_nand2_1 _16717_ (.Y(_10739_),
    .A(\top_ihp.oisc.regs[15][6] ),
    .B(net716));
 sg13g2_o21ai_1 _16718_ (.B1(_10739_),
    .Y(_00672_),
    .A1(net140),
    .A2(_10730_));
 sg13g2_nand2_1 _16719_ (.Y(_10740_),
    .A(\top_ihp.oisc.regs[15][7] ),
    .B(net716));
 sg13g2_o21ai_1 _16720_ (.B1(_10740_),
    .Y(_00673_),
    .A1(net518),
    .A2(net644));
 sg13g2_nand2_1 _16721_ (.Y(_10741_),
    .A(\top_ihp.oisc.regs[15][8] ),
    .B(_10704_));
 sg13g2_o21ai_1 _16722_ (.B1(_10741_),
    .Y(_00674_),
    .A1(net316),
    .A2(_10706_));
 sg13g2_nand2_1 _16723_ (.Y(_10742_),
    .A(\top_ihp.oisc.regs[15][9] ),
    .B(net716));
 sg13g2_o21ai_1 _16724_ (.B1(_10742_),
    .Y(_00675_),
    .A1(net138),
    .A2(_10706_));
 sg13g2_buf_1 _16725_ (.A(\top_ihp.oisc.regs[16][0] ),
    .X(_00676_));
 sg13g2_buf_1 _16726_ (.A(\top_ihp.oisc.regs[16][10] ),
    .X(_00677_));
 sg13g2_buf_1 _16727_ (.A(\top_ihp.oisc.regs[16][11] ),
    .X(_00678_));
 sg13g2_buf_1 _16728_ (.A(\top_ihp.oisc.regs[16][12] ),
    .X(_00679_));
 sg13g2_buf_1 _16729_ (.A(\top_ihp.oisc.regs[16][13] ),
    .X(_00680_));
 sg13g2_buf_1 _16730_ (.A(\top_ihp.oisc.regs[16][14] ),
    .X(_00681_));
 sg13g2_buf_1 _16731_ (.A(\top_ihp.oisc.regs[16][15] ),
    .X(_00682_));
 sg13g2_buf_1 _16732_ (.A(\top_ihp.oisc.regs[16][16] ),
    .X(_00683_));
 sg13g2_buf_1 _16733_ (.A(\top_ihp.oisc.regs[16][17] ),
    .X(_00684_));
 sg13g2_buf_1 _16734_ (.A(\top_ihp.oisc.regs[16][18] ),
    .X(_00685_));
 sg13g2_buf_1 _16735_ (.A(\top_ihp.oisc.regs[16][19] ),
    .X(_00686_));
 sg13g2_buf_1 _16736_ (.A(\top_ihp.oisc.regs[16][1] ),
    .X(_00687_));
 sg13g2_buf_1 _16737_ (.A(\top_ihp.oisc.regs[16][20] ),
    .X(_00688_));
 sg13g2_buf_1 _16738_ (.A(\top_ihp.oisc.regs[16][21] ),
    .X(_00689_));
 sg13g2_buf_1 _16739_ (.A(\top_ihp.oisc.regs[16][22] ),
    .X(_00690_));
 sg13g2_buf_1 _16740_ (.A(\top_ihp.oisc.regs[16][23] ),
    .X(_00691_));
 sg13g2_buf_1 _16741_ (.A(\top_ihp.oisc.regs[16][24] ),
    .X(_00692_));
 sg13g2_buf_1 _16742_ (.A(\top_ihp.oisc.regs[16][25] ),
    .X(_00693_));
 sg13g2_buf_1 _16743_ (.A(\top_ihp.oisc.regs[16][26] ),
    .X(_00694_));
 sg13g2_buf_1 _16744_ (.A(\top_ihp.oisc.regs[16][27] ),
    .X(_00695_));
 sg13g2_buf_1 _16745_ (.A(\top_ihp.oisc.regs[16][28] ),
    .X(_00696_));
 sg13g2_buf_1 _16746_ (.A(\top_ihp.oisc.regs[16][29] ),
    .X(_00697_));
 sg13g2_buf_1 _16747_ (.A(\top_ihp.oisc.regs[16][2] ),
    .X(_00698_));
 sg13g2_buf_1 _16748_ (.A(\top_ihp.oisc.regs[16][30] ),
    .X(_00699_));
 sg13g2_buf_1 _16749_ (.A(\top_ihp.oisc.regs[16][31] ),
    .X(_00700_));
 sg13g2_buf_1 _16750_ (.A(\top_ihp.oisc.regs[16][3] ),
    .X(_00701_));
 sg13g2_buf_1 _16751_ (.A(\top_ihp.oisc.regs[16][4] ),
    .X(_00702_));
 sg13g2_buf_1 _16752_ (.A(\top_ihp.oisc.regs[16][5] ),
    .X(_00703_));
 sg13g2_buf_1 _16753_ (.A(\top_ihp.oisc.regs[16][6] ),
    .X(_00704_));
 sg13g2_buf_1 _16754_ (.A(\top_ihp.oisc.regs[16][7] ),
    .X(_00705_));
 sg13g2_buf_1 _16755_ (.A(\top_ihp.oisc.regs[16][8] ),
    .X(_00706_));
 sg13g2_buf_1 _16756_ (.A(\top_ihp.oisc.regs[16][9] ),
    .X(_00707_));
 sg13g2_buf_1 _16757_ (.A(\top_ihp.oisc.regs[17][0] ),
    .X(_00708_));
 sg13g2_buf_1 _16758_ (.A(\top_ihp.oisc.regs[17][10] ),
    .X(_00709_));
 sg13g2_buf_1 _16759_ (.A(\top_ihp.oisc.regs[17][11] ),
    .X(_00710_));
 sg13g2_buf_1 _16760_ (.A(\top_ihp.oisc.regs[17][12] ),
    .X(_00711_));
 sg13g2_buf_1 _16761_ (.A(\top_ihp.oisc.regs[17][13] ),
    .X(_00712_));
 sg13g2_buf_1 _16762_ (.A(\top_ihp.oisc.regs[17][14] ),
    .X(_00713_));
 sg13g2_buf_1 _16763_ (.A(\top_ihp.oisc.regs[17][15] ),
    .X(_00714_));
 sg13g2_buf_1 _16764_ (.A(\top_ihp.oisc.regs[17][16] ),
    .X(_00715_));
 sg13g2_buf_1 _16765_ (.A(\top_ihp.oisc.regs[17][17] ),
    .X(_00716_));
 sg13g2_buf_1 _16766_ (.A(\top_ihp.oisc.regs[17][18] ),
    .X(_00717_));
 sg13g2_buf_1 _16767_ (.A(\top_ihp.oisc.regs[17][19] ),
    .X(_00718_));
 sg13g2_buf_1 _16768_ (.A(\top_ihp.oisc.regs[17][1] ),
    .X(_00719_));
 sg13g2_buf_1 _16769_ (.A(\top_ihp.oisc.regs[17][20] ),
    .X(_00720_));
 sg13g2_buf_1 _16770_ (.A(\top_ihp.oisc.regs[17][21] ),
    .X(_00721_));
 sg13g2_buf_1 _16771_ (.A(\top_ihp.oisc.regs[17][22] ),
    .X(_00722_));
 sg13g2_buf_1 _16772_ (.A(\top_ihp.oisc.regs[17][23] ),
    .X(_00723_));
 sg13g2_buf_1 _16773_ (.A(\top_ihp.oisc.regs[17][24] ),
    .X(_00724_));
 sg13g2_buf_1 _16774_ (.A(\top_ihp.oisc.regs[17][25] ),
    .X(_00725_));
 sg13g2_buf_1 _16775_ (.A(\top_ihp.oisc.regs[17][26] ),
    .X(_00726_));
 sg13g2_buf_1 _16776_ (.A(\top_ihp.oisc.regs[17][27] ),
    .X(_00727_));
 sg13g2_buf_1 _16777_ (.A(\top_ihp.oisc.regs[17][28] ),
    .X(_00728_));
 sg13g2_buf_1 _16778_ (.A(\top_ihp.oisc.regs[17][29] ),
    .X(_00729_));
 sg13g2_buf_1 _16779_ (.A(\top_ihp.oisc.regs[17][2] ),
    .X(_00730_));
 sg13g2_buf_1 _16780_ (.A(\top_ihp.oisc.regs[17][30] ),
    .X(_00731_));
 sg13g2_buf_1 _16781_ (.A(\top_ihp.oisc.regs[17][31] ),
    .X(_00732_));
 sg13g2_buf_1 _16782_ (.A(\top_ihp.oisc.regs[17][3] ),
    .X(_00733_));
 sg13g2_buf_1 _16783_ (.A(\top_ihp.oisc.regs[17][4] ),
    .X(_00734_));
 sg13g2_buf_1 _16784_ (.A(\top_ihp.oisc.regs[17][5] ),
    .X(_00735_));
 sg13g2_buf_1 _16785_ (.A(\top_ihp.oisc.regs[17][6] ),
    .X(_00736_));
 sg13g2_buf_1 _16786_ (.A(\top_ihp.oisc.regs[17][7] ),
    .X(_00737_));
 sg13g2_buf_1 _16787_ (.A(\top_ihp.oisc.regs[17][8] ),
    .X(_00738_));
 sg13g2_buf_1 _16788_ (.A(\top_ihp.oisc.regs[17][9] ),
    .X(_00739_));
 sg13g2_buf_1 _16789_ (.A(\top_ihp.oisc.regs[18][0] ),
    .X(_00740_));
 sg13g2_buf_1 _16790_ (.A(\top_ihp.oisc.regs[18][10] ),
    .X(_00741_));
 sg13g2_buf_1 _16791_ (.A(\top_ihp.oisc.regs[18][11] ),
    .X(_00742_));
 sg13g2_buf_1 _16792_ (.A(\top_ihp.oisc.regs[18][12] ),
    .X(_00743_));
 sg13g2_buf_1 _16793_ (.A(\top_ihp.oisc.regs[18][13] ),
    .X(_00744_));
 sg13g2_buf_1 _16794_ (.A(\top_ihp.oisc.regs[18][14] ),
    .X(_00745_));
 sg13g2_buf_1 _16795_ (.A(\top_ihp.oisc.regs[18][15] ),
    .X(_00746_));
 sg13g2_buf_1 _16796_ (.A(\top_ihp.oisc.regs[18][16] ),
    .X(_00747_));
 sg13g2_buf_1 _16797_ (.A(\top_ihp.oisc.regs[18][17] ),
    .X(_00748_));
 sg13g2_buf_1 _16798_ (.A(\top_ihp.oisc.regs[18][18] ),
    .X(_00749_));
 sg13g2_buf_1 _16799_ (.A(\top_ihp.oisc.regs[18][19] ),
    .X(_00750_));
 sg13g2_buf_1 _16800_ (.A(\top_ihp.oisc.regs[18][1] ),
    .X(_00751_));
 sg13g2_buf_1 _16801_ (.A(\top_ihp.oisc.regs[18][20] ),
    .X(_00752_));
 sg13g2_buf_1 _16802_ (.A(\top_ihp.oisc.regs[18][21] ),
    .X(_00753_));
 sg13g2_buf_1 _16803_ (.A(\top_ihp.oisc.regs[18][22] ),
    .X(_00754_));
 sg13g2_buf_1 _16804_ (.A(\top_ihp.oisc.regs[18][23] ),
    .X(_00755_));
 sg13g2_buf_1 _16805_ (.A(\top_ihp.oisc.regs[18][24] ),
    .X(_00756_));
 sg13g2_buf_1 _16806_ (.A(\top_ihp.oisc.regs[18][25] ),
    .X(_00757_));
 sg13g2_buf_1 _16807_ (.A(\top_ihp.oisc.regs[18][26] ),
    .X(_00758_));
 sg13g2_buf_1 _16808_ (.A(\top_ihp.oisc.regs[18][27] ),
    .X(_00759_));
 sg13g2_buf_1 _16809_ (.A(\top_ihp.oisc.regs[18][28] ),
    .X(_00760_));
 sg13g2_buf_1 _16810_ (.A(\top_ihp.oisc.regs[18][29] ),
    .X(_00761_));
 sg13g2_buf_1 _16811_ (.A(\top_ihp.oisc.regs[18][2] ),
    .X(_00762_));
 sg13g2_buf_1 _16812_ (.A(\top_ihp.oisc.regs[18][30] ),
    .X(_00763_));
 sg13g2_buf_1 _16813_ (.A(\top_ihp.oisc.regs[18][31] ),
    .X(_00764_));
 sg13g2_buf_1 _16814_ (.A(\top_ihp.oisc.regs[18][3] ),
    .X(_00765_));
 sg13g2_buf_1 _16815_ (.A(\top_ihp.oisc.regs[18][4] ),
    .X(_00766_));
 sg13g2_buf_1 _16816_ (.A(\top_ihp.oisc.regs[18][5] ),
    .X(_00767_));
 sg13g2_buf_1 _16817_ (.A(\top_ihp.oisc.regs[18][6] ),
    .X(_00768_));
 sg13g2_buf_1 _16818_ (.A(\top_ihp.oisc.regs[18][7] ),
    .X(_00769_));
 sg13g2_buf_1 _16819_ (.A(\top_ihp.oisc.regs[18][8] ),
    .X(_00770_));
 sg13g2_buf_1 _16820_ (.A(\top_ihp.oisc.regs[18][9] ),
    .X(_00771_));
 sg13g2_buf_1 _16821_ (.A(\top_ihp.oisc.regs[19][0] ),
    .X(_00772_));
 sg13g2_buf_1 _16822_ (.A(\top_ihp.oisc.regs[19][10] ),
    .X(_00773_));
 sg13g2_buf_1 _16823_ (.A(\top_ihp.oisc.regs[19][11] ),
    .X(_00774_));
 sg13g2_buf_1 _16824_ (.A(\top_ihp.oisc.regs[19][12] ),
    .X(_00775_));
 sg13g2_buf_1 _16825_ (.A(\top_ihp.oisc.regs[19][13] ),
    .X(_00776_));
 sg13g2_buf_1 _16826_ (.A(\top_ihp.oisc.regs[19][14] ),
    .X(_00777_));
 sg13g2_buf_1 _16827_ (.A(\top_ihp.oisc.regs[19][15] ),
    .X(_00778_));
 sg13g2_buf_1 _16828_ (.A(\top_ihp.oisc.regs[19][16] ),
    .X(_00779_));
 sg13g2_buf_1 _16829_ (.A(\top_ihp.oisc.regs[19][17] ),
    .X(_00780_));
 sg13g2_buf_1 _16830_ (.A(\top_ihp.oisc.regs[19][18] ),
    .X(_00781_));
 sg13g2_buf_1 _16831_ (.A(\top_ihp.oisc.regs[19][19] ),
    .X(_00782_));
 sg13g2_buf_1 _16832_ (.A(\top_ihp.oisc.regs[19][1] ),
    .X(_00783_));
 sg13g2_buf_1 _16833_ (.A(\top_ihp.oisc.regs[19][20] ),
    .X(_00784_));
 sg13g2_buf_1 _16834_ (.A(\top_ihp.oisc.regs[19][21] ),
    .X(_00785_));
 sg13g2_buf_1 _16835_ (.A(\top_ihp.oisc.regs[19][22] ),
    .X(_00786_));
 sg13g2_buf_1 _16836_ (.A(\top_ihp.oisc.regs[19][23] ),
    .X(_00787_));
 sg13g2_buf_1 _16837_ (.A(\top_ihp.oisc.regs[19][24] ),
    .X(_00788_));
 sg13g2_buf_1 _16838_ (.A(\top_ihp.oisc.regs[19][25] ),
    .X(_00789_));
 sg13g2_buf_1 _16839_ (.A(\top_ihp.oisc.regs[19][26] ),
    .X(_00790_));
 sg13g2_buf_1 _16840_ (.A(\top_ihp.oisc.regs[19][27] ),
    .X(_00791_));
 sg13g2_buf_1 _16841_ (.A(\top_ihp.oisc.regs[19][28] ),
    .X(_00792_));
 sg13g2_buf_1 _16842_ (.A(\top_ihp.oisc.regs[19][29] ),
    .X(_00793_));
 sg13g2_buf_1 _16843_ (.A(\top_ihp.oisc.regs[19][2] ),
    .X(_00794_));
 sg13g2_buf_1 _16844_ (.A(\top_ihp.oisc.regs[19][30] ),
    .X(_00795_));
 sg13g2_buf_1 _16845_ (.A(\top_ihp.oisc.regs[19][31] ),
    .X(_00796_));
 sg13g2_buf_1 _16846_ (.A(\top_ihp.oisc.regs[19][3] ),
    .X(_00797_));
 sg13g2_buf_1 _16847_ (.A(\top_ihp.oisc.regs[19][4] ),
    .X(_00798_));
 sg13g2_buf_1 _16848_ (.A(\top_ihp.oisc.regs[19][5] ),
    .X(_00799_));
 sg13g2_buf_1 _16849_ (.A(\top_ihp.oisc.regs[19][6] ),
    .X(_00800_));
 sg13g2_buf_1 _16850_ (.A(\top_ihp.oisc.regs[19][7] ),
    .X(_00801_));
 sg13g2_buf_1 _16851_ (.A(\top_ihp.oisc.regs[19][8] ),
    .X(_00802_));
 sg13g2_buf_1 _16852_ (.A(\top_ihp.oisc.regs[19][9] ),
    .X(_00803_));
 sg13g2_nand2_1 _16853_ (.Y(_10743_),
    .A(net767),
    .B(_10651_));
 sg13g2_buf_1 _16854_ (.A(_10743_),
    .X(_10744_));
 sg13g2_buf_1 _16855_ (.A(net734),
    .X(_10745_));
 sg13g2_buf_1 _16856_ (.A(net734),
    .X(_10746_));
 sg13g2_nand2_1 _16857_ (.Y(_10747_),
    .A(\top_ihp.oisc.regs[1][0] ),
    .B(net713));
 sg13g2_o21ai_1 _16858_ (.B1(_10747_),
    .Y(_00804_),
    .A1(net53),
    .A2(net714));
 sg13g2_nand2_1 _16859_ (.Y(_10748_),
    .A(\top_ihp.oisc.regs[1][10] ),
    .B(net713));
 sg13g2_o21ai_1 _16860_ (.B1(_10748_),
    .Y(_00805_),
    .A1(net155),
    .A2(net714));
 sg13g2_nand2_1 _16861_ (.Y(_10749_),
    .A(\top_ihp.oisc.regs[1][11] ),
    .B(net713));
 sg13g2_o21ai_1 _16862_ (.B1(_10749_),
    .Y(_00806_),
    .A1(net154),
    .A2(net714));
 sg13g2_nand2_1 _16863_ (.Y(_10750_),
    .A(\top_ihp.oisc.regs[1][12] ),
    .B(net713));
 sg13g2_o21ai_1 _16864_ (.B1(_10750_),
    .Y(_00807_),
    .A1(net137),
    .A2(net714));
 sg13g2_nand2_1 _16865_ (.Y(_10751_),
    .A(\top_ihp.oisc.regs[1][13] ),
    .B(net713));
 sg13g2_o21ai_1 _16866_ (.B1(_10751_),
    .Y(_00808_),
    .A1(net331),
    .A2(net714));
 sg13g2_nand2_1 _16867_ (.Y(_10752_),
    .A(\top_ihp.oisc.regs[1][14] ),
    .B(net713));
 sg13g2_o21ai_1 _16868_ (.B1(_10752_),
    .Y(_00809_),
    .A1(net136),
    .A2(_10745_));
 sg13g2_nand2_1 _16869_ (.Y(_10753_),
    .A(\top_ihp.oisc.regs[1][15] ),
    .B(net713));
 sg13g2_o21ai_1 _16870_ (.B1(_10753_),
    .Y(_00810_),
    .A1(net135),
    .A2(net714));
 sg13g2_nand2_1 _16871_ (.Y(_10754_),
    .A(\top_ihp.oisc.regs[1][16] ),
    .B(_10746_));
 sg13g2_o21ai_1 _16872_ (.B1(_10754_),
    .Y(_00811_),
    .A1(net150),
    .A2(_10745_));
 sg13g2_buf_1 _16873_ (.A(net734),
    .X(_10755_));
 sg13g2_nand2_1 _16874_ (.Y(_10756_),
    .A(\top_ihp.oisc.regs[1][17] ),
    .B(net712));
 sg13g2_o21ai_1 _16875_ (.B1(_10756_),
    .Y(_00812_),
    .A1(net328),
    .A2(net714));
 sg13g2_nand2_1 _16876_ (.Y(_10757_),
    .A(\top_ihp.oisc.regs[1][18] ),
    .B(net712));
 sg13g2_o21ai_1 _16877_ (.B1(_10757_),
    .Y(_00813_),
    .A1(net327),
    .A2(net714));
 sg13g2_buf_1 _16878_ (.A(net734),
    .X(_10758_));
 sg13g2_nand2_1 _16879_ (.Y(_10759_),
    .A(\top_ihp.oisc.regs[1][19] ),
    .B(net712));
 sg13g2_o21ai_1 _16880_ (.B1(_10759_),
    .Y(_00814_),
    .A1(net326),
    .A2(net711));
 sg13g2_nand2_1 _16881_ (.Y(_10760_),
    .A(\top_ihp.oisc.regs[1][1] ),
    .B(net712));
 sg13g2_o21ai_1 _16882_ (.B1(_10760_),
    .Y(_00815_),
    .A1(net134),
    .A2(net711));
 sg13g2_nand2_1 _16883_ (.Y(_10761_),
    .A(\top_ihp.oisc.regs[1][20] ),
    .B(_10755_));
 sg13g2_o21ai_1 _16884_ (.B1(_10761_),
    .Y(_00816_),
    .A1(net653),
    .A2(_10758_));
 sg13g2_nand2_1 _16885_ (.Y(_10762_),
    .A(\top_ihp.oisc.regs[1][21] ),
    .B(net712));
 sg13g2_o21ai_1 _16886_ (.B1(_10762_),
    .Y(_00817_),
    .A1(net323),
    .A2(net711));
 sg13g2_nand2_1 _16887_ (.Y(_10763_),
    .A(\top_ihp.oisc.regs[1][22] ),
    .B(net712));
 sg13g2_o21ai_1 _16888_ (.B1(_10763_),
    .Y(_00818_),
    .A1(net133),
    .A2(net711));
 sg13g2_nand2_1 _16889_ (.Y(_10764_),
    .A(\top_ihp.oisc.regs[1][23] ),
    .B(net712));
 sg13g2_o21ai_1 _16890_ (.B1(_10764_),
    .Y(_00819_),
    .A1(net321),
    .A2(net711));
 sg13g2_nand2_1 _16891_ (.Y(_10765_),
    .A(\top_ihp.oisc.regs[1][24] ),
    .B(_10755_));
 sg13g2_o21ai_1 _16892_ (.B1(_10765_),
    .Y(_00820_),
    .A1(net320),
    .A2(_10758_));
 sg13g2_nand2_1 _16893_ (.Y(_10766_),
    .A(\top_ihp.oisc.regs[1][25] ),
    .B(net712));
 sg13g2_o21ai_1 _16894_ (.B1(_10766_),
    .Y(_00821_),
    .A1(net132),
    .A2(net711));
 sg13g2_buf_1 _16895_ (.A(net734),
    .X(_10767_));
 sg13g2_nand2_1 _16896_ (.Y(_10768_),
    .A(\top_ihp.oisc.regs[1][26] ),
    .B(net710));
 sg13g2_o21ai_1 _16897_ (.B1(_10768_),
    .Y(_00822_),
    .A1(net146),
    .A2(net711));
 sg13g2_nand2_1 _16898_ (.Y(_10769_),
    .A(\top_ihp.oisc.regs[1][27] ),
    .B(net710));
 sg13g2_o21ai_1 _16899_ (.B1(_10769_),
    .Y(_00823_),
    .A1(net318),
    .A2(net711));
 sg13g2_buf_1 _16900_ (.A(net734),
    .X(_10770_));
 sg13g2_nand2_1 _16901_ (.Y(_10771_),
    .A(\top_ihp.oisc.regs[1][28] ),
    .B(net710));
 sg13g2_o21ai_1 _16902_ (.B1(_10771_),
    .Y(_00824_),
    .A1(net525),
    .A2(net709));
 sg13g2_nand2_1 _16903_ (.Y(_10772_),
    .A(\top_ihp.oisc.regs[1][29] ),
    .B(net710));
 sg13g2_o21ai_1 _16904_ (.B1(_10772_),
    .Y(_00825_),
    .A1(net317),
    .A2(net709));
 sg13g2_nand2_1 _16905_ (.Y(_10773_),
    .A(\top_ihp.oisc.regs[1][2] ),
    .B(_10767_));
 sg13g2_o21ai_1 _16906_ (.B1(_10773_),
    .Y(_00826_),
    .A1(net145),
    .A2(_10770_));
 sg13g2_mux2_1 _16907_ (.A0(_10643_),
    .A1(_00303_),
    .S(net713),
    .X(_00827_));
 sg13g2_nand2_1 _16908_ (.Y(_10774_),
    .A(\top_ihp.oisc.regs[1][31] ),
    .B(net710));
 sg13g2_o21ai_1 _16909_ (.B1(_10774_),
    .Y(_00828_),
    .A1(net315),
    .A2(net709));
 sg13g2_nand2_1 _16910_ (.Y(_10775_),
    .A(\top_ihp.oisc.regs[1][3] ),
    .B(net710));
 sg13g2_o21ai_1 _16911_ (.B1(_10775_),
    .Y(_00829_),
    .A1(net143),
    .A2(net709));
 sg13g2_nand2_1 _16912_ (.Y(_10776_),
    .A(\top_ihp.oisc.regs[1][4] ),
    .B(net710));
 sg13g2_o21ai_1 _16913_ (.B1(_10776_),
    .Y(_00830_),
    .A1(net142),
    .A2(net709));
 sg13g2_nand2_1 _16914_ (.Y(_10777_),
    .A(\top_ihp.oisc.regs[1][5] ),
    .B(net710));
 sg13g2_o21ai_1 _16915_ (.B1(_10777_),
    .Y(_00831_),
    .A1(net141),
    .A2(net709));
 sg13g2_nand2_1 _16916_ (.Y(_10778_),
    .A(\top_ihp.oisc.regs[1][6] ),
    .B(_10767_));
 sg13g2_o21ai_1 _16917_ (.B1(_10778_),
    .Y(_00832_),
    .A1(net140),
    .A2(net709));
 sg13g2_nand2_1 _16918_ (.Y(_10779_),
    .A(\top_ihp.oisc.regs[1][7] ),
    .B(net734));
 sg13g2_o21ai_1 _16919_ (.B1(_10779_),
    .Y(_00833_),
    .A1(net518),
    .A2(_10770_));
 sg13g2_nand2_1 _16920_ (.Y(_10780_),
    .A(\top_ihp.oisc.regs[1][8] ),
    .B(_10744_));
 sg13g2_o21ai_1 _16921_ (.B1(_10780_),
    .Y(_00834_),
    .A1(net316),
    .A2(net709));
 sg13g2_nand2_1 _16922_ (.Y(_10781_),
    .A(\top_ihp.oisc.regs[1][9] ),
    .B(net734));
 sg13g2_o21ai_1 _16923_ (.B1(_10781_),
    .Y(_00835_),
    .A1(net138),
    .A2(_10746_));
 sg13g2_buf_1 _16924_ (.A(\top_ihp.oisc.regs[20][0] ),
    .X(_00836_));
 sg13g2_buf_1 _16925_ (.A(\top_ihp.oisc.regs[20][10] ),
    .X(_00837_));
 sg13g2_buf_1 _16926_ (.A(\top_ihp.oisc.regs[20][11] ),
    .X(_00838_));
 sg13g2_buf_1 _16927_ (.A(\top_ihp.oisc.regs[20][12] ),
    .X(_00839_));
 sg13g2_buf_1 _16928_ (.A(\top_ihp.oisc.regs[20][13] ),
    .X(_00840_));
 sg13g2_buf_1 _16929_ (.A(\top_ihp.oisc.regs[20][14] ),
    .X(_00841_));
 sg13g2_buf_1 _16930_ (.A(\top_ihp.oisc.regs[20][15] ),
    .X(_00842_));
 sg13g2_buf_1 _16931_ (.A(\top_ihp.oisc.regs[20][16] ),
    .X(_00843_));
 sg13g2_buf_1 _16932_ (.A(\top_ihp.oisc.regs[20][17] ),
    .X(_00844_));
 sg13g2_buf_1 _16933_ (.A(\top_ihp.oisc.regs[20][18] ),
    .X(_00845_));
 sg13g2_buf_1 _16934_ (.A(\top_ihp.oisc.regs[20][19] ),
    .X(_00846_));
 sg13g2_buf_1 _16935_ (.A(\top_ihp.oisc.regs[20][1] ),
    .X(_00847_));
 sg13g2_buf_1 _16936_ (.A(\top_ihp.oisc.regs[20][20] ),
    .X(_00848_));
 sg13g2_buf_1 _16937_ (.A(\top_ihp.oisc.regs[20][21] ),
    .X(_00849_));
 sg13g2_buf_1 _16938_ (.A(\top_ihp.oisc.regs[20][22] ),
    .X(_00850_));
 sg13g2_buf_1 _16939_ (.A(\top_ihp.oisc.regs[20][23] ),
    .X(_00851_));
 sg13g2_buf_1 _16940_ (.A(\top_ihp.oisc.regs[20][24] ),
    .X(_00852_));
 sg13g2_buf_1 _16941_ (.A(\top_ihp.oisc.regs[20][25] ),
    .X(_00853_));
 sg13g2_buf_1 _16942_ (.A(\top_ihp.oisc.regs[20][26] ),
    .X(_00854_));
 sg13g2_buf_1 _16943_ (.A(\top_ihp.oisc.regs[20][27] ),
    .X(_00855_));
 sg13g2_buf_1 _16944_ (.A(\top_ihp.oisc.regs[20][28] ),
    .X(_00856_));
 sg13g2_buf_1 _16945_ (.A(\top_ihp.oisc.regs[20][29] ),
    .X(_00857_));
 sg13g2_buf_1 _16946_ (.A(\top_ihp.oisc.regs[20][2] ),
    .X(_00858_));
 sg13g2_buf_1 _16947_ (.A(\top_ihp.oisc.regs[20][30] ),
    .X(_00859_));
 sg13g2_buf_1 _16948_ (.A(\top_ihp.oisc.regs[20][31] ),
    .X(_00860_));
 sg13g2_buf_1 _16949_ (.A(\top_ihp.oisc.regs[20][3] ),
    .X(_00861_));
 sg13g2_buf_1 _16950_ (.A(\top_ihp.oisc.regs[20][4] ),
    .X(_00862_));
 sg13g2_buf_1 _16951_ (.A(\top_ihp.oisc.regs[20][5] ),
    .X(_00863_));
 sg13g2_buf_1 _16952_ (.A(\top_ihp.oisc.regs[20][6] ),
    .X(_00864_));
 sg13g2_buf_1 _16953_ (.A(\top_ihp.oisc.regs[20][7] ),
    .X(_00865_));
 sg13g2_buf_1 _16954_ (.A(\top_ihp.oisc.regs[20][8] ),
    .X(_00866_));
 sg13g2_buf_1 _16955_ (.A(\top_ihp.oisc.regs[20][9] ),
    .X(_00867_));
 sg13g2_buf_1 _16956_ (.A(\top_ihp.oisc.regs[21][0] ),
    .X(_00868_));
 sg13g2_buf_1 _16957_ (.A(\top_ihp.oisc.regs[21][10] ),
    .X(_00869_));
 sg13g2_buf_1 _16958_ (.A(\top_ihp.oisc.regs[21][11] ),
    .X(_00870_));
 sg13g2_buf_1 _16959_ (.A(\top_ihp.oisc.regs[21][12] ),
    .X(_00871_));
 sg13g2_buf_1 _16960_ (.A(\top_ihp.oisc.regs[21][13] ),
    .X(_00872_));
 sg13g2_buf_1 _16961_ (.A(\top_ihp.oisc.regs[21][14] ),
    .X(_00873_));
 sg13g2_buf_1 _16962_ (.A(\top_ihp.oisc.regs[21][15] ),
    .X(_00874_));
 sg13g2_buf_1 _16963_ (.A(\top_ihp.oisc.regs[21][16] ),
    .X(_00875_));
 sg13g2_buf_1 _16964_ (.A(\top_ihp.oisc.regs[21][17] ),
    .X(_00876_));
 sg13g2_buf_1 _16965_ (.A(\top_ihp.oisc.regs[21][18] ),
    .X(_00877_));
 sg13g2_buf_1 _16966_ (.A(\top_ihp.oisc.regs[21][19] ),
    .X(_00878_));
 sg13g2_buf_1 _16967_ (.A(\top_ihp.oisc.regs[21][1] ),
    .X(_00879_));
 sg13g2_buf_1 _16968_ (.A(\top_ihp.oisc.regs[21][20] ),
    .X(_00880_));
 sg13g2_buf_1 _16969_ (.A(\top_ihp.oisc.regs[21][21] ),
    .X(_00881_));
 sg13g2_buf_1 _16970_ (.A(\top_ihp.oisc.regs[21][22] ),
    .X(_00882_));
 sg13g2_buf_1 _16971_ (.A(\top_ihp.oisc.regs[21][23] ),
    .X(_00883_));
 sg13g2_buf_1 _16972_ (.A(\top_ihp.oisc.regs[21][24] ),
    .X(_00884_));
 sg13g2_buf_1 _16973_ (.A(\top_ihp.oisc.regs[21][25] ),
    .X(_00885_));
 sg13g2_buf_1 _16974_ (.A(\top_ihp.oisc.regs[21][26] ),
    .X(_00886_));
 sg13g2_buf_1 _16975_ (.A(\top_ihp.oisc.regs[21][27] ),
    .X(_00887_));
 sg13g2_buf_1 _16976_ (.A(\top_ihp.oisc.regs[21][28] ),
    .X(_00888_));
 sg13g2_buf_1 _16977_ (.A(\top_ihp.oisc.regs[21][29] ),
    .X(_00889_));
 sg13g2_buf_1 _16978_ (.A(\top_ihp.oisc.regs[21][2] ),
    .X(_00890_));
 sg13g2_buf_1 _16979_ (.A(\top_ihp.oisc.regs[21][30] ),
    .X(_00891_));
 sg13g2_buf_1 _16980_ (.A(\top_ihp.oisc.regs[21][31] ),
    .X(_00892_));
 sg13g2_buf_1 _16981_ (.A(\top_ihp.oisc.regs[21][3] ),
    .X(_00893_));
 sg13g2_buf_1 _16982_ (.A(\top_ihp.oisc.regs[21][4] ),
    .X(_00894_));
 sg13g2_buf_1 _16983_ (.A(\top_ihp.oisc.regs[21][5] ),
    .X(_00895_));
 sg13g2_buf_1 _16984_ (.A(\top_ihp.oisc.regs[21][6] ),
    .X(_00896_));
 sg13g2_buf_1 _16985_ (.A(\top_ihp.oisc.regs[21][7] ),
    .X(_00897_));
 sg13g2_buf_1 _16986_ (.A(\top_ihp.oisc.regs[21][8] ),
    .X(_00898_));
 sg13g2_buf_1 _16987_ (.A(\top_ihp.oisc.regs[21][9] ),
    .X(_00899_));
 sg13g2_buf_1 _16988_ (.A(\top_ihp.oisc.regs[22][0] ),
    .X(_00900_));
 sg13g2_buf_1 _16989_ (.A(\top_ihp.oisc.regs[22][10] ),
    .X(_00901_));
 sg13g2_buf_1 _16990_ (.A(\top_ihp.oisc.regs[22][11] ),
    .X(_00902_));
 sg13g2_buf_1 _16991_ (.A(\top_ihp.oisc.regs[22][12] ),
    .X(_00903_));
 sg13g2_buf_1 _16992_ (.A(\top_ihp.oisc.regs[22][13] ),
    .X(_00904_));
 sg13g2_buf_1 _16993_ (.A(\top_ihp.oisc.regs[22][14] ),
    .X(_00905_));
 sg13g2_buf_1 _16994_ (.A(\top_ihp.oisc.regs[22][15] ),
    .X(_00906_));
 sg13g2_buf_1 _16995_ (.A(\top_ihp.oisc.regs[22][16] ),
    .X(_00907_));
 sg13g2_buf_1 _16996_ (.A(\top_ihp.oisc.regs[22][17] ),
    .X(_00908_));
 sg13g2_buf_1 _16997_ (.A(\top_ihp.oisc.regs[22][18] ),
    .X(_00909_));
 sg13g2_buf_1 _16998_ (.A(\top_ihp.oisc.regs[22][19] ),
    .X(_00910_));
 sg13g2_buf_1 _16999_ (.A(\top_ihp.oisc.regs[22][1] ),
    .X(_00911_));
 sg13g2_buf_1 _17000_ (.A(\top_ihp.oisc.regs[22][20] ),
    .X(_00912_));
 sg13g2_buf_1 _17001_ (.A(\top_ihp.oisc.regs[22][21] ),
    .X(_00913_));
 sg13g2_buf_1 _17002_ (.A(\top_ihp.oisc.regs[22][22] ),
    .X(_00914_));
 sg13g2_buf_1 _17003_ (.A(\top_ihp.oisc.regs[22][23] ),
    .X(_00915_));
 sg13g2_buf_1 _17004_ (.A(\top_ihp.oisc.regs[22][24] ),
    .X(_00916_));
 sg13g2_buf_1 _17005_ (.A(\top_ihp.oisc.regs[22][25] ),
    .X(_00917_));
 sg13g2_buf_1 _17006_ (.A(\top_ihp.oisc.regs[22][26] ),
    .X(_00918_));
 sg13g2_buf_1 _17007_ (.A(\top_ihp.oisc.regs[22][27] ),
    .X(_00919_));
 sg13g2_buf_1 _17008_ (.A(\top_ihp.oisc.regs[22][28] ),
    .X(_00920_));
 sg13g2_buf_1 _17009_ (.A(\top_ihp.oisc.regs[22][29] ),
    .X(_00921_));
 sg13g2_buf_1 _17010_ (.A(\top_ihp.oisc.regs[22][2] ),
    .X(_00922_));
 sg13g2_buf_1 _17011_ (.A(\top_ihp.oisc.regs[22][30] ),
    .X(_00923_));
 sg13g2_buf_1 _17012_ (.A(\top_ihp.oisc.regs[22][31] ),
    .X(_00924_));
 sg13g2_buf_1 _17013_ (.A(\top_ihp.oisc.regs[22][3] ),
    .X(_00925_));
 sg13g2_buf_1 _17014_ (.A(\top_ihp.oisc.regs[22][4] ),
    .X(_00926_));
 sg13g2_buf_1 _17015_ (.A(\top_ihp.oisc.regs[22][5] ),
    .X(_00927_));
 sg13g2_buf_1 _17016_ (.A(\top_ihp.oisc.regs[22][6] ),
    .X(_00928_));
 sg13g2_buf_1 _17017_ (.A(\top_ihp.oisc.regs[22][7] ),
    .X(_00929_));
 sg13g2_buf_1 _17018_ (.A(\top_ihp.oisc.regs[22][8] ),
    .X(_00930_));
 sg13g2_buf_1 _17019_ (.A(\top_ihp.oisc.regs[22][9] ),
    .X(_00931_));
 sg13g2_buf_1 _17020_ (.A(\top_ihp.oisc.regs[23][0] ),
    .X(_00932_));
 sg13g2_buf_1 _17021_ (.A(\top_ihp.oisc.regs[23][10] ),
    .X(_00933_));
 sg13g2_buf_1 _17022_ (.A(\top_ihp.oisc.regs[23][11] ),
    .X(_00934_));
 sg13g2_buf_1 _17023_ (.A(\top_ihp.oisc.regs[23][12] ),
    .X(_00935_));
 sg13g2_buf_1 _17024_ (.A(\top_ihp.oisc.regs[23][13] ),
    .X(_00936_));
 sg13g2_buf_1 _17025_ (.A(\top_ihp.oisc.regs[23][14] ),
    .X(_00937_));
 sg13g2_buf_1 _17026_ (.A(\top_ihp.oisc.regs[23][15] ),
    .X(_00938_));
 sg13g2_buf_1 _17027_ (.A(\top_ihp.oisc.regs[23][16] ),
    .X(_00939_));
 sg13g2_buf_1 _17028_ (.A(\top_ihp.oisc.regs[23][17] ),
    .X(_00940_));
 sg13g2_buf_1 _17029_ (.A(\top_ihp.oisc.regs[23][18] ),
    .X(_00941_));
 sg13g2_buf_1 _17030_ (.A(\top_ihp.oisc.regs[23][19] ),
    .X(_00942_));
 sg13g2_buf_1 _17031_ (.A(\top_ihp.oisc.regs[23][1] ),
    .X(_00943_));
 sg13g2_buf_1 _17032_ (.A(\top_ihp.oisc.regs[23][20] ),
    .X(_00944_));
 sg13g2_buf_1 _17033_ (.A(\top_ihp.oisc.regs[23][21] ),
    .X(_00945_));
 sg13g2_buf_1 _17034_ (.A(\top_ihp.oisc.regs[23][22] ),
    .X(_00946_));
 sg13g2_buf_1 _17035_ (.A(\top_ihp.oisc.regs[23][23] ),
    .X(_00947_));
 sg13g2_buf_1 _17036_ (.A(\top_ihp.oisc.regs[23][24] ),
    .X(_00948_));
 sg13g2_buf_1 _17037_ (.A(\top_ihp.oisc.regs[23][25] ),
    .X(_00949_));
 sg13g2_buf_1 _17038_ (.A(\top_ihp.oisc.regs[23][26] ),
    .X(_00950_));
 sg13g2_buf_1 _17039_ (.A(\top_ihp.oisc.regs[23][27] ),
    .X(_00951_));
 sg13g2_buf_1 _17040_ (.A(\top_ihp.oisc.regs[23][28] ),
    .X(_00952_));
 sg13g2_buf_1 _17041_ (.A(\top_ihp.oisc.regs[23][29] ),
    .X(_00953_));
 sg13g2_buf_1 _17042_ (.A(\top_ihp.oisc.regs[23][2] ),
    .X(_00954_));
 sg13g2_buf_1 _17043_ (.A(\top_ihp.oisc.regs[23][30] ),
    .X(_00955_));
 sg13g2_buf_1 _17044_ (.A(\top_ihp.oisc.regs[23][31] ),
    .X(_00956_));
 sg13g2_buf_1 _17045_ (.A(\top_ihp.oisc.regs[23][3] ),
    .X(_00957_));
 sg13g2_buf_1 _17046_ (.A(\top_ihp.oisc.regs[23][4] ),
    .X(_00958_));
 sg13g2_buf_1 _17047_ (.A(\top_ihp.oisc.regs[23][5] ),
    .X(_00959_));
 sg13g2_buf_1 _17048_ (.A(\top_ihp.oisc.regs[23][6] ),
    .X(_00960_));
 sg13g2_buf_1 _17049_ (.A(\top_ihp.oisc.regs[23][7] ),
    .X(_00961_));
 sg13g2_buf_1 _17050_ (.A(\top_ihp.oisc.regs[23][8] ),
    .X(_00962_));
 sg13g2_buf_1 _17051_ (.A(\top_ihp.oisc.regs[23][9] ),
    .X(_00963_));
 sg13g2_buf_1 _17052_ (.A(\top_ihp.oisc.regs[24][0] ),
    .X(_00964_));
 sg13g2_buf_1 _17053_ (.A(\top_ihp.oisc.regs[24][10] ),
    .X(_00965_));
 sg13g2_buf_1 _17054_ (.A(\top_ihp.oisc.regs[24][11] ),
    .X(_00966_));
 sg13g2_buf_1 _17055_ (.A(\top_ihp.oisc.regs[24][12] ),
    .X(_00967_));
 sg13g2_buf_1 _17056_ (.A(\top_ihp.oisc.regs[24][13] ),
    .X(_00968_));
 sg13g2_buf_1 _17057_ (.A(\top_ihp.oisc.regs[24][14] ),
    .X(_00969_));
 sg13g2_buf_1 _17058_ (.A(\top_ihp.oisc.regs[24][15] ),
    .X(_00970_));
 sg13g2_buf_1 _17059_ (.A(\top_ihp.oisc.regs[24][16] ),
    .X(_00971_));
 sg13g2_buf_1 _17060_ (.A(\top_ihp.oisc.regs[24][17] ),
    .X(_00972_));
 sg13g2_buf_1 _17061_ (.A(\top_ihp.oisc.regs[24][18] ),
    .X(_00973_));
 sg13g2_buf_1 _17062_ (.A(\top_ihp.oisc.regs[24][19] ),
    .X(_00974_));
 sg13g2_buf_1 _17063_ (.A(\top_ihp.oisc.regs[24][1] ),
    .X(_00975_));
 sg13g2_buf_1 _17064_ (.A(\top_ihp.oisc.regs[24][20] ),
    .X(_00976_));
 sg13g2_buf_1 _17065_ (.A(\top_ihp.oisc.regs[24][21] ),
    .X(_00977_));
 sg13g2_buf_1 _17066_ (.A(\top_ihp.oisc.regs[24][22] ),
    .X(_00978_));
 sg13g2_buf_1 _17067_ (.A(\top_ihp.oisc.regs[24][23] ),
    .X(_00979_));
 sg13g2_buf_1 _17068_ (.A(\top_ihp.oisc.regs[24][24] ),
    .X(_00980_));
 sg13g2_buf_1 _17069_ (.A(\top_ihp.oisc.regs[24][25] ),
    .X(_00981_));
 sg13g2_buf_1 _17070_ (.A(\top_ihp.oisc.regs[24][26] ),
    .X(_00982_));
 sg13g2_buf_1 _17071_ (.A(\top_ihp.oisc.regs[24][27] ),
    .X(_00983_));
 sg13g2_buf_1 _17072_ (.A(\top_ihp.oisc.regs[24][28] ),
    .X(_00984_));
 sg13g2_buf_1 _17073_ (.A(\top_ihp.oisc.regs[24][29] ),
    .X(_00985_));
 sg13g2_buf_1 _17074_ (.A(\top_ihp.oisc.regs[24][2] ),
    .X(_00986_));
 sg13g2_buf_1 _17075_ (.A(\top_ihp.oisc.regs[24][30] ),
    .X(_00987_));
 sg13g2_buf_1 _17076_ (.A(\top_ihp.oisc.regs[24][31] ),
    .X(_00988_));
 sg13g2_buf_1 _17077_ (.A(\top_ihp.oisc.regs[24][3] ),
    .X(_00989_));
 sg13g2_buf_1 _17078_ (.A(\top_ihp.oisc.regs[24][4] ),
    .X(_00990_));
 sg13g2_buf_1 _17079_ (.A(\top_ihp.oisc.regs[24][5] ),
    .X(_00991_));
 sg13g2_buf_1 _17080_ (.A(\top_ihp.oisc.regs[24][6] ),
    .X(_00992_));
 sg13g2_buf_1 _17081_ (.A(\top_ihp.oisc.regs[24][7] ),
    .X(_00993_));
 sg13g2_buf_1 _17082_ (.A(\top_ihp.oisc.regs[24][8] ),
    .X(_00994_));
 sg13g2_buf_1 _17083_ (.A(\top_ihp.oisc.regs[24][9] ),
    .X(_00995_));
 sg13g2_buf_1 _17084_ (.A(\top_ihp.oisc.regs[25][0] ),
    .X(_00996_));
 sg13g2_buf_1 _17085_ (.A(\top_ihp.oisc.regs[25][10] ),
    .X(_00997_));
 sg13g2_buf_1 _17086_ (.A(\top_ihp.oisc.regs[25][11] ),
    .X(_00998_));
 sg13g2_buf_1 _17087_ (.A(\top_ihp.oisc.regs[25][12] ),
    .X(_00999_));
 sg13g2_buf_1 _17088_ (.A(\top_ihp.oisc.regs[25][13] ),
    .X(_01000_));
 sg13g2_buf_1 _17089_ (.A(\top_ihp.oisc.regs[25][14] ),
    .X(_01001_));
 sg13g2_buf_1 _17090_ (.A(\top_ihp.oisc.regs[25][15] ),
    .X(_01002_));
 sg13g2_buf_1 _17091_ (.A(\top_ihp.oisc.regs[25][16] ),
    .X(_01003_));
 sg13g2_buf_1 _17092_ (.A(\top_ihp.oisc.regs[25][17] ),
    .X(_01004_));
 sg13g2_buf_1 _17093_ (.A(\top_ihp.oisc.regs[25][18] ),
    .X(_01005_));
 sg13g2_buf_1 _17094_ (.A(\top_ihp.oisc.regs[25][19] ),
    .X(_01006_));
 sg13g2_buf_1 _17095_ (.A(\top_ihp.oisc.regs[25][1] ),
    .X(_01007_));
 sg13g2_buf_1 _17096_ (.A(\top_ihp.oisc.regs[25][20] ),
    .X(_01008_));
 sg13g2_buf_1 _17097_ (.A(\top_ihp.oisc.regs[25][21] ),
    .X(_01009_));
 sg13g2_buf_1 _17098_ (.A(\top_ihp.oisc.regs[25][22] ),
    .X(_01010_));
 sg13g2_buf_1 _17099_ (.A(\top_ihp.oisc.regs[25][23] ),
    .X(_01011_));
 sg13g2_buf_1 _17100_ (.A(\top_ihp.oisc.regs[25][24] ),
    .X(_01012_));
 sg13g2_buf_1 _17101_ (.A(\top_ihp.oisc.regs[25][25] ),
    .X(_01013_));
 sg13g2_buf_1 _17102_ (.A(\top_ihp.oisc.regs[25][26] ),
    .X(_01014_));
 sg13g2_buf_1 _17103_ (.A(\top_ihp.oisc.regs[25][27] ),
    .X(_01015_));
 sg13g2_buf_1 _17104_ (.A(\top_ihp.oisc.regs[25][28] ),
    .X(_01016_));
 sg13g2_buf_1 _17105_ (.A(\top_ihp.oisc.regs[25][29] ),
    .X(_01017_));
 sg13g2_buf_1 _17106_ (.A(\top_ihp.oisc.regs[25][2] ),
    .X(_01018_));
 sg13g2_buf_1 _17107_ (.A(\top_ihp.oisc.regs[25][30] ),
    .X(_01019_));
 sg13g2_buf_1 _17108_ (.A(\top_ihp.oisc.regs[25][31] ),
    .X(_01020_));
 sg13g2_buf_1 _17109_ (.A(\top_ihp.oisc.regs[25][3] ),
    .X(_01021_));
 sg13g2_buf_1 _17110_ (.A(\top_ihp.oisc.regs[25][4] ),
    .X(_01022_));
 sg13g2_buf_1 _17111_ (.A(\top_ihp.oisc.regs[25][5] ),
    .X(_01023_));
 sg13g2_buf_1 _17112_ (.A(\top_ihp.oisc.regs[25][6] ),
    .X(_01024_));
 sg13g2_buf_1 _17113_ (.A(\top_ihp.oisc.regs[25][7] ),
    .X(_01025_));
 sg13g2_buf_1 _17114_ (.A(\top_ihp.oisc.regs[25][8] ),
    .X(_01026_));
 sg13g2_buf_1 _17115_ (.A(\top_ihp.oisc.regs[25][9] ),
    .X(_01027_));
 sg13g2_buf_1 _17116_ (.A(\top_ihp.oisc.regs[26][0] ),
    .X(_01028_));
 sg13g2_buf_1 _17117_ (.A(\top_ihp.oisc.regs[26][10] ),
    .X(_01029_));
 sg13g2_buf_1 _17118_ (.A(\top_ihp.oisc.regs[26][11] ),
    .X(_01030_));
 sg13g2_buf_1 _17119_ (.A(\top_ihp.oisc.regs[26][12] ),
    .X(_01031_));
 sg13g2_buf_1 _17120_ (.A(\top_ihp.oisc.regs[26][13] ),
    .X(_01032_));
 sg13g2_buf_1 _17121_ (.A(\top_ihp.oisc.regs[26][14] ),
    .X(_01033_));
 sg13g2_buf_1 _17122_ (.A(\top_ihp.oisc.regs[26][15] ),
    .X(_01034_));
 sg13g2_buf_1 _17123_ (.A(\top_ihp.oisc.regs[26][16] ),
    .X(_01035_));
 sg13g2_buf_1 _17124_ (.A(\top_ihp.oisc.regs[26][17] ),
    .X(_01036_));
 sg13g2_buf_1 _17125_ (.A(\top_ihp.oisc.regs[26][18] ),
    .X(_01037_));
 sg13g2_buf_1 _17126_ (.A(\top_ihp.oisc.regs[26][19] ),
    .X(_01038_));
 sg13g2_buf_1 _17127_ (.A(\top_ihp.oisc.regs[26][1] ),
    .X(_01039_));
 sg13g2_buf_1 _17128_ (.A(\top_ihp.oisc.regs[26][20] ),
    .X(_01040_));
 sg13g2_buf_1 _17129_ (.A(\top_ihp.oisc.regs[26][21] ),
    .X(_01041_));
 sg13g2_buf_1 _17130_ (.A(\top_ihp.oisc.regs[26][22] ),
    .X(_01042_));
 sg13g2_buf_1 _17131_ (.A(\top_ihp.oisc.regs[26][23] ),
    .X(_01043_));
 sg13g2_buf_1 _17132_ (.A(\top_ihp.oisc.regs[26][24] ),
    .X(_01044_));
 sg13g2_buf_1 _17133_ (.A(\top_ihp.oisc.regs[26][25] ),
    .X(_01045_));
 sg13g2_buf_1 _17134_ (.A(\top_ihp.oisc.regs[26][26] ),
    .X(_01046_));
 sg13g2_buf_1 _17135_ (.A(\top_ihp.oisc.regs[26][27] ),
    .X(_01047_));
 sg13g2_buf_1 _17136_ (.A(\top_ihp.oisc.regs[26][28] ),
    .X(_01048_));
 sg13g2_buf_1 _17137_ (.A(\top_ihp.oisc.regs[26][29] ),
    .X(_01049_));
 sg13g2_buf_1 _17138_ (.A(\top_ihp.oisc.regs[26][2] ),
    .X(_01050_));
 sg13g2_buf_1 _17139_ (.A(\top_ihp.oisc.regs[26][30] ),
    .X(_01051_));
 sg13g2_buf_1 _17140_ (.A(\top_ihp.oisc.regs[26][31] ),
    .X(_01052_));
 sg13g2_buf_1 _17141_ (.A(\top_ihp.oisc.regs[26][3] ),
    .X(_01053_));
 sg13g2_buf_1 _17142_ (.A(\top_ihp.oisc.regs[26][4] ),
    .X(_01054_));
 sg13g2_buf_1 _17143_ (.A(\top_ihp.oisc.regs[26][5] ),
    .X(_01055_));
 sg13g2_buf_1 _17144_ (.A(\top_ihp.oisc.regs[26][6] ),
    .X(_01056_));
 sg13g2_buf_1 _17145_ (.A(\top_ihp.oisc.regs[26][7] ),
    .X(_01057_));
 sg13g2_buf_1 _17146_ (.A(\top_ihp.oisc.regs[26][8] ),
    .X(_01058_));
 sg13g2_buf_1 _17147_ (.A(\top_ihp.oisc.regs[26][9] ),
    .X(_01059_));
 sg13g2_buf_1 _17148_ (.A(\top_ihp.oisc.regs[27][0] ),
    .X(_01060_));
 sg13g2_buf_1 _17149_ (.A(\top_ihp.oisc.regs[27][10] ),
    .X(_01061_));
 sg13g2_buf_1 _17150_ (.A(\top_ihp.oisc.regs[27][11] ),
    .X(_01062_));
 sg13g2_buf_1 _17151_ (.A(\top_ihp.oisc.regs[27][12] ),
    .X(_01063_));
 sg13g2_buf_1 _17152_ (.A(\top_ihp.oisc.regs[27][13] ),
    .X(_01064_));
 sg13g2_buf_1 _17153_ (.A(\top_ihp.oisc.regs[27][14] ),
    .X(_01065_));
 sg13g2_buf_1 _17154_ (.A(\top_ihp.oisc.regs[27][15] ),
    .X(_01066_));
 sg13g2_buf_1 _17155_ (.A(\top_ihp.oisc.regs[27][16] ),
    .X(_01067_));
 sg13g2_buf_1 _17156_ (.A(\top_ihp.oisc.regs[27][17] ),
    .X(_01068_));
 sg13g2_buf_1 _17157_ (.A(\top_ihp.oisc.regs[27][18] ),
    .X(_01069_));
 sg13g2_buf_1 _17158_ (.A(\top_ihp.oisc.regs[27][19] ),
    .X(_01070_));
 sg13g2_buf_1 _17159_ (.A(\top_ihp.oisc.regs[27][1] ),
    .X(_01071_));
 sg13g2_buf_1 _17160_ (.A(\top_ihp.oisc.regs[27][20] ),
    .X(_01072_));
 sg13g2_buf_1 _17161_ (.A(\top_ihp.oisc.regs[27][21] ),
    .X(_01073_));
 sg13g2_buf_1 _17162_ (.A(\top_ihp.oisc.regs[27][22] ),
    .X(_01074_));
 sg13g2_buf_1 _17163_ (.A(\top_ihp.oisc.regs[27][23] ),
    .X(_01075_));
 sg13g2_buf_1 _17164_ (.A(\top_ihp.oisc.regs[27][24] ),
    .X(_01076_));
 sg13g2_buf_1 _17165_ (.A(\top_ihp.oisc.regs[27][25] ),
    .X(_01077_));
 sg13g2_buf_1 _17166_ (.A(\top_ihp.oisc.regs[27][26] ),
    .X(_01078_));
 sg13g2_buf_1 _17167_ (.A(\top_ihp.oisc.regs[27][27] ),
    .X(_01079_));
 sg13g2_buf_1 _17168_ (.A(\top_ihp.oisc.regs[27][28] ),
    .X(_01080_));
 sg13g2_buf_1 _17169_ (.A(\top_ihp.oisc.regs[27][29] ),
    .X(_01081_));
 sg13g2_buf_1 _17170_ (.A(\top_ihp.oisc.regs[27][2] ),
    .X(_01082_));
 sg13g2_buf_1 _17171_ (.A(\top_ihp.oisc.regs[27][30] ),
    .X(_01083_));
 sg13g2_buf_1 _17172_ (.A(\top_ihp.oisc.regs[27][31] ),
    .X(_01084_));
 sg13g2_buf_1 _17173_ (.A(\top_ihp.oisc.regs[27][3] ),
    .X(_01085_));
 sg13g2_buf_1 _17174_ (.A(\top_ihp.oisc.regs[27][4] ),
    .X(_01086_));
 sg13g2_buf_1 _17175_ (.A(\top_ihp.oisc.regs[27][5] ),
    .X(_01087_));
 sg13g2_buf_1 _17176_ (.A(\top_ihp.oisc.regs[27][6] ),
    .X(_01088_));
 sg13g2_buf_1 _17177_ (.A(\top_ihp.oisc.regs[27][7] ),
    .X(_01089_));
 sg13g2_buf_1 _17178_ (.A(\top_ihp.oisc.regs[27][8] ),
    .X(_01090_));
 sg13g2_buf_1 _17179_ (.A(\top_ihp.oisc.regs[27][9] ),
    .X(_01091_));
 sg13g2_buf_1 _17180_ (.A(\top_ihp.oisc.regs[28][0] ),
    .X(_01092_));
 sg13g2_buf_1 _17181_ (.A(\top_ihp.oisc.regs[28][10] ),
    .X(_01093_));
 sg13g2_buf_1 _17182_ (.A(\top_ihp.oisc.regs[28][11] ),
    .X(_01094_));
 sg13g2_buf_1 _17183_ (.A(\top_ihp.oisc.regs[28][12] ),
    .X(_01095_));
 sg13g2_buf_1 _17184_ (.A(\top_ihp.oisc.regs[28][13] ),
    .X(_01096_));
 sg13g2_buf_1 _17185_ (.A(\top_ihp.oisc.regs[28][14] ),
    .X(_01097_));
 sg13g2_buf_1 _17186_ (.A(\top_ihp.oisc.regs[28][15] ),
    .X(_01098_));
 sg13g2_buf_1 _17187_ (.A(\top_ihp.oisc.regs[28][16] ),
    .X(_01099_));
 sg13g2_buf_1 _17188_ (.A(\top_ihp.oisc.regs[28][17] ),
    .X(_01100_));
 sg13g2_buf_1 _17189_ (.A(\top_ihp.oisc.regs[28][18] ),
    .X(_01101_));
 sg13g2_buf_1 _17190_ (.A(\top_ihp.oisc.regs[28][19] ),
    .X(_01102_));
 sg13g2_buf_1 _17191_ (.A(\top_ihp.oisc.regs[28][1] ),
    .X(_01103_));
 sg13g2_buf_1 _17192_ (.A(\top_ihp.oisc.regs[28][20] ),
    .X(_01104_));
 sg13g2_buf_1 _17193_ (.A(\top_ihp.oisc.regs[28][21] ),
    .X(_01105_));
 sg13g2_buf_1 _17194_ (.A(\top_ihp.oisc.regs[28][22] ),
    .X(_01106_));
 sg13g2_buf_1 _17195_ (.A(\top_ihp.oisc.regs[28][23] ),
    .X(_01107_));
 sg13g2_buf_1 _17196_ (.A(\top_ihp.oisc.regs[28][24] ),
    .X(_01108_));
 sg13g2_buf_1 _17197_ (.A(\top_ihp.oisc.regs[28][25] ),
    .X(_01109_));
 sg13g2_buf_1 _17198_ (.A(\top_ihp.oisc.regs[28][26] ),
    .X(_01110_));
 sg13g2_buf_1 _17199_ (.A(\top_ihp.oisc.regs[28][27] ),
    .X(_01111_));
 sg13g2_buf_1 _17200_ (.A(\top_ihp.oisc.regs[28][28] ),
    .X(_01112_));
 sg13g2_buf_1 _17201_ (.A(\top_ihp.oisc.regs[28][29] ),
    .X(_01113_));
 sg13g2_buf_1 _17202_ (.A(\top_ihp.oisc.regs[28][2] ),
    .X(_01114_));
 sg13g2_buf_1 _17203_ (.A(\top_ihp.oisc.regs[28][30] ),
    .X(_01115_));
 sg13g2_buf_1 _17204_ (.A(\top_ihp.oisc.regs[28][31] ),
    .X(_01116_));
 sg13g2_buf_1 _17205_ (.A(\top_ihp.oisc.regs[28][3] ),
    .X(_01117_));
 sg13g2_buf_1 _17206_ (.A(\top_ihp.oisc.regs[28][4] ),
    .X(_01118_));
 sg13g2_buf_1 _17207_ (.A(\top_ihp.oisc.regs[28][5] ),
    .X(_01119_));
 sg13g2_buf_1 _17208_ (.A(\top_ihp.oisc.regs[28][6] ),
    .X(_01120_));
 sg13g2_buf_1 _17209_ (.A(\top_ihp.oisc.regs[28][7] ),
    .X(_01121_));
 sg13g2_buf_1 _17210_ (.A(\top_ihp.oisc.regs[28][8] ),
    .X(_01122_));
 sg13g2_buf_1 _17211_ (.A(\top_ihp.oisc.regs[28][9] ),
    .X(_01123_));
 sg13g2_buf_1 _17212_ (.A(\top_ihp.oisc.regs[29][0] ),
    .X(_01124_));
 sg13g2_buf_1 _17213_ (.A(\top_ihp.oisc.regs[29][10] ),
    .X(_01125_));
 sg13g2_buf_1 _17214_ (.A(\top_ihp.oisc.regs[29][11] ),
    .X(_01126_));
 sg13g2_buf_1 _17215_ (.A(\top_ihp.oisc.regs[29][12] ),
    .X(_01127_));
 sg13g2_buf_1 _17216_ (.A(\top_ihp.oisc.regs[29][13] ),
    .X(_01128_));
 sg13g2_buf_1 _17217_ (.A(\top_ihp.oisc.regs[29][14] ),
    .X(_01129_));
 sg13g2_buf_1 _17218_ (.A(\top_ihp.oisc.regs[29][15] ),
    .X(_01130_));
 sg13g2_buf_1 _17219_ (.A(\top_ihp.oisc.regs[29][16] ),
    .X(_01131_));
 sg13g2_buf_1 _17220_ (.A(\top_ihp.oisc.regs[29][17] ),
    .X(_01132_));
 sg13g2_buf_1 _17221_ (.A(\top_ihp.oisc.regs[29][18] ),
    .X(_01133_));
 sg13g2_buf_1 _17222_ (.A(\top_ihp.oisc.regs[29][19] ),
    .X(_01134_));
 sg13g2_buf_1 _17223_ (.A(\top_ihp.oisc.regs[29][1] ),
    .X(_01135_));
 sg13g2_buf_1 _17224_ (.A(\top_ihp.oisc.regs[29][20] ),
    .X(_01136_));
 sg13g2_buf_1 _17225_ (.A(\top_ihp.oisc.regs[29][21] ),
    .X(_01137_));
 sg13g2_buf_1 _17226_ (.A(\top_ihp.oisc.regs[29][22] ),
    .X(_01138_));
 sg13g2_buf_1 _17227_ (.A(\top_ihp.oisc.regs[29][23] ),
    .X(_01139_));
 sg13g2_buf_1 _17228_ (.A(\top_ihp.oisc.regs[29][24] ),
    .X(_01140_));
 sg13g2_buf_1 _17229_ (.A(\top_ihp.oisc.regs[29][25] ),
    .X(_01141_));
 sg13g2_buf_1 _17230_ (.A(\top_ihp.oisc.regs[29][26] ),
    .X(_01142_));
 sg13g2_buf_1 _17231_ (.A(\top_ihp.oisc.regs[29][27] ),
    .X(_01143_));
 sg13g2_buf_1 _17232_ (.A(\top_ihp.oisc.regs[29][28] ),
    .X(_01144_));
 sg13g2_buf_1 _17233_ (.A(\top_ihp.oisc.regs[29][29] ),
    .X(_01145_));
 sg13g2_buf_1 _17234_ (.A(\top_ihp.oisc.regs[29][2] ),
    .X(_01146_));
 sg13g2_buf_1 _17235_ (.A(\top_ihp.oisc.regs[29][30] ),
    .X(_01147_));
 sg13g2_buf_1 _17236_ (.A(\top_ihp.oisc.regs[29][31] ),
    .X(_01148_));
 sg13g2_buf_1 _17237_ (.A(\top_ihp.oisc.regs[29][3] ),
    .X(_01149_));
 sg13g2_buf_1 _17238_ (.A(\top_ihp.oisc.regs[29][4] ),
    .X(_01150_));
 sg13g2_buf_1 _17239_ (.A(\top_ihp.oisc.regs[29][5] ),
    .X(_01151_));
 sg13g2_buf_1 _17240_ (.A(\top_ihp.oisc.regs[29][6] ),
    .X(_01152_));
 sg13g2_buf_1 _17241_ (.A(\top_ihp.oisc.regs[29][7] ),
    .X(_01153_));
 sg13g2_buf_1 _17242_ (.A(\top_ihp.oisc.regs[29][8] ),
    .X(_01154_));
 sg13g2_buf_1 _17243_ (.A(\top_ihp.oisc.regs[29][9] ),
    .X(_01155_));
 sg13g2_nand2_1 _17244_ (.Y(_10782_),
    .A(net767),
    .B(_10524_));
 sg13g2_buf_1 _17245_ (.A(_10782_),
    .X(_10783_));
 sg13g2_buf_1 _17246_ (.A(net643),
    .X(_10784_));
 sg13g2_buf_1 _17247_ (.A(_10782_),
    .X(_10785_));
 sg13g2_nand2_1 _17248_ (.Y(_10786_),
    .A(\top_ihp.oisc.regs[2][0] ),
    .B(net642));
 sg13g2_o21ai_1 _17249_ (.B1(_10786_),
    .Y(_01156_),
    .A1(net53),
    .A2(net508));
 sg13g2_nand2_1 _17250_ (.Y(_10787_),
    .A(\top_ihp.oisc.regs[2][10] ),
    .B(net642));
 sg13g2_o21ai_1 _17251_ (.B1(_10787_),
    .Y(_01157_),
    .A1(net155),
    .A2(net508));
 sg13g2_nand2_1 _17252_ (.Y(_10788_),
    .A(\top_ihp.oisc.regs[2][11] ),
    .B(net642));
 sg13g2_o21ai_1 _17253_ (.B1(_10788_),
    .Y(_01158_),
    .A1(net154),
    .A2(net508));
 sg13g2_nand2_1 _17254_ (.Y(_10789_),
    .A(\top_ihp.oisc.regs[2][12] ),
    .B(net642));
 sg13g2_o21ai_1 _17255_ (.B1(_10789_),
    .Y(_01159_),
    .A1(net137),
    .A2(_10784_));
 sg13g2_nand2_1 _17256_ (.Y(_10790_),
    .A(\top_ihp.oisc.regs[2][13] ),
    .B(net642));
 sg13g2_o21ai_1 _17257_ (.B1(_10790_),
    .Y(_01160_),
    .A1(net331),
    .A2(net508));
 sg13g2_nand2_1 _17258_ (.Y(_10791_),
    .A(\top_ihp.oisc.regs[2][14] ),
    .B(net642));
 sg13g2_o21ai_1 _17259_ (.B1(_10791_),
    .Y(_01161_),
    .A1(net136),
    .A2(net508));
 sg13g2_nand2_1 _17260_ (.Y(_10792_),
    .A(\top_ihp.oisc.regs[2][15] ),
    .B(net642));
 sg13g2_o21ai_1 _17261_ (.B1(_10792_),
    .Y(_01162_),
    .A1(net135),
    .A2(_10784_));
 sg13g2_nand2_1 _17262_ (.Y(_10793_),
    .A(\top_ihp.oisc.regs[2][16] ),
    .B(net642));
 sg13g2_o21ai_1 _17263_ (.B1(_10793_),
    .Y(_01163_),
    .A1(net150),
    .A2(net508));
 sg13g2_buf_1 _17264_ (.A(net643),
    .X(_10794_));
 sg13g2_nand2_1 _17265_ (.Y(_10795_),
    .A(\top_ihp.oisc.regs[2][17] ),
    .B(net507));
 sg13g2_o21ai_1 _17266_ (.B1(_10795_),
    .Y(_01164_),
    .A1(net328),
    .A2(net508));
 sg13g2_nand2_1 _17267_ (.Y(_10796_),
    .A(\top_ihp.oisc.regs[2][18] ),
    .B(net507));
 sg13g2_o21ai_1 _17268_ (.B1(_10796_),
    .Y(_01165_),
    .A1(net327),
    .A2(net508));
 sg13g2_buf_1 _17269_ (.A(net643),
    .X(_10797_));
 sg13g2_nand2_1 _17270_ (.Y(_10798_),
    .A(\top_ihp.oisc.regs[2][19] ),
    .B(net507));
 sg13g2_o21ai_1 _17271_ (.B1(_10798_),
    .Y(_01166_),
    .A1(net326),
    .A2(net506));
 sg13g2_nand2_1 _17272_ (.Y(_10799_),
    .A(\top_ihp.oisc.regs[2][1] ),
    .B(net507));
 sg13g2_o21ai_1 _17273_ (.B1(_10799_),
    .Y(_01167_),
    .A1(net134),
    .A2(net506));
 sg13g2_nand2_1 _17274_ (.Y(_10800_),
    .A(\top_ihp.oisc.regs[2][20] ),
    .B(_10794_));
 sg13g2_o21ai_1 _17275_ (.B1(_10800_),
    .Y(_01168_),
    .A1(net324),
    .A2(_10797_));
 sg13g2_nand2_1 _17276_ (.Y(_10801_),
    .A(\top_ihp.oisc.regs[2][21] ),
    .B(net507));
 sg13g2_o21ai_1 _17277_ (.B1(_10801_),
    .Y(_01169_),
    .A1(net323),
    .A2(net506));
 sg13g2_nand2_1 _17278_ (.Y(_10802_),
    .A(\top_ihp.oisc.regs[2][22] ),
    .B(_10794_));
 sg13g2_o21ai_1 _17279_ (.B1(_10802_),
    .Y(_01170_),
    .A1(net133),
    .A2(net506));
 sg13g2_nand2_1 _17280_ (.Y(_10803_),
    .A(\top_ihp.oisc.regs[2][23] ),
    .B(net507));
 sg13g2_o21ai_1 _17281_ (.B1(_10803_),
    .Y(_01171_),
    .A1(net321),
    .A2(net506));
 sg13g2_nand2_1 _17282_ (.Y(_10804_),
    .A(\top_ihp.oisc.regs[2][24] ),
    .B(net507));
 sg13g2_o21ai_1 _17283_ (.B1(_10804_),
    .Y(_01172_),
    .A1(net320),
    .A2(_10797_));
 sg13g2_nand2_1 _17284_ (.Y(_10805_),
    .A(\top_ihp.oisc.regs[2][25] ),
    .B(net507));
 sg13g2_o21ai_1 _17285_ (.B1(_10805_),
    .Y(_01173_),
    .A1(net132),
    .A2(net506));
 sg13g2_buf_8 _17286_ (.A(net643),
    .X(_10806_));
 sg13g2_nand2_1 _17287_ (.Y(_10807_),
    .A(\top_ihp.oisc.regs[2][26] ),
    .B(net505));
 sg13g2_o21ai_1 _17288_ (.B1(_10807_),
    .Y(_01174_),
    .A1(net146),
    .A2(net506));
 sg13g2_nand2_1 _17289_ (.Y(_10808_),
    .A(\top_ihp.oisc.regs[2][27] ),
    .B(net505));
 sg13g2_o21ai_1 _17290_ (.B1(_10808_),
    .Y(_01175_),
    .A1(net318),
    .A2(net506));
 sg13g2_buf_8 _17291_ (.A(net643),
    .X(_10809_));
 sg13g2_nand2_1 _17292_ (.Y(_10810_),
    .A(\top_ihp.oisc.regs[2][28] ),
    .B(net505));
 sg13g2_o21ai_1 _17293_ (.B1(_10810_),
    .Y(_01176_),
    .A1(net525),
    .A2(net504));
 sg13g2_nand2_1 _17294_ (.Y(_10811_),
    .A(\top_ihp.oisc.regs[2][29] ),
    .B(net505));
 sg13g2_o21ai_1 _17295_ (.B1(_10811_),
    .Y(_01177_),
    .A1(net317),
    .A2(net504));
 sg13g2_nand2_1 _17296_ (.Y(_10812_),
    .A(\top_ihp.oisc.regs[2][2] ),
    .B(_10806_));
 sg13g2_o21ai_1 _17297_ (.B1(_10812_),
    .Y(_01178_),
    .A1(net145),
    .A2(_10809_));
 sg13g2_nand2_1 _17298_ (.Y(_10813_),
    .A(\top_ihp.oisc.regs[2][30] ),
    .B(net505));
 sg13g2_o21ai_1 _17299_ (.B1(_10813_),
    .Y(_01179_),
    .A1(net144),
    .A2(net504));
 sg13g2_nand2_1 _17300_ (.Y(_10814_),
    .A(\top_ihp.oisc.regs[2][31] ),
    .B(net505));
 sg13g2_o21ai_1 _17301_ (.B1(_10814_),
    .Y(_01180_),
    .A1(net52),
    .A2(net504));
 sg13g2_nand2_1 _17302_ (.Y(_10815_),
    .A(\top_ihp.oisc.regs[2][3] ),
    .B(net505));
 sg13g2_o21ai_1 _17303_ (.B1(_10815_),
    .Y(_01181_),
    .A1(net143),
    .A2(net504));
 sg13g2_nand2_1 _17304_ (.Y(_10816_),
    .A(\top_ihp.oisc.regs[2][4] ),
    .B(net505));
 sg13g2_o21ai_1 _17305_ (.B1(_10816_),
    .Y(_01182_),
    .A1(net142),
    .A2(net504));
 sg13g2_nand2_1 _17306_ (.Y(_10817_),
    .A(\top_ihp.oisc.regs[2][5] ),
    .B(_10806_));
 sg13g2_o21ai_1 _17307_ (.B1(_10817_),
    .Y(_01183_),
    .A1(net141),
    .A2(net504));
 sg13g2_nand2_1 _17308_ (.Y(_10818_),
    .A(\top_ihp.oisc.regs[2][6] ),
    .B(net643));
 sg13g2_o21ai_1 _17309_ (.B1(_10818_),
    .Y(_01184_),
    .A1(net140),
    .A2(net504));
 sg13g2_nand2_1 _17310_ (.Y(_10819_),
    .A(\top_ihp.oisc.regs[2][7] ),
    .B(net643));
 sg13g2_o21ai_1 _17311_ (.B1(_10819_),
    .Y(_01185_),
    .A1(net139),
    .A2(_10809_));
 sg13g2_nand2_1 _17312_ (.Y(_10820_),
    .A(\top_ihp.oisc.regs[2][8] ),
    .B(_10783_));
 sg13g2_o21ai_1 _17313_ (.B1(_10820_),
    .Y(_01186_),
    .A1(net316),
    .A2(_10785_));
 sg13g2_nand2_1 _17314_ (.Y(_10821_),
    .A(\top_ihp.oisc.regs[2][9] ),
    .B(net643));
 sg13g2_o21ai_1 _17315_ (.B1(_10821_),
    .Y(_01187_),
    .A1(net138),
    .A2(_10785_));
 sg13g2_buf_1 _17316_ (.A(\top_ihp.oisc.regs[30][0] ),
    .X(_01188_));
 sg13g2_buf_1 _17317_ (.A(\top_ihp.oisc.regs[30][10] ),
    .X(_01189_));
 sg13g2_buf_1 _17318_ (.A(\top_ihp.oisc.regs[30][11] ),
    .X(_01190_));
 sg13g2_buf_1 _17319_ (.A(\top_ihp.oisc.regs[30][12] ),
    .X(_01191_));
 sg13g2_buf_1 _17320_ (.A(\top_ihp.oisc.regs[30][13] ),
    .X(_01192_));
 sg13g2_buf_1 _17321_ (.A(\top_ihp.oisc.regs[30][14] ),
    .X(_01193_));
 sg13g2_buf_1 _17322_ (.A(\top_ihp.oisc.regs[30][15] ),
    .X(_01194_));
 sg13g2_buf_1 _17323_ (.A(\top_ihp.oisc.regs[30][16] ),
    .X(_01195_));
 sg13g2_buf_1 _17324_ (.A(\top_ihp.oisc.regs[30][17] ),
    .X(_01196_));
 sg13g2_buf_1 _17325_ (.A(\top_ihp.oisc.regs[30][18] ),
    .X(_01197_));
 sg13g2_buf_1 _17326_ (.A(\top_ihp.oisc.regs[30][19] ),
    .X(_01198_));
 sg13g2_buf_1 _17327_ (.A(\top_ihp.oisc.regs[30][1] ),
    .X(_01199_));
 sg13g2_buf_1 _17328_ (.A(\top_ihp.oisc.regs[30][20] ),
    .X(_01200_));
 sg13g2_buf_1 _17329_ (.A(\top_ihp.oisc.regs[30][21] ),
    .X(_01201_));
 sg13g2_buf_1 _17330_ (.A(\top_ihp.oisc.regs[30][22] ),
    .X(_01202_));
 sg13g2_buf_1 _17331_ (.A(\top_ihp.oisc.regs[30][23] ),
    .X(_01203_));
 sg13g2_buf_1 _17332_ (.A(\top_ihp.oisc.regs[30][24] ),
    .X(_01204_));
 sg13g2_buf_1 _17333_ (.A(\top_ihp.oisc.regs[30][25] ),
    .X(_01205_));
 sg13g2_buf_1 _17334_ (.A(\top_ihp.oisc.regs[30][26] ),
    .X(_01206_));
 sg13g2_buf_1 _17335_ (.A(\top_ihp.oisc.regs[30][27] ),
    .X(_01207_));
 sg13g2_buf_1 _17336_ (.A(\top_ihp.oisc.regs[30][28] ),
    .X(_01208_));
 sg13g2_buf_1 _17337_ (.A(\top_ihp.oisc.regs[30][29] ),
    .X(_01209_));
 sg13g2_buf_1 _17338_ (.A(\top_ihp.oisc.regs[30][2] ),
    .X(_01210_));
 sg13g2_buf_1 _17339_ (.A(\top_ihp.oisc.regs[30][30] ),
    .X(_01211_));
 sg13g2_buf_1 _17340_ (.A(\top_ihp.oisc.regs[30][31] ),
    .X(_01212_));
 sg13g2_buf_1 _17341_ (.A(\top_ihp.oisc.regs[30][3] ),
    .X(_01213_));
 sg13g2_buf_1 _17342_ (.A(\top_ihp.oisc.regs[30][4] ),
    .X(_01214_));
 sg13g2_buf_1 _17343_ (.A(\top_ihp.oisc.regs[30][5] ),
    .X(_01215_));
 sg13g2_buf_1 _17344_ (.A(\top_ihp.oisc.regs[30][6] ),
    .X(_01216_));
 sg13g2_buf_1 _17345_ (.A(\top_ihp.oisc.regs[30][7] ),
    .X(_01217_));
 sg13g2_buf_1 _17346_ (.A(\top_ihp.oisc.regs[30][8] ),
    .X(_01218_));
 sg13g2_buf_1 _17347_ (.A(\top_ihp.oisc.regs[30][9] ),
    .X(_01219_));
 sg13g2_buf_1 _17348_ (.A(\top_ihp.oisc.regs[31][0] ),
    .X(_01220_));
 sg13g2_buf_1 _17349_ (.A(\top_ihp.oisc.regs[31][10] ),
    .X(_01221_));
 sg13g2_buf_1 _17350_ (.A(\top_ihp.oisc.regs[31][11] ),
    .X(_01222_));
 sg13g2_buf_1 _17351_ (.A(\top_ihp.oisc.regs[31][12] ),
    .X(_01223_));
 sg13g2_buf_1 _17352_ (.A(\top_ihp.oisc.regs[31][13] ),
    .X(_01224_));
 sg13g2_buf_1 _17353_ (.A(\top_ihp.oisc.regs[31][14] ),
    .X(_01225_));
 sg13g2_buf_1 _17354_ (.A(\top_ihp.oisc.regs[31][15] ),
    .X(_01226_));
 sg13g2_buf_1 _17355_ (.A(\top_ihp.oisc.regs[31][16] ),
    .X(_01227_));
 sg13g2_buf_1 _17356_ (.A(\top_ihp.oisc.regs[31][17] ),
    .X(_01228_));
 sg13g2_buf_1 _17357_ (.A(\top_ihp.oisc.regs[31][18] ),
    .X(_01229_));
 sg13g2_buf_1 _17358_ (.A(\top_ihp.oisc.regs[31][19] ),
    .X(_01230_));
 sg13g2_buf_1 _17359_ (.A(\top_ihp.oisc.regs[31][1] ),
    .X(_01231_));
 sg13g2_buf_1 _17360_ (.A(\top_ihp.oisc.regs[31][20] ),
    .X(_01232_));
 sg13g2_buf_1 _17361_ (.A(\top_ihp.oisc.regs[31][21] ),
    .X(_01233_));
 sg13g2_buf_1 _17362_ (.A(\top_ihp.oisc.regs[31][22] ),
    .X(_01234_));
 sg13g2_buf_1 _17363_ (.A(\top_ihp.oisc.regs[31][23] ),
    .X(_01235_));
 sg13g2_buf_1 _17364_ (.A(\top_ihp.oisc.regs[31][24] ),
    .X(_01236_));
 sg13g2_buf_1 _17365_ (.A(\top_ihp.oisc.regs[31][25] ),
    .X(_01237_));
 sg13g2_buf_1 _17366_ (.A(\top_ihp.oisc.regs[31][26] ),
    .X(_01238_));
 sg13g2_buf_1 _17367_ (.A(\top_ihp.oisc.regs[31][27] ),
    .X(_01239_));
 sg13g2_buf_1 _17368_ (.A(\top_ihp.oisc.regs[31][28] ),
    .X(_01240_));
 sg13g2_buf_1 _17369_ (.A(\top_ihp.oisc.regs[31][29] ),
    .X(_01241_));
 sg13g2_buf_1 _17370_ (.A(\top_ihp.oisc.regs[31][2] ),
    .X(_01242_));
 sg13g2_buf_1 _17371_ (.A(\top_ihp.oisc.regs[31][30] ),
    .X(_01243_));
 sg13g2_buf_1 _17372_ (.A(\top_ihp.oisc.regs[31][31] ),
    .X(_01244_));
 sg13g2_buf_1 _17373_ (.A(\top_ihp.oisc.regs[31][3] ),
    .X(_01245_));
 sg13g2_buf_1 _17374_ (.A(\top_ihp.oisc.regs[31][4] ),
    .X(_01246_));
 sg13g2_buf_1 _17375_ (.A(\top_ihp.oisc.regs[31][5] ),
    .X(_01247_));
 sg13g2_buf_1 _17376_ (.A(\top_ihp.oisc.regs[31][6] ),
    .X(_01248_));
 sg13g2_buf_1 _17377_ (.A(\top_ihp.oisc.regs[31][7] ),
    .X(_01249_));
 sg13g2_buf_1 _17378_ (.A(\top_ihp.oisc.regs[31][8] ),
    .X(_01250_));
 sg13g2_buf_1 _17379_ (.A(\top_ihp.oisc.regs[31][9] ),
    .X(_01251_));
 sg13g2_buf_1 _17380_ (.A(\top_ihp.oisc.regs[32][0] ),
    .X(_01252_));
 sg13g2_buf_1 _17381_ (.A(\top_ihp.oisc.regs[32][10] ),
    .X(_01253_));
 sg13g2_buf_1 _17382_ (.A(\top_ihp.oisc.regs[32][11] ),
    .X(_01254_));
 sg13g2_buf_1 _17383_ (.A(\top_ihp.oisc.regs[32][12] ),
    .X(_01255_));
 sg13g2_buf_1 _17384_ (.A(\top_ihp.oisc.regs[32][13] ),
    .X(_01256_));
 sg13g2_buf_1 _17385_ (.A(\top_ihp.oisc.regs[32][14] ),
    .X(_01257_));
 sg13g2_buf_1 _17386_ (.A(\top_ihp.oisc.regs[32][15] ),
    .X(_01258_));
 sg13g2_buf_1 _17387_ (.A(\top_ihp.oisc.regs[32][16] ),
    .X(_01259_));
 sg13g2_buf_1 _17388_ (.A(\top_ihp.oisc.regs[32][17] ),
    .X(_01260_));
 sg13g2_buf_1 _17389_ (.A(\top_ihp.oisc.regs[32][18] ),
    .X(_01261_));
 sg13g2_buf_1 _17390_ (.A(\top_ihp.oisc.regs[32][19] ),
    .X(_01262_));
 sg13g2_buf_1 _17391_ (.A(\top_ihp.oisc.regs[32][1] ),
    .X(_01263_));
 sg13g2_buf_1 _17392_ (.A(\top_ihp.oisc.regs[32][20] ),
    .X(_01264_));
 sg13g2_buf_1 _17393_ (.A(\top_ihp.oisc.regs[32][21] ),
    .X(_01265_));
 sg13g2_buf_1 _17394_ (.A(\top_ihp.oisc.regs[32][22] ),
    .X(_01266_));
 sg13g2_buf_1 _17395_ (.A(\top_ihp.oisc.regs[32][23] ),
    .X(_01267_));
 sg13g2_buf_1 _17396_ (.A(\top_ihp.oisc.regs[32][24] ),
    .X(_01268_));
 sg13g2_buf_1 _17397_ (.A(\top_ihp.oisc.regs[32][25] ),
    .X(_01269_));
 sg13g2_buf_1 _17398_ (.A(\top_ihp.oisc.regs[32][26] ),
    .X(_01270_));
 sg13g2_buf_1 _17399_ (.A(\top_ihp.oisc.regs[32][27] ),
    .X(_01271_));
 sg13g2_buf_1 _17400_ (.A(\top_ihp.oisc.regs[32][28] ),
    .X(_01272_));
 sg13g2_buf_1 _17401_ (.A(\top_ihp.oisc.regs[32][29] ),
    .X(_01273_));
 sg13g2_buf_1 _17402_ (.A(\top_ihp.oisc.regs[32][2] ),
    .X(_01274_));
 sg13g2_buf_1 _17403_ (.A(\top_ihp.oisc.regs[32][30] ),
    .X(_01275_));
 sg13g2_buf_1 _17404_ (.A(\top_ihp.oisc.regs[32][31] ),
    .X(_01276_));
 sg13g2_buf_1 _17405_ (.A(\top_ihp.oisc.regs[32][3] ),
    .X(_01277_));
 sg13g2_buf_1 _17406_ (.A(\top_ihp.oisc.regs[32][4] ),
    .X(_01278_));
 sg13g2_buf_1 _17407_ (.A(\top_ihp.oisc.regs[32][5] ),
    .X(_01279_));
 sg13g2_buf_1 _17408_ (.A(\top_ihp.oisc.regs[32][6] ),
    .X(_01280_));
 sg13g2_buf_1 _17409_ (.A(\top_ihp.oisc.regs[32][7] ),
    .X(_01281_));
 sg13g2_buf_1 _17410_ (.A(\top_ihp.oisc.regs[32][8] ),
    .X(_01282_));
 sg13g2_buf_1 _17411_ (.A(\top_ihp.oisc.regs[32][9] ),
    .X(_01283_));
 sg13g2_buf_1 _17412_ (.A(_10649_),
    .X(_10822_));
 sg13g2_nand2b_2 _17413_ (.Y(_10823_),
    .B(_09738_),
    .A_N(_09729_));
 sg13g2_a21oi_1 _17414_ (.A1(_09725_),
    .A2(net766),
    .Y(_10824_),
    .B1(_10823_));
 sg13g2_buf_2 _17415_ (.A(_10824_),
    .X(_10825_));
 sg13g2_buf_8 _17416_ (.A(_10825_),
    .X(_10826_));
 sg13g2_nand3_1 _17417_ (.B(net784),
    .C(net708),
    .A(_09725_),
    .Y(_10827_));
 sg13g2_buf_1 _17418_ (.A(_10827_),
    .X(_10828_));
 sg13g2_buf_1 _17419_ (.A(_10828_),
    .X(_10829_));
 sg13g2_buf_1 _17420_ (.A(net304),
    .X(_10830_));
 sg13g2_buf_8 _17421_ (.A(_10825_),
    .X(_10831_));
 sg13g2_nand3_1 _17422_ (.B(net784),
    .C(_10831_),
    .A(net767),
    .Y(_10832_));
 sg13g2_buf_2 _17423_ (.A(_10832_),
    .X(_10833_));
 sg13g2_buf_1 _17424_ (.A(_10833_),
    .X(_10834_));
 sg13g2_nand2_1 _17425_ (.Y(_10835_),
    .A(\top_ihp.oisc.regs[33][0] ),
    .B(net303));
 sg13g2_o21ai_1 _17426_ (.B1(_10835_),
    .Y(_01284_),
    .A1(net53),
    .A2(_10830_));
 sg13g2_nand2_1 _17427_ (.Y(_10836_),
    .A(\top_ihp.oisc.regs[33][10] ),
    .B(net303));
 sg13g2_o21ai_1 _17428_ (.B1(_10836_),
    .Y(_01285_),
    .A1(net155),
    .A2(net120));
 sg13g2_nand2_1 _17429_ (.Y(_10837_),
    .A(\top_ihp.oisc.regs[33][11] ),
    .B(net303));
 sg13g2_o21ai_1 _17430_ (.B1(_10837_),
    .Y(_01286_),
    .A1(net154),
    .A2(net120));
 sg13g2_nand2_1 _17431_ (.Y(_10838_),
    .A(\top_ihp.oisc.regs[33][12] ),
    .B(net304));
 sg13g2_o21ai_1 _17432_ (.B1(_10838_),
    .Y(_01287_),
    .A1(net137),
    .A2(net120));
 sg13g2_nand2_1 _17433_ (.Y(_10839_),
    .A(\top_ihp.oisc.regs[33][13] ),
    .B(net303));
 sg13g2_o21ai_1 _17434_ (.B1(_10839_),
    .Y(_01288_),
    .A1(net331),
    .A2(net120));
 sg13g2_nand2_1 _17435_ (.Y(_10840_),
    .A(\top_ihp.oisc.regs[33][14] ),
    .B(net304));
 sg13g2_o21ai_1 _17436_ (.B1(_10840_),
    .Y(_01289_),
    .A1(net136),
    .A2(net120));
 sg13g2_nand2_1 _17437_ (.Y(_10841_),
    .A(\top_ihp.oisc.regs[33][15] ),
    .B(net304));
 sg13g2_o21ai_1 _17438_ (.B1(_10841_),
    .Y(_01290_),
    .A1(_10536_),
    .A2(net120));
 sg13g2_nand2_1 _17439_ (.Y(_10842_),
    .A(\top_ihp.oisc.regs[33][16] ),
    .B(net303));
 sg13g2_o21ai_1 _17440_ (.B1(_10842_),
    .Y(_01291_),
    .A1(_10015_),
    .A2(net120));
 sg13g2_nand2_1 _17441_ (.Y(_10843_),
    .A(\top_ihp.oisc.regs[33][17] ),
    .B(net303));
 sg13g2_o21ai_1 _17442_ (.B1(_10843_),
    .Y(_01292_),
    .A1(net328),
    .A2(_10830_));
 sg13g2_nand2_1 _17443_ (.Y(_10844_),
    .A(\top_ihp.oisc.regs[33][18] ),
    .B(net303));
 sg13g2_o21ai_1 _17444_ (.B1(_10844_),
    .Y(_01293_),
    .A1(net327),
    .A2(net120));
 sg13g2_buf_1 _17445_ (.A(net304),
    .X(_10845_));
 sg13g2_nand2_1 _17446_ (.Y(_10846_),
    .A(\top_ihp.oisc.regs[33][19] ),
    .B(net303));
 sg13g2_o21ai_1 _17447_ (.B1(_10846_),
    .Y(_01294_),
    .A1(net326),
    .A2(net119));
 sg13g2_nand2_1 _17448_ (.Y(_10847_),
    .A(\top_ihp.oisc.regs[33][1] ),
    .B(net304));
 sg13g2_o21ai_1 _17449_ (.B1(_10847_),
    .Y(_01295_),
    .A1(net134),
    .A2(net119));
 sg13g2_buf_1 _17450_ (.A(_10833_),
    .X(_10848_));
 sg13g2_nand2_1 _17451_ (.Y(_10849_),
    .A(\top_ihp.oisc.regs[33][20] ),
    .B(_10848_));
 sg13g2_o21ai_1 _17452_ (.B1(_10849_),
    .Y(_01296_),
    .A1(net653),
    .A2(_10834_));
 sg13g2_nand2_1 _17453_ (.Y(_10850_),
    .A(\top_ihp.oisc.regs[33][21] ),
    .B(net302));
 sg13g2_o21ai_1 _17454_ (.B1(_10850_),
    .Y(_01297_),
    .A1(net323),
    .A2(net119));
 sg13g2_nand2_1 _17455_ (.Y(_10851_),
    .A(\top_ihp.oisc.regs[33][22] ),
    .B(net304));
 sg13g2_o21ai_1 _17456_ (.B1(_10851_),
    .Y(_01298_),
    .A1(net133),
    .A2(net119));
 sg13g2_nand2_1 _17457_ (.Y(_10852_),
    .A(\top_ihp.oisc.regs[33][23] ),
    .B(_10829_));
 sg13g2_o21ai_1 _17458_ (.B1(_10852_),
    .Y(_01299_),
    .A1(_10204_),
    .A2(net119));
 sg13g2_nand2_1 _17459_ (.Y(_10853_),
    .A(\top_ihp.oisc.regs[33][24] ),
    .B(net302));
 sg13g2_o21ai_1 _17460_ (.B1(_10853_),
    .Y(_01300_),
    .A1(net320),
    .A2(net119));
 sg13g2_nand2_1 _17461_ (.Y(_10854_),
    .A(\top_ihp.oisc.regs[33][25] ),
    .B(net304));
 sg13g2_o21ai_1 _17462_ (.B1(_10854_),
    .Y(_01301_),
    .A1(net132),
    .A2(net119));
 sg13g2_nand2_1 _17463_ (.Y(_10855_),
    .A(\top_ihp.oisc.regs[33][26] ),
    .B(net302));
 sg13g2_o21ai_1 _17464_ (.B1(_10855_),
    .Y(_01302_),
    .A1(net146),
    .A2(_10845_));
 sg13g2_nand2_1 _17465_ (.Y(_10856_),
    .A(\top_ihp.oisc.regs[33][27] ),
    .B(net302));
 sg13g2_o21ai_1 _17466_ (.B1(_10856_),
    .Y(_01303_),
    .A1(net318),
    .A2(_10845_));
 sg13g2_nand2_1 _17467_ (.Y(_10857_),
    .A(\top_ihp.oisc.regs[33][28] ),
    .B(net302));
 sg13g2_o21ai_1 _17468_ (.B1(_10857_),
    .Y(_01304_),
    .A1(net525),
    .A2(net119));
 sg13g2_buf_1 _17469_ (.A(_10828_),
    .X(_10858_));
 sg13g2_nand2_1 _17470_ (.Y(_10859_),
    .A(\top_ihp.oisc.regs[33][29] ),
    .B(net302));
 sg13g2_o21ai_1 _17471_ (.B1(_10859_),
    .Y(_01305_),
    .A1(net317),
    .A2(_10858_));
 sg13g2_nand2_1 _17472_ (.Y(_10860_),
    .A(\top_ihp.oisc.regs[33][2] ),
    .B(_10848_));
 sg13g2_o21ai_1 _17473_ (.B1(_10860_),
    .Y(_01306_),
    .A1(net145),
    .A2(net301));
 sg13g2_nand2_1 _17474_ (.Y(_10861_),
    .A(\top_ihp.oisc.regs[33][30] ),
    .B(net302));
 sg13g2_o21ai_1 _17475_ (.B1(_10861_),
    .Y(_01307_),
    .A1(net144),
    .A2(_10858_));
 sg13g2_nand2_1 _17476_ (.Y(_10862_),
    .A(\top_ihp.oisc.regs[33][31] ),
    .B(_10829_));
 sg13g2_o21ai_1 _17477_ (.B1(_10862_),
    .Y(_01308_),
    .A1(net315),
    .A2(net301));
 sg13g2_nand2_1 _17478_ (.Y(_10863_),
    .A(\top_ihp.oisc.regs[33][3] ),
    .B(net302));
 sg13g2_o21ai_1 _17479_ (.B1(_10863_),
    .Y(_01309_),
    .A1(net143),
    .A2(net301));
 sg13g2_nand2_1 _17480_ (.Y(_10864_),
    .A(\top_ihp.oisc.regs[33][4] ),
    .B(_10833_));
 sg13g2_o21ai_1 _17481_ (.B1(_10864_),
    .Y(_01310_),
    .A1(net142),
    .A2(net301));
 sg13g2_nand2_1 _17482_ (.Y(_10865_),
    .A(\top_ihp.oisc.regs[33][5] ),
    .B(_10833_));
 sg13g2_o21ai_1 _17483_ (.B1(_10865_),
    .Y(_01311_),
    .A1(net141),
    .A2(net301));
 sg13g2_nand2_1 _17484_ (.Y(_10866_),
    .A(\top_ihp.oisc.regs[33][6] ),
    .B(_10833_));
 sg13g2_o21ai_1 _17485_ (.B1(_10866_),
    .Y(_01312_),
    .A1(net140),
    .A2(net301));
 sg13g2_nand2_1 _17486_ (.Y(_10867_),
    .A(\top_ihp.oisc.regs[33][7] ),
    .B(_10833_));
 sg13g2_o21ai_1 _17487_ (.B1(_10867_),
    .Y(_01313_),
    .A1(net518),
    .A2(_10834_));
 sg13g2_nand2_1 _17488_ (.Y(_10868_),
    .A(\top_ihp.oisc.regs[33][8] ),
    .B(_10833_));
 sg13g2_o21ai_1 _17489_ (.B1(_10868_),
    .Y(_01314_),
    .A1(net316),
    .A2(net301));
 sg13g2_nand2_1 _17490_ (.Y(_10869_),
    .A(\top_ihp.oisc.regs[33][9] ),
    .B(_10833_));
 sg13g2_o21ai_1 _17491_ (.B1(_10869_),
    .Y(_01315_),
    .A1(net138),
    .A2(net301));
 sg13g2_buf_1 _17492_ (.A(_10522_),
    .X(_10870_));
 sg13g2_nand3_1 _17493_ (.B(net741),
    .C(net708),
    .A(net767),
    .Y(_10871_));
 sg13g2_buf_1 _17494_ (.A(_10871_),
    .X(_10872_));
 sg13g2_buf_1 _17495_ (.A(_10872_),
    .X(_10873_));
 sg13g2_buf_1 _17496_ (.A(_10872_),
    .X(_10874_));
 sg13g2_nand2_1 _17497_ (.Y(_10875_),
    .A(\top_ihp.oisc.regs[34][0] ),
    .B(net299));
 sg13g2_o21ai_1 _17498_ (.B1(_10875_),
    .Y(_01316_),
    .A1(net53),
    .A2(net300));
 sg13g2_nand2_1 _17499_ (.Y(_10876_),
    .A(\top_ihp.oisc.regs[34][10] ),
    .B(net299));
 sg13g2_o21ai_1 _17500_ (.B1(_10876_),
    .Y(_01317_),
    .A1(_09825_),
    .A2(net300));
 sg13g2_nand2_1 _17501_ (.Y(_10877_),
    .A(\top_ihp.oisc.regs[34][11] ),
    .B(net299));
 sg13g2_o21ai_1 _17502_ (.B1(_10877_),
    .Y(_01318_),
    .A1(_09861_),
    .A2(_10873_));
 sg13g2_nand2_1 _17503_ (.Y(_10878_),
    .A(\top_ihp.oisc.regs[34][12] ),
    .B(net299));
 sg13g2_o21ai_1 _17504_ (.B1(_10878_),
    .Y(_01319_),
    .A1(net137),
    .A2(net300));
 sg13g2_nand2_1 _17505_ (.Y(_10879_),
    .A(\top_ihp.oisc.regs[34][13] ),
    .B(net299));
 sg13g2_o21ai_1 _17506_ (.B1(_10879_),
    .Y(_01320_),
    .A1(_09942_),
    .A2(net300));
 sg13g2_nand2_1 _17507_ (.Y(_10880_),
    .A(\top_ihp.oisc.regs[34][14] ),
    .B(net299));
 sg13g2_o21ai_1 _17508_ (.B1(_10880_),
    .Y(_01321_),
    .A1(net136),
    .A2(net300));
 sg13g2_buf_8 _17509_ (.A(_10825_),
    .X(_10881_));
 sg13g2_nand2_2 _17510_ (.Y(_10882_),
    .A(net741),
    .B(net706));
 sg13g2_nor2b_2 _17511_ (.A(_10882_),
    .B_N(net767),
    .Y(_10883_));
 sg13g2_mux2_1 _17512_ (.A0(_00304_),
    .A1(net329),
    .S(_10883_),
    .X(_01322_));
 sg13g2_nand2_1 _17513_ (.Y(_10884_),
    .A(\top_ihp.oisc.regs[34][16] ),
    .B(_10874_));
 sg13g2_o21ai_1 _17514_ (.B1(_10884_),
    .Y(_01323_),
    .A1(_10015_),
    .A2(net300));
 sg13g2_nand2_1 _17515_ (.Y(_10885_),
    .A(\top_ihp.oisc.regs[34][17] ),
    .B(net299));
 sg13g2_o21ai_1 _17516_ (.B1(_10885_),
    .Y(_01324_),
    .A1(_10039_),
    .A2(net300));
 sg13g2_nand2_1 _17517_ (.Y(_10886_),
    .A(\top_ihp.oisc.regs[34][18] ),
    .B(_10874_));
 sg13g2_o21ai_1 _17518_ (.B1(_10886_),
    .Y(_01325_),
    .A1(_10060_),
    .A2(_10873_));
 sg13g2_nand2_1 _17519_ (.Y(_10887_),
    .A(\top_ihp.oisc.regs[34][19] ),
    .B(net299));
 sg13g2_o21ai_1 _17520_ (.B1(_10887_),
    .Y(_01326_),
    .A1(_10085_),
    .A2(net300));
 sg13g2_buf_2 _17521_ (.A(_10872_),
    .X(_10888_));
 sg13g2_buf_1 _17522_ (.A(_10872_),
    .X(_10889_));
 sg13g2_nand2_1 _17523_ (.Y(_10890_),
    .A(\top_ihp.oisc.regs[34][1] ),
    .B(net297));
 sg13g2_o21ai_1 _17524_ (.B1(_10890_),
    .Y(_01327_),
    .A1(net134),
    .A2(net298));
 sg13g2_nand2_1 _17525_ (.Y(_10891_),
    .A(\top_ihp.oisc.regs[34][20] ),
    .B(net297));
 sg13g2_o21ai_1 _17526_ (.B1(_10891_),
    .Y(_01328_),
    .A1(net324),
    .A2(net298));
 sg13g2_nand2_1 _17527_ (.Y(_10892_),
    .A(\top_ihp.oisc.regs[34][21] ),
    .B(_10889_));
 sg13g2_o21ai_1 _17528_ (.B1(_10892_),
    .Y(_01329_),
    .A1(_10169_),
    .A2(_10888_));
 sg13g2_nand2_1 _17529_ (.Y(_10893_),
    .A(\top_ihp.oisc.regs[34][22] ),
    .B(net297));
 sg13g2_o21ai_1 _17530_ (.B1(_10893_),
    .Y(_01330_),
    .A1(net133),
    .A2(net298));
 sg13g2_nand2_1 _17531_ (.Y(_10894_),
    .A(\top_ihp.oisc.regs[34][23] ),
    .B(net297));
 sg13g2_o21ai_1 _17532_ (.B1(_10894_),
    .Y(_01331_),
    .A1(_10204_),
    .A2(net298));
 sg13g2_nand2_1 _17533_ (.Y(_10895_),
    .A(\top_ihp.oisc.regs[34][24] ),
    .B(net297));
 sg13g2_o21ai_1 _17534_ (.B1(_10895_),
    .Y(_01332_),
    .A1(_10217_),
    .A2(net298));
 sg13g2_nand2_1 _17535_ (.Y(_10896_),
    .A(\top_ihp.oisc.regs[34][25] ),
    .B(net297));
 sg13g2_o21ai_1 _17536_ (.B1(_10896_),
    .Y(_01333_),
    .A1(net132),
    .A2(net298));
 sg13g2_nand2_1 _17537_ (.Y(_10897_),
    .A(\top_ihp.oisc.regs[34][26] ),
    .B(net297));
 sg13g2_o21ai_1 _17538_ (.B1(_10897_),
    .Y(_01334_),
    .A1(_10248_),
    .A2(net298));
 sg13g2_nand2_1 _17539_ (.Y(_10898_),
    .A(\top_ihp.oisc.regs[34][27] ),
    .B(_10889_));
 sg13g2_o21ai_1 _17540_ (.B1(_10898_),
    .Y(_01335_),
    .A1(_10260_),
    .A2(_10888_));
 sg13g2_nand2_1 _17541_ (.Y(_10899_),
    .A(\top_ihp.oisc.regs[34][28] ),
    .B(net297));
 sg13g2_o21ai_1 _17542_ (.B1(_10899_),
    .Y(_01336_),
    .A1(_10269_),
    .A2(net298));
 sg13g2_buf_1 _17543_ (.A(_10872_),
    .X(_10900_));
 sg13g2_buf_1 _17544_ (.A(_10872_),
    .X(_10901_));
 sg13g2_nand2_1 _17545_ (.Y(_10902_),
    .A(\top_ihp.oisc.regs[34][29] ),
    .B(net295));
 sg13g2_o21ai_1 _17546_ (.B1(_10902_),
    .Y(_01337_),
    .A1(_10281_),
    .A2(net296));
 sg13g2_nand2_1 _17547_ (.Y(_10903_),
    .A(\top_ihp.oisc.regs[34][2] ),
    .B(net295));
 sg13g2_o21ai_1 _17548_ (.B1(_10903_),
    .Y(_01338_),
    .A1(net145),
    .A2(net296));
 sg13g2_nand2_1 _17549_ (.Y(_10904_),
    .A(\top_ihp.oisc.regs[34][30] ),
    .B(net295));
 sg13g2_o21ai_1 _17550_ (.B1(_10904_),
    .Y(_01339_),
    .A1(net144),
    .A2(net296));
 sg13g2_mux2_1 _17551_ (.A0(_00305_),
    .A1(_10348_),
    .S(_10883_),
    .X(_01340_));
 sg13g2_nand2_1 _17552_ (.Y(_10905_),
    .A(\top_ihp.oisc.regs[34][3] ),
    .B(_10901_));
 sg13g2_o21ai_1 _17553_ (.B1(_10905_),
    .Y(_01341_),
    .A1(net143),
    .A2(_10900_));
 sg13g2_nand2_1 _17554_ (.Y(_10906_),
    .A(\top_ihp.oisc.regs[34][4] ),
    .B(net295));
 sg13g2_o21ai_1 _17555_ (.B1(_10906_),
    .Y(_01342_),
    .A1(net142),
    .A2(net296));
 sg13g2_nand2_1 _17556_ (.Y(_10907_),
    .A(\top_ihp.oisc.regs[34][5] ),
    .B(net295));
 sg13g2_o21ai_1 _17557_ (.B1(_10907_),
    .Y(_01343_),
    .A1(_10440_),
    .A2(net296));
 sg13g2_nand2_1 _17558_ (.Y(_10908_),
    .A(\top_ihp.oisc.regs[34][6] ),
    .B(net295));
 sg13g2_o21ai_1 _17559_ (.B1(_10908_),
    .Y(_01344_),
    .A1(_10469_),
    .A2(net296));
 sg13g2_nand2_1 _17560_ (.Y(_10909_),
    .A(\top_ihp.oisc.regs[34][7] ),
    .B(_10901_));
 sg13g2_o21ai_1 _17561_ (.B1(_10909_),
    .Y(_01345_),
    .A1(net139),
    .A2(_10900_));
 sg13g2_nand2_1 _17562_ (.Y(_10910_),
    .A(\top_ihp.oisc.regs[34][8] ),
    .B(net295));
 sg13g2_o21ai_1 _17563_ (.B1(_10910_),
    .Y(_01346_),
    .A1(_10499_),
    .A2(net296));
 sg13g2_nand2_1 _17564_ (.Y(_10911_),
    .A(\top_ihp.oisc.regs[34][9] ),
    .B(net295));
 sg13g2_o21ai_1 _17565_ (.B1(_10911_),
    .Y(_01347_),
    .A1(net138),
    .A2(net296));
 sg13g2_nand3_1 _17566_ (.B(net785),
    .C(net708),
    .A(net767),
    .Y(_10912_));
 sg13g2_buf_2 _17567_ (.A(_10912_),
    .X(_10913_));
 sg13g2_buf_1 _17568_ (.A(_10913_),
    .X(_10914_));
 sg13g2_buf_1 _17569_ (.A(_10913_),
    .X(_10915_));
 sg13g2_nand2_1 _17570_ (.Y(_10916_),
    .A(\top_ihp.oisc.regs[35][0] ),
    .B(net293));
 sg13g2_o21ai_1 _17571_ (.B1(_10916_),
    .Y(_01348_),
    .A1(_09698_),
    .A2(net294));
 sg13g2_nand2_1 _17572_ (.Y(_10917_),
    .A(\top_ihp.oisc.regs[35][10] ),
    .B(net293));
 sg13g2_o21ai_1 _17573_ (.B1(_10917_),
    .Y(_01349_),
    .A1(_09825_),
    .A2(net294));
 sg13g2_mux2_1 _17574_ (.A0(net127),
    .A1(_00306_),
    .S(net293),
    .X(_01350_));
 sg13g2_nand2_1 _17575_ (.Y(_10918_),
    .A(\top_ihp.oisc.regs[35][12] ),
    .B(net293));
 sg13g2_o21ai_1 _17576_ (.B1(_10918_),
    .Y(_01351_),
    .A1(_10531_),
    .A2(net294));
 sg13g2_nand2_1 _17577_ (.Y(_10919_),
    .A(\top_ihp.oisc.regs[35][13] ),
    .B(net293));
 sg13g2_o21ai_1 _17578_ (.B1(_10919_),
    .Y(_01352_),
    .A1(_09942_),
    .A2(_10914_));
 sg13g2_nand2_1 _17579_ (.Y(_10920_),
    .A(\top_ihp.oisc.regs[35][14] ),
    .B(net293));
 sg13g2_o21ai_1 _17580_ (.B1(_10920_),
    .Y(_01353_),
    .A1(_10534_),
    .A2(net294));
 sg13g2_nand2_1 _17581_ (.Y(_10921_),
    .A(\top_ihp.oisc.regs[35][15] ),
    .B(_10915_));
 sg13g2_o21ai_1 _17582_ (.B1(_10921_),
    .Y(_01354_),
    .A1(net135),
    .A2(net294));
 sg13g2_nand2_1 _17583_ (.Y(_10922_),
    .A(\top_ihp.oisc.regs[35][16] ),
    .B(net293));
 sg13g2_o21ai_1 _17584_ (.B1(_10922_),
    .Y(_01355_),
    .A1(net150),
    .A2(net294));
 sg13g2_nand2_1 _17585_ (.Y(_10923_),
    .A(\top_ihp.oisc.regs[35][17] ),
    .B(net293));
 sg13g2_o21ai_1 _17586_ (.B1(_10923_),
    .Y(_01356_),
    .A1(_10039_),
    .A2(_10914_));
 sg13g2_buf_1 _17587_ (.A(_10913_),
    .X(_10924_));
 sg13g2_nand2_1 _17588_ (.Y(_10925_),
    .A(\top_ihp.oisc.regs[35][18] ),
    .B(net292));
 sg13g2_o21ai_1 _17589_ (.B1(_10925_),
    .Y(_01357_),
    .A1(_10060_),
    .A2(net294));
 sg13g2_nand2_1 _17590_ (.Y(_10926_),
    .A(\top_ihp.oisc.regs[35][19] ),
    .B(net292));
 sg13g2_o21ai_1 _17591_ (.B1(_10926_),
    .Y(_01358_),
    .A1(_10085_),
    .A2(net294));
 sg13g2_buf_1 _17592_ (.A(_10913_),
    .X(_10927_));
 sg13g2_nand2_1 _17593_ (.Y(_10928_),
    .A(\top_ihp.oisc.regs[35][1] ),
    .B(net292));
 sg13g2_o21ai_1 _17594_ (.B1(_10928_),
    .Y(_01359_),
    .A1(_10543_),
    .A2(net291));
 sg13g2_nand2_1 _17595_ (.Y(_10929_),
    .A(\top_ihp.oisc.regs[35][20] ),
    .B(net292));
 sg13g2_o21ai_1 _17596_ (.B1(_10929_),
    .Y(_01360_),
    .A1(net653),
    .A2(net291));
 sg13g2_nand2_1 _17597_ (.Y(_10930_),
    .A(\top_ihp.oisc.regs[35][21] ),
    .B(net292));
 sg13g2_o21ai_1 _17598_ (.B1(_10930_),
    .Y(_01361_),
    .A1(_10169_),
    .A2(_10927_));
 sg13g2_nand2_1 _17599_ (.Y(_10931_),
    .A(\top_ihp.oisc.regs[35][22] ),
    .B(net292));
 sg13g2_o21ai_1 _17600_ (.B1(_10931_),
    .Y(_01362_),
    .A1(_10548_),
    .A2(net291));
 sg13g2_nand2_1 _17601_ (.Y(_10932_),
    .A(\top_ihp.oisc.regs[35][23] ),
    .B(net292));
 sg13g2_o21ai_1 _17602_ (.B1(_10932_),
    .Y(_01363_),
    .A1(net321),
    .A2(net291));
 sg13g2_nand2_1 _17603_ (.Y(_10933_),
    .A(\top_ihp.oisc.regs[35][24] ),
    .B(net292));
 sg13g2_o21ai_1 _17604_ (.B1(_10933_),
    .Y(_01364_),
    .A1(_10217_),
    .A2(net291));
 sg13g2_nand2_1 _17605_ (.Y(_10934_),
    .A(\top_ihp.oisc.regs[35][25] ),
    .B(_10924_));
 sg13g2_o21ai_1 _17606_ (.B1(_10934_),
    .Y(_01365_),
    .A1(_10597_),
    .A2(_10927_));
 sg13g2_nand2_1 _17607_ (.Y(_10935_),
    .A(\top_ihp.oisc.regs[35][26] ),
    .B(_10924_));
 sg13g2_o21ai_1 _17608_ (.B1(_10935_),
    .Y(_01366_),
    .A1(_10248_),
    .A2(net291));
 sg13g2_buf_1 _17609_ (.A(_10913_),
    .X(_10936_));
 sg13g2_nand2_1 _17610_ (.Y(_10937_),
    .A(\top_ihp.oisc.regs[35][27] ),
    .B(net290));
 sg13g2_o21ai_1 _17611_ (.B1(_10937_),
    .Y(_01367_),
    .A1(_10260_),
    .A2(net291));
 sg13g2_nand2_1 _17612_ (.Y(_10938_),
    .A(\top_ihp.oisc.regs[35][28] ),
    .B(net290));
 sg13g2_o21ai_1 _17613_ (.B1(_10938_),
    .Y(_01368_),
    .A1(_10269_),
    .A2(net291));
 sg13g2_buf_1 _17614_ (.A(_10913_),
    .X(_10939_));
 sg13g2_nand2_1 _17615_ (.Y(_10940_),
    .A(\top_ihp.oisc.regs[35][29] ),
    .B(net290));
 sg13g2_o21ai_1 _17616_ (.B1(_10940_),
    .Y(_01369_),
    .A1(_10281_),
    .A2(net289));
 sg13g2_nand2_1 _17617_ (.Y(_10941_),
    .A(\top_ihp.oisc.regs[35][2] ),
    .B(net290));
 sg13g2_o21ai_1 _17618_ (.B1(_10941_),
    .Y(_01370_),
    .A1(_10315_),
    .A2(net289));
 sg13g2_nand2_1 _17619_ (.Y(_10942_),
    .A(\top_ihp.oisc.regs[35][30] ),
    .B(net290));
 sg13g2_o21ai_1 _17620_ (.B1(_10942_),
    .Y(_01371_),
    .A1(_10327_),
    .A2(net289));
 sg13g2_mux2_1 _17621_ (.A0(_10345_),
    .A1(_00307_),
    .S(_10915_),
    .X(_01372_));
 sg13g2_nand2_1 _17622_ (.Y(_10943_),
    .A(\top_ihp.oisc.regs[35][3] ),
    .B(_10936_));
 sg13g2_o21ai_1 _17623_ (.B1(_10943_),
    .Y(_01373_),
    .A1(_10381_),
    .A2(_10939_));
 sg13g2_nand2_1 _17624_ (.Y(_10944_),
    .A(\top_ihp.oisc.regs[35][4] ),
    .B(net290));
 sg13g2_o21ai_1 _17625_ (.B1(_10944_),
    .Y(_01374_),
    .A1(_10413_),
    .A2(net289));
 sg13g2_nand2_1 _17626_ (.Y(_10945_),
    .A(\top_ihp.oisc.regs[35][5] ),
    .B(_10936_));
 sg13g2_o21ai_1 _17627_ (.B1(_10945_),
    .Y(_01375_),
    .A1(_10440_),
    .A2(_10939_));
 sg13g2_nand2_1 _17628_ (.Y(_10946_),
    .A(\top_ihp.oisc.regs[35][6] ),
    .B(net290));
 sg13g2_o21ai_1 _17629_ (.B1(_10946_),
    .Y(_01376_),
    .A1(_10469_),
    .A2(net289));
 sg13g2_nand2_1 _17630_ (.Y(_10947_),
    .A(\top_ihp.oisc.regs[35][7] ),
    .B(net290));
 sg13g2_o21ai_1 _17631_ (.B1(_10947_),
    .Y(_01377_),
    .A1(net518),
    .A2(net289));
 sg13g2_nand2_1 _17632_ (.Y(_10948_),
    .A(\top_ihp.oisc.regs[35][8] ),
    .B(_10913_));
 sg13g2_o21ai_1 _17633_ (.B1(_10948_),
    .Y(_01378_),
    .A1(_10499_),
    .A2(net289));
 sg13g2_nand2_1 _17634_ (.Y(_10949_),
    .A(\top_ihp.oisc.regs[35][9] ),
    .B(_10913_));
 sg13g2_o21ai_1 _17635_ (.B1(_10949_),
    .Y(_01379_),
    .A1(_10514_),
    .A2(net289));
 sg13g2_nand2_1 _17636_ (.Y(_10950_),
    .A(_09494_),
    .B(_09702_));
 sg13g2_nand2_1 _17637_ (.Y(_10951_),
    .A(_09532_),
    .B(_09714_));
 sg13g2_and4_1 _17638_ (.A(_09723_),
    .B(_09722_),
    .C(_10950_),
    .D(_10951_),
    .X(_10952_));
 sg13g2_buf_2 _17639_ (.A(_10952_),
    .X(_10953_));
 sg13g2_nand3_1 _17640_ (.B(net708),
    .C(_10953_),
    .A(net766),
    .Y(_10954_));
 sg13g2_buf_1 _17641_ (.A(_10954_),
    .X(_10955_));
 sg13g2_buf_8 _17642_ (.A(_10955_),
    .X(_10956_));
 sg13g2_buf_1 _17643_ (.A(_10956_),
    .X(_10957_));
 sg13g2_buf_2 _17644_ (.A(_10955_),
    .X(_10958_));
 sg13g2_nand2_1 _17645_ (.Y(_10959_),
    .A(\top_ihp.oisc.regs[36][0] ),
    .B(net287));
 sg13g2_o21ai_1 _17646_ (.B1(_10959_),
    .Y(_01380_),
    .A1(_09698_),
    .A2(net118));
 sg13g2_buf_8 _17647_ (.A(net128),
    .X(_10960_));
 sg13g2_nand2_1 _17648_ (.Y(_10961_),
    .A(\top_ihp.oisc.regs[36][10] ),
    .B(net287));
 sg13g2_o21ai_1 _17649_ (.B1(_10961_),
    .Y(_01381_),
    .A1(_10960_),
    .A2(_10957_));
 sg13g2_nand2_1 _17650_ (.Y(_10962_),
    .A(\top_ihp.oisc.regs[36][11] ),
    .B(net287));
 sg13g2_o21ai_1 _17651_ (.B1(_10962_),
    .Y(_01382_),
    .A1(_09861_),
    .A2(net118));
 sg13g2_nand4_1 _17652_ (.B(_09722_),
    .C(_10950_),
    .A(_09723_),
    .Y(_10963_),
    .D(_10951_));
 sg13g2_buf_2 _17653_ (.A(_10963_),
    .X(_10964_));
 sg13g2_nand2_2 _17654_ (.Y(_10965_),
    .A(net766),
    .B(net707));
 sg13g2_nor2_2 _17655_ (.A(_10964_),
    .B(_10965_),
    .Y(_10966_));
 sg13g2_buf_8 _17656_ (.A(_10966_),
    .X(_10967_));
 sg13g2_nor2_1 _17657_ (.A(\top_ihp.oisc.regs[36][12] ),
    .B(net286),
    .Y(_10968_));
 sg13g2_a21oi_1 _17658_ (.A1(net153),
    .A2(net286),
    .Y(_01383_),
    .B1(_10968_));
 sg13g2_buf_8 _17659_ (.A(net314),
    .X(_10969_));
 sg13g2_nand2_1 _17660_ (.Y(_10970_),
    .A(\top_ihp.oisc.regs[36][13] ),
    .B(net287));
 sg13g2_o21ai_1 _17661_ (.B1(_10970_),
    .Y(_01384_),
    .A1(net117),
    .A2(net118));
 sg13g2_nor2_1 _17662_ (.A(\top_ihp.oisc.regs[36][14] ),
    .B(net286),
    .Y(_10971_));
 sg13g2_a21oi_1 _17663_ (.A1(net152),
    .A2(net286),
    .Y(_01385_),
    .B1(_10971_));
 sg13g2_nor2_1 _17664_ (.A(\top_ihp.oisc.regs[36][15] ),
    .B(net286),
    .Y(_10972_));
 sg13g2_a21oi_1 _17665_ (.A1(net151),
    .A2(net286),
    .Y(_01386_),
    .B1(_10972_));
 sg13g2_buf_8 _17666_ (.A(net126),
    .X(_10973_));
 sg13g2_nand2_1 _17667_ (.Y(_10974_),
    .A(\top_ihp.oisc.regs[36][16] ),
    .B(net287));
 sg13g2_o21ai_1 _17668_ (.B1(_10974_),
    .Y(_01387_),
    .A1(net50),
    .A2(net118));
 sg13g2_buf_1 _17669_ (.A(_10629_),
    .X(_10975_));
 sg13g2_nand2_1 _17670_ (.Y(_10976_),
    .A(\top_ihp.oisc.regs[36][17] ),
    .B(net287));
 sg13g2_o21ai_1 _17671_ (.B1(_10976_),
    .Y(_01388_),
    .A1(net116),
    .A2(net118));
 sg13g2_buf_1 _17672_ (.A(_10630_),
    .X(_10977_));
 sg13g2_nand2_1 _17673_ (.Y(_10978_),
    .A(\top_ihp.oisc.regs[36][18] ),
    .B(_10958_));
 sg13g2_o21ai_1 _17674_ (.B1(_10978_),
    .Y(_01389_),
    .A1(net115),
    .A2(net118));
 sg13g2_buf_8 _17675_ (.A(net311),
    .X(_10979_));
 sg13g2_buf_1 _17676_ (.A(_10956_),
    .X(_10980_));
 sg13g2_nand2_1 _17677_ (.Y(_10981_),
    .A(\top_ihp.oisc.regs[36][19] ),
    .B(net113));
 sg13g2_o21ai_1 _17678_ (.B1(_10981_),
    .Y(_01390_),
    .A1(_10979_),
    .A2(_10957_));
 sg13g2_nor2_1 _17679_ (.A(\top_ihp.oisc.regs[36][1] ),
    .B(net286),
    .Y(_10982_));
 sg13g2_a21oi_1 _17680_ (.A1(net149),
    .A2(_10967_),
    .Y(_01391_),
    .B1(_10982_));
 sg13g2_nand2_1 _17681_ (.Y(_10983_),
    .A(\top_ihp.oisc.regs[36][20] ),
    .B(net113));
 sg13g2_o21ai_1 _17682_ (.B1(_10983_),
    .Y(_01392_),
    .A1(_10591_),
    .A2(net118));
 sg13g2_buf_8 _17683_ (.A(_10633_),
    .X(_10984_));
 sg13g2_nand2_1 _17684_ (.Y(_10985_),
    .A(\top_ihp.oisc.regs[36][21] ),
    .B(net113));
 sg13g2_o21ai_1 _17685_ (.B1(_10985_),
    .Y(_01393_),
    .A1(net112),
    .A2(net118));
 sg13g2_nor2_1 _17686_ (.A(\top_ihp.oisc.regs[36][22] ),
    .B(_10966_),
    .Y(_10986_));
 sg13g2_a21oi_1 _17687_ (.A1(_10189_),
    .A2(net286),
    .Y(_01394_),
    .B1(_10986_));
 sg13g2_buf_8 _17688_ (.A(net528),
    .X(_10987_));
 sg13g2_buf_1 _17689_ (.A(_10953_),
    .X(_10988_));
 sg13g2_nand3_1 _17690_ (.B(net706),
    .C(net762),
    .A(net766),
    .Y(_10989_));
 sg13g2_buf_2 _17691_ (.A(_10989_),
    .X(_10990_));
 sg13g2_nand2_1 _17692_ (.Y(_10991_),
    .A(\top_ihp.oisc.regs[36][23] ),
    .B(_10990_));
 sg13g2_o21ai_1 _17693_ (.B1(_10991_),
    .Y(_01395_),
    .A1(net285),
    .A2(_10990_));
 sg13g2_buf_1 _17694_ (.A(net309),
    .X(_10992_));
 sg13g2_buf_1 _17695_ (.A(net288),
    .X(_10993_));
 sg13g2_nand2_1 _17696_ (.Y(_10994_),
    .A(\top_ihp.oisc.regs[36][24] ),
    .B(_10980_));
 sg13g2_o21ai_1 _17697_ (.B1(_10994_),
    .Y(_01396_),
    .A1(net111),
    .A2(_10993_));
 sg13g2_nor2_1 _17698_ (.A(\top_ihp.oisc.regs[36][25] ),
    .B(_10966_),
    .Y(_10995_));
 sg13g2_a21oi_1 _17699_ (.A1(net147),
    .A2(_10967_),
    .Y(_01397_),
    .B1(_10995_));
 sg13g2_buf_1 _17700_ (.A(net125),
    .X(_10996_));
 sg13g2_nand2_1 _17701_ (.Y(_10997_),
    .A(\top_ihp.oisc.regs[36][26] ),
    .B(net113));
 sg13g2_o21ai_1 _17702_ (.B1(_10997_),
    .Y(_01398_),
    .A1(net49),
    .A2(net110));
 sg13g2_buf_1 _17703_ (.A(net308),
    .X(_10998_));
 sg13g2_nand2_1 _17704_ (.Y(_10999_),
    .A(\top_ihp.oisc.regs[36][27] ),
    .B(_10980_));
 sg13g2_o21ai_1 _17705_ (.B1(_10999_),
    .Y(_01399_),
    .A1(net109),
    .A2(_10993_));
 sg13g2_buf_8 _17706_ (.A(net515),
    .X(_11000_));
 sg13g2_nand2_1 _17707_ (.Y(_11001_),
    .A(\top_ihp.oisc.regs[36][28] ),
    .B(net113));
 sg13g2_o21ai_1 _17708_ (.B1(_11001_),
    .Y(_01400_),
    .A1(_11000_),
    .A2(_10990_));
 sg13g2_buf_8 _17709_ (.A(net307),
    .X(_11002_));
 sg13g2_nand2_1 _17710_ (.Y(_11003_),
    .A(\top_ihp.oisc.regs[36][29] ),
    .B(net113));
 sg13g2_o21ai_1 _17711_ (.B1(_11003_),
    .Y(_01401_),
    .A1(net108),
    .A2(net110));
 sg13g2_nand2_1 _17712_ (.Y(_11004_),
    .A(\top_ihp.oisc.regs[36][2] ),
    .B(net113));
 sg13g2_o21ai_1 _17713_ (.B1(_11004_),
    .Y(_01402_),
    .A1(_10315_),
    .A2(net110));
 sg13g2_nand2_1 _17714_ (.Y(_11005_),
    .A(\top_ihp.oisc.regs[36][30] ),
    .B(net113));
 sg13g2_o21ai_1 _17715_ (.B1(_11005_),
    .Y(_01403_),
    .A1(_10327_),
    .A2(net110));
 sg13g2_nand2_1 _17716_ (.Y(_11006_),
    .A(\top_ihp.oisc.regs[36][31] ),
    .B(_10990_));
 sg13g2_o21ai_1 _17717_ (.B1(_11006_),
    .Y(_01404_),
    .A1(net315),
    .A2(_10990_));
 sg13g2_nand2_1 _17718_ (.Y(_11007_),
    .A(\top_ihp.oisc.regs[36][3] ),
    .B(net288));
 sg13g2_o21ai_1 _17719_ (.B1(_11007_),
    .Y(_01405_),
    .A1(_10381_),
    .A2(net110));
 sg13g2_nand2_1 _17720_ (.Y(_11008_),
    .A(\top_ihp.oisc.regs[36][4] ),
    .B(net288));
 sg13g2_o21ai_1 _17721_ (.B1(_11008_),
    .Y(_01406_),
    .A1(_10413_),
    .A2(net110));
 sg13g2_buf_1 _17722_ (.A(net123),
    .X(_11009_));
 sg13g2_nand2_1 _17723_ (.Y(_11010_),
    .A(\top_ihp.oisc.regs[36][5] ),
    .B(net288));
 sg13g2_o21ai_1 _17724_ (.B1(_11010_),
    .Y(_01407_),
    .A1(net48),
    .A2(net110));
 sg13g2_buf_1 _17725_ (.A(net122),
    .X(_11011_));
 sg13g2_nand2_1 _17726_ (.Y(_11012_),
    .A(\top_ihp.oisc.regs[36][6] ),
    .B(net288));
 sg13g2_o21ai_1 _17727_ (.B1(_11012_),
    .Y(_01408_),
    .A1(net47),
    .A2(net110));
 sg13g2_nand2_1 _17728_ (.Y(_11013_),
    .A(\top_ihp.oisc.regs[36][7] ),
    .B(net288));
 sg13g2_o21ai_1 _17729_ (.B1(_11013_),
    .Y(_01409_),
    .A1(net518),
    .A2(net287));
 sg13g2_buf_8 _17730_ (.A(net305),
    .X(_11014_));
 sg13g2_nand2_1 _17731_ (.Y(_11015_),
    .A(\top_ihp.oisc.regs[36][8] ),
    .B(net288));
 sg13g2_o21ai_1 _17732_ (.B1(_11015_),
    .Y(_01410_),
    .A1(net107),
    .A2(net287));
 sg13g2_buf_8 _17733_ (.A(net121),
    .X(_11016_));
 sg13g2_nand2_1 _17734_ (.Y(_11017_),
    .A(\top_ihp.oisc.regs[36][9] ),
    .B(net288));
 sg13g2_o21ai_1 _17735_ (.B1(_11017_),
    .Y(_01411_),
    .A1(net46),
    .A2(_10958_));
 sg13g2_buf_1 _17736_ (.A(net156),
    .X(_11018_));
 sg13g2_nand3_1 _17737_ (.B(net706),
    .C(net762),
    .A(net784),
    .Y(_11019_));
 sg13g2_buf_2 _17738_ (.A(_11019_),
    .X(_11020_));
 sg13g2_buf_1 _17739_ (.A(_11020_),
    .X(_11021_));
 sg13g2_nand3_1 _17740_ (.B(net707),
    .C(_10953_),
    .A(_10822_),
    .Y(_11022_));
 sg13g2_buf_1 _17741_ (.A(_11022_),
    .X(_11023_));
 sg13g2_buf_1 _17742_ (.A(net503),
    .X(_11024_));
 sg13g2_nand2_1 _17743_ (.Y(_11025_),
    .A(\top_ihp.oisc.regs[37][0] ),
    .B(net282));
 sg13g2_o21ai_1 _17744_ (.B1(_11025_),
    .Y(_01412_),
    .A1(net45),
    .A2(net283));
 sg13g2_nand2_1 _17745_ (.Y(_11026_),
    .A(\top_ihp.oisc.regs[37][10] ),
    .B(net282));
 sg13g2_o21ai_1 _17746_ (.B1(_11026_),
    .Y(_01413_),
    .A1(_10960_),
    .A2(net283));
 sg13g2_buf_8 _17747_ (.A(_10624_),
    .X(_11027_));
 sg13g2_nand2_1 _17748_ (.Y(_11028_),
    .A(\top_ihp.oisc.regs[37][11] ),
    .B(net282));
 sg13g2_o21ai_1 _17749_ (.B1(_11028_),
    .Y(_01414_),
    .A1(net44),
    .A2(net283));
 sg13g2_nand2_1 _17750_ (.Y(_11029_),
    .A(net784),
    .B(net707));
 sg13g2_nor2_1 _17751_ (.A(_11029_),
    .B(_10964_),
    .Y(_11030_));
 sg13g2_buf_1 _17752_ (.A(_11030_),
    .X(_11031_));
 sg13g2_nor2_1 _17753_ (.A(\top_ihp.oisc.regs[37][12] ),
    .B(net281),
    .Y(_11032_));
 sg13g2_a21oi_1 _17754_ (.A1(net153),
    .A2(net281),
    .Y(_01415_),
    .B1(_11032_));
 sg13g2_nand2_1 _17755_ (.Y(_11033_),
    .A(\top_ihp.oisc.regs[37][13] ),
    .B(net282));
 sg13g2_o21ai_1 _17756_ (.B1(_11033_),
    .Y(_01416_),
    .A1(net117),
    .A2(net283));
 sg13g2_nor2_1 _17757_ (.A(\top_ihp.oisc.regs[37][14] ),
    .B(net281),
    .Y(_11034_));
 sg13g2_a21oi_1 _17758_ (.A1(net152),
    .A2(net281),
    .Y(_01417_),
    .B1(_11034_));
 sg13g2_nor2_1 _17759_ (.A(\top_ihp.oisc.regs[37][15] ),
    .B(_11031_),
    .Y(_11035_));
 sg13g2_a21oi_1 _17760_ (.A1(net151),
    .A2(_11031_),
    .Y(_01418_),
    .B1(_11035_));
 sg13g2_nand2_1 _17761_ (.Y(_11036_),
    .A(\top_ihp.oisc.regs[37][16] ),
    .B(net282));
 sg13g2_o21ai_1 _17762_ (.B1(_11036_),
    .Y(_01419_),
    .A1(net50),
    .A2(net283));
 sg13g2_nand2_1 _17763_ (.Y(_11037_),
    .A(\top_ihp.oisc.regs[37][17] ),
    .B(net282));
 sg13g2_o21ai_1 _17764_ (.B1(_11037_),
    .Y(_01420_),
    .A1(net116),
    .A2(net283));
 sg13g2_nand2_1 _17765_ (.Y(_11038_),
    .A(\top_ihp.oisc.regs[37][18] ),
    .B(net282));
 sg13g2_o21ai_1 _17766_ (.B1(_11038_),
    .Y(_01421_),
    .A1(net115),
    .A2(net283));
 sg13g2_nand2_1 _17767_ (.Y(_11039_),
    .A(\top_ihp.oisc.regs[37][19] ),
    .B(_11024_));
 sg13g2_o21ai_1 _17768_ (.B1(_11039_),
    .Y(_01422_),
    .A1(net114),
    .A2(_11021_));
 sg13g2_nor2_1 _17769_ (.A(\top_ihp.oisc.regs[37][1] ),
    .B(net281),
    .Y(_11040_));
 sg13g2_a21oi_1 _17770_ (.A1(net149),
    .A2(net281),
    .Y(_01423_),
    .B1(_11040_));
 sg13g2_buf_1 _17771_ (.A(net503),
    .X(_11041_));
 sg13g2_nand2_1 _17772_ (.Y(_11042_),
    .A(\top_ihp.oisc.regs[37][20] ),
    .B(net280));
 sg13g2_o21ai_1 _17773_ (.B1(_11042_),
    .Y(_01424_),
    .A1(net653),
    .A2(_11024_));
 sg13g2_nand2_1 _17774_ (.Y(_11043_),
    .A(\top_ihp.oisc.regs[37][21] ),
    .B(net280));
 sg13g2_o21ai_1 _17775_ (.B1(_11043_),
    .Y(_01425_),
    .A1(net112),
    .A2(_11021_));
 sg13g2_nor2_1 _17776_ (.A(\top_ihp.oisc.regs[37][22] ),
    .B(_11030_),
    .Y(_11044_));
 sg13g2_a21oi_1 _17777_ (.A1(net148),
    .A2(net281),
    .Y(_01426_),
    .B1(_11044_));
 sg13g2_nand2_1 _17778_ (.Y(_11045_),
    .A(\top_ihp.oisc.regs[37][23] ),
    .B(net280));
 sg13g2_o21ai_1 _17779_ (.B1(_11045_),
    .Y(_01427_),
    .A1(net285),
    .A2(net283));
 sg13g2_buf_1 _17780_ (.A(_11020_),
    .X(_11046_));
 sg13g2_nand2_1 _17781_ (.Y(_11047_),
    .A(\top_ihp.oisc.regs[37][24] ),
    .B(net280));
 sg13g2_o21ai_1 _17782_ (.B1(_11047_),
    .Y(_01428_),
    .A1(net111),
    .A2(net279));
 sg13g2_nor2_1 _17783_ (.A(\top_ihp.oisc.regs[37][25] ),
    .B(_11030_),
    .Y(_11048_));
 sg13g2_a21oi_1 _17784_ (.A1(net147),
    .A2(net281),
    .Y(_01429_),
    .B1(_11048_));
 sg13g2_nand2_1 _17785_ (.Y(_11049_),
    .A(\top_ihp.oisc.regs[37][26] ),
    .B(net280));
 sg13g2_o21ai_1 _17786_ (.B1(_11049_),
    .Y(_01430_),
    .A1(_10996_),
    .A2(net279));
 sg13g2_nand2_1 _17787_ (.Y(_11050_),
    .A(\top_ihp.oisc.regs[37][27] ),
    .B(_11041_));
 sg13g2_o21ai_1 _17788_ (.B1(_11050_),
    .Y(_01431_),
    .A1(net109),
    .A2(net279));
 sg13g2_nand2_1 _17789_ (.Y(_11051_),
    .A(\top_ihp.oisc.regs[37][28] ),
    .B(net280));
 sg13g2_o21ai_1 _17790_ (.B1(_11051_),
    .Y(_01432_),
    .A1(net284),
    .A2(net279));
 sg13g2_nand2_1 _17791_ (.Y(_11052_),
    .A(\top_ihp.oisc.regs[37][29] ),
    .B(net280));
 sg13g2_o21ai_1 _17792_ (.B1(_11052_),
    .Y(_01433_),
    .A1(net108),
    .A2(net279));
 sg13g2_buf_1 _17793_ (.A(net131),
    .X(_11053_));
 sg13g2_nand2_1 _17794_ (.Y(_11054_),
    .A(\top_ihp.oisc.regs[37][2] ),
    .B(_11041_));
 sg13g2_o21ai_1 _17795_ (.B1(_11054_),
    .Y(_01434_),
    .A1(net43),
    .A2(_11046_));
 sg13g2_buf_8 _17796_ (.A(net124),
    .X(_11055_));
 sg13g2_nand2_1 _17797_ (.Y(_11056_),
    .A(\top_ihp.oisc.regs[37][30] ),
    .B(net280));
 sg13g2_o21ai_1 _17798_ (.B1(_11056_),
    .Y(_01435_),
    .A1(net42),
    .A2(_11046_));
 sg13g2_nand2_1 _17799_ (.Y(_11057_),
    .A(\top_ihp.oisc.regs[37][31] ),
    .B(_11020_));
 sg13g2_o21ai_1 _17800_ (.B1(_11057_),
    .Y(_01436_),
    .A1(net315),
    .A2(net279));
 sg13g2_buf_2 _17801_ (.A(net130),
    .X(_11058_));
 sg13g2_nand2_1 _17802_ (.Y(_11059_),
    .A(\top_ihp.oisc.regs[37][3] ),
    .B(net503));
 sg13g2_o21ai_1 _17803_ (.B1(_11059_),
    .Y(_01437_),
    .A1(net41),
    .A2(net279));
 sg13g2_buf_1 _17804_ (.A(net129),
    .X(_11060_));
 sg13g2_nand2_1 _17805_ (.Y(_11061_),
    .A(\top_ihp.oisc.regs[37][4] ),
    .B(net503));
 sg13g2_o21ai_1 _17806_ (.B1(_11061_),
    .Y(_01438_),
    .A1(net40),
    .A2(net279));
 sg13g2_nand2_1 _17807_ (.Y(_11062_),
    .A(\top_ihp.oisc.regs[37][5] ),
    .B(net503));
 sg13g2_o21ai_1 _17808_ (.B1(_11062_),
    .Y(_01439_),
    .A1(net48),
    .A2(_11020_));
 sg13g2_nand2_1 _17809_ (.Y(_11063_),
    .A(\top_ihp.oisc.regs[37][6] ),
    .B(net503));
 sg13g2_o21ai_1 _17810_ (.B1(_11063_),
    .Y(_01440_),
    .A1(net47),
    .A2(_11020_));
 sg13g2_nand2_1 _17811_ (.Y(_11064_),
    .A(\top_ihp.oisc.regs[37][7] ),
    .B(net503));
 sg13g2_o21ai_1 _17812_ (.B1(_11064_),
    .Y(_01441_),
    .A1(net518),
    .A2(net282));
 sg13g2_nand2_1 _17813_ (.Y(_11065_),
    .A(\top_ihp.oisc.regs[37][8] ),
    .B(_11023_));
 sg13g2_o21ai_1 _17814_ (.B1(_11065_),
    .Y(_01442_),
    .A1(net107),
    .A2(_11020_));
 sg13g2_nand2_1 _17815_ (.Y(_11066_),
    .A(\top_ihp.oisc.regs[37][9] ),
    .B(net503));
 sg13g2_o21ai_1 _17816_ (.B1(_11066_),
    .Y(_01443_),
    .A1(net46),
    .A2(_11020_));
 sg13g2_nand3_1 _17817_ (.B(net706),
    .C(net762),
    .A(net741),
    .Y(_11067_));
 sg13g2_buf_8 _17818_ (.A(_11067_),
    .X(_11068_));
 sg13g2_buf_1 _17819_ (.A(net502),
    .X(_11069_));
 sg13g2_nand3_1 _17820_ (.B(net707),
    .C(net762),
    .A(net741),
    .Y(_11070_));
 sg13g2_buf_2 _17821_ (.A(_11070_),
    .X(_11071_));
 sg13g2_buf_1 _17822_ (.A(_11071_),
    .X(_11072_));
 sg13g2_nand2_1 _17823_ (.Y(_11073_),
    .A(\top_ihp.oisc.regs[38][0] ),
    .B(net277));
 sg13g2_o21ai_1 _17824_ (.B1(_11073_),
    .Y(_01444_),
    .A1(net45),
    .A2(net278));
 sg13g2_nand2_1 _17825_ (.Y(_11074_),
    .A(\top_ihp.oisc.regs[38][10] ),
    .B(net277));
 sg13g2_o21ai_1 _17826_ (.B1(_11074_),
    .Y(_01445_),
    .A1(net51),
    .A2(net278));
 sg13g2_nand2_1 _17827_ (.Y(_11075_),
    .A(\top_ihp.oisc.regs[38][11] ),
    .B(net277));
 sg13g2_o21ai_1 _17828_ (.B1(_11075_),
    .Y(_01446_),
    .A1(net44),
    .A2(net278));
 sg13g2_nor2_2 _17829_ (.A(_10882_),
    .B(_10964_),
    .Y(_11076_));
 sg13g2_buf_8 _17830_ (.A(_11076_),
    .X(_11077_));
 sg13g2_nor2_1 _17831_ (.A(\top_ihp.oisc.regs[38][12] ),
    .B(net276),
    .Y(_11078_));
 sg13g2_a21oi_1 _17832_ (.A1(net153),
    .A2(net276),
    .Y(_01447_),
    .B1(_11078_));
 sg13g2_nand2_1 _17833_ (.Y(_11079_),
    .A(\top_ihp.oisc.regs[38][13] ),
    .B(net277));
 sg13g2_o21ai_1 _17834_ (.B1(_11079_),
    .Y(_01448_),
    .A1(net117),
    .A2(net278));
 sg13g2_nor2_1 _17835_ (.A(\top_ihp.oisc.regs[38][14] ),
    .B(net276),
    .Y(_11080_));
 sg13g2_a21oi_1 _17836_ (.A1(net152),
    .A2(net276),
    .Y(_01449_),
    .B1(_11080_));
 sg13g2_nor2_1 _17837_ (.A(\top_ihp.oisc.regs[38][15] ),
    .B(net276),
    .Y(_11081_));
 sg13g2_a21oi_1 _17838_ (.A1(_09993_),
    .A2(net276),
    .Y(_01450_),
    .B1(_11081_));
 sg13g2_nand2_1 _17839_ (.Y(_11082_),
    .A(\top_ihp.oisc.regs[38][16] ),
    .B(net277));
 sg13g2_o21ai_1 _17840_ (.B1(_11082_),
    .Y(_01451_),
    .A1(net50),
    .A2(net278));
 sg13g2_nand2_1 _17841_ (.Y(_11083_),
    .A(\top_ihp.oisc.regs[38][17] ),
    .B(net277));
 sg13g2_o21ai_1 _17842_ (.B1(_11083_),
    .Y(_01452_),
    .A1(net116),
    .A2(net278));
 sg13g2_nand2_1 _17843_ (.Y(_11084_),
    .A(\top_ihp.oisc.regs[38][18] ),
    .B(_11072_));
 sg13g2_o21ai_1 _17844_ (.B1(_11084_),
    .Y(_01453_),
    .A1(_10977_),
    .A2(_11069_));
 sg13g2_nand2_1 _17845_ (.Y(_11085_),
    .A(\top_ihp.oisc.regs[38][19] ),
    .B(net277));
 sg13g2_o21ai_1 _17846_ (.B1(_11085_),
    .Y(_01454_),
    .A1(net114),
    .A2(net278));
 sg13g2_nor2_1 _17847_ (.A(\top_ihp.oisc.regs[38][1] ),
    .B(net276),
    .Y(_11086_));
 sg13g2_a21oi_1 _17848_ (.A1(net149),
    .A2(net276),
    .Y(_01455_),
    .B1(_11086_));
 sg13g2_nand2_1 _17849_ (.Y(_11087_),
    .A(\top_ihp.oisc.regs[38][20] ),
    .B(_11072_));
 sg13g2_o21ai_1 _17850_ (.B1(_11087_),
    .Y(_01456_),
    .A1(net324),
    .A2(_11069_));
 sg13g2_nand2_1 _17851_ (.Y(_11088_),
    .A(\top_ihp.oisc.regs[38][21] ),
    .B(net277));
 sg13g2_o21ai_1 _17852_ (.B1(_11088_),
    .Y(_01457_),
    .A1(net112),
    .A2(net278));
 sg13g2_nor2_1 _17853_ (.A(\top_ihp.oisc.regs[38][22] ),
    .B(_11076_),
    .Y(_11089_));
 sg13g2_a21oi_1 _17854_ (.A1(net148),
    .A2(_11077_),
    .Y(_01458_),
    .B1(_11089_));
 sg13g2_buf_8 _17855_ (.A(net502),
    .X(_11090_));
 sg13g2_buf_1 _17856_ (.A(_11071_),
    .X(_11091_));
 sg13g2_nand2_1 _17857_ (.Y(_11092_),
    .A(\top_ihp.oisc.regs[38][23] ),
    .B(net274));
 sg13g2_o21ai_1 _17858_ (.B1(_11092_),
    .Y(_01459_),
    .A1(net285),
    .A2(net275));
 sg13g2_nand2_1 _17859_ (.Y(_11093_),
    .A(\top_ihp.oisc.regs[38][24] ),
    .B(net274));
 sg13g2_o21ai_1 _17860_ (.B1(_11093_),
    .Y(_01460_),
    .A1(net111),
    .A2(net275));
 sg13g2_nor2_1 _17861_ (.A(\top_ihp.oisc.regs[38][25] ),
    .B(_11076_),
    .Y(_11094_));
 sg13g2_a21oi_1 _17862_ (.A1(net147),
    .A2(_11077_),
    .Y(_01461_),
    .B1(_11094_));
 sg13g2_nand2_1 _17863_ (.Y(_11095_),
    .A(\top_ihp.oisc.regs[38][26] ),
    .B(net274));
 sg13g2_o21ai_1 _17864_ (.B1(_11095_),
    .Y(_01462_),
    .A1(net49),
    .A2(net275));
 sg13g2_nand2_1 _17865_ (.Y(_11096_),
    .A(\top_ihp.oisc.regs[38][27] ),
    .B(net274));
 sg13g2_o21ai_1 _17866_ (.B1(_11096_),
    .Y(_01463_),
    .A1(net109),
    .A2(net275));
 sg13g2_nand2_1 _17867_ (.Y(_11097_),
    .A(\top_ihp.oisc.regs[38][28] ),
    .B(net274));
 sg13g2_o21ai_1 _17868_ (.B1(_11097_),
    .Y(_01464_),
    .A1(net284),
    .A2(net275));
 sg13g2_nand2_1 _17869_ (.Y(_11098_),
    .A(\top_ihp.oisc.regs[38][29] ),
    .B(net274));
 sg13g2_o21ai_1 _17870_ (.B1(_11098_),
    .Y(_01465_),
    .A1(net108),
    .A2(net275));
 sg13g2_nand2_1 _17871_ (.Y(_11099_),
    .A(\top_ihp.oisc.regs[38][2] ),
    .B(net274));
 sg13g2_o21ai_1 _17872_ (.B1(_11099_),
    .Y(_01466_),
    .A1(net43),
    .A2(net275));
 sg13g2_nand2_1 _17873_ (.Y(_11100_),
    .A(\top_ihp.oisc.regs[38][30] ),
    .B(_11091_));
 sg13g2_o21ai_1 _17874_ (.B1(_11100_),
    .Y(_01467_),
    .A1(_11055_),
    .A2(_11090_));
 sg13g2_nand2_1 _17875_ (.Y(_11101_),
    .A(\top_ihp.oisc.regs[38][31] ),
    .B(net502));
 sg13g2_o21ai_1 _17876_ (.B1(_11101_),
    .Y(_01468_),
    .A1(net52),
    .A2(net275));
 sg13g2_nand2_1 _17877_ (.Y(_11102_),
    .A(\top_ihp.oisc.regs[38][3] ),
    .B(_11091_));
 sg13g2_o21ai_1 _17878_ (.B1(_11102_),
    .Y(_01469_),
    .A1(net41),
    .A2(_11090_));
 sg13g2_nand2_1 _17879_ (.Y(_11103_),
    .A(\top_ihp.oisc.regs[38][4] ),
    .B(net274));
 sg13g2_o21ai_1 _17880_ (.B1(_11103_),
    .Y(_01470_),
    .A1(_11060_),
    .A2(net502));
 sg13g2_nand2_1 _17881_ (.Y(_11104_),
    .A(\top_ihp.oisc.regs[38][5] ),
    .B(_11071_));
 sg13g2_o21ai_1 _17882_ (.B1(_11104_),
    .Y(_01471_),
    .A1(net48),
    .A2(net502));
 sg13g2_nand2_1 _17883_ (.Y(_11105_),
    .A(\top_ihp.oisc.regs[38][6] ),
    .B(_11071_));
 sg13g2_o21ai_1 _17884_ (.B1(_11105_),
    .Y(_01472_),
    .A1(net47),
    .A2(net502));
 sg13g2_nand2_1 _17885_ (.Y(_11106_),
    .A(\top_ihp.oisc.regs[38][7] ),
    .B(_11071_));
 sg13g2_o21ai_1 _17886_ (.B1(_11106_),
    .Y(_01473_),
    .A1(net139),
    .A2(net502));
 sg13g2_nand2_1 _17887_ (.Y(_11107_),
    .A(\top_ihp.oisc.regs[38][8] ),
    .B(_11071_));
 sg13g2_o21ai_1 _17888_ (.B1(_11107_),
    .Y(_01474_),
    .A1(net107),
    .A2(net502));
 sg13g2_nand2_1 _17889_ (.Y(_11108_),
    .A(\top_ihp.oisc.regs[38][9] ),
    .B(_11071_));
 sg13g2_o21ai_1 _17890_ (.B1(_11108_),
    .Y(_01475_),
    .A1(net46),
    .A2(_11068_));
 sg13g2_nand3_1 _17891_ (.B(_10826_),
    .C(_10953_),
    .A(net785),
    .Y(_11109_));
 sg13g2_buf_1 _17892_ (.A(_11109_),
    .X(_11110_));
 sg13g2_buf_1 _17893_ (.A(_11110_),
    .X(_11111_));
 sg13g2_buf_1 _17894_ (.A(net273),
    .X(_11112_));
 sg13g2_nand3_1 _17895_ (.B(net707),
    .C(_10953_),
    .A(net785),
    .Y(_11113_));
 sg13g2_buf_2 _17896_ (.A(_11113_),
    .X(_11114_));
 sg13g2_buf_1 _17897_ (.A(_11114_),
    .X(_11115_));
 sg13g2_nand2_1 _17898_ (.Y(_11116_),
    .A(\top_ihp.oisc.regs[39][0] ),
    .B(net272));
 sg13g2_o21ai_1 _17899_ (.B1(_11116_),
    .Y(_01476_),
    .A1(_11018_),
    .A2(net106));
 sg13g2_nand2_1 _17900_ (.Y(_11117_),
    .A(\top_ihp.oisc.regs[39][10] ),
    .B(net272));
 sg13g2_o21ai_1 _17901_ (.B1(_11117_),
    .Y(_01477_),
    .A1(net51),
    .A2(net106));
 sg13g2_nand2_1 _17902_ (.Y(_11118_),
    .A(\top_ihp.oisc.regs[39][11] ),
    .B(net272));
 sg13g2_o21ai_1 _17903_ (.B1(_11118_),
    .Y(_01478_),
    .A1(_11027_),
    .A2(net106));
 sg13g2_nand2_1 _17904_ (.Y(_11119_),
    .A(\top_ihp.oisc.regs[39][12] ),
    .B(net273));
 sg13g2_o21ai_1 _17905_ (.B1(_11119_),
    .Y(_01479_),
    .A1(_10531_),
    .A2(net106));
 sg13g2_nand2_1 _17906_ (.Y(_11120_),
    .A(\top_ihp.oisc.regs[39][13] ),
    .B(net272));
 sg13g2_o21ai_1 _17907_ (.B1(_11120_),
    .Y(_01480_),
    .A1(net117),
    .A2(_11112_));
 sg13g2_nand2_1 _17908_ (.Y(_11121_),
    .A(\top_ihp.oisc.regs[39][14] ),
    .B(net273));
 sg13g2_o21ai_1 _17909_ (.B1(_11121_),
    .Y(_01481_),
    .A1(_10534_),
    .A2(net106));
 sg13g2_nand2_1 _17910_ (.Y(_11122_),
    .A(\top_ihp.oisc.regs[39][15] ),
    .B(net273));
 sg13g2_o21ai_1 _17911_ (.B1(_11122_),
    .Y(_01482_),
    .A1(_10536_),
    .A2(net106));
 sg13g2_nand2_1 _17912_ (.Y(_11123_),
    .A(\top_ihp.oisc.regs[39][16] ),
    .B(net272));
 sg13g2_o21ai_1 _17913_ (.B1(_11123_),
    .Y(_01483_),
    .A1(net50),
    .A2(_11112_));
 sg13g2_nand2_1 _17914_ (.Y(_11124_),
    .A(\top_ihp.oisc.regs[39][17] ),
    .B(net272));
 sg13g2_o21ai_1 _17915_ (.B1(_11124_),
    .Y(_01484_),
    .A1(net116),
    .A2(net106));
 sg13g2_nand2_1 _17916_ (.Y(_11125_),
    .A(\top_ihp.oisc.regs[39][18] ),
    .B(net272));
 sg13g2_o21ai_1 _17917_ (.B1(_11125_),
    .Y(_01485_),
    .A1(net115),
    .A2(net106));
 sg13g2_buf_1 _17918_ (.A(net273),
    .X(_11126_));
 sg13g2_nand2_1 _17919_ (.Y(_11127_),
    .A(\top_ihp.oisc.regs[39][19] ),
    .B(_11115_));
 sg13g2_o21ai_1 _17920_ (.B1(_11127_),
    .Y(_01486_),
    .A1(net114),
    .A2(net105));
 sg13g2_nand2_1 _17921_ (.Y(_11128_),
    .A(\top_ihp.oisc.regs[39][1] ),
    .B(net273));
 sg13g2_o21ai_1 _17922_ (.B1(_11128_),
    .Y(_01487_),
    .A1(_10543_),
    .A2(net105));
 sg13g2_buf_1 _17923_ (.A(_11114_),
    .X(_11129_));
 sg13g2_nand2_1 _17924_ (.Y(_11130_),
    .A(\top_ihp.oisc.regs[39][20] ),
    .B(net271));
 sg13g2_o21ai_1 _17925_ (.B1(_11130_),
    .Y(_01488_),
    .A1(net653),
    .A2(_11115_));
 sg13g2_nand2_1 _17926_ (.Y(_11131_),
    .A(\top_ihp.oisc.regs[39][21] ),
    .B(net271));
 sg13g2_o21ai_1 _17927_ (.B1(_11131_),
    .Y(_01489_),
    .A1(net112),
    .A2(net105));
 sg13g2_nand2_1 _17928_ (.Y(_11132_),
    .A(\top_ihp.oisc.regs[39][22] ),
    .B(net273));
 sg13g2_o21ai_1 _17929_ (.B1(_11132_),
    .Y(_01490_),
    .A1(_10548_),
    .A2(net105));
 sg13g2_nand2_1 _17930_ (.Y(_11133_),
    .A(\top_ihp.oisc.regs[39][23] ),
    .B(_11111_));
 sg13g2_o21ai_1 _17931_ (.B1(_11133_),
    .Y(_01491_),
    .A1(net285),
    .A2(net105));
 sg13g2_nand2_1 _17932_ (.Y(_11134_),
    .A(\top_ihp.oisc.regs[39][24] ),
    .B(net271));
 sg13g2_o21ai_1 _17933_ (.B1(_11134_),
    .Y(_01492_),
    .A1(net111),
    .A2(net105));
 sg13g2_nand2_1 _17934_ (.Y(_11135_),
    .A(\top_ihp.oisc.regs[39][25] ),
    .B(net273));
 sg13g2_o21ai_1 _17935_ (.B1(_11135_),
    .Y(_01493_),
    .A1(_10597_),
    .A2(net105));
 sg13g2_nand2_1 _17936_ (.Y(_11136_),
    .A(\top_ihp.oisc.regs[39][26] ),
    .B(net271));
 sg13g2_o21ai_1 _17937_ (.B1(_11136_),
    .Y(_01494_),
    .A1(net49),
    .A2(net105));
 sg13g2_nand2_1 _17938_ (.Y(_11137_),
    .A(\top_ihp.oisc.regs[39][27] ),
    .B(net271));
 sg13g2_o21ai_1 _17939_ (.B1(_11137_),
    .Y(_01495_),
    .A1(net109),
    .A2(_11126_));
 sg13g2_nand2_1 _17940_ (.Y(_11138_),
    .A(\top_ihp.oisc.regs[39][28] ),
    .B(_11129_));
 sg13g2_o21ai_1 _17941_ (.B1(_11138_),
    .Y(_01496_),
    .A1(_11000_),
    .A2(_11126_));
 sg13g2_buf_2 _17942_ (.A(_11110_),
    .X(_11139_));
 sg13g2_nand2_1 _17943_ (.Y(_11140_),
    .A(\top_ihp.oisc.regs[39][29] ),
    .B(net271));
 sg13g2_o21ai_1 _17944_ (.B1(_11140_),
    .Y(_01497_),
    .A1(net108),
    .A2(net270));
 sg13g2_nand2_1 _17945_ (.Y(_11141_),
    .A(\top_ihp.oisc.regs[39][2] ),
    .B(net271));
 sg13g2_o21ai_1 _17946_ (.B1(_11141_),
    .Y(_01498_),
    .A1(net43),
    .A2(net270));
 sg13g2_nand2_1 _17947_ (.Y(_11142_),
    .A(\top_ihp.oisc.regs[39][30] ),
    .B(_11129_));
 sg13g2_o21ai_1 _17948_ (.B1(_11142_),
    .Y(_01499_),
    .A1(net42),
    .A2(net270));
 sg13g2_nand2_1 _17949_ (.Y(_11143_),
    .A(\top_ihp.oisc.regs[39][31] ),
    .B(_11111_));
 sg13g2_o21ai_1 _17950_ (.B1(_11143_),
    .Y(_01500_),
    .A1(net315),
    .A2(net270));
 sg13g2_nand2_1 _17951_ (.Y(_11144_),
    .A(\top_ihp.oisc.regs[39][3] ),
    .B(net271));
 sg13g2_o21ai_1 _17952_ (.B1(_11144_),
    .Y(_01501_),
    .A1(net41),
    .A2(net270));
 sg13g2_nand2_1 _17953_ (.Y(_11145_),
    .A(\top_ihp.oisc.regs[39][4] ),
    .B(_11114_));
 sg13g2_o21ai_1 _17954_ (.B1(_11145_),
    .Y(_01502_),
    .A1(net40),
    .A2(net270));
 sg13g2_nand2_1 _17955_ (.Y(_11146_),
    .A(\top_ihp.oisc.regs[39][5] ),
    .B(_11114_));
 sg13g2_o21ai_1 _17956_ (.B1(_11146_),
    .Y(_01503_),
    .A1(_11009_),
    .A2(_11139_));
 sg13g2_nand2_1 _17957_ (.Y(_11147_),
    .A(\top_ihp.oisc.regs[39][6] ),
    .B(_11114_));
 sg13g2_o21ai_1 _17958_ (.B1(_11147_),
    .Y(_01504_),
    .A1(net47),
    .A2(_11139_));
 sg13g2_nand2_1 _17959_ (.Y(_11148_),
    .A(\top_ihp.oisc.regs[39][7] ),
    .B(_11114_));
 sg13g2_o21ai_1 _17960_ (.B1(_11148_),
    .Y(_01505_),
    .A1(_10612_),
    .A2(net272));
 sg13g2_nand2_1 _17961_ (.Y(_11149_),
    .A(\top_ihp.oisc.regs[39][8] ),
    .B(_11114_));
 sg13g2_o21ai_1 _17962_ (.B1(_11149_),
    .Y(_01506_),
    .A1(net107),
    .A2(net270));
 sg13g2_nand2_1 _17963_ (.Y(_11150_),
    .A(\top_ihp.oisc.regs[39][9] ),
    .B(_11114_));
 sg13g2_o21ai_1 _17964_ (.B1(_11150_),
    .Y(_01507_),
    .A1(net46),
    .A2(net270));
 sg13g2_nand2_1 _17965_ (.Y(_11151_),
    .A(net767),
    .B(_10572_));
 sg13g2_buf_1 _17966_ (.A(_11151_),
    .X(_11152_));
 sg13g2_buf_1 _17967_ (.A(net705),
    .X(_11153_));
 sg13g2_buf_1 _17968_ (.A(_11151_),
    .X(_11154_));
 sg13g2_nand2_1 _17969_ (.Y(_11155_),
    .A(\top_ihp.oisc.regs[3][0] ),
    .B(net704));
 sg13g2_o21ai_1 _17970_ (.B1(_11155_),
    .Y(_01508_),
    .A1(_11018_),
    .A2(net641));
 sg13g2_nand2_1 _17971_ (.Y(_11156_),
    .A(\top_ihp.oisc.regs[3][10] ),
    .B(net704));
 sg13g2_o21ai_1 _17972_ (.B1(_11156_),
    .Y(_01509_),
    .A1(net51),
    .A2(_11153_));
 sg13g2_nand2_1 _17973_ (.Y(_11157_),
    .A(\top_ihp.oisc.regs[3][11] ),
    .B(net704));
 sg13g2_o21ai_1 _17974_ (.B1(_11157_),
    .Y(_01510_),
    .A1(_11027_),
    .A2(net641));
 sg13g2_buf_8 _17975_ (.A(net332),
    .X(_11158_));
 sg13g2_nand2_1 _17976_ (.Y(_11159_),
    .A(\top_ihp.oisc.regs[3][12] ),
    .B(net704));
 sg13g2_o21ai_1 _17977_ (.B1(_11159_),
    .Y(_01511_),
    .A1(net104),
    .A2(net641));
 sg13g2_nand2_1 _17978_ (.Y(_11160_),
    .A(\top_ihp.oisc.regs[3][13] ),
    .B(net704));
 sg13g2_o21ai_1 _17979_ (.B1(_11160_),
    .Y(_01512_),
    .A1(_10969_),
    .A2(net641));
 sg13g2_buf_8 _17980_ (.A(net330),
    .X(_11161_));
 sg13g2_nand2_1 _17981_ (.Y(_11162_),
    .A(\top_ihp.oisc.regs[3][14] ),
    .B(net704));
 sg13g2_o21ai_1 _17982_ (.B1(_11162_),
    .Y(_01513_),
    .A1(net103),
    .A2(net641));
 sg13g2_nand2_1 _17983_ (.Y(_11163_),
    .A(\top_ihp.oisc.regs[3][15] ),
    .B(net704));
 sg13g2_o21ai_1 _17984_ (.B1(_11163_),
    .Y(_01514_),
    .A1(net135),
    .A2(net641));
 sg13g2_nand2_1 _17985_ (.Y(_11164_),
    .A(\top_ihp.oisc.regs[3][16] ),
    .B(net704));
 sg13g2_o21ai_1 _17986_ (.B1(_11164_),
    .Y(_01515_),
    .A1(net50),
    .A2(net641));
 sg13g2_buf_1 _17987_ (.A(net705),
    .X(_11165_));
 sg13g2_nand2_1 _17988_ (.Y(_11166_),
    .A(\top_ihp.oisc.regs[3][17] ),
    .B(net640));
 sg13g2_o21ai_1 _17989_ (.B1(_11166_),
    .Y(_01516_),
    .A1(net116),
    .A2(net641));
 sg13g2_nand2_1 _17990_ (.Y(_11167_),
    .A(\top_ihp.oisc.regs[3][18] ),
    .B(net640));
 sg13g2_o21ai_1 _17991_ (.B1(_11167_),
    .Y(_01517_),
    .A1(_10977_),
    .A2(_11153_));
 sg13g2_buf_1 _17992_ (.A(_11152_),
    .X(_11168_));
 sg13g2_nand2_1 _17993_ (.Y(_11169_),
    .A(\top_ihp.oisc.regs[3][19] ),
    .B(net640));
 sg13g2_o21ai_1 _17994_ (.B1(_11169_),
    .Y(_01518_),
    .A1(_10979_),
    .A2(net639));
 sg13g2_buf_2 _17995_ (.A(net325),
    .X(_11170_));
 sg13g2_nand2_1 _17996_ (.Y(_11171_),
    .A(\top_ihp.oisc.regs[3][1] ),
    .B(net640));
 sg13g2_o21ai_1 _17997_ (.B1(_11171_),
    .Y(_01519_),
    .A1(net102),
    .A2(net639));
 sg13g2_nand2_1 _17998_ (.Y(_11172_),
    .A(\top_ihp.oisc.regs[3][20] ),
    .B(_11165_));
 sg13g2_o21ai_1 _17999_ (.B1(_11172_),
    .Y(_01520_),
    .A1(net653),
    .A2(_11168_));
 sg13g2_nand2_1 _18000_ (.Y(_11173_),
    .A(\top_ihp.oisc.regs[3][21] ),
    .B(net640));
 sg13g2_o21ai_1 _18001_ (.B1(_11173_),
    .Y(_01521_),
    .A1(net112),
    .A2(net639));
 sg13g2_buf_8 _18002_ (.A(net322),
    .X(_11174_));
 sg13g2_nand2_1 _18003_ (.Y(_11175_),
    .A(\top_ihp.oisc.regs[3][22] ),
    .B(net640));
 sg13g2_o21ai_1 _18004_ (.B1(_11175_),
    .Y(_01522_),
    .A1(net101),
    .A2(net639));
 sg13g2_nand2_1 _18005_ (.Y(_11176_),
    .A(\top_ihp.oisc.regs[3][23] ),
    .B(net640));
 sg13g2_o21ai_1 _18006_ (.B1(_11176_),
    .Y(_01523_),
    .A1(_10987_),
    .A2(net639));
 sg13g2_nand2_1 _18007_ (.Y(_11177_),
    .A(\top_ihp.oisc.regs[3][24] ),
    .B(_11165_));
 sg13g2_o21ai_1 _18008_ (.B1(_11177_),
    .Y(_01524_),
    .A1(net111),
    .A2(_11168_));
 sg13g2_nand2_1 _18009_ (.Y(_11178_),
    .A(\top_ihp.oisc.regs[3][25] ),
    .B(net640));
 sg13g2_o21ai_1 _18010_ (.B1(_11178_),
    .Y(_01525_),
    .A1(net132),
    .A2(net639));
 sg13g2_buf_1 _18011_ (.A(net705),
    .X(_11179_));
 sg13g2_nand2_1 _18012_ (.Y(_11180_),
    .A(\top_ihp.oisc.regs[3][26] ),
    .B(net638));
 sg13g2_o21ai_1 _18013_ (.B1(_11180_),
    .Y(_01526_),
    .A1(net49),
    .A2(net639));
 sg13g2_nand2_1 _18014_ (.Y(_11181_),
    .A(\top_ihp.oisc.regs[3][27] ),
    .B(_11179_));
 sg13g2_o21ai_1 _18015_ (.B1(_11181_),
    .Y(_01527_),
    .A1(_10998_),
    .A2(net639));
 sg13g2_buf_1 _18016_ (.A(net705),
    .X(_11182_));
 sg13g2_nand2_1 _18017_ (.Y(_11183_),
    .A(\top_ihp.oisc.regs[3][28] ),
    .B(net638));
 sg13g2_o21ai_1 _18018_ (.B1(_11183_),
    .Y(_01528_),
    .A1(net284),
    .A2(net637));
 sg13g2_nand2_1 _18019_ (.Y(_11184_),
    .A(\top_ihp.oisc.regs[3][29] ),
    .B(net638));
 sg13g2_o21ai_1 _18020_ (.B1(_11184_),
    .Y(_01529_),
    .A1(net108),
    .A2(_11182_));
 sg13g2_nand2_1 _18021_ (.Y(_11185_),
    .A(\top_ihp.oisc.regs[3][2] ),
    .B(net638));
 sg13g2_o21ai_1 _18022_ (.B1(_11185_),
    .Y(_01530_),
    .A1(net43),
    .A2(net637));
 sg13g2_nand2_1 _18023_ (.Y(_11186_),
    .A(\top_ihp.oisc.regs[3][30] ),
    .B(net638));
 sg13g2_o21ai_1 _18024_ (.B1(_11186_),
    .Y(_01531_),
    .A1(_11055_),
    .A2(net637));
 sg13g2_nand2_1 _18025_ (.Y(_11187_),
    .A(\top_ihp.oisc.regs[3][31] ),
    .B(net638));
 sg13g2_o21ai_1 _18026_ (.B1(_11187_),
    .Y(_01532_),
    .A1(net315),
    .A2(net637));
 sg13g2_nand2_1 _18027_ (.Y(_11188_),
    .A(\top_ihp.oisc.regs[3][3] ),
    .B(net638));
 sg13g2_o21ai_1 _18028_ (.B1(_11188_),
    .Y(_01533_),
    .A1(_11058_),
    .A2(net637));
 sg13g2_nand2_1 _18029_ (.Y(_11189_),
    .A(\top_ihp.oisc.regs[3][4] ),
    .B(net638));
 sg13g2_o21ai_1 _18030_ (.B1(_11189_),
    .Y(_01534_),
    .A1(net40),
    .A2(net637));
 sg13g2_nand2_1 _18031_ (.Y(_11190_),
    .A(\top_ihp.oisc.regs[3][5] ),
    .B(_11179_));
 sg13g2_o21ai_1 _18032_ (.B1(_11190_),
    .Y(_01535_),
    .A1(net48),
    .A2(_11182_));
 sg13g2_nand2_1 _18033_ (.Y(_11191_),
    .A(\top_ihp.oisc.regs[3][6] ),
    .B(net705));
 sg13g2_o21ai_1 _18034_ (.B1(_11191_),
    .Y(_01536_),
    .A1(net47),
    .A2(net637));
 sg13g2_nand2_1 _18035_ (.Y(_11192_),
    .A(\top_ihp.oisc.regs[3][7] ),
    .B(net705));
 sg13g2_o21ai_1 _18036_ (.B1(_11192_),
    .Y(_01537_),
    .A1(net518),
    .A2(net637));
 sg13g2_nand2_1 _18037_ (.Y(_11193_),
    .A(\top_ihp.oisc.regs[3][8] ),
    .B(net705));
 sg13g2_o21ai_1 _18038_ (.B1(_11193_),
    .Y(_01538_),
    .A1(_11014_),
    .A2(_11154_));
 sg13g2_nand2_1 _18039_ (.Y(_11194_),
    .A(\top_ihp.oisc.regs[3][9] ),
    .B(net705));
 sg13g2_o21ai_1 _18040_ (.B1(_11194_),
    .Y(_01539_),
    .A1(net46),
    .A2(_11154_));
 sg13g2_nand3_1 _18041_ (.B(_10519_),
    .C(net708),
    .A(net766),
    .Y(_11195_));
 sg13g2_buf_1 _18042_ (.A(_11195_),
    .X(_11196_));
 sg13g2_buf_1 _18043_ (.A(_11196_),
    .X(_11197_));
 sg13g2_buf_8 _18044_ (.A(net269),
    .X(_11198_));
 sg13g2_buf_2 _18045_ (.A(_11196_),
    .X(_11199_));
 sg13g2_nand2_1 _18046_ (.Y(_11200_),
    .A(\top_ihp.oisc.regs[40][0] ),
    .B(net268));
 sg13g2_o21ai_1 _18047_ (.B1(_11200_),
    .Y(_01540_),
    .A1(net45),
    .A2(net100));
 sg13g2_nand2_1 _18048_ (.Y(_11201_),
    .A(\top_ihp.oisc.regs[40][10] ),
    .B(net268));
 sg13g2_o21ai_1 _18049_ (.B1(_11201_),
    .Y(_01541_),
    .A1(net51),
    .A2(net100));
 sg13g2_nand2_1 _18050_ (.Y(_11202_),
    .A(\top_ihp.oisc.regs[40][11] ),
    .B(net268));
 sg13g2_o21ai_1 _18051_ (.B1(_11202_),
    .Y(_01542_),
    .A1(net44),
    .A2(net100));
 sg13g2_nand2b_2 _18052_ (.Y(_11203_),
    .B(_09723_),
    .A_N(_10517_));
 sg13g2_nor2_2 _18053_ (.A(_11203_),
    .B(_10965_),
    .Y(_11204_));
 sg13g2_buf_8 _18054_ (.A(_11204_),
    .X(_11205_));
 sg13g2_nor2_1 _18055_ (.A(\top_ihp.oisc.regs[40][12] ),
    .B(net267),
    .Y(_11206_));
 sg13g2_a21oi_1 _18056_ (.A1(net153),
    .A2(net267),
    .Y(_01543_),
    .B1(_11206_));
 sg13g2_nand2_1 _18057_ (.Y(_11207_),
    .A(\top_ihp.oisc.regs[40][13] ),
    .B(net268));
 sg13g2_o21ai_1 _18058_ (.B1(_11207_),
    .Y(_01544_),
    .A1(net117),
    .A2(net100));
 sg13g2_nor2_1 _18059_ (.A(\top_ihp.oisc.regs[40][14] ),
    .B(net267),
    .Y(_11208_));
 sg13g2_a21oi_1 _18060_ (.A1(net152),
    .A2(net267),
    .Y(_01545_),
    .B1(_11208_));
 sg13g2_nor2_1 _18061_ (.A(\top_ihp.oisc.regs[40][15] ),
    .B(net267),
    .Y(_11209_));
 sg13g2_a21oi_1 _18062_ (.A1(net151),
    .A2(net267),
    .Y(_01546_),
    .B1(_11209_));
 sg13g2_nand2_1 _18063_ (.Y(_11210_),
    .A(\top_ihp.oisc.regs[40][16] ),
    .B(net268));
 sg13g2_o21ai_1 _18064_ (.B1(_11210_),
    .Y(_01547_),
    .A1(net50),
    .A2(net100));
 sg13g2_nand2_1 _18065_ (.Y(_11211_),
    .A(\top_ihp.oisc.regs[40][17] ),
    .B(_11199_));
 sg13g2_o21ai_1 _18066_ (.B1(_11211_),
    .Y(_01548_),
    .A1(net116),
    .A2(net100));
 sg13g2_nand2_1 _18067_ (.Y(_11212_),
    .A(\top_ihp.oisc.regs[40][18] ),
    .B(_11199_));
 sg13g2_o21ai_1 _18068_ (.B1(_11212_),
    .Y(_01549_),
    .A1(net115),
    .A2(net100));
 sg13g2_buf_1 _18069_ (.A(_11196_),
    .X(_11213_));
 sg13g2_nand2_1 _18070_ (.Y(_11214_),
    .A(\top_ihp.oisc.regs[40][19] ),
    .B(net266));
 sg13g2_o21ai_1 _18071_ (.B1(_11214_),
    .Y(_01550_),
    .A1(net114),
    .A2(_11198_));
 sg13g2_nor2_1 _18072_ (.A(\top_ihp.oisc.regs[40][1] ),
    .B(net267),
    .Y(_11215_));
 sg13g2_a21oi_1 _18073_ (.A1(net149),
    .A2(_11205_),
    .Y(_01551_),
    .B1(_11215_));
 sg13g2_nand2_1 _18074_ (.Y(_11216_),
    .A(\top_ihp.oisc.regs[40][20] ),
    .B(net266));
 sg13g2_o21ai_1 _18075_ (.B1(_11216_),
    .Y(_01552_),
    .A1(_10591_),
    .A2(_11198_));
 sg13g2_nand2_1 _18076_ (.Y(_11217_),
    .A(\top_ihp.oisc.regs[40][21] ),
    .B(net266));
 sg13g2_o21ai_1 _18077_ (.B1(_11217_),
    .Y(_01553_),
    .A1(net112),
    .A2(net100));
 sg13g2_nor2_1 _18078_ (.A(\top_ihp.oisc.regs[40][22] ),
    .B(_11204_),
    .Y(_11218_));
 sg13g2_a21oi_1 _18079_ (.A1(net148),
    .A2(net267),
    .Y(_01554_),
    .B1(_11218_));
 sg13g2_nand3_1 _18080_ (.B(net764),
    .C(net706),
    .A(net766),
    .Y(_11219_));
 sg13g2_buf_1 _18081_ (.A(_11219_),
    .X(_11220_));
 sg13g2_nand2_1 _18082_ (.Y(_11221_),
    .A(\top_ihp.oisc.regs[40][23] ),
    .B(net266));
 sg13g2_o21ai_1 _18083_ (.B1(_11221_),
    .Y(_01555_),
    .A1(net285),
    .A2(_11220_));
 sg13g2_buf_8 _18084_ (.A(net269),
    .X(_11222_));
 sg13g2_nand2_1 _18085_ (.Y(_11223_),
    .A(\top_ihp.oisc.regs[40][24] ),
    .B(net266));
 sg13g2_o21ai_1 _18086_ (.B1(_11223_),
    .Y(_01556_),
    .A1(net111),
    .A2(net99));
 sg13g2_nor2_1 _18087_ (.A(\top_ihp.oisc.regs[40][25] ),
    .B(_11204_),
    .Y(_11224_));
 sg13g2_a21oi_1 _18088_ (.A1(net147),
    .A2(_11205_),
    .Y(_01557_),
    .B1(_11224_));
 sg13g2_nand2_1 _18089_ (.Y(_11225_),
    .A(\top_ihp.oisc.regs[40][26] ),
    .B(net266));
 sg13g2_o21ai_1 _18090_ (.B1(_11225_),
    .Y(_01558_),
    .A1(net49),
    .A2(net99));
 sg13g2_nand2_1 _18091_ (.Y(_11226_),
    .A(\top_ihp.oisc.regs[40][27] ),
    .B(_11213_));
 sg13g2_o21ai_1 _18092_ (.B1(_11226_),
    .Y(_01559_),
    .A1(net109),
    .A2(net99));
 sg13g2_nand2_1 _18093_ (.Y(_11227_),
    .A(\top_ihp.oisc.regs[40][28] ),
    .B(net266));
 sg13g2_o21ai_1 _18094_ (.B1(_11227_),
    .Y(_01560_),
    .A1(net284),
    .A2(_11220_));
 sg13g2_nand2_1 _18095_ (.Y(_11228_),
    .A(\top_ihp.oisc.regs[40][29] ),
    .B(net266));
 sg13g2_o21ai_1 _18096_ (.B1(_11228_),
    .Y(_01561_),
    .A1(net108),
    .A2(net99));
 sg13g2_nand2_1 _18097_ (.Y(_11229_),
    .A(\top_ihp.oisc.regs[40][2] ),
    .B(_11213_));
 sg13g2_o21ai_1 _18098_ (.B1(_11229_),
    .Y(_01562_),
    .A1(net43),
    .A2(net99));
 sg13g2_nand2_1 _18099_ (.Y(_11230_),
    .A(\top_ihp.oisc.regs[40][30] ),
    .B(_11197_));
 sg13g2_o21ai_1 _18100_ (.B1(_11230_),
    .Y(_01563_),
    .A1(net42),
    .A2(net99));
 sg13g2_nand2_1 _18101_ (.Y(_11231_),
    .A(\top_ihp.oisc.regs[40][31] ),
    .B(_11220_));
 sg13g2_o21ai_1 _18102_ (.B1(_11231_),
    .Y(_01564_),
    .A1(_10606_),
    .A2(_11220_));
 sg13g2_nand2_1 _18103_ (.Y(_11232_),
    .A(\top_ihp.oisc.regs[40][3] ),
    .B(net269));
 sg13g2_o21ai_1 _18104_ (.B1(_11232_),
    .Y(_01565_),
    .A1(net41),
    .A2(_11222_));
 sg13g2_nand2_1 _18105_ (.Y(_11233_),
    .A(\top_ihp.oisc.regs[40][4] ),
    .B(net269));
 sg13g2_o21ai_1 _18106_ (.B1(_11233_),
    .Y(_01566_),
    .A1(net40),
    .A2(_11222_));
 sg13g2_nand2_1 _18107_ (.Y(_11234_),
    .A(\top_ihp.oisc.regs[40][5] ),
    .B(net269));
 sg13g2_o21ai_1 _18108_ (.B1(_11234_),
    .Y(_01567_),
    .A1(net48),
    .A2(net99));
 sg13g2_nand2_1 _18109_ (.Y(_11235_),
    .A(\top_ihp.oisc.regs[40][6] ),
    .B(_11197_));
 sg13g2_o21ai_1 _18110_ (.B1(_11235_),
    .Y(_01568_),
    .A1(net47),
    .A2(net99));
 sg13g2_nand2_1 _18111_ (.Y(_11236_),
    .A(\top_ihp.oisc.regs[40][7] ),
    .B(net269));
 sg13g2_o21ai_1 _18112_ (.B1(_11236_),
    .Y(_01569_),
    .A1(_10612_),
    .A2(net268));
 sg13g2_nand2_1 _18113_ (.Y(_11237_),
    .A(\top_ihp.oisc.regs[40][8] ),
    .B(net269));
 sg13g2_o21ai_1 _18114_ (.B1(_11237_),
    .Y(_01570_),
    .A1(net107),
    .A2(net268));
 sg13g2_nand2_1 _18115_ (.Y(_11238_),
    .A(\top_ihp.oisc.regs[40][9] ),
    .B(net269));
 sg13g2_o21ai_1 _18116_ (.B1(_11238_),
    .Y(_01571_),
    .A1(net46),
    .A2(net268));
 sg13g2_nand3_1 _18117_ (.B(net784),
    .C(_10881_),
    .A(net764),
    .Y(_11239_));
 sg13g2_buf_2 _18118_ (.A(_11239_),
    .X(_11240_));
 sg13g2_buf_1 _18119_ (.A(_11240_),
    .X(_11241_));
 sg13g2_nand3_1 _18120_ (.B(net784),
    .C(net707),
    .A(net764),
    .Y(_11242_));
 sg13g2_buf_2 _18121_ (.A(_11242_),
    .X(_11243_));
 sg13g2_buf_1 _18122_ (.A(_11243_),
    .X(_11244_));
 sg13g2_nand2_1 _18123_ (.Y(_11245_),
    .A(\top_ihp.oisc.regs[41][0] ),
    .B(net264));
 sg13g2_o21ai_1 _18124_ (.B1(_11245_),
    .Y(_01572_),
    .A1(net45),
    .A2(net265));
 sg13g2_nand2_1 _18125_ (.Y(_11246_),
    .A(\top_ihp.oisc.regs[41][10] ),
    .B(net264));
 sg13g2_o21ai_1 _18126_ (.B1(_11246_),
    .Y(_01573_),
    .A1(net51),
    .A2(net265));
 sg13g2_nand2_1 _18127_ (.Y(_11247_),
    .A(\top_ihp.oisc.regs[41][11] ),
    .B(net264));
 sg13g2_o21ai_1 _18128_ (.B1(_11247_),
    .Y(_01574_),
    .A1(net44),
    .A2(net265));
 sg13g2_nor2_1 _18129_ (.A(_11203_),
    .B(_11029_),
    .Y(_11248_));
 sg13g2_buf_1 _18130_ (.A(_11248_),
    .X(_11249_));
 sg13g2_nor2_1 _18131_ (.A(\top_ihp.oisc.regs[41][12] ),
    .B(net263),
    .Y(_11250_));
 sg13g2_a21oi_1 _18132_ (.A1(net153),
    .A2(net263),
    .Y(_01575_),
    .B1(_11250_));
 sg13g2_nand2_1 _18133_ (.Y(_11251_),
    .A(\top_ihp.oisc.regs[41][13] ),
    .B(net264));
 sg13g2_o21ai_1 _18134_ (.B1(_11251_),
    .Y(_01576_),
    .A1(net117),
    .A2(net265));
 sg13g2_nor2_1 _18135_ (.A(\top_ihp.oisc.regs[41][14] ),
    .B(net263),
    .Y(_11252_));
 sg13g2_a21oi_1 _18136_ (.A1(net152),
    .A2(net263),
    .Y(_01577_),
    .B1(_11252_));
 sg13g2_nor2_1 _18137_ (.A(\top_ihp.oisc.regs[41][15] ),
    .B(net263),
    .Y(_11253_));
 sg13g2_a21oi_1 _18138_ (.A1(net151),
    .A2(net263),
    .Y(_01578_),
    .B1(_11253_));
 sg13g2_nand2_1 _18139_ (.Y(_11254_),
    .A(\top_ihp.oisc.regs[41][16] ),
    .B(net264));
 sg13g2_o21ai_1 _18140_ (.B1(_11254_),
    .Y(_01579_),
    .A1(net50),
    .A2(net265));
 sg13g2_nand2_1 _18141_ (.Y(_02838_),
    .A(\top_ihp.oisc.regs[41][17] ),
    .B(net264));
 sg13g2_o21ai_1 _18142_ (.B1(_02838_),
    .Y(_01580_),
    .A1(net116),
    .A2(_11241_));
 sg13g2_nand2_1 _18143_ (.Y(_02839_),
    .A(\top_ihp.oisc.regs[41][18] ),
    .B(net264));
 sg13g2_o21ai_1 _18144_ (.B1(_02839_),
    .Y(_01581_),
    .A1(net115),
    .A2(net265));
 sg13g2_nand2_1 _18145_ (.Y(_02840_),
    .A(\top_ihp.oisc.regs[41][19] ),
    .B(net264));
 sg13g2_o21ai_1 _18146_ (.B1(_02840_),
    .Y(_01582_),
    .A1(net114),
    .A2(_11241_));
 sg13g2_nor2_1 _18147_ (.A(\top_ihp.oisc.regs[41][1] ),
    .B(_11249_),
    .Y(_02841_));
 sg13g2_a21oi_1 _18148_ (.A1(net149),
    .A2(_11249_),
    .Y(_01583_),
    .B1(_02841_));
 sg13g2_buf_1 _18149_ (.A(_10144_),
    .X(_02842_));
 sg13g2_buf_1 _18150_ (.A(_11243_),
    .X(_02843_));
 sg13g2_nand2_1 _18151_ (.Y(_02844_),
    .A(\top_ihp.oisc.regs[41][20] ),
    .B(net262));
 sg13g2_o21ai_1 _18152_ (.B1(_02844_),
    .Y(_01584_),
    .A1(net636),
    .A2(_11244_));
 sg13g2_nand2_1 _18153_ (.Y(_02845_),
    .A(\top_ihp.oisc.regs[41][21] ),
    .B(net262));
 sg13g2_o21ai_1 _18154_ (.B1(_02845_),
    .Y(_01585_),
    .A1(net112),
    .A2(net265));
 sg13g2_nor2_1 _18155_ (.A(\top_ihp.oisc.regs[41][22] ),
    .B(_11248_),
    .Y(_02846_));
 sg13g2_a21oi_1 _18156_ (.A1(net148),
    .A2(net263),
    .Y(_01586_),
    .B1(_02846_));
 sg13g2_nand2_1 _18157_ (.Y(_02847_),
    .A(\top_ihp.oisc.regs[41][23] ),
    .B(_11240_));
 sg13g2_o21ai_1 _18158_ (.B1(_02847_),
    .Y(_01587_),
    .A1(net285),
    .A2(net265));
 sg13g2_buf_1 _18159_ (.A(_11240_),
    .X(_02848_));
 sg13g2_nand2_1 _18160_ (.Y(_02849_),
    .A(\top_ihp.oisc.regs[41][24] ),
    .B(net262));
 sg13g2_o21ai_1 _18161_ (.B1(_02849_),
    .Y(_01588_),
    .A1(net111),
    .A2(net261));
 sg13g2_nor2_1 _18162_ (.A(\top_ihp.oisc.regs[41][25] ),
    .B(_11248_),
    .Y(_02850_));
 sg13g2_a21oi_1 _18163_ (.A1(net147),
    .A2(net263),
    .Y(_01589_),
    .B1(_02850_));
 sg13g2_nand2_1 _18164_ (.Y(_02851_),
    .A(\top_ihp.oisc.regs[41][26] ),
    .B(net262));
 sg13g2_o21ai_1 _18165_ (.B1(_02851_),
    .Y(_01590_),
    .A1(net49),
    .A2(net261));
 sg13g2_nand2_1 _18166_ (.Y(_02852_),
    .A(\top_ihp.oisc.regs[41][27] ),
    .B(_02843_));
 sg13g2_o21ai_1 _18167_ (.B1(_02852_),
    .Y(_01591_),
    .A1(net109),
    .A2(_02848_));
 sg13g2_nand2_1 _18168_ (.Y(_02853_),
    .A(\top_ihp.oisc.regs[41][28] ),
    .B(_02843_));
 sg13g2_o21ai_1 _18169_ (.B1(_02853_),
    .Y(_01592_),
    .A1(net284),
    .A2(net261));
 sg13g2_nand2_1 _18170_ (.Y(_02854_),
    .A(\top_ihp.oisc.regs[41][29] ),
    .B(net262));
 sg13g2_o21ai_1 _18171_ (.B1(_02854_),
    .Y(_01593_),
    .A1(net108),
    .A2(net261));
 sg13g2_nand2_1 _18172_ (.Y(_02855_),
    .A(\top_ihp.oisc.regs[41][2] ),
    .B(net262));
 sg13g2_o21ai_1 _18173_ (.B1(_02855_),
    .Y(_01594_),
    .A1(net43),
    .A2(net261));
 sg13g2_nand2_1 _18174_ (.Y(_02856_),
    .A(\top_ihp.oisc.regs[41][30] ),
    .B(net262));
 sg13g2_o21ai_1 _18175_ (.B1(_02856_),
    .Y(_01595_),
    .A1(net42),
    .A2(net261));
 sg13g2_nand2_1 _18176_ (.Y(_02857_),
    .A(\top_ihp.oisc.regs[41][31] ),
    .B(_11240_));
 sg13g2_o21ai_1 _18177_ (.B1(_02857_),
    .Y(_01596_),
    .A1(_10606_),
    .A2(net261));
 sg13g2_nand2_1 _18178_ (.Y(_02858_),
    .A(\top_ihp.oisc.regs[41][3] ),
    .B(net262));
 sg13g2_o21ai_1 _18179_ (.B1(_02858_),
    .Y(_01597_),
    .A1(_11058_),
    .A2(net261));
 sg13g2_nand2_1 _18180_ (.Y(_02859_),
    .A(\top_ihp.oisc.regs[41][4] ),
    .B(_11243_));
 sg13g2_o21ai_1 _18181_ (.B1(_02859_),
    .Y(_01598_),
    .A1(net40),
    .A2(_02848_));
 sg13g2_nand2_1 _18182_ (.Y(_02860_),
    .A(\top_ihp.oisc.regs[41][5] ),
    .B(_11243_));
 sg13g2_o21ai_1 _18183_ (.B1(_02860_),
    .Y(_01599_),
    .A1(net48),
    .A2(_11240_));
 sg13g2_nand2_1 _18184_ (.Y(_02861_),
    .A(\top_ihp.oisc.regs[41][6] ),
    .B(_11243_));
 sg13g2_o21ai_1 _18185_ (.B1(_02861_),
    .Y(_01600_),
    .A1(_11011_),
    .A2(_11240_));
 sg13g2_buf_2 _18186_ (.A(_10480_),
    .X(_02862_));
 sg13g2_nand2_1 _18187_ (.Y(_02863_),
    .A(\top_ihp.oisc.regs[41][7] ),
    .B(_11243_));
 sg13g2_o21ai_1 _18188_ (.B1(_02863_),
    .Y(_01601_),
    .A1(net501),
    .A2(_11244_));
 sg13g2_nand2_1 _18189_ (.Y(_02864_),
    .A(\top_ihp.oisc.regs[41][8] ),
    .B(_11243_));
 sg13g2_o21ai_1 _18190_ (.B1(_02864_),
    .Y(_01602_),
    .A1(net107),
    .A2(_11240_));
 sg13g2_nand2_1 _18191_ (.Y(_02865_),
    .A(\top_ihp.oisc.regs[41][9] ),
    .B(_11243_));
 sg13g2_o21ai_1 _18192_ (.B1(_02865_),
    .Y(_01603_),
    .A1(net46),
    .A2(_11240_));
 sg13g2_nand3_1 _18193_ (.B(net741),
    .C(net708),
    .A(_10519_),
    .Y(_02866_));
 sg13g2_buf_1 _18194_ (.A(_02866_),
    .X(_02867_));
 sg13g2_buf_1 _18195_ (.A(net500),
    .X(_02868_));
 sg13g2_buf_1 _18196_ (.A(net500),
    .X(_02869_));
 sg13g2_nand2_1 _18197_ (.Y(_02870_),
    .A(\top_ihp.oisc.regs[42][0] ),
    .B(net259));
 sg13g2_o21ai_1 _18198_ (.B1(_02870_),
    .Y(_01604_),
    .A1(net45),
    .A2(net260));
 sg13g2_nand2_1 _18199_ (.Y(_02871_),
    .A(\top_ihp.oisc.regs[42][10] ),
    .B(net259));
 sg13g2_o21ai_1 _18200_ (.B1(_02871_),
    .Y(_01605_),
    .A1(net51),
    .A2(net260));
 sg13g2_nand2_1 _18201_ (.Y(_02872_),
    .A(\top_ihp.oisc.regs[42][11] ),
    .B(net259));
 sg13g2_o21ai_1 _18202_ (.B1(_02872_),
    .Y(_01606_),
    .A1(net44),
    .A2(net260));
 sg13g2_nand3_1 _18203_ (.B(net741),
    .C(net706),
    .A(net764),
    .Y(_02873_));
 sg13g2_buf_8 _18204_ (.A(_02873_),
    .X(_02874_));
 sg13g2_buf_8 _18205_ (.A(net499),
    .X(_02875_));
 sg13g2_nand2_1 _18206_ (.Y(_02876_),
    .A(\top_ihp.oisc.regs[42][12] ),
    .B(net499));
 sg13g2_o21ai_1 _18207_ (.B1(_02876_),
    .Y(_01607_),
    .A1(net104),
    .A2(net258));
 sg13g2_nand2_1 _18208_ (.Y(_02877_),
    .A(\top_ihp.oisc.regs[42][13] ),
    .B(net259));
 sg13g2_o21ai_1 _18209_ (.B1(_02877_),
    .Y(_01608_),
    .A1(net117),
    .A2(net260));
 sg13g2_nand2_1 _18210_ (.Y(_02878_),
    .A(\top_ihp.oisc.regs[42][14] ),
    .B(net499));
 sg13g2_o21ai_1 _18211_ (.B1(_02878_),
    .Y(_01609_),
    .A1(_11161_),
    .A2(net258));
 sg13g2_buf_8 _18212_ (.A(net329),
    .X(_02879_));
 sg13g2_nand2_1 _18213_ (.Y(_02880_),
    .A(\top_ihp.oisc.regs[42][15] ),
    .B(net499));
 sg13g2_o21ai_1 _18214_ (.B1(_02880_),
    .Y(_01610_),
    .A1(net98),
    .A2(net258));
 sg13g2_nand2_1 _18215_ (.Y(_02881_),
    .A(\top_ihp.oisc.regs[42][16] ),
    .B(net259));
 sg13g2_o21ai_1 _18216_ (.B1(_02881_),
    .Y(_01611_),
    .A1(net50),
    .A2(net260));
 sg13g2_nand2_1 _18217_ (.Y(_02882_),
    .A(\top_ihp.oisc.regs[42][17] ),
    .B(net259));
 sg13g2_o21ai_1 _18218_ (.B1(_02882_),
    .Y(_01612_),
    .A1(net116),
    .A2(net260));
 sg13g2_nand2_1 _18219_ (.Y(_02883_),
    .A(\top_ihp.oisc.regs[42][18] ),
    .B(net259));
 sg13g2_o21ai_1 _18220_ (.B1(_02883_),
    .Y(_01613_),
    .A1(net115),
    .A2(net260));
 sg13g2_nand2_1 _18221_ (.Y(_02884_),
    .A(\top_ihp.oisc.regs[42][19] ),
    .B(net259));
 sg13g2_o21ai_1 _18222_ (.B1(_02884_),
    .Y(_01614_),
    .A1(net114),
    .A2(net260));
 sg13g2_nand2_1 _18223_ (.Y(_02885_),
    .A(\top_ihp.oisc.regs[42][1] ),
    .B(net499));
 sg13g2_o21ai_1 _18224_ (.B1(_02885_),
    .Y(_01615_),
    .A1(net102),
    .A2(net258));
 sg13g2_nand2_1 _18225_ (.Y(_02886_),
    .A(\top_ihp.oisc.regs[42][20] ),
    .B(_02869_));
 sg13g2_o21ai_1 _18226_ (.B1(_02886_),
    .Y(_01616_),
    .A1(net324),
    .A2(_02875_));
 sg13g2_buf_1 _18227_ (.A(net500),
    .X(_02887_));
 sg13g2_nand2_1 _18228_ (.Y(_02888_),
    .A(\top_ihp.oisc.regs[42][21] ),
    .B(net257));
 sg13g2_o21ai_1 _18229_ (.B1(_02888_),
    .Y(_01617_),
    .A1(net112),
    .A2(_02868_));
 sg13g2_nand2_1 _18230_ (.Y(_02889_),
    .A(\top_ihp.oisc.regs[42][22] ),
    .B(net499));
 sg13g2_o21ai_1 _18231_ (.B1(_02889_),
    .Y(_01618_),
    .A1(net101),
    .A2(net258));
 sg13g2_nand2_1 _18232_ (.Y(_02890_),
    .A(\top_ihp.oisc.regs[42][23] ),
    .B(_02874_));
 sg13g2_o21ai_1 _18233_ (.B1(_02890_),
    .Y(_01619_),
    .A1(net285),
    .A2(_02875_));
 sg13g2_nand2_1 _18234_ (.Y(_02891_),
    .A(\top_ihp.oisc.regs[42][24] ),
    .B(net257));
 sg13g2_o21ai_1 _18235_ (.B1(_02891_),
    .Y(_01620_),
    .A1(net111),
    .A2(_02868_));
 sg13g2_buf_1 _18236_ (.A(net319),
    .X(_02892_));
 sg13g2_nand2_1 _18237_ (.Y(_02893_),
    .A(\top_ihp.oisc.regs[42][25] ),
    .B(net499));
 sg13g2_o21ai_1 _18238_ (.B1(_02893_),
    .Y(_01621_),
    .A1(net97),
    .A2(net258));
 sg13g2_buf_1 _18239_ (.A(net500),
    .X(_02894_));
 sg13g2_nand2_1 _18240_ (.Y(_02895_),
    .A(\top_ihp.oisc.regs[42][26] ),
    .B(net257));
 sg13g2_o21ai_1 _18241_ (.B1(_02895_),
    .Y(_01622_),
    .A1(net49),
    .A2(net256));
 sg13g2_nand2_1 _18242_ (.Y(_02896_),
    .A(\top_ihp.oisc.regs[42][27] ),
    .B(net257));
 sg13g2_o21ai_1 _18243_ (.B1(_02896_),
    .Y(_01623_),
    .A1(net109),
    .A2(net256));
 sg13g2_nand2_1 _18244_ (.Y(_02897_),
    .A(\top_ihp.oisc.regs[42][28] ),
    .B(net257));
 sg13g2_o21ai_1 _18245_ (.B1(_02897_),
    .Y(_01624_),
    .A1(net284),
    .A2(net258));
 sg13g2_nand2_1 _18246_ (.Y(_02898_),
    .A(\top_ihp.oisc.regs[42][29] ),
    .B(net257));
 sg13g2_o21ai_1 _18247_ (.B1(_02898_),
    .Y(_01625_),
    .A1(net108),
    .A2(net256));
 sg13g2_nand2_1 _18248_ (.Y(_02899_),
    .A(\top_ihp.oisc.regs[42][2] ),
    .B(net257));
 sg13g2_o21ai_1 _18249_ (.B1(_02899_),
    .Y(_01626_),
    .A1(net43),
    .A2(_02894_));
 sg13g2_nand2_1 _18250_ (.Y(_02900_),
    .A(\top_ihp.oisc.regs[42][30] ),
    .B(net257));
 sg13g2_o21ai_1 _18251_ (.B1(_02900_),
    .Y(_01627_),
    .A1(net42),
    .A2(net256));
 sg13g2_nand2_1 _18252_ (.Y(_02901_),
    .A(\top_ihp.oisc.regs[42][31] ),
    .B(net499));
 sg13g2_o21ai_1 _18253_ (.B1(_02901_),
    .Y(_01628_),
    .A1(net52),
    .A2(net258));
 sg13g2_nand2_1 _18254_ (.Y(_02902_),
    .A(\top_ihp.oisc.regs[42][3] ),
    .B(_02887_));
 sg13g2_o21ai_1 _18255_ (.B1(_02902_),
    .Y(_01629_),
    .A1(net41),
    .A2(_02894_));
 sg13g2_nand2_1 _18256_ (.Y(_02903_),
    .A(\top_ihp.oisc.regs[42][4] ),
    .B(_02887_));
 sg13g2_o21ai_1 _18257_ (.B1(_02903_),
    .Y(_01630_),
    .A1(net40),
    .A2(net256));
 sg13g2_nand2_1 _18258_ (.Y(_02904_),
    .A(\top_ihp.oisc.regs[42][5] ),
    .B(_02867_));
 sg13g2_o21ai_1 _18259_ (.B1(_02904_),
    .Y(_01631_),
    .A1(net48),
    .A2(net256));
 sg13g2_nand2_1 _18260_ (.Y(_02905_),
    .A(\top_ihp.oisc.regs[42][6] ),
    .B(net500));
 sg13g2_o21ai_1 _18261_ (.B1(_02905_),
    .Y(_01632_),
    .A1(_11011_),
    .A2(net256));
 sg13g2_nand2_1 _18262_ (.Y(_02906_),
    .A(\top_ihp.oisc.regs[42][7] ),
    .B(net500));
 sg13g2_o21ai_1 _18263_ (.B1(_02906_),
    .Y(_01633_),
    .A1(_10484_),
    .A2(_02874_));
 sg13g2_nand2_1 _18264_ (.Y(_02907_),
    .A(\top_ihp.oisc.regs[42][8] ),
    .B(net500));
 sg13g2_o21ai_1 _18265_ (.B1(_02907_),
    .Y(_01634_),
    .A1(net107),
    .A2(net256));
 sg13g2_nand2_1 _18266_ (.Y(_02908_),
    .A(\top_ihp.oisc.regs[42][9] ),
    .B(net500));
 sg13g2_o21ai_1 _18267_ (.B1(_02908_),
    .Y(_01635_),
    .A1(_11016_),
    .A2(_02869_));
 sg13g2_nand3_1 _18268_ (.B(net785),
    .C(net708),
    .A(_10519_),
    .Y(_02909_));
 sg13g2_buf_1 _18269_ (.A(_02909_),
    .X(_02910_));
 sg13g2_buf_1 _18270_ (.A(_02910_),
    .X(_02911_));
 sg13g2_buf_1 _18271_ (.A(net255),
    .X(_02912_));
 sg13g2_nand3_1 _18272_ (.B(net785),
    .C(net707),
    .A(_10519_),
    .Y(_02913_));
 sg13g2_buf_2 _18273_ (.A(_02913_),
    .X(_02914_));
 sg13g2_buf_1 _18274_ (.A(_02914_),
    .X(_02915_));
 sg13g2_nand2_1 _18275_ (.Y(_02916_),
    .A(\top_ihp.oisc.regs[43][0] ),
    .B(net254));
 sg13g2_o21ai_1 _18276_ (.B1(_02916_),
    .Y(_01636_),
    .A1(net45),
    .A2(net96));
 sg13g2_nand2_1 _18277_ (.Y(_02917_),
    .A(\top_ihp.oisc.regs[43][10] ),
    .B(net254));
 sg13g2_o21ai_1 _18278_ (.B1(_02917_),
    .Y(_01637_),
    .A1(net51),
    .A2(net96));
 sg13g2_nand2_1 _18279_ (.Y(_02918_),
    .A(\top_ihp.oisc.regs[43][11] ),
    .B(net254));
 sg13g2_o21ai_1 _18280_ (.B1(_02918_),
    .Y(_01638_),
    .A1(net44),
    .A2(net96));
 sg13g2_nand2_1 _18281_ (.Y(_02919_),
    .A(\top_ihp.oisc.regs[43][12] ),
    .B(net255));
 sg13g2_o21ai_1 _18282_ (.B1(_02919_),
    .Y(_01639_),
    .A1(net104),
    .A2(net96));
 sg13g2_nand2_1 _18283_ (.Y(_02920_),
    .A(\top_ihp.oisc.regs[43][13] ),
    .B(_02915_));
 sg13g2_o21ai_1 _18284_ (.B1(_02920_),
    .Y(_01640_),
    .A1(net117),
    .A2(net96));
 sg13g2_nand2_1 _18285_ (.Y(_02921_),
    .A(\top_ihp.oisc.regs[43][14] ),
    .B(net255));
 sg13g2_o21ai_1 _18286_ (.B1(_02921_),
    .Y(_01641_),
    .A1(net103),
    .A2(net96));
 sg13g2_nand2_1 _18287_ (.Y(_02922_),
    .A(\top_ihp.oisc.regs[43][15] ),
    .B(net255));
 sg13g2_o21ai_1 _18288_ (.B1(_02922_),
    .Y(_01642_),
    .A1(net98),
    .A2(net96));
 sg13g2_nand2_1 _18289_ (.Y(_02923_),
    .A(\top_ihp.oisc.regs[43][16] ),
    .B(_02915_));
 sg13g2_o21ai_1 _18290_ (.B1(_02923_),
    .Y(_01643_),
    .A1(_10973_),
    .A2(net96));
 sg13g2_nand2_1 _18291_ (.Y(_02924_),
    .A(\top_ihp.oisc.regs[43][17] ),
    .B(net254));
 sg13g2_o21ai_1 _18292_ (.B1(_02924_),
    .Y(_01644_),
    .A1(_10975_),
    .A2(_02912_));
 sg13g2_nand2_1 _18293_ (.Y(_02925_),
    .A(\top_ihp.oisc.regs[43][18] ),
    .B(net254));
 sg13g2_o21ai_1 _18294_ (.B1(_02925_),
    .Y(_01645_),
    .A1(net115),
    .A2(_02912_));
 sg13g2_buf_1 _18295_ (.A(_02911_),
    .X(_02926_));
 sg13g2_nand2_1 _18296_ (.Y(_02927_),
    .A(\top_ihp.oisc.regs[43][19] ),
    .B(net254));
 sg13g2_o21ai_1 _18297_ (.B1(_02927_),
    .Y(_01646_),
    .A1(net114),
    .A2(net95));
 sg13g2_nand2_1 _18298_ (.Y(_02928_),
    .A(\top_ihp.oisc.regs[43][1] ),
    .B(_02911_));
 sg13g2_o21ai_1 _18299_ (.B1(_02928_),
    .Y(_01647_),
    .A1(net102),
    .A2(_02926_));
 sg13g2_buf_1 _18300_ (.A(_02914_),
    .X(_02929_));
 sg13g2_nand2_1 _18301_ (.Y(_02930_),
    .A(\top_ihp.oisc.regs[43][20] ),
    .B(net253));
 sg13g2_o21ai_1 _18302_ (.B1(_02930_),
    .Y(_01648_),
    .A1(net636),
    .A2(net254));
 sg13g2_nand2_1 _18303_ (.Y(_02931_),
    .A(\top_ihp.oisc.regs[43][21] ),
    .B(net253));
 sg13g2_o21ai_1 _18304_ (.B1(_02931_),
    .Y(_01649_),
    .A1(_10984_),
    .A2(net95));
 sg13g2_nand2_1 _18305_ (.Y(_02932_),
    .A(\top_ihp.oisc.regs[43][22] ),
    .B(net255));
 sg13g2_o21ai_1 _18306_ (.B1(_02932_),
    .Y(_01650_),
    .A1(net101),
    .A2(net95));
 sg13g2_nand2_1 _18307_ (.Y(_02933_),
    .A(\top_ihp.oisc.regs[43][23] ),
    .B(net255));
 sg13g2_o21ai_1 _18308_ (.B1(_02933_),
    .Y(_01651_),
    .A1(_10987_),
    .A2(_02926_));
 sg13g2_nand2_1 _18309_ (.Y(_02934_),
    .A(\top_ihp.oisc.regs[43][24] ),
    .B(net253));
 sg13g2_o21ai_1 _18310_ (.B1(_02934_),
    .Y(_01652_),
    .A1(_10992_),
    .A2(net95));
 sg13g2_nand2_1 _18311_ (.Y(_02935_),
    .A(\top_ihp.oisc.regs[43][25] ),
    .B(net255));
 sg13g2_o21ai_1 _18312_ (.B1(_02935_),
    .Y(_01653_),
    .A1(net97),
    .A2(net95));
 sg13g2_nand2_1 _18313_ (.Y(_02936_),
    .A(\top_ihp.oisc.regs[43][26] ),
    .B(net253));
 sg13g2_o21ai_1 _18314_ (.B1(_02936_),
    .Y(_01654_),
    .A1(net49),
    .A2(net95));
 sg13g2_nand2_1 _18315_ (.Y(_02937_),
    .A(\top_ihp.oisc.regs[43][27] ),
    .B(_02929_));
 sg13g2_o21ai_1 _18316_ (.B1(_02937_),
    .Y(_01655_),
    .A1(net109),
    .A2(net95));
 sg13g2_nand2_1 _18317_ (.Y(_02938_),
    .A(\top_ihp.oisc.regs[43][28] ),
    .B(net253));
 sg13g2_o21ai_1 _18318_ (.B1(_02938_),
    .Y(_01656_),
    .A1(net284),
    .A2(net95));
 sg13g2_buf_2 _18319_ (.A(_02910_),
    .X(_02939_));
 sg13g2_nand2_1 _18320_ (.Y(_02940_),
    .A(\top_ihp.oisc.regs[43][29] ),
    .B(net253));
 sg13g2_o21ai_1 _18321_ (.B1(_02940_),
    .Y(_01657_),
    .A1(_11002_),
    .A2(net252));
 sg13g2_nand2_1 _18322_ (.Y(_02941_),
    .A(\top_ihp.oisc.regs[43][2] ),
    .B(net253));
 sg13g2_o21ai_1 _18323_ (.B1(_02941_),
    .Y(_01658_),
    .A1(_11053_),
    .A2(net252));
 sg13g2_nand2_1 _18324_ (.Y(_02942_),
    .A(\top_ihp.oisc.regs[43][30] ),
    .B(net253));
 sg13g2_o21ai_1 _18325_ (.B1(_02942_),
    .Y(_01659_),
    .A1(net42),
    .A2(net252));
 sg13g2_buf_1 _18326_ (.A(_10345_),
    .X(_02943_));
 sg13g2_nand2_1 _18327_ (.Y(_02944_),
    .A(\top_ihp.oisc.regs[43][31] ),
    .B(net255));
 sg13g2_o21ai_1 _18328_ (.B1(_02944_),
    .Y(_01660_),
    .A1(net251),
    .A2(net252));
 sg13g2_nand2_1 _18329_ (.Y(_02945_),
    .A(\top_ihp.oisc.regs[43][3] ),
    .B(_02929_));
 sg13g2_o21ai_1 _18330_ (.B1(_02945_),
    .Y(_01661_),
    .A1(net41),
    .A2(_02939_));
 sg13g2_nand2_1 _18331_ (.Y(_02946_),
    .A(\top_ihp.oisc.regs[43][4] ),
    .B(_02914_));
 sg13g2_o21ai_1 _18332_ (.B1(_02946_),
    .Y(_01662_),
    .A1(net40),
    .A2(net252));
 sg13g2_nand2_1 _18333_ (.Y(_02947_),
    .A(\top_ihp.oisc.regs[43][5] ),
    .B(_02914_));
 sg13g2_o21ai_1 _18334_ (.B1(_02947_),
    .Y(_01663_),
    .A1(net48),
    .A2(_02939_));
 sg13g2_nand2_1 _18335_ (.Y(_02948_),
    .A(\top_ihp.oisc.regs[43][6] ),
    .B(_02914_));
 sg13g2_o21ai_1 _18336_ (.B1(_02948_),
    .Y(_01664_),
    .A1(net47),
    .A2(net252));
 sg13g2_nand2_1 _18337_ (.Y(_02949_),
    .A(\top_ihp.oisc.regs[43][7] ),
    .B(_02914_));
 sg13g2_o21ai_1 _18338_ (.B1(_02949_),
    .Y(_01665_),
    .A1(net501),
    .A2(net254));
 sg13g2_nand2_1 _18339_ (.Y(_02950_),
    .A(\top_ihp.oisc.regs[43][8] ),
    .B(_02914_));
 sg13g2_o21ai_1 _18340_ (.B1(_02950_),
    .Y(_01666_),
    .A1(_11014_),
    .A2(net252));
 sg13g2_nand2_1 _18341_ (.Y(_02951_),
    .A(\top_ihp.oisc.regs[43][9] ),
    .B(_02914_));
 sg13g2_o21ai_1 _18342_ (.B1(_02951_),
    .Y(_01667_),
    .A1(_11016_),
    .A2(net252));
 sg13g2_nand3_1 _18343_ (.B(_10618_),
    .C(_10826_),
    .A(net766),
    .Y(_02952_));
 sg13g2_buf_1 _18344_ (.A(_02952_),
    .X(_02953_));
 sg13g2_buf_2 _18345_ (.A(_02953_),
    .X(_02954_));
 sg13g2_buf_8 _18346_ (.A(net250),
    .X(_02955_));
 sg13g2_buf_2 _18347_ (.A(_02953_),
    .X(_02956_));
 sg13g2_nand2_1 _18348_ (.Y(_02957_),
    .A(\top_ihp.oisc.regs[44][0] ),
    .B(net249));
 sg13g2_o21ai_1 _18349_ (.B1(_02957_),
    .Y(_01668_),
    .A1(net45),
    .A2(net94));
 sg13g2_nand2_1 _18350_ (.Y(_02958_),
    .A(\top_ihp.oisc.regs[44][10] ),
    .B(net249));
 sg13g2_o21ai_1 _18351_ (.B1(_02958_),
    .Y(_01669_),
    .A1(net51),
    .A2(net94));
 sg13g2_nand2_1 _18352_ (.Y(_02959_),
    .A(\top_ihp.oisc.regs[44][11] ),
    .B(net249));
 sg13g2_o21ai_1 _18353_ (.B1(_02959_),
    .Y(_01670_),
    .A1(net44),
    .A2(net94));
 sg13g2_nand4_1 _18354_ (.B(_09723_),
    .C(_09714_),
    .A(_09532_),
    .Y(_02960_),
    .D(_09720_));
 sg13g2_buf_2 _18355_ (.A(_02960_),
    .X(_02961_));
 sg13g2_nor2_2 _18356_ (.A(_02961_),
    .B(_10965_),
    .Y(_02962_));
 sg13g2_buf_8 _18357_ (.A(_02962_),
    .X(_02963_));
 sg13g2_nor2_1 _18358_ (.A(\top_ihp.oisc.regs[44][12] ),
    .B(net248),
    .Y(_02964_));
 sg13g2_a21oi_1 _18359_ (.A1(_09906_),
    .A2(net248),
    .Y(_01671_),
    .B1(_02964_));
 sg13g2_nand2_1 _18360_ (.Y(_02965_),
    .A(\top_ihp.oisc.regs[44][13] ),
    .B(net249));
 sg13g2_o21ai_1 _18361_ (.B1(_02965_),
    .Y(_01672_),
    .A1(_10969_),
    .A2(net94));
 sg13g2_nor2_1 _18362_ (.A(\top_ihp.oisc.regs[44][14] ),
    .B(net248),
    .Y(_02966_));
 sg13g2_a21oi_1 _18363_ (.A1(net152),
    .A2(net248),
    .Y(_01673_),
    .B1(_02966_));
 sg13g2_nor2_1 _18364_ (.A(\top_ihp.oisc.regs[44][15] ),
    .B(net248),
    .Y(_02967_));
 sg13g2_a21oi_1 _18365_ (.A1(net151),
    .A2(net248),
    .Y(_01674_),
    .B1(_02967_));
 sg13g2_nand2_1 _18366_ (.Y(_02968_),
    .A(\top_ihp.oisc.regs[44][16] ),
    .B(net249));
 sg13g2_o21ai_1 _18367_ (.B1(_02968_),
    .Y(_01675_),
    .A1(_10973_),
    .A2(net94));
 sg13g2_nand2_1 _18368_ (.Y(_02969_),
    .A(\top_ihp.oisc.regs[44][17] ),
    .B(_02956_));
 sg13g2_o21ai_1 _18369_ (.B1(_02969_),
    .Y(_01676_),
    .A1(_10975_),
    .A2(net94));
 sg13g2_nand2_1 _18370_ (.Y(_02970_),
    .A(\top_ihp.oisc.regs[44][18] ),
    .B(_02956_));
 sg13g2_o21ai_1 _18371_ (.B1(_02970_),
    .Y(_01677_),
    .A1(net115),
    .A2(_02955_));
 sg13g2_buf_8 _18372_ (.A(net250),
    .X(_02971_));
 sg13g2_nand2_1 _18373_ (.Y(_02972_),
    .A(\top_ihp.oisc.regs[44][19] ),
    .B(net93));
 sg13g2_o21ai_1 _18374_ (.B1(_02972_),
    .Y(_01678_),
    .A1(net114),
    .A2(_02955_));
 sg13g2_nor2_1 _18375_ (.A(\top_ihp.oisc.regs[44][1] ),
    .B(net248),
    .Y(_02973_));
 sg13g2_a21oi_1 _18376_ (.A1(net149),
    .A2(net248),
    .Y(_01679_),
    .B1(_02973_));
 sg13g2_nand2_1 _18377_ (.Y(_02974_),
    .A(\top_ihp.oisc.regs[44][20] ),
    .B(net93));
 sg13g2_o21ai_1 _18378_ (.B1(_02974_),
    .Y(_01680_),
    .A1(net636),
    .A2(net94));
 sg13g2_nand2_1 _18379_ (.Y(_02975_),
    .A(\top_ihp.oisc.regs[44][21] ),
    .B(net93));
 sg13g2_o21ai_1 _18380_ (.B1(_02975_),
    .Y(_01681_),
    .A1(_10984_),
    .A2(net94));
 sg13g2_nor2_1 _18381_ (.A(\top_ihp.oisc.regs[44][22] ),
    .B(_02962_),
    .Y(_02976_));
 sg13g2_a21oi_1 _18382_ (.A1(net148),
    .A2(_02963_),
    .Y(_01682_),
    .B1(_02976_));
 sg13g2_nand3_1 _18383_ (.B(net763),
    .C(net706),
    .A(_09752_),
    .Y(_02977_));
 sg13g2_buf_2 _18384_ (.A(_02977_),
    .X(_02978_));
 sg13g2_nand2_1 _18385_ (.Y(_02979_),
    .A(\top_ihp.oisc.regs[44][23] ),
    .B(_02978_));
 sg13g2_o21ai_1 _18386_ (.B1(_02979_),
    .Y(_01683_),
    .A1(net285),
    .A2(_02978_));
 sg13g2_buf_8 _18387_ (.A(_02954_),
    .X(_02980_));
 sg13g2_nand2_1 _18388_ (.Y(_02981_),
    .A(\top_ihp.oisc.regs[44][24] ),
    .B(net93));
 sg13g2_o21ai_1 _18389_ (.B1(_02981_),
    .Y(_01684_),
    .A1(_10992_),
    .A2(net92));
 sg13g2_nor2_1 _18390_ (.A(\top_ihp.oisc.regs[44][25] ),
    .B(_02962_),
    .Y(_02982_));
 sg13g2_a21oi_1 _18391_ (.A1(net147),
    .A2(_02963_),
    .Y(_01685_),
    .B1(_02982_));
 sg13g2_nand2_1 _18392_ (.Y(_02983_),
    .A(\top_ihp.oisc.regs[44][26] ),
    .B(net93));
 sg13g2_o21ai_1 _18393_ (.B1(_02983_),
    .Y(_01686_),
    .A1(_10996_),
    .A2(net92));
 sg13g2_nand2_1 _18394_ (.Y(_02984_),
    .A(\top_ihp.oisc.regs[44][27] ),
    .B(_02971_));
 sg13g2_o21ai_1 _18395_ (.B1(_02984_),
    .Y(_01687_),
    .A1(_10998_),
    .A2(net92));
 sg13g2_nand2_1 _18396_ (.Y(_02985_),
    .A(\top_ihp.oisc.regs[44][28] ),
    .B(net93));
 sg13g2_o21ai_1 _18397_ (.B1(_02985_),
    .Y(_01688_),
    .A1(net284),
    .A2(_02978_));
 sg13g2_nand2_1 _18398_ (.Y(_02986_),
    .A(\top_ihp.oisc.regs[44][29] ),
    .B(_02971_));
 sg13g2_o21ai_1 _18399_ (.B1(_02986_),
    .Y(_01689_),
    .A1(_11002_),
    .A2(net92));
 sg13g2_nand2_1 _18400_ (.Y(_02987_),
    .A(\top_ihp.oisc.regs[44][2] ),
    .B(net93));
 sg13g2_o21ai_1 _18401_ (.B1(_02987_),
    .Y(_01690_),
    .A1(_11053_),
    .A2(net92));
 sg13g2_nand2_1 _18402_ (.Y(_02988_),
    .A(\top_ihp.oisc.regs[44][30] ),
    .B(net93));
 sg13g2_o21ai_1 _18403_ (.B1(_02988_),
    .Y(_01691_),
    .A1(net42),
    .A2(_02980_));
 sg13g2_nand2_1 _18404_ (.Y(_02989_),
    .A(\top_ihp.oisc.regs[44][31] ),
    .B(_02978_));
 sg13g2_o21ai_1 _18405_ (.B1(_02989_),
    .Y(_01692_),
    .A1(net251),
    .A2(_02978_));
 sg13g2_nand2_1 _18406_ (.Y(_02990_),
    .A(\top_ihp.oisc.regs[44][3] ),
    .B(net250));
 sg13g2_o21ai_1 _18407_ (.B1(_02990_),
    .Y(_01693_),
    .A1(net41),
    .A2(net92));
 sg13g2_nand2_1 _18408_ (.Y(_02991_),
    .A(\top_ihp.oisc.regs[44][4] ),
    .B(net250));
 sg13g2_o21ai_1 _18409_ (.B1(_02991_),
    .Y(_01694_),
    .A1(_11060_),
    .A2(net92));
 sg13g2_nand2_1 _18410_ (.Y(_02992_),
    .A(\top_ihp.oisc.regs[44][5] ),
    .B(_02954_));
 sg13g2_o21ai_1 _18411_ (.B1(_02992_),
    .Y(_01695_),
    .A1(_11009_),
    .A2(_02980_));
 sg13g2_nand2_1 _18412_ (.Y(_02993_),
    .A(\top_ihp.oisc.regs[44][6] ),
    .B(net250));
 sg13g2_o21ai_1 _18413_ (.B1(_02993_),
    .Y(_01696_),
    .A1(net47),
    .A2(net92));
 sg13g2_nand2_1 _18414_ (.Y(_02994_),
    .A(\top_ihp.oisc.regs[44][7] ),
    .B(net250));
 sg13g2_o21ai_1 _18415_ (.B1(_02994_),
    .Y(_01697_),
    .A1(net501),
    .A2(net249));
 sg13g2_nand2_1 _18416_ (.Y(_02995_),
    .A(\top_ihp.oisc.regs[44][8] ),
    .B(net250));
 sg13g2_o21ai_1 _18417_ (.B1(_02995_),
    .Y(_01698_),
    .A1(net107),
    .A2(net249));
 sg13g2_nand2_1 _18418_ (.Y(_02996_),
    .A(\top_ihp.oisc.regs[44][9] ),
    .B(net250));
 sg13g2_o21ai_1 _18419_ (.B1(_02996_),
    .Y(_01699_),
    .A1(net46),
    .A2(net249));
 sg13g2_nand3_1 _18420_ (.B(_10822_),
    .C(net706),
    .A(net763),
    .Y(_02997_));
 sg13g2_buf_2 _18421_ (.A(_02997_),
    .X(_02998_));
 sg13g2_buf_1 _18422_ (.A(_02998_),
    .X(_02999_));
 sg13g2_nand3_1 _18423_ (.B(net784),
    .C(net707),
    .A(net763),
    .Y(_03000_));
 sg13g2_buf_1 _18424_ (.A(_03000_),
    .X(_03001_));
 sg13g2_buf_1 _18425_ (.A(net498),
    .X(_03002_));
 sg13g2_nand2_1 _18426_ (.Y(_03003_),
    .A(\top_ihp.oisc.regs[45][0] ),
    .B(net246));
 sg13g2_o21ai_1 _18427_ (.B1(_03003_),
    .Y(_01700_),
    .A1(net45),
    .A2(net247));
 sg13g2_buf_8 _18428_ (.A(_10623_),
    .X(_03004_));
 sg13g2_nand2_1 _18429_ (.Y(_03005_),
    .A(\top_ihp.oisc.regs[45][10] ),
    .B(net246));
 sg13g2_o21ai_1 _18430_ (.B1(_03005_),
    .Y(_01701_),
    .A1(net39),
    .A2(net247));
 sg13g2_nand2_1 _18431_ (.Y(_03006_),
    .A(\top_ihp.oisc.regs[45][11] ),
    .B(net246));
 sg13g2_o21ai_1 _18432_ (.B1(_03006_),
    .Y(_01702_),
    .A1(net44),
    .A2(net247));
 sg13g2_nor2_1 _18433_ (.A(_02961_),
    .B(_11029_),
    .Y(_03007_));
 sg13g2_buf_1 _18434_ (.A(_03007_),
    .X(_03008_));
 sg13g2_nor2_1 _18435_ (.A(\top_ihp.oisc.regs[45][12] ),
    .B(net245),
    .Y(_03009_));
 sg13g2_a21oi_1 _18436_ (.A1(net153),
    .A2(net245),
    .Y(_01703_),
    .B1(_03009_));
 sg13g2_buf_8 _18437_ (.A(net314),
    .X(_03010_));
 sg13g2_nand2_1 _18438_ (.Y(_03011_),
    .A(\top_ihp.oisc.regs[45][13] ),
    .B(net246));
 sg13g2_o21ai_1 _18439_ (.B1(_03011_),
    .Y(_01704_),
    .A1(net91),
    .A2(net247));
 sg13g2_nor2_1 _18440_ (.A(\top_ihp.oisc.regs[45][14] ),
    .B(net245),
    .Y(_03012_));
 sg13g2_a21oi_1 _18441_ (.A1(net152),
    .A2(net245),
    .Y(_01705_),
    .B1(_03012_));
 sg13g2_nor2_1 _18442_ (.A(\top_ihp.oisc.regs[45][15] ),
    .B(net245),
    .Y(_03013_));
 sg13g2_a21oi_1 _18443_ (.A1(net151),
    .A2(net245),
    .Y(_01706_),
    .B1(_03013_));
 sg13g2_buf_8 _18444_ (.A(net126),
    .X(_03014_));
 sg13g2_nand2_1 _18445_ (.Y(_03015_),
    .A(\top_ihp.oisc.regs[45][16] ),
    .B(net246));
 sg13g2_o21ai_1 _18446_ (.B1(_03015_),
    .Y(_01707_),
    .A1(net38),
    .A2(net247));
 sg13g2_buf_1 _18447_ (.A(net313),
    .X(_03016_));
 sg13g2_nand2_1 _18448_ (.Y(_03017_),
    .A(\top_ihp.oisc.regs[45][17] ),
    .B(net246));
 sg13g2_o21ai_1 _18449_ (.B1(_03017_),
    .Y(_01708_),
    .A1(net90),
    .A2(net247));
 sg13g2_buf_1 _18450_ (.A(net312),
    .X(_03018_));
 sg13g2_nand2_1 _18451_ (.Y(_03019_),
    .A(\top_ihp.oisc.regs[45][18] ),
    .B(net246));
 sg13g2_o21ai_1 _18452_ (.B1(_03019_),
    .Y(_01709_),
    .A1(net89),
    .A2(net247));
 sg13g2_buf_8 _18453_ (.A(net311),
    .X(_03020_));
 sg13g2_nand2_1 _18454_ (.Y(_03021_),
    .A(\top_ihp.oisc.regs[45][19] ),
    .B(net246));
 sg13g2_o21ai_1 _18455_ (.B1(_03021_),
    .Y(_01710_),
    .A1(net88),
    .A2(net247));
 sg13g2_nor2_1 _18456_ (.A(\top_ihp.oisc.regs[45][1] ),
    .B(net245),
    .Y(_03022_));
 sg13g2_a21oi_1 _18457_ (.A1(net149),
    .A2(_03008_),
    .Y(_01711_),
    .B1(_03022_));
 sg13g2_buf_1 _18458_ (.A(net498),
    .X(_03023_));
 sg13g2_nand2_1 _18459_ (.Y(_03024_),
    .A(\top_ihp.oisc.regs[45][20] ),
    .B(net244));
 sg13g2_o21ai_1 _18460_ (.B1(_03024_),
    .Y(_01712_),
    .A1(_02842_),
    .A2(_03002_));
 sg13g2_buf_8 _18461_ (.A(_10633_),
    .X(_03025_));
 sg13g2_nand2_1 _18462_ (.Y(_03026_),
    .A(\top_ihp.oisc.regs[45][21] ),
    .B(net244));
 sg13g2_o21ai_1 _18463_ (.B1(_03026_),
    .Y(_01713_),
    .A1(net87),
    .A2(_02999_));
 sg13g2_nor2_1 _18464_ (.A(\top_ihp.oisc.regs[45][22] ),
    .B(_03007_),
    .Y(_03027_));
 sg13g2_a21oi_1 _18465_ (.A1(_10189_),
    .A2(net245),
    .Y(_01714_),
    .B1(_03027_));
 sg13g2_buf_8 _18466_ (.A(net528),
    .X(_03028_));
 sg13g2_nand2_1 _18467_ (.Y(_03029_),
    .A(\top_ihp.oisc.regs[45][23] ),
    .B(net244));
 sg13g2_o21ai_1 _18468_ (.B1(_03029_),
    .Y(_01715_),
    .A1(net243),
    .A2(_02999_));
 sg13g2_buf_1 _18469_ (.A(net309),
    .X(_03030_));
 sg13g2_buf_1 _18470_ (.A(_02998_),
    .X(_03031_));
 sg13g2_nand2_1 _18471_ (.Y(_03032_),
    .A(\top_ihp.oisc.regs[45][24] ),
    .B(net244));
 sg13g2_o21ai_1 _18472_ (.B1(_03032_),
    .Y(_01716_),
    .A1(net86),
    .A2(net242));
 sg13g2_nor2_1 _18473_ (.A(\top_ihp.oisc.regs[45][25] ),
    .B(_03007_),
    .Y(_03033_));
 sg13g2_a21oi_1 _18474_ (.A1(_10237_),
    .A2(_03008_),
    .Y(_01717_),
    .B1(_03033_));
 sg13g2_buf_1 _18475_ (.A(net125),
    .X(_03034_));
 sg13g2_nand2_1 _18476_ (.Y(_03035_),
    .A(\top_ihp.oisc.regs[45][26] ),
    .B(net244));
 sg13g2_o21ai_1 _18477_ (.B1(_03035_),
    .Y(_01718_),
    .A1(net37),
    .A2(net242));
 sg13g2_buf_1 _18478_ (.A(_10639_),
    .X(_03036_));
 sg13g2_nand2_1 _18479_ (.Y(_03037_),
    .A(\top_ihp.oisc.regs[45][27] ),
    .B(_03023_));
 sg13g2_o21ai_1 _18480_ (.B1(_03037_),
    .Y(_01719_),
    .A1(net85),
    .A2(net242));
 sg13g2_buf_8 _18481_ (.A(net515),
    .X(_03038_));
 sg13g2_nand2_1 _18482_ (.Y(_03039_),
    .A(\top_ihp.oisc.regs[45][28] ),
    .B(net244));
 sg13g2_o21ai_1 _18483_ (.B1(_03039_),
    .Y(_01720_),
    .A1(net241),
    .A2(net242));
 sg13g2_buf_8 _18484_ (.A(_10642_),
    .X(_03040_));
 sg13g2_nand2_1 _18485_ (.Y(_03041_),
    .A(\top_ihp.oisc.regs[45][29] ),
    .B(net244));
 sg13g2_o21ai_1 _18486_ (.B1(_03041_),
    .Y(_01721_),
    .A1(net84),
    .A2(net242));
 sg13g2_nand2_1 _18487_ (.Y(_03042_),
    .A(\top_ihp.oisc.regs[45][2] ),
    .B(net244));
 sg13g2_o21ai_1 _18488_ (.B1(_03042_),
    .Y(_01722_),
    .A1(net43),
    .A2(net242));
 sg13g2_nand2_1 _18489_ (.Y(_03043_),
    .A(\top_ihp.oisc.regs[45][30] ),
    .B(_03023_));
 sg13g2_o21ai_1 _18490_ (.B1(_03043_),
    .Y(_01723_),
    .A1(net42),
    .A2(net242));
 sg13g2_nand2_1 _18491_ (.Y(_03044_),
    .A(\top_ihp.oisc.regs[45][31] ),
    .B(_02998_));
 sg13g2_o21ai_1 _18492_ (.B1(_03044_),
    .Y(_01724_),
    .A1(net251),
    .A2(_03031_));
 sg13g2_nand2_1 _18493_ (.Y(_03045_),
    .A(\top_ihp.oisc.regs[45][3] ),
    .B(_03001_));
 sg13g2_o21ai_1 _18494_ (.B1(_03045_),
    .Y(_01725_),
    .A1(net41),
    .A2(_03031_));
 sg13g2_nand2_1 _18495_ (.Y(_03046_),
    .A(\top_ihp.oisc.regs[45][4] ),
    .B(net498));
 sg13g2_o21ai_1 _18496_ (.B1(_03046_),
    .Y(_01726_),
    .A1(net40),
    .A2(net242));
 sg13g2_buf_1 _18497_ (.A(_10645_),
    .X(_03047_));
 sg13g2_nand2_1 _18498_ (.Y(_03048_),
    .A(\top_ihp.oisc.regs[45][5] ),
    .B(net498));
 sg13g2_o21ai_1 _18499_ (.B1(_03048_),
    .Y(_01727_),
    .A1(net36),
    .A2(_02998_));
 sg13g2_buf_1 _18500_ (.A(net122),
    .X(_03049_));
 sg13g2_nand2_1 _18501_ (.Y(_03050_),
    .A(\top_ihp.oisc.regs[45][6] ),
    .B(net498));
 sg13g2_o21ai_1 _18502_ (.B1(_03050_),
    .Y(_01728_),
    .A1(net35),
    .A2(_02998_));
 sg13g2_nand2_1 _18503_ (.Y(_03051_),
    .A(\top_ihp.oisc.regs[45][7] ),
    .B(net498));
 sg13g2_o21ai_1 _18504_ (.B1(_03051_),
    .Y(_01729_),
    .A1(_02862_),
    .A2(_03002_));
 sg13g2_buf_8 _18505_ (.A(net305),
    .X(_03052_));
 sg13g2_nand2_1 _18506_ (.Y(_03053_),
    .A(\top_ihp.oisc.regs[45][8] ),
    .B(net498));
 sg13g2_o21ai_1 _18507_ (.B1(_03053_),
    .Y(_01730_),
    .A1(net83),
    .A2(_02998_));
 sg13g2_buf_8 _18508_ (.A(net121),
    .X(_03054_));
 sg13g2_nand2_1 _18509_ (.Y(_03055_),
    .A(\top_ihp.oisc.regs[45][9] ),
    .B(net498));
 sg13g2_o21ai_1 _18510_ (.B1(_03055_),
    .Y(_01731_),
    .A1(net34),
    .A2(_02998_));
 sg13g2_buf_2 _18511_ (.A(_09696_),
    .X(_03056_));
 sg13g2_nand3_1 _18512_ (.B(_10618_),
    .C(net708),
    .A(net741),
    .Y(_03057_));
 sg13g2_buf_1 _18513_ (.A(_03057_),
    .X(_03058_));
 sg13g2_buf_1 _18514_ (.A(net497),
    .X(_03059_));
 sg13g2_buf_1 _18515_ (.A(net497),
    .X(_03060_));
 sg13g2_nand2_1 _18516_ (.Y(_03061_),
    .A(\top_ihp.oisc.regs[46][0] ),
    .B(net239));
 sg13g2_o21ai_1 _18517_ (.B1(_03061_),
    .Y(_01732_),
    .A1(net82),
    .A2(net240));
 sg13g2_nand2_1 _18518_ (.Y(_03062_),
    .A(\top_ihp.oisc.regs[46][10] ),
    .B(_03060_));
 sg13g2_o21ai_1 _18519_ (.B1(_03062_),
    .Y(_01733_),
    .A1(net39),
    .A2(net240));
 sg13g2_buf_8 _18520_ (.A(net127),
    .X(_03063_));
 sg13g2_nand2_1 _18521_ (.Y(_03064_),
    .A(\top_ihp.oisc.regs[46][11] ),
    .B(_03060_));
 sg13g2_o21ai_1 _18522_ (.B1(_03064_),
    .Y(_01734_),
    .A1(net33),
    .A2(net240));
 sg13g2_nor2_1 _18523_ (.A(_02961_),
    .B(_10882_),
    .Y(_03065_));
 sg13g2_buf_1 _18524_ (.A(_03065_),
    .X(_03066_));
 sg13g2_nor2_1 _18525_ (.A(\top_ihp.oisc.regs[46][12] ),
    .B(net238),
    .Y(_03067_));
 sg13g2_a21oi_1 _18526_ (.A1(net153),
    .A2(net238),
    .Y(_01735_),
    .B1(_03067_));
 sg13g2_buf_1 _18527_ (.A(net497),
    .X(_03068_));
 sg13g2_nand2_1 _18528_ (.Y(_03069_),
    .A(\top_ihp.oisc.regs[46][13] ),
    .B(_03068_));
 sg13g2_o21ai_1 _18529_ (.B1(_03069_),
    .Y(_01736_),
    .A1(net91),
    .A2(net240));
 sg13g2_nor2_1 _18530_ (.A(\top_ihp.oisc.regs[46][14] ),
    .B(net238),
    .Y(_03070_));
 sg13g2_a21oi_1 _18531_ (.A1(_09978_),
    .A2(net238),
    .Y(_01737_),
    .B1(_03070_));
 sg13g2_nor2_1 _18532_ (.A(\top_ihp.oisc.regs[46][15] ),
    .B(net238),
    .Y(_03071_));
 sg13g2_a21oi_1 _18533_ (.A1(_09993_),
    .A2(net238),
    .Y(_01738_),
    .B1(_03071_));
 sg13g2_nand2_1 _18534_ (.Y(_03072_),
    .A(\top_ihp.oisc.regs[46][16] ),
    .B(net237));
 sg13g2_o21ai_1 _18535_ (.B1(_03072_),
    .Y(_01739_),
    .A1(net38),
    .A2(net240));
 sg13g2_nand2_1 _18536_ (.Y(_03073_),
    .A(\top_ihp.oisc.regs[46][17] ),
    .B(net237));
 sg13g2_o21ai_1 _18537_ (.B1(_03073_),
    .Y(_01740_),
    .A1(net90),
    .A2(net240));
 sg13g2_nand2_1 _18538_ (.Y(_03074_),
    .A(\top_ihp.oisc.regs[46][18] ),
    .B(net237));
 sg13g2_o21ai_1 _18539_ (.B1(_03074_),
    .Y(_01741_),
    .A1(net89),
    .A2(net240));
 sg13g2_nand2_1 _18540_ (.Y(_03075_),
    .A(\top_ihp.oisc.regs[46][19] ),
    .B(net237));
 sg13g2_o21ai_1 _18541_ (.B1(_03075_),
    .Y(_01742_),
    .A1(net88),
    .A2(_03059_));
 sg13g2_nor2_1 _18542_ (.A(\top_ihp.oisc.regs[46][1] ),
    .B(net238),
    .Y(_03076_));
 sg13g2_a21oi_1 _18543_ (.A1(_10128_),
    .A2(net238),
    .Y(_01743_),
    .B1(_03076_));
 sg13g2_nand2_1 _18544_ (.Y(_03077_),
    .A(\top_ihp.oisc.regs[46][20] ),
    .B(net237));
 sg13g2_o21ai_1 _18545_ (.B1(_03077_),
    .Y(_01744_),
    .A1(_10153_),
    .A2(_03059_));
 sg13g2_nand2_1 _18546_ (.Y(_03078_),
    .A(\top_ihp.oisc.regs[46][21] ),
    .B(net237));
 sg13g2_o21ai_1 _18547_ (.B1(_03078_),
    .Y(_01745_),
    .A1(_03025_),
    .A2(net240));
 sg13g2_nor2_1 _18548_ (.A(\top_ihp.oisc.regs[46][22] ),
    .B(_03066_),
    .Y(_03079_));
 sg13g2_a21oi_1 _18549_ (.A1(net148),
    .A2(_03066_),
    .Y(_01746_),
    .B1(_03079_));
 sg13g2_buf_8 _18550_ (.A(net497),
    .X(_03080_));
 sg13g2_nand2_1 _18551_ (.Y(_03081_),
    .A(\top_ihp.oisc.regs[46][23] ),
    .B(net237));
 sg13g2_o21ai_1 _18552_ (.B1(_03081_),
    .Y(_01747_),
    .A1(net243),
    .A2(net236));
 sg13g2_nand2_1 _18553_ (.Y(_03082_),
    .A(\top_ihp.oisc.regs[46][24] ),
    .B(_03068_));
 sg13g2_o21ai_1 _18554_ (.B1(_03082_),
    .Y(_01748_),
    .A1(net86),
    .A2(net236));
 sg13g2_nand2_1 _18555_ (.Y(_03083_),
    .A(\top_ihp.oisc.regs[46][25] ),
    .B(net237));
 sg13g2_o21ai_1 _18556_ (.B1(_03083_),
    .Y(_01749_),
    .A1(net97),
    .A2(net236));
 sg13g2_buf_8 _18557_ (.A(net497),
    .X(_03084_));
 sg13g2_nand2_1 _18558_ (.Y(_03085_),
    .A(\top_ihp.oisc.regs[46][26] ),
    .B(net235));
 sg13g2_o21ai_1 _18559_ (.B1(_03085_),
    .Y(_01750_),
    .A1(net37),
    .A2(net236));
 sg13g2_nand2_1 _18560_ (.Y(_03086_),
    .A(\top_ihp.oisc.regs[46][27] ),
    .B(net235));
 sg13g2_o21ai_1 _18561_ (.B1(_03086_),
    .Y(_01751_),
    .A1(net85),
    .A2(net236));
 sg13g2_nand2_1 _18562_ (.Y(_03087_),
    .A(\top_ihp.oisc.regs[46][28] ),
    .B(net235));
 sg13g2_o21ai_1 _18563_ (.B1(_03087_),
    .Y(_01752_),
    .A1(net241),
    .A2(_03080_));
 sg13g2_nand2_1 _18564_ (.Y(_03088_),
    .A(\top_ihp.oisc.regs[46][29] ),
    .B(net235));
 sg13g2_o21ai_1 _18565_ (.B1(_03088_),
    .Y(_01753_),
    .A1(net84),
    .A2(net236));
 sg13g2_buf_1 _18566_ (.A(net131),
    .X(_03089_));
 sg13g2_nand2_1 _18567_ (.Y(_03090_),
    .A(\top_ihp.oisc.regs[46][2] ),
    .B(net235));
 sg13g2_o21ai_1 _18568_ (.B1(_03090_),
    .Y(_01754_),
    .A1(net32),
    .A2(net236));
 sg13g2_buf_8 _18569_ (.A(net124),
    .X(_03091_));
 sg13g2_nand2_1 _18570_ (.Y(_03092_),
    .A(\top_ihp.oisc.regs[46][30] ),
    .B(_03084_));
 sg13g2_o21ai_1 _18571_ (.B1(_03092_),
    .Y(_01755_),
    .A1(net31),
    .A2(_03080_));
 sg13g2_nand2_1 _18572_ (.Y(_03093_),
    .A(\top_ihp.oisc.regs[46][31] ),
    .B(net235));
 sg13g2_o21ai_1 _18573_ (.B1(_03093_),
    .Y(_01756_),
    .A1(net52),
    .A2(net236));
 sg13g2_buf_2 _18574_ (.A(net130),
    .X(_03094_));
 sg13g2_nand2_1 _18575_ (.Y(_03095_),
    .A(\top_ihp.oisc.regs[46][3] ),
    .B(net235));
 sg13g2_o21ai_1 _18576_ (.B1(_03095_),
    .Y(_01757_),
    .A1(net30),
    .A2(net239));
 sg13g2_buf_1 _18577_ (.A(net129),
    .X(_03096_));
 sg13g2_nand2_1 _18578_ (.Y(_03097_),
    .A(\top_ihp.oisc.regs[46][4] ),
    .B(net235));
 sg13g2_o21ai_1 _18579_ (.B1(_03097_),
    .Y(_01758_),
    .A1(net29),
    .A2(net239));
 sg13g2_nand2_1 _18580_ (.Y(_03098_),
    .A(\top_ihp.oisc.regs[46][5] ),
    .B(_03084_));
 sg13g2_o21ai_1 _18581_ (.B1(_03098_),
    .Y(_01759_),
    .A1(net36),
    .A2(net239));
 sg13g2_nand2_1 _18582_ (.Y(_03099_),
    .A(\top_ihp.oisc.regs[46][6] ),
    .B(_03058_));
 sg13g2_o21ai_1 _18583_ (.B1(_03099_),
    .Y(_01760_),
    .A1(net35),
    .A2(net239));
 sg13g2_nand2_1 _18584_ (.Y(_03100_),
    .A(\top_ihp.oisc.regs[46][7] ),
    .B(net497));
 sg13g2_o21ai_1 _18585_ (.B1(_03100_),
    .Y(_01761_),
    .A1(net139),
    .A2(net239));
 sg13g2_nand2_1 _18586_ (.Y(_03101_),
    .A(\top_ihp.oisc.regs[46][8] ),
    .B(net497));
 sg13g2_o21ai_1 _18587_ (.B1(_03101_),
    .Y(_01762_),
    .A1(_03052_),
    .A2(net239));
 sg13g2_nand2_1 _18588_ (.Y(_03102_),
    .A(\top_ihp.oisc.regs[46][9] ),
    .B(net497));
 sg13g2_o21ai_1 _18589_ (.B1(_03102_),
    .Y(_01763_),
    .A1(net34),
    .A2(net239));
 sg13g2_nand3_1 _18590_ (.B(net763),
    .C(_10881_),
    .A(net785),
    .Y(_03103_));
 sg13g2_buf_2 _18591_ (.A(_03103_),
    .X(_03104_));
 sg13g2_buf_1 _18592_ (.A(_03104_),
    .X(_03105_));
 sg13g2_nand3_1 _18593_ (.B(_10618_),
    .C(_10831_),
    .A(_10570_),
    .Y(_03106_));
 sg13g2_buf_1 _18594_ (.A(_03106_),
    .X(_03107_));
 sg13g2_buf_1 _18595_ (.A(net496),
    .X(_03108_));
 sg13g2_nand2_1 _18596_ (.Y(_03109_),
    .A(\top_ihp.oisc.regs[47][0] ),
    .B(net233));
 sg13g2_o21ai_1 _18597_ (.B1(_03109_),
    .Y(_01764_),
    .A1(net82),
    .A2(net234));
 sg13g2_nand2_1 _18598_ (.Y(_03110_),
    .A(\top_ihp.oisc.regs[47][10] ),
    .B(net233));
 sg13g2_o21ai_1 _18599_ (.B1(_03110_),
    .Y(_01765_),
    .A1(net39),
    .A2(net234));
 sg13g2_nand2_1 _18600_ (.Y(_03111_),
    .A(\top_ihp.oisc.regs[47][11] ),
    .B(net233));
 sg13g2_o21ai_1 _18601_ (.B1(_03111_),
    .Y(_01766_),
    .A1(net33),
    .A2(net234));
 sg13g2_nor4_2 _18602_ (.A(_09750_),
    .B(_09743_),
    .C(_02961_),
    .Y(_03112_),
    .D(_10823_));
 sg13g2_buf_1 _18603_ (.A(_03112_),
    .X(_03113_));
 sg13g2_nor2_1 _18604_ (.A(\top_ihp.oisc.regs[47][12] ),
    .B(net761),
    .Y(_03114_));
 sg13g2_a21oi_1 _18605_ (.A1(net153),
    .A2(net761),
    .Y(_01767_),
    .B1(_03114_));
 sg13g2_nand2_1 _18606_ (.Y(_03115_),
    .A(\top_ihp.oisc.regs[47][13] ),
    .B(net233));
 sg13g2_o21ai_1 _18607_ (.B1(_03115_),
    .Y(_01768_),
    .A1(net91),
    .A2(net234));
 sg13g2_nor2_1 _18608_ (.A(\top_ihp.oisc.regs[47][14] ),
    .B(net761),
    .Y(_03116_));
 sg13g2_a21oi_1 _18609_ (.A1(_09978_),
    .A2(net761),
    .Y(_01769_),
    .B1(_03116_));
 sg13g2_nor2_1 _18610_ (.A(\top_ihp.oisc.regs[47][15] ),
    .B(net761),
    .Y(_03117_));
 sg13g2_a21oi_1 _18611_ (.A1(net151),
    .A2(net761),
    .Y(_01770_),
    .B1(_03117_));
 sg13g2_nand2_1 _18612_ (.Y(_03118_),
    .A(\top_ihp.oisc.regs[47][16] ),
    .B(net233));
 sg13g2_o21ai_1 _18613_ (.B1(_03118_),
    .Y(_01771_),
    .A1(net38),
    .A2(net234));
 sg13g2_nand2_1 _18614_ (.Y(_03119_),
    .A(\top_ihp.oisc.regs[47][17] ),
    .B(net233));
 sg13g2_o21ai_1 _18615_ (.B1(_03119_),
    .Y(_01772_),
    .A1(net90),
    .A2(net234));
 sg13g2_nand2_1 _18616_ (.Y(_03120_),
    .A(\top_ihp.oisc.regs[47][18] ),
    .B(net233));
 sg13g2_o21ai_1 _18617_ (.B1(_03120_),
    .Y(_01773_),
    .A1(net89),
    .A2(net234));
 sg13g2_nand2_1 _18618_ (.Y(_03121_),
    .A(\top_ihp.oisc.regs[47][19] ),
    .B(net233));
 sg13g2_o21ai_1 _18619_ (.B1(_03121_),
    .Y(_01774_),
    .A1(net88),
    .A2(net234));
 sg13g2_nor2_1 _18620_ (.A(\top_ihp.oisc.regs[47][1] ),
    .B(_03113_),
    .Y(_03122_));
 sg13g2_a21oi_1 _18621_ (.A1(_10128_),
    .A2(_03113_),
    .Y(_01775_),
    .B1(_03122_));
 sg13g2_buf_1 _18622_ (.A(net496),
    .X(_03123_));
 sg13g2_nand2_1 _18623_ (.Y(_03124_),
    .A(\top_ihp.oisc.regs[47][20] ),
    .B(net232));
 sg13g2_o21ai_1 _18624_ (.B1(_03124_),
    .Y(_01776_),
    .A1(_02842_),
    .A2(_03108_));
 sg13g2_nand2_1 _18625_ (.Y(_03125_),
    .A(\top_ihp.oisc.regs[47][21] ),
    .B(net232));
 sg13g2_o21ai_1 _18626_ (.B1(_03125_),
    .Y(_01777_),
    .A1(net87),
    .A2(_03105_));
 sg13g2_nor2_1 _18627_ (.A(\top_ihp.oisc.regs[47][22] ),
    .B(_03112_),
    .Y(_03126_));
 sg13g2_a21oi_1 _18628_ (.A1(net148),
    .A2(net761),
    .Y(_01778_),
    .B1(_03126_));
 sg13g2_nand2_1 _18629_ (.Y(_03127_),
    .A(\top_ihp.oisc.regs[47][23] ),
    .B(net232));
 sg13g2_o21ai_1 _18630_ (.B1(_03127_),
    .Y(_01779_),
    .A1(net243),
    .A2(_03105_));
 sg13g2_buf_1 _18631_ (.A(_03104_),
    .X(_03128_));
 sg13g2_nand2_1 _18632_ (.Y(_03129_),
    .A(\top_ihp.oisc.regs[47][24] ),
    .B(net232));
 sg13g2_o21ai_1 _18633_ (.B1(_03129_),
    .Y(_01780_),
    .A1(net86),
    .A2(net231));
 sg13g2_nor2_1 _18634_ (.A(\top_ihp.oisc.regs[47][25] ),
    .B(_03112_),
    .Y(_03130_));
 sg13g2_a21oi_1 _18635_ (.A1(_10237_),
    .A2(net761),
    .Y(_01781_),
    .B1(_03130_));
 sg13g2_nand2_1 _18636_ (.Y(_03131_),
    .A(\top_ihp.oisc.regs[47][26] ),
    .B(net232));
 sg13g2_o21ai_1 _18637_ (.B1(_03131_),
    .Y(_01782_),
    .A1(net37),
    .A2(_03128_));
 sg13g2_nand2_1 _18638_ (.Y(_03132_),
    .A(\top_ihp.oisc.regs[47][27] ),
    .B(net232));
 sg13g2_o21ai_1 _18639_ (.B1(_03132_),
    .Y(_01783_),
    .A1(net85),
    .A2(net231));
 sg13g2_nand2_1 _18640_ (.Y(_03133_),
    .A(\top_ihp.oisc.regs[47][28] ),
    .B(net232));
 sg13g2_o21ai_1 _18641_ (.B1(_03133_),
    .Y(_01784_),
    .A1(net241),
    .A2(net231));
 sg13g2_nand2_1 _18642_ (.Y(_03134_),
    .A(\top_ihp.oisc.regs[47][29] ),
    .B(_03123_));
 sg13g2_o21ai_1 _18643_ (.B1(_03134_),
    .Y(_01785_),
    .A1(net84),
    .A2(net231));
 sg13g2_nand2_1 _18644_ (.Y(_03135_),
    .A(\top_ihp.oisc.regs[47][2] ),
    .B(net232));
 sg13g2_o21ai_1 _18645_ (.B1(_03135_),
    .Y(_01786_),
    .A1(net32),
    .A2(net231));
 sg13g2_nand2_1 _18646_ (.Y(_03136_),
    .A(\top_ihp.oisc.regs[47][30] ),
    .B(_03123_));
 sg13g2_o21ai_1 _18647_ (.B1(_03136_),
    .Y(_01787_),
    .A1(net31),
    .A2(_03128_));
 sg13g2_nand2_1 _18648_ (.Y(_03137_),
    .A(\top_ihp.oisc.regs[47][31] ),
    .B(_03104_));
 sg13g2_o21ai_1 _18649_ (.B1(_03137_),
    .Y(_01788_),
    .A1(net251),
    .A2(net231));
 sg13g2_nand2_1 _18650_ (.Y(_03138_),
    .A(\top_ihp.oisc.regs[47][3] ),
    .B(net496));
 sg13g2_o21ai_1 _18651_ (.B1(_03138_),
    .Y(_01789_),
    .A1(net30),
    .A2(net231));
 sg13g2_nand2_1 _18652_ (.Y(_03139_),
    .A(\top_ihp.oisc.regs[47][4] ),
    .B(net496));
 sg13g2_o21ai_1 _18653_ (.B1(_03139_),
    .Y(_01790_),
    .A1(_03096_),
    .A2(net231));
 sg13g2_nand2_1 _18654_ (.Y(_03140_),
    .A(\top_ihp.oisc.regs[47][5] ),
    .B(net496));
 sg13g2_o21ai_1 _18655_ (.B1(_03140_),
    .Y(_01791_),
    .A1(net36),
    .A2(_03104_));
 sg13g2_nand2_1 _18656_ (.Y(_03141_),
    .A(\top_ihp.oisc.regs[47][6] ),
    .B(_03107_));
 sg13g2_o21ai_1 _18657_ (.B1(_03141_),
    .Y(_01792_),
    .A1(net35),
    .A2(_03104_));
 sg13g2_nand2_1 _18658_ (.Y(_03142_),
    .A(\top_ihp.oisc.regs[47][7] ),
    .B(net496));
 sg13g2_o21ai_1 _18659_ (.B1(_03142_),
    .Y(_01793_),
    .A1(_02862_),
    .A2(_03108_));
 sg13g2_nand2_1 _18660_ (.Y(_03143_),
    .A(\top_ihp.oisc.regs[47][8] ),
    .B(net496));
 sg13g2_o21ai_1 _18661_ (.B1(_03143_),
    .Y(_01794_),
    .A1(net83),
    .A2(_03104_));
 sg13g2_nand2_1 _18662_ (.Y(_03144_),
    .A(\top_ihp.oisc.regs[47][9] ),
    .B(net496));
 sg13g2_o21ai_1 _18663_ (.B1(_03144_),
    .Y(_01795_),
    .A1(net34),
    .A2(_03104_));
 sg13g2_nor2b_1 _18664_ (.A(_09731_),
    .B_N(_09737_),
    .Y(_03145_));
 sg13g2_buf_2 _18665_ (.A(_03145_),
    .X(_03146_));
 sg13g2_and2_1 _18666_ (.A(_09752_),
    .B(_03146_),
    .X(_03147_));
 sg13g2_buf_1 _18667_ (.A(_03147_),
    .X(_03148_));
 sg13g2_nand2_1 _18668_ (.Y(_03149_),
    .A(_09726_),
    .B(_03148_));
 sg13g2_buf_1 _18669_ (.A(_03149_),
    .X(_03150_));
 sg13g2_buf_1 _18670_ (.A(net635),
    .X(_03151_));
 sg13g2_buf_1 _18671_ (.A(_03149_),
    .X(_03152_));
 sg13g2_nand2_1 _18672_ (.Y(_03153_),
    .A(\top_ihp.oisc.regs[48][0] ),
    .B(_03152_));
 sg13g2_o21ai_1 _18673_ (.B1(_03153_),
    .Y(_01796_),
    .A1(net82),
    .A2(_03151_));
 sg13g2_nand2_1 _18674_ (.Y(_03154_),
    .A(\top_ihp.oisc.regs[48][10] ),
    .B(net634));
 sg13g2_o21ai_1 _18675_ (.B1(_03154_),
    .Y(_01797_),
    .A1(net39),
    .A2(net495));
 sg13g2_nand2_1 _18676_ (.Y(_03155_),
    .A(\top_ihp.oisc.regs[48][11] ),
    .B(net634));
 sg13g2_o21ai_1 _18677_ (.B1(_03155_),
    .Y(_01798_),
    .A1(_03063_),
    .A2(net495));
 sg13g2_nand2_1 _18678_ (.Y(_03156_),
    .A(\top_ihp.oisc.regs[48][12] ),
    .B(_03152_));
 sg13g2_o21ai_1 _18679_ (.B1(_03156_),
    .Y(_01799_),
    .A1(net104),
    .A2(_03151_));
 sg13g2_nand2_1 _18680_ (.Y(_03157_),
    .A(\top_ihp.oisc.regs[48][13] ),
    .B(net634));
 sg13g2_o21ai_1 _18681_ (.B1(_03157_),
    .Y(_01800_),
    .A1(net91),
    .A2(net495));
 sg13g2_nand2_1 _18682_ (.Y(_03158_),
    .A(\top_ihp.oisc.regs[48][14] ),
    .B(net634));
 sg13g2_o21ai_1 _18683_ (.B1(_03158_),
    .Y(_01801_),
    .A1(net103),
    .A2(net495));
 sg13g2_nand2_1 _18684_ (.Y(_03159_),
    .A(\top_ihp.oisc.regs[48][15] ),
    .B(net634));
 sg13g2_o21ai_1 _18685_ (.B1(_03159_),
    .Y(_01802_),
    .A1(net98),
    .A2(net495));
 sg13g2_nand2_1 _18686_ (.Y(_03160_),
    .A(\top_ihp.oisc.regs[48][16] ),
    .B(net634));
 sg13g2_o21ai_1 _18687_ (.B1(_03160_),
    .Y(_01803_),
    .A1(net38),
    .A2(net495));
 sg13g2_buf_1 _18688_ (.A(net635),
    .X(_03161_));
 sg13g2_nand2_1 _18689_ (.Y(_03162_),
    .A(\top_ihp.oisc.regs[48][17] ),
    .B(net494));
 sg13g2_o21ai_1 _18690_ (.B1(_03162_),
    .Y(_01804_),
    .A1(net90),
    .A2(net495));
 sg13g2_nand2_1 _18691_ (.Y(_03163_),
    .A(\top_ihp.oisc.regs[48][18] ),
    .B(_03161_));
 sg13g2_o21ai_1 _18692_ (.B1(_03163_),
    .Y(_01805_),
    .A1(net89),
    .A2(net495));
 sg13g2_buf_1 _18693_ (.A(net635),
    .X(_03164_));
 sg13g2_nand2_1 _18694_ (.Y(_03165_),
    .A(\top_ihp.oisc.regs[48][19] ),
    .B(net494));
 sg13g2_o21ai_1 _18695_ (.B1(_03165_),
    .Y(_01806_),
    .A1(net88),
    .A2(net493));
 sg13g2_nand2_1 _18696_ (.Y(_03166_),
    .A(\top_ihp.oisc.regs[48][1] ),
    .B(net494));
 sg13g2_o21ai_1 _18697_ (.B1(_03166_),
    .Y(_01807_),
    .A1(net102),
    .A2(net493));
 sg13g2_nand2_1 _18698_ (.Y(_03167_),
    .A(\top_ihp.oisc.regs[48][20] ),
    .B(net494));
 sg13g2_o21ai_1 _18699_ (.B1(_03167_),
    .Y(_01808_),
    .A1(net636),
    .A2(net493));
 sg13g2_nand2_1 _18700_ (.Y(_03168_),
    .A(\top_ihp.oisc.regs[48][21] ),
    .B(net494));
 sg13g2_o21ai_1 _18701_ (.B1(_03168_),
    .Y(_01809_),
    .A1(net87),
    .A2(net493));
 sg13g2_nand2_1 _18702_ (.Y(_03169_),
    .A(\top_ihp.oisc.regs[48][22] ),
    .B(net494));
 sg13g2_o21ai_1 _18703_ (.B1(_03169_),
    .Y(_01810_),
    .A1(net101),
    .A2(net493));
 sg13g2_nand2_1 _18704_ (.Y(_03170_),
    .A(\top_ihp.oisc.regs[48][23] ),
    .B(net494));
 sg13g2_o21ai_1 _18705_ (.B1(_03170_),
    .Y(_01811_),
    .A1(net243),
    .A2(_03164_));
 sg13g2_nand2_1 _18706_ (.Y(_03171_),
    .A(\top_ihp.oisc.regs[48][24] ),
    .B(_03161_));
 sg13g2_o21ai_1 _18707_ (.B1(_03171_),
    .Y(_01812_),
    .A1(net86),
    .A2(_03164_));
 sg13g2_nand2_1 _18708_ (.Y(_03172_),
    .A(\top_ihp.oisc.regs[48][25] ),
    .B(net494));
 sg13g2_o21ai_1 _18709_ (.B1(_03172_),
    .Y(_01813_),
    .A1(net97),
    .A2(net493));
 sg13g2_buf_1 _18710_ (.A(net635),
    .X(_03173_));
 sg13g2_nand2_1 _18711_ (.Y(_03174_),
    .A(\top_ihp.oisc.regs[48][26] ),
    .B(net492));
 sg13g2_o21ai_1 _18712_ (.B1(_03174_),
    .Y(_01814_),
    .A1(net37),
    .A2(net493));
 sg13g2_nand2_1 _18713_ (.Y(_03175_),
    .A(\top_ihp.oisc.regs[48][27] ),
    .B(net492));
 sg13g2_o21ai_1 _18714_ (.B1(_03175_),
    .Y(_01815_),
    .A1(net85),
    .A2(net493));
 sg13g2_buf_1 _18715_ (.A(net635),
    .X(_03176_));
 sg13g2_nand2_1 _18716_ (.Y(_03177_),
    .A(\top_ihp.oisc.regs[48][28] ),
    .B(net492));
 sg13g2_o21ai_1 _18717_ (.B1(_03177_),
    .Y(_01816_),
    .A1(net241),
    .A2(net491));
 sg13g2_nand2_1 _18718_ (.Y(_03178_),
    .A(\top_ihp.oisc.regs[48][29] ),
    .B(_03173_));
 sg13g2_o21ai_1 _18719_ (.B1(_03178_),
    .Y(_01817_),
    .A1(net84),
    .A2(net491));
 sg13g2_nand2_1 _18720_ (.Y(_03179_),
    .A(\top_ihp.oisc.regs[48][2] ),
    .B(_03173_));
 sg13g2_o21ai_1 _18721_ (.B1(_03179_),
    .Y(_01818_),
    .A1(net32),
    .A2(_03176_));
 sg13g2_nand2_1 _18722_ (.Y(_03180_),
    .A(\top_ihp.oisc.regs[48][30] ),
    .B(net492));
 sg13g2_o21ai_1 _18723_ (.B1(_03180_),
    .Y(_01819_),
    .A1(net31),
    .A2(net491));
 sg13g2_nand2_1 _18724_ (.Y(_03181_),
    .A(\top_ihp.oisc.regs[48][31] ),
    .B(net492));
 sg13g2_o21ai_1 _18725_ (.B1(_03181_),
    .Y(_01820_),
    .A1(net251),
    .A2(net491));
 sg13g2_nand2_1 _18726_ (.Y(_03182_),
    .A(\top_ihp.oisc.regs[48][3] ),
    .B(net492));
 sg13g2_o21ai_1 _18727_ (.B1(_03182_),
    .Y(_01821_),
    .A1(net30),
    .A2(net491));
 sg13g2_nand2_1 _18728_ (.Y(_03183_),
    .A(\top_ihp.oisc.regs[48][4] ),
    .B(net492));
 sg13g2_o21ai_1 _18729_ (.B1(_03183_),
    .Y(_01822_),
    .A1(_03096_),
    .A2(net491));
 sg13g2_nand2_1 _18730_ (.Y(_03184_),
    .A(\top_ihp.oisc.regs[48][5] ),
    .B(net492));
 sg13g2_o21ai_1 _18731_ (.B1(_03184_),
    .Y(_01823_),
    .A1(net36),
    .A2(net491));
 sg13g2_nand2_1 _18732_ (.Y(_03185_),
    .A(\top_ihp.oisc.regs[48][6] ),
    .B(net635));
 sg13g2_o21ai_1 _18733_ (.B1(_03185_),
    .Y(_01824_),
    .A1(net35),
    .A2(net491));
 sg13g2_nand2_1 _18734_ (.Y(_03186_),
    .A(\top_ihp.oisc.regs[48][7] ),
    .B(_03150_));
 sg13g2_o21ai_1 _18735_ (.B1(_03186_),
    .Y(_01825_),
    .A1(net501),
    .A2(_03176_));
 sg13g2_nand2_1 _18736_ (.Y(_03187_),
    .A(\top_ihp.oisc.regs[48][8] ),
    .B(net635));
 sg13g2_o21ai_1 _18737_ (.B1(_03187_),
    .Y(_01826_),
    .A1(net83),
    .A2(net634));
 sg13g2_nand2_1 _18738_ (.Y(_03188_),
    .A(\top_ihp.oisc.regs[48][9] ),
    .B(net635));
 sg13g2_o21ai_1 _18739_ (.B1(_03188_),
    .Y(_01827_),
    .A1(net34),
    .A2(net634));
 sg13g2_nand2_1 _18740_ (.Y(_03189_),
    .A(net784),
    .B(_03146_));
 sg13g2_nand2b_1 _18741_ (.Y(_03190_),
    .B(_09725_),
    .A_N(_03189_));
 sg13g2_buf_1 _18742_ (.A(_03190_),
    .X(_03191_));
 sg13g2_buf_1 _18743_ (.A(_03191_),
    .X(_03192_));
 sg13g2_buf_1 _18744_ (.A(net703),
    .X(_03193_));
 sg13g2_buf_1 _18745_ (.A(_03191_),
    .X(_03194_));
 sg13g2_nand2_1 _18746_ (.Y(_03195_),
    .A(\top_ihp.oisc.regs[49][0] ),
    .B(net702));
 sg13g2_o21ai_1 _18747_ (.B1(_03195_),
    .Y(_01828_),
    .A1(net82),
    .A2(_03193_));
 sg13g2_nand2_1 _18748_ (.Y(_03196_),
    .A(\top_ihp.oisc.regs[49][10] ),
    .B(_03194_));
 sg13g2_o21ai_1 _18749_ (.B1(_03196_),
    .Y(_01829_),
    .A1(net39),
    .A2(net633));
 sg13g2_nand2_1 _18750_ (.Y(_03197_),
    .A(\top_ihp.oisc.regs[49][11] ),
    .B(net702));
 sg13g2_o21ai_1 _18751_ (.B1(_03197_),
    .Y(_01830_),
    .A1(net33),
    .A2(net633));
 sg13g2_nand2_1 _18752_ (.Y(_03198_),
    .A(\top_ihp.oisc.regs[49][12] ),
    .B(net702));
 sg13g2_o21ai_1 _18753_ (.B1(_03198_),
    .Y(_01831_),
    .A1(net104),
    .A2(net633));
 sg13g2_nand2_1 _18754_ (.Y(_03199_),
    .A(\top_ihp.oisc.regs[49][13] ),
    .B(net702));
 sg13g2_o21ai_1 _18755_ (.B1(_03199_),
    .Y(_01832_),
    .A1(net91),
    .A2(net633));
 sg13g2_nand2_1 _18756_ (.Y(_03200_),
    .A(\top_ihp.oisc.regs[49][14] ),
    .B(net702));
 sg13g2_o21ai_1 _18757_ (.B1(_03200_),
    .Y(_01833_),
    .A1(net103),
    .A2(net633));
 sg13g2_nand2_1 _18758_ (.Y(_03201_),
    .A(\top_ihp.oisc.regs[49][15] ),
    .B(net702));
 sg13g2_o21ai_1 _18759_ (.B1(_03201_),
    .Y(_01834_),
    .A1(_02879_),
    .A2(net633));
 sg13g2_nand2_1 _18760_ (.Y(_03202_),
    .A(\top_ihp.oisc.regs[49][16] ),
    .B(_03194_));
 sg13g2_o21ai_1 _18761_ (.B1(_03202_),
    .Y(_01835_),
    .A1(net38),
    .A2(net633));
 sg13g2_buf_1 _18762_ (.A(net703),
    .X(_03203_));
 sg13g2_nand2_1 _18763_ (.Y(_03204_),
    .A(\top_ihp.oisc.regs[49][17] ),
    .B(net632));
 sg13g2_o21ai_1 _18764_ (.B1(_03204_),
    .Y(_01836_),
    .A1(net90),
    .A2(net633));
 sg13g2_nand2_1 _18765_ (.Y(_03205_),
    .A(\top_ihp.oisc.regs[49][18] ),
    .B(_03203_));
 sg13g2_o21ai_1 _18766_ (.B1(_03205_),
    .Y(_01837_),
    .A1(net89),
    .A2(_03193_));
 sg13g2_buf_2 _18767_ (.A(net703),
    .X(_03206_));
 sg13g2_nand2_1 _18768_ (.Y(_03207_),
    .A(\top_ihp.oisc.regs[49][19] ),
    .B(net632));
 sg13g2_o21ai_1 _18769_ (.B1(_03207_),
    .Y(_01838_),
    .A1(net88),
    .A2(net631));
 sg13g2_nand2_1 _18770_ (.Y(_03208_),
    .A(\top_ihp.oisc.regs[49][1] ),
    .B(net632));
 sg13g2_o21ai_1 _18771_ (.B1(_03208_),
    .Y(_01839_),
    .A1(net102),
    .A2(net631));
 sg13g2_nand2_1 _18772_ (.Y(_03209_),
    .A(\top_ihp.oisc.regs[49][20] ),
    .B(net632));
 sg13g2_o21ai_1 _18773_ (.B1(_03209_),
    .Y(_01840_),
    .A1(net636),
    .A2(net631));
 sg13g2_nand2_1 _18774_ (.Y(_03210_),
    .A(\top_ihp.oisc.regs[49][21] ),
    .B(net632));
 sg13g2_o21ai_1 _18775_ (.B1(_03210_),
    .Y(_01841_),
    .A1(net87),
    .A2(net631));
 sg13g2_nand2_1 _18776_ (.Y(_03211_),
    .A(\top_ihp.oisc.regs[49][22] ),
    .B(net632));
 sg13g2_o21ai_1 _18777_ (.B1(_03211_),
    .Y(_01842_),
    .A1(net101),
    .A2(net631));
 sg13g2_nand2_1 _18778_ (.Y(_03212_),
    .A(\top_ihp.oisc.regs[49][23] ),
    .B(net632));
 sg13g2_o21ai_1 _18779_ (.B1(_03212_),
    .Y(_01843_),
    .A1(net243),
    .A2(net631));
 sg13g2_nand2_1 _18780_ (.Y(_03213_),
    .A(\top_ihp.oisc.regs[49][24] ),
    .B(_03203_));
 sg13g2_o21ai_1 _18781_ (.B1(_03213_),
    .Y(_01844_),
    .A1(net86),
    .A2(net631));
 sg13g2_nand2_1 _18782_ (.Y(_03214_),
    .A(\top_ihp.oisc.regs[49][25] ),
    .B(net632));
 sg13g2_o21ai_1 _18783_ (.B1(_03214_),
    .Y(_01845_),
    .A1(net97),
    .A2(_03206_));
 sg13g2_buf_1 _18784_ (.A(net703),
    .X(_03215_));
 sg13g2_nand2_1 _18785_ (.Y(_03216_),
    .A(\top_ihp.oisc.regs[49][26] ),
    .B(_03215_));
 sg13g2_o21ai_1 _18786_ (.B1(_03216_),
    .Y(_01846_),
    .A1(net37),
    .A2(_03206_));
 sg13g2_nand2_1 _18787_ (.Y(_03217_),
    .A(\top_ihp.oisc.regs[49][27] ),
    .B(_03215_));
 sg13g2_o21ai_1 _18788_ (.B1(_03217_),
    .Y(_01847_),
    .A1(net85),
    .A2(net631));
 sg13g2_buf_1 _18789_ (.A(net703),
    .X(_03218_));
 sg13g2_nand2_1 _18790_ (.Y(_03219_),
    .A(\top_ihp.oisc.regs[49][28] ),
    .B(net630));
 sg13g2_o21ai_1 _18791_ (.B1(_03219_),
    .Y(_01848_),
    .A1(net241),
    .A2(net629));
 sg13g2_nand2_1 _18792_ (.Y(_03220_),
    .A(\top_ihp.oisc.regs[49][29] ),
    .B(net630));
 sg13g2_o21ai_1 _18793_ (.B1(_03220_),
    .Y(_01849_),
    .A1(net84),
    .A2(net629));
 sg13g2_nand2_1 _18794_ (.Y(_03221_),
    .A(\top_ihp.oisc.regs[49][2] ),
    .B(net630));
 sg13g2_o21ai_1 _18795_ (.B1(_03221_),
    .Y(_01850_),
    .A1(net32),
    .A2(net629));
 sg13g2_nand2_1 _18796_ (.Y(_03222_),
    .A(\top_ihp.oisc.regs[49][30] ),
    .B(net630));
 sg13g2_o21ai_1 _18797_ (.B1(_03222_),
    .Y(_01851_),
    .A1(net31),
    .A2(_03218_));
 sg13g2_nand2_1 _18798_ (.Y(_03223_),
    .A(\top_ihp.oisc.regs[49][31] ),
    .B(net630));
 sg13g2_o21ai_1 _18799_ (.B1(_03223_),
    .Y(_01852_),
    .A1(net251),
    .A2(_03218_));
 sg13g2_nand2_1 _18800_ (.Y(_03224_),
    .A(\top_ihp.oisc.regs[49][3] ),
    .B(net630));
 sg13g2_o21ai_1 _18801_ (.B1(_03224_),
    .Y(_01853_),
    .A1(net30),
    .A2(net629));
 sg13g2_nand2_1 _18802_ (.Y(_03225_),
    .A(\top_ihp.oisc.regs[49][4] ),
    .B(net630));
 sg13g2_o21ai_1 _18803_ (.B1(_03225_),
    .Y(_01854_),
    .A1(net29),
    .A2(net629));
 sg13g2_nand2_1 _18804_ (.Y(_03226_),
    .A(\top_ihp.oisc.regs[49][5] ),
    .B(net630));
 sg13g2_o21ai_1 _18805_ (.B1(_03226_),
    .Y(_01855_),
    .A1(net36),
    .A2(net629));
 sg13g2_nand2_1 _18806_ (.Y(_03227_),
    .A(\top_ihp.oisc.regs[49][6] ),
    .B(net703));
 sg13g2_o21ai_1 _18807_ (.B1(_03227_),
    .Y(_01856_),
    .A1(net35),
    .A2(net629));
 sg13g2_nand2_1 _18808_ (.Y(_03228_),
    .A(\top_ihp.oisc.regs[49][7] ),
    .B(net703));
 sg13g2_o21ai_1 _18809_ (.B1(_03228_),
    .Y(_01857_),
    .A1(net501),
    .A2(net629));
 sg13g2_nand2_1 _18810_ (.Y(_03229_),
    .A(\top_ihp.oisc.regs[49][8] ),
    .B(_03192_));
 sg13g2_o21ai_1 _18811_ (.B1(_03229_),
    .Y(_01858_),
    .A1(net83),
    .A2(net702));
 sg13g2_nand2_1 _18812_ (.Y(_03230_),
    .A(\top_ihp.oisc.regs[49][9] ),
    .B(net703));
 sg13g2_o21ai_1 _18813_ (.B1(_03230_),
    .Y(_01859_),
    .A1(net34),
    .A2(net702));
 sg13g2_nand2_1 _18814_ (.Y(_03231_),
    .A(_09754_),
    .B(net762));
 sg13g2_buf_1 _18815_ (.A(_03231_),
    .X(_03232_));
 sg13g2_buf_1 _18816_ (.A(net628),
    .X(_03233_));
 sg13g2_buf_1 _18817_ (.A(_03231_),
    .X(_03234_));
 sg13g2_nand2_1 _18818_ (.Y(_03235_),
    .A(\top_ihp.oisc.regs[4][0] ),
    .B(net627));
 sg13g2_o21ai_1 _18819_ (.B1(_03235_),
    .Y(_01860_),
    .A1(_03056_),
    .A2(net490));
 sg13g2_nand2_1 _18820_ (.Y(_03236_),
    .A(\top_ihp.oisc.regs[4][10] ),
    .B(net627));
 sg13g2_o21ai_1 _18821_ (.B1(_03236_),
    .Y(_01861_),
    .A1(net39),
    .A2(net490));
 sg13g2_nand2_1 _18822_ (.Y(_03237_),
    .A(\top_ihp.oisc.regs[4][11] ),
    .B(net627));
 sg13g2_o21ai_1 _18823_ (.B1(_03237_),
    .Y(_01862_),
    .A1(_03063_),
    .A2(net490));
 sg13g2_nand2_1 _18824_ (.Y(_03238_),
    .A(\top_ihp.oisc.regs[4][12] ),
    .B(net627));
 sg13g2_o21ai_1 _18825_ (.B1(_03238_),
    .Y(_01863_),
    .A1(net104),
    .A2(net490));
 sg13g2_nand2_1 _18826_ (.Y(_03239_),
    .A(\top_ihp.oisc.regs[4][13] ),
    .B(net627));
 sg13g2_o21ai_1 _18827_ (.B1(_03239_),
    .Y(_01864_),
    .A1(net91),
    .A2(net490));
 sg13g2_nand2_1 _18828_ (.Y(_03240_),
    .A(\top_ihp.oisc.regs[4][14] ),
    .B(net627));
 sg13g2_o21ai_1 _18829_ (.B1(_03240_),
    .Y(_01865_),
    .A1(net103),
    .A2(net490));
 sg13g2_nand2_1 _18830_ (.Y(_03241_),
    .A(\top_ihp.oisc.regs[4][15] ),
    .B(net627));
 sg13g2_o21ai_1 _18831_ (.B1(_03241_),
    .Y(_01866_),
    .A1(net98),
    .A2(net490));
 sg13g2_nand2_1 _18832_ (.Y(_03242_),
    .A(\top_ihp.oisc.regs[4][16] ),
    .B(net627));
 sg13g2_o21ai_1 _18833_ (.B1(_03242_),
    .Y(_01867_),
    .A1(net38),
    .A2(net490));
 sg13g2_buf_1 _18834_ (.A(net628),
    .X(_03243_));
 sg13g2_nand2_1 _18835_ (.Y(_03244_),
    .A(\top_ihp.oisc.regs[4][17] ),
    .B(net489));
 sg13g2_o21ai_1 _18836_ (.B1(_03244_),
    .Y(_01868_),
    .A1(_03016_),
    .A2(_03233_));
 sg13g2_nand2_1 _18837_ (.Y(_03245_),
    .A(\top_ihp.oisc.regs[4][18] ),
    .B(net489));
 sg13g2_o21ai_1 _18838_ (.B1(_03245_),
    .Y(_01869_),
    .A1(_03018_),
    .A2(_03233_));
 sg13g2_buf_1 _18839_ (.A(net628),
    .X(_03246_));
 sg13g2_nand2_1 _18840_ (.Y(_03247_),
    .A(\top_ihp.oisc.regs[4][19] ),
    .B(net489));
 sg13g2_o21ai_1 _18841_ (.B1(_03247_),
    .Y(_01870_),
    .A1(net88),
    .A2(net488));
 sg13g2_nand2_1 _18842_ (.Y(_03248_),
    .A(\top_ihp.oisc.regs[4][1] ),
    .B(net489));
 sg13g2_o21ai_1 _18843_ (.B1(_03248_),
    .Y(_01871_),
    .A1(net102),
    .A2(net488));
 sg13g2_nand2_1 _18844_ (.Y(_03249_),
    .A(\top_ihp.oisc.regs[4][20] ),
    .B(net489));
 sg13g2_o21ai_1 _18845_ (.B1(_03249_),
    .Y(_01872_),
    .A1(net324),
    .A2(net488));
 sg13g2_nand2_1 _18846_ (.Y(_03250_),
    .A(\top_ihp.oisc.regs[4][21] ),
    .B(net489));
 sg13g2_o21ai_1 _18847_ (.B1(_03250_),
    .Y(_01873_),
    .A1(net87),
    .A2(net488));
 sg13g2_nand2_1 _18848_ (.Y(_03251_),
    .A(\top_ihp.oisc.regs[4][22] ),
    .B(net489));
 sg13g2_o21ai_1 _18849_ (.B1(_03251_),
    .Y(_01874_),
    .A1(net101),
    .A2(net488));
 sg13g2_nand2_1 _18850_ (.Y(_03252_),
    .A(\top_ihp.oisc.regs[4][23] ),
    .B(_03243_));
 sg13g2_o21ai_1 _18851_ (.B1(_03252_),
    .Y(_01875_),
    .A1(net243),
    .A2(net488));
 sg13g2_nand2_1 _18852_ (.Y(_03253_),
    .A(\top_ihp.oisc.regs[4][24] ),
    .B(net489));
 sg13g2_o21ai_1 _18853_ (.B1(_03253_),
    .Y(_01876_),
    .A1(_03030_),
    .A2(_03246_));
 sg13g2_nand2_1 _18854_ (.Y(_03254_),
    .A(\top_ihp.oisc.regs[4][25] ),
    .B(_03243_));
 sg13g2_o21ai_1 _18855_ (.B1(_03254_),
    .Y(_01877_),
    .A1(_02892_),
    .A2(net488));
 sg13g2_buf_8 _18856_ (.A(net628),
    .X(_03255_));
 sg13g2_nand2_1 _18857_ (.Y(_03256_),
    .A(\top_ihp.oisc.regs[4][26] ),
    .B(net487));
 sg13g2_o21ai_1 _18858_ (.B1(_03256_),
    .Y(_01878_),
    .A1(net37),
    .A2(_03246_));
 sg13g2_nand2_1 _18859_ (.Y(_03257_),
    .A(\top_ihp.oisc.regs[4][27] ),
    .B(net487));
 sg13g2_o21ai_1 _18860_ (.B1(_03257_),
    .Y(_01879_),
    .A1(net85),
    .A2(net488));
 sg13g2_buf_1 _18861_ (.A(net628),
    .X(_03258_));
 sg13g2_nand2_1 _18862_ (.Y(_03259_),
    .A(\top_ihp.oisc.regs[4][28] ),
    .B(net487));
 sg13g2_o21ai_1 _18863_ (.B1(_03259_),
    .Y(_01880_),
    .A1(net241),
    .A2(net486));
 sg13g2_nand2_1 _18864_ (.Y(_03260_),
    .A(\top_ihp.oisc.regs[4][29] ),
    .B(_03255_));
 sg13g2_o21ai_1 _18865_ (.B1(_03260_),
    .Y(_01881_),
    .A1(net84),
    .A2(_03258_));
 sg13g2_nand2_1 _18866_ (.Y(_03261_),
    .A(\top_ihp.oisc.regs[4][2] ),
    .B(net487));
 sg13g2_o21ai_1 _18867_ (.B1(_03261_),
    .Y(_01882_),
    .A1(net32),
    .A2(net486));
 sg13g2_nand2_1 _18868_ (.Y(_03262_),
    .A(\top_ihp.oisc.regs[4][30] ),
    .B(net487));
 sg13g2_o21ai_1 _18869_ (.B1(_03262_),
    .Y(_01883_),
    .A1(_03091_),
    .A2(net486));
 sg13g2_nand2_1 _18870_ (.Y(_03263_),
    .A(\top_ihp.oisc.regs[4][31] ),
    .B(net487));
 sg13g2_o21ai_1 _18871_ (.B1(_03263_),
    .Y(_01884_),
    .A1(net52),
    .A2(net486));
 sg13g2_nand2_1 _18872_ (.Y(_03264_),
    .A(\top_ihp.oisc.regs[4][3] ),
    .B(net487));
 sg13g2_o21ai_1 _18873_ (.B1(_03264_),
    .Y(_01885_),
    .A1(net30),
    .A2(net486));
 sg13g2_nand2_1 _18874_ (.Y(_03265_),
    .A(\top_ihp.oisc.regs[4][4] ),
    .B(net487));
 sg13g2_o21ai_1 _18875_ (.B1(_03265_),
    .Y(_01886_),
    .A1(net29),
    .A2(net486));
 sg13g2_nand2_1 _18876_ (.Y(_03266_),
    .A(\top_ihp.oisc.regs[4][5] ),
    .B(_03255_));
 sg13g2_o21ai_1 _18877_ (.B1(_03266_),
    .Y(_01887_),
    .A1(net36),
    .A2(_03258_));
 sg13g2_nand2_1 _18878_ (.Y(_03267_),
    .A(\top_ihp.oisc.regs[4][6] ),
    .B(net628));
 sg13g2_o21ai_1 _18879_ (.B1(_03267_),
    .Y(_01888_),
    .A1(net35),
    .A2(net486));
 sg13g2_nand2_1 _18880_ (.Y(_03268_),
    .A(\top_ihp.oisc.regs[4][7] ),
    .B(net628));
 sg13g2_o21ai_1 _18881_ (.B1(_03268_),
    .Y(_01889_),
    .A1(net139),
    .A2(net486));
 sg13g2_nand2_1 _18882_ (.Y(_03269_),
    .A(\top_ihp.oisc.regs[4][8] ),
    .B(_03232_));
 sg13g2_o21ai_1 _18883_ (.B1(_03269_),
    .Y(_01890_),
    .A1(net83),
    .A2(_03234_));
 sg13g2_nand2_1 _18884_ (.Y(_03270_),
    .A(\top_ihp.oisc.regs[4][9] ),
    .B(net628));
 sg13g2_o21ai_1 _18885_ (.B1(_03270_),
    .Y(_01891_),
    .A1(net34),
    .A2(_03234_));
 sg13g2_nand3_1 _18886_ (.B(net741),
    .C(_03146_),
    .A(_09725_),
    .Y(_03271_));
 sg13g2_buf_1 _18887_ (.A(_03271_),
    .X(_03272_));
 sg13g2_buf_8 _18888_ (.A(_03272_),
    .X(_03273_));
 sg13g2_buf_1 _18889_ (.A(net626),
    .X(_03274_));
 sg13g2_buf_1 _18890_ (.A(_03272_),
    .X(_03275_));
 sg13g2_nand2_1 _18891_ (.Y(_03276_),
    .A(\top_ihp.oisc.regs[50][0] ),
    .B(net625));
 sg13g2_o21ai_1 _18892_ (.B1(_03276_),
    .Y(_01892_),
    .A1(net82),
    .A2(net485));
 sg13g2_nand2_1 _18893_ (.Y(_03277_),
    .A(\top_ihp.oisc.regs[50][10] ),
    .B(net625));
 sg13g2_o21ai_1 _18894_ (.B1(_03277_),
    .Y(_01893_),
    .A1(net39),
    .A2(net485));
 sg13g2_nand2_1 _18895_ (.Y(_03278_),
    .A(\top_ihp.oisc.regs[50][11] ),
    .B(_03275_));
 sg13g2_o21ai_1 _18896_ (.B1(_03278_),
    .Y(_01894_),
    .A1(net33),
    .A2(net485));
 sg13g2_nand2_1 _18897_ (.Y(_03279_),
    .A(\top_ihp.oisc.regs[50][12] ),
    .B(net625));
 sg13g2_o21ai_1 _18898_ (.B1(_03279_),
    .Y(_01895_),
    .A1(net104),
    .A2(net485));
 sg13g2_nand2_1 _18899_ (.Y(_03280_),
    .A(\top_ihp.oisc.regs[50][13] ),
    .B(_03275_));
 sg13g2_o21ai_1 _18900_ (.B1(_03280_),
    .Y(_01896_),
    .A1(net91),
    .A2(net485));
 sg13g2_nand2_1 _18901_ (.Y(_03281_),
    .A(\top_ihp.oisc.regs[50][14] ),
    .B(net625));
 sg13g2_o21ai_1 _18902_ (.B1(_03281_),
    .Y(_01897_),
    .A1(net103),
    .A2(net485));
 sg13g2_nand2_1 _18903_ (.Y(_03282_),
    .A(\top_ihp.oisc.regs[50][15] ),
    .B(net625));
 sg13g2_o21ai_1 _18904_ (.B1(_03282_),
    .Y(_01898_),
    .A1(net98),
    .A2(net485));
 sg13g2_nand2_1 _18905_ (.Y(_03283_),
    .A(\top_ihp.oisc.regs[50][16] ),
    .B(net625));
 sg13g2_o21ai_1 _18906_ (.B1(_03283_),
    .Y(_01899_),
    .A1(net38),
    .A2(net485));
 sg13g2_buf_1 _18907_ (.A(_03273_),
    .X(_03284_));
 sg13g2_nand2_1 _18908_ (.Y(_03285_),
    .A(\top_ihp.oisc.regs[50][17] ),
    .B(_03284_));
 sg13g2_o21ai_1 _18909_ (.B1(_03285_),
    .Y(_01900_),
    .A1(net90),
    .A2(_03274_));
 sg13g2_nand2_1 _18910_ (.Y(_03286_),
    .A(\top_ihp.oisc.regs[50][18] ),
    .B(_03284_));
 sg13g2_o21ai_1 _18911_ (.B1(_03286_),
    .Y(_01901_),
    .A1(net89),
    .A2(_03274_));
 sg13g2_buf_1 _18912_ (.A(net626),
    .X(_03287_));
 sg13g2_nand2_1 _18913_ (.Y(_03288_),
    .A(\top_ihp.oisc.regs[50][19] ),
    .B(net484));
 sg13g2_o21ai_1 _18914_ (.B1(_03288_),
    .Y(_01902_),
    .A1(net88),
    .A2(net483));
 sg13g2_nand2_1 _18915_ (.Y(_03289_),
    .A(\top_ihp.oisc.regs[50][1] ),
    .B(net484));
 sg13g2_o21ai_1 _18916_ (.B1(_03289_),
    .Y(_01903_),
    .A1(net102),
    .A2(net483));
 sg13g2_nand2_1 _18917_ (.Y(_03290_),
    .A(\top_ihp.oisc.regs[50][20] ),
    .B(net484));
 sg13g2_o21ai_1 _18918_ (.B1(_03290_),
    .Y(_01904_),
    .A1(_10153_),
    .A2(net483));
 sg13g2_nand2_1 _18919_ (.Y(_03291_),
    .A(\top_ihp.oisc.regs[50][21] ),
    .B(net484));
 sg13g2_o21ai_1 _18920_ (.B1(_03291_),
    .Y(_01905_),
    .A1(net87),
    .A2(net483));
 sg13g2_nand2_1 _18921_ (.Y(_03292_),
    .A(\top_ihp.oisc.regs[50][22] ),
    .B(net484));
 sg13g2_o21ai_1 _18922_ (.B1(_03292_),
    .Y(_01906_),
    .A1(net101),
    .A2(net483));
 sg13g2_nand2_1 _18923_ (.Y(_03293_),
    .A(\top_ihp.oisc.regs[50][23] ),
    .B(net484));
 sg13g2_o21ai_1 _18924_ (.B1(_03293_),
    .Y(_01907_),
    .A1(net243),
    .A2(_03287_));
 sg13g2_nand2_1 _18925_ (.Y(_03294_),
    .A(\top_ihp.oisc.regs[50][24] ),
    .B(net484));
 sg13g2_o21ai_1 _18926_ (.B1(_03294_),
    .Y(_01908_),
    .A1(net86),
    .A2(_03287_));
 sg13g2_nand2_1 _18927_ (.Y(_03295_),
    .A(\top_ihp.oisc.regs[50][25] ),
    .B(net484));
 sg13g2_o21ai_1 _18928_ (.B1(_03295_),
    .Y(_01909_),
    .A1(net97),
    .A2(net483));
 sg13g2_buf_1 _18929_ (.A(net626),
    .X(_03296_));
 sg13g2_nand2_1 _18930_ (.Y(_03297_),
    .A(\top_ihp.oisc.regs[50][26] ),
    .B(net482));
 sg13g2_o21ai_1 _18931_ (.B1(_03297_),
    .Y(_01910_),
    .A1(net37),
    .A2(net483));
 sg13g2_nand2_1 _18932_ (.Y(_03298_),
    .A(\top_ihp.oisc.regs[50][27] ),
    .B(net482));
 sg13g2_o21ai_1 _18933_ (.B1(_03298_),
    .Y(_01911_),
    .A1(net85),
    .A2(net483));
 sg13g2_buf_1 _18934_ (.A(net626),
    .X(_03299_));
 sg13g2_nand2_1 _18935_ (.Y(_03300_),
    .A(\top_ihp.oisc.regs[50][28] ),
    .B(net482));
 sg13g2_o21ai_1 _18936_ (.B1(_03300_),
    .Y(_01912_),
    .A1(net241),
    .A2(net481));
 sg13g2_nand2_1 _18937_ (.Y(_03301_),
    .A(\top_ihp.oisc.regs[50][29] ),
    .B(net482));
 sg13g2_o21ai_1 _18938_ (.B1(_03301_),
    .Y(_01913_),
    .A1(net84),
    .A2(net481));
 sg13g2_nand2_1 _18939_ (.Y(_03302_),
    .A(\top_ihp.oisc.regs[50][2] ),
    .B(net482));
 sg13g2_o21ai_1 _18940_ (.B1(_03302_),
    .Y(_01914_),
    .A1(net32),
    .A2(net481));
 sg13g2_nand2_1 _18941_ (.Y(_03303_),
    .A(\top_ihp.oisc.regs[50][30] ),
    .B(net482));
 sg13g2_o21ai_1 _18942_ (.B1(_03303_),
    .Y(_01915_),
    .A1(net31),
    .A2(net481));
 sg13g2_nand2_1 _18943_ (.Y(_03304_),
    .A(\top_ihp.oisc.regs[50][31] ),
    .B(net482));
 sg13g2_o21ai_1 _18944_ (.B1(_03304_),
    .Y(_01916_),
    .A1(_10349_),
    .A2(net481));
 sg13g2_nand2_1 _18945_ (.Y(_03305_),
    .A(\top_ihp.oisc.regs[50][3] ),
    .B(_03296_));
 sg13g2_o21ai_1 _18946_ (.B1(_03305_),
    .Y(_01917_),
    .A1(net30),
    .A2(_03299_));
 sg13g2_nand2_1 _18947_ (.Y(_03306_),
    .A(\top_ihp.oisc.regs[50][4] ),
    .B(net482));
 sg13g2_o21ai_1 _18948_ (.B1(_03306_),
    .Y(_01918_),
    .A1(net29),
    .A2(net481));
 sg13g2_nand2_1 _18949_ (.Y(_03307_),
    .A(\top_ihp.oisc.regs[50][5] ),
    .B(_03296_));
 sg13g2_o21ai_1 _18950_ (.B1(_03307_),
    .Y(_01919_),
    .A1(net36),
    .A2(_03299_));
 sg13g2_nand2_1 _18951_ (.Y(_03308_),
    .A(\top_ihp.oisc.regs[50][6] ),
    .B(net626));
 sg13g2_o21ai_1 _18952_ (.B1(_03308_),
    .Y(_01920_),
    .A1(net35),
    .A2(net481));
 sg13g2_nand2_1 _18953_ (.Y(_03309_),
    .A(\top_ihp.oisc.regs[50][7] ),
    .B(net626));
 sg13g2_o21ai_1 _18954_ (.B1(_03309_),
    .Y(_01921_),
    .A1(_10484_),
    .A2(net481));
 sg13g2_nand2_1 _18955_ (.Y(_03310_),
    .A(\top_ihp.oisc.regs[50][8] ),
    .B(net626));
 sg13g2_o21ai_1 _18956_ (.B1(_03310_),
    .Y(_01922_),
    .A1(net83),
    .A2(net625));
 sg13g2_nand2_1 _18957_ (.Y(_03311_),
    .A(\top_ihp.oisc.regs[50][9] ),
    .B(net626));
 sg13g2_o21ai_1 _18958_ (.B1(_03311_),
    .Y(_01923_),
    .A1(net34),
    .A2(net625));
 sg13g2_and2_1 _18959_ (.A(net785),
    .B(_03146_),
    .X(_03312_));
 sg13g2_buf_1 _18960_ (.A(_03312_),
    .X(_03313_));
 sg13g2_nand2_1 _18961_ (.Y(_03314_),
    .A(_09726_),
    .B(_03313_));
 sg13g2_buf_1 _18962_ (.A(_03314_),
    .X(_03315_));
 sg13g2_buf_1 _18963_ (.A(net701),
    .X(_03316_));
 sg13g2_buf_1 _18964_ (.A(_03314_),
    .X(_03317_));
 sg13g2_nand2_1 _18965_ (.Y(_03318_),
    .A(\top_ihp.oisc.regs[51][0] ),
    .B(net700));
 sg13g2_o21ai_1 _18966_ (.B1(_03318_),
    .Y(_01924_),
    .A1(_03056_),
    .A2(net624));
 sg13g2_nand2_1 _18967_ (.Y(_03319_),
    .A(\top_ihp.oisc.regs[51][10] ),
    .B(net700));
 sg13g2_o21ai_1 _18968_ (.B1(_03319_),
    .Y(_01925_),
    .A1(net39),
    .A2(net624));
 sg13g2_nand2_1 _18969_ (.Y(_03320_),
    .A(\top_ihp.oisc.regs[51][11] ),
    .B(net700));
 sg13g2_o21ai_1 _18970_ (.B1(_03320_),
    .Y(_01926_),
    .A1(net33),
    .A2(net624));
 sg13g2_nand2_1 _18971_ (.Y(_03321_),
    .A(\top_ihp.oisc.regs[51][12] ),
    .B(net700));
 sg13g2_o21ai_1 _18972_ (.B1(_03321_),
    .Y(_01927_),
    .A1(_11158_),
    .A2(net624));
 sg13g2_nand2_1 _18973_ (.Y(_03322_),
    .A(\top_ihp.oisc.regs[51][13] ),
    .B(_03317_));
 sg13g2_o21ai_1 _18974_ (.B1(_03322_),
    .Y(_01928_),
    .A1(_03010_),
    .A2(net624));
 sg13g2_nand2_1 _18975_ (.Y(_03323_),
    .A(\top_ihp.oisc.regs[51][14] ),
    .B(net700));
 sg13g2_o21ai_1 _18976_ (.B1(_03323_),
    .Y(_01929_),
    .A1(net103),
    .A2(net624));
 sg13g2_nand2_1 _18977_ (.Y(_03324_),
    .A(\top_ihp.oisc.regs[51][15] ),
    .B(net700));
 sg13g2_o21ai_1 _18978_ (.B1(_03324_),
    .Y(_01930_),
    .A1(net98),
    .A2(net624));
 sg13g2_nand2_1 _18979_ (.Y(_03325_),
    .A(\top_ihp.oisc.regs[51][16] ),
    .B(_03317_));
 sg13g2_o21ai_1 _18980_ (.B1(_03325_),
    .Y(_01931_),
    .A1(_03014_),
    .A2(net624));
 sg13g2_buf_1 _18981_ (.A(net701),
    .X(_03326_));
 sg13g2_nand2_1 _18982_ (.Y(_03327_),
    .A(\top_ihp.oisc.regs[51][17] ),
    .B(_03326_));
 sg13g2_o21ai_1 _18983_ (.B1(_03327_),
    .Y(_01932_),
    .A1(net90),
    .A2(_03316_));
 sg13g2_nand2_1 _18984_ (.Y(_03328_),
    .A(\top_ihp.oisc.regs[51][18] ),
    .B(_03326_));
 sg13g2_o21ai_1 _18985_ (.B1(_03328_),
    .Y(_01933_),
    .A1(_03018_),
    .A2(_03316_));
 sg13g2_buf_1 _18986_ (.A(net701),
    .X(_03329_));
 sg13g2_nand2_1 _18987_ (.Y(_03330_),
    .A(\top_ihp.oisc.regs[51][19] ),
    .B(net623));
 sg13g2_o21ai_1 _18988_ (.B1(_03330_),
    .Y(_01934_),
    .A1(net88),
    .A2(net622));
 sg13g2_nand2_1 _18989_ (.Y(_03331_),
    .A(\top_ihp.oisc.regs[51][1] ),
    .B(net623));
 sg13g2_o21ai_1 _18990_ (.B1(_03331_),
    .Y(_01935_),
    .A1(_11170_),
    .A2(net622));
 sg13g2_nand2_1 _18991_ (.Y(_03332_),
    .A(\top_ihp.oisc.regs[51][20] ),
    .B(net623));
 sg13g2_o21ai_1 _18992_ (.B1(_03332_),
    .Y(_01936_),
    .A1(net636),
    .A2(net622));
 sg13g2_nand2_1 _18993_ (.Y(_03333_),
    .A(\top_ihp.oisc.regs[51][21] ),
    .B(net623));
 sg13g2_o21ai_1 _18994_ (.B1(_03333_),
    .Y(_01937_),
    .A1(net87),
    .A2(_03329_));
 sg13g2_nand2_1 _18995_ (.Y(_03334_),
    .A(\top_ihp.oisc.regs[51][22] ),
    .B(net623));
 sg13g2_o21ai_1 _18996_ (.B1(_03334_),
    .Y(_01938_),
    .A1(net101),
    .A2(net622));
 sg13g2_nand2_1 _18997_ (.Y(_03335_),
    .A(\top_ihp.oisc.regs[51][23] ),
    .B(net623));
 sg13g2_o21ai_1 _18998_ (.B1(_03335_),
    .Y(_01939_),
    .A1(_03028_),
    .A2(_03329_));
 sg13g2_nand2_1 _18999_ (.Y(_03336_),
    .A(\top_ihp.oisc.regs[51][24] ),
    .B(net623));
 sg13g2_o21ai_1 _19000_ (.B1(_03336_),
    .Y(_01940_),
    .A1(net86),
    .A2(net622));
 sg13g2_nand2_1 _19001_ (.Y(_03337_),
    .A(\top_ihp.oisc.regs[51][25] ),
    .B(net623));
 sg13g2_o21ai_1 _19002_ (.B1(_03337_),
    .Y(_01941_),
    .A1(net97),
    .A2(net622));
 sg13g2_buf_1 _19003_ (.A(net701),
    .X(_03338_));
 sg13g2_nand2_1 _19004_ (.Y(_03339_),
    .A(\top_ihp.oisc.regs[51][26] ),
    .B(net621));
 sg13g2_o21ai_1 _19005_ (.B1(_03339_),
    .Y(_01942_),
    .A1(net37),
    .A2(net622));
 sg13g2_nand2_1 _19006_ (.Y(_03340_),
    .A(\top_ihp.oisc.regs[51][27] ),
    .B(net621));
 sg13g2_o21ai_1 _19007_ (.B1(_03340_),
    .Y(_01943_),
    .A1(net85),
    .A2(net622));
 sg13g2_buf_1 _19008_ (.A(net701),
    .X(_03341_));
 sg13g2_nand2_1 _19009_ (.Y(_03342_),
    .A(\top_ihp.oisc.regs[51][28] ),
    .B(net621));
 sg13g2_o21ai_1 _19010_ (.B1(_03342_),
    .Y(_01944_),
    .A1(net241),
    .A2(net620));
 sg13g2_nand2_1 _19011_ (.Y(_03343_),
    .A(\top_ihp.oisc.regs[51][29] ),
    .B(net621));
 sg13g2_o21ai_1 _19012_ (.B1(_03343_),
    .Y(_01945_),
    .A1(_03040_),
    .A2(net620));
 sg13g2_nand2_1 _19013_ (.Y(_03344_),
    .A(\top_ihp.oisc.regs[51][2] ),
    .B(net621));
 sg13g2_o21ai_1 _19014_ (.B1(_03344_),
    .Y(_01946_),
    .A1(net32),
    .A2(net620));
 sg13g2_nand2_1 _19015_ (.Y(_03345_),
    .A(\top_ihp.oisc.regs[51][30] ),
    .B(net621));
 sg13g2_o21ai_1 _19016_ (.B1(_03345_),
    .Y(_01947_),
    .A1(net31),
    .A2(_03341_));
 sg13g2_nand2_1 _19017_ (.Y(_03346_),
    .A(\top_ihp.oisc.regs[51][31] ),
    .B(net621));
 sg13g2_o21ai_1 _19018_ (.B1(_03346_),
    .Y(_01948_),
    .A1(net251),
    .A2(net620));
 sg13g2_nand2_1 _19019_ (.Y(_03347_),
    .A(\top_ihp.oisc.regs[51][3] ),
    .B(net621));
 sg13g2_o21ai_1 _19020_ (.B1(_03347_),
    .Y(_01949_),
    .A1(net30),
    .A2(net620));
 sg13g2_nand2_1 _19021_ (.Y(_03348_),
    .A(\top_ihp.oisc.regs[51][4] ),
    .B(_03338_));
 sg13g2_o21ai_1 _19022_ (.B1(_03348_),
    .Y(_01950_),
    .A1(net29),
    .A2(_03341_));
 sg13g2_nand2_1 _19023_ (.Y(_03349_),
    .A(\top_ihp.oisc.regs[51][5] ),
    .B(_03338_));
 sg13g2_o21ai_1 _19024_ (.B1(_03349_),
    .Y(_01951_),
    .A1(net36),
    .A2(net620));
 sg13g2_nand2_1 _19025_ (.Y(_03350_),
    .A(\top_ihp.oisc.regs[51][6] ),
    .B(net701));
 sg13g2_o21ai_1 _19026_ (.B1(_03350_),
    .Y(_01952_),
    .A1(_03049_),
    .A2(net620));
 sg13g2_nand2_1 _19027_ (.Y(_03351_),
    .A(\top_ihp.oisc.regs[51][7] ),
    .B(net701));
 sg13g2_o21ai_1 _19028_ (.B1(_03351_),
    .Y(_01953_),
    .A1(net501),
    .A2(net620));
 sg13g2_nand2_1 _19029_ (.Y(_03352_),
    .A(\top_ihp.oisc.regs[51][8] ),
    .B(_03315_));
 sg13g2_o21ai_1 _19030_ (.B1(_03352_),
    .Y(_01954_),
    .A1(_03052_),
    .A2(net700));
 sg13g2_nand2_1 _19031_ (.Y(_03353_),
    .A(\top_ihp.oisc.regs[51][9] ),
    .B(net701));
 sg13g2_o21ai_1 _19032_ (.B1(_03353_),
    .Y(_01955_),
    .A1(_03054_),
    .A2(net700));
 sg13g2_nand2_1 _19033_ (.Y(_03354_),
    .A(_10988_),
    .B(_03148_));
 sg13g2_buf_1 _19034_ (.A(_03354_),
    .X(_03355_));
 sg13g2_buf_1 _19035_ (.A(net619),
    .X(_03356_));
 sg13g2_buf_1 _19036_ (.A(_03354_),
    .X(_03357_));
 sg13g2_nand2_1 _19037_ (.Y(_03358_),
    .A(\top_ihp.oisc.regs[52][0] ),
    .B(_03357_));
 sg13g2_o21ai_1 _19038_ (.B1(_03358_),
    .Y(_01956_),
    .A1(net82),
    .A2(_03356_));
 sg13g2_nand2_1 _19039_ (.Y(_03359_),
    .A(\top_ihp.oisc.regs[52][10] ),
    .B(net618));
 sg13g2_o21ai_1 _19040_ (.B1(_03359_),
    .Y(_01957_),
    .A1(_03004_),
    .A2(net480));
 sg13g2_nand2_1 _19041_ (.Y(_03360_),
    .A(\top_ihp.oisc.regs[52][11] ),
    .B(net618));
 sg13g2_o21ai_1 _19042_ (.B1(_03360_),
    .Y(_01958_),
    .A1(net33),
    .A2(net480));
 sg13g2_nand2_1 _19043_ (.Y(_03361_),
    .A(\top_ihp.oisc.regs[52][12] ),
    .B(net618));
 sg13g2_o21ai_1 _19044_ (.B1(_03361_),
    .Y(_01959_),
    .A1(net104),
    .A2(net480));
 sg13g2_nand2_1 _19045_ (.Y(_03362_),
    .A(\top_ihp.oisc.regs[52][13] ),
    .B(_03357_));
 sg13g2_o21ai_1 _19046_ (.B1(_03362_),
    .Y(_01960_),
    .A1(_03010_),
    .A2(net480));
 sg13g2_nand2_1 _19047_ (.Y(_03363_),
    .A(\top_ihp.oisc.regs[52][14] ),
    .B(net618));
 sg13g2_o21ai_1 _19048_ (.B1(_03363_),
    .Y(_01961_),
    .A1(net103),
    .A2(net480));
 sg13g2_nand2_1 _19049_ (.Y(_03364_),
    .A(\top_ihp.oisc.regs[52][15] ),
    .B(net618));
 sg13g2_o21ai_1 _19050_ (.B1(_03364_),
    .Y(_01962_),
    .A1(net98),
    .A2(net480));
 sg13g2_nand2_1 _19051_ (.Y(_03365_),
    .A(\top_ihp.oisc.regs[52][16] ),
    .B(net618));
 sg13g2_o21ai_1 _19052_ (.B1(_03365_),
    .Y(_01963_),
    .A1(_03014_),
    .A2(net480));
 sg13g2_buf_2 _19053_ (.A(net619),
    .X(_03366_));
 sg13g2_nand2_1 _19054_ (.Y(_03367_),
    .A(\top_ihp.oisc.regs[52][17] ),
    .B(net479));
 sg13g2_o21ai_1 _19055_ (.B1(_03367_),
    .Y(_01964_),
    .A1(net90),
    .A2(net480));
 sg13g2_nand2_1 _19056_ (.Y(_03368_),
    .A(\top_ihp.oisc.regs[52][18] ),
    .B(net479));
 sg13g2_o21ai_1 _19057_ (.B1(_03368_),
    .Y(_01965_),
    .A1(net89),
    .A2(_03356_));
 sg13g2_buf_2 _19058_ (.A(net619),
    .X(_03369_));
 sg13g2_nand2_1 _19059_ (.Y(_03370_),
    .A(\top_ihp.oisc.regs[52][19] ),
    .B(net479));
 sg13g2_o21ai_1 _19060_ (.B1(_03370_),
    .Y(_01966_),
    .A1(_03020_),
    .A2(net478));
 sg13g2_nand2_1 _19061_ (.Y(_03371_),
    .A(\top_ihp.oisc.regs[52][1] ),
    .B(net479));
 sg13g2_o21ai_1 _19062_ (.B1(_03371_),
    .Y(_01967_),
    .A1(net102),
    .A2(net478));
 sg13g2_nand2_1 _19063_ (.Y(_03372_),
    .A(\top_ihp.oisc.regs[52][20] ),
    .B(net479));
 sg13g2_o21ai_1 _19064_ (.B1(_03372_),
    .Y(_01968_),
    .A1(net636),
    .A2(net478));
 sg13g2_nand2_1 _19065_ (.Y(_03373_),
    .A(\top_ihp.oisc.regs[52][21] ),
    .B(_03366_));
 sg13g2_o21ai_1 _19066_ (.B1(_03373_),
    .Y(_01969_),
    .A1(net87),
    .A2(net478));
 sg13g2_nand2_1 _19067_ (.Y(_03374_),
    .A(\top_ihp.oisc.regs[52][22] ),
    .B(net479));
 sg13g2_o21ai_1 _19068_ (.B1(_03374_),
    .Y(_01970_),
    .A1(_11174_),
    .A2(net478));
 sg13g2_nand2_1 _19069_ (.Y(_03375_),
    .A(\top_ihp.oisc.regs[52][23] ),
    .B(net479));
 sg13g2_o21ai_1 _19070_ (.B1(_03375_),
    .Y(_01971_),
    .A1(net243),
    .A2(net478));
 sg13g2_nand2_1 _19071_ (.Y(_03376_),
    .A(\top_ihp.oisc.regs[52][24] ),
    .B(_03366_));
 sg13g2_o21ai_1 _19072_ (.B1(_03376_),
    .Y(_01972_),
    .A1(net86),
    .A2(_03369_));
 sg13g2_nand2_1 _19073_ (.Y(_03377_),
    .A(\top_ihp.oisc.regs[52][25] ),
    .B(net479));
 sg13g2_o21ai_1 _19074_ (.B1(_03377_),
    .Y(_01973_),
    .A1(net97),
    .A2(net478));
 sg13g2_buf_2 _19075_ (.A(net619),
    .X(_03378_));
 sg13g2_nand2_1 _19076_ (.Y(_03379_),
    .A(\top_ihp.oisc.regs[52][26] ),
    .B(net477));
 sg13g2_o21ai_1 _19077_ (.B1(_03379_),
    .Y(_01974_),
    .A1(_03034_),
    .A2(_03369_));
 sg13g2_nand2_1 _19078_ (.Y(_03380_),
    .A(\top_ihp.oisc.regs[52][27] ),
    .B(_03378_));
 sg13g2_o21ai_1 _19079_ (.B1(_03380_),
    .Y(_01975_),
    .A1(_03036_),
    .A2(net478));
 sg13g2_buf_1 _19080_ (.A(net619),
    .X(_03381_));
 sg13g2_nand2_1 _19081_ (.Y(_03382_),
    .A(\top_ihp.oisc.regs[52][28] ),
    .B(net477));
 sg13g2_o21ai_1 _19082_ (.B1(_03382_),
    .Y(_01976_),
    .A1(_03038_),
    .A2(net476));
 sg13g2_nand2_1 _19083_ (.Y(_03383_),
    .A(\top_ihp.oisc.regs[52][29] ),
    .B(net477));
 sg13g2_o21ai_1 _19084_ (.B1(_03383_),
    .Y(_01977_),
    .A1(net84),
    .A2(net476));
 sg13g2_nand2_1 _19085_ (.Y(_03384_),
    .A(\top_ihp.oisc.regs[52][2] ),
    .B(net477));
 sg13g2_o21ai_1 _19086_ (.B1(_03384_),
    .Y(_01978_),
    .A1(net32),
    .A2(net476));
 sg13g2_nand2_1 _19087_ (.Y(_03385_),
    .A(\top_ihp.oisc.regs[52][30] ),
    .B(net477));
 sg13g2_o21ai_1 _19088_ (.B1(_03385_),
    .Y(_01979_),
    .A1(net31),
    .A2(net476));
 sg13g2_nand2_1 _19089_ (.Y(_03386_),
    .A(\top_ihp.oisc.regs[52][31] ),
    .B(net477));
 sg13g2_o21ai_1 _19090_ (.B1(_03386_),
    .Y(_01980_),
    .A1(net251),
    .A2(net476));
 sg13g2_nand2_1 _19091_ (.Y(_03387_),
    .A(\top_ihp.oisc.regs[52][3] ),
    .B(net477));
 sg13g2_o21ai_1 _19092_ (.B1(_03387_),
    .Y(_01981_),
    .A1(net30),
    .A2(_03381_));
 sg13g2_nand2_1 _19093_ (.Y(_03388_),
    .A(\top_ihp.oisc.regs[52][4] ),
    .B(_03378_));
 sg13g2_o21ai_1 _19094_ (.B1(_03388_),
    .Y(_01982_),
    .A1(net29),
    .A2(_03381_));
 sg13g2_nand2_1 _19095_ (.Y(_03389_),
    .A(\top_ihp.oisc.regs[52][5] ),
    .B(net477));
 sg13g2_o21ai_1 _19096_ (.B1(_03389_),
    .Y(_01983_),
    .A1(_03047_),
    .A2(net476));
 sg13g2_nand2_1 _19097_ (.Y(_03390_),
    .A(\top_ihp.oisc.regs[52][6] ),
    .B(net619));
 sg13g2_o21ai_1 _19098_ (.B1(_03390_),
    .Y(_01984_),
    .A1(net35),
    .A2(net476));
 sg13g2_nand2_1 _19099_ (.Y(_03391_),
    .A(\top_ihp.oisc.regs[52][7] ),
    .B(_03355_));
 sg13g2_o21ai_1 _19100_ (.B1(_03391_),
    .Y(_01985_),
    .A1(net501),
    .A2(net476));
 sg13g2_nand2_1 _19101_ (.Y(_03392_),
    .A(\top_ihp.oisc.regs[52][8] ),
    .B(net619));
 sg13g2_o21ai_1 _19102_ (.B1(_03392_),
    .Y(_01986_),
    .A1(net83),
    .A2(net618));
 sg13g2_nand2_1 _19103_ (.Y(_03393_),
    .A(\top_ihp.oisc.regs[52][9] ),
    .B(net619));
 sg13g2_o21ai_1 _19104_ (.B1(_03393_),
    .Y(_01987_),
    .A1(net34),
    .A2(net618));
 sg13g2_or2_1 _19105_ (.X(_03394_),
    .B(_03189_),
    .A(_10964_));
 sg13g2_buf_1 _19106_ (.A(_03394_),
    .X(_03395_));
 sg13g2_buf_1 _19107_ (.A(_03395_),
    .X(_03396_));
 sg13g2_buf_1 _19108_ (.A(net699),
    .X(_03397_));
 sg13g2_buf_1 _19109_ (.A(_03395_),
    .X(_03398_));
 sg13g2_nand2_1 _19110_ (.Y(_03399_),
    .A(\top_ihp.oisc.regs[53][0] ),
    .B(_03398_));
 sg13g2_o21ai_1 _19111_ (.B1(_03399_),
    .Y(_01988_),
    .A1(net82),
    .A2(net617));
 sg13g2_nand2_1 _19112_ (.Y(_03400_),
    .A(\top_ihp.oisc.regs[53][10] ),
    .B(net698));
 sg13g2_o21ai_1 _19113_ (.B1(_03400_),
    .Y(_01989_),
    .A1(_03004_),
    .A2(net617));
 sg13g2_nand2_1 _19114_ (.Y(_03401_),
    .A(\top_ihp.oisc.regs[53][11] ),
    .B(_03398_));
 sg13g2_o21ai_1 _19115_ (.B1(_03401_),
    .Y(_01990_),
    .A1(net33),
    .A2(_03397_));
 sg13g2_nand2_1 _19116_ (.Y(_03402_),
    .A(\top_ihp.oisc.regs[53][12] ),
    .B(net698));
 sg13g2_o21ai_1 _19117_ (.B1(_03402_),
    .Y(_01991_),
    .A1(_11158_),
    .A2(net617));
 sg13g2_nand2_1 _19118_ (.Y(_03403_),
    .A(\top_ihp.oisc.regs[53][13] ),
    .B(net698));
 sg13g2_o21ai_1 _19119_ (.B1(_03403_),
    .Y(_01992_),
    .A1(net91),
    .A2(net617));
 sg13g2_nand2_1 _19120_ (.Y(_03404_),
    .A(\top_ihp.oisc.regs[53][14] ),
    .B(net698));
 sg13g2_o21ai_1 _19121_ (.B1(_03404_),
    .Y(_01993_),
    .A1(_11161_),
    .A2(net617));
 sg13g2_nand2_1 _19122_ (.Y(_03405_),
    .A(\top_ihp.oisc.regs[53][15] ),
    .B(net698));
 sg13g2_o21ai_1 _19123_ (.B1(_03405_),
    .Y(_01994_),
    .A1(net98),
    .A2(net617));
 sg13g2_nand2_1 _19124_ (.Y(_03406_),
    .A(\top_ihp.oisc.regs[53][16] ),
    .B(net698));
 sg13g2_o21ai_1 _19125_ (.B1(_03406_),
    .Y(_01995_),
    .A1(net38),
    .A2(net617));
 sg13g2_buf_1 _19126_ (.A(net699),
    .X(_03407_));
 sg13g2_nand2_1 _19127_ (.Y(_03408_),
    .A(\top_ihp.oisc.regs[53][17] ),
    .B(net616));
 sg13g2_o21ai_1 _19128_ (.B1(_03408_),
    .Y(_01996_),
    .A1(_03016_),
    .A2(_03397_));
 sg13g2_nand2_1 _19129_ (.Y(_03409_),
    .A(\top_ihp.oisc.regs[53][18] ),
    .B(net616));
 sg13g2_o21ai_1 _19130_ (.B1(_03409_),
    .Y(_01997_),
    .A1(net89),
    .A2(net617));
 sg13g2_buf_1 _19131_ (.A(net699),
    .X(_03410_));
 sg13g2_nand2_1 _19132_ (.Y(_03411_),
    .A(\top_ihp.oisc.regs[53][19] ),
    .B(net616));
 sg13g2_o21ai_1 _19133_ (.B1(_03411_),
    .Y(_01998_),
    .A1(_03020_),
    .A2(net615));
 sg13g2_nand2_1 _19134_ (.Y(_03412_),
    .A(\top_ihp.oisc.regs[53][1] ),
    .B(net616));
 sg13g2_o21ai_1 _19135_ (.B1(_03412_),
    .Y(_01999_),
    .A1(_11170_),
    .A2(net615));
 sg13g2_nand2_1 _19136_ (.Y(_03413_),
    .A(\top_ihp.oisc.regs[53][20] ),
    .B(net616));
 sg13g2_o21ai_1 _19137_ (.B1(_03413_),
    .Y(_02000_),
    .A1(net636),
    .A2(net615));
 sg13g2_nand2_1 _19138_ (.Y(_03414_),
    .A(\top_ihp.oisc.regs[53][21] ),
    .B(_03407_));
 sg13g2_o21ai_1 _19139_ (.B1(_03414_),
    .Y(_02001_),
    .A1(_03025_),
    .A2(_03410_));
 sg13g2_nand2_1 _19140_ (.Y(_03415_),
    .A(\top_ihp.oisc.regs[53][22] ),
    .B(net616));
 sg13g2_o21ai_1 _19141_ (.B1(_03415_),
    .Y(_02002_),
    .A1(_11174_),
    .A2(net615));
 sg13g2_nand2_1 _19142_ (.Y(_03416_),
    .A(\top_ihp.oisc.regs[53][23] ),
    .B(_03407_));
 sg13g2_o21ai_1 _19143_ (.B1(_03416_),
    .Y(_02003_),
    .A1(_03028_),
    .A2(_03410_));
 sg13g2_nand2_1 _19144_ (.Y(_03417_),
    .A(\top_ihp.oisc.regs[53][24] ),
    .B(net616));
 sg13g2_o21ai_1 _19145_ (.B1(_03417_),
    .Y(_02004_),
    .A1(_03030_),
    .A2(net615));
 sg13g2_nand2_1 _19146_ (.Y(_03418_),
    .A(\top_ihp.oisc.regs[53][25] ),
    .B(net616));
 sg13g2_o21ai_1 _19147_ (.B1(_03418_),
    .Y(_02005_),
    .A1(_02892_),
    .A2(net615));
 sg13g2_buf_1 _19148_ (.A(_03396_),
    .X(_03419_));
 sg13g2_nand2_1 _19149_ (.Y(_03420_),
    .A(\top_ihp.oisc.regs[53][26] ),
    .B(_03419_));
 sg13g2_o21ai_1 _19150_ (.B1(_03420_),
    .Y(_02006_),
    .A1(_03034_),
    .A2(net615));
 sg13g2_nand2_1 _19151_ (.Y(_03421_),
    .A(\top_ihp.oisc.regs[53][27] ),
    .B(net614));
 sg13g2_o21ai_1 _19152_ (.B1(_03421_),
    .Y(_02007_),
    .A1(_03036_),
    .A2(net615));
 sg13g2_buf_1 _19153_ (.A(net699),
    .X(_03422_));
 sg13g2_nand2_1 _19154_ (.Y(_03423_),
    .A(\top_ihp.oisc.regs[53][28] ),
    .B(net614));
 sg13g2_o21ai_1 _19155_ (.B1(_03423_),
    .Y(_02008_),
    .A1(_03038_),
    .A2(net613));
 sg13g2_nand2_1 _19156_ (.Y(_03424_),
    .A(\top_ihp.oisc.regs[53][29] ),
    .B(net614));
 sg13g2_o21ai_1 _19157_ (.B1(_03424_),
    .Y(_02009_),
    .A1(_03040_),
    .A2(net613));
 sg13g2_nand2_1 _19158_ (.Y(_03425_),
    .A(\top_ihp.oisc.regs[53][2] ),
    .B(net614));
 sg13g2_o21ai_1 _19159_ (.B1(_03425_),
    .Y(_02010_),
    .A1(_03089_),
    .A2(net613));
 sg13g2_nand2_1 _19160_ (.Y(_03426_),
    .A(\top_ihp.oisc.regs[53][30] ),
    .B(_03419_));
 sg13g2_o21ai_1 _19161_ (.B1(_03426_),
    .Y(_02011_),
    .A1(_03091_),
    .A2(net613));
 sg13g2_nand2_1 _19162_ (.Y(_03427_),
    .A(\top_ihp.oisc.regs[53][31] ),
    .B(net614));
 sg13g2_o21ai_1 _19163_ (.B1(_03427_),
    .Y(_02012_),
    .A1(_02943_),
    .A2(net613));
 sg13g2_nand2_1 _19164_ (.Y(_03428_),
    .A(\top_ihp.oisc.regs[53][3] ),
    .B(net614));
 sg13g2_o21ai_1 _19165_ (.B1(_03428_),
    .Y(_02013_),
    .A1(_03094_),
    .A2(net613));
 sg13g2_nand2_1 _19166_ (.Y(_03429_),
    .A(\top_ihp.oisc.regs[53][4] ),
    .B(net614));
 sg13g2_o21ai_1 _19167_ (.B1(_03429_),
    .Y(_02014_),
    .A1(net29),
    .A2(_03422_));
 sg13g2_nand2_1 _19168_ (.Y(_03430_),
    .A(\top_ihp.oisc.regs[53][5] ),
    .B(net614));
 sg13g2_o21ai_1 _19169_ (.B1(_03430_),
    .Y(_02015_),
    .A1(_03047_),
    .A2(_03422_));
 sg13g2_nand2_1 _19170_ (.Y(_03431_),
    .A(\top_ihp.oisc.regs[53][6] ),
    .B(net699));
 sg13g2_o21ai_1 _19171_ (.B1(_03431_),
    .Y(_02016_),
    .A1(_03049_),
    .A2(net613));
 sg13g2_nand2_1 _19172_ (.Y(_03432_),
    .A(\top_ihp.oisc.regs[53][7] ),
    .B(net699));
 sg13g2_o21ai_1 _19173_ (.B1(_03432_),
    .Y(_02017_),
    .A1(net501),
    .A2(net613));
 sg13g2_nand2_1 _19174_ (.Y(_03433_),
    .A(\top_ihp.oisc.regs[53][8] ),
    .B(net699));
 sg13g2_o21ai_1 _19175_ (.B1(_03433_),
    .Y(_02018_),
    .A1(net83),
    .A2(net698));
 sg13g2_nand2_1 _19176_ (.Y(_03434_),
    .A(\top_ihp.oisc.regs[53][9] ),
    .B(net699));
 sg13g2_o21ai_1 _19177_ (.B1(_03434_),
    .Y(_02019_),
    .A1(_03054_),
    .A2(net698));
 sg13g2_nand3_1 _19178_ (.B(_10953_),
    .C(_03146_),
    .A(_10870_),
    .Y(_03435_));
 sg13g2_buf_1 _19179_ (.A(_03435_),
    .X(_03436_));
 sg13g2_buf_8 _19180_ (.A(_03436_),
    .X(_03437_));
 sg13g2_buf_1 _19181_ (.A(net612),
    .X(_03438_));
 sg13g2_buf_1 _19182_ (.A(_03436_),
    .X(_03439_));
 sg13g2_nand2_1 _19183_ (.Y(_03440_),
    .A(\top_ihp.oisc.regs[54][0] ),
    .B(net611));
 sg13g2_o21ai_1 _19184_ (.B1(_03440_),
    .Y(_02020_),
    .A1(net82),
    .A2(_03438_));
 sg13g2_buf_2 _19185_ (.A(_09824_),
    .X(_03441_));
 sg13g2_nand2_1 _19186_ (.Y(_03442_),
    .A(\top_ihp.oisc.regs[54][10] ),
    .B(net611));
 sg13g2_o21ai_1 _19187_ (.B1(_03442_),
    .Y(_02021_),
    .A1(net81),
    .A2(net475));
 sg13g2_nand2_1 _19188_ (.Y(_03443_),
    .A(\top_ihp.oisc.regs[54][11] ),
    .B(net611));
 sg13g2_o21ai_1 _19189_ (.B1(_03443_),
    .Y(_02022_),
    .A1(net33),
    .A2(net475));
 sg13g2_buf_8 _19190_ (.A(net332),
    .X(_03444_));
 sg13g2_nand2_1 _19191_ (.Y(_03445_),
    .A(\top_ihp.oisc.regs[54][12] ),
    .B(net611));
 sg13g2_o21ai_1 _19192_ (.B1(_03445_),
    .Y(_02023_),
    .A1(net80),
    .A2(net475));
 sg13g2_buf_8 _19193_ (.A(_10626_),
    .X(_03446_));
 sg13g2_nand2_1 _19194_ (.Y(_03447_),
    .A(\top_ihp.oisc.regs[54][13] ),
    .B(net611));
 sg13g2_o21ai_1 _19195_ (.B1(_03447_),
    .Y(_02024_),
    .A1(net79),
    .A2(net475));
 sg13g2_buf_1 _19196_ (.A(_09976_),
    .X(_03448_));
 sg13g2_nand2_1 _19197_ (.Y(_03449_),
    .A(\top_ihp.oisc.regs[54][14] ),
    .B(net611));
 sg13g2_o21ai_1 _19198_ (.B1(_03449_),
    .Y(_02025_),
    .A1(net230),
    .A2(net475));
 sg13g2_nand2_1 _19199_ (.Y(_03450_),
    .A(\top_ihp.oisc.regs[54][15] ),
    .B(net611));
 sg13g2_o21ai_1 _19200_ (.B1(_03450_),
    .Y(_02026_),
    .A1(_02879_),
    .A2(net475));
 sg13g2_buf_1 _19201_ (.A(_10014_),
    .X(_03451_));
 sg13g2_nand2_1 _19202_ (.Y(_03452_),
    .A(\top_ihp.oisc.regs[54][16] ),
    .B(net611));
 sg13g2_o21ai_1 _19203_ (.B1(_03452_),
    .Y(_02027_),
    .A1(net78),
    .A2(net475));
 sg13g2_buf_2 _19204_ (.A(_10038_),
    .X(_03453_));
 sg13g2_buf_1 _19205_ (.A(net612),
    .X(_03454_));
 sg13g2_nand2_1 _19206_ (.Y(_03455_),
    .A(\top_ihp.oisc.regs[54][17] ),
    .B(_03454_));
 sg13g2_o21ai_1 _19207_ (.B1(_03455_),
    .Y(_02028_),
    .A1(net229),
    .A2(net475));
 sg13g2_buf_2 _19208_ (.A(_10059_),
    .X(_03456_));
 sg13g2_nand2_1 _19209_ (.Y(_03457_),
    .A(\top_ihp.oisc.regs[54][18] ),
    .B(net474));
 sg13g2_o21ai_1 _19210_ (.B1(_03457_),
    .Y(_02029_),
    .A1(net228),
    .A2(_03438_));
 sg13g2_buf_8 _19211_ (.A(_10631_),
    .X(_03458_));
 sg13g2_buf_2 _19212_ (.A(net612),
    .X(_03459_));
 sg13g2_nand2_1 _19213_ (.Y(_03460_),
    .A(\top_ihp.oisc.regs[54][19] ),
    .B(net474));
 sg13g2_o21ai_1 _19214_ (.B1(_03460_),
    .Y(_02030_),
    .A1(net77),
    .A2(net473));
 sg13g2_buf_1 _19215_ (.A(net325),
    .X(_03461_));
 sg13g2_nand2_1 _19216_ (.Y(_03462_),
    .A(\top_ihp.oisc.regs[54][1] ),
    .B(net474));
 sg13g2_o21ai_1 _19217_ (.B1(_03462_),
    .Y(_02031_),
    .A1(net76),
    .A2(net473));
 sg13g2_nand2_1 _19218_ (.Y(_03463_),
    .A(\top_ihp.oisc.regs[54][20] ),
    .B(net474));
 sg13g2_o21ai_1 _19219_ (.B1(_03463_),
    .Y(_02032_),
    .A1(_10152_),
    .A2(net473));
 sg13g2_buf_2 _19220_ (.A(_10168_),
    .X(_03464_));
 sg13g2_nand2_1 _19221_ (.Y(_03465_),
    .A(\top_ihp.oisc.regs[54][21] ),
    .B(net474));
 sg13g2_o21ai_1 _19222_ (.B1(_03465_),
    .Y(_02033_),
    .A1(net227),
    .A2(net473));
 sg13g2_buf_8 _19223_ (.A(net322),
    .X(_03466_));
 sg13g2_nand2_1 _19224_ (.Y(_03467_),
    .A(\top_ihp.oisc.regs[54][22] ),
    .B(net474));
 sg13g2_o21ai_1 _19225_ (.B1(_03467_),
    .Y(_02034_),
    .A1(net75),
    .A2(net473));
 sg13g2_buf_8 _19226_ (.A(net528),
    .X(_03468_));
 sg13g2_nand2_1 _19227_ (.Y(_03469_),
    .A(\top_ihp.oisc.regs[54][23] ),
    .B(net474));
 sg13g2_o21ai_1 _19228_ (.B1(_03469_),
    .Y(_02035_),
    .A1(net226),
    .A2(_03459_));
 sg13g2_buf_2 _19229_ (.A(_10216_),
    .X(_03470_));
 sg13g2_nand2_1 _19230_ (.Y(_03471_),
    .A(\top_ihp.oisc.regs[54][24] ),
    .B(_03454_));
 sg13g2_o21ai_1 _19231_ (.B1(_03471_),
    .Y(_02036_),
    .A1(net225),
    .A2(net473));
 sg13g2_buf_1 _19232_ (.A(net319),
    .X(_03472_));
 sg13g2_nand2_1 _19233_ (.Y(_03473_),
    .A(\top_ihp.oisc.regs[54][25] ),
    .B(net474));
 sg13g2_o21ai_1 _19234_ (.B1(_03473_),
    .Y(_02037_),
    .A1(net74),
    .A2(net473));
 sg13g2_buf_1 _19235_ (.A(_10638_),
    .X(_03474_));
 sg13g2_buf_1 _19236_ (.A(net612),
    .X(_03475_));
 sg13g2_nand2_1 _19237_ (.Y(_03476_),
    .A(\top_ihp.oisc.regs[54][26] ),
    .B(net472));
 sg13g2_o21ai_1 _19238_ (.B1(_03476_),
    .Y(_02038_),
    .A1(net28),
    .A2(net473));
 sg13g2_buf_2 _19239_ (.A(_10259_),
    .X(_03477_));
 sg13g2_nand2_1 _19240_ (.Y(_03478_),
    .A(\top_ihp.oisc.regs[54][27] ),
    .B(net472));
 sg13g2_o21ai_1 _19241_ (.B1(_03478_),
    .Y(_02039_),
    .A1(net224),
    .A2(_03459_));
 sg13g2_buf_8 _19242_ (.A(_10640_),
    .X(_03479_));
 sg13g2_buf_1 _19243_ (.A(net612),
    .X(_03480_));
 sg13g2_nand2_1 _19244_ (.Y(_03481_),
    .A(\top_ihp.oisc.regs[54][28] ),
    .B(net472));
 sg13g2_o21ai_1 _19245_ (.B1(_03481_),
    .Y(_02040_),
    .A1(_03479_),
    .A2(net471));
 sg13g2_buf_1 _19246_ (.A(_10280_),
    .X(_03482_));
 sg13g2_nand2_1 _19247_ (.Y(_03483_),
    .A(\top_ihp.oisc.regs[54][29] ),
    .B(net472));
 sg13g2_o21ai_1 _19248_ (.B1(_03483_),
    .Y(_02041_),
    .A1(net222),
    .A2(net471));
 sg13g2_nand2_1 _19249_ (.Y(_03484_),
    .A(\top_ihp.oisc.regs[54][2] ),
    .B(net472));
 sg13g2_o21ai_1 _19250_ (.B1(_03484_),
    .Y(_02042_),
    .A1(_03089_),
    .A2(net471));
 sg13g2_nand2_1 _19251_ (.Y(_03485_),
    .A(\top_ihp.oisc.regs[54][30] ),
    .B(net472));
 sg13g2_o21ai_1 _19252_ (.B1(_03485_),
    .Y(_02043_),
    .A1(net31),
    .A2(net471));
 sg13g2_nand2_1 _19253_ (.Y(_03486_),
    .A(\top_ihp.oisc.regs[54][31] ),
    .B(_03475_));
 sg13g2_o21ai_1 _19254_ (.B1(_03486_),
    .Y(_02044_),
    .A1(_10349_),
    .A2(_03480_));
 sg13g2_nand2_1 _19255_ (.Y(_03487_),
    .A(\top_ihp.oisc.regs[54][3] ),
    .B(net472));
 sg13g2_o21ai_1 _19256_ (.B1(_03487_),
    .Y(_02045_),
    .A1(_03094_),
    .A2(_03480_));
 sg13g2_nand2_1 _19257_ (.Y(_03488_),
    .A(\top_ihp.oisc.regs[54][4] ),
    .B(net472));
 sg13g2_o21ai_1 _19258_ (.B1(_03488_),
    .Y(_02046_),
    .A1(net29),
    .A2(net471));
 sg13g2_buf_2 _19259_ (.A(_10439_),
    .X(_03489_));
 sg13g2_nand2_1 _19260_ (.Y(_03490_),
    .A(\top_ihp.oisc.regs[54][5] ),
    .B(_03475_));
 sg13g2_o21ai_1 _19261_ (.B1(_03490_),
    .Y(_02047_),
    .A1(net73),
    .A2(net471));
 sg13g2_buf_1 _19262_ (.A(_10468_),
    .X(_03491_));
 sg13g2_nand2_1 _19263_ (.Y(_03492_),
    .A(\top_ihp.oisc.regs[54][6] ),
    .B(net612));
 sg13g2_o21ai_1 _19264_ (.B1(_03492_),
    .Y(_02048_),
    .A1(net72),
    .A2(net471));
 sg13g2_nand2_1 _19265_ (.Y(_03493_),
    .A(\top_ihp.oisc.regs[54][7] ),
    .B(_03437_));
 sg13g2_o21ai_1 _19266_ (.B1(_03493_),
    .Y(_02049_),
    .A1(_10483_),
    .A2(net471));
 sg13g2_buf_8 _19267_ (.A(_10498_),
    .X(_03494_));
 sg13g2_nand2_1 _19268_ (.Y(_03495_),
    .A(\top_ihp.oisc.regs[54][8] ),
    .B(net612));
 sg13g2_o21ai_1 _19269_ (.B1(_03495_),
    .Y(_02050_),
    .A1(_03494_),
    .A2(_03439_));
 sg13g2_buf_1 _19270_ (.A(_10513_),
    .X(_03496_));
 sg13g2_nand2_1 _19271_ (.Y(_03497_),
    .A(\top_ihp.oisc.regs[54][9] ),
    .B(net612));
 sg13g2_o21ai_1 _19272_ (.B1(_03497_),
    .Y(_02051_),
    .A1(net71),
    .A2(_03439_));
 sg13g2_buf_2 _19273_ (.A(_09696_),
    .X(_03498_));
 sg13g2_nand2_1 _19274_ (.Y(_03499_),
    .A(_10988_),
    .B(_03313_));
 sg13g2_buf_1 _19275_ (.A(_03499_),
    .X(_03500_));
 sg13g2_buf_1 _19276_ (.A(net697),
    .X(_03501_));
 sg13g2_buf_1 _19277_ (.A(_03499_),
    .X(_03502_));
 sg13g2_nand2_1 _19278_ (.Y(_03503_),
    .A(\top_ihp.oisc.regs[55][0] ),
    .B(net696));
 sg13g2_o21ai_1 _19279_ (.B1(_03503_),
    .Y(_02052_),
    .A1(net70),
    .A2(net610));
 sg13g2_nand2_1 _19280_ (.Y(_03504_),
    .A(\top_ihp.oisc.regs[55][10] ),
    .B(net696));
 sg13g2_o21ai_1 _19281_ (.B1(_03504_),
    .Y(_02053_),
    .A1(net81),
    .A2(net610));
 sg13g2_buf_2 _19282_ (.A(_09860_),
    .X(_03505_));
 sg13g2_nand2_1 _19283_ (.Y(_03506_),
    .A(\top_ihp.oisc.regs[55][11] ),
    .B(net696));
 sg13g2_o21ai_1 _19284_ (.B1(_03506_),
    .Y(_02054_),
    .A1(_03505_),
    .A2(net610));
 sg13g2_nand2_1 _19285_ (.Y(_03507_),
    .A(\top_ihp.oisc.regs[55][12] ),
    .B(net696));
 sg13g2_o21ai_1 _19286_ (.B1(_03507_),
    .Y(_02055_),
    .A1(net80),
    .A2(net610));
 sg13g2_nand2_1 _19287_ (.Y(_03508_),
    .A(\top_ihp.oisc.regs[55][13] ),
    .B(net696));
 sg13g2_o21ai_1 _19288_ (.B1(_03508_),
    .Y(_02056_),
    .A1(net79),
    .A2(net610));
 sg13g2_nand2_1 _19289_ (.Y(_03509_),
    .A(\top_ihp.oisc.regs[55][14] ),
    .B(net696));
 sg13g2_o21ai_1 _19290_ (.B1(_03509_),
    .Y(_02057_),
    .A1(_03448_),
    .A2(net610));
 sg13g2_buf_2 _19291_ (.A(_09991_),
    .X(_03510_));
 sg13g2_nand2_1 _19292_ (.Y(_03511_),
    .A(\top_ihp.oisc.regs[55][15] ),
    .B(net696));
 sg13g2_o21ai_1 _19293_ (.B1(_03511_),
    .Y(_02058_),
    .A1(net220),
    .A2(net610));
 sg13g2_nand2_1 _19294_ (.Y(_03512_),
    .A(\top_ihp.oisc.regs[55][16] ),
    .B(net696));
 sg13g2_o21ai_1 _19295_ (.B1(_03512_),
    .Y(_02059_),
    .A1(net78),
    .A2(net610));
 sg13g2_buf_1 _19296_ (.A(net697),
    .X(_03513_));
 sg13g2_nand2_1 _19297_ (.Y(_03514_),
    .A(\top_ihp.oisc.regs[55][17] ),
    .B(_03513_));
 sg13g2_o21ai_1 _19298_ (.B1(_03514_),
    .Y(_02060_),
    .A1(net229),
    .A2(_03501_));
 sg13g2_nand2_1 _19299_ (.Y(_03515_),
    .A(\top_ihp.oisc.regs[55][18] ),
    .B(net609));
 sg13g2_o21ai_1 _19300_ (.B1(_03515_),
    .Y(_02061_),
    .A1(net228),
    .A2(_03501_));
 sg13g2_buf_1 _19301_ (.A(net697),
    .X(_03516_));
 sg13g2_nand2_1 _19302_ (.Y(_03517_),
    .A(\top_ihp.oisc.regs[55][19] ),
    .B(_03513_));
 sg13g2_o21ai_1 _19303_ (.B1(_03517_),
    .Y(_02062_),
    .A1(net77),
    .A2(net608));
 sg13g2_nand2_1 _19304_ (.Y(_03518_),
    .A(\top_ihp.oisc.regs[55][1] ),
    .B(net609));
 sg13g2_o21ai_1 _19305_ (.B1(_03518_),
    .Y(_02063_),
    .A1(net76),
    .A2(net608));
 sg13g2_buf_1 _19306_ (.A(_10144_),
    .X(_03519_));
 sg13g2_nand2_1 _19307_ (.Y(_03520_),
    .A(\top_ihp.oisc.regs[55][20] ),
    .B(net609));
 sg13g2_o21ai_1 _19308_ (.B1(_03520_),
    .Y(_02064_),
    .A1(net607),
    .A2(net608));
 sg13g2_nand2_1 _19309_ (.Y(_03521_),
    .A(\top_ihp.oisc.regs[55][21] ),
    .B(net609));
 sg13g2_o21ai_1 _19310_ (.B1(_03521_),
    .Y(_02065_),
    .A1(net227),
    .A2(net608));
 sg13g2_nand2_1 _19311_ (.Y(_03522_),
    .A(\top_ihp.oisc.regs[55][22] ),
    .B(net609));
 sg13g2_o21ai_1 _19312_ (.B1(_03522_),
    .Y(_02066_),
    .A1(net75),
    .A2(net608));
 sg13g2_nand2_1 _19313_ (.Y(_03523_),
    .A(\top_ihp.oisc.regs[55][23] ),
    .B(net609));
 sg13g2_o21ai_1 _19314_ (.B1(_03523_),
    .Y(_02067_),
    .A1(net226),
    .A2(_03516_));
 sg13g2_nand2_1 _19315_ (.Y(_03524_),
    .A(\top_ihp.oisc.regs[55][24] ),
    .B(net609));
 sg13g2_o21ai_1 _19316_ (.B1(_03524_),
    .Y(_02068_),
    .A1(net225),
    .A2(_03516_));
 sg13g2_nand2_1 _19317_ (.Y(_03525_),
    .A(\top_ihp.oisc.regs[55][25] ),
    .B(net609));
 sg13g2_o21ai_1 _19318_ (.B1(_03525_),
    .Y(_02069_),
    .A1(net74),
    .A2(net608));
 sg13g2_buf_1 _19319_ (.A(net697),
    .X(_03526_));
 sg13g2_nand2_1 _19320_ (.Y(_03527_),
    .A(\top_ihp.oisc.regs[55][26] ),
    .B(net606));
 sg13g2_o21ai_1 _19321_ (.B1(_03527_),
    .Y(_02070_),
    .A1(net28),
    .A2(net608));
 sg13g2_nand2_1 _19322_ (.Y(_03528_),
    .A(\top_ihp.oisc.regs[55][27] ),
    .B(_03526_));
 sg13g2_o21ai_1 _19323_ (.B1(_03528_),
    .Y(_02071_),
    .A1(net224),
    .A2(net608));
 sg13g2_buf_1 _19324_ (.A(net697),
    .X(_03529_));
 sg13g2_nand2_1 _19325_ (.Y(_03530_),
    .A(\top_ihp.oisc.regs[55][28] ),
    .B(net606));
 sg13g2_o21ai_1 _19326_ (.B1(_03530_),
    .Y(_02072_),
    .A1(net223),
    .A2(net605));
 sg13g2_nand2_1 _19327_ (.Y(_03531_),
    .A(\top_ihp.oisc.regs[55][29] ),
    .B(net606));
 sg13g2_o21ai_1 _19328_ (.B1(_03531_),
    .Y(_02073_),
    .A1(_03482_),
    .A2(net605));
 sg13g2_buf_2 _19329_ (.A(_10314_),
    .X(_03532_));
 sg13g2_nand2_1 _19330_ (.Y(_03533_),
    .A(\top_ihp.oisc.regs[55][2] ),
    .B(net606));
 sg13g2_o21ai_1 _19331_ (.B1(_03533_),
    .Y(_02074_),
    .A1(net68),
    .A2(net605));
 sg13g2_buf_1 _19332_ (.A(_10326_),
    .X(_03534_));
 sg13g2_nand2_1 _19333_ (.Y(_03535_),
    .A(\top_ihp.oisc.regs[55][30] ),
    .B(net606));
 sg13g2_o21ai_1 _19334_ (.B1(_03535_),
    .Y(_02075_),
    .A1(net67),
    .A2(_03529_));
 sg13g2_nand2_1 _19335_ (.Y(_03536_),
    .A(\top_ihp.oisc.regs[55][31] ),
    .B(_03526_));
 sg13g2_o21ai_1 _19336_ (.B1(_03536_),
    .Y(_02076_),
    .A1(_02943_),
    .A2(_03529_));
 sg13g2_buf_2 _19337_ (.A(_10380_),
    .X(_03537_));
 sg13g2_nand2_1 _19338_ (.Y(_03538_),
    .A(\top_ihp.oisc.regs[55][3] ),
    .B(net606));
 sg13g2_o21ai_1 _19339_ (.B1(_03538_),
    .Y(_02077_),
    .A1(net66),
    .A2(net605));
 sg13g2_buf_2 _19340_ (.A(_10412_),
    .X(_03539_));
 sg13g2_nand2_1 _19341_ (.Y(_03540_),
    .A(\top_ihp.oisc.regs[55][4] ),
    .B(net606));
 sg13g2_o21ai_1 _19342_ (.B1(_03540_),
    .Y(_02078_),
    .A1(net65),
    .A2(net605));
 sg13g2_nand2_1 _19343_ (.Y(_03541_),
    .A(\top_ihp.oisc.regs[55][5] ),
    .B(net606));
 sg13g2_o21ai_1 _19344_ (.B1(_03541_),
    .Y(_02079_),
    .A1(net73),
    .A2(net605));
 sg13g2_nand2_1 _19345_ (.Y(_03542_),
    .A(\top_ihp.oisc.regs[55][6] ),
    .B(net697));
 sg13g2_o21ai_1 _19346_ (.B1(_03542_),
    .Y(_02080_),
    .A1(net72),
    .A2(net605));
 sg13g2_buf_2 _19347_ (.A(_10480_),
    .X(_03543_));
 sg13g2_nand2_1 _19348_ (.Y(_03544_),
    .A(\top_ihp.oisc.regs[55][7] ),
    .B(net697));
 sg13g2_o21ai_1 _19349_ (.B1(_03544_),
    .Y(_02081_),
    .A1(net470),
    .A2(net605));
 sg13g2_nand2_1 _19350_ (.Y(_03545_),
    .A(\top_ihp.oisc.regs[55][8] ),
    .B(_03500_));
 sg13g2_o21ai_1 _19351_ (.B1(_03545_),
    .Y(_02082_),
    .A1(net221),
    .A2(_03502_));
 sg13g2_nand2_1 _19352_ (.Y(_03546_),
    .A(\top_ihp.oisc.regs[55][9] ),
    .B(net697));
 sg13g2_o21ai_1 _19353_ (.B1(_03546_),
    .Y(_02083_),
    .A1(net71),
    .A2(_03502_));
 sg13g2_nand2_1 _19354_ (.Y(_03547_),
    .A(_10520_),
    .B(_03148_));
 sg13g2_buf_1 _19355_ (.A(_03547_),
    .X(_03548_));
 sg13g2_buf_1 _19356_ (.A(net604),
    .X(_03549_));
 sg13g2_buf_1 _19357_ (.A(_03547_),
    .X(_03550_));
 sg13g2_nand2_1 _19358_ (.Y(_03551_),
    .A(\top_ihp.oisc.regs[56][0] ),
    .B(net603));
 sg13g2_o21ai_1 _19359_ (.B1(_03551_),
    .Y(_02084_),
    .A1(net70),
    .A2(net469));
 sg13g2_nand2_1 _19360_ (.Y(_03552_),
    .A(\top_ihp.oisc.regs[56][10] ),
    .B(net603));
 sg13g2_o21ai_1 _19361_ (.B1(_03552_),
    .Y(_02085_),
    .A1(net81),
    .A2(net469));
 sg13g2_nand2_1 _19362_ (.Y(_03553_),
    .A(\top_ihp.oisc.regs[56][11] ),
    .B(net603));
 sg13g2_o21ai_1 _19363_ (.B1(_03553_),
    .Y(_02086_),
    .A1(net69),
    .A2(net469));
 sg13g2_nand2_1 _19364_ (.Y(_03554_),
    .A(\top_ihp.oisc.regs[56][12] ),
    .B(net603));
 sg13g2_o21ai_1 _19365_ (.B1(_03554_),
    .Y(_02087_),
    .A1(net80),
    .A2(net469));
 sg13g2_nand2_1 _19366_ (.Y(_03555_),
    .A(\top_ihp.oisc.regs[56][13] ),
    .B(_03550_));
 sg13g2_o21ai_1 _19367_ (.B1(_03555_),
    .Y(_02088_),
    .A1(net79),
    .A2(_03549_));
 sg13g2_nand2_1 _19368_ (.Y(_03556_),
    .A(\top_ihp.oisc.regs[56][14] ),
    .B(net603));
 sg13g2_o21ai_1 _19369_ (.B1(_03556_),
    .Y(_02089_),
    .A1(net230),
    .A2(net469));
 sg13g2_nand2_1 _19370_ (.Y(_03557_),
    .A(\top_ihp.oisc.regs[56][15] ),
    .B(net603));
 sg13g2_o21ai_1 _19371_ (.B1(_03557_),
    .Y(_02090_),
    .A1(net220),
    .A2(net469));
 sg13g2_nand2_1 _19372_ (.Y(_03558_),
    .A(\top_ihp.oisc.regs[56][16] ),
    .B(_03550_));
 sg13g2_o21ai_1 _19373_ (.B1(_03558_),
    .Y(_02091_),
    .A1(net78),
    .A2(net469));
 sg13g2_buf_1 _19374_ (.A(net604),
    .X(_03559_));
 sg13g2_nand2_1 _19375_ (.Y(_03560_),
    .A(\top_ihp.oisc.regs[56][17] ),
    .B(_03559_));
 sg13g2_o21ai_1 _19376_ (.B1(_03560_),
    .Y(_02092_),
    .A1(net229),
    .A2(net469));
 sg13g2_nand2_1 _19377_ (.Y(_03561_),
    .A(\top_ihp.oisc.regs[56][18] ),
    .B(_03559_));
 sg13g2_o21ai_1 _19378_ (.B1(_03561_),
    .Y(_02093_),
    .A1(net228),
    .A2(_03549_));
 sg13g2_buf_1 _19379_ (.A(net604),
    .X(_03562_));
 sg13g2_nand2_1 _19380_ (.Y(_03563_),
    .A(\top_ihp.oisc.regs[56][19] ),
    .B(net468));
 sg13g2_o21ai_1 _19381_ (.B1(_03563_),
    .Y(_02094_),
    .A1(_03458_),
    .A2(net467));
 sg13g2_nand2_1 _19382_ (.Y(_03564_),
    .A(\top_ihp.oisc.regs[56][1] ),
    .B(net468));
 sg13g2_o21ai_1 _19383_ (.B1(_03564_),
    .Y(_02095_),
    .A1(net76),
    .A2(net467));
 sg13g2_nand2_1 _19384_ (.Y(_03565_),
    .A(\top_ihp.oisc.regs[56][20] ),
    .B(net468));
 sg13g2_o21ai_1 _19385_ (.B1(_03565_),
    .Y(_02096_),
    .A1(net607),
    .A2(net467));
 sg13g2_nand2_1 _19386_ (.Y(_03566_),
    .A(\top_ihp.oisc.regs[56][21] ),
    .B(net468));
 sg13g2_o21ai_1 _19387_ (.B1(_03566_),
    .Y(_02097_),
    .A1(net227),
    .A2(net467));
 sg13g2_nand2_1 _19388_ (.Y(_03567_),
    .A(\top_ihp.oisc.regs[56][22] ),
    .B(net468));
 sg13g2_o21ai_1 _19389_ (.B1(_03567_),
    .Y(_02098_),
    .A1(net75),
    .A2(net467));
 sg13g2_nand2_1 _19390_ (.Y(_03568_),
    .A(\top_ihp.oisc.regs[56][23] ),
    .B(net468));
 sg13g2_o21ai_1 _19391_ (.B1(_03568_),
    .Y(_02099_),
    .A1(net226),
    .A2(net467));
 sg13g2_nand2_1 _19392_ (.Y(_03569_),
    .A(\top_ihp.oisc.regs[56][24] ),
    .B(net468));
 sg13g2_o21ai_1 _19393_ (.B1(_03569_),
    .Y(_02100_),
    .A1(net225),
    .A2(_03562_));
 sg13g2_nand2_1 _19394_ (.Y(_03570_),
    .A(\top_ihp.oisc.regs[56][25] ),
    .B(net468));
 sg13g2_o21ai_1 _19395_ (.B1(_03570_),
    .Y(_02101_),
    .A1(net74),
    .A2(net467));
 sg13g2_buf_2 _19396_ (.A(net604),
    .X(_03571_));
 sg13g2_nand2_1 _19397_ (.Y(_03572_),
    .A(\top_ihp.oisc.regs[56][26] ),
    .B(net466));
 sg13g2_o21ai_1 _19398_ (.B1(_03572_),
    .Y(_02102_),
    .A1(net28),
    .A2(net467));
 sg13g2_nand2_1 _19399_ (.Y(_03573_),
    .A(\top_ihp.oisc.regs[56][27] ),
    .B(net466));
 sg13g2_o21ai_1 _19400_ (.B1(_03573_),
    .Y(_02103_),
    .A1(net224),
    .A2(_03562_));
 sg13g2_buf_1 _19401_ (.A(net604),
    .X(_03574_));
 sg13g2_nand2_1 _19402_ (.Y(_03575_),
    .A(\top_ihp.oisc.regs[56][28] ),
    .B(net466));
 sg13g2_o21ai_1 _19403_ (.B1(_03575_),
    .Y(_02104_),
    .A1(net223),
    .A2(net465));
 sg13g2_nand2_1 _19404_ (.Y(_03576_),
    .A(\top_ihp.oisc.regs[56][29] ),
    .B(net466));
 sg13g2_o21ai_1 _19405_ (.B1(_03576_),
    .Y(_02105_),
    .A1(net222),
    .A2(net465));
 sg13g2_nand2_1 _19406_ (.Y(_03577_),
    .A(\top_ihp.oisc.regs[56][2] ),
    .B(net466));
 sg13g2_o21ai_1 _19407_ (.B1(_03577_),
    .Y(_02106_),
    .A1(net68),
    .A2(net465));
 sg13g2_nand2_1 _19408_ (.Y(_03578_),
    .A(\top_ihp.oisc.regs[56][30] ),
    .B(net466));
 sg13g2_o21ai_1 _19409_ (.B1(_03578_),
    .Y(_02107_),
    .A1(_03534_),
    .A2(net465));
 sg13g2_nand2_1 _19410_ (.Y(_03579_),
    .A(\top_ihp.oisc.regs[56][31] ),
    .B(net466));
 sg13g2_o21ai_1 _19411_ (.B1(_03579_),
    .Y(_02108_),
    .A1(net306),
    .A2(net465));
 sg13g2_nand2_1 _19412_ (.Y(_03580_),
    .A(\top_ihp.oisc.regs[56][3] ),
    .B(net466));
 sg13g2_o21ai_1 _19413_ (.B1(_03580_),
    .Y(_02109_),
    .A1(net66),
    .A2(net465));
 sg13g2_nand2_1 _19414_ (.Y(_03581_),
    .A(\top_ihp.oisc.regs[56][4] ),
    .B(_03571_));
 sg13g2_o21ai_1 _19415_ (.B1(_03581_),
    .Y(_02110_),
    .A1(net65),
    .A2(_03574_));
 sg13g2_nand2_1 _19416_ (.Y(_03582_),
    .A(\top_ihp.oisc.regs[56][5] ),
    .B(_03571_));
 sg13g2_o21ai_1 _19417_ (.B1(_03582_),
    .Y(_02111_),
    .A1(net73),
    .A2(_03574_));
 sg13g2_nand2_1 _19418_ (.Y(_03583_),
    .A(\top_ihp.oisc.regs[56][6] ),
    .B(_03548_));
 sg13g2_o21ai_1 _19419_ (.B1(_03583_),
    .Y(_02112_),
    .A1(net72),
    .A2(net465));
 sg13g2_nand2_1 _19420_ (.Y(_03584_),
    .A(\top_ihp.oisc.regs[56][7] ),
    .B(net604));
 sg13g2_o21ai_1 _19421_ (.B1(_03584_),
    .Y(_02113_),
    .A1(net470),
    .A2(net465));
 sg13g2_nand2_1 _19422_ (.Y(_03585_),
    .A(\top_ihp.oisc.regs[56][8] ),
    .B(net604));
 sg13g2_o21ai_1 _19423_ (.B1(_03585_),
    .Y(_02114_),
    .A1(net221),
    .A2(net603));
 sg13g2_nand2_1 _19424_ (.Y(_03586_),
    .A(\top_ihp.oisc.regs[56][9] ),
    .B(net604));
 sg13g2_o21ai_1 _19425_ (.B1(_03586_),
    .Y(_02115_),
    .A1(net71),
    .A2(net603));
 sg13g2_or2_1 _19426_ (.X(_03587_),
    .B(_03189_),
    .A(_11203_));
 sg13g2_buf_1 _19427_ (.A(_03587_),
    .X(_03588_));
 sg13g2_buf_1 _19428_ (.A(_03588_),
    .X(_03589_));
 sg13g2_buf_1 _19429_ (.A(net695),
    .X(_03590_));
 sg13g2_buf_1 _19430_ (.A(_03588_),
    .X(_03591_));
 sg13g2_nand2_1 _19431_ (.Y(_03592_),
    .A(\top_ihp.oisc.regs[57][0] ),
    .B(_03591_));
 sg13g2_o21ai_1 _19432_ (.B1(_03592_),
    .Y(_02116_),
    .A1(net70),
    .A2(_03590_));
 sg13g2_nand2_1 _19433_ (.Y(_03593_),
    .A(\top_ihp.oisc.regs[57][10] ),
    .B(net694));
 sg13g2_o21ai_1 _19434_ (.B1(_03593_),
    .Y(_02117_),
    .A1(net81),
    .A2(net602));
 sg13g2_nand2_1 _19435_ (.Y(_03594_),
    .A(\top_ihp.oisc.regs[57][11] ),
    .B(net694));
 sg13g2_o21ai_1 _19436_ (.B1(_03594_),
    .Y(_02118_),
    .A1(net69),
    .A2(net602));
 sg13g2_nand2_1 _19437_ (.Y(_03595_),
    .A(\top_ihp.oisc.regs[57][12] ),
    .B(net694));
 sg13g2_o21ai_1 _19438_ (.B1(_03595_),
    .Y(_02119_),
    .A1(net80),
    .A2(net602));
 sg13g2_nand2_1 _19439_ (.Y(_03596_),
    .A(\top_ihp.oisc.regs[57][13] ),
    .B(net694));
 sg13g2_o21ai_1 _19440_ (.B1(_03596_),
    .Y(_02120_),
    .A1(net79),
    .A2(net602));
 sg13g2_nand2_1 _19441_ (.Y(_03597_),
    .A(\top_ihp.oisc.regs[57][14] ),
    .B(net694));
 sg13g2_o21ai_1 _19442_ (.B1(_03597_),
    .Y(_02121_),
    .A1(net230),
    .A2(net602));
 sg13g2_nand2_1 _19443_ (.Y(_03598_),
    .A(\top_ihp.oisc.regs[57][15] ),
    .B(net694));
 sg13g2_o21ai_1 _19444_ (.B1(_03598_),
    .Y(_02122_),
    .A1(net220),
    .A2(net602));
 sg13g2_nand2_1 _19445_ (.Y(_03599_),
    .A(\top_ihp.oisc.regs[57][16] ),
    .B(_03591_));
 sg13g2_o21ai_1 _19446_ (.B1(_03599_),
    .Y(_02123_),
    .A1(net78),
    .A2(net602));
 sg13g2_buf_1 _19447_ (.A(net695),
    .X(_03600_));
 sg13g2_nand2_1 _19448_ (.Y(_03601_),
    .A(\top_ihp.oisc.regs[57][17] ),
    .B(net601));
 sg13g2_o21ai_1 _19449_ (.B1(_03601_),
    .Y(_02124_),
    .A1(net229),
    .A2(net602));
 sg13g2_nand2_1 _19450_ (.Y(_03602_),
    .A(\top_ihp.oisc.regs[57][18] ),
    .B(net601));
 sg13g2_o21ai_1 _19451_ (.B1(_03602_),
    .Y(_02125_),
    .A1(net228),
    .A2(_03590_));
 sg13g2_buf_1 _19452_ (.A(net695),
    .X(_03603_));
 sg13g2_nand2_1 _19453_ (.Y(_03604_),
    .A(\top_ihp.oisc.regs[57][19] ),
    .B(net601));
 sg13g2_o21ai_1 _19454_ (.B1(_03604_),
    .Y(_02126_),
    .A1(net77),
    .A2(net600));
 sg13g2_nand2_1 _19455_ (.Y(_03605_),
    .A(\top_ihp.oisc.regs[57][1] ),
    .B(net601));
 sg13g2_o21ai_1 _19456_ (.B1(_03605_),
    .Y(_02127_),
    .A1(net76),
    .A2(net600));
 sg13g2_nand2_1 _19457_ (.Y(_03606_),
    .A(\top_ihp.oisc.regs[57][20] ),
    .B(net601));
 sg13g2_o21ai_1 _19458_ (.B1(_03606_),
    .Y(_02128_),
    .A1(net607),
    .A2(net600));
 sg13g2_nand2_1 _19459_ (.Y(_03607_),
    .A(\top_ihp.oisc.regs[57][21] ),
    .B(_03600_));
 sg13g2_o21ai_1 _19460_ (.B1(_03607_),
    .Y(_02129_),
    .A1(net227),
    .A2(net600));
 sg13g2_nand2_1 _19461_ (.Y(_03608_),
    .A(\top_ihp.oisc.regs[57][22] ),
    .B(net601));
 sg13g2_o21ai_1 _19462_ (.B1(_03608_),
    .Y(_02130_),
    .A1(net75),
    .A2(net600));
 sg13g2_nand2_1 _19463_ (.Y(_03609_),
    .A(\top_ihp.oisc.regs[57][23] ),
    .B(_03600_));
 sg13g2_o21ai_1 _19464_ (.B1(_03609_),
    .Y(_02131_),
    .A1(net226),
    .A2(_03603_));
 sg13g2_nand2_1 _19465_ (.Y(_03610_),
    .A(\top_ihp.oisc.regs[57][24] ),
    .B(net601));
 sg13g2_o21ai_1 _19466_ (.B1(_03610_),
    .Y(_02132_),
    .A1(net225),
    .A2(net600));
 sg13g2_nand2_1 _19467_ (.Y(_03611_),
    .A(\top_ihp.oisc.regs[57][25] ),
    .B(net601));
 sg13g2_o21ai_1 _19468_ (.B1(_03611_),
    .Y(_02133_),
    .A1(net74),
    .A2(net600));
 sg13g2_buf_1 _19469_ (.A(net695),
    .X(_03612_));
 sg13g2_nand2_1 _19470_ (.Y(_03613_),
    .A(\top_ihp.oisc.regs[57][26] ),
    .B(_03612_));
 sg13g2_o21ai_1 _19471_ (.B1(_03613_),
    .Y(_02134_),
    .A1(net28),
    .A2(net600));
 sg13g2_nand2_1 _19472_ (.Y(_03614_),
    .A(\top_ihp.oisc.regs[57][27] ),
    .B(net599));
 sg13g2_o21ai_1 _19473_ (.B1(_03614_),
    .Y(_02135_),
    .A1(net224),
    .A2(_03603_));
 sg13g2_buf_1 _19474_ (.A(net695),
    .X(_03615_));
 sg13g2_nand2_1 _19475_ (.Y(_03616_),
    .A(\top_ihp.oisc.regs[57][28] ),
    .B(net599));
 sg13g2_o21ai_1 _19476_ (.B1(_03616_),
    .Y(_02136_),
    .A1(net223),
    .A2(net598));
 sg13g2_nand2_1 _19477_ (.Y(_03617_),
    .A(\top_ihp.oisc.regs[57][29] ),
    .B(net599));
 sg13g2_o21ai_1 _19478_ (.B1(_03617_),
    .Y(_02137_),
    .A1(net222),
    .A2(net598));
 sg13g2_nand2_1 _19479_ (.Y(_03618_),
    .A(\top_ihp.oisc.regs[57][2] ),
    .B(net599));
 sg13g2_o21ai_1 _19480_ (.B1(_03618_),
    .Y(_02138_),
    .A1(net68),
    .A2(_03615_));
 sg13g2_nand2_1 _19481_ (.Y(_03619_),
    .A(\top_ihp.oisc.regs[57][30] ),
    .B(net599));
 sg13g2_o21ai_1 _19482_ (.B1(_03619_),
    .Y(_02139_),
    .A1(net67),
    .A2(net598));
 sg13g2_nand2_1 _19483_ (.Y(_03620_),
    .A(\top_ihp.oisc.regs[57][31] ),
    .B(net599));
 sg13g2_o21ai_1 _19484_ (.B1(_03620_),
    .Y(_02140_),
    .A1(net306),
    .A2(net598));
 sg13g2_nand2_1 _19485_ (.Y(_03621_),
    .A(\top_ihp.oisc.regs[57][3] ),
    .B(net599));
 sg13g2_o21ai_1 _19486_ (.B1(_03621_),
    .Y(_02141_),
    .A1(net66),
    .A2(net598));
 sg13g2_nand2_1 _19487_ (.Y(_03622_),
    .A(\top_ihp.oisc.regs[57][4] ),
    .B(net599));
 sg13g2_o21ai_1 _19488_ (.B1(_03622_),
    .Y(_02142_),
    .A1(net65),
    .A2(net598));
 sg13g2_nand2_1 _19489_ (.Y(_03623_),
    .A(\top_ihp.oisc.regs[57][5] ),
    .B(_03612_));
 sg13g2_o21ai_1 _19490_ (.B1(_03623_),
    .Y(_02143_),
    .A1(net73),
    .A2(_03615_));
 sg13g2_nand2_1 _19491_ (.Y(_03624_),
    .A(\top_ihp.oisc.regs[57][6] ),
    .B(net695));
 sg13g2_o21ai_1 _19492_ (.B1(_03624_),
    .Y(_02144_),
    .A1(net72),
    .A2(net598));
 sg13g2_nand2_1 _19493_ (.Y(_03625_),
    .A(\top_ihp.oisc.regs[57][7] ),
    .B(net695));
 sg13g2_o21ai_1 _19494_ (.B1(_03625_),
    .Y(_02145_),
    .A1(net470),
    .A2(net598));
 sg13g2_nand2_1 _19495_ (.Y(_03626_),
    .A(\top_ihp.oisc.regs[57][8] ),
    .B(_03589_));
 sg13g2_o21ai_1 _19496_ (.B1(_03626_),
    .Y(_02146_),
    .A1(net221),
    .A2(net694));
 sg13g2_nand2_1 _19497_ (.Y(_03627_),
    .A(\top_ihp.oisc.regs[57][9] ),
    .B(net695));
 sg13g2_o21ai_1 _19498_ (.B1(_03627_),
    .Y(_02147_),
    .A1(net71),
    .A2(net694));
 sg13g2_nand3_1 _19499_ (.B(_10522_),
    .C(_03146_),
    .A(_10519_),
    .Y(_03628_));
 sg13g2_buf_1 _19500_ (.A(_03628_),
    .X(_03629_));
 sg13g2_buf_1 _19501_ (.A(_03629_),
    .X(_03630_));
 sg13g2_buf_1 _19502_ (.A(net693),
    .X(_03631_));
 sg13g2_buf_1 _19503_ (.A(_03629_),
    .X(_03632_));
 sg13g2_nand2_1 _19504_ (.Y(_03633_),
    .A(\top_ihp.oisc.regs[58][0] ),
    .B(net692));
 sg13g2_o21ai_1 _19505_ (.B1(_03633_),
    .Y(_02148_),
    .A1(net70),
    .A2(net597));
 sg13g2_nand2_1 _19506_ (.Y(_03634_),
    .A(\top_ihp.oisc.regs[58][10] ),
    .B(net692));
 sg13g2_o21ai_1 _19507_ (.B1(_03634_),
    .Y(_02149_),
    .A1(net81),
    .A2(net597));
 sg13g2_nand2_1 _19508_ (.Y(_03635_),
    .A(\top_ihp.oisc.regs[58][11] ),
    .B(net692));
 sg13g2_o21ai_1 _19509_ (.B1(_03635_),
    .Y(_02150_),
    .A1(net69),
    .A2(net597));
 sg13g2_nand2_1 _19510_ (.Y(_03636_),
    .A(\top_ihp.oisc.regs[58][12] ),
    .B(net692));
 sg13g2_o21ai_1 _19511_ (.B1(_03636_),
    .Y(_02151_),
    .A1(net80),
    .A2(net597));
 sg13g2_nand2_1 _19512_ (.Y(_03637_),
    .A(\top_ihp.oisc.regs[58][13] ),
    .B(net692));
 sg13g2_o21ai_1 _19513_ (.B1(_03637_),
    .Y(_02152_),
    .A1(net79),
    .A2(net597));
 sg13g2_nand2_1 _19514_ (.Y(_03638_),
    .A(\top_ihp.oisc.regs[58][14] ),
    .B(net692));
 sg13g2_o21ai_1 _19515_ (.B1(_03638_),
    .Y(_02153_),
    .A1(net230),
    .A2(net597));
 sg13g2_nand2_1 _19516_ (.Y(_03639_),
    .A(\top_ihp.oisc.regs[58][15] ),
    .B(net692));
 sg13g2_o21ai_1 _19517_ (.B1(_03639_),
    .Y(_02154_),
    .A1(_03510_),
    .A2(net597));
 sg13g2_nand2_1 _19518_ (.Y(_03640_),
    .A(\top_ihp.oisc.regs[58][16] ),
    .B(_03632_));
 sg13g2_o21ai_1 _19519_ (.B1(_03640_),
    .Y(_02155_),
    .A1(net78),
    .A2(net597));
 sg13g2_buf_1 _19520_ (.A(net693),
    .X(_03641_));
 sg13g2_nand2_1 _19521_ (.Y(_03642_),
    .A(\top_ihp.oisc.regs[58][17] ),
    .B(net596));
 sg13g2_o21ai_1 _19522_ (.B1(_03642_),
    .Y(_02156_),
    .A1(_03453_),
    .A2(_03631_));
 sg13g2_nand2_1 _19523_ (.Y(_03643_),
    .A(\top_ihp.oisc.regs[58][18] ),
    .B(net596));
 sg13g2_o21ai_1 _19524_ (.B1(_03643_),
    .Y(_02157_),
    .A1(net228),
    .A2(_03631_));
 sg13g2_buf_1 _19525_ (.A(net693),
    .X(_03644_));
 sg13g2_nand2_1 _19526_ (.Y(_03645_),
    .A(\top_ihp.oisc.regs[58][19] ),
    .B(net596));
 sg13g2_o21ai_1 _19527_ (.B1(_03645_),
    .Y(_02158_),
    .A1(net77),
    .A2(net595));
 sg13g2_nand2_1 _19528_ (.Y(_03646_),
    .A(\top_ihp.oisc.regs[58][1] ),
    .B(_03641_));
 sg13g2_o21ai_1 _19529_ (.B1(_03646_),
    .Y(_02159_),
    .A1(net76),
    .A2(net595));
 sg13g2_nand2_1 _19530_ (.Y(_03647_),
    .A(\top_ihp.oisc.regs[58][20] ),
    .B(net596));
 sg13g2_o21ai_1 _19531_ (.B1(_03647_),
    .Y(_02160_),
    .A1(_10152_),
    .A2(net595));
 sg13g2_nand2_1 _19532_ (.Y(_03648_),
    .A(\top_ihp.oisc.regs[58][21] ),
    .B(net596));
 sg13g2_o21ai_1 _19533_ (.B1(_03648_),
    .Y(_02161_),
    .A1(net227),
    .A2(net595));
 sg13g2_nand2_1 _19534_ (.Y(_03649_),
    .A(\top_ihp.oisc.regs[58][22] ),
    .B(net596));
 sg13g2_o21ai_1 _19535_ (.B1(_03649_),
    .Y(_02162_),
    .A1(net75),
    .A2(net595));
 sg13g2_nand2_1 _19536_ (.Y(_03650_),
    .A(\top_ihp.oisc.regs[58][23] ),
    .B(net596));
 sg13g2_o21ai_1 _19537_ (.B1(_03650_),
    .Y(_02163_),
    .A1(net226),
    .A2(net595));
 sg13g2_nand2_1 _19538_ (.Y(_03651_),
    .A(\top_ihp.oisc.regs[58][24] ),
    .B(_03641_));
 sg13g2_o21ai_1 _19539_ (.B1(_03651_),
    .Y(_02164_),
    .A1(_03470_),
    .A2(_03644_));
 sg13g2_nand2_1 _19540_ (.Y(_03652_),
    .A(\top_ihp.oisc.regs[58][25] ),
    .B(net596));
 sg13g2_o21ai_1 _19541_ (.B1(_03652_),
    .Y(_02165_),
    .A1(net74),
    .A2(net595));
 sg13g2_buf_1 _19542_ (.A(net693),
    .X(_03653_));
 sg13g2_nand2_1 _19543_ (.Y(_03654_),
    .A(\top_ihp.oisc.regs[58][26] ),
    .B(net594));
 sg13g2_o21ai_1 _19544_ (.B1(_03654_),
    .Y(_02166_),
    .A1(net28),
    .A2(net595));
 sg13g2_nand2_1 _19545_ (.Y(_03655_),
    .A(\top_ihp.oisc.regs[58][27] ),
    .B(net594));
 sg13g2_o21ai_1 _19546_ (.B1(_03655_),
    .Y(_02167_),
    .A1(net224),
    .A2(_03644_));
 sg13g2_buf_1 _19547_ (.A(net693),
    .X(_03656_));
 sg13g2_nand2_1 _19548_ (.Y(_03657_),
    .A(\top_ihp.oisc.regs[58][28] ),
    .B(net594));
 sg13g2_o21ai_1 _19549_ (.B1(_03657_),
    .Y(_02168_),
    .A1(net223),
    .A2(net593));
 sg13g2_nand2_1 _19550_ (.Y(_03658_),
    .A(\top_ihp.oisc.regs[58][29] ),
    .B(_03653_));
 sg13g2_o21ai_1 _19551_ (.B1(_03658_),
    .Y(_02169_),
    .A1(_03482_),
    .A2(_03656_));
 sg13g2_nand2_1 _19552_ (.Y(_03659_),
    .A(\top_ihp.oisc.regs[58][2] ),
    .B(net594));
 sg13g2_o21ai_1 _19553_ (.B1(_03659_),
    .Y(_02170_),
    .A1(_03532_),
    .A2(net593));
 sg13g2_nand2_1 _19554_ (.Y(_03660_),
    .A(\top_ihp.oisc.regs[58][30] ),
    .B(net594));
 sg13g2_o21ai_1 _19555_ (.B1(_03660_),
    .Y(_02171_),
    .A1(net67),
    .A2(net593));
 sg13g2_nand2_1 _19556_ (.Y(_03661_),
    .A(\top_ihp.oisc.regs[58][31] ),
    .B(net594));
 sg13g2_o21ai_1 _19557_ (.B1(_03661_),
    .Y(_02172_),
    .A1(_10348_),
    .A2(net593));
 sg13g2_nand2_1 _19558_ (.Y(_03662_),
    .A(\top_ihp.oisc.regs[58][3] ),
    .B(net594));
 sg13g2_o21ai_1 _19559_ (.B1(_03662_),
    .Y(_02173_),
    .A1(net66),
    .A2(net593));
 sg13g2_nand2_1 _19560_ (.Y(_03663_),
    .A(\top_ihp.oisc.regs[58][4] ),
    .B(net594));
 sg13g2_o21ai_1 _19561_ (.B1(_03663_),
    .Y(_02174_),
    .A1(net65),
    .A2(net593));
 sg13g2_nand2_1 _19562_ (.Y(_03664_),
    .A(\top_ihp.oisc.regs[58][5] ),
    .B(_03653_));
 sg13g2_o21ai_1 _19563_ (.B1(_03664_),
    .Y(_02175_),
    .A1(net73),
    .A2(net593));
 sg13g2_nand2_1 _19564_ (.Y(_03665_),
    .A(\top_ihp.oisc.regs[58][6] ),
    .B(net693));
 sg13g2_o21ai_1 _19565_ (.B1(_03665_),
    .Y(_02176_),
    .A1(net72),
    .A2(net593));
 sg13g2_nand2_1 _19566_ (.Y(_03666_),
    .A(\top_ihp.oisc.regs[58][7] ),
    .B(_03630_));
 sg13g2_o21ai_1 _19567_ (.B1(_03666_),
    .Y(_02177_),
    .A1(_10483_),
    .A2(_03656_));
 sg13g2_nand2_1 _19568_ (.Y(_03667_),
    .A(\top_ihp.oisc.regs[58][8] ),
    .B(net693));
 sg13g2_o21ai_1 _19569_ (.B1(_03667_),
    .Y(_02178_),
    .A1(net221),
    .A2(_03632_));
 sg13g2_nand2_1 _19570_ (.Y(_03668_),
    .A(\top_ihp.oisc.regs[58][9] ),
    .B(net693));
 sg13g2_o21ai_1 _19571_ (.B1(_03668_),
    .Y(_02179_),
    .A1(net71),
    .A2(net692));
 sg13g2_nand2_1 _19572_ (.Y(_03669_),
    .A(_10520_),
    .B(_03313_));
 sg13g2_buf_1 _19573_ (.A(_03669_),
    .X(_03670_));
 sg13g2_buf_1 _19574_ (.A(net691),
    .X(_03671_));
 sg13g2_buf_1 _19575_ (.A(_03669_),
    .X(_03672_));
 sg13g2_nand2_1 _19576_ (.Y(_03673_),
    .A(\top_ihp.oisc.regs[59][0] ),
    .B(_03672_));
 sg13g2_o21ai_1 _19577_ (.B1(_03673_),
    .Y(_02180_),
    .A1(net70),
    .A2(net592));
 sg13g2_nand2_1 _19578_ (.Y(_03674_),
    .A(\top_ihp.oisc.regs[59][10] ),
    .B(net690));
 sg13g2_o21ai_1 _19579_ (.B1(_03674_),
    .Y(_02181_),
    .A1(net81),
    .A2(net592));
 sg13g2_nand2_1 _19580_ (.Y(_03675_),
    .A(\top_ihp.oisc.regs[59][11] ),
    .B(_03672_));
 sg13g2_o21ai_1 _19581_ (.B1(_03675_),
    .Y(_02182_),
    .A1(net69),
    .A2(_03671_));
 sg13g2_nand2_1 _19582_ (.Y(_03676_),
    .A(\top_ihp.oisc.regs[59][12] ),
    .B(net690));
 sg13g2_o21ai_1 _19583_ (.B1(_03676_),
    .Y(_02183_),
    .A1(net80),
    .A2(net592));
 sg13g2_nand2_1 _19584_ (.Y(_03677_),
    .A(\top_ihp.oisc.regs[59][13] ),
    .B(net690));
 sg13g2_o21ai_1 _19585_ (.B1(_03677_),
    .Y(_02184_),
    .A1(net79),
    .A2(net592));
 sg13g2_nand2_1 _19586_ (.Y(_03678_),
    .A(\top_ihp.oisc.regs[59][14] ),
    .B(net690));
 sg13g2_o21ai_1 _19587_ (.B1(_03678_),
    .Y(_02185_),
    .A1(net230),
    .A2(net592));
 sg13g2_nand2_1 _19588_ (.Y(_03679_),
    .A(\top_ihp.oisc.regs[59][15] ),
    .B(net690));
 sg13g2_o21ai_1 _19589_ (.B1(_03679_),
    .Y(_02186_),
    .A1(net220),
    .A2(net592));
 sg13g2_nand2_1 _19590_ (.Y(_03680_),
    .A(\top_ihp.oisc.regs[59][16] ),
    .B(net690));
 sg13g2_o21ai_1 _19591_ (.B1(_03680_),
    .Y(_02187_),
    .A1(net78),
    .A2(net592));
 sg13g2_buf_1 _19592_ (.A(net691),
    .X(_03681_));
 sg13g2_nand2_1 _19593_ (.Y(_03682_),
    .A(\top_ihp.oisc.regs[59][17] ),
    .B(net591));
 sg13g2_o21ai_1 _19594_ (.B1(_03682_),
    .Y(_02188_),
    .A1(net229),
    .A2(net592));
 sg13g2_nand2_1 _19595_ (.Y(_03683_),
    .A(\top_ihp.oisc.regs[59][18] ),
    .B(net591));
 sg13g2_o21ai_1 _19596_ (.B1(_03683_),
    .Y(_02189_),
    .A1(_03456_),
    .A2(_03671_));
 sg13g2_buf_1 _19597_ (.A(net691),
    .X(_03684_));
 sg13g2_nand2_1 _19598_ (.Y(_03685_),
    .A(\top_ihp.oisc.regs[59][19] ),
    .B(_03681_));
 sg13g2_o21ai_1 _19599_ (.B1(_03685_),
    .Y(_02190_),
    .A1(net77),
    .A2(_03684_));
 sg13g2_nand2_1 _19600_ (.Y(_03686_),
    .A(\top_ihp.oisc.regs[59][1] ),
    .B(net591));
 sg13g2_o21ai_1 _19601_ (.B1(_03686_),
    .Y(_02191_),
    .A1(net76),
    .A2(net590));
 sg13g2_nand2_1 _19602_ (.Y(_03687_),
    .A(\top_ihp.oisc.regs[59][20] ),
    .B(_03681_));
 sg13g2_o21ai_1 _19603_ (.B1(_03687_),
    .Y(_02192_),
    .A1(net607),
    .A2(_03684_));
 sg13g2_nand2_1 _19604_ (.Y(_03688_),
    .A(\top_ihp.oisc.regs[59][21] ),
    .B(net591));
 sg13g2_o21ai_1 _19605_ (.B1(_03688_),
    .Y(_02193_),
    .A1(net227),
    .A2(net590));
 sg13g2_nand2_1 _19606_ (.Y(_03689_),
    .A(\top_ihp.oisc.regs[59][22] ),
    .B(net591));
 sg13g2_o21ai_1 _19607_ (.B1(_03689_),
    .Y(_02194_),
    .A1(net75),
    .A2(net590));
 sg13g2_nand2_1 _19608_ (.Y(_03690_),
    .A(\top_ihp.oisc.regs[59][23] ),
    .B(net591));
 sg13g2_o21ai_1 _19609_ (.B1(_03690_),
    .Y(_02195_),
    .A1(net226),
    .A2(net590));
 sg13g2_nand2_1 _19610_ (.Y(_03691_),
    .A(\top_ihp.oisc.regs[59][24] ),
    .B(net591));
 sg13g2_o21ai_1 _19611_ (.B1(_03691_),
    .Y(_02196_),
    .A1(net225),
    .A2(net590));
 sg13g2_nand2_1 _19612_ (.Y(_03692_),
    .A(\top_ihp.oisc.regs[59][25] ),
    .B(net591));
 sg13g2_o21ai_1 _19613_ (.B1(_03692_),
    .Y(_02197_),
    .A1(net74),
    .A2(net590));
 sg13g2_buf_1 _19614_ (.A(net691),
    .X(_03693_));
 sg13g2_nand2_1 _19615_ (.Y(_03694_),
    .A(\top_ihp.oisc.regs[59][26] ),
    .B(net589));
 sg13g2_o21ai_1 _19616_ (.B1(_03694_),
    .Y(_02198_),
    .A1(net28),
    .A2(net590));
 sg13g2_nand2_1 _19617_ (.Y(_03695_),
    .A(\top_ihp.oisc.regs[59][27] ),
    .B(net589));
 sg13g2_o21ai_1 _19618_ (.B1(_03695_),
    .Y(_02199_),
    .A1(net224),
    .A2(net590));
 sg13g2_buf_1 _19619_ (.A(net691),
    .X(_03696_));
 sg13g2_nand2_1 _19620_ (.Y(_03697_),
    .A(\top_ihp.oisc.regs[59][28] ),
    .B(net589));
 sg13g2_o21ai_1 _19621_ (.B1(_03697_),
    .Y(_02200_),
    .A1(net223),
    .A2(net588));
 sg13g2_nand2_1 _19622_ (.Y(_03698_),
    .A(\top_ihp.oisc.regs[59][29] ),
    .B(net589));
 sg13g2_o21ai_1 _19623_ (.B1(_03698_),
    .Y(_02201_),
    .A1(net222),
    .A2(net588));
 sg13g2_nand2_1 _19624_ (.Y(_03699_),
    .A(\top_ihp.oisc.regs[59][2] ),
    .B(net589));
 sg13g2_o21ai_1 _19625_ (.B1(_03699_),
    .Y(_02202_),
    .A1(net68),
    .A2(_03696_));
 sg13g2_nand2_1 _19626_ (.Y(_03700_),
    .A(\top_ihp.oisc.regs[59][30] ),
    .B(_03693_));
 sg13g2_o21ai_1 _19627_ (.B1(_03700_),
    .Y(_02203_),
    .A1(net67),
    .A2(_03696_));
 sg13g2_nand2_1 _19628_ (.Y(_03701_),
    .A(\top_ihp.oisc.regs[59][31] ),
    .B(net589));
 sg13g2_o21ai_1 _19629_ (.B1(_03701_),
    .Y(_02204_),
    .A1(net306),
    .A2(net588));
 sg13g2_nand2_1 _19630_ (.Y(_03702_),
    .A(\top_ihp.oisc.regs[59][3] ),
    .B(net589));
 sg13g2_o21ai_1 _19631_ (.B1(_03702_),
    .Y(_02205_),
    .A1(net66),
    .A2(net588));
 sg13g2_nand2_1 _19632_ (.Y(_03703_),
    .A(\top_ihp.oisc.regs[59][4] ),
    .B(net589));
 sg13g2_o21ai_1 _19633_ (.B1(_03703_),
    .Y(_02206_),
    .A1(net65),
    .A2(net588));
 sg13g2_nand2_1 _19634_ (.Y(_03704_),
    .A(\top_ihp.oisc.regs[59][5] ),
    .B(_03693_));
 sg13g2_o21ai_1 _19635_ (.B1(_03704_),
    .Y(_02207_),
    .A1(net73),
    .A2(net588));
 sg13g2_nand2_1 _19636_ (.Y(_03705_),
    .A(\top_ihp.oisc.regs[59][6] ),
    .B(net691));
 sg13g2_o21ai_1 _19637_ (.B1(_03705_),
    .Y(_02208_),
    .A1(net72),
    .A2(net588));
 sg13g2_nand2_1 _19638_ (.Y(_03706_),
    .A(\top_ihp.oisc.regs[59][7] ),
    .B(net691));
 sg13g2_o21ai_1 _19639_ (.B1(_03706_),
    .Y(_02209_),
    .A1(net470),
    .A2(net588));
 sg13g2_nand2_1 _19640_ (.Y(_03707_),
    .A(\top_ihp.oisc.regs[59][8] ),
    .B(_03670_));
 sg13g2_o21ai_1 _19641_ (.B1(_03707_),
    .Y(_02210_),
    .A1(net221),
    .A2(net690));
 sg13g2_nand2_1 _19642_ (.Y(_03708_),
    .A(\top_ihp.oisc.regs[59][9] ),
    .B(net691));
 sg13g2_o21ai_1 _19643_ (.B1(_03708_),
    .Y(_02211_),
    .A1(_03496_),
    .A2(net690));
 sg13g2_nand2_1 _19644_ (.Y(_03709_),
    .A(_10651_),
    .B(net762));
 sg13g2_buf_1 _19645_ (.A(_03709_),
    .X(_03710_));
 sg13g2_buf_1 _19646_ (.A(net733),
    .X(_03711_));
 sg13g2_buf_1 _19647_ (.A(_03709_),
    .X(_03712_));
 sg13g2_nand2_1 _19648_ (.Y(_03713_),
    .A(\top_ihp.oisc.regs[5][0] ),
    .B(net732));
 sg13g2_o21ai_1 _19649_ (.B1(_03713_),
    .Y(_02212_),
    .A1(net70),
    .A2(net689));
 sg13g2_nand2_1 _19650_ (.Y(_03714_),
    .A(\top_ihp.oisc.regs[5][10] ),
    .B(net732));
 sg13g2_o21ai_1 _19651_ (.B1(_03714_),
    .Y(_02213_),
    .A1(_03441_),
    .A2(net689));
 sg13g2_nand2_1 _19652_ (.Y(_03715_),
    .A(\top_ihp.oisc.regs[5][11] ),
    .B(net732));
 sg13g2_o21ai_1 _19653_ (.B1(_03715_),
    .Y(_02214_),
    .A1(_03505_),
    .A2(net689));
 sg13g2_nand2_1 _19654_ (.Y(_03716_),
    .A(\top_ihp.oisc.regs[5][12] ),
    .B(net732));
 sg13g2_o21ai_1 _19655_ (.B1(_03716_),
    .Y(_02215_),
    .A1(_03444_),
    .A2(net689));
 sg13g2_nand2_1 _19656_ (.Y(_03717_),
    .A(\top_ihp.oisc.regs[5][13] ),
    .B(net732));
 sg13g2_o21ai_1 _19657_ (.B1(_03717_),
    .Y(_02216_),
    .A1(_03446_),
    .A2(_03711_));
 sg13g2_nand2_1 _19658_ (.Y(_03718_),
    .A(\top_ihp.oisc.regs[5][14] ),
    .B(net732));
 sg13g2_o21ai_1 _19659_ (.B1(_03718_),
    .Y(_02217_),
    .A1(_03448_),
    .A2(net689));
 sg13g2_nand2_1 _19660_ (.Y(_03719_),
    .A(\top_ihp.oisc.regs[5][15] ),
    .B(net732));
 sg13g2_o21ai_1 _19661_ (.B1(_03719_),
    .Y(_02218_),
    .A1(_03510_),
    .A2(net689));
 sg13g2_nand2_1 _19662_ (.Y(_03720_),
    .A(\top_ihp.oisc.regs[5][16] ),
    .B(net732));
 sg13g2_o21ai_1 _19663_ (.B1(_03720_),
    .Y(_02219_),
    .A1(_03451_),
    .A2(_03711_));
 sg13g2_buf_1 _19664_ (.A(net733),
    .X(_03721_));
 sg13g2_nand2_1 _19665_ (.Y(_03722_),
    .A(\top_ihp.oisc.regs[5][17] ),
    .B(net688));
 sg13g2_o21ai_1 _19666_ (.B1(_03722_),
    .Y(_02220_),
    .A1(_03453_),
    .A2(net689));
 sg13g2_nand2_1 _19667_ (.Y(_03723_),
    .A(\top_ihp.oisc.regs[5][18] ),
    .B(net688));
 sg13g2_o21ai_1 _19668_ (.B1(_03723_),
    .Y(_02221_),
    .A1(_03456_),
    .A2(net689));
 sg13g2_buf_1 _19669_ (.A(net733),
    .X(_03724_));
 sg13g2_nand2_1 _19670_ (.Y(_03725_),
    .A(\top_ihp.oisc.regs[5][19] ),
    .B(net688));
 sg13g2_o21ai_1 _19671_ (.B1(_03725_),
    .Y(_02222_),
    .A1(net77),
    .A2(net687));
 sg13g2_nand2_1 _19672_ (.Y(_03726_),
    .A(\top_ihp.oisc.regs[5][1] ),
    .B(net688));
 sg13g2_o21ai_1 _19673_ (.B1(_03726_),
    .Y(_02223_),
    .A1(net76),
    .A2(net687));
 sg13g2_nand2_1 _19674_ (.Y(_03727_),
    .A(\top_ihp.oisc.regs[5][20] ),
    .B(net688));
 sg13g2_o21ai_1 _19675_ (.B1(_03727_),
    .Y(_02224_),
    .A1(net607),
    .A2(net687));
 sg13g2_nand2_1 _19676_ (.Y(_03728_),
    .A(\top_ihp.oisc.regs[5][21] ),
    .B(net688));
 sg13g2_o21ai_1 _19677_ (.B1(_03728_),
    .Y(_02225_),
    .A1(_03464_),
    .A2(net687));
 sg13g2_nand2_1 _19678_ (.Y(_03729_),
    .A(\top_ihp.oisc.regs[5][22] ),
    .B(net688));
 sg13g2_o21ai_1 _19679_ (.B1(_03729_),
    .Y(_02226_),
    .A1(net75),
    .A2(net687));
 sg13g2_nand2_1 _19680_ (.Y(_03730_),
    .A(\top_ihp.oisc.regs[5][23] ),
    .B(net688));
 sg13g2_o21ai_1 _19681_ (.B1(_03730_),
    .Y(_02227_),
    .A1(net226),
    .A2(net687));
 sg13g2_nand2_1 _19682_ (.Y(_03731_),
    .A(\top_ihp.oisc.regs[5][24] ),
    .B(_03721_));
 sg13g2_o21ai_1 _19683_ (.B1(_03731_),
    .Y(_02228_),
    .A1(net225),
    .A2(_03724_));
 sg13g2_nand2_1 _19684_ (.Y(_03732_),
    .A(\top_ihp.oisc.regs[5][25] ),
    .B(_03721_));
 sg13g2_o21ai_1 _19685_ (.B1(_03732_),
    .Y(_02229_),
    .A1(net74),
    .A2(net687));
 sg13g2_buf_1 _19686_ (.A(net733),
    .X(_03733_));
 sg13g2_nand2_1 _19687_ (.Y(_03734_),
    .A(\top_ihp.oisc.regs[5][26] ),
    .B(net686));
 sg13g2_o21ai_1 _19688_ (.B1(_03734_),
    .Y(_02230_),
    .A1(net28),
    .A2(_03724_));
 sg13g2_nand2_1 _19689_ (.Y(_03735_),
    .A(\top_ihp.oisc.regs[5][27] ),
    .B(net686));
 sg13g2_o21ai_1 _19690_ (.B1(_03735_),
    .Y(_02231_),
    .A1(_03477_),
    .A2(net687));
 sg13g2_buf_1 _19691_ (.A(net733),
    .X(_03736_));
 sg13g2_nand2_1 _19692_ (.Y(_03737_),
    .A(\top_ihp.oisc.regs[5][28] ),
    .B(_03733_));
 sg13g2_o21ai_1 _19693_ (.B1(_03737_),
    .Y(_02232_),
    .A1(net223),
    .A2(net685));
 sg13g2_nand2_1 _19694_ (.Y(_03738_),
    .A(\top_ihp.oisc.regs[5][29] ),
    .B(_03733_));
 sg13g2_o21ai_1 _19695_ (.B1(_03738_),
    .Y(_02233_),
    .A1(net222),
    .A2(_03736_));
 sg13g2_nand2_1 _19696_ (.Y(_03739_),
    .A(\top_ihp.oisc.regs[5][2] ),
    .B(net686));
 sg13g2_o21ai_1 _19697_ (.B1(_03739_),
    .Y(_02234_),
    .A1(net68),
    .A2(_03736_));
 sg13g2_nand2_1 _19698_ (.Y(_03740_),
    .A(\top_ihp.oisc.regs[5][30] ),
    .B(net686));
 sg13g2_o21ai_1 _19699_ (.B1(_03740_),
    .Y(_02235_),
    .A1(net67),
    .A2(net685));
 sg13g2_nand2_1 _19700_ (.Y(_03741_),
    .A(\top_ihp.oisc.regs[5][31] ),
    .B(net686));
 sg13g2_o21ai_1 _19701_ (.B1(_03741_),
    .Y(_02236_),
    .A1(net306),
    .A2(net685));
 sg13g2_nand2_1 _19702_ (.Y(_03742_),
    .A(\top_ihp.oisc.regs[5][3] ),
    .B(net686));
 sg13g2_o21ai_1 _19703_ (.B1(_03742_),
    .Y(_02237_),
    .A1(_03537_),
    .A2(net685));
 sg13g2_nand2_1 _19704_ (.Y(_03743_),
    .A(\top_ihp.oisc.regs[5][4] ),
    .B(net686));
 sg13g2_o21ai_1 _19705_ (.B1(_03743_),
    .Y(_02238_),
    .A1(net65),
    .A2(net685));
 sg13g2_nand2_1 _19706_ (.Y(_03744_),
    .A(\top_ihp.oisc.regs[5][5] ),
    .B(net686));
 sg13g2_o21ai_1 _19707_ (.B1(_03744_),
    .Y(_02239_),
    .A1(_03489_),
    .A2(net685));
 sg13g2_nand2_1 _19708_ (.Y(_03745_),
    .A(\top_ihp.oisc.regs[5][6] ),
    .B(net733));
 sg13g2_o21ai_1 _19709_ (.B1(_03745_),
    .Y(_02240_),
    .A1(net72),
    .A2(net685));
 sg13g2_nand2_1 _19710_ (.Y(_03746_),
    .A(\top_ihp.oisc.regs[5][7] ),
    .B(net733));
 sg13g2_o21ai_1 _19711_ (.B1(_03746_),
    .Y(_02241_),
    .A1(net470),
    .A2(net685));
 sg13g2_nand2_1 _19712_ (.Y(_03747_),
    .A(\top_ihp.oisc.regs[5][8] ),
    .B(_03710_));
 sg13g2_o21ai_1 _19713_ (.B1(_03747_),
    .Y(_02242_),
    .A1(_03494_),
    .A2(_03712_));
 sg13g2_nand2_1 _19714_ (.Y(_03748_),
    .A(\top_ihp.oisc.regs[5][9] ),
    .B(net733));
 sg13g2_o21ai_1 _19715_ (.B1(_03748_),
    .Y(_02243_),
    .A1(_03496_),
    .A2(_03712_));
 sg13g2_nand2_1 _19716_ (.Y(_03749_),
    .A(_10619_),
    .B(_03148_));
 sg13g2_buf_1 _19717_ (.A(_03749_),
    .X(_03750_));
 sg13g2_buf_1 _19718_ (.A(net587),
    .X(_03751_));
 sg13g2_buf_2 _19719_ (.A(_03749_),
    .X(_03752_));
 sg13g2_nand2_1 _19720_ (.Y(_03753_),
    .A(\top_ihp.oisc.regs[60][0] ),
    .B(net586));
 sg13g2_o21ai_1 _19721_ (.B1(_03753_),
    .Y(_02244_),
    .A1(net70),
    .A2(net464));
 sg13g2_nand2_1 _19722_ (.Y(_03754_),
    .A(\top_ihp.oisc.regs[60][10] ),
    .B(net586));
 sg13g2_o21ai_1 _19723_ (.B1(_03754_),
    .Y(_02245_),
    .A1(net81),
    .A2(net464));
 sg13g2_nand2_1 _19724_ (.Y(_03755_),
    .A(\top_ihp.oisc.regs[60][11] ),
    .B(net586));
 sg13g2_o21ai_1 _19725_ (.B1(_03755_),
    .Y(_02246_),
    .A1(net69),
    .A2(net464));
 sg13g2_nand2_1 _19726_ (.Y(_03756_),
    .A(\top_ihp.oisc.regs[60][12] ),
    .B(net586));
 sg13g2_o21ai_1 _19727_ (.B1(_03756_),
    .Y(_02247_),
    .A1(net80),
    .A2(net464));
 sg13g2_nand2_1 _19728_ (.Y(_03757_),
    .A(\top_ihp.oisc.regs[60][13] ),
    .B(_03752_));
 sg13g2_o21ai_1 _19729_ (.B1(_03757_),
    .Y(_02248_),
    .A1(_03446_),
    .A2(net464));
 sg13g2_nand2_1 _19730_ (.Y(_03758_),
    .A(\top_ihp.oisc.regs[60][14] ),
    .B(net586));
 sg13g2_o21ai_1 _19731_ (.B1(_03758_),
    .Y(_02249_),
    .A1(net230),
    .A2(net464));
 sg13g2_nand2_1 _19732_ (.Y(_03759_),
    .A(\top_ihp.oisc.regs[60][15] ),
    .B(net586));
 sg13g2_o21ai_1 _19733_ (.B1(_03759_),
    .Y(_02250_),
    .A1(net220),
    .A2(net464));
 sg13g2_nand2_1 _19734_ (.Y(_03760_),
    .A(\top_ihp.oisc.regs[60][16] ),
    .B(_03752_));
 sg13g2_o21ai_1 _19735_ (.B1(_03760_),
    .Y(_02251_),
    .A1(_03451_),
    .A2(net464));
 sg13g2_buf_1 _19736_ (.A(net587),
    .X(_03761_));
 sg13g2_nand2_1 _19737_ (.Y(_03762_),
    .A(\top_ihp.oisc.regs[60][17] ),
    .B(net463));
 sg13g2_o21ai_1 _19738_ (.B1(_03762_),
    .Y(_02252_),
    .A1(net229),
    .A2(_03751_));
 sg13g2_nand2_1 _19739_ (.Y(_03763_),
    .A(\top_ihp.oisc.regs[60][18] ),
    .B(net463));
 sg13g2_o21ai_1 _19740_ (.B1(_03763_),
    .Y(_02253_),
    .A1(net228),
    .A2(_03751_));
 sg13g2_buf_1 _19741_ (.A(net587),
    .X(_03764_));
 sg13g2_nand2_1 _19742_ (.Y(_03765_),
    .A(\top_ihp.oisc.regs[60][19] ),
    .B(net463));
 sg13g2_o21ai_1 _19743_ (.B1(_03765_),
    .Y(_02254_),
    .A1(net77),
    .A2(net462));
 sg13g2_nand2_1 _19744_ (.Y(_03766_),
    .A(\top_ihp.oisc.regs[60][1] ),
    .B(net463));
 sg13g2_o21ai_1 _19745_ (.B1(_03766_),
    .Y(_02255_),
    .A1(_03461_),
    .A2(net462));
 sg13g2_nand2_1 _19746_ (.Y(_03767_),
    .A(\top_ihp.oisc.regs[60][20] ),
    .B(net463));
 sg13g2_o21ai_1 _19747_ (.B1(_03767_),
    .Y(_02256_),
    .A1(_03519_),
    .A2(net462));
 sg13g2_nand2_1 _19748_ (.Y(_03768_),
    .A(\top_ihp.oisc.regs[60][21] ),
    .B(net463));
 sg13g2_o21ai_1 _19749_ (.B1(_03768_),
    .Y(_02257_),
    .A1(net227),
    .A2(net462));
 sg13g2_nand2_1 _19750_ (.Y(_03769_),
    .A(\top_ihp.oisc.regs[60][22] ),
    .B(net463));
 sg13g2_o21ai_1 _19751_ (.B1(_03769_),
    .Y(_02258_),
    .A1(net75),
    .A2(net462));
 sg13g2_nand2_1 _19752_ (.Y(_03770_),
    .A(\top_ihp.oisc.regs[60][23] ),
    .B(_03761_));
 sg13g2_o21ai_1 _19753_ (.B1(_03770_),
    .Y(_02259_),
    .A1(net226),
    .A2(_03764_));
 sg13g2_nand2_1 _19754_ (.Y(_03771_),
    .A(\top_ihp.oisc.regs[60][24] ),
    .B(_03761_));
 sg13g2_o21ai_1 _19755_ (.B1(_03771_),
    .Y(_02260_),
    .A1(net225),
    .A2(_03764_));
 sg13g2_nand2_1 _19756_ (.Y(_03772_),
    .A(\top_ihp.oisc.regs[60][25] ),
    .B(net463));
 sg13g2_o21ai_1 _19757_ (.B1(_03772_),
    .Y(_02261_),
    .A1(net74),
    .A2(net462));
 sg13g2_buf_1 _19758_ (.A(net587),
    .X(_03773_));
 sg13g2_nand2_1 _19759_ (.Y(_03774_),
    .A(\top_ihp.oisc.regs[60][26] ),
    .B(net461));
 sg13g2_o21ai_1 _19760_ (.B1(_03774_),
    .Y(_02262_),
    .A1(net28),
    .A2(net462));
 sg13g2_nand2_1 _19761_ (.Y(_03775_),
    .A(\top_ihp.oisc.regs[60][27] ),
    .B(net461));
 sg13g2_o21ai_1 _19762_ (.B1(_03775_),
    .Y(_02263_),
    .A1(net224),
    .A2(net462));
 sg13g2_buf_1 _19763_ (.A(net587),
    .X(_03776_));
 sg13g2_nand2_1 _19764_ (.Y(_03777_),
    .A(\top_ihp.oisc.regs[60][28] ),
    .B(net461));
 sg13g2_o21ai_1 _19765_ (.B1(_03777_),
    .Y(_02264_),
    .A1(net223),
    .A2(net460));
 sg13g2_nand2_1 _19766_ (.Y(_03778_),
    .A(\top_ihp.oisc.regs[60][29] ),
    .B(_03773_));
 sg13g2_o21ai_1 _19767_ (.B1(_03778_),
    .Y(_02265_),
    .A1(net222),
    .A2(_03776_));
 sg13g2_nand2_1 _19768_ (.Y(_03779_),
    .A(\top_ihp.oisc.regs[60][2] ),
    .B(net461));
 sg13g2_o21ai_1 _19769_ (.B1(_03779_),
    .Y(_02266_),
    .A1(net68),
    .A2(net460));
 sg13g2_nand2_1 _19770_ (.Y(_03780_),
    .A(\top_ihp.oisc.regs[60][30] ),
    .B(net461));
 sg13g2_o21ai_1 _19771_ (.B1(_03780_),
    .Y(_02267_),
    .A1(net67),
    .A2(net460));
 sg13g2_nand2_1 _19772_ (.Y(_03781_),
    .A(\top_ihp.oisc.regs[60][31] ),
    .B(net461));
 sg13g2_o21ai_1 _19773_ (.B1(_03781_),
    .Y(_02268_),
    .A1(net306),
    .A2(net460));
 sg13g2_nand2_1 _19774_ (.Y(_03782_),
    .A(\top_ihp.oisc.regs[60][3] ),
    .B(net461));
 sg13g2_o21ai_1 _19775_ (.B1(_03782_),
    .Y(_02269_),
    .A1(net66),
    .A2(net460));
 sg13g2_nand2_1 _19776_ (.Y(_03783_),
    .A(\top_ihp.oisc.regs[60][4] ),
    .B(net461));
 sg13g2_o21ai_1 _19777_ (.B1(_03783_),
    .Y(_02270_),
    .A1(net65),
    .A2(net460));
 sg13g2_nand2_1 _19778_ (.Y(_03784_),
    .A(\top_ihp.oisc.regs[60][5] ),
    .B(_03773_));
 sg13g2_o21ai_1 _19779_ (.B1(_03784_),
    .Y(_02271_),
    .A1(_03489_),
    .A2(_03776_));
 sg13g2_nand2_1 _19780_ (.Y(_03785_),
    .A(\top_ihp.oisc.regs[60][6] ),
    .B(net587));
 sg13g2_o21ai_1 _19781_ (.B1(_03785_),
    .Y(_02272_),
    .A1(_03491_),
    .A2(net460));
 sg13g2_nand2_1 _19782_ (.Y(_03786_),
    .A(\top_ihp.oisc.regs[60][7] ),
    .B(_03750_));
 sg13g2_o21ai_1 _19783_ (.B1(_03786_),
    .Y(_02273_),
    .A1(_03543_),
    .A2(net460));
 sg13g2_nand2_1 _19784_ (.Y(_03787_),
    .A(\top_ihp.oisc.regs[60][8] ),
    .B(net587));
 sg13g2_o21ai_1 _19785_ (.B1(_03787_),
    .Y(_02274_),
    .A1(net221),
    .A2(net586));
 sg13g2_nand2_1 _19786_ (.Y(_03788_),
    .A(\top_ihp.oisc.regs[60][9] ),
    .B(net587));
 sg13g2_o21ai_1 _19787_ (.B1(_03788_),
    .Y(_02275_),
    .A1(net71),
    .A2(net586));
 sg13g2_or2_1 _19788_ (.X(_03789_),
    .B(_03189_),
    .A(_02961_));
 sg13g2_buf_1 _19789_ (.A(_03789_),
    .X(_03790_));
 sg13g2_buf_1 _19790_ (.A(_03790_),
    .X(_03791_));
 sg13g2_buf_2 _19791_ (.A(net684),
    .X(_03792_));
 sg13g2_buf_1 _19792_ (.A(_03790_),
    .X(_03793_));
 sg13g2_nand2_1 _19793_ (.Y(_03794_),
    .A(\top_ihp.oisc.regs[61][0] ),
    .B(net683));
 sg13g2_o21ai_1 _19794_ (.B1(_03794_),
    .Y(_02276_),
    .A1(_03498_),
    .A2(net585));
 sg13g2_nand2_1 _19795_ (.Y(_03795_),
    .A(\top_ihp.oisc.regs[61][10] ),
    .B(net683));
 sg13g2_o21ai_1 _19796_ (.B1(_03795_),
    .Y(_02277_),
    .A1(net81),
    .A2(net585));
 sg13g2_nand2_1 _19797_ (.Y(_03796_),
    .A(\top_ihp.oisc.regs[61][11] ),
    .B(net683));
 sg13g2_o21ai_1 _19798_ (.B1(_03796_),
    .Y(_02278_),
    .A1(net69),
    .A2(net585));
 sg13g2_nand2_1 _19799_ (.Y(_03797_),
    .A(\top_ihp.oisc.regs[61][12] ),
    .B(net683));
 sg13g2_o21ai_1 _19800_ (.B1(_03797_),
    .Y(_02279_),
    .A1(_03444_),
    .A2(net585));
 sg13g2_nand2_1 _19801_ (.Y(_03798_),
    .A(\top_ihp.oisc.regs[61][13] ),
    .B(_03793_));
 sg13g2_o21ai_1 _19802_ (.B1(_03798_),
    .Y(_02280_),
    .A1(net79),
    .A2(_03792_));
 sg13g2_nand2_1 _19803_ (.Y(_03799_),
    .A(\top_ihp.oisc.regs[61][14] ),
    .B(net683));
 sg13g2_o21ai_1 _19804_ (.B1(_03799_),
    .Y(_02281_),
    .A1(net230),
    .A2(net585));
 sg13g2_nand2_1 _19805_ (.Y(_03800_),
    .A(\top_ihp.oisc.regs[61][15] ),
    .B(net683));
 sg13g2_o21ai_1 _19806_ (.B1(_03800_),
    .Y(_02282_),
    .A1(net220),
    .A2(net585));
 sg13g2_nand2_1 _19807_ (.Y(_03801_),
    .A(\top_ihp.oisc.regs[61][16] ),
    .B(_03793_));
 sg13g2_o21ai_1 _19808_ (.B1(_03801_),
    .Y(_02283_),
    .A1(net78),
    .A2(net585));
 sg13g2_buf_1 _19809_ (.A(net684),
    .X(_03802_));
 sg13g2_nand2_1 _19810_ (.Y(_03803_),
    .A(\top_ihp.oisc.regs[61][17] ),
    .B(net584));
 sg13g2_o21ai_1 _19811_ (.B1(_03803_),
    .Y(_02284_),
    .A1(net229),
    .A2(net585));
 sg13g2_nand2_1 _19812_ (.Y(_03804_),
    .A(\top_ihp.oisc.regs[61][18] ),
    .B(net584));
 sg13g2_o21ai_1 _19813_ (.B1(_03804_),
    .Y(_02285_),
    .A1(net228),
    .A2(_03792_));
 sg13g2_buf_1 _19814_ (.A(net684),
    .X(_03805_));
 sg13g2_nand2_1 _19815_ (.Y(_03806_),
    .A(\top_ihp.oisc.regs[61][19] ),
    .B(net584));
 sg13g2_o21ai_1 _19816_ (.B1(_03806_),
    .Y(_02286_),
    .A1(_03458_),
    .A2(net583));
 sg13g2_nand2_1 _19817_ (.Y(_03807_),
    .A(\top_ihp.oisc.regs[61][1] ),
    .B(net584));
 sg13g2_o21ai_1 _19818_ (.B1(_03807_),
    .Y(_02287_),
    .A1(net76),
    .A2(net583));
 sg13g2_nand2_1 _19819_ (.Y(_03808_),
    .A(\top_ihp.oisc.regs[61][20] ),
    .B(net584));
 sg13g2_o21ai_1 _19820_ (.B1(_03808_),
    .Y(_02288_),
    .A1(_03519_),
    .A2(net583));
 sg13g2_nand2_1 _19821_ (.Y(_03809_),
    .A(\top_ihp.oisc.regs[61][21] ),
    .B(net584));
 sg13g2_o21ai_1 _19822_ (.B1(_03809_),
    .Y(_02289_),
    .A1(net227),
    .A2(net583));
 sg13g2_nand2_1 _19823_ (.Y(_03810_),
    .A(\top_ihp.oisc.regs[61][22] ),
    .B(net584));
 sg13g2_o21ai_1 _19824_ (.B1(_03810_),
    .Y(_02290_),
    .A1(_03466_),
    .A2(net583));
 sg13g2_nand2_1 _19825_ (.Y(_03811_),
    .A(\top_ihp.oisc.regs[61][23] ),
    .B(net584));
 sg13g2_o21ai_1 _19826_ (.B1(_03811_),
    .Y(_02291_),
    .A1(_03468_),
    .A2(net583));
 sg13g2_nand2_1 _19827_ (.Y(_03812_),
    .A(\top_ihp.oisc.regs[61][24] ),
    .B(_03802_));
 sg13g2_o21ai_1 _19828_ (.B1(_03812_),
    .Y(_02292_),
    .A1(net225),
    .A2(_03805_));
 sg13g2_nand2_1 _19829_ (.Y(_03813_),
    .A(\top_ihp.oisc.regs[61][25] ),
    .B(_03802_));
 sg13g2_o21ai_1 _19830_ (.B1(_03813_),
    .Y(_02293_),
    .A1(_03472_),
    .A2(_03805_));
 sg13g2_buf_1 _19831_ (.A(net684),
    .X(_03814_));
 sg13g2_nand2_1 _19832_ (.Y(_03815_),
    .A(\top_ihp.oisc.regs[61][26] ),
    .B(net582));
 sg13g2_o21ai_1 _19833_ (.B1(_03815_),
    .Y(_02294_),
    .A1(_03474_),
    .A2(net583));
 sg13g2_nand2_1 _19834_ (.Y(_03816_),
    .A(\top_ihp.oisc.regs[61][27] ),
    .B(net582));
 sg13g2_o21ai_1 _19835_ (.B1(_03816_),
    .Y(_02295_),
    .A1(_03477_),
    .A2(net583));
 sg13g2_buf_1 _19836_ (.A(_03791_),
    .X(_03817_));
 sg13g2_nand2_1 _19837_ (.Y(_03818_),
    .A(\top_ihp.oisc.regs[61][28] ),
    .B(_03814_));
 sg13g2_o21ai_1 _19838_ (.B1(_03818_),
    .Y(_02296_),
    .A1(_03479_),
    .A2(net581));
 sg13g2_nand2_1 _19839_ (.Y(_03819_),
    .A(\top_ihp.oisc.regs[61][29] ),
    .B(net582));
 sg13g2_o21ai_1 _19840_ (.B1(_03819_),
    .Y(_02297_),
    .A1(net222),
    .A2(net581));
 sg13g2_nand2_1 _19841_ (.Y(_03820_),
    .A(\top_ihp.oisc.regs[61][2] ),
    .B(net582));
 sg13g2_o21ai_1 _19842_ (.B1(_03820_),
    .Y(_02298_),
    .A1(net68),
    .A2(net581));
 sg13g2_nand2_1 _19843_ (.Y(_03821_),
    .A(\top_ihp.oisc.regs[61][30] ),
    .B(net582));
 sg13g2_o21ai_1 _19844_ (.B1(_03821_),
    .Y(_02299_),
    .A1(_03534_),
    .A2(net581));
 sg13g2_nand2_1 _19845_ (.Y(_03822_),
    .A(\top_ihp.oisc.regs[61][31] ),
    .B(net582));
 sg13g2_o21ai_1 _19846_ (.B1(_03822_),
    .Y(_02300_),
    .A1(_10644_),
    .A2(net581));
 sg13g2_nand2_1 _19847_ (.Y(_03823_),
    .A(\top_ihp.oisc.regs[61][3] ),
    .B(_03814_));
 sg13g2_o21ai_1 _19848_ (.B1(_03823_),
    .Y(_02301_),
    .A1(_03537_),
    .A2(_03817_));
 sg13g2_nand2_1 _19849_ (.Y(_03824_),
    .A(\top_ihp.oisc.regs[61][4] ),
    .B(net582));
 sg13g2_o21ai_1 _19850_ (.B1(_03824_),
    .Y(_02302_),
    .A1(_03539_),
    .A2(net581));
 sg13g2_nand2_1 _19851_ (.Y(_03825_),
    .A(\top_ihp.oisc.regs[61][5] ),
    .B(net582));
 sg13g2_o21ai_1 _19852_ (.B1(_03825_),
    .Y(_02303_),
    .A1(net73),
    .A2(net581));
 sg13g2_nand2_1 _19853_ (.Y(_03826_),
    .A(\top_ihp.oisc.regs[61][6] ),
    .B(net684));
 sg13g2_o21ai_1 _19854_ (.B1(_03826_),
    .Y(_02304_),
    .A1(net72),
    .A2(net581));
 sg13g2_nand2_1 _19855_ (.Y(_03827_),
    .A(\top_ihp.oisc.regs[61][7] ),
    .B(net684));
 sg13g2_o21ai_1 _19856_ (.B1(_03827_),
    .Y(_02305_),
    .A1(_03543_),
    .A2(_03817_));
 sg13g2_nand2_1 _19857_ (.Y(_03828_),
    .A(\top_ihp.oisc.regs[61][8] ),
    .B(net684));
 sg13g2_o21ai_1 _19858_ (.B1(_03828_),
    .Y(_02306_),
    .A1(net221),
    .A2(net683));
 sg13g2_nand2_1 _19859_ (.Y(_03829_),
    .A(\top_ihp.oisc.regs[61][9] ),
    .B(net684));
 sg13g2_o21ai_1 _19860_ (.B1(_03829_),
    .Y(_02307_),
    .A1(net71),
    .A2(net683));
 sg13g2_nand3_1 _19861_ (.B(_10618_),
    .C(_03146_),
    .A(_10870_),
    .Y(_03830_));
 sg13g2_buf_1 _19862_ (.A(_03830_),
    .X(_03831_));
 sg13g2_buf_1 _19863_ (.A(_03831_),
    .X(_03832_));
 sg13g2_buf_1 _19864_ (.A(net580),
    .X(_03833_));
 sg13g2_buf_1 _19865_ (.A(_03831_),
    .X(_03834_));
 sg13g2_nand2_1 _19866_ (.Y(_03835_),
    .A(\top_ihp.oisc.regs[62][0] ),
    .B(net579));
 sg13g2_o21ai_1 _19867_ (.B1(_03835_),
    .Y(_02308_),
    .A1(_03498_),
    .A2(net459));
 sg13g2_nand2_1 _19868_ (.Y(_03836_),
    .A(\top_ihp.oisc.regs[62][10] ),
    .B(net579));
 sg13g2_o21ai_1 _19869_ (.B1(_03836_),
    .Y(_02309_),
    .A1(_03441_),
    .A2(net459));
 sg13g2_nand2_1 _19870_ (.Y(_03837_),
    .A(\top_ihp.oisc.regs[62][11] ),
    .B(net579));
 sg13g2_o21ai_1 _19871_ (.B1(_03837_),
    .Y(_02310_),
    .A1(net69),
    .A2(net459));
 sg13g2_nand2_1 _19872_ (.Y(_03838_),
    .A(\top_ihp.oisc.regs[62][12] ),
    .B(net579));
 sg13g2_o21ai_1 _19873_ (.B1(_03838_),
    .Y(_02311_),
    .A1(net80),
    .A2(net459));
 sg13g2_nand2_1 _19874_ (.Y(_03839_),
    .A(\top_ihp.oisc.regs[62][13] ),
    .B(net579));
 sg13g2_o21ai_1 _19875_ (.B1(_03839_),
    .Y(_02312_),
    .A1(net79),
    .A2(net459));
 sg13g2_nand2_1 _19876_ (.Y(_03840_),
    .A(\top_ihp.oisc.regs[62][14] ),
    .B(net579));
 sg13g2_o21ai_1 _19877_ (.B1(_03840_),
    .Y(_02313_),
    .A1(net230),
    .A2(net459));
 sg13g2_nand2_1 _19878_ (.Y(_03841_),
    .A(\top_ihp.oisc.regs[62][15] ),
    .B(net579));
 sg13g2_o21ai_1 _19879_ (.B1(_03841_),
    .Y(_02314_),
    .A1(net220),
    .A2(net459));
 sg13g2_nand2_1 _19880_ (.Y(_03842_),
    .A(\top_ihp.oisc.regs[62][16] ),
    .B(net579));
 sg13g2_o21ai_1 _19881_ (.B1(_03842_),
    .Y(_02315_),
    .A1(net78),
    .A2(_03833_));
 sg13g2_buf_1 _19882_ (.A(net580),
    .X(_03843_));
 sg13g2_nand2_1 _19883_ (.Y(_03844_),
    .A(\top_ihp.oisc.regs[62][17] ),
    .B(net458));
 sg13g2_o21ai_1 _19884_ (.B1(_03844_),
    .Y(_02316_),
    .A1(net229),
    .A2(net459));
 sg13g2_nand2_1 _19885_ (.Y(_03845_),
    .A(\top_ihp.oisc.regs[62][18] ),
    .B(net458));
 sg13g2_o21ai_1 _19886_ (.B1(_03845_),
    .Y(_02317_),
    .A1(net228),
    .A2(_03833_));
 sg13g2_buf_1 _19887_ (.A(net580),
    .X(_03846_));
 sg13g2_nand2_1 _19888_ (.Y(_03847_),
    .A(\top_ihp.oisc.regs[62][19] ),
    .B(net458));
 sg13g2_o21ai_1 _19889_ (.B1(_03847_),
    .Y(_02318_),
    .A1(net77),
    .A2(net457));
 sg13g2_nand2_1 _19890_ (.Y(_03848_),
    .A(\top_ihp.oisc.regs[62][1] ),
    .B(net458));
 sg13g2_o21ai_1 _19891_ (.B1(_03848_),
    .Y(_02319_),
    .A1(_03461_),
    .A2(net457));
 sg13g2_nand2_1 _19892_ (.Y(_03849_),
    .A(\top_ihp.oisc.regs[62][20] ),
    .B(net458));
 sg13g2_o21ai_1 _19893_ (.B1(_03849_),
    .Y(_02320_),
    .A1(_10152_),
    .A2(net457));
 sg13g2_nand2_1 _19894_ (.Y(_03850_),
    .A(\top_ihp.oisc.regs[62][21] ),
    .B(net458));
 sg13g2_o21ai_1 _19895_ (.B1(_03850_),
    .Y(_02321_),
    .A1(_03464_),
    .A2(net457));
 sg13g2_nand2_1 _19896_ (.Y(_03851_),
    .A(\top_ihp.oisc.regs[62][22] ),
    .B(net458));
 sg13g2_o21ai_1 _19897_ (.B1(_03851_),
    .Y(_02322_),
    .A1(_03466_),
    .A2(net457));
 sg13g2_nand2_1 _19898_ (.Y(_03852_),
    .A(\top_ihp.oisc.regs[62][23] ),
    .B(_03843_));
 sg13g2_o21ai_1 _19899_ (.B1(_03852_),
    .Y(_02323_),
    .A1(_03468_),
    .A2(net457));
 sg13g2_nand2_1 _19900_ (.Y(_03853_),
    .A(\top_ihp.oisc.regs[62][24] ),
    .B(_03843_));
 sg13g2_o21ai_1 _19901_ (.B1(_03853_),
    .Y(_02324_),
    .A1(_03470_),
    .A2(_03846_));
 sg13g2_nand2_1 _19902_ (.Y(_03854_),
    .A(\top_ihp.oisc.regs[62][25] ),
    .B(net458));
 sg13g2_o21ai_1 _19903_ (.B1(_03854_),
    .Y(_02325_),
    .A1(_03472_),
    .A2(net457));
 sg13g2_buf_1 _19904_ (.A(net580),
    .X(_03855_));
 sg13g2_nand2_1 _19905_ (.Y(_03856_),
    .A(\top_ihp.oisc.regs[62][26] ),
    .B(net456));
 sg13g2_o21ai_1 _19906_ (.B1(_03856_),
    .Y(_02326_),
    .A1(_03474_),
    .A2(_03846_));
 sg13g2_nand2_1 _19907_ (.Y(_03857_),
    .A(\top_ihp.oisc.regs[62][27] ),
    .B(net456));
 sg13g2_o21ai_1 _19908_ (.B1(_03857_),
    .Y(_02327_),
    .A1(net224),
    .A2(net457));
 sg13g2_buf_1 _19909_ (.A(net580),
    .X(_03858_));
 sg13g2_nand2_1 _19910_ (.Y(_03859_),
    .A(\top_ihp.oisc.regs[62][28] ),
    .B(net456));
 sg13g2_o21ai_1 _19911_ (.B1(_03859_),
    .Y(_02328_),
    .A1(net223),
    .A2(net455));
 sg13g2_nand2_1 _19912_ (.Y(_03860_),
    .A(\top_ihp.oisc.regs[62][29] ),
    .B(net456));
 sg13g2_o21ai_1 _19913_ (.B1(_03860_),
    .Y(_02329_),
    .A1(net222),
    .A2(net455));
 sg13g2_nand2_1 _19914_ (.Y(_03861_),
    .A(\top_ihp.oisc.regs[62][2] ),
    .B(net456));
 sg13g2_o21ai_1 _19915_ (.B1(_03861_),
    .Y(_02330_),
    .A1(_03532_),
    .A2(net455));
 sg13g2_nand2_1 _19916_ (.Y(_03862_),
    .A(\top_ihp.oisc.regs[62][30] ),
    .B(_03855_));
 sg13g2_o21ai_1 _19917_ (.B1(_03862_),
    .Y(_02331_),
    .A1(net67),
    .A2(_03858_));
 sg13g2_nand2_1 _19918_ (.Y(_03863_),
    .A(\top_ihp.oisc.regs[62][31] ),
    .B(net456));
 sg13g2_o21ai_1 _19919_ (.B1(_03863_),
    .Y(_02332_),
    .A1(_10348_),
    .A2(net455));
 sg13g2_nand2_1 _19920_ (.Y(_03864_),
    .A(\top_ihp.oisc.regs[62][3] ),
    .B(net456));
 sg13g2_o21ai_1 _19921_ (.B1(_03864_),
    .Y(_02333_),
    .A1(net66),
    .A2(net455));
 sg13g2_nand2_1 _19922_ (.Y(_03865_),
    .A(\top_ihp.oisc.regs[62][4] ),
    .B(net456));
 sg13g2_o21ai_1 _19923_ (.B1(_03865_),
    .Y(_02334_),
    .A1(_03539_),
    .A2(net455));
 sg13g2_nand2_1 _19924_ (.Y(_03866_),
    .A(\top_ihp.oisc.regs[62][5] ),
    .B(_03855_));
 sg13g2_o21ai_1 _19925_ (.B1(_03866_),
    .Y(_02335_),
    .A1(net73),
    .A2(_03858_));
 sg13g2_nand2_1 _19926_ (.Y(_03867_),
    .A(\top_ihp.oisc.regs[62][6] ),
    .B(net580));
 sg13g2_o21ai_1 _19927_ (.B1(_03867_),
    .Y(_02336_),
    .A1(_03491_),
    .A2(net455));
 sg13g2_nand2_1 _19928_ (.Y(_03868_),
    .A(\top_ihp.oisc.regs[62][7] ),
    .B(net580));
 sg13g2_o21ai_1 _19929_ (.B1(_03868_),
    .Y(_02337_),
    .A1(_10483_),
    .A2(net455));
 sg13g2_nand2_1 _19930_ (.Y(_03869_),
    .A(\top_ihp.oisc.regs[62][8] ),
    .B(_03832_));
 sg13g2_o21ai_1 _19931_ (.B1(_03869_),
    .Y(_02338_),
    .A1(net221),
    .A2(_03834_));
 sg13g2_nand2_1 _19932_ (.Y(_03870_),
    .A(\top_ihp.oisc.regs[62][9] ),
    .B(net580));
 sg13g2_o21ai_1 _19933_ (.B1(_03870_),
    .Y(_02339_),
    .A1(net71),
    .A2(_03834_));
 sg13g2_nand2_1 _19934_ (.Y(_03871_),
    .A(_10619_),
    .B(_03313_));
 sg13g2_buf_1 _19935_ (.A(_03871_),
    .X(_03872_));
 sg13g2_buf_1 _19936_ (.A(net682),
    .X(_03873_));
 sg13g2_buf_1 _19937_ (.A(_03871_),
    .X(_03874_));
 sg13g2_nand2_1 _19938_ (.Y(_03875_),
    .A(\top_ihp.oisc.regs[63][0] ),
    .B(net681));
 sg13g2_o21ai_1 _19939_ (.B1(_03875_),
    .Y(_02340_),
    .A1(net70),
    .A2(net578));
 sg13g2_nand2_1 _19940_ (.Y(_03876_),
    .A(\top_ihp.oisc.regs[63][10] ),
    .B(net681));
 sg13g2_o21ai_1 _19941_ (.B1(_03876_),
    .Y(_02341_),
    .A1(_10623_),
    .A2(net578));
 sg13g2_nand2_1 _19942_ (.Y(_03877_),
    .A(\top_ihp.oisc.regs[63][11] ),
    .B(net681));
 sg13g2_o21ai_1 _19943_ (.B1(_03877_),
    .Y(_02342_),
    .A1(net69),
    .A2(net578));
 sg13g2_nand2_1 _19944_ (.Y(_03878_),
    .A(\top_ihp.oisc.regs[63][12] ),
    .B(net681));
 sg13g2_o21ai_1 _19945_ (.B1(_03878_),
    .Y(_02343_),
    .A1(net332),
    .A2(net578));
 sg13g2_nand2_1 _19946_ (.Y(_03879_),
    .A(\top_ihp.oisc.regs[63][13] ),
    .B(net681));
 sg13g2_o21ai_1 _19947_ (.B1(_03879_),
    .Y(_02344_),
    .A1(_10626_),
    .A2(net578));
 sg13g2_nand2_1 _19948_ (.Y(_03880_),
    .A(\top_ihp.oisc.regs[63][14] ),
    .B(net681));
 sg13g2_o21ai_1 _19949_ (.B1(_03880_),
    .Y(_02345_),
    .A1(_09977_),
    .A2(net578));
 sg13g2_nand2_1 _19950_ (.Y(_03881_),
    .A(\top_ihp.oisc.regs[63][15] ),
    .B(net681));
 sg13g2_o21ai_1 _19951_ (.B1(_03881_),
    .Y(_02346_),
    .A1(net220),
    .A2(net578));
 sg13g2_nand2_1 _19952_ (.Y(_03882_),
    .A(\top_ihp.oisc.regs[63][16] ),
    .B(net681));
 sg13g2_o21ai_1 _19953_ (.B1(_03882_),
    .Y(_02347_),
    .A1(_10628_),
    .A2(net578));
 sg13g2_buf_1 _19954_ (.A(net682),
    .X(_03883_));
 sg13g2_nand2_1 _19955_ (.Y(_03884_),
    .A(\top_ihp.oisc.regs[63][17] ),
    .B(net577));
 sg13g2_o21ai_1 _19956_ (.B1(_03884_),
    .Y(_02348_),
    .A1(_10629_),
    .A2(_03873_));
 sg13g2_nand2_1 _19957_ (.Y(_03885_),
    .A(\top_ihp.oisc.regs[63][18] ),
    .B(net577));
 sg13g2_o21ai_1 _19958_ (.B1(_03885_),
    .Y(_02349_),
    .A1(_10630_),
    .A2(_03873_));
 sg13g2_buf_1 _19959_ (.A(net682),
    .X(_03886_));
 sg13g2_nand2_1 _19960_ (.Y(_03887_),
    .A(\top_ihp.oisc.regs[63][19] ),
    .B(net577));
 sg13g2_o21ai_1 _19961_ (.B1(_03887_),
    .Y(_02350_),
    .A1(_10631_),
    .A2(net576));
 sg13g2_nand2_1 _19962_ (.Y(_03888_),
    .A(\top_ihp.oisc.regs[63][1] ),
    .B(net577));
 sg13g2_o21ai_1 _19963_ (.B1(_03888_),
    .Y(_02351_),
    .A1(_10127_),
    .A2(net576));
 sg13g2_nand2_1 _19964_ (.Y(_03889_),
    .A(\top_ihp.oisc.regs[63][20] ),
    .B(_03883_));
 sg13g2_o21ai_1 _19965_ (.B1(_03889_),
    .Y(_02352_),
    .A1(net607),
    .A2(net576));
 sg13g2_nand2_1 _19966_ (.Y(_03890_),
    .A(\top_ihp.oisc.regs[63][21] ),
    .B(net577));
 sg13g2_o21ai_1 _19967_ (.B1(_03890_),
    .Y(_02353_),
    .A1(net310),
    .A2(net576));
 sg13g2_nand2_1 _19968_ (.Y(_03891_),
    .A(\top_ihp.oisc.regs[63][22] ),
    .B(net577));
 sg13g2_o21ai_1 _19969_ (.B1(_03891_),
    .Y(_02354_),
    .A1(net322),
    .A2(net576));
 sg13g2_nand2_1 _19970_ (.Y(_03892_),
    .A(\top_ihp.oisc.regs[63][23] ),
    .B(net577));
 sg13g2_o21ai_1 _19971_ (.B1(_03892_),
    .Y(_02355_),
    .A1(_10203_),
    .A2(net576));
 sg13g2_nand2_1 _19972_ (.Y(_03893_),
    .A(\top_ihp.oisc.regs[63][24] ),
    .B(_03883_));
 sg13g2_o21ai_1 _19973_ (.B1(_03893_),
    .Y(_02356_),
    .A1(_10636_),
    .A2(_03886_));
 sg13g2_nand2_1 _19974_ (.Y(_03894_),
    .A(\top_ihp.oisc.regs[63][25] ),
    .B(net577));
 sg13g2_o21ai_1 _19975_ (.B1(_03894_),
    .Y(_02357_),
    .A1(net319),
    .A2(net576));
 sg13g2_buf_1 _19976_ (.A(net682),
    .X(_03895_));
 sg13g2_nand2_1 _19977_ (.Y(_03896_),
    .A(\top_ihp.oisc.regs[63][26] ),
    .B(net575));
 sg13g2_o21ai_1 _19978_ (.B1(_03896_),
    .Y(_02358_),
    .A1(_10638_),
    .A2(_03886_));
 sg13g2_nand2_1 _19979_ (.Y(_03897_),
    .A(\top_ihp.oisc.regs[63][27] ),
    .B(net575));
 sg13g2_o21ai_1 _19980_ (.B1(_03897_),
    .Y(_02359_),
    .A1(_10639_),
    .A2(net576));
 sg13g2_buf_1 _19981_ (.A(net682),
    .X(_03898_));
 sg13g2_nand2_1 _19982_ (.Y(_03899_),
    .A(\top_ihp.oisc.regs[63][28] ),
    .B(net575));
 sg13g2_o21ai_1 _19983_ (.B1(_03899_),
    .Y(_02360_),
    .A1(_10640_),
    .A2(net574));
 sg13g2_nand2_1 _19984_ (.Y(_03900_),
    .A(\top_ihp.oisc.regs[63][29] ),
    .B(net575));
 sg13g2_o21ai_1 _19985_ (.B1(_03900_),
    .Y(_02361_),
    .A1(net307),
    .A2(net574));
 sg13g2_nand2_1 _19986_ (.Y(_03901_),
    .A(\top_ihp.oisc.regs[63][2] ),
    .B(net575));
 sg13g2_o21ai_1 _19987_ (.B1(_03901_),
    .Y(_02362_),
    .A1(net68),
    .A2(_03898_));
 sg13g2_nand2_1 _19988_ (.Y(_03902_),
    .A(\top_ihp.oisc.regs[63][30] ),
    .B(net575));
 sg13g2_o21ai_1 _19989_ (.B1(_03902_),
    .Y(_02363_),
    .A1(net67),
    .A2(net574));
 sg13g2_nand2_1 _19990_ (.Y(_03903_),
    .A(\top_ihp.oisc.regs[63][31] ),
    .B(_03895_));
 sg13g2_o21ai_1 _19991_ (.B1(_03903_),
    .Y(_02364_),
    .A1(_10644_),
    .A2(net574));
 sg13g2_nand2_1 _19992_ (.Y(_03904_),
    .A(\top_ihp.oisc.regs[63][3] ),
    .B(net575));
 sg13g2_o21ai_1 _19993_ (.B1(_03904_),
    .Y(_02365_),
    .A1(net66),
    .A2(net574));
 sg13g2_nand2_1 _19994_ (.Y(_03905_),
    .A(\top_ihp.oisc.regs[63][4] ),
    .B(_03895_));
 sg13g2_o21ai_1 _19995_ (.B1(_03905_),
    .Y(_02366_),
    .A1(net65),
    .A2(net574));
 sg13g2_nand2_1 _19996_ (.Y(_03906_),
    .A(\top_ihp.oisc.regs[63][5] ),
    .B(net575));
 sg13g2_o21ai_1 _19997_ (.B1(_03906_),
    .Y(_02367_),
    .A1(net123),
    .A2(_03898_));
 sg13g2_nand2_1 _19998_ (.Y(_03907_),
    .A(\top_ihp.oisc.regs[63][6] ),
    .B(net682));
 sg13g2_o21ai_1 _19999_ (.B1(_03907_),
    .Y(_02368_),
    .A1(net122),
    .A2(net574));
 sg13g2_nand2_1 _20000_ (.Y(_03908_),
    .A(\top_ihp.oisc.regs[63][7] ),
    .B(net682));
 sg13g2_o21ai_1 _20001_ (.B1(_03908_),
    .Y(_02369_),
    .A1(net470),
    .A2(net574));
 sg13g2_nand2_1 _20002_ (.Y(_03909_),
    .A(\top_ihp.oisc.regs[63][8] ),
    .B(_03872_));
 sg13g2_o21ai_1 _20003_ (.B1(_03909_),
    .Y(_02370_),
    .A1(net305),
    .A2(_03874_));
 sg13g2_nand2_1 _20004_ (.Y(_03910_),
    .A(\top_ihp.oisc.regs[63][9] ),
    .B(net682));
 sg13g2_o21ai_1 _20005_ (.B1(_03910_),
    .Y(_02371_),
    .A1(net121),
    .A2(_03874_));
 sg13g2_nand2_1 _20006_ (.Y(_03911_),
    .A(_10524_),
    .B(net762));
 sg13g2_buf_1 _20007_ (.A(_03911_),
    .X(_03912_));
 sg13g2_buf_1 _20008_ (.A(net573),
    .X(_03913_));
 sg13g2_buf_1 _20009_ (.A(_03911_),
    .X(_03914_));
 sg13g2_nand2_1 _20010_ (.Y(_03915_),
    .A(\top_ihp.oisc.regs[6][0] ),
    .B(net572));
 sg13g2_o21ai_1 _20011_ (.B1(_03915_),
    .Y(_02372_),
    .A1(_09697_),
    .A2(_03913_));
 sg13g2_nand2_1 _20012_ (.Y(_03916_),
    .A(\top_ihp.oisc.regs[6][10] ),
    .B(net572));
 sg13g2_o21ai_1 _20013_ (.B1(_03916_),
    .Y(_02373_),
    .A1(net128),
    .A2(net454));
 sg13g2_nand2_1 _20014_ (.Y(_03917_),
    .A(\top_ihp.oisc.regs[6][11] ),
    .B(net572));
 sg13g2_o21ai_1 _20015_ (.B1(_03917_),
    .Y(_02374_),
    .A1(net127),
    .A2(net454));
 sg13g2_nand2_1 _20016_ (.Y(_03918_),
    .A(\top_ihp.oisc.regs[6][12] ),
    .B(net572));
 sg13g2_o21ai_1 _20017_ (.B1(_03918_),
    .Y(_02375_),
    .A1(net332),
    .A2(net454));
 sg13g2_nand2_1 _20018_ (.Y(_03919_),
    .A(\top_ihp.oisc.regs[6][13] ),
    .B(net572));
 sg13g2_o21ai_1 _20019_ (.B1(_03919_),
    .Y(_02376_),
    .A1(net314),
    .A2(net454));
 sg13g2_nand2_1 _20020_ (.Y(_03920_),
    .A(\top_ihp.oisc.regs[6][14] ),
    .B(net572));
 sg13g2_o21ai_1 _20021_ (.B1(_03920_),
    .Y(_02377_),
    .A1(net330),
    .A2(net454));
 sg13g2_nand2_1 _20022_ (.Y(_03921_),
    .A(\top_ihp.oisc.regs[6][15] ),
    .B(net572));
 sg13g2_o21ai_1 _20023_ (.B1(_03921_),
    .Y(_02378_),
    .A1(net329),
    .A2(net454));
 sg13g2_nand2_1 _20024_ (.Y(_03922_),
    .A(\top_ihp.oisc.regs[6][16] ),
    .B(net572));
 sg13g2_o21ai_1 _20025_ (.B1(_03922_),
    .Y(_02379_),
    .A1(net126),
    .A2(_03913_));
 sg13g2_buf_1 _20026_ (.A(net573),
    .X(_03923_));
 sg13g2_nand2_1 _20027_ (.Y(_03924_),
    .A(\top_ihp.oisc.regs[6][17] ),
    .B(_03923_));
 sg13g2_o21ai_1 _20028_ (.B1(_03924_),
    .Y(_02380_),
    .A1(net313),
    .A2(net454));
 sg13g2_nand2_1 _20029_ (.Y(_03925_),
    .A(\top_ihp.oisc.regs[6][18] ),
    .B(net453));
 sg13g2_o21ai_1 _20030_ (.B1(_03925_),
    .Y(_02381_),
    .A1(net312),
    .A2(net454));
 sg13g2_buf_1 _20031_ (.A(net573),
    .X(_03926_));
 sg13g2_nand2_1 _20032_ (.Y(_03927_),
    .A(\top_ihp.oisc.regs[6][19] ),
    .B(net453));
 sg13g2_o21ai_1 _20033_ (.B1(_03927_),
    .Y(_02382_),
    .A1(net311),
    .A2(net452));
 sg13g2_nand2_1 _20034_ (.Y(_03928_),
    .A(\top_ihp.oisc.regs[6][1] ),
    .B(net453));
 sg13g2_o21ai_1 _20035_ (.B1(_03928_),
    .Y(_02383_),
    .A1(net325),
    .A2(net452));
 sg13g2_nand2_1 _20036_ (.Y(_03929_),
    .A(\top_ihp.oisc.regs[6][20] ),
    .B(net453));
 sg13g2_o21ai_1 _20037_ (.B1(_03929_),
    .Y(_02384_),
    .A1(_10152_),
    .A2(net452));
 sg13g2_nand2_1 _20038_ (.Y(_03930_),
    .A(\top_ihp.oisc.regs[6][21] ),
    .B(net453));
 sg13g2_o21ai_1 _20039_ (.B1(_03930_),
    .Y(_02385_),
    .A1(net310),
    .A2(net452));
 sg13g2_nand2_1 _20040_ (.Y(_03931_),
    .A(\top_ihp.oisc.regs[6][22] ),
    .B(_03923_));
 sg13g2_o21ai_1 _20041_ (.B1(_03931_),
    .Y(_02386_),
    .A1(net322),
    .A2(_03926_));
 sg13g2_nand2_1 _20042_ (.Y(_03932_),
    .A(\top_ihp.oisc.regs[6][23] ),
    .B(net453));
 sg13g2_o21ai_1 _20043_ (.B1(_03932_),
    .Y(_02387_),
    .A1(net528),
    .A2(_03926_));
 sg13g2_nand2_1 _20044_ (.Y(_03933_),
    .A(\top_ihp.oisc.regs[6][24] ),
    .B(net453));
 sg13g2_o21ai_1 _20045_ (.B1(_03933_),
    .Y(_02388_),
    .A1(net309),
    .A2(net452));
 sg13g2_nand2_1 _20046_ (.Y(_03934_),
    .A(\top_ihp.oisc.regs[6][25] ),
    .B(net453));
 sg13g2_o21ai_1 _20047_ (.B1(_03934_),
    .Y(_02389_),
    .A1(net319),
    .A2(net452));
 sg13g2_buf_1 _20048_ (.A(net573),
    .X(_03935_));
 sg13g2_nand2_1 _20049_ (.Y(_03936_),
    .A(\top_ihp.oisc.regs[6][26] ),
    .B(net451));
 sg13g2_o21ai_1 _20050_ (.B1(_03936_),
    .Y(_02390_),
    .A1(net125),
    .A2(net452));
 sg13g2_nand2_1 _20051_ (.Y(_03937_),
    .A(\top_ihp.oisc.regs[6][27] ),
    .B(net451));
 sg13g2_o21ai_1 _20052_ (.B1(_03937_),
    .Y(_02391_),
    .A1(net308),
    .A2(net452));
 sg13g2_buf_1 _20053_ (.A(net573),
    .X(_03938_));
 sg13g2_nand2_1 _20054_ (.Y(_03939_),
    .A(\top_ihp.oisc.regs[6][28] ),
    .B(_03935_));
 sg13g2_o21ai_1 _20055_ (.B1(_03939_),
    .Y(_02392_),
    .A1(net515),
    .A2(net450));
 sg13g2_nand2_1 _20056_ (.Y(_03940_),
    .A(\top_ihp.oisc.regs[6][29] ),
    .B(_03935_));
 sg13g2_o21ai_1 _20057_ (.B1(_03940_),
    .Y(_02393_),
    .A1(net307),
    .A2(_03938_));
 sg13g2_nand2_1 _20058_ (.Y(_03941_),
    .A(\top_ihp.oisc.regs[6][2] ),
    .B(net451));
 sg13g2_o21ai_1 _20059_ (.B1(_03941_),
    .Y(_02394_),
    .A1(net131),
    .A2(_03938_));
 sg13g2_nand2_1 _20060_ (.Y(_03942_),
    .A(\top_ihp.oisc.regs[6][30] ),
    .B(net451));
 sg13g2_o21ai_1 _20061_ (.B1(_03942_),
    .Y(_02395_),
    .A1(net124),
    .A2(net450));
 sg13g2_nand2_1 _20062_ (.Y(_03943_),
    .A(\top_ihp.oisc.regs[6][31] ),
    .B(net451));
 sg13g2_o21ai_1 _20063_ (.B1(_03943_),
    .Y(_02396_),
    .A1(_10348_),
    .A2(net450));
 sg13g2_nand2_1 _20064_ (.Y(_03944_),
    .A(\top_ihp.oisc.regs[6][3] ),
    .B(net451));
 sg13g2_o21ai_1 _20065_ (.B1(_03944_),
    .Y(_02397_),
    .A1(_10608_),
    .A2(net450));
 sg13g2_nand2_1 _20066_ (.Y(_03945_),
    .A(\top_ihp.oisc.regs[6][4] ),
    .B(net451));
 sg13g2_o21ai_1 _20067_ (.B1(_03945_),
    .Y(_02398_),
    .A1(net129),
    .A2(net450));
 sg13g2_nand2_1 _20068_ (.Y(_03946_),
    .A(\top_ihp.oisc.regs[6][5] ),
    .B(net451));
 sg13g2_o21ai_1 _20069_ (.B1(_03946_),
    .Y(_02399_),
    .A1(_10645_),
    .A2(net450));
 sg13g2_nand2_1 _20070_ (.Y(_03947_),
    .A(\top_ihp.oisc.regs[6][6] ),
    .B(net573));
 sg13g2_o21ai_1 _20071_ (.B1(_03947_),
    .Y(_02400_),
    .A1(net122),
    .A2(net450));
 sg13g2_nand2_1 _20072_ (.Y(_03948_),
    .A(\top_ihp.oisc.regs[6][7] ),
    .B(net573));
 sg13g2_o21ai_1 _20073_ (.B1(_03948_),
    .Y(_02401_),
    .A1(_10483_),
    .A2(net450));
 sg13g2_nand2_1 _20074_ (.Y(_03949_),
    .A(\top_ihp.oisc.regs[6][8] ),
    .B(_03912_));
 sg13g2_o21ai_1 _20075_ (.B1(_03949_),
    .Y(_02402_),
    .A1(net305),
    .A2(_03914_));
 sg13g2_nand2_1 _20076_ (.Y(_03950_),
    .A(\top_ihp.oisc.regs[6][9] ),
    .B(net573));
 sg13g2_o21ai_1 _20077_ (.B1(_03950_),
    .Y(_02403_),
    .A1(net121),
    .A2(_03914_));
 sg13g2_nand2_1 _20078_ (.Y(_03951_),
    .A(_10572_),
    .B(net762));
 sg13g2_buf_1 _20079_ (.A(_03951_),
    .X(_03952_));
 sg13g2_buf_1 _20080_ (.A(net680),
    .X(_03953_));
 sg13g2_buf_1 _20081_ (.A(_03951_),
    .X(_03954_));
 sg13g2_nand2_1 _20082_ (.Y(_03955_),
    .A(\top_ihp.oisc.regs[7][0] ),
    .B(net679));
 sg13g2_o21ai_1 _20083_ (.B1(_03955_),
    .Y(_02404_),
    .A1(net156),
    .A2(net571));
 sg13g2_nand2_1 _20084_ (.Y(_03956_),
    .A(\top_ihp.oisc.regs[7][10] ),
    .B(net679));
 sg13g2_o21ai_1 _20085_ (.B1(_03956_),
    .Y(_02405_),
    .A1(net128),
    .A2(net571));
 sg13g2_nand2_1 _20086_ (.Y(_03957_),
    .A(\top_ihp.oisc.regs[7][11] ),
    .B(net679));
 sg13g2_o21ai_1 _20087_ (.B1(_03957_),
    .Y(_02406_),
    .A1(net127),
    .A2(net571));
 sg13g2_nand2_1 _20088_ (.Y(_03958_),
    .A(\top_ihp.oisc.regs[7][12] ),
    .B(net679));
 sg13g2_o21ai_1 _20089_ (.B1(_03958_),
    .Y(_02407_),
    .A1(net332),
    .A2(net571));
 sg13g2_nand2_1 _20090_ (.Y(_03959_),
    .A(\top_ihp.oisc.regs[7][13] ),
    .B(net679));
 sg13g2_o21ai_1 _20091_ (.B1(_03959_),
    .Y(_02408_),
    .A1(net314),
    .A2(net571));
 sg13g2_nand2_1 _20092_ (.Y(_03960_),
    .A(\top_ihp.oisc.regs[7][14] ),
    .B(net679));
 sg13g2_o21ai_1 _20093_ (.B1(_03960_),
    .Y(_02409_),
    .A1(net330),
    .A2(net571));
 sg13g2_nand2_1 _20094_ (.Y(_03961_),
    .A(\top_ihp.oisc.regs[7][15] ),
    .B(net679));
 sg13g2_o21ai_1 _20095_ (.B1(_03961_),
    .Y(_02410_),
    .A1(net329),
    .A2(_03953_));
 sg13g2_nand2_1 _20096_ (.Y(_03962_),
    .A(\top_ihp.oisc.regs[7][16] ),
    .B(net679));
 sg13g2_o21ai_1 _20097_ (.B1(_03962_),
    .Y(_02411_),
    .A1(net126),
    .A2(_03953_));
 sg13g2_buf_1 _20098_ (.A(net680),
    .X(_03963_));
 sg13g2_nand2_1 _20099_ (.Y(_03964_),
    .A(\top_ihp.oisc.regs[7][17] ),
    .B(net570));
 sg13g2_o21ai_1 _20100_ (.B1(_03964_),
    .Y(_02412_),
    .A1(net313),
    .A2(net571));
 sg13g2_nand2_1 _20101_ (.Y(_03965_),
    .A(\top_ihp.oisc.regs[7][18] ),
    .B(net570));
 sg13g2_o21ai_1 _20102_ (.B1(_03965_),
    .Y(_02413_),
    .A1(net312),
    .A2(net571));
 sg13g2_buf_1 _20103_ (.A(net680),
    .X(_03966_));
 sg13g2_nand2_1 _20104_ (.Y(_03967_),
    .A(\top_ihp.oisc.regs[7][19] ),
    .B(net570));
 sg13g2_o21ai_1 _20105_ (.B1(_03967_),
    .Y(_02414_),
    .A1(net311),
    .A2(net569));
 sg13g2_nand2_1 _20106_ (.Y(_03968_),
    .A(\top_ihp.oisc.regs[7][1] ),
    .B(_03963_));
 sg13g2_o21ai_1 _20107_ (.B1(_03968_),
    .Y(_02415_),
    .A1(net325),
    .A2(_03966_));
 sg13g2_nand2_1 _20108_ (.Y(_03969_),
    .A(\top_ihp.oisc.regs[7][20] ),
    .B(net570));
 sg13g2_o21ai_1 _20109_ (.B1(_03969_),
    .Y(_02416_),
    .A1(net607),
    .A2(net569));
 sg13g2_nand2_1 _20110_ (.Y(_03970_),
    .A(\top_ihp.oisc.regs[7][21] ),
    .B(net570));
 sg13g2_o21ai_1 _20111_ (.B1(_03970_),
    .Y(_02417_),
    .A1(net310),
    .A2(net569));
 sg13g2_nand2_1 _20112_ (.Y(_03971_),
    .A(\top_ihp.oisc.regs[7][22] ),
    .B(net570));
 sg13g2_o21ai_1 _20113_ (.B1(_03971_),
    .Y(_02418_),
    .A1(net322),
    .A2(net569));
 sg13g2_nand2_1 _20114_ (.Y(_03972_),
    .A(\top_ihp.oisc.regs[7][23] ),
    .B(_03963_));
 sg13g2_o21ai_1 _20115_ (.B1(_03972_),
    .Y(_02419_),
    .A1(net528),
    .A2(_03966_));
 sg13g2_nand2_1 _20116_ (.Y(_03973_),
    .A(\top_ihp.oisc.regs[7][24] ),
    .B(net570));
 sg13g2_o21ai_1 _20117_ (.B1(_03973_),
    .Y(_02420_),
    .A1(net309),
    .A2(net569));
 sg13g2_nand2_1 _20118_ (.Y(_03974_),
    .A(\top_ihp.oisc.regs[7][25] ),
    .B(net570));
 sg13g2_o21ai_1 _20119_ (.B1(_03974_),
    .Y(_02421_),
    .A1(net319),
    .A2(net569));
 sg13g2_buf_1 _20120_ (.A(net680),
    .X(_03975_));
 sg13g2_nand2_1 _20121_ (.Y(_03976_),
    .A(\top_ihp.oisc.regs[7][26] ),
    .B(net568));
 sg13g2_o21ai_1 _20122_ (.B1(_03976_),
    .Y(_02422_),
    .A1(net125),
    .A2(net569));
 sg13g2_nand2_1 _20123_ (.Y(_03977_),
    .A(\top_ihp.oisc.regs[7][27] ),
    .B(net568));
 sg13g2_o21ai_1 _20124_ (.B1(_03977_),
    .Y(_02423_),
    .A1(net308),
    .A2(net569));
 sg13g2_buf_1 _20125_ (.A(net680),
    .X(_03978_));
 sg13g2_nand2_1 _20126_ (.Y(_03979_),
    .A(\top_ihp.oisc.regs[7][28] ),
    .B(_03975_));
 sg13g2_o21ai_1 _20127_ (.B1(_03979_),
    .Y(_02424_),
    .A1(net515),
    .A2(_03978_));
 sg13g2_nand2_1 _20128_ (.Y(_03980_),
    .A(\top_ihp.oisc.regs[7][29] ),
    .B(_03975_));
 sg13g2_o21ai_1 _20129_ (.B1(_03980_),
    .Y(_02425_),
    .A1(net307),
    .A2(_03978_));
 sg13g2_nand2_1 _20130_ (.Y(_03981_),
    .A(\top_ihp.oisc.regs[7][2] ),
    .B(net568));
 sg13g2_o21ai_1 _20131_ (.B1(_03981_),
    .Y(_02426_),
    .A1(net131),
    .A2(net567));
 sg13g2_nand2_1 _20132_ (.Y(_03982_),
    .A(\top_ihp.oisc.regs[7][30] ),
    .B(net568));
 sg13g2_o21ai_1 _20133_ (.B1(_03982_),
    .Y(_02427_),
    .A1(net124),
    .A2(net567));
 sg13g2_nand2_1 _20134_ (.Y(_03983_),
    .A(\top_ihp.oisc.regs[7][31] ),
    .B(net568));
 sg13g2_o21ai_1 _20135_ (.B1(_03983_),
    .Y(_02428_),
    .A1(net306),
    .A2(net567));
 sg13g2_nand2_1 _20136_ (.Y(_03984_),
    .A(\top_ihp.oisc.regs[7][3] ),
    .B(net568));
 sg13g2_o21ai_1 _20137_ (.B1(_03984_),
    .Y(_02429_),
    .A1(net130),
    .A2(net567));
 sg13g2_nand2_1 _20138_ (.Y(_03985_),
    .A(\top_ihp.oisc.regs[7][4] ),
    .B(net568));
 sg13g2_o21ai_1 _20139_ (.B1(_03985_),
    .Y(_02430_),
    .A1(_10609_),
    .A2(net567));
 sg13g2_nand2_1 _20140_ (.Y(_03986_),
    .A(\top_ihp.oisc.regs[7][5] ),
    .B(net568));
 sg13g2_o21ai_1 _20141_ (.B1(_03986_),
    .Y(_02431_),
    .A1(net123),
    .A2(net567));
 sg13g2_nand2_1 _20142_ (.Y(_03987_),
    .A(\top_ihp.oisc.regs[7][6] ),
    .B(net680));
 sg13g2_o21ai_1 _20143_ (.B1(_03987_),
    .Y(_02432_),
    .A1(net122),
    .A2(net567));
 sg13g2_nand2_1 _20144_ (.Y(_03988_),
    .A(\top_ihp.oisc.regs[7][7] ),
    .B(net680));
 sg13g2_o21ai_1 _20145_ (.B1(_03988_),
    .Y(_02433_),
    .A1(net470),
    .A2(net567));
 sg13g2_nand2_1 _20146_ (.Y(_03989_),
    .A(\top_ihp.oisc.regs[7][8] ),
    .B(_03952_));
 sg13g2_o21ai_1 _20147_ (.B1(_03989_),
    .Y(_02434_),
    .A1(net305),
    .A2(_03954_));
 sg13g2_nand2_1 _20148_ (.Y(_03990_),
    .A(\top_ihp.oisc.regs[7][9] ),
    .B(net680));
 sg13g2_o21ai_1 _20149_ (.B1(_03990_),
    .Y(_02435_),
    .A1(net121),
    .A2(_03954_));
 sg13g2_nand2_1 _20150_ (.Y(_03991_),
    .A(_09754_),
    .B(net764));
 sg13g2_buf_1 _20151_ (.A(_03991_),
    .X(_03992_));
 sg13g2_buf_1 _20152_ (.A(net566),
    .X(_03993_));
 sg13g2_buf_1 _20153_ (.A(_03991_),
    .X(_03994_));
 sg13g2_nand2_1 _20154_ (.Y(_03995_),
    .A(\top_ihp.oisc.regs[8][0] ),
    .B(net565));
 sg13g2_o21ai_1 _20155_ (.B1(_03995_),
    .Y(_02436_),
    .A1(net156),
    .A2(net449));
 sg13g2_nand2_1 _20156_ (.Y(_03996_),
    .A(\top_ihp.oisc.regs[8][10] ),
    .B(net565));
 sg13g2_o21ai_1 _20157_ (.B1(_03996_),
    .Y(_02437_),
    .A1(net128),
    .A2(net449));
 sg13g2_nand2_1 _20158_ (.Y(_03997_),
    .A(\top_ihp.oisc.regs[8][11] ),
    .B(net565));
 sg13g2_o21ai_1 _20159_ (.B1(_03997_),
    .Y(_02438_),
    .A1(_10624_),
    .A2(net449));
 sg13g2_nand2_1 _20160_ (.Y(_03998_),
    .A(\top_ihp.oisc.regs[8][12] ),
    .B(net565));
 sg13g2_o21ai_1 _20161_ (.B1(_03998_),
    .Y(_02439_),
    .A1(net332),
    .A2(net449));
 sg13g2_nand2_1 _20162_ (.Y(_03999_),
    .A(\top_ihp.oisc.regs[8][13] ),
    .B(net565));
 sg13g2_o21ai_1 _20163_ (.B1(_03999_),
    .Y(_02440_),
    .A1(net314),
    .A2(net449));
 sg13g2_nand2_1 _20164_ (.Y(_04000_),
    .A(\top_ihp.oisc.regs[8][14] ),
    .B(net565));
 sg13g2_o21ai_1 _20165_ (.B1(_04000_),
    .Y(_02441_),
    .A1(net330),
    .A2(_03993_));
 sg13g2_nand2_1 _20166_ (.Y(_04001_),
    .A(\top_ihp.oisc.regs[8][15] ),
    .B(net565));
 sg13g2_o21ai_1 _20167_ (.B1(_04001_),
    .Y(_02442_),
    .A1(net329),
    .A2(net449));
 sg13g2_nand2_1 _20168_ (.Y(_04002_),
    .A(\top_ihp.oisc.regs[8][16] ),
    .B(net565));
 sg13g2_o21ai_1 _20169_ (.B1(_04002_),
    .Y(_02443_),
    .A1(net126),
    .A2(_03993_));
 sg13g2_buf_1 _20170_ (.A(net566),
    .X(_04003_));
 sg13g2_nand2_1 _20171_ (.Y(_04004_),
    .A(\top_ihp.oisc.regs[8][17] ),
    .B(net448));
 sg13g2_o21ai_1 _20172_ (.B1(_04004_),
    .Y(_02444_),
    .A1(net313),
    .A2(net449));
 sg13g2_nand2_1 _20173_ (.Y(_04005_),
    .A(\top_ihp.oisc.regs[8][18] ),
    .B(net448));
 sg13g2_o21ai_1 _20174_ (.B1(_04005_),
    .Y(_02445_),
    .A1(net312),
    .A2(net449));
 sg13g2_buf_1 _20175_ (.A(net566),
    .X(_04006_));
 sg13g2_nand2_1 _20176_ (.Y(_04007_),
    .A(\top_ihp.oisc.regs[8][19] ),
    .B(net448));
 sg13g2_o21ai_1 _20177_ (.B1(_04007_),
    .Y(_02446_),
    .A1(net311),
    .A2(net447));
 sg13g2_nand2_1 _20178_ (.Y(_04008_),
    .A(\top_ihp.oisc.regs[8][1] ),
    .B(net448));
 sg13g2_o21ai_1 _20179_ (.B1(_04008_),
    .Y(_02447_),
    .A1(net325),
    .A2(net447));
 sg13g2_nand2_1 _20180_ (.Y(_04009_),
    .A(\top_ihp.oisc.regs[8][20] ),
    .B(net448));
 sg13g2_o21ai_1 _20181_ (.B1(_04009_),
    .Y(_02448_),
    .A1(_10152_),
    .A2(_04006_));
 sg13g2_nand2_1 _20182_ (.Y(_04010_),
    .A(\top_ihp.oisc.regs[8][21] ),
    .B(net448));
 sg13g2_o21ai_1 _20183_ (.B1(_04010_),
    .Y(_02449_),
    .A1(net310),
    .A2(net447));
 sg13g2_nand2_1 _20184_ (.Y(_04011_),
    .A(\top_ihp.oisc.regs[8][22] ),
    .B(_04003_));
 sg13g2_o21ai_1 _20185_ (.B1(_04011_),
    .Y(_02450_),
    .A1(net322),
    .A2(_04006_));
 sg13g2_nand2_1 _20186_ (.Y(_04012_),
    .A(\top_ihp.oisc.regs[8][23] ),
    .B(net448));
 sg13g2_o21ai_1 _20187_ (.B1(_04012_),
    .Y(_02451_),
    .A1(net528),
    .A2(net447));
 sg13g2_nand2_1 _20188_ (.Y(_04013_),
    .A(\top_ihp.oisc.regs[8][24] ),
    .B(_04003_));
 sg13g2_o21ai_1 _20189_ (.B1(_04013_),
    .Y(_02452_),
    .A1(net309),
    .A2(net447));
 sg13g2_nand2_1 _20190_ (.Y(_04014_),
    .A(\top_ihp.oisc.regs[8][25] ),
    .B(net448));
 sg13g2_o21ai_1 _20191_ (.B1(_04014_),
    .Y(_02453_),
    .A1(net319),
    .A2(net447));
 sg13g2_buf_1 _20192_ (.A(net566),
    .X(_04015_));
 sg13g2_nand2_1 _20193_ (.Y(_04016_),
    .A(\top_ihp.oisc.regs[8][26] ),
    .B(_04015_));
 sg13g2_o21ai_1 _20194_ (.B1(_04016_),
    .Y(_02454_),
    .A1(net125),
    .A2(net447));
 sg13g2_nand2_1 _20195_ (.Y(_04017_),
    .A(\top_ihp.oisc.regs[8][27] ),
    .B(net446));
 sg13g2_o21ai_1 _20196_ (.B1(_04017_),
    .Y(_02455_),
    .A1(net308),
    .A2(net447));
 sg13g2_buf_1 _20197_ (.A(net566),
    .X(_04018_));
 sg13g2_nand2_1 _20198_ (.Y(_04019_),
    .A(\top_ihp.oisc.regs[8][28] ),
    .B(net446));
 sg13g2_o21ai_1 _20199_ (.B1(_04019_),
    .Y(_02456_),
    .A1(net515),
    .A2(net445));
 sg13g2_nand2_1 _20200_ (.Y(_04020_),
    .A(\top_ihp.oisc.regs[8][29] ),
    .B(_04015_));
 sg13g2_o21ai_1 _20201_ (.B1(_04020_),
    .Y(_02457_),
    .A1(net307),
    .A2(net445));
 sg13g2_nand2_1 _20202_ (.Y(_04021_),
    .A(\top_ihp.oisc.regs[8][2] ),
    .B(net446));
 sg13g2_o21ai_1 _20203_ (.B1(_04021_),
    .Y(_02458_),
    .A1(net131),
    .A2(_04018_));
 sg13g2_nand2_1 _20204_ (.Y(_04022_),
    .A(\top_ihp.oisc.regs[8][30] ),
    .B(net446));
 sg13g2_o21ai_1 _20205_ (.B1(_04022_),
    .Y(_02459_),
    .A1(net124),
    .A2(net445));
 sg13g2_nand2_1 _20206_ (.Y(_04023_),
    .A(\top_ihp.oisc.regs[8][31] ),
    .B(net446));
 sg13g2_o21ai_1 _20207_ (.B1(_04023_),
    .Y(_02460_),
    .A1(_10348_),
    .A2(net445));
 sg13g2_nand2_1 _20208_ (.Y(_04024_),
    .A(\top_ihp.oisc.regs[8][3] ),
    .B(net446));
 sg13g2_o21ai_1 _20209_ (.B1(_04024_),
    .Y(_02461_),
    .A1(net130),
    .A2(net445));
 sg13g2_nand2_1 _20210_ (.Y(_04025_),
    .A(\top_ihp.oisc.regs[8][4] ),
    .B(net446));
 sg13g2_o21ai_1 _20211_ (.B1(_04025_),
    .Y(_02462_),
    .A1(net129),
    .A2(net445));
 sg13g2_nand2_1 _20212_ (.Y(_04026_),
    .A(\top_ihp.oisc.regs[8][5] ),
    .B(net446));
 sg13g2_o21ai_1 _20213_ (.B1(_04026_),
    .Y(_02463_),
    .A1(net123),
    .A2(net445));
 sg13g2_nand2_1 _20214_ (.Y(_04027_),
    .A(\top_ihp.oisc.regs[8][6] ),
    .B(net566));
 sg13g2_o21ai_1 _20215_ (.B1(_04027_),
    .Y(_02464_),
    .A1(net122),
    .A2(net445));
 sg13g2_nand2_1 _20216_ (.Y(_04028_),
    .A(\top_ihp.oisc.regs[8][7] ),
    .B(net566));
 sg13g2_o21ai_1 _20217_ (.B1(_04028_),
    .Y(_02465_),
    .A1(_10483_),
    .A2(_04018_));
 sg13g2_nand2_1 _20218_ (.Y(_04029_),
    .A(\top_ihp.oisc.regs[8][8] ),
    .B(_03992_));
 sg13g2_o21ai_1 _20219_ (.B1(_04029_),
    .Y(_02466_),
    .A1(_10647_),
    .A2(_03994_));
 sg13g2_nand2_1 _20220_ (.Y(_04030_),
    .A(\top_ihp.oisc.regs[8][9] ),
    .B(net566));
 sg13g2_o21ai_1 _20221_ (.B1(_04030_),
    .Y(_02467_),
    .A1(net121),
    .A2(_03994_));
 sg13g2_nand2_1 _20222_ (.Y(_04031_),
    .A(net764),
    .B(_10651_));
 sg13g2_buf_1 _20223_ (.A(_04031_),
    .X(_04032_));
 sg13g2_buf_1 _20224_ (.A(net731),
    .X(_04033_));
 sg13g2_buf_1 _20225_ (.A(_04031_),
    .X(_04034_));
 sg13g2_nand2_1 _20226_ (.Y(_04035_),
    .A(\top_ihp.oisc.regs[9][0] ),
    .B(net730));
 sg13g2_o21ai_1 _20227_ (.B1(_04035_),
    .Y(_02468_),
    .A1(net156),
    .A2(net678));
 sg13g2_nand2_1 _20228_ (.Y(_04036_),
    .A(\top_ihp.oisc.regs[9][10] ),
    .B(net730));
 sg13g2_o21ai_1 _20229_ (.B1(_04036_),
    .Y(_02469_),
    .A1(net128),
    .A2(net678));
 sg13g2_nand2_1 _20230_ (.Y(_04037_),
    .A(\top_ihp.oisc.regs[9][11] ),
    .B(net730));
 sg13g2_o21ai_1 _20231_ (.B1(_04037_),
    .Y(_02470_),
    .A1(net127),
    .A2(net678));
 sg13g2_nand2_1 _20232_ (.Y(_04038_),
    .A(\top_ihp.oisc.regs[9][12] ),
    .B(net730));
 sg13g2_o21ai_1 _20233_ (.B1(_04038_),
    .Y(_02471_),
    .A1(_09905_),
    .A2(net678));
 sg13g2_nand2_1 _20234_ (.Y(_04039_),
    .A(\top_ihp.oisc.regs[9][13] ),
    .B(net730));
 sg13g2_o21ai_1 _20235_ (.B1(_04039_),
    .Y(_02472_),
    .A1(net314),
    .A2(net678));
 sg13g2_nand2_1 _20236_ (.Y(_04040_),
    .A(\top_ihp.oisc.regs[9][14] ),
    .B(net730));
 sg13g2_o21ai_1 _20237_ (.B1(_04040_),
    .Y(_02473_),
    .A1(net330),
    .A2(net678));
 sg13g2_nand2_1 _20238_ (.Y(_04041_),
    .A(\top_ihp.oisc.regs[9][15] ),
    .B(net730));
 sg13g2_o21ai_1 _20239_ (.B1(_04041_),
    .Y(_02474_),
    .A1(net329),
    .A2(_04033_));
 sg13g2_nand2_1 _20240_ (.Y(_04042_),
    .A(\top_ihp.oisc.regs[9][16] ),
    .B(net730));
 sg13g2_o21ai_1 _20241_ (.B1(_04042_),
    .Y(_02475_),
    .A1(net126),
    .A2(_04033_));
 sg13g2_buf_1 _20242_ (.A(net731),
    .X(_04043_));
 sg13g2_nand2_1 _20243_ (.Y(_04044_),
    .A(\top_ihp.oisc.regs[9][17] ),
    .B(net677));
 sg13g2_o21ai_1 _20244_ (.B1(_04044_),
    .Y(_02476_),
    .A1(net313),
    .A2(net678));
 sg13g2_nand2_1 _20245_ (.Y(_04045_),
    .A(\top_ihp.oisc.regs[9][18] ),
    .B(net677));
 sg13g2_o21ai_1 _20246_ (.B1(_04045_),
    .Y(_02477_),
    .A1(net312),
    .A2(net678));
 sg13g2_buf_1 _20247_ (.A(net731),
    .X(_04046_));
 sg13g2_nand2_1 _20248_ (.Y(_04047_),
    .A(\top_ihp.oisc.regs[9][19] ),
    .B(net677));
 sg13g2_o21ai_1 _20249_ (.B1(_04047_),
    .Y(_02478_),
    .A1(net311),
    .A2(net676));
 sg13g2_nand2_1 _20250_ (.Y(_04048_),
    .A(\top_ihp.oisc.regs[9][1] ),
    .B(_04043_));
 sg13g2_o21ai_1 _20251_ (.B1(_04048_),
    .Y(_02479_),
    .A1(net325),
    .A2(_04046_));
 sg13g2_nand2_1 _20252_ (.Y(_04049_),
    .A(\top_ihp.oisc.regs[9][20] ),
    .B(net677));
 sg13g2_o21ai_1 _20253_ (.B1(_04049_),
    .Y(_02480_),
    .A1(net607),
    .A2(net676));
 sg13g2_nand2_1 _20254_ (.Y(_04050_),
    .A(\top_ihp.oisc.regs[9][21] ),
    .B(net677));
 sg13g2_o21ai_1 _20255_ (.B1(_04050_),
    .Y(_02481_),
    .A1(net310),
    .A2(net676));
 sg13g2_nand2_1 _20256_ (.Y(_04051_),
    .A(\top_ihp.oisc.regs[9][22] ),
    .B(net677));
 sg13g2_o21ai_1 _20257_ (.B1(_04051_),
    .Y(_02482_),
    .A1(net322),
    .A2(net676));
 sg13g2_nand2_1 _20258_ (.Y(_04052_),
    .A(\top_ihp.oisc.regs[9][23] ),
    .B(net677));
 sg13g2_o21ai_1 _20259_ (.B1(_04052_),
    .Y(_02483_),
    .A1(net528),
    .A2(net676));
 sg13g2_nand2_1 _20260_ (.Y(_04053_),
    .A(\top_ihp.oisc.regs[9][24] ),
    .B(_04043_));
 sg13g2_o21ai_1 _20261_ (.B1(_04053_),
    .Y(_02484_),
    .A1(net309),
    .A2(_04046_));
 sg13g2_nand2_1 _20262_ (.Y(_04054_),
    .A(\top_ihp.oisc.regs[9][25] ),
    .B(net677));
 sg13g2_o21ai_1 _20263_ (.B1(_04054_),
    .Y(_02485_),
    .A1(net319),
    .A2(net676));
 sg13g2_buf_1 _20264_ (.A(net731),
    .X(_04055_));
 sg13g2_nand2_1 _20265_ (.Y(_04056_),
    .A(\top_ihp.oisc.regs[9][26] ),
    .B(_04055_));
 sg13g2_o21ai_1 _20266_ (.B1(_04056_),
    .Y(_02486_),
    .A1(net125),
    .A2(net676));
 sg13g2_nand2_1 _20267_ (.Y(_04057_),
    .A(\top_ihp.oisc.regs[9][27] ),
    .B(net675));
 sg13g2_o21ai_1 _20268_ (.B1(_04057_),
    .Y(_02487_),
    .A1(net308),
    .A2(net676));
 sg13g2_buf_1 _20269_ (.A(net731),
    .X(_04058_));
 sg13g2_nand2_1 _20270_ (.Y(_04059_),
    .A(\top_ihp.oisc.regs[9][28] ),
    .B(net675));
 sg13g2_o21ai_1 _20271_ (.B1(_04059_),
    .Y(_02488_),
    .A1(net515),
    .A2(net674));
 sg13g2_nand2_1 _20272_ (.Y(_04060_),
    .A(\top_ihp.oisc.regs[9][29] ),
    .B(net675));
 sg13g2_o21ai_1 _20273_ (.B1(_04060_),
    .Y(_02489_),
    .A1(net307),
    .A2(net674));
 sg13g2_nand2_1 _20274_ (.Y(_04061_),
    .A(\top_ihp.oisc.regs[9][2] ),
    .B(_04055_));
 sg13g2_o21ai_1 _20275_ (.B1(_04061_),
    .Y(_02490_),
    .A1(net131),
    .A2(_04058_));
 sg13g2_nand2_1 _20276_ (.Y(_04062_),
    .A(\top_ihp.oisc.regs[9][30] ),
    .B(net675));
 sg13g2_o21ai_1 _20277_ (.B1(_04062_),
    .Y(_02491_),
    .A1(_10643_),
    .A2(net674));
 sg13g2_nand2_1 _20278_ (.Y(_04063_),
    .A(\top_ihp.oisc.regs[9][31] ),
    .B(net675));
 sg13g2_o21ai_1 _20279_ (.B1(_04063_),
    .Y(_02492_),
    .A1(net306),
    .A2(net674));
 sg13g2_nand2_1 _20280_ (.Y(_04064_),
    .A(\top_ihp.oisc.regs[9][3] ),
    .B(net675));
 sg13g2_o21ai_1 _20281_ (.B1(_04064_),
    .Y(_02493_),
    .A1(net130),
    .A2(net674));
 sg13g2_nand2_1 _20282_ (.Y(_04065_),
    .A(\top_ihp.oisc.regs[9][4] ),
    .B(net675));
 sg13g2_o21ai_1 _20283_ (.B1(_04065_),
    .Y(_02494_),
    .A1(net129),
    .A2(net674));
 sg13g2_nand2_1 _20284_ (.Y(_04066_),
    .A(\top_ihp.oisc.regs[9][5] ),
    .B(net675));
 sg13g2_o21ai_1 _20285_ (.B1(_04066_),
    .Y(_02495_),
    .A1(net123),
    .A2(net674));
 sg13g2_nand2_1 _20286_ (.Y(_04067_),
    .A(\top_ihp.oisc.regs[9][6] ),
    .B(net731));
 sg13g2_o21ai_1 _20287_ (.B1(_04067_),
    .Y(_02496_),
    .A1(net122),
    .A2(_04058_));
 sg13g2_nand2_1 _20288_ (.Y(_04068_),
    .A(\top_ihp.oisc.regs[9][7] ),
    .B(net731));
 sg13g2_o21ai_1 _20289_ (.B1(_04068_),
    .Y(_02497_),
    .A1(net470),
    .A2(net674));
 sg13g2_nand2_1 _20290_ (.Y(_04069_),
    .A(\top_ihp.oisc.regs[9][8] ),
    .B(_04032_));
 sg13g2_o21ai_1 _20291_ (.B1(_04069_),
    .Y(_02498_),
    .A1(net305),
    .A2(_04034_));
 sg13g2_nand2_1 _20292_ (.Y(_04070_),
    .A(\top_ihp.oisc.regs[9][9] ),
    .B(net731));
 sg13g2_o21ai_1 _20293_ (.B1(_04070_),
    .Y(_02499_),
    .A1(net121),
    .A2(_04034_));
 sg13g2_a21oi_1 _20294_ (.A1(_07958_),
    .A2(net856),
    .Y(_04071_),
    .B1(net1058));
 sg13g2_nand2_1 _20295_ (.Y(_04072_),
    .A(net922),
    .B(_04071_));
 sg13g2_o21ai_1 _20296_ (.B1(_04072_),
    .Y(_04073_),
    .A1(_13600_),
    .A2(net922));
 sg13g2_nand2_1 _20297_ (.Y(_04074_),
    .A(_07985_),
    .B(_08825_));
 sg13g2_buf_1 _20298_ (.A(_04074_),
    .X(_04075_));
 sg13g2_inv_1 _20299_ (.Y(_04076_),
    .A(_08823_));
 sg13g2_a221oi_1 _20300_ (.B2(_04076_),
    .C1(net1049),
    .B1(_04075_),
    .A1(_13600_),
    .Y(_04077_),
    .A2(_08825_));
 sg13g2_a21oi_1 _20301_ (.A1(net1049),
    .A2(_04073_),
    .Y(_02500_),
    .B1(_04077_));
 sg13g2_buf_2 _20302_ (.A(_09735_),
    .X(_04078_));
 sg13g2_buf_1 _20303_ (.A(net1021),
    .X(_04079_));
 sg13g2_buf_1 _20304_ (.A(_00073_),
    .X(_04080_));
 sg13g2_nand3_1 _20305_ (.B(_04080_),
    .C(net806),
    .A(_04079_),
    .Y(_04081_));
 sg13g2_nor2_1 _20306_ (.A(_07973_),
    .B(_04081_),
    .Y(_04082_));
 sg13g2_a21oi_1 _20307_ (.A1(net939),
    .A2(_07973_),
    .Y(_04083_),
    .B1(_04082_));
 sg13g2_nor2_1 _20308_ (.A(_08310_),
    .B(_08802_),
    .Y(_04084_));
 sg13g2_buf_1 _20309_ (.A(_04084_),
    .X(_04085_));
 sg13g2_buf_2 _20310_ (.A(net835),
    .X(_04086_));
 sg13g2_buf_1 _20311_ (.A(_04086_),
    .X(_04087_));
 sg13g2_buf_1 _20312_ (.A(net783),
    .X(_04088_));
 sg13g2_nor2_1 _20313_ (.A(net1049),
    .B(net760),
    .Y(_04089_));
 sg13g2_a22oi_1 _20314_ (.Y(_02501_),
    .B1(_04089_),
    .B2(_04081_),
    .A2(_04083_),
    .A1(net1049));
 sg13g2_o21ai_1 _20315_ (.B1(_08821_),
    .Y(_04090_),
    .A1(_07960_),
    .A2(net806));
 sg13g2_nor2_1 _20316_ (.A(_08220_),
    .B(net856),
    .Y(_04091_));
 sg13g2_buf_8 _20317_ (.A(_04091_),
    .X(_04092_));
 sg13g2_buf_1 _20318_ (.A(_04092_),
    .X(_04093_));
 sg13g2_nand2_1 _20319_ (.Y(_04094_),
    .A(_04080_),
    .B(_04093_));
 sg13g2_nand2_1 _20320_ (.Y(_04095_),
    .A(net1052),
    .B(_04090_));
 sg13g2_o21ai_1 _20321_ (.B1(_04095_),
    .Y(_02502_),
    .A1(_04090_),
    .A2(_04094_));
 sg13g2_nand3_1 _20322_ (.B(_04080_),
    .C(net806),
    .A(net1052),
    .Y(_04096_));
 sg13g2_o21ai_1 _20323_ (.B1(_04096_),
    .Y(_04097_),
    .A1(_09532_),
    .A2(net806));
 sg13g2_nand4_1 _20324_ (.B(_04080_),
    .C(net922),
    .A(net1052),
    .Y(_04098_),
    .D(net806));
 sg13g2_o21ai_1 _20325_ (.B1(_04098_),
    .Y(_04099_),
    .A1(_09532_),
    .A2(_08821_));
 sg13g2_a21o_1 _20326_ (.A2(_04097_),
    .A1(_07961_),
    .B1(_04099_),
    .X(_02503_));
 sg13g2_nand3_1 _20327_ (.B(_04080_),
    .C(net806),
    .A(_09495_),
    .Y(_04100_));
 sg13g2_o21ai_1 _20328_ (.B1(_04100_),
    .Y(_04101_),
    .A1(_09596_),
    .A2(net806));
 sg13g2_nand4_1 _20329_ (.B(_04080_),
    .C(net922),
    .A(net1031),
    .Y(_04102_),
    .D(_08827_));
 sg13g2_o21ai_1 _20330_ (.B1(_04102_),
    .Y(_04103_),
    .A1(net995),
    .A2(_08821_));
 sg13g2_a21o_1 _20331_ (.A2(_04101_),
    .A1(_07961_),
    .B1(_04103_),
    .X(_02504_));
 sg13g2_nand2b_1 _20332_ (.Y(_04104_),
    .B(_07974_),
    .A_N(_04071_));
 sg13g2_o21ai_1 _20333_ (.B1(_08821_),
    .Y(_04105_),
    .A1(net1049),
    .A2(_08802_));
 sg13g2_nand2_1 _20334_ (.Y(_04106_),
    .A(_08823_),
    .B(_04105_));
 sg13g2_nand2_1 _20335_ (.Y(_02505_),
    .A(_04104_),
    .B(_04106_));
 sg13g2_nand2_1 _20336_ (.Y(_04107_),
    .A(_07958_),
    .B(_09495_));
 sg13g2_buf_1 _20337_ (.A(_04107_),
    .X(_04108_));
 sg13g2_buf_1 _20338_ (.A(_04108_),
    .X(_04109_));
 sg13g2_buf_1 _20339_ (.A(\top_ihp.oisc.wb_dat_o[0] ),
    .X(_04110_));
 sg13g2_buf_1 _20340_ (.A(_04108_),
    .X(_04111_));
 sg13g2_nand2_1 _20341_ (.Y(_04112_),
    .A(net1050),
    .B(net910));
 sg13g2_o21ai_1 _20342_ (.B1(_04112_),
    .Y(_02506_),
    .A1(_09697_),
    .A2(_04109_));
 sg13g2_buf_2 _20343_ (.A(\top_ihp.oisc.wb_dat_o[10] ),
    .X(_04113_));
 sg13g2_nand2_1 _20344_ (.Y(_04114_),
    .A(_04113_),
    .B(net910));
 sg13g2_o21ai_1 _20345_ (.B1(_04114_),
    .Y(_02507_),
    .A1(net128),
    .A2(net911));
 sg13g2_buf_2 _20346_ (.A(\top_ihp.oisc.wb_dat_o[11] ),
    .X(_04115_));
 sg13g2_nand2_1 _20347_ (.Y(_04116_),
    .A(_04115_),
    .B(net910));
 sg13g2_o21ai_1 _20348_ (.B1(_04116_),
    .Y(_02508_),
    .A1(net127),
    .A2(net911));
 sg13g2_buf_2 _20349_ (.A(\top_ihp.oisc.wb_dat_o[12] ),
    .X(_04117_));
 sg13g2_nand2_1 _20350_ (.Y(_04118_),
    .A(_04117_),
    .B(net910));
 sg13g2_o21ai_1 _20351_ (.B1(_04118_),
    .Y(_02509_),
    .A1(net332),
    .A2(net911));
 sg13g2_buf_2 _20352_ (.A(\top_ihp.oisc.wb_dat_o[13] ),
    .X(_04119_));
 sg13g2_nand2_1 _20353_ (.Y(_04120_),
    .A(_04119_),
    .B(net910));
 sg13g2_o21ai_1 _20354_ (.B1(_04120_),
    .Y(_02510_),
    .A1(_08234_),
    .A2(net911));
 sg13g2_buf_2 _20355_ (.A(\top_ihp.oisc.wb_dat_o[14] ),
    .X(_04121_));
 sg13g2_buf_1 _20356_ (.A(_04108_),
    .X(_04122_));
 sg13g2_mux2_1 _20357_ (.A0(net1067),
    .A1(_04121_),
    .S(net909),
    .X(_02511_));
 sg13g2_inv_1 _20358_ (.Y(_04123_),
    .A(net1068));
 sg13g2_buf_2 _20359_ (.A(\top_ihp.oisc.wb_dat_o[15] ),
    .X(_04124_));
 sg13g2_nand2_1 _20360_ (.Y(_04125_),
    .A(_04124_),
    .B(net910));
 sg13g2_o21ai_1 _20361_ (.B1(_04125_),
    .Y(_02512_),
    .A1(_04123_),
    .A2(net911));
 sg13g2_buf_2 _20362_ (.A(\top_ihp.oisc.wb_dat_o[16] ),
    .X(_04126_));
 sg13g2_nand2_1 _20363_ (.Y(_04127_),
    .A(_04126_),
    .B(net910));
 sg13g2_o21ai_1 _20364_ (.B1(_04127_),
    .Y(_02513_),
    .A1(_10628_),
    .A2(net911));
 sg13g2_buf_2 _20365_ (.A(\top_ihp.oisc.wb_dat_o[17] ),
    .X(_04128_));
 sg13g2_nand2_1 _20366_ (.Y(_04129_),
    .A(_04128_),
    .B(net910));
 sg13g2_o21ai_1 _20367_ (.B1(_04129_),
    .Y(_02514_),
    .A1(net313),
    .A2(net911));
 sg13g2_buf_2 _20368_ (.A(\top_ihp.oisc.wb_dat_o[18] ),
    .X(_04130_));
 sg13g2_buf_1 _20369_ (.A(_04108_),
    .X(_04131_));
 sg13g2_nand2_1 _20370_ (.Y(_04132_),
    .A(_04130_),
    .B(net908));
 sg13g2_o21ai_1 _20371_ (.B1(_04132_),
    .Y(_02515_),
    .A1(net312),
    .A2(net911));
 sg13g2_buf_1 _20372_ (.A(_04108_),
    .X(_04133_));
 sg13g2_buf_1 _20373_ (.A(\top_ihp.oisc.wb_dat_o[19] ),
    .X(_04134_));
 sg13g2_nand2_1 _20374_ (.Y(_04135_),
    .A(_04134_),
    .B(net908));
 sg13g2_o21ai_1 _20375_ (.B1(_04135_),
    .Y(_02516_),
    .A1(_08000_),
    .A2(net907));
 sg13g2_buf_2 _20376_ (.A(\top_ihp.oisc.wb_dat_o[1] ),
    .X(_04136_));
 sg13g2_nand2_1 _20377_ (.Y(_04137_),
    .A(_04136_),
    .B(net908));
 sg13g2_o21ai_1 _20378_ (.B1(_04137_),
    .Y(_02517_),
    .A1(_10127_),
    .A2(net907));
 sg13g2_buf_1 _20379_ (.A(\top_ihp.oisc.wb_dat_o[20] ),
    .X(_04138_));
 sg13g2_nand2_1 _20380_ (.Y(_04139_),
    .A(_04138_),
    .B(net908));
 sg13g2_o21ai_1 _20381_ (.B1(_04139_),
    .Y(_02518_),
    .A1(_10150_),
    .A2(net907));
 sg13g2_buf_1 _20382_ (.A(\top_ihp.oisc.wb_dat_o[21] ),
    .X(_04140_));
 sg13g2_nand2_1 _20383_ (.Y(_04141_),
    .A(_04140_),
    .B(_04131_));
 sg13g2_o21ai_1 _20384_ (.B1(_04141_),
    .Y(_02519_),
    .A1(net310),
    .A2(_04133_));
 sg13g2_buf_1 _20385_ (.A(\top_ihp.oisc.wb_dat_o[22] ),
    .X(_04142_));
 sg13g2_nand2_1 _20386_ (.Y(_04143_),
    .A(_04142_),
    .B(net908));
 sg13g2_o21ai_1 _20387_ (.B1(_04143_),
    .Y(_02520_),
    .A1(_10188_),
    .A2(net907));
 sg13g2_buf_1 _20388_ (.A(\top_ihp.oisc.wb_dat_o[23] ),
    .X(_04144_));
 sg13g2_inv_1 _20389_ (.Y(_04145_),
    .A(_04144_));
 sg13g2_buf_1 _20390_ (.A(_04108_),
    .X(_04146_));
 sg13g2_a21oi_1 _20391_ (.A1(net1061),
    .A2(net898),
    .Y(_04147_),
    .B1(_04146_));
 sg13g2_a21oi_1 _20392_ (.A1(_04145_),
    .A2(_04109_),
    .Y(_02521_),
    .B1(_04147_));
 sg13g2_buf_1 _20393_ (.A(\top_ihp.oisc.wb_dat_o[24] ),
    .X(_04148_));
 sg13g2_nand2_1 _20394_ (.Y(_04149_),
    .A(_04148_),
    .B(_04131_));
 sg13g2_o21ai_1 _20395_ (.B1(_04149_),
    .Y(_02522_),
    .A1(_10636_),
    .A2(net907));
 sg13g2_buf_1 _20396_ (.A(\top_ihp.oisc.wb_dat_o[25] ),
    .X(_04150_));
 sg13g2_mux2_1 _20397_ (.A0(_08157_),
    .A1(_04150_),
    .S(net909),
    .X(_02523_));
 sg13g2_buf_1 _20398_ (.A(\top_ihp.oisc.wb_dat_o[26] ),
    .X(_04151_));
 sg13g2_nand2_1 _20399_ (.Y(_04152_),
    .A(_04151_),
    .B(net908));
 sg13g2_o21ai_1 _20400_ (.B1(_04152_),
    .Y(_02524_),
    .A1(net974),
    .A2(net907));
 sg13g2_buf_1 _20401_ (.A(\top_ihp.oisc.wb_dat_o[27] ),
    .X(_04153_));
 sg13g2_nand2_1 _20402_ (.Y(_04154_),
    .A(_04153_),
    .B(net908));
 sg13g2_o21ai_1 _20403_ (.B1(_04154_),
    .Y(_02525_),
    .A1(net308),
    .A2(net907));
 sg13g2_buf_1 _20404_ (.A(\top_ihp.oisc.wb_dat_o[28] ),
    .X(_04155_));
 sg13g2_mux2_1 _20405_ (.A0(net1057),
    .A1(_04155_),
    .S(_04111_),
    .X(_02526_));
 sg13g2_buf_1 _20406_ (.A(\top_ihp.oisc.wb_dat_o[29] ),
    .X(_04156_));
 sg13g2_nand2_1 _20407_ (.Y(_04157_),
    .A(_04156_),
    .B(net908));
 sg13g2_o21ai_1 _20408_ (.B1(_04157_),
    .Y(_02527_),
    .A1(net307),
    .A2(_04133_));
 sg13g2_buf_2 _20409_ (.A(\top_ihp.oisc.wb_dat_o[2] ),
    .X(_04158_));
 sg13g2_nand2_1 _20410_ (.Y(_04159_),
    .A(_04158_),
    .B(net906));
 sg13g2_o21ai_1 _20411_ (.B1(_04159_),
    .Y(_02528_),
    .A1(_10604_),
    .A2(net907));
 sg13g2_buf_1 _20412_ (.A(\top_ihp.oisc.wb_dat_o[30] ),
    .X(_04160_));
 sg13g2_nand2_1 _20413_ (.Y(_04161_),
    .A(_04160_),
    .B(net906));
 sg13g2_o21ai_1 _20414_ (.B1(_04161_),
    .Y(_02529_),
    .A1(net124),
    .A2(net909));
 sg13g2_buf_1 _20415_ (.A(\top_ihp.oisc.wb_dat_o[31] ),
    .X(_04162_));
 sg13g2_mux2_1 _20416_ (.A0(_09497_),
    .A1(_04162_),
    .S(_04111_),
    .X(_02530_));
 sg13g2_buf_2 _20417_ (.A(\top_ihp.oisc.wb_dat_o[3] ),
    .X(_04163_));
 sg13g2_nand2_1 _20418_ (.Y(_04164_),
    .A(_04163_),
    .B(net906));
 sg13g2_o21ai_1 _20419_ (.B1(_04164_),
    .Y(_02531_),
    .A1(_10608_),
    .A2(net909));
 sg13g2_buf_2 _20420_ (.A(\top_ihp.oisc.wb_dat_o[4] ),
    .X(_04165_));
 sg13g2_nand2_1 _20421_ (.Y(_04166_),
    .A(_04165_),
    .B(net906));
 sg13g2_o21ai_1 _20422_ (.B1(_04166_),
    .Y(_02532_),
    .A1(_10609_),
    .A2(net909));
 sg13g2_buf_2 _20423_ (.A(\top_ihp.oisc.wb_dat_o[5] ),
    .X(_04167_));
 sg13g2_nand2_1 _20424_ (.Y(_04168_),
    .A(_04167_),
    .B(net906));
 sg13g2_o21ai_1 _20425_ (.B1(_04168_),
    .Y(_02533_),
    .A1(net123),
    .A2(net909));
 sg13g2_buf_2 _20426_ (.A(\top_ihp.oisc.wb_dat_o[6] ),
    .X(_04169_));
 sg13g2_nand2_1 _20427_ (.Y(_04170_),
    .A(_04169_),
    .B(net906));
 sg13g2_o21ai_1 _20428_ (.B1(_04170_),
    .Y(_02534_),
    .A1(_10646_),
    .A2(_04122_));
 sg13g2_buf_2 _20429_ (.A(\top_ihp.oisc.wb_dat_o[7] ),
    .X(_04171_));
 sg13g2_nand2_1 _20430_ (.Y(_04172_),
    .A(_04171_),
    .B(net906));
 sg13g2_o21ai_1 _20431_ (.B1(_04172_),
    .Y(_02535_),
    .A1(_10481_),
    .A2(_04122_));
 sg13g2_buf_2 _20432_ (.A(\top_ihp.oisc.wb_dat_o[8] ),
    .X(_04173_));
 sg13g2_nand2_1 _20433_ (.Y(_04174_),
    .A(_04173_),
    .B(net906));
 sg13g2_o21ai_1 _20434_ (.B1(_04174_),
    .Y(_02536_),
    .A1(_10647_),
    .A2(net909));
 sg13g2_buf_2 _20435_ (.A(\top_ihp.oisc.wb_dat_o[9] ),
    .X(_04175_));
 sg13g2_nand2_1 _20436_ (.Y(_04176_),
    .A(_04175_),
    .B(_04146_));
 sg13g2_o21ai_1 _20437_ (.B1(_04176_),
    .Y(_02537_),
    .A1(_10648_),
    .A2(net909));
 sg13g2_inv_1 _20438_ (.Y(_04177_),
    .A(\top_ihp.wb_coproc.opa[0] ));
 sg13g2_inv_1 _20439_ (.Y(_04178_),
    .A(_08087_));
 sg13g2_xnor2_1 _20440_ (.Y(_04179_),
    .A(_04178_),
    .B(_10366_));
 sg13g2_nor2_1 _20441_ (.A(_08086_),
    .B(_08223_),
    .Y(_04180_));
 sg13g2_o21ai_1 _20442_ (.B1(net1017),
    .Y(_04181_),
    .A1(_08223_),
    .A2(_04179_));
 sg13g2_and2_1 _20443_ (.A(_08086_),
    .B(_04181_),
    .X(_04182_));
 sg13g2_a21oi_2 _20444_ (.B1(_04182_),
    .Y(_04183_),
    .A2(_04180_),
    .A1(_04179_));
 sg13g2_o21ai_1 _20445_ (.B1(net1017),
    .Y(_04184_),
    .A1(_08210_),
    .A2(_10397_));
 sg13g2_nor2_1 _20446_ (.A(_08109_),
    .B(_08223_),
    .Y(_04185_));
 sg13g2_a22oi_1 _20447_ (.Y(_04186_),
    .B1(_04185_),
    .B2(_10397_),
    .A2(_04184_),
    .A1(_08109_));
 sg13g2_buf_2 _20448_ (.A(_04186_),
    .X(_04187_));
 sg13g2_inv_1 _20449_ (.Y(_04188_),
    .A(_04187_));
 sg13g2_inv_1 _20450_ (.Y(_04189_),
    .A(_09508_));
 sg13g2_or2_1 _20451_ (.X(_04190_),
    .B(_08082_),
    .A(_08078_));
 sg13g2_a22oi_1 _20452_ (.Y(_04191_),
    .B1(_04190_),
    .B2(net1047),
    .A2(_04189_),
    .A1(_08212_));
 sg13g2_buf_1 _20453_ (.A(_04191_),
    .X(_04192_));
 sg13g2_nand3_1 _20454_ (.B(_04188_),
    .C(_04192_),
    .A(_04183_),
    .Y(_04193_));
 sg13g2_buf_2 _20455_ (.A(_04193_),
    .X(_04194_));
 sg13g2_buf_1 _20456_ (.A(_04194_),
    .X(_04195_));
 sg13g2_a21o_1 _20457_ (.A2(_04180_),
    .A1(_04179_),
    .B1(_04182_),
    .X(_04196_));
 sg13g2_buf_1 _20458_ (.A(_04196_),
    .X(_04197_));
 sg13g2_xor2_1 _20459_ (.B(_10299_),
    .A(_08091_),
    .X(_04198_));
 sg13g2_a21o_1 _20460_ (.A2(_04198_),
    .A1(_08212_),
    .B1(net1047),
    .X(_04199_));
 sg13g2_nor3_1 _20461_ (.A(_08090_),
    .B(_08223_),
    .C(_04198_),
    .Y(_04200_));
 sg13g2_a21o_1 _20462_ (.A2(_04199_),
    .A1(_08090_),
    .B1(_04200_),
    .X(_04201_));
 sg13g2_buf_2 _20463_ (.A(_04201_),
    .X(_04202_));
 sg13g2_nand4_1 _20464_ (.B(_04187_),
    .C(_04192_),
    .A(_04197_),
    .Y(_04203_),
    .D(_04202_));
 sg13g2_buf_2 _20465_ (.A(_04203_),
    .X(_04204_));
 sg13g2_buf_1 _20466_ (.A(_04204_),
    .X(_04205_));
 sg13g2_mux2_1 _20467_ (.A0(net564),
    .A1(net563),
    .S(\top_ihp.wb_coproc.opb[0] ),
    .X(_04206_));
 sg13g2_inv_1 _20468_ (.Y(_04207_),
    .A(_04192_));
 sg13g2_nor3_1 _20469_ (.A(_04197_),
    .B(_04187_),
    .C(_04207_),
    .Y(_04208_));
 sg13g2_buf_2 _20470_ (.A(_04208_),
    .X(_04209_));
 sg13g2_buf_1 _20471_ (.A(_04209_),
    .X(_04210_));
 sg13g2_buf_1 _20472_ (.A(_04202_),
    .X(_04211_));
 sg13g2_nand2_1 _20473_ (.Y(_04212_),
    .A(\top_ihp.wb_coproc.opa[0] ),
    .B(net740));
 sg13g2_nand3_1 _20474_ (.B(net562),
    .C(_04212_),
    .A(\top_ihp.wb_coproc.opb[0] ),
    .Y(_04213_));
 sg13g2_o21ai_1 _20475_ (.B1(_04213_),
    .Y(_04214_),
    .A1(_04177_),
    .A2(_04206_));
 sg13g2_and2_1 _20476_ (.A(_08207_),
    .B(_00003_),
    .X(_04215_));
 sg13g2_buf_2 _20477_ (.A(_04215_),
    .X(_04216_));
 sg13g2_buf_8 _20478_ (.A(_04216_),
    .X(_04217_));
 sg13g2_mux2_1 _20479_ (.A0(\top_ihp.wb_coproc.dat_o[0] ),
    .A1(_04214_),
    .S(_04217_),
    .X(_02538_));
 sg13g2_inv_1 _20480_ (.Y(_04218_),
    .A(\top_ihp.wb_coproc.opa[10] ));
 sg13g2_mux2_1 _20481_ (.A0(_04195_),
    .A1(_04205_),
    .S(\top_ihp.wb_coproc.opb[10] ),
    .X(_04219_));
 sg13g2_nand2_1 _20482_ (.Y(_04220_),
    .A(\top_ihp.wb_coproc.opa[10] ),
    .B(_04211_));
 sg13g2_nand3_1 _20483_ (.B(_04210_),
    .C(_04220_),
    .A(\top_ihp.wb_coproc.opb[10] ),
    .Y(_04221_));
 sg13g2_o21ai_1 _20484_ (.B1(_04221_),
    .Y(_04222_),
    .A1(_04218_),
    .A2(_04219_));
 sg13g2_mux2_1 _20485_ (.A0(\top_ihp.wb_coproc.dat_o[10] ),
    .A1(_04222_),
    .S(net219),
    .X(_02539_));
 sg13g2_inv_1 _20486_ (.Y(_04223_),
    .A(\top_ihp.wb_coproc.opa[11] ));
 sg13g2_mux2_1 _20487_ (.A0(net564),
    .A1(net563),
    .S(\top_ihp.wb_coproc.opb[11] ),
    .X(_04224_));
 sg13g2_nand2_1 _20488_ (.Y(_04225_),
    .A(\top_ihp.wb_coproc.opa[11] ),
    .B(net740));
 sg13g2_nand3_1 _20489_ (.B(net562),
    .C(_04225_),
    .A(\top_ihp.wb_coproc.opb[11] ),
    .Y(_04226_));
 sg13g2_o21ai_1 _20490_ (.B1(_04226_),
    .Y(_04227_),
    .A1(_04223_),
    .A2(_04224_));
 sg13g2_mux2_1 _20491_ (.A0(\top_ihp.wb_coproc.dat_o[11] ),
    .A1(_04227_),
    .S(net219),
    .X(_02540_));
 sg13g2_inv_1 _20492_ (.Y(_04228_),
    .A(\top_ihp.wb_coproc.opa[12] ));
 sg13g2_mux2_1 _20493_ (.A0(net564),
    .A1(net563),
    .S(\top_ihp.wb_coproc.opb[12] ),
    .X(_04229_));
 sg13g2_nand2_1 _20494_ (.Y(_04230_),
    .A(\top_ihp.wb_coproc.opa[12] ),
    .B(net740));
 sg13g2_nand3_1 _20495_ (.B(net562),
    .C(_04230_),
    .A(\top_ihp.wb_coproc.opb[12] ),
    .Y(_04231_));
 sg13g2_o21ai_1 _20496_ (.B1(_04231_),
    .Y(_04232_),
    .A1(_04228_),
    .A2(_04229_));
 sg13g2_mux2_1 _20497_ (.A0(\top_ihp.wb_coproc.dat_o[12] ),
    .A1(_04232_),
    .S(net219),
    .X(_02541_));
 sg13g2_inv_1 _20498_ (.Y(_04233_),
    .A(\top_ihp.wb_coproc.opa[13] ));
 sg13g2_mux2_1 _20499_ (.A0(net564),
    .A1(net563),
    .S(\top_ihp.wb_coproc.opb[13] ),
    .X(_04234_));
 sg13g2_nand2_1 _20500_ (.Y(_04235_),
    .A(\top_ihp.wb_coproc.opa[13] ),
    .B(net740));
 sg13g2_nand3_1 _20501_ (.B(net562),
    .C(_04235_),
    .A(\top_ihp.wb_coproc.opb[13] ),
    .Y(_04236_));
 sg13g2_o21ai_1 _20502_ (.B1(_04236_),
    .Y(_04237_),
    .A1(_04233_),
    .A2(_04234_));
 sg13g2_mux2_1 _20503_ (.A0(\top_ihp.wb_coproc.dat_o[13] ),
    .A1(_04237_),
    .S(_04217_),
    .X(_02542_));
 sg13g2_inv_1 _20504_ (.Y(_04238_),
    .A(\top_ihp.wb_coproc.opa[14] ));
 sg13g2_mux2_1 _20505_ (.A0(net564),
    .A1(net563),
    .S(\top_ihp.wb_coproc.opb[14] ),
    .X(_04239_));
 sg13g2_nand2_1 _20506_ (.Y(_04240_),
    .A(\top_ihp.wb_coproc.opa[14] ),
    .B(net740));
 sg13g2_nand3_1 _20507_ (.B(net562),
    .C(_04240_),
    .A(\top_ihp.wb_coproc.opb[14] ),
    .Y(_04241_));
 sg13g2_o21ai_1 _20508_ (.B1(_04241_),
    .Y(_04242_),
    .A1(_04238_),
    .A2(_04239_));
 sg13g2_mux2_1 _20509_ (.A0(\top_ihp.wb_coproc.dat_o[14] ),
    .A1(_04242_),
    .S(net219),
    .X(_02543_));
 sg13g2_inv_1 _20510_ (.Y(_04243_),
    .A(\top_ihp.wb_coproc.opa[15] ));
 sg13g2_mux2_1 _20511_ (.A0(_04195_),
    .A1(_04205_),
    .S(\top_ihp.wb_coproc.opb[15] ),
    .X(_04244_));
 sg13g2_nand2_1 _20512_ (.Y(_04245_),
    .A(\top_ihp.wb_coproc.opa[15] ),
    .B(net740));
 sg13g2_nand3_1 _20513_ (.B(_04210_),
    .C(_04245_),
    .A(\top_ihp.wb_coproc.opb[15] ),
    .Y(_04246_));
 sg13g2_o21ai_1 _20514_ (.B1(_04246_),
    .Y(_04247_),
    .A1(_04243_),
    .A2(_04244_));
 sg13g2_mux2_1 _20515_ (.A0(\top_ihp.wb_coproc.dat_o[15] ),
    .A1(_04247_),
    .S(net219),
    .X(_02544_));
 sg13g2_inv_1 _20516_ (.Y(_04248_),
    .A(\top_ihp.wb_coproc.opa[16] ));
 sg13g2_mux2_1 _20517_ (.A0(net564),
    .A1(net563),
    .S(\top_ihp.wb_coproc.opb[16] ),
    .X(_04249_));
 sg13g2_nand2_1 _20518_ (.Y(_04250_),
    .A(\top_ihp.wb_coproc.opa[16] ),
    .B(net740));
 sg13g2_nand3_1 _20519_ (.B(net562),
    .C(_04250_),
    .A(\top_ihp.wb_coproc.opb[16] ),
    .Y(_04251_));
 sg13g2_o21ai_1 _20520_ (.B1(_04251_),
    .Y(_04252_),
    .A1(_04248_),
    .A2(_04249_));
 sg13g2_mux2_1 _20521_ (.A0(\top_ihp.wb_coproc.dat_o[16] ),
    .A1(_04252_),
    .S(net219),
    .X(_02545_));
 sg13g2_inv_1 _20522_ (.Y(_04253_),
    .A(\top_ihp.wb_coproc.opa[17] ));
 sg13g2_mux2_1 _20523_ (.A0(net564),
    .A1(net563),
    .S(\top_ihp.wb_coproc.opb[17] ),
    .X(_04254_));
 sg13g2_nand2_1 _20524_ (.Y(_04255_),
    .A(\top_ihp.wb_coproc.opa[17] ),
    .B(_04211_));
 sg13g2_nand3_1 _20525_ (.B(net562),
    .C(_04255_),
    .A(\top_ihp.wb_coproc.opb[17] ),
    .Y(_04256_));
 sg13g2_o21ai_1 _20526_ (.B1(_04256_),
    .Y(_04257_),
    .A1(_04253_),
    .A2(_04254_));
 sg13g2_mux2_1 _20527_ (.A0(\top_ihp.wb_coproc.dat_o[17] ),
    .A1(_04257_),
    .S(net219),
    .X(_02546_));
 sg13g2_inv_1 _20528_ (.Y(_04258_),
    .A(\top_ihp.wb_coproc.opa[18] ));
 sg13g2_mux2_1 _20529_ (.A0(net564),
    .A1(net563),
    .S(\top_ihp.wb_coproc.opb[18] ),
    .X(_04259_));
 sg13g2_nand2_1 _20530_ (.Y(_04260_),
    .A(\top_ihp.wb_coproc.opa[18] ),
    .B(net740));
 sg13g2_nand3_1 _20531_ (.B(net562),
    .C(_04260_),
    .A(\top_ihp.wb_coproc.opb[18] ),
    .Y(_04261_));
 sg13g2_o21ai_1 _20532_ (.B1(_04261_),
    .Y(_04262_),
    .A1(_04258_),
    .A2(_04259_));
 sg13g2_mux2_1 _20533_ (.A0(\top_ihp.wb_coproc.dat_o[18] ),
    .A1(_04262_),
    .S(net219),
    .X(_02547_));
 sg13g2_inv_1 _20534_ (.Y(_04263_),
    .A(\top_ihp.wb_coproc.opa[19] ));
 sg13g2_buf_1 _20535_ (.A(_04194_),
    .X(_04264_));
 sg13g2_buf_1 _20536_ (.A(_04204_),
    .X(_04265_));
 sg13g2_mux2_1 _20537_ (.A0(net561),
    .A1(net560),
    .S(\top_ihp.wb_coproc.opb[19] ),
    .X(_04266_));
 sg13g2_buf_1 _20538_ (.A(_04209_),
    .X(_04267_));
 sg13g2_buf_1 _20539_ (.A(_04202_),
    .X(_04268_));
 sg13g2_nand2_1 _20540_ (.Y(_04269_),
    .A(\top_ihp.wb_coproc.opa[19] ),
    .B(net739));
 sg13g2_nand3_1 _20541_ (.B(net559),
    .C(_04269_),
    .A(\top_ihp.wb_coproc.opb[19] ),
    .Y(_04270_));
 sg13g2_o21ai_1 _20542_ (.B1(_04270_),
    .Y(_04271_),
    .A1(_04263_),
    .A2(_04266_));
 sg13g2_buf_8 _20543_ (.A(_04216_),
    .X(_04272_));
 sg13g2_mux2_1 _20544_ (.A0(\top_ihp.wb_coproc.dat_o[19] ),
    .A1(_04271_),
    .S(_04272_),
    .X(_02548_));
 sg13g2_inv_1 _20545_ (.Y(_04273_),
    .A(\top_ihp.wb_coproc.opa[1] ));
 sg13g2_mux2_1 _20546_ (.A0(net561),
    .A1(net560),
    .S(\top_ihp.wb_coproc.opb[1] ),
    .X(_04274_));
 sg13g2_nand2_1 _20547_ (.Y(_04275_),
    .A(\top_ihp.wb_coproc.opa[1] ),
    .B(net739));
 sg13g2_nand3_1 _20548_ (.B(net559),
    .C(_04275_),
    .A(\top_ihp.wb_coproc.opb[1] ),
    .Y(_04276_));
 sg13g2_o21ai_1 _20549_ (.B1(_04276_),
    .Y(_04277_),
    .A1(_04273_),
    .A2(_04274_));
 sg13g2_mux2_1 _20550_ (.A0(\top_ihp.wb_coproc.dat_o[1] ),
    .A1(_04277_),
    .S(net218),
    .X(_02549_));
 sg13g2_inv_1 _20551_ (.Y(_04278_),
    .A(\top_ihp.wb_coproc.opa[20] ));
 sg13g2_mux2_1 _20552_ (.A0(net561),
    .A1(net560),
    .S(\top_ihp.wb_coproc.opb[20] ),
    .X(_04279_));
 sg13g2_nand2_1 _20553_ (.Y(_04280_),
    .A(\top_ihp.wb_coproc.opa[20] ),
    .B(net739));
 sg13g2_nand3_1 _20554_ (.B(net559),
    .C(_04280_),
    .A(\top_ihp.wb_coproc.opb[20] ),
    .Y(_04281_));
 sg13g2_o21ai_1 _20555_ (.B1(_04281_),
    .Y(_04282_),
    .A1(_04278_),
    .A2(_04279_));
 sg13g2_mux2_1 _20556_ (.A0(\top_ihp.wb_coproc.dat_o[20] ),
    .A1(_04282_),
    .S(net218),
    .X(_02550_));
 sg13g2_inv_1 _20557_ (.Y(_04283_),
    .A(\top_ihp.wb_coproc.opa[21] ));
 sg13g2_mux2_1 _20558_ (.A0(net561),
    .A1(net560),
    .S(\top_ihp.wb_coproc.opb[21] ),
    .X(_04284_));
 sg13g2_nand2_1 _20559_ (.Y(_04285_),
    .A(\top_ihp.wb_coproc.opa[21] ),
    .B(net739));
 sg13g2_nand3_1 _20560_ (.B(net559),
    .C(_04285_),
    .A(\top_ihp.wb_coproc.opb[21] ),
    .Y(_04286_));
 sg13g2_o21ai_1 _20561_ (.B1(_04286_),
    .Y(_04287_),
    .A1(_04283_),
    .A2(_04284_));
 sg13g2_mux2_1 _20562_ (.A0(\top_ihp.wb_coproc.dat_o[21] ),
    .A1(_04287_),
    .S(net218),
    .X(_02551_));
 sg13g2_inv_1 _20563_ (.Y(_04288_),
    .A(\top_ihp.wb_coproc.opa[22] ));
 sg13g2_mux2_1 _20564_ (.A0(net561),
    .A1(net560),
    .S(\top_ihp.wb_coproc.opb[22] ),
    .X(_04289_));
 sg13g2_nand2_1 _20565_ (.Y(_04290_),
    .A(\top_ihp.wb_coproc.opa[22] ),
    .B(net739));
 sg13g2_nand3_1 _20566_ (.B(net559),
    .C(_04290_),
    .A(\top_ihp.wb_coproc.opb[22] ),
    .Y(_04291_));
 sg13g2_o21ai_1 _20567_ (.B1(_04291_),
    .Y(_04292_),
    .A1(_04288_),
    .A2(_04289_));
 sg13g2_mux2_1 _20568_ (.A0(\top_ihp.wb_coproc.dat_o[22] ),
    .A1(_04292_),
    .S(net218),
    .X(_02552_));
 sg13g2_inv_1 _20569_ (.Y(_04293_),
    .A(\top_ihp.wb_coproc.opa[23] ));
 sg13g2_mux2_1 _20570_ (.A0(net561),
    .A1(net560),
    .S(\top_ihp.wb_coproc.opb[23] ),
    .X(_04294_));
 sg13g2_nand2_1 _20571_ (.Y(_04295_),
    .A(\top_ihp.wb_coproc.opa[23] ),
    .B(net739));
 sg13g2_nand3_1 _20572_ (.B(net559),
    .C(_04295_),
    .A(\top_ihp.wb_coproc.opb[23] ),
    .Y(_04296_));
 sg13g2_o21ai_1 _20573_ (.B1(_04296_),
    .Y(_04297_),
    .A1(_04293_),
    .A2(_04294_));
 sg13g2_mux2_1 _20574_ (.A0(\top_ihp.wb_coproc.dat_o[23] ),
    .A1(_04297_),
    .S(net218),
    .X(_02553_));
 sg13g2_inv_1 _20575_ (.Y(_04298_),
    .A(\top_ihp.wb_coproc.opa[24] ));
 sg13g2_mux2_1 _20576_ (.A0(_04264_),
    .A1(_04265_),
    .S(\top_ihp.wb_coproc.opb[24] ),
    .X(_04299_));
 sg13g2_nand2_1 _20577_ (.Y(_04300_),
    .A(\top_ihp.wb_coproc.opa[24] ),
    .B(net739));
 sg13g2_nand3_1 _20578_ (.B(_04267_),
    .C(_04300_),
    .A(\top_ihp.wb_coproc.opb[24] ),
    .Y(_04301_));
 sg13g2_o21ai_1 _20579_ (.B1(_04301_),
    .Y(_04302_),
    .A1(_04298_),
    .A2(_04299_));
 sg13g2_mux2_1 _20580_ (.A0(\top_ihp.wb_coproc.dat_o[24] ),
    .A1(_04302_),
    .S(_04272_),
    .X(_02554_));
 sg13g2_inv_1 _20581_ (.Y(_04303_),
    .A(\top_ihp.wb_coproc.opa[25] ));
 sg13g2_mux2_1 _20582_ (.A0(net561),
    .A1(net560),
    .S(\top_ihp.wb_coproc.opb[25] ),
    .X(_04304_));
 sg13g2_nand2_1 _20583_ (.Y(_04305_),
    .A(\top_ihp.wb_coproc.opa[25] ),
    .B(_04268_));
 sg13g2_nand3_1 _20584_ (.B(net559),
    .C(_04305_),
    .A(\top_ihp.wb_coproc.opb[25] ),
    .Y(_04306_));
 sg13g2_o21ai_1 _20585_ (.B1(_04306_),
    .Y(_04307_),
    .A1(_04303_),
    .A2(_04304_));
 sg13g2_mux2_1 _20586_ (.A0(\top_ihp.wb_coproc.dat_o[25] ),
    .A1(_04307_),
    .S(net218),
    .X(_02555_));
 sg13g2_inv_1 _20587_ (.Y(_04308_),
    .A(\top_ihp.wb_coproc.opa[26] ));
 sg13g2_mux2_1 _20588_ (.A0(net561),
    .A1(net560),
    .S(\top_ihp.wb_coproc.opb[26] ),
    .X(_04309_));
 sg13g2_nand2_1 _20589_ (.Y(_04310_),
    .A(\top_ihp.wb_coproc.opa[26] ),
    .B(net739));
 sg13g2_nand3_1 _20590_ (.B(net559),
    .C(_04310_),
    .A(\top_ihp.wb_coproc.opb[26] ),
    .Y(_04311_));
 sg13g2_o21ai_1 _20591_ (.B1(_04311_),
    .Y(_04312_),
    .A1(_04308_),
    .A2(_04309_));
 sg13g2_mux2_1 _20592_ (.A0(\top_ihp.wb_coproc.dat_o[26] ),
    .A1(_04312_),
    .S(net218),
    .X(_02556_));
 sg13g2_inv_1 _20593_ (.Y(_04313_),
    .A(\top_ihp.wb_coproc.opa[27] ));
 sg13g2_mux2_1 _20594_ (.A0(_04264_),
    .A1(_04265_),
    .S(\top_ihp.wb_coproc.opb[27] ),
    .X(_04314_));
 sg13g2_nand2_1 _20595_ (.Y(_04315_),
    .A(\top_ihp.wb_coproc.opa[27] ),
    .B(_04268_));
 sg13g2_nand3_1 _20596_ (.B(_04267_),
    .C(_04315_),
    .A(\top_ihp.wb_coproc.opb[27] ),
    .Y(_04316_));
 sg13g2_o21ai_1 _20597_ (.B1(_04316_),
    .Y(_04317_),
    .A1(_04313_),
    .A2(_04314_));
 sg13g2_mux2_1 _20598_ (.A0(\top_ihp.wb_coproc.dat_o[27] ),
    .A1(_04317_),
    .S(net218),
    .X(_02557_));
 sg13g2_inv_1 _20599_ (.Y(_04318_),
    .A(\top_ihp.wb_coproc.opa[28] ));
 sg13g2_buf_1 _20600_ (.A(_04194_),
    .X(_04319_));
 sg13g2_buf_1 _20601_ (.A(_04204_),
    .X(_04320_));
 sg13g2_mux2_1 _20602_ (.A0(_04319_),
    .A1(_04320_),
    .S(\top_ihp.wb_coproc.opb[28] ),
    .X(_04321_));
 sg13g2_buf_1 _20603_ (.A(_04209_),
    .X(_04322_));
 sg13g2_buf_1 _20604_ (.A(_04202_),
    .X(_04323_));
 sg13g2_nand2_1 _20605_ (.Y(_04324_),
    .A(\top_ihp.wb_coproc.opa[28] ),
    .B(_04323_));
 sg13g2_nand3_1 _20606_ (.B(net556),
    .C(_04324_),
    .A(\top_ihp.wb_coproc.opb[28] ),
    .Y(_04325_));
 sg13g2_o21ai_1 _20607_ (.B1(_04325_),
    .Y(_04326_),
    .A1(_04318_),
    .A2(_04321_));
 sg13g2_buf_8 _20608_ (.A(_04216_),
    .X(_04327_));
 sg13g2_mux2_1 _20609_ (.A0(\top_ihp.wb_coproc.dat_o[28] ),
    .A1(_04326_),
    .S(net217),
    .X(_02558_));
 sg13g2_inv_1 _20610_ (.Y(_04328_),
    .A(\top_ihp.wb_coproc.opa[29] ));
 sg13g2_mux2_1 _20611_ (.A0(_04319_),
    .A1(_04320_),
    .S(\top_ihp.wb_coproc.opb[29] ),
    .X(_04329_));
 sg13g2_nand2_1 _20612_ (.Y(_04330_),
    .A(\top_ihp.wb_coproc.opa[29] ),
    .B(net738));
 sg13g2_nand3_1 _20613_ (.B(net556),
    .C(_04330_),
    .A(\top_ihp.wb_coproc.opb[29] ),
    .Y(_04331_));
 sg13g2_o21ai_1 _20614_ (.B1(_04331_),
    .Y(_04332_),
    .A1(_04328_),
    .A2(_04329_));
 sg13g2_mux2_1 _20615_ (.A0(\top_ihp.wb_coproc.dat_o[29] ),
    .A1(_04332_),
    .S(_04327_),
    .X(_02559_));
 sg13g2_inv_1 _20616_ (.Y(_04333_),
    .A(\top_ihp.wb_coproc.opa[2] ));
 sg13g2_mux2_1 _20617_ (.A0(net558),
    .A1(net557),
    .S(\top_ihp.wb_coproc.opb[2] ),
    .X(_04334_));
 sg13g2_nand2_1 _20618_ (.Y(_04335_),
    .A(\top_ihp.wb_coproc.opa[2] ),
    .B(net738));
 sg13g2_nand3_1 _20619_ (.B(net556),
    .C(_04335_),
    .A(\top_ihp.wb_coproc.opb[2] ),
    .Y(_04336_));
 sg13g2_o21ai_1 _20620_ (.B1(_04336_),
    .Y(_04337_),
    .A1(_04333_),
    .A2(_04334_));
 sg13g2_mux2_1 _20621_ (.A0(\top_ihp.wb_coproc.dat_o[2] ),
    .A1(_04337_),
    .S(net217),
    .X(_02560_));
 sg13g2_inv_1 _20622_ (.Y(_04338_),
    .A(\top_ihp.wb_coproc.opa[30] ));
 sg13g2_mux2_1 _20623_ (.A0(net558),
    .A1(net557),
    .S(\top_ihp.wb_coproc.opb[30] ),
    .X(_04339_));
 sg13g2_nand2_1 _20624_ (.Y(_04340_),
    .A(\top_ihp.wb_coproc.opa[30] ),
    .B(_04323_));
 sg13g2_nand3_1 _20625_ (.B(_04322_),
    .C(_04340_),
    .A(\top_ihp.wb_coproc.opb[30] ),
    .Y(_04341_));
 sg13g2_o21ai_1 _20626_ (.B1(_04341_),
    .Y(_04342_),
    .A1(_04338_),
    .A2(_04339_));
 sg13g2_mux2_1 _20627_ (.A0(\top_ihp.wb_coproc.dat_o[30] ),
    .A1(_04342_),
    .S(_04327_),
    .X(_02561_));
 sg13g2_inv_1 _20628_ (.Y(_04343_),
    .A(\top_ihp.wb_coproc.opa[31] ));
 sg13g2_mux2_1 _20629_ (.A0(net558),
    .A1(net557),
    .S(\top_ihp.wb_coproc.opb[31] ),
    .X(_04344_));
 sg13g2_nand2_1 _20630_ (.Y(_04345_),
    .A(\top_ihp.wb_coproc.opa[31] ),
    .B(net738));
 sg13g2_nand3_1 _20631_ (.B(_04322_),
    .C(_04345_),
    .A(\top_ihp.wb_coproc.opb[31] ),
    .Y(_04346_));
 sg13g2_o21ai_1 _20632_ (.B1(_04346_),
    .Y(_04347_),
    .A1(_04343_),
    .A2(_04344_));
 sg13g2_mux2_1 _20633_ (.A0(\top_ihp.wb_coproc.dat_o[31] ),
    .A1(_04347_),
    .S(net217),
    .X(_02562_));
 sg13g2_inv_1 _20634_ (.Y(_04348_),
    .A(\top_ihp.wb_coproc.opa[3] ));
 sg13g2_mux2_1 _20635_ (.A0(net558),
    .A1(net557),
    .S(\top_ihp.wb_coproc.opb[3] ),
    .X(_04349_));
 sg13g2_nand2_1 _20636_ (.Y(_04350_),
    .A(\top_ihp.wb_coproc.opa[3] ),
    .B(net738));
 sg13g2_nand3_1 _20637_ (.B(net556),
    .C(_04350_),
    .A(\top_ihp.wb_coproc.opb[3] ),
    .Y(_04351_));
 sg13g2_o21ai_1 _20638_ (.B1(_04351_),
    .Y(_04352_),
    .A1(_04348_),
    .A2(_04349_));
 sg13g2_mux2_1 _20639_ (.A0(\top_ihp.wb_coproc.dat_o[3] ),
    .A1(_04352_),
    .S(net217),
    .X(_02563_));
 sg13g2_inv_1 _20640_ (.Y(_04353_),
    .A(\top_ihp.wb_coproc.opa[4] ));
 sg13g2_mux2_1 _20641_ (.A0(net558),
    .A1(net557),
    .S(\top_ihp.wb_coproc.opb[4] ),
    .X(_04354_));
 sg13g2_nand2_1 _20642_ (.Y(_04355_),
    .A(\top_ihp.wb_coproc.opa[4] ),
    .B(net738));
 sg13g2_nand3_1 _20643_ (.B(net556),
    .C(_04355_),
    .A(\top_ihp.wb_coproc.opb[4] ),
    .Y(_04356_));
 sg13g2_o21ai_1 _20644_ (.B1(_04356_),
    .Y(_04357_),
    .A1(_04353_),
    .A2(_04354_));
 sg13g2_mux2_1 _20645_ (.A0(\top_ihp.wb_coproc.dat_o[4] ),
    .A1(_04357_),
    .S(net217),
    .X(_02564_));
 sg13g2_inv_1 _20646_ (.Y(_04358_),
    .A(\top_ihp.wb_coproc.opa[5] ));
 sg13g2_mux2_1 _20647_ (.A0(net558),
    .A1(net557),
    .S(\top_ihp.wb_coproc.opb[5] ),
    .X(_04359_));
 sg13g2_nand2_1 _20648_ (.Y(_04360_),
    .A(\top_ihp.wb_coproc.opa[5] ),
    .B(net738));
 sg13g2_nand3_1 _20649_ (.B(net556),
    .C(_04360_),
    .A(\top_ihp.wb_coproc.opb[5] ),
    .Y(_04361_));
 sg13g2_o21ai_1 _20650_ (.B1(_04361_),
    .Y(_04362_),
    .A1(_04358_),
    .A2(_04359_));
 sg13g2_mux2_1 _20651_ (.A0(\top_ihp.wb_coproc.dat_o[5] ),
    .A1(_04362_),
    .S(net217),
    .X(_02565_));
 sg13g2_inv_1 _20652_ (.Y(_04363_),
    .A(\top_ihp.wb_coproc.opa[6] ));
 sg13g2_mux2_1 _20653_ (.A0(net558),
    .A1(net557),
    .S(\top_ihp.wb_coproc.opb[6] ),
    .X(_04364_));
 sg13g2_nand2_1 _20654_ (.Y(_04365_),
    .A(\top_ihp.wb_coproc.opa[6] ),
    .B(net738));
 sg13g2_nand3_1 _20655_ (.B(net556),
    .C(_04365_),
    .A(\top_ihp.wb_coproc.opb[6] ),
    .Y(_04366_));
 sg13g2_o21ai_1 _20656_ (.B1(_04366_),
    .Y(_04367_),
    .A1(_04363_),
    .A2(_04364_));
 sg13g2_mux2_1 _20657_ (.A0(\top_ihp.wb_coproc.dat_o[6] ),
    .A1(_04367_),
    .S(net217),
    .X(_02566_));
 sg13g2_inv_1 _20658_ (.Y(_04368_),
    .A(\top_ihp.wb_coproc.opa[7] ));
 sg13g2_mux2_1 _20659_ (.A0(net558),
    .A1(net557),
    .S(\top_ihp.wb_coproc.opb[7] ),
    .X(_04369_));
 sg13g2_nand2_1 _20660_ (.Y(_04370_),
    .A(\top_ihp.wb_coproc.opa[7] ),
    .B(net738));
 sg13g2_nand3_1 _20661_ (.B(net556),
    .C(_04370_),
    .A(\top_ihp.wb_coproc.opb[7] ),
    .Y(_04371_));
 sg13g2_o21ai_1 _20662_ (.B1(_04371_),
    .Y(_04372_),
    .A1(_04368_),
    .A2(_04369_));
 sg13g2_mux2_1 _20663_ (.A0(\top_ihp.wb_coproc.dat_o[7] ),
    .A1(_04372_),
    .S(net217),
    .X(_02567_));
 sg13g2_inv_1 _20664_ (.Y(_04373_),
    .A(\top_ihp.wb_coproc.opa[8] ));
 sg13g2_mux2_1 _20665_ (.A0(_04194_),
    .A1(_04204_),
    .S(\top_ihp.wb_coproc.opb[8] ),
    .X(_04374_));
 sg13g2_nand2_1 _20666_ (.Y(_04375_),
    .A(\top_ihp.wb_coproc.opa[8] ),
    .B(_04202_));
 sg13g2_nand3_1 _20667_ (.B(_04209_),
    .C(_04375_),
    .A(\top_ihp.wb_coproc.opb[8] ),
    .Y(_04376_));
 sg13g2_o21ai_1 _20668_ (.B1(_04376_),
    .Y(_04377_),
    .A1(_04373_),
    .A2(_04374_));
 sg13g2_mux2_1 _20669_ (.A0(\top_ihp.wb_coproc.dat_o[8] ),
    .A1(_04377_),
    .S(_04216_),
    .X(_02568_));
 sg13g2_inv_1 _20670_ (.Y(_04378_),
    .A(\top_ihp.wb_coproc.opa[9] ));
 sg13g2_mux2_1 _20671_ (.A0(_04194_),
    .A1(_04204_),
    .S(\top_ihp.wb_coproc.opb[9] ),
    .X(_04379_));
 sg13g2_nand2_1 _20672_ (.Y(_04380_),
    .A(\top_ihp.wb_coproc.opa[9] ),
    .B(_04202_));
 sg13g2_nand3_1 _20673_ (.B(_04209_),
    .C(_04380_),
    .A(\top_ihp.wb_coproc.opb[9] ),
    .Y(_04381_));
 sg13g2_o21ai_1 _20674_ (.B1(_04381_),
    .Y(_04382_),
    .A1(_04378_),
    .A2(_04379_));
 sg13g2_mux2_1 _20675_ (.A0(\top_ihp.wb_coproc.dat_o[9] ),
    .A1(_04382_),
    .S(_04216_),
    .X(_02569_));
 sg13g2_inv_1 _20676_ (.Y(_04383_),
    .A(_04202_));
 sg13g2_nor4_1 _20677_ (.A(net883),
    .B(_04197_),
    .C(_04188_),
    .D(_04207_),
    .Y(_04384_));
 sg13g2_nand3_1 _20678_ (.B(_04383_),
    .C(_04384_),
    .A(_00003_),
    .Y(_04385_));
 sg13g2_buf_2 _20679_ (.A(_04385_),
    .X(_04386_));
 sg13g2_buf_1 _20680_ (.A(_04386_),
    .X(_04387_));
 sg13g2_mux2_1 _20681_ (.A0(net1050),
    .A1(\top_ihp.wb_coproc.opa[0] ),
    .S(net216),
    .X(_02570_));
 sg13g2_mux2_1 _20682_ (.A0(_04113_),
    .A1(\top_ihp.wb_coproc.opa[10] ),
    .S(_04387_),
    .X(_02571_));
 sg13g2_mux2_1 _20683_ (.A0(_04115_),
    .A1(\top_ihp.wb_coproc.opa[11] ),
    .S(net216),
    .X(_02572_));
 sg13g2_mux2_1 _20684_ (.A0(_04117_),
    .A1(\top_ihp.wb_coproc.opa[12] ),
    .S(net216),
    .X(_02573_));
 sg13g2_mux2_1 _20685_ (.A0(_04119_),
    .A1(\top_ihp.wb_coproc.opa[13] ),
    .S(net216),
    .X(_02574_));
 sg13g2_mux2_1 _20686_ (.A0(_04121_),
    .A1(\top_ihp.wb_coproc.opa[14] ),
    .S(net216),
    .X(_02575_));
 sg13g2_mux2_1 _20687_ (.A0(_04124_),
    .A1(\top_ihp.wb_coproc.opa[15] ),
    .S(net216),
    .X(_02576_));
 sg13g2_mux2_1 _20688_ (.A0(_04126_),
    .A1(\top_ihp.wb_coproc.opa[16] ),
    .S(net216),
    .X(_02577_));
 sg13g2_mux2_1 _20689_ (.A0(_04128_),
    .A1(\top_ihp.wb_coproc.opa[17] ),
    .S(_04387_),
    .X(_02578_));
 sg13g2_mux2_1 _20690_ (.A0(_04130_),
    .A1(\top_ihp.wb_coproc.opa[18] ),
    .S(net216),
    .X(_02579_));
 sg13g2_buf_1 _20691_ (.A(_04386_),
    .X(_04388_));
 sg13g2_mux2_1 _20692_ (.A0(_04134_),
    .A1(\top_ihp.wb_coproc.opa[19] ),
    .S(net215),
    .X(_02580_));
 sg13g2_mux2_1 _20693_ (.A0(_04136_),
    .A1(\top_ihp.wb_coproc.opa[1] ),
    .S(net215),
    .X(_02581_));
 sg13g2_mux2_1 _20694_ (.A0(_04138_),
    .A1(\top_ihp.wb_coproc.opa[20] ),
    .S(net215),
    .X(_02582_));
 sg13g2_mux2_1 _20695_ (.A0(_04140_),
    .A1(\top_ihp.wb_coproc.opa[21] ),
    .S(net215),
    .X(_02583_));
 sg13g2_mux2_1 _20696_ (.A0(_04142_),
    .A1(\top_ihp.wb_coproc.opa[22] ),
    .S(net215),
    .X(_02584_));
 sg13g2_mux2_1 _20697_ (.A0(_04144_),
    .A1(\top_ihp.wb_coproc.opa[23] ),
    .S(net215),
    .X(_02585_));
 sg13g2_mux2_1 _20698_ (.A0(_04148_),
    .A1(\top_ihp.wb_coproc.opa[24] ),
    .S(net215),
    .X(_02586_));
 sg13g2_mux2_1 _20699_ (.A0(_04150_),
    .A1(\top_ihp.wb_coproc.opa[25] ),
    .S(_04388_),
    .X(_02587_));
 sg13g2_mux2_1 _20700_ (.A0(_04151_),
    .A1(\top_ihp.wb_coproc.opa[26] ),
    .S(net215),
    .X(_02588_));
 sg13g2_mux2_1 _20701_ (.A0(_04153_),
    .A1(\top_ihp.wb_coproc.opa[27] ),
    .S(_04388_),
    .X(_02589_));
 sg13g2_buf_8 _20702_ (.A(_04386_),
    .X(_04389_));
 sg13g2_mux2_1 _20703_ (.A0(_04155_),
    .A1(\top_ihp.wb_coproc.opa[28] ),
    .S(net214),
    .X(_02590_));
 sg13g2_mux2_1 _20704_ (.A0(_04156_),
    .A1(\top_ihp.wb_coproc.opa[29] ),
    .S(net214),
    .X(_02591_));
 sg13g2_mux2_1 _20705_ (.A0(_04158_),
    .A1(\top_ihp.wb_coproc.opa[2] ),
    .S(net214),
    .X(_02592_));
 sg13g2_mux2_1 _20706_ (.A0(_04160_),
    .A1(\top_ihp.wb_coproc.opa[30] ),
    .S(_04389_),
    .X(_02593_));
 sg13g2_mux2_1 _20707_ (.A0(_04162_),
    .A1(\top_ihp.wb_coproc.opa[31] ),
    .S(_04389_),
    .X(_02594_));
 sg13g2_mux2_1 _20708_ (.A0(_04163_),
    .A1(\top_ihp.wb_coproc.opa[3] ),
    .S(net214),
    .X(_02595_));
 sg13g2_mux2_1 _20709_ (.A0(_04165_),
    .A1(\top_ihp.wb_coproc.opa[4] ),
    .S(net214),
    .X(_02596_));
 sg13g2_mux2_1 _20710_ (.A0(_04167_),
    .A1(\top_ihp.wb_coproc.opa[5] ),
    .S(net214),
    .X(_02597_));
 sg13g2_mux2_1 _20711_ (.A0(_04169_),
    .A1(\top_ihp.wb_coproc.opa[6] ),
    .S(net214),
    .X(_02598_));
 sg13g2_mux2_1 _20712_ (.A0(_04171_),
    .A1(\top_ihp.wb_coproc.opa[7] ),
    .S(net214),
    .X(_02599_));
 sg13g2_mux2_1 _20713_ (.A0(_04173_),
    .A1(\top_ihp.wb_coproc.opa[8] ),
    .S(_04386_),
    .X(_02600_));
 sg13g2_mux2_1 _20714_ (.A0(_04175_),
    .A1(\top_ihp.wb_coproc.opa[9] ),
    .S(_04386_),
    .X(_02601_));
 sg13g2_nand3_1 _20715_ (.B(_04202_),
    .C(_04384_),
    .A(_00003_),
    .Y(_04390_));
 sg13g2_buf_8 _20716_ (.A(_04390_),
    .X(_04391_));
 sg13g2_buf_8 _20717_ (.A(_04391_),
    .X(_04392_));
 sg13g2_mux2_1 _20718_ (.A0(net1050),
    .A1(\top_ihp.wb_coproc.opb[0] ),
    .S(net213),
    .X(_02602_));
 sg13g2_mux2_1 _20719_ (.A0(_04113_),
    .A1(\top_ihp.wb_coproc.opb[10] ),
    .S(_04392_),
    .X(_02603_));
 sg13g2_mux2_1 _20720_ (.A0(_04115_),
    .A1(\top_ihp.wb_coproc.opb[11] ),
    .S(net213),
    .X(_02604_));
 sg13g2_mux2_1 _20721_ (.A0(_04117_),
    .A1(\top_ihp.wb_coproc.opb[12] ),
    .S(net213),
    .X(_02605_));
 sg13g2_mux2_1 _20722_ (.A0(_04119_),
    .A1(\top_ihp.wb_coproc.opb[13] ),
    .S(net213),
    .X(_02606_));
 sg13g2_mux2_1 _20723_ (.A0(_04121_),
    .A1(\top_ihp.wb_coproc.opb[14] ),
    .S(net213),
    .X(_02607_));
 sg13g2_mux2_1 _20724_ (.A0(_04124_),
    .A1(\top_ihp.wb_coproc.opb[15] ),
    .S(net213),
    .X(_02608_));
 sg13g2_mux2_1 _20725_ (.A0(_04126_),
    .A1(\top_ihp.wb_coproc.opb[16] ),
    .S(net213),
    .X(_02609_));
 sg13g2_mux2_1 _20726_ (.A0(_04128_),
    .A1(\top_ihp.wb_coproc.opb[17] ),
    .S(_04392_),
    .X(_02610_));
 sg13g2_mux2_1 _20727_ (.A0(_04130_),
    .A1(\top_ihp.wb_coproc.opb[18] ),
    .S(net213),
    .X(_02611_));
 sg13g2_buf_1 _20728_ (.A(_04391_),
    .X(_04393_));
 sg13g2_mux2_1 _20729_ (.A0(_04134_),
    .A1(\top_ihp.wb_coproc.opb[19] ),
    .S(net212),
    .X(_02612_));
 sg13g2_mux2_1 _20730_ (.A0(_04136_),
    .A1(\top_ihp.wb_coproc.opb[1] ),
    .S(net212),
    .X(_02613_));
 sg13g2_mux2_1 _20731_ (.A0(_04138_),
    .A1(\top_ihp.wb_coproc.opb[20] ),
    .S(net212),
    .X(_02614_));
 sg13g2_mux2_1 _20732_ (.A0(_04140_),
    .A1(\top_ihp.wb_coproc.opb[21] ),
    .S(net212),
    .X(_02615_));
 sg13g2_mux2_1 _20733_ (.A0(_04142_),
    .A1(\top_ihp.wb_coproc.opb[22] ),
    .S(net212),
    .X(_02616_));
 sg13g2_mux2_1 _20734_ (.A0(_04144_),
    .A1(\top_ihp.wb_coproc.opb[23] ),
    .S(net212),
    .X(_02617_));
 sg13g2_mux2_1 _20735_ (.A0(_04148_),
    .A1(\top_ihp.wb_coproc.opb[24] ),
    .S(_04393_),
    .X(_02618_));
 sg13g2_mux2_1 _20736_ (.A0(_04150_),
    .A1(\top_ihp.wb_coproc.opb[25] ),
    .S(net212),
    .X(_02619_));
 sg13g2_mux2_1 _20737_ (.A0(_04151_),
    .A1(\top_ihp.wb_coproc.opb[26] ),
    .S(net212),
    .X(_02620_));
 sg13g2_mux2_1 _20738_ (.A0(_04153_),
    .A1(\top_ihp.wb_coproc.opb[27] ),
    .S(_04393_),
    .X(_02621_));
 sg13g2_buf_8 _20739_ (.A(_04391_),
    .X(_04394_));
 sg13g2_mux2_1 _20740_ (.A0(_04155_),
    .A1(\top_ihp.wb_coproc.opb[28] ),
    .S(net211),
    .X(_02622_));
 sg13g2_mux2_1 _20741_ (.A0(_04156_),
    .A1(\top_ihp.wb_coproc.opb[29] ),
    .S(net211),
    .X(_02623_));
 sg13g2_mux2_1 _20742_ (.A0(_04158_),
    .A1(\top_ihp.wb_coproc.opb[2] ),
    .S(net211),
    .X(_02624_));
 sg13g2_mux2_1 _20743_ (.A0(_04160_),
    .A1(\top_ihp.wb_coproc.opb[30] ),
    .S(net211),
    .X(_02625_));
 sg13g2_mux2_1 _20744_ (.A0(_04162_),
    .A1(\top_ihp.wb_coproc.opb[31] ),
    .S(net211),
    .X(_02626_));
 sg13g2_mux2_1 _20745_ (.A0(_04163_),
    .A1(\top_ihp.wb_coproc.opb[3] ),
    .S(net211),
    .X(_02627_));
 sg13g2_mux2_1 _20746_ (.A0(_04165_),
    .A1(\top_ihp.wb_coproc.opb[4] ),
    .S(net211),
    .X(_02628_));
 sg13g2_mux2_1 _20747_ (.A0(_04167_),
    .A1(\top_ihp.wb_coproc.opb[5] ),
    .S(_04394_),
    .X(_02629_));
 sg13g2_mux2_1 _20748_ (.A0(_04169_),
    .A1(\top_ihp.wb_coproc.opb[6] ),
    .S(net211),
    .X(_02630_));
 sg13g2_mux2_1 _20749_ (.A0(_04171_),
    .A1(\top_ihp.wb_coproc.opb[7] ),
    .S(_04394_),
    .X(_02631_));
 sg13g2_mux2_1 _20750_ (.A0(_04173_),
    .A1(\top_ihp.wb_coproc.opb[8] ),
    .S(_04391_),
    .X(_02632_));
 sg13g2_mux2_1 _20751_ (.A0(_04175_),
    .A1(\top_ihp.wb_coproc.opb[9] ),
    .S(_04391_),
    .X(_02633_));
 sg13g2_inv_1 _20752_ (.Y(_04395_),
    .A(_00232_));
 sg13g2_buf_1 _20753_ (.A(_08775_),
    .X(_04396_));
 sg13g2_nand2_2 _20754_ (.Y(_04397_),
    .A(_08774_),
    .B(_04396_));
 sg13g2_nand2_1 _20755_ (.Y(_04398_),
    .A(_08778_),
    .B(_08779_));
 sg13g2_nand2b_1 _20756_ (.Y(_04399_),
    .B(_04398_),
    .A_N(_04397_));
 sg13g2_buf_1 _20757_ (.A(_04399_),
    .X(_04400_));
 sg13g2_buf_1 _20758_ (.A(\top_ihp.wb_emem.bit_counter[0] ),
    .X(_04401_));
 sg13g2_inv_1 _20759_ (.Y(_04402_),
    .A(_08774_));
 sg13g2_inv_1 _20760_ (.Y(_04403_),
    .A(_08775_));
 sg13g2_nand2_1 _20761_ (.Y(_04404_),
    .A(net982),
    .B(_04403_));
 sg13g2_buf_1 _20762_ (.A(_04404_),
    .X(_04405_));
 sg13g2_nand3_1 _20763_ (.B(_04405_),
    .C(net897),
    .A(_04401_),
    .Y(_04406_));
 sg13g2_o21ai_1 _20764_ (.B1(_04406_),
    .Y(_02634_),
    .A1(_04395_),
    .A2(net897));
 sg13g2_buf_1 _20765_ (.A(\top_ihp.wb_emem.bit_counter[1] ),
    .X(_04407_));
 sg13g2_nor2_2 _20766_ (.A(net913),
    .B(_04397_),
    .Y(_04408_));
 sg13g2_nand2_1 _20767_ (.Y(_04409_),
    .A(_04401_),
    .B(_04408_));
 sg13g2_nor2_1 _20768_ (.A(net914),
    .B(_04408_),
    .Y(_04410_));
 sg13g2_buf_1 _20769_ (.A(_04410_),
    .X(_04411_));
 sg13g2_nor2_1 _20770_ (.A(_04401_),
    .B(net897),
    .Y(_04412_));
 sg13g2_o21ai_1 _20771_ (.B1(_04407_),
    .Y(_04413_),
    .A1(_04411_),
    .A2(_04412_));
 sg13g2_o21ai_1 _20772_ (.B1(_04413_),
    .Y(_02635_),
    .A1(_04407_),
    .A2(_04409_));
 sg13g2_nand2_1 _20773_ (.Y(_04414_),
    .A(_04407_),
    .B(_04401_));
 sg13g2_xor2_1 _20774_ (.B(_04414_),
    .A(\top_ihp.wb_emem.bit_counter[2] ),
    .X(_04415_));
 sg13g2_nand3_1 _20775_ (.B(_04405_),
    .C(net897),
    .A(\top_ihp.wb_emem.bit_counter[2] ),
    .Y(_04416_));
 sg13g2_o21ai_1 _20776_ (.B1(_04416_),
    .Y(_02636_),
    .A1(net897),
    .A2(_04415_));
 sg13g2_buf_1 _20777_ (.A(\top_ihp.wb_emem.bit_counter[3] ),
    .X(_04417_));
 sg13g2_and3_1 _20778_ (.X(_04418_),
    .A(_04407_),
    .B(_04401_),
    .C(\top_ihp.wb_emem.bit_counter[2] ));
 sg13g2_buf_1 _20779_ (.A(_04418_),
    .X(_04419_));
 sg13g2_nand2_1 _20780_ (.Y(_04420_),
    .A(_04408_),
    .B(_04419_));
 sg13g2_nor2_1 _20781_ (.A(net897),
    .B(_04419_),
    .Y(_04421_));
 sg13g2_o21ai_1 _20782_ (.B1(_04417_),
    .Y(_04422_),
    .A1(_04411_),
    .A2(_04421_));
 sg13g2_o21ai_1 _20783_ (.B1(_04422_),
    .Y(_02637_),
    .A1(_04417_),
    .A2(_04420_));
 sg13g2_buf_1 _20784_ (.A(\top_ihp.wb_emem.bit_counter[4] ),
    .X(_04423_));
 sg13g2_nand2b_1 _20785_ (.Y(_04424_),
    .B(_04417_),
    .A_N(_04423_));
 sg13g2_a21oi_1 _20786_ (.A1(_04417_),
    .A2(_04419_),
    .Y(_04425_),
    .B1(net897));
 sg13g2_o21ai_1 _20787_ (.B1(_04423_),
    .Y(_04426_),
    .A1(_04411_),
    .A2(_04425_));
 sg13g2_o21ai_1 _20788_ (.B1(_04426_),
    .Y(_02638_),
    .A1(_04420_),
    .A2(_04424_));
 sg13g2_buf_1 _20789_ (.A(\top_ihp.wb_emem.bit_counter[5] ),
    .X(_04427_));
 sg13g2_and3_1 _20790_ (.X(_04428_),
    .A(_04417_),
    .B(_04423_),
    .C(_04419_));
 sg13g2_buf_1 _20791_ (.A(_04428_),
    .X(_04429_));
 sg13g2_nand2_1 _20792_ (.Y(_04430_),
    .A(_04408_),
    .B(_04429_));
 sg13g2_nor2_1 _20793_ (.A(net897),
    .B(_04429_),
    .Y(_04431_));
 sg13g2_o21ai_1 _20794_ (.B1(_04427_),
    .Y(_04432_),
    .A1(_04411_),
    .A2(_04431_));
 sg13g2_o21ai_1 _20795_ (.B1(_04432_),
    .Y(_02639_),
    .A1(_04427_),
    .A2(_04430_));
 sg13g2_nand3_1 _20796_ (.B(_04408_),
    .C(_04429_),
    .A(_04427_),
    .Y(_04433_));
 sg13g2_a21oi_1 _20797_ (.A1(_04427_),
    .A2(_04429_),
    .Y(_04434_),
    .B1(_04400_));
 sg13g2_o21ai_1 _20798_ (.B1(\top_ihp.wb_emem.bit_counter[6] ),
    .Y(_04435_),
    .A1(_04411_),
    .A2(_04434_));
 sg13g2_o21ai_1 _20799_ (.B1(_04435_),
    .Y(_02640_),
    .A1(\top_ihp.wb_emem.bit_counter[6] ),
    .A2(_04433_));
 sg13g2_nand2_1 _20800_ (.Y(_04436_),
    .A(\top_ihp.wb_emem.bit_counter[7] ),
    .B(_04405_));
 sg13g2_inv_1 _20801_ (.Y(_04437_),
    .A(\top_ihp.wb_emem.bit_counter[6] ));
 sg13g2_or2_1 _20802_ (.X(_04438_),
    .B(_04433_),
    .A(_04437_));
 sg13g2_mux2_1 _20803_ (.A0(\top_ihp.wb_emem.bit_counter[7] ),
    .A1(_04436_),
    .S(_04438_),
    .X(_04439_));
 sg13g2_inv_1 _20804_ (.Y(_02641_),
    .A(_04439_));
 sg13g2_a21oi_1 _20805_ (.A1(_04403_),
    .A2(net913),
    .Y(_04440_),
    .B1(_08774_));
 sg13g2_buf_1 _20806_ (.A(_04440_),
    .X(_04441_));
 sg13g2_buf_1 _20807_ (.A(_04441_),
    .X(_04442_));
 sg13g2_buf_1 _20808_ (.A(net876),
    .X(_04443_));
 sg13g2_nand2_1 _20809_ (.Y(_04444_),
    .A(_09869_),
    .B(net913));
 sg13g2_buf_1 _20810_ (.A(_04444_),
    .X(_04445_));
 sg13g2_buf_1 _20811_ (.A(_04445_),
    .X(_04446_));
 sg13g2_nand2_1 _20812_ (.Y(_04447_),
    .A(net4),
    .B(_04446_));
 sg13g2_nor2_1 _20813_ (.A(_04405_),
    .B(_04398_),
    .Y(_04448_));
 sg13g2_buf_1 _20814_ (.A(_04448_),
    .X(_04449_));
 sg13g2_buf_1 _20815_ (.A(_04449_),
    .X(_04450_));
 sg13g2_nand3_1 _20816_ (.B(net837),
    .C(net874),
    .A(_04148_),
    .Y(_04451_));
 sg13g2_buf_1 _20817_ (.A(_04441_),
    .X(_04452_));
 sg13g2_a21oi_1 _20818_ (.A1(_04447_),
    .A2(_04451_),
    .Y(_04453_),
    .B1(net873));
 sg13g2_a21o_1 _20819_ (.A2(net853),
    .A1(\top_ihp.wb_dati_ram[24] ),
    .B1(_04453_),
    .X(_02642_));
 sg13g2_nand2_1 _20820_ (.Y(_04454_),
    .A(\top_ihp.wb_dati_ram[17] ),
    .B(net875));
 sg13g2_buf_1 _20821_ (.A(_04449_),
    .X(_04455_));
 sg13g2_nand3_1 _20822_ (.B(_07978_),
    .C(net872),
    .A(_04130_),
    .Y(_04456_));
 sg13g2_a21oi_1 _20823_ (.A1(_04454_),
    .A2(_04456_),
    .Y(_04457_),
    .B1(net873));
 sg13g2_a21o_1 _20824_ (.A2(net853),
    .A1(\top_ihp.wb_dati_ram[18] ),
    .B1(_04457_),
    .X(_02643_));
 sg13g2_nand2_1 _20825_ (.Y(_04458_),
    .A(\top_ihp.wb_dati_ram[18] ),
    .B(net875));
 sg13g2_buf_1 _20826_ (.A(_07977_),
    .X(_04459_));
 sg13g2_nand3_1 _20827_ (.B(net834),
    .C(net872),
    .A(_04134_),
    .Y(_04460_));
 sg13g2_a21oi_1 _20828_ (.A1(_04458_),
    .A2(_04460_),
    .Y(_04461_),
    .B1(net873));
 sg13g2_a21o_1 _20829_ (.A2(net853),
    .A1(\top_ihp.wb_dati_ram[19] ),
    .B1(_04461_),
    .X(_02644_));
 sg13g2_nand2_1 _20830_ (.Y(_04462_),
    .A(\top_ihp.wb_dati_ram[19] ),
    .B(net875));
 sg13g2_nand3_1 _20831_ (.B(net834),
    .C(net872),
    .A(_04138_),
    .Y(_04463_));
 sg13g2_a21oi_1 _20832_ (.A1(_04462_),
    .A2(_04463_),
    .Y(_04464_),
    .B1(net873));
 sg13g2_a21o_1 _20833_ (.A2(net853),
    .A1(\top_ihp.wb_dati_ram[20] ),
    .B1(_04464_),
    .X(_02645_));
 sg13g2_nand2_1 _20834_ (.Y(_04465_),
    .A(\top_ihp.wb_dati_ram[20] ),
    .B(_04446_));
 sg13g2_nand3_1 _20835_ (.B(net834),
    .C(net872),
    .A(_04140_),
    .Y(_04466_));
 sg13g2_a21oi_1 _20836_ (.A1(_04465_),
    .A2(_04466_),
    .Y(_04467_),
    .B1(net873));
 sg13g2_a21o_1 _20837_ (.A2(_04443_),
    .A1(\top_ihp.wb_dati_ram[21] ),
    .B1(_04467_),
    .X(_02646_));
 sg13g2_buf_1 _20838_ (.A(_04445_),
    .X(_04468_));
 sg13g2_buf_1 _20839_ (.A(net871),
    .X(_04469_));
 sg13g2_nand2_1 _20840_ (.Y(_04470_),
    .A(\top_ihp.wb_dati_ram[21] ),
    .B(net852));
 sg13g2_nand3_1 _20841_ (.B(net834),
    .C(net872),
    .A(_04142_),
    .Y(_04471_));
 sg13g2_a21oi_1 _20842_ (.A1(_04470_),
    .A2(_04471_),
    .Y(_04472_),
    .B1(net873));
 sg13g2_a21o_1 _20843_ (.A2(_04443_),
    .A1(\top_ihp.wb_dati_ram[22] ),
    .B1(_04472_),
    .X(_02647_));
 sg13g2_buf_1 _20844_ (.A(net876),
    .X(_04473_));
 sg13g2_nand2_1 _20845_ (.Y(_04474_),
    .A(\top_ihp.wb_dati_ram[22] ),
    .B(net852));
 sg13g2_nand3_1 _20846_ (.B(net834),
    .C(net872),
    .A(_04144_),
    .Y(_04475_));
 sg13g2_a21oi_1 _20847_ (.A1(_04474_),
    .A2(_04475_),
    .Y(_04476_),
    .B1(net873));
 sg13g2_a21o_1 _20848_ (.A2(net851),
    .A1(\top_ihp.wb_dati_ram[23] ),
    .B1(_04476_),
    .X(_02648_));
 sg13g2_nand2_1 _20849_ (.Y(_04477_),
    .A(\top_ihp.wb_dati_ram[23] ),
    .B(net852));
 sg13g2_nand3_1 _20850_ (.B(_04459_),
    .C(_04455_),
    .A(_04173_),
    .Y(_04478_));
 sg13g2_a21oi_1 _20851_ (.A1(_04477_),
    .A2(_04478_),
    .Y(_04479_),
    .B1(_04452_));
 sg13g2_a21o_1 _20852_ (.A2(net851),
    .A1(\top_ihp.wb_dati_ram[8] ),
    .B1(_04479_),
    .X(_02649_));
 sg13g2_nand2_1 _20853_ (.Y(_04480_),
    .A(\top_ihp.wb_dati_ram[8] ),
    .B(_04469_));
 sg13g2_nand3_1 _20854_ (.B(_04459_),
    .C(_04455_),
    .A(_04175_),
    .Y(_04481_));
 sg13g2_a21oi_1 _20855_ (.A1(_04480_),
    .A2(_04481_),
    .Y(_04482_),
    .B1(_04452_));
 sg13g2_a21o_1 _20856_ (.A2(net851),
    .A1(\top_ihp.wb_dati_ram[9] ),
    .B1(_04482_),
    .X(_02650_));
 sg13g2_nand2_1 _20857_ (.Y(_04483_),
    .A(\top_ihp.wb_dati_ram[9] ),
    .B(_04469_));
 sg13g2_nand3_1 _20858_ (.B(net834),
    .C(net872),
    .A(_04113_),
    .Y(_04484_));
 sg13g2_a21oi_1 _20859_ (.A1(_04483_),
    .A2(_04484_),
    .Y(_04485_),
    .B1(net873));
 sg13g2_a21o_1 _20860_ (.A2(_04473_),
    .A1(\top_ihp.wb_dati_ram[10] ),
    .B1(_04485_),
    .X(_02651_));
 sg13g2_nand2_1 _20861_ (.Y(_04486_),
    .A(\top_ihp.wb_dati_ram[10] ),
    .B(net852));
 sg13g2_nand3_1 _20862_ (.B(net834),
    .C(net872),
    .A(_04115_),
    .Y(_04487_));
 sg13g2_buf_1 _20863_ (.A(_04441_),
    .X(_04488_));
 sg13g2_a21oi_1 _20864_ (.A1(_04486_),
    .A2(_04487_),
    .Y(_04489_),
    .B1(net870));
 sg13g2_a21o_1 _20865_ (.A2(net851),
    .A1(\top_ihp.wb_dati_ram[11] ),
    .B1(_04489_),
    .X(_02652_));
 sg13g2_nand2_1 _20866_ (.Y(_04490_),
    .A(\top_ihp.wb_dati_ram[24] ),
    .B(net852));
 sg13g2_buf_1 _20867_ (.A(_04449_),
    .X(_04491_));
 sg13g2_nand3_1 _20868_ (.B(net834),
    .C(net869),
    .A(_04150_),
    .Y(_04492_));
 sg13g2_a21oi_1 _20869_ (.A1(_04490_),
    .A2(_04492_),
    .Y(_04493_),
    .B1(net870));
 sg13g2_a21o_1 _20870_ (.A2(net851),
    .A1(\top_ihp.wb_dati_ram[25] ),
    .B1(_04493_),
    .X(_02653_));
 sg13g2_nand2_1 _20871_ (.Y(_04494_),
    .A(\top_ihp.wb_dati_ram[11] ),
    .B(net852));
 sg13g2_buf_1 _20872_ (.A(net857),
    .X(_04495_));
 sg13g2_nand3_1 _20873_ (.B(net833),
    .C(_04491_),
    .A(_04117_),
    .Y(_04496_));
 sg13g2_a21oi_1 _20874_ (.A1(_04494_),
    .A2(_04496_),
    .Y(_04497_),
    .B1(net870));
 sg13g2_a21o_1 _20875_ (.A2(net851),
    .A1(\top_ihp.wb_dati_ram[12] ),
    .B1(_04497_),
    .X(_02654_));
 sg13g2_nand2_1 _20876_ (.Y(_04498_),
    .A(\top_ihp.wb_dati_ram[12] ),
    .B(net852));
 sg13g2_nand3_1 _20877_ (.B(net833),
    .C(net869),
    .A(_04119_),
    .Y(_04499_));
 sg13g2_a21oi_1 _20878_ (.A1(_04498_),
    .A2(_04499_),
    .Y(_04500_),
    .B1(_04488_));
 sg13g2_a21o_1 _20879_ (.A2(net851),
    .A1(\top_ihp.wb_dati_ram[13] ),
    .B1(_04500_),
    .X(_02655_));
 sg13g2_nand2_1 _20880_ (.Y(_04501_),
    .A(\top_ihp.wb_dati_ram[13] ),
    .B(net852));
 sg13g2_nand3_1 _20881_ (.B(net833),
    .C(net869),
    .A(_04121_),
    .Y(_04502_));
 sg13g2_a21oi_1 _20882_ (.A1(_04501_),
    .A2(_04502_),
    .Y(_04503_),
    .B1(net870));
 sg13g2_a21o_1 _20883_ (.A2(net851),
    .A1(\top_ihp.wb_dati_ram[14] ),
    .B1(_04503_),
    .X(_02656_));
 sg13g2_buf_1 _20884_ (.A(net871),
    .X(_04504_));
 sg13g2_nand2_1 _20885_ (.Y(_04505_),
    .A(\top_ihp.wb_dati_ram[14] ),
    .B(net850));
 sg13g2_nand3_1 _20886_ (.B(_04495_),
    .C(_04491_),
    .A(_04124_),
    .Y(_04506_));
 sg13g2_a21oi_1 _20887_ (.A1(_04505_),
    .A2(_04506_),
    .Y(_04507_),
    .B1(_04488_));
 sg13g2_a21o_1 _20888_ (.A2(_04473_),
    .A1(\top_ihp.wb_dati_ram[15] ),
    .B1(_04507_),
    .X(_02657_));
 sg13g2_buf_1 _20889_ (.A(_04468_),
    .X(_04508_));
 sg13g2_and2_1 _20890_ (.A(net1050),
    .B(_04449_),
    .X(_04509_));
 sg13g2_buf_1 _20891_ (.A(_04441_),
    .X(_04510_));
 sg13g2_a221oi_1 _20892_ (.B2(net837),
    .C1(net868),
    .B1(_04509_),
    .A1(\top_ihp.wb_dati_ram[15] ),
    .Y(_04511_),
    .A2(net849));
 sg13g2_a21oi_1 _20893_ (.A1(_09662_),
    .A2(net853),
    .Y(_02658_),
    .B1(_04511_));
 sg13g2_nand3_1 _20894_ (.B(_07978_),
    .C(net874),
    .A(_04136_),
    .Y(_04512_));
 sg13g2_o21ai_1 _20895_ (.B1(_04512_),
    .Y(_04513_),
    .A1(_09662_),
    .A2(net874));
 sg13g2_o21ai_1 _20896_ (.B1(net982),
    .Y(_04514_),
    .A1(net983),
    .A2(_04398_));
 sg13g2_buf_1 _20897_ (.A(_04514_),
    .X(_04515_));
 sg13g2_mux2_1 _20898_ (.A0(\top_ihp.wb_dati_ram[1] ),
    .A1(_04513_),
    .S(_04515_),
    .X(_02659_));
 sg13g2_buf_1 _20899_ (.A(_04442_),
    .X(_04516_));
 sg13g2_nand2_1 _20900_ (.Y(_04517_),
    .A(\top_ihp.wb_dati_ram[1] ),
    .B(net850));
 sg13g2_nand3_1 _20901_ (.B(net833),
    .C(net869),
    .A(_04158_),
    .Y(_04518_));
 sg13g2_a21oi_1 _20902_ (.A1(_04517_),
    .A2(_04518_),
    .Y(_04519_),
    .B1(net870));
 sg13g2_a21o_1 _20903_ (.A2(net848),
    .A1(\top_ihp.wb_dati_ram[2] ),
    .B1(_04519_),
    .X(_02660_));
 sg13g2_nand2_1 _20904_ (.Y(_04520_),
    .A(\top_ihp.wb_dati_ram[2] ),
    .B(net850));
 sg13g2_nand3_1 _20905_ (.B(net833),
    .C(net869),
    .A(_04163_),
    .Y(_04521_));
 sg13g2_a21oi_1 _20906_ (.A1(_04520_),
    .A2(_04521_),
    .Y(_04522_),
    .B1(net870));
 sg13g2_a21o_1 _20907_ (.A2(net848),
    .A1(\top_ihp.wb_dati_ram[3] ),
    .B1(_04522_),
    .X(_02661_));
 sg13g2_nand2_1 _20908_ (.Y(_04523_),
    .A(\top_ihp.wb_dati_ram[3] ),
    .B(net850));
 sg13g2_nand3_1 _20909_ (.B(net833),
    .C(net869),
    .A(_04165_),
    .Y(_04524_));
 sg13g2_a21oi_1 _20910_ (.A1(_04523_),
    .A2(_04524_),
    .Y(_04525_),
    .B1(net870));
 sg13g2_a21o_1 _20911_ (.A2(net848),
    .A1(\top_ihp.wb_dati_ram[4] ),
    .B1(_04525_),
    .X(_02662_));
 sg13g2_nand2_1 _20912_ (.Y(_04526_),
    .A(\top_ihp.wb_dati_ram[4] ),
    .B(net850));
 sg13g2_nand3_1 _20913_ (.B(net833),
    .C(net869),
    .A(_04167_),
    .Y(_04527_));
 sg13g2_a21oi_1 _20914_ (.A1(_04526_),
    .A2(_04527_),
    .Y(_04528_),
    .B1(net870));
 sg13g2_a21o_1 _20915_ (.A2(net848),
    .A1(\top_ihp.wb_dati_ram[5] ),
    .B1(_04528_),
    .X(_02663_));
 sg13g2_nand2_1 _20916_ (.Y(_04529_),
    .A(\top_ihp.wb_dati_ram[25] ),
    .B(net850));
 sg13g2_nand3_1 _20917_ (.B(_04495_),
    .C(net869),
    .A(_04151_),
    .Y(_04530_));
 sg13g2_buf_1 _20918_ (.A(_04441_),
    .X(_04531_));
 sg13g2_a21oi_1 _20919_ (.A1(_04529_),
    .A2(_04530_),
    .Y(_04532_),
    .B1(net867));
 sg13g2_a21o_1 _20920_ (.A2(net848),
    .A1(\top_ihp.wb_dati_ram[26] ),
    .B1(_04532_),
    .X(_02664_));
 sg13g2_nand2_1 _20921_ (.Y(_04533_),
    .A(\top_ihp.wb_dati_ram[5] ),
    .B(net850));
 sg13g2_buf_1 _20922_ (.A(_04449_),
    .X(_04534_));
 sg13g2_nand3_1 _20923_ (.B(net833),
    .C(net866),
    .A(_04169_),
    .Y(_04535_));
 sg13g2_a21oi_1 _20924_ (.A1(_04533_),
    .A2(_04535_),
    .Y(_04536_),
    .B1(net867));
 sg13g2_a21o_1 _20925_ (.A2(net848),
    .A1(\top_ihp.wb_dati_ram[6] ),
    .B1(_04536_),
    .X(_02665_));
 sg13g2_nand2_1 _20926_ (.Y(_04537_),
    .A(\top_ihp.wb_dati_ram[6] ),
    .B(net850));
 sg13g2_nand3_1 _20927_ (.B(_08640_),
    .C(net866),
    .A(_04171_),
    .Y(_04538_));
 sg13g2_a21oi_1 _20928_ (.A1(_04537_),
    .A2(_04538_),
    .Y(_04539_),
    .B1(_04531_));
 sg13g2_a21o_1 _20929_ (.A2(net848),
    .A1(\top_ihp.wb_dati_ram[7] ),
    .B1(_04539_),
    .X(_02666_));
 sg13g2_and2_1 _20930_ (.A(\top_ihp.oisc.wb_adr_o[0] ),
    .B(net866),
    .X(_04540_));
 sg13g2_a21oi_1 _20931_ (.A1(\top_ihp.wb_dati_ram[7] ),
    .A2(net849),
    .Y(_04541_),
    .B1(_04540_));
 sg13g2_buf_1 _20932_ (.A(_04441_),
    .X(_04542_));
 sg13g2_nand2_1 _20933_ (.Y(_04543_),
    .A(\top_ihp.wb_emem.cmd[32] ),
    .B(net865));
 sg13g2_o21ai_1 _20934_ (.B1(_04543_),
    .Y(_02667_),
    .A1(net853),
    .A2(_04541_));
 sg13g2_nor2_1 _20935_ (.A(_08457_),
    .B(net875),
    .Y(_04544_));
 sg13g2_a21oi_1 _20936_ (.A1(\top_ihp.wb_emem.cmd[32] ),
    .A2(net849),
    .Y(_04545_),
    .B1(_04544_));
 sg13g2_nand2_1 _20937_ (.Y(_04546_),
    .A(\top_ihp.wb_emem.cmd[33] ),
    .B(net865));
 sg13g2_o21ai_1 _20938_ (.B1(_04546_),
    .Y(_02668_),
    .A1(net853),
    .A2(_04545_));
 sg13g2_nor2_1 _20939_ (.A(net875),
    .B(_04383_),
    .Y(_04547_));
 sg13g2_a21oi_1 _20940_ (.A1(\top_ihp.wb_emem.cmd[33] ),
    .A2(net849),
    .Y(_04548_),
    .B1(_04547_));
 sg13g2_nand2_1 _20941_ (.Y(_04549_),
    .A(\top_ihp.wb_emem.cmd[34] ),
    .B(net865));
 sg13g2_o21ai_1 _20942_ (.B1(_04549_),
    .Y(_02669_),
    .A1(net853),
    .A2(_04548_));
 sg13g2_inv_1 _20943_ (.Y(_04550_),
    .A(\top_ihp.wb_emem.cmd[35] ));
 sg13g2_nand2_1 _20944_ (.Y(_04551_),
    .A(\top_ihp.wb_emem.cmd[34] ),
    .B(_04468_));
 sg13g2_o21ai_1 _20945_ (.B1(_04551_),
    .Y(_04552_),
    .A1(net875),
    .A2(_04183_));
 sg13g2_nand2_1 _20946_ (.Y(_04553_),
    .A(_04515_),
    .B(_04552_));
 sg13g2_o21ai_1 _20947_ (.B1(_04553_),
    .Y(_02670_),
    .A1(_04550_),
    .A2(_04515_));
 sg13g2_a221oi_1 _20948_ (.B2(net982),
    .C1(net876),
    .B1(_04187_),
    .A1(_04550_),
    .Y(_04554_),
    .A2(net849));
 sg13g2_a21o_1 _20949_ (.A2(_04516_),
    .A1(\top_ihp.wb_emem.cmd[36] ),
    .B1(_04554_),
    .X(_02671_));
 sg13g2_inv_1 _20950_ (.Y(_04555_),
    .A(\top_ihp.wb_emem.cmd[36] ));
 sg13g2_a21o_1 _20951_ (.A2(_10416_),
    .A1(_08214_),
    .B1(_07986_),
    .X(_04556_));
 sg13g2_nor3_1 _20952_ (.A(_08126_),
    .B(_08224_),
    .C(_10416_),
    .Y(_04557_));
 sg13g2_a21oi_2 _20953_ (.B1(_04557_),
    .Y(_04558_),
    .A2(_04556_),
    .A1(_08126_));
 sg13g2_a221oi_1 _20954_ (.B2(net982),
    .C1(_04442_),
    .B1(_04558_),
    .A1(_04555_),
    .Y(_04559_),
    .A2(net875));
 sg13g2_a21o_1 _20955_ (.A2(_04516_),
    .A1(\top_ihp.wb_emem.cmd[37] ),
    .B1(_04559_),
    .X(_02672_));
 sg13g2_nand2_1 _20956_ (.Y(_04560_),
    .A(_08214_),
    .B(_10446_));
 sg13g2_o21ai_1 _20957_ (.B1(_08310_),
    .Y(_04561_),
    .A1(net808),
    .A2(_10446_));
 sg13g2_nand2_1 _20958_ (.Y(_04562_),
    .A(net1045),
    .B(_04561_));
 sg13g2_o21ai_1 _20959_ (.B1(_04562_),
    .Y(_04563_),
    .A1(net1045),
    .A2(_04560_));
 sg13g2_nand2_1 _20960_ (.Y(_04564_),
    .A(net874),
    .B(_04563_));
 sg13g2_buf_1 _20961_ (.A(_08774_),
    .X(_04565_));
 sg13g2_buf_1 _20962_ (.A(net981),
    .X(_04566_));
 sg13g2_a22oi_1 _20963_ (.Y(_04567_),
    .B1(\top_ihp.wb_emem.cmd[38] ),
    .B2(net865),
    .A2(\top_ihp.wb_emem.cmd[37] ),
    .A1(net943));
 sg13g2_nand2_1 _20964_ (.Y(_02673_),
    .A(_04564_),
    .B(_04567_));
 sg13g2_buf_1 _20965_ (.A(net849),
    .X(_04568_));
 sg13g2_buf_1 _20966_ (.A(_08213_),
    .X(_04569_));
 sg13g2_a22oi_1 _20967_ (.Y(_04570_),
    .B1(_04569_),
    .B2(_10477_),
    .A2(_08116_),
    .A1(_07987_));
 sg13g2_a22oi_1 _20968_ (.Y(_04571_),
    .B1(\top_ihp.wb_emem.cmd[39] ),
    .B2(net865),
    .A2(\top_ihp.wb_emem.cmd[38] ),
    .A1(net943));
 sg13g2_o21ai_1 _20969_ (.B1(_04571_),
    .Y(_02674_),
    .A1(net832),
    .A2(_04570_));
 sg13g2_nand2_1 _20970_ (.Y(_04572_),
    .A(\top_ihp.wb_dati_ram[26] ),
    .B(_04504_));
 sg13g2_nand3_1 _20971_ (.B(net836),
    .C(net866),
    .A(_04153_),
    .Y(_04573_));
 sg13g2_a21oi_1 _20972_ (.A1(_04572_),
    .A2(_04573_),
    .Y(_04574_),
    .B1(_04531_));
 sg13g2_a21o_1 _20973_ (.A2(net848),
    .A1(\top_ihp.wb_dati_ram[27] ),
    .B1(_04574_),
    .X(_02675_));
 sg13g2_a21o_1 _20974_ (.A2(_10491_),
    .A1(_04569_),
    .B1(net939),
    .X(_04575_));
 sg13g2_buf_1 _20975_ (.A(_08224_),
    .X(_04576_));
 sg13g2_nor3_1 _20976_ (.A(_08100_),
    .B(_04576_),
    .C(_10491_),
    .Y(_04577_));
 sg13g2_a21oi_1 _20977_ (.A1(_08100_),
    .A2(_04575_),
    .Y(_04578_),
    .B1(_04577_));
 sg13g2_a22oi_1 _20978_ (.Y(_04579_),
    .B1(\top_ihp.wb_emem.cmd[40] ),
    .B2(net865),
    .A2(\top_ihp.wb_emem.cmd[39] ),
    .A1(_04566_));
 sg13g2_o21ai_1 _20979_ (.B1(_04579_),
    .Y(_02676_),
    .A1(net832),
    .A2(_04578_));
 sg13g2_a21o_1 _20980_ (.A2(_10507_),
    .A1(net781),
    .B1(net939),
    .X(_04580_));
 sg13g2_nor3_1 _20981_ (.A(_08103_),
    .B(_04576_),
    .C(_10507_),
    .Y(_04581_));
 sg13g2_a21oi_1 _20982_ (.A1(_08103_),
    .A2(_04580_),
    .Y(_04582_),
    .B1(_04581_));
 sg13g2_buf_1 _20983_ (.A(net981),
    .X(_04583_));
 sg13g2_a22oi_1 _20984_ (.Y(_04584_),
    .B1(\top_ihp.wb_emem.cmd[41] ),
    .B2(net865),
    .A2(\top_ihp.wb_emem.cmd[40] ),
    .A1(net942));
 sg13g2_o21ai_1 _20985_ (.B1(_04584_),
    .Y(_02677_),
    .A1(net832),
    .A2(_04582_));
 sg13g2_a21o_1 _20986_ (.A2(_09817_),
    .A1(net790),
    .B1(net973),
    .X(_04585_));
 sg13g2_nor3_1 _20987_ (.A(net1065),
    .B(net780),
    .C(_09817_),
    .Y(_04586_));
 sg13g2_a21oi_1 _20988_ (.A1(net1065),
    .A2(_04585_),
    .Y(_04587_),
    .B1(_04586_));
 sg13g2_a22oi_1 _20989_ (.Y(_04588_),
    .B1(\top_ihp.wb_emem.cmd[42] ),
    .B2(_04542_),
    .A2(\top_ihp.wb_emem.cmd[41] ),
    .A1(net942));
 sg13g2_o21ai_1 _20990_ (.B1(_04588_),
    .Y(_02678_),
    .A1(net832),
    .A2(_04587_));
 sg13g2_xor2_1 _20991_ (.B(_09846_),
    .A(_08028_),
    .X(_04589_));
 sg13g2_a21o_1 _20992_ (.A2(_04589_),
    .A1(net790),
    .B1(net973),
    .X(_04590_));
 sg13g2_nor3_1 _20993_ (.A(net1063),
    .B(net780),
    .C(_04589_),
    .Y(_04591_));
 sg13g2_a21oi_1 _20994_ (.A1(net1063),
    .A2(_04590_),
    .Y(_04592_),
    .B1(_04591_));
 sg13g2_a22oi_1 _20995_ (.Y(_04593_),
    .B1(\top_ihp.wb_emem.cmd[43] ),
    .B2(_04542_),
    .A2(\top_ihp.wb_emem.cmd[42] ),
    .A1(net942));
 sg13g2_o21ai_1 _20996_ (.B1(_04593_),
    .Y(_02679_),
    .A1(net832),
    .A2(_04592_));
 sg13g2_inv_1 _20997_ (.Y(_04594_),
    .A(_08032_));
 sg13g2_xnor2_1 _20998_ (.Y(_04595_),
    .A(_04594_),
    .B(_08230_));
 sg13g2_a21o_1 _20999_ (.A2(_04595_),
    .A1(net790),
    .B1(net973),
    .X(_04596_));
 sg13g2_nor3_1 _21000_ (.A(net1064),
    .B(net780),
    .C(_04595_),
    .Y(_04597_));
 sg13g2_a21oi_1 _21001_ (.A1(net1064),
    .A2(_04596_),
    .Y(_04598_),
    .B1(_04597_));
 sg13g2_a22oi_1 _21002_ (.Y(_04599_),
    .B1(\top_ihp.wb_emem.cmd[44] ),
    .B2(net868),
    .A2(\top_ihp.wb_emem.cmd[43] ),
    .A1(net942));
 sg13g2_o21ai_1 _21003_ (.B1(_04599_),
    .Y(_02680_),
    .A1(net832),
    .A2(_04598_));
 sg13g2_a21o_1 _21004_ (.A2(_09934_),
    .A1(net790),
    .B1(net973),
    .X(_04600_));
 sg13g2_nor3_1 _21005_ (.A(_08046_),
    .B(net780),
    .C(_09934_),
    .Y(_04601_));
 sg13g2_a21oi_1 _21006_ (.A1(_08046_),
    .A2(_04600_),
    .Y(_04602_),
    .B1(_04601_));
 sg13g2_a22oi_1 _21007_ (.Y(_04603_),
    .B1(\top_ihp.wb_emem.cmd[45] ),
    .B2(net868),
    .A2(\top_ihp.wb_emem.cmd[44] ),
    .A1(net942));
 sg13g2_o21ai_1 _21008_ (.B1(_04603_),
    .Y(_02681_),
    .A1(net832),
    .A2(_04602_));
 sg13g2_a21o_1 _21009_ (.A2(_09969_),
    .A1(net790),
    .B1(net973),
    .X(_04604_));
 sg13g2_nor3_1 _21010_ (.A(net1067),
    .B(net780),
    .C(_09969_),
    .Y(_04605_));
 sg13g2_a21oi_1 _21011_ (.A1(net1067),
    .A2(_04604_),
    .Y(_04606_),
    .B1(_04605_));
 sg13g2_a22oi_1 _21012_ (.Y(_04607_),
    .B1(\top_ihp.wb_emem.cmd[46] ),
    .B2(net868),
    .A2(\top_ihp.wb_emem.cmd[45] ),
    .A1(net942));
 sg13g2_o21ai_1 _21013_ (.B1(_04607_),
    .Y(_02682_),
    .A1(net832),
    .A2(_04606_));
 sg13g2_a22oi_1 _21014_ (.Y(_04608_),
    .B1(net781),
    .B2(_09982_),
    .A2(net1068),
    .A1(net939));
 sg13g2_a22oi_1 _21015_ (.Y(_04609_),
    .B1(\top_ihp.wb_emem.cmd[47] ),
    .B2(net868),
    .A2(\top_ihp.wb_emem.cmd[46] ),
    .A1(_04583_));
 sg13g2_o21ai_1 _21016_ (.B1(_04609_),
    .Y(_02683_),
    .A1(_04568_),
    .A2(_04608_));
 sg13g2_o21ai_1 _21017_ (.B1(net971),
    .Y(_04610_),
    .A1(net808),
    .A2(_10005_));
 sg13g2_nand2_1 _21018_ (.Y(_04611_),
    .A(net1069),
    .B(_04610_));
 sg13g2_nand3_1 _21019_ (.B(net781),
    .C(_10005_),
    .A(_08428_),
    .Y(_04612_));
 sg13g2_nand2_1 _21020_ (.Y(_04613_),
    .A(_04611_),
    .B(_04612_));
 sg13g2_inv_1 _21021_ (.Y(_04614_),
    .A(\top_ihp.wb_emem.cmd[47] ));
 sg13g2_a22oi_1 _21022_ (.Y(_04615_),
    .B1(_00308_),
    .B2(_04510_),
    .A2(_04614_),
    .A1(net942));
 sg13g2_o21ai_1 _21023_ (.B1(_04615_),
    .Y(_02684_),
    .A1(_04568_),
    .A2(_04613_));
 sg13g2_xor2_1 _21024_ (.B(_10021_),
    .A(_08006_),
    .X(_04616_));
 sg13g2_a21o_1 _21025_ (.A2(_04616_),
    .A1(net790),
    .B1(net973),
    .X(_04617_));
 sg13g2_nor3_1 _21026_ (.A(_08005_),
    .B(net780),
    .C(_04616_),
    .Y(_04618_));
 sg13g2_a21oi_1 _21027_ (.A1(_08005_),
    .A2(_04617_),
    .Y(_04619_),
    .B1(_04618_));
 sg13g2_a22oi_1 _21028_ (.Y(_04620_),
    .B1(\top_ihp.wb_emem.cmd[49] ),
    .B2(_04510_),
    .A2(\top_ihp.wb_emem.cmd[48] ),
    .A1(net942));
 sg13g2_o21ai_1 _21029_ (.B1(_04620_),
    .Y(_02685_),
    .A1(_04508_),
    .A2(_04619_));
 sg13g2_buf_1 _21030_ (.A(net876),
    .X(_04621_));
 sg13g2_nand2_1 _21031_ (.Y(_04622_),
    .A(\top_ihp.wb_dati_ram[27] ),
    .B(_04504_));
 sg13g2_nand3_1 _21032_ (.B(net836),
    .C(net866),
    .A(_04155_),
    .Y(_04623_));
 sg13g2_a21oi_1 _21033_ (.A1(_04622_),
    .A2(_04623_),
    .Y(_04624_),
    .B1(net867));
 sg13g2_a21o_1 _21034_ (.A2(net847),
    .A1(\top_ihp.wb_dati_ram[28] ),
    .B1(_04624_),
    .X(_02686_));
 sg13g2_a22oi_1 _21035_ (.Y(_04625_),
    .B1(net781),
    .B2(_10052_),
    .A2(net1070),
    .A1(net939));
 sg13g2_a22oi_1 _21036_ (.Y(_04626_),
    .B1(\top_ihp.wb_emem.cmd[50] ),
    .B2(net868),
    .A2(\top_ihp.wb_emem.cmd[49] ),
    .A1(_04583_));
 sg13g2_o21ai_1 _21037_ (.B1(_04626_),
    .Y(_02687_),
    .A1(_04508_),
    .A2(_04625_));
 sg13g2_a21oi_1 _21038_ (.A1(net781),
    .A2(_10065_),
    .Y(_04627_),
    .B1(_07999_));
 sg13g2_nor2_1 _21039_ (.A(net973),
    .B(_08000_),
    .Y(_04628_));
 sg13g2_o21ai_1 _21040_ (.B1(_04628_),
    .Y(_04629_),
    .A1(net780),
    .A2(_10065_));
 sg13g2_nand2b_1 _21041_ (.Y(_04630_),
    .B(_04629_),
    .A_N(_04627_));
 sg13g2_nand2_1 _21042_ (.Y(_04631_),
    .A(_00309_),
    .B(_04441_));
 sg13g2_o21ai_1 _21043_ (.B1(_04631_),
    .Y(_04632_),
    .A1(net982),
    .A2(\top_ihp.wb_emem.cmd[50] ));
 sg13g2_a21o_1 _21044_ (.A2(_04630_),
    .A1(_04450_),
    .B1(_04632_),
    .X(_02688_));
 sg13g2_nand2_1 _21045_ (.Y(_04633_),
    .A(net939),
    .B(_07990_));
 sg13g2_o21ai_1 _21046_ (.B1(_04633_),
    .Y(_04634_),
    .A1(net780),
    .A2(_10141_));
 sg13g2_inv_1 _21047_ (.Y(_04635_),
    .A(\top_ihp.wb_emem.cmd[51] ));
 sg13g2_a22oi_1 _21048_ (.Y(_04636_),
    .B1(_00310_),
    .B2(net868),
    .A2(_04635_),
    .A1(_04565_));
 sg13g2_o21ai_1 _21049_ (.B1(_04636_),
    .Y(_02689_),
    .A1(net849),
    .A2(_04634_));
 sg13g2_xor2_1 _21050_ (.B(_08464_),
    .A(_08153_),
    .X(_04637_));
 sg13g2_o21ai_1 _21051_ (.B1(net971),
    .Y(_04638_),
    .A1(net808),
    .A2(_04637_));
 sg13g2_nor2_1 _21052_ (.A(net1060),
    .B(net808),
    .Y(_04639_));
 sg13g2_a22oi_1 _21053_ (.Y(_04640_),
    .B1(_04639_),
    .B2(_04637_),
    .A2(_04638_),
    .A1(net1060));
 sg13g2_a22oi_1 _21054_ (.Y(_04641_),
    .B1(\top_ihp.wb_emem.cmd[53] ),
    .B2(net868),
    .A2(\top_ihp.wb_emem.cmd[52] ),
    .A1(_04565_));
 sg13g2_o21ai_1 _21055_ (.B1(_04641_),
    .Y(_02690_),
    .A1(net849),
    .A2(_04640_));
 sg13g2_xnor2_1 _21056_ (.Y(_04642_),
    .A(_08393_),
    .B(_10171_));
 sg13g2_a21oi_1 _21057_ (.A1(net781),
    .A2(_04642_),
    .Y(_04643_),
    .B1(_08160_));
 sg13g2_nor2_1 _21058_ (.A(net973),
    .B(_08180_),
    .Y(_04644_));
 sg13g2_o21ai_1 _21059_ (.B1(_04644_),
    .Y(_04645_),
    .A1(net808),
    .A2(_04642_));
 sg13g2_nor2b_1 _21060_ (.A(_04643_),
    .B_N(_04645_),
    .Y(_04646_));
 sg13g2_nand2_1 _21061_ (.Y(_04647_),
    .A(net874),
    .B(_04646_));
 sg13g2_a22oi_1 _21062_ (.Y(_04648_),
    .B1(\top_ihp.wb_emem.cmd[54] ),
    .B2(net865),
    .A2(\top_ihp.wb_emem.cmd[53] ),
    .A1(_04566_));
 sg13g2_nand2_1 _21063_ (.Y(_02691_),
    .A(_04647_),
    .B(_04648_));
 sg13g2_a22oi_1 _21064_ (.Y(_04649_),
    .B1(net781),
    .B2(_10192_),
    .A2(net1061),
    .A1(net939));
 sg13g2_nor2_1 _21065_ (.A(_04402_),
    .B(\top_ihp.wb_emem.cmd[54] ),
    .Y(_04650_));
 sg13g2_a221oi_1 _21066_ (.B2(_04450_),
    .C1(_04650_),
    .B1(_04649_),
    .A1(_00311_),
    .Y(_04651_),
    .A2(net876));
 sg13g2_inv_1 _21067_ (.Y(_02692_),
    .A(_04651_));
 sg13g2_inv_1 _21068_ (.Y(_04652_),
    .A(\top_ihp.wb_emem.cmd[56] ));
 sg13g2_nand2_1 _21069_ (.Y(_04653_),
    .A(\top_ihp.wb_emem.cmd[55] ),
    .B(net871));
 sg13g2_o21ai_1 _21070_ (.B1(_04653_),
    .Y(_04654_),
    .A1(net837),
    .A2(net875));
 sg13g2_nand2_1 _21071_ (.Y(_04655_),
    .A(_04515_),
    .B(_04654_));
 sg13g2_o21ai_1 _21072_ (.B1(_04655_),
    .Y(_02693_),
    .A1(_04652_),
    .A2(_04515_));
 sg13g2_a22oi_1 _21073_ (.Y(_04656_),
    .B1(_00312_),
    .B2(net847),
    .A2(_04652_),
    .A1(net943));
 sg13g2_inv_1 _21074_ (.Y(_02694_),
    .A(_04656_));
 sg13g2_inv_1 _21075_ (.Y(_04657_),
    .A(\top_ihp.wb_emem.cmd[57] ));
 sg13g2_a221oi_1 _21076_ (.B2(net876),
    .C1(net874),
    .B1(_00313_),
    .A1(net981),
    .Y(_04658_),
    .A2(_04657_));
 sg13g2_inv_1 _21077_ (.Y(_02695_),
    .A(_04658_));
 sg13g2_a22oi_1 _21078_ (.Y(_04659_),
    .B1(\top_ihp.wb_emem.cmd[59] ),
    .B2(net847),
    .A2(\top_ihp.wb_emem.cmd[58] ),
    .A1(net943));
 sg13g2_inv_1 _21079_ (.Y(_02696_),
    .A(_04659_));
 sg13g2_nand2_1 _21080_ (.Y(_04660_),
    .A(\top_ihp.wb_dati_ram[28] ),
    .B(net871));
 sg13g2_nand3_1 _21081_ (.B(net836),
    .C(net866),
    .A(_04156_),
    .Y(_04661_));
 sg13g2_a21oi_1 _21082_ (.A1(_04660_),
    .A2(_04661_),
    .Y(_04662_),
    .B1(net867));
 sg13g2_a21o_1 _21083_ (.A2(net847),
    .A1(\top_ihp.wb_dati_ram[29] ),
    .B1(_04662_),
    .X(_02697_));
 sg13g2_a22oi_1 _21084_ (.Y(_04663_),
    .B1(\top_ihp.wb_emem.cmd[60] ),
    .B2(_04621_),
    .A2(\top_ihp.wb_emem.cmd[59] ),
    .A1(net943));
 sg13g2_inv_1 _21085_ (.Y(_02698_),
    .A(_04663_));
 sg13g2_inv_1 _21086_ (.Y(_04664_),
    .A(\top_ihp.wb_emem.cmd[60] ));
 sg13g2_a221oi_1 _21087_ (.B2(net876),
    .C1(net874),
    .B1(_00314_),
    .A1(net981),
    .Y(_04665_),
    .A2(_04664_));
 sg13g2_inv_1 _21088_ (.Y(_02699_),
    .A(_04665_));
 sg13g2_inv_1 _21089_ (.Y(_04666_),
    .A(\top_ihp.wb_emem.cmd[61] ));
 sg13g2_a221oi_1 _21090_ (.B2(net876),
    .C1(net874),
    .B1(_00315_),
    .A1(net981),
    .Y(_04667_),
    .A2(_04666_));
 sg13g2_inv_1 _21091_ (.Y(_02700_),
    .A(_04667_));
 sg13g2_a22oi_1 _21092_ (.Y(_04668_),
    .B1(\top_ihp.wb_emem.cmd[63] ),
    .B2(_04621_),
    .A2(\top_ihp.wb_emem.cmd[62] ),
    .A1(net943));
 sg13g2_inv_1 _21093_ (.Y(_02701_),
    .A(_04668_));
 sg13g2_nand2_1 _21094_ (.Y(_04669_),
    .A(\top_ihp.wb_dati_ram[29] ),
    .B(net871));
 sg13g2_nand3_1 _21095_ (.B(net836),
    .C(net866),
    .A(_04160_),
    .Y(_04670_));
 sg13g2_a21oi_1 _21096_ (.A1(_04669_),
    .A2(_04670_),
    .Y(_04671_),
    .B1(net867));
 sg13g2_a21o_1 _21097_ (.A2(net847),
    .A1(\top_ihp.wb_dati_ram[30] ),
    .B1(_04671_),
    .X(_02702_));
 sg13g2_nand2_1 _21098_ (.Y(_04672_),
    .A(\top_ihp.wb_dati_ram[30] ),
    .B(net871));
 sg13g2_nand3_1 _21099_ (.B(net836),
    .C(net866),
    .A(_04162_),
    .Y(_04673_));
 sg13g2_a21oi_1 _21100_ (.A1(_04672_),
    .A2(_04673_),
    .Y(_04674_),
    .B1(net867));
 sg13g2_a21o_1 _21101_ (.A2(net847),
    .A1(\top_ihp.wb_dati_ram[31] ),
    .B1(_04674_),
    .X(_02703_));
 sg13g2_nand2_1 _21102_ (.Y(_04675_),
    .A(\top_ihp.wb_dati_ram[31] ),
    .B(net871));
 sg13g2_nand3_1 _21103_ (.B(net836),
    .C(_04534_),
    .A(_04126_),
    .Y(_04676_));
 sg13g2_a21oi_1 _21104_ (.A1(_04675_),
    .A2(_04676_),
    .Y(_04677_),
    .B1(net867));
 sg13g2_a21o_1 _21105_ (.A2(net847),
    .A1(\top_ihp.wb_dati_ram[16] ),
    .B1(_04677_),
    .X(_02704_));
 sg13g2_nand2_1 _21106_ (.Y(_04678_),
    .A(\top_ihp.wb_dati_ram[16] ),
    .B(net871));
 sg13g2_nand3_1 _21107_ (.B(net836),
    .C(_04534_),
    .A(_04128_),
    .Y(_04679_));
 sg13g2_a21oi_1 _21108_ (.A1(_04678_),
    .A2(_04679_),
    .Y(_04680_),
    .B1(net867));
 sg13g2_a21o_1 _21109_ (.A2(net847),
    .A1(\top_ihp.wb_dati_ram[17] ),
    .B1(_04680_),
    .X(_02705_));
 sg13g2_buf_1 _21110_ (.A(\top_ihp.wb_emem.nbits[5] ),
    .X(_04681_));
 sg13g2_buf_2 _21111_ (.A(\top_ihp.wb_emem.nbits[3] ),
    .X(_04682_));
 sg13g2_buf_1 _21112_ (.A(\top_ihp.wb_emem.nbits[4] ),
    .X(_04683_));
 sg13g2_nor2_1 _21113_ (.A(_04682_),
    .B(_04683_),
    .Y(_04684_));
 sg13g2_xnor2_1 _21114_ (.Y(_04685_),
    .A(_04681_),
    .B(_04684_));
 sg13g2_buf_1 _21115_ (.A(\top_ihp.wb_emem.nbits[6] ),
    .X(_04686_));
 sg13g2_nand3b_1 _21116_ (.B(_04686_),
    .C(_04684_),
    .Y(_04687_),
    .A_N(_04681_));
 sg13g2_o21ai_1 _21117_ (.B1(_04681_),
    .Y(_04688_),
    .A1(_04682_),
    .A2(_04683_));
 sg13g2_nand3_1 _21118_ (.B(_04687_),
    .C(_04688_),
    .A(_04427_),
    .Y(_04689_));
 sg13g2_o21ai_1 _21119_ (.B1(_04689_),
    .Y(_04690_),
    .A1(_04427_),
    .A2(_04685_));
 sg13g2_nor3_1 _21120_ (.A(_04682_),
    .B(_04683_),
    .C(_04681_),
    .Y(_04691_));
 sg13g2_nand2_1 _21121_ (.Y(_04692_),
    .A(_04437_),
    .B(_04686_));
 sg13g2_o21ai_1 _21122_ (.B1(_04423_),
    .Y(_04693_),
    .A1(_04691_),
    .A2(_04692_));
 sg13g2_xor2_1 _21123_ (.B(_04683_),
    .A(_04682_),
    .X(_04694_));
 sg13g2_nand2_1 _21124_ (.Y(_04695_),
    .A(_04692_),
    .B(_04694_));
 sg13g2_nand2_1 _21125_ (.Y(_04696_),
    .A(_04693_),
    .B(_04695_));
 sg13g2_nand2_1 _21126_ (.Y(_04697_),
    .A(_04682_),
    .B(_04683_));
 sg13g2_o21ai_1 _21127_ (.B1(_04684_),
    .Y(_04698_),
    .A1(_04437_),
    .A2(_04681_));
 sg13g2_nand3_1 _21128_ (.B(_04697_),
    .C(_04698_),
    .A(_04423_),
    .Y(_04699_));
 sg13g2_xor2_1 _21129_ (.B(_04682_),
    .A(_04417_),
    .X(_04700_));
 sg13g2_o21ai_1 _21130_ (.B1(_04700_),
    .Y(_04701_),
    .A1(_04437_),
    .A2(_04686_));
 sg13g2_nor3_1 _21131_ (.A(\top_ihp.wb_emem.bit_counter[7] ),
    .B(_04420_),
    .C(_04701_),
    .Y(_04702_));
 sg13g2_nand3_1 _21132_ (.B(_04699_),
    .C(_04702_),
    .A(_04696_),
    .Y(_04703_));
 sg13g2_nand2_1 _21133_ (.Y(_04704_),
    .A(net1024),
    .B(_04411_));
 sg13g2_o21ai_1 _21134_ (.B1(_04704_),
    .Y(_02706_),
    .A1(_04690_),
    .A2(_04703_));
 sg13g2_inv_1 _21135_ (.Y(_04705_),
    .A(\top_ihp.wb_emem.last_wait ));
 sg13g2_xor2_1 _21136_ (.B(_08779_),
    .A(_08778_),
    .X(_04706_));
 sg13g2_and2_1 _21137_ (.A(net914),
    .B(_04706_),
    .X(_04707_));
 sg13g2_buf_2 _21138_ (.A(_04707_),
    .X(_04708_));
 sg13g2_inv_1 _21139_ (.Y(_04709_),
    .A(\top_ihp.wb_emem.wait_counter[3] ));
 sg13g2_buf_1 _21140_ (.A(\top_ihp.wb_emem.wait_counter[1] ),
    .X(_04710_));
 sg13g2_buf_2 _21141_ (.A(\top_ihp.wb_emem.wait_counter[0] ),
    .X(_04711_));
 sg13g2_nand3_1 _21142_ (.B(_04711_),
    .C(\top_ihp.wb_emem.wait_counter[2] ),
    .A(_04710_),
    .Y(_04712_));
 sg13g2_nor2_1 _21143_ (.A(_04709_),
    .B(_04712_),
    .Y(_04713_));
 sg13g2_buf_1 _21144_ (.A(\top_ihp.wb_emem.wait_counter[5] ),
    .X(_04714_));
 sg13g2_buf_1 _21145_ (.A(\top_ihp.wb_emem.wait_counter[4] ),
    .X(_04715_));
 sg13g2_buf_1 _21146_ (.A(\top_ihp.wb_emem.wait_counter[6] ),
    .X(_04716_));
 sg13g2_nor4_1 _21147_ (.A(_04714_),
    .B(_04715_),
    .C(\top_ihp.wb_emem.wait_counter[7] ),
    .D(_04716_),
    .Y(_04717_));
 sg13g2_nand3_1 _21148_ (.B(_04717_),
    .C(_04708_),
    .A(_04713_),
    .Y(_04718_));
 sg13g2_o21ai_1 _21149_ (.B1(_04718_),
    .Y(_02707_),
    .A1(_04705_),
    .A2(_04708_));
 sg13g2_inv_1 _21150_ (.Y(_04719_),
    .A(_04682_));
 sg13g2_inv_1 _21151_ (.Y(_04720_),
    .A(_08778_));
 sg13g2_nand2_1 _21152_ (.Y(_04721_),
    .A(_04720_),
    .B(_08779_));
 sg13g2_nand3_1 _21153_ (.B(net914),
    .C(_04721_),
    .A(_09490_),
    .Y(_04722_));
 sg13g2_buf_1 _21154_ (.A(_04722_),
    .X(_04723_));
 sg13g2_nand2_1 _21155_ (.Y(_04724_),
    .A(_09490_),
    .B(_04449_));
 sg13g2_inv_1 _21156_ (.Y(_04725_),
    .A(_04724_));
 sg13g2_nand3_1 _21157_ (.B(net837),
    .C(_09639_),
    .A(_08476_),
    .Y(_04726_));
 sg13g2_a22oi_1 _21158_ (.Y(_02708_),
    .B1(_04725_),
    .B2(_04726_),
    .A2(_04723_),
    .A1(_04719_));
 sg13g2_nand3_1 _21159_ (.B(_08478_),
    .C(_08481_),
    .A(net1023),
    .Y(_04727_));
 sg13g2_nor3_1 _21160_ (.A(net883),
    .B(_04724_),
    .C(_04727_),
    .Y(_04728_));
 sg13g2_a21o_1 _21161_ (.A2(_04723_),
    .A1(_04683_),
    .B1(_04728_),
    .X(_02709_));
 sg13g2_nand2_1 _21162_ (.Y(_04729_),
    .A(net837),
    .B(_08478_));
 sg13g2_nand2_1 _21163_ (.Y(_04730_),
    .A(_04681_),
    .B(_04723_));
 sg13g2_o21ai_1 _21164_ (.B1(_04730_),
    .Y(_02710_),
    .A1(_04724_),
    .A2(_04729_));
 sg13g2_a21oi_1 _21165_ (.A1(net837),
    .A2(_08478_),
    .Y(_04731_),
    .B1(_04724_));
 sg13g2_a21o_1 _21166_ (.A2(_04723_),
    .A1(_04686_),
    .B1(_04731_),
    .X(_02711_));
 sg13g2_nor2_1 _21167_ (.A(_08779_),
    .B(_04397_),
    .Y(_04732_));
 sg13g2_a21oi_1 _21168_ (.A1(net1019),
    .A2(_09497_),
    .Y(_04733_),
    .B1(_04445_));
 sg13g2_nor3_1 _21169_ (.A(net1043),
    .B(_08223_),
    .C(_10330_),
    .Y(_04734_));
 sg13g2_nor3_1 _21170_ (.A(_08315_),
    .B(_08223_),
    .C(_10330_),
    .Y(_04735_));
 sg13g2_o21ai_1 _21171_ (.B1(_08351_),
    .Y(_04736_),
    .A1(_04734_),
    .A2(_04735_));
 sg13g2_nand3_1 _21172_ (.B(net809),
    .C(_10330_),
    .A(net1043),
    .Y(_04737_));
 sg13g2_nand3_1 _21173_ (.B(net809),
    .C(_10330_),
    .A(_08315_),
    .Y(_04738_));
 sg13g2_a21o_1 _21174_ (.A2(_04738_),
    .A1(_04737_),
    .B1(_08351_),
    .X(_04739_));
 sg13g2_nor3_1 _21175_ (.A(_08315_),
    .B(net1043),
    .C(_10330_),
    .Y(_04740_));
 sg13g2_nor3_1 _21176_ (.A(_08312_),
    .B(_08311_),
    .C(_09503_),
    .Y(_04741_));
 sg13g2_o21ai_1 _21177_ (.B1(net809),
    .Y(_04742_),
    .A1(_04740_),
    .A2(_04741_));
 sg13g2_nand4_1 _21178_ (.B(_04736_),
    .C(_04739_),
    .A(_04733_),
    .Y(_04743_),
    .D(_04742_));
 sg13g2_inv_1 _21179_ (.Y(_04744_),
    .A(_08779_));
 sg13g2_nor2_1 _21180_ (.A(_08778_),
    .B(_04744_),
    .Y(_04745_));
 sg13g2_nor2_1 _21181_ (.A(net983),
    .B(\top_ihp.wb_emem.last_wait ),
    .Y(_04746_));
 sg13g2_mux2_1 _21182_ (.A0(net983),
    .A1(_04746_),
    .S(_04744_),
    .X(_04747_));
 sg13g2_a21oi_1 _21183_ (.A1(_04396_),
    .A2(net1024),
    .Y(_04748_),
    .B1(net982));
 sg13g2_a221oi_1 _21184_ (.B2(_08778_),
    .C1(_04748_),
    .B1(_04747_),
    .A1(_04745_),
    .Y(_04749_),
    .A2(_04746_));
 sg13g2_and2_1 _21185_ (.A(_04743_),
    .B(_04749_),
    .X(_04750_));
 sg13g2_buf_1 _21186_ (.A(_04750_),
    .X(_04751_));
 sg13g2_nor2b_1 _21187_ (.A(_04732_),
    .B_N(_04751_),
    .Y(_04752_));
 sg13g2_nor2_1 _21188_ (.A(_08779_),
    .B(net983),
    .Y(_04753_));
 sg13g2_nor3_1 _21189_ (.A(_08778_),
    .B(net981),
    .C(_04753_),
    .Y(_04754_));
 sg13g2_nor2_1 _21190_ (.A(_04720_),
    .B(net981),
    .Y(_04755_));
 sg13g2_a22oi_1 _21191_ (.Y(_04756_),
    .B1(_04755_),
    .B2(_04753_),
    .A2(_04754_),
    .A1(_04751_));
 sg13g2_o21ai_1 _21192_ (.B1(_04756_),
    .Y(_02712_),
    .A1(_04720_),
    .A2(_04752_));
 sg13g2_a21o_1 _21193_ (.A2(_04755_),
    .A1(net983),
    .B1(_08779_),
    .X(_02713_));
 sg13g2_a21oi_1 _21194_ (.A1(_04751_),
    .A2(_04753_),
    .Y(_04757_),
    .B1(_04748_));
 sg13g2_o21ai_1 _21195_ (.B1(net913),
    .Y(_04758_),
    .A1(net943),
    .A2(_04751_));
 sg13g2_nand2_1 _21196_ (.Y(_02714_),
    .A(_04757_),
    .B(_04758_));
 sg13g2_nand2_1 _21197_ (.Y(_04759_),
    .A(_04744_),
    .B(net983));
 sg13g2_a21oi_1 _21198_ (.A1(_04721_),
    .A2(_04759_),
    .Y(_04760_),
    .B1(net981));
 sg13g2_nor2_1 _21199_ (.A(net983),
    .B(_04751_),
    .Y(_04761_));
 sg13g2_a21oi_1 _21200_ (.A1(_04751_),
    .A2(_04760_),
    .Y(_02715_),
    .B1(_04761_));
 sg13g2_inv_1 _21201_ (.Y(_04762_),
    .A(_04711_));
 sg13g2_o21ai_1 _21202_ (.B1(_04706_),
    .Y(_04763_),
    .A1(_00233_),
    .A2(_04405_));
 sg13g2_or2_1 _21203_ (.X(_04764_),
    .B(_04706_),
    .A(_04762_));
 sg13g2_a21oi_1 _21204_ (.A1(_04711_),
    .A2(_04759_),
    .Y(_04765_),
    .B1(net982));
 sg13g2_a221oi_1 _21205_ (.B2(_04764_),
    .C1(_04765_),
    .B1(_04763_),
    .A1(net983),
    .Y(_02716_),
    .A2(_04762_));
 sg13g2_nand2_1 _21206_ (.Y(_04766_),
    .A(_04711_),
    .B(_04708_));
 sg13g2_o21ai_1 _21207_ (.B1(_04397_),
    .Y(_04767_),
    .A1(_04720_),
    .A2(_04405_));
 sg13g2_a22oi_1 _21208_ (.Y(_04768_),
    .B1(_04767_),
    .B2(_04744_),
    .A2(_04745_),
    .A1(net914));
 sg13g2_buf_1 _21209_ (.A(_04768_),
    .X(_04769_));
 sg13g2_nand2_1 _21210_ (.Y(_04770_),
    .A(net914),
    .B(_04706_));
 sg13g2_buf_1 _21211_ (.A(_04770_),
    .X(_04771_));
 sg13g2_nor2_1 _21212_ (.A(_04711_),
    .B(_04771_),
    .Y(_04772_));
 sg13g2_o21ai_1 _21213_ (.B1(_04710_),
    .Y(_04773_),
    .A1(_04769_),
    .A2(_04772_));
 sg13g2_o21ai_1 _21214_ (.B1(_04773_),
    .Y(_02717_),
    .A1(_04710_),
    .A2(_04766_));
 sg13g2_nand3_1 _21215_ (.B(_04711_),
    .C(_04708_),
    .A(_04710_),
    .Y(_04774_));
 sg13g2_a21oi_1 _21216_ (.A1(_04710_),
    .A2(_04711_),
    .Y(_04775_),
    .B1(_04771_));
 sg13g2_o21ai_1 _21217_ (.B1(\top_ihp.wb_emem.wait_counter[2] ),
    .Y(_04776_),
    .A1(_04769_),
    .A2(_04775_));
 sg13g2_o21ai_1 _21218_ (.B1(_04776_),
    .Y(_02718_),
    .A1(\top_ihp.wb_emem.wait_counter[2] ),
    .A2(_04774_));
 sg13g2_xnor2_1 _21219_ (.Y(_04777_),
    .A(_04709_),
    .B(_04712_));
 sg13g2_nand2_1 _21220_ (.Y(_04778_),
    .A(\top_ihp.wb_emem.wait_counter[3] ),
    .B(_04769_));
 sg13g2_o21ai_1 _21221_ (.B1(_04778_),
    .Y(_02719_),
    .A1(_04771_),
    .A2(_04777_));
 sg13g2_nand2_1 _21222_ (.Y(_04779_),
    .A(_04713_),
    .B(_04708_));
 sg13g2_nor2_1 _21223_ (.A(_04713_),
    .B(_04771_),
    .Y(_04780_));
 sg13g2_o21ai_1 _21224_ (.B1(_04715_),
    .Y(_04781_),
    .A1(_04769_),
    .A2(_04780_));
 sg13g2_o21ai_1 _21225_ (.B1(_04781_),
    .Y(_02720_),
    .A1(_04715_),
    .A2(_04779_));
 sg13g2_and2_1 _21226_ (.A(_04715_),
    .B(_04713_),
    .X(_04782_));
 sg13g2_buf_1 _21227_ (.A(_04782_),
    .X(_04783_));
 sg13g2_nand2_1 _21228_ (.Y(_04784_),
    .A(_04708_),
    .B(_04783_));
 sg13g2_nor2_1 _21229_ (.A(_04771_),
    .B(_04783_),
    .Y(_04785_));
 sg13g2_o21ai_1 _21230_ (.B1(_04714_),
    .Y(_04786_),
    .A1(_04769_),
    .A2(_04785_));
 sg13g2_o21ai_1 _21231_ (.B1(_04786_),
    .Y(_02721_),
    .A1(_04714_),
    .A2(_04784_));
 sg13g2_nand2_1 _21232_ (.Y(_04787_),
    .A(_04714_),
    .B(_04783_));
 sg13g2_xor2_1 _21233_ (.B(_04787_),
    .A(_04716_),
    .X(_04788_));
 sg13g2_nand2_1 _21234_ (.Y(_04789_),
    .A(_04716_),
    .B(_04769_));
 sg13g2_o21ai_1 _21235_ (.B1(_04789_),
    .Y(_02722_),
    .A1(_04771_),
    .A2(_04788_));
 sg13g2_nand4_1 _21236_ (.B(_04716_),
    .C(_04708_),
    .A(_04714_),
    .Y(_04790_),
    .D(_04783_));
 sg13g2_nand3b_1 _21237_ (.B(_04790_),
    .C(\top_ihp.wb_emem.wait_counter[7] ),
    .Y(_04791_),
    .A_N(_04732_));
 sg13g2_o21ai_1 _21238_ (.B1(_04791_),
    .Y(_02723_),
    .A1(\top_ihp.wb_emem.wait_counter[7] ),
    .A2(_04790_));
 sg13g2_mux4_1 _21239_ (.S0(\top_ihp.oisc.wb_adr_o[0] ),
    .A0(net6),
    .A1(net7),
    .A2(net8),
    .A3(net9),
    .S1(\top_ihp.oisc.wb_adr_o[1] ),
    .X(_04792_));
 sg13g2_nand3_1 _21240_ (.B(net883),
    .C(_08303_),
    .A(_08219_),
    .Y(_04793_));
 sg13g2_mux2_1 _21241_ (.A0(_04792_),
    .A1(\top_ihp.wb_dati_gpio[0] ),
    .S(_04793_),
    .X(_02724_));
 sg13g2_and3_1 _21242_ (.X(_04794_),
    .A(_08219_),
    .B(_08640_),
    .C(_08303_));
 sg13g2_buf_1 _21243_ (.A(_04794_),
    .X(_04795_));
 sg13g2_and2_1 _21244_ (.A(net1050),
    .B(_04192_),
    .X(_04796_));
 sg13g2_nand3_1 _21245_ (.B(net857),
    .C(net781),
    .A(_08219_),
    .Y(_04797_));
 sg13g2_nand4_1 _21246_ (.B(net1057),
    .C(_08219_),
    .A(_07987_),
    .Y(_04798_),
    .D(net857));
 sg13g2_o21ai_1 _21247_ (.B1(_04798_),
    .Y(_04799_),
    .A1(_08301_),
    .A2(_04797_));
 sg13g2_inv_1 _21248_ (.Y(_04800_),
    .A(\top_ihp.gpio_o_1 ));
 sg13g2_a21oi_1 _21249_ (.A1(_04192_),
    .A2(_04799_),
    .Y(_04801_),
    .B1(_04800_));
 sg13g2_a21o_1 _21250_ (.A2(_04796_),
    .A1(_04795_),
    .B1(_04801_),
    .X(_02725_));
 sg13g2_nand2_1 _21251_ (.Y(_04802_),
    .A(_08457_),
    .B(\top_ihp.oisc.wb_adr_o[0] ));
 sg13g2_mux2_1 _21252_ (.A0(net1050),
    .A1(\top_ihp.gpio_o_2 ),
    .S(_04802_),
    .X(_04803_));
 sg13g2_inv_1 _21253_ (.Y(_04804_),
    .A(_04803_));
 sg13g2_mux2_1 _21254_ (.A0(_00316_),
    .A1(_04804_),
    .S(_04795_),
    .X(_02726_));
 sg13g2_nor3_1 _21255_ (.A(_00185_),
    .B(_08457_),
    .C(\top_ihp.oisc.wb_adr_o[0] ),
    .Y(_04805_));
 sg13g2_nor2_1 _21256_ (.A(_08457_),
    .B(\top_ihp.oisc.wb_adr_o[0] ),
    .Y(_04806_));
 sg13g2_inv_1 _21257_ (.Y(_04807_),
    .A(\top_ihp.gpio_o_3 ));
 sg13g2_a21oi_1 _21258_ (.A1(_04799_),
    .A2(_04806_),
    .Y(_04808_),
    .B1(_04807_));
 sg13g2_a21o_1 _21259_ (.A2(_04805_),
    .A1(_04795_),
    .B1(_04808_),
    .X(_02727_));
 sg13g2_nand2_1 _21260_ (.Y(_04809_),
    .A(\top_ihp.oisc.wb_adr_o[1] ),
    .B(\top_ihp.oisc.wb_adr_o[0] ));
 sg13g2_mux2_1 _21261_ (.A0(_04110_),
    .A1(\top_ihp.gpio_o_4 ),
    .S(_04809_),
    .X(_04810_));
 sg13g2_inv_1 _21262_ (.Y(_04811_),
    .A(_04810_));
 sg13g2_mux2_1 _21263_ (.A0(_00317_),
    .A1(_04811_),
    .S(_04795_),
    .X(_02728_));
 sg13g2_inv_1 _21264_ (.Y(_04812_),
    .A(_08360_));
 sg13g2_nor2_1 _21265_ (.A(_09631_),
    .B(_08366_),
    .Y(_04813_));
 sg13g2_buf_1 _21266_ (.A(_04813_),
    .X(_04814_));
 sg13g2_buf_1 _21267_ (.A(_04814_),
    .X(_04815_));
 sg13g2_a21oi_1 _21268_ (.A1(_08304_),
    .A2(_08359_),
    .Y(_04816_),
    .B1(net896));
 sg13g2_buf_1 _21269_ (.A(_04816_),
    .X(_04817_));
 sg13g2_mux2_1 _21270_ (.A0(_08309_),
    .A1(_04814_),
    .S(_08305_),
    .X(_04818_));
 sg13g2_a21oi_1 _21271_ (.A1(_08304_),
    .A2(_08357_),
    .Y(_04819_),
    .B1(_04818_));
 sg13g2_buf_2 _21272_ (.A(_04819_),
    .X(_04820_));
 sg13g2_buf_1 _21273_ (.A(_04820_),
    .X(_04821_));
 sg13g2_nor2_1 _21274_ (.A(_04812_),
    .B(net210),
    .Y(_04822_));
 sg13g2_a21o_1 _21275_ (.A2(net64),
    .A1(_04812_),
    .B1(_04822_),
    .X(_02729_));
 sg13g2_buf_8 _21276_ (.A(_04820_),
    .X(_04823_));
 sg13g2_inv_1 _21277_ (.Y(_04824_),
    .A(_08368_));
 sg13g2_a21oi_1 _21278_ (.A1(net992),
    .A2(_04824_),
    .Y(_04825_),
    .B1(_08366_));
 sg13g2_nand2b_1 _21279_ (.Y(_04826_),
    .B(_08360_),
    .A_N(_04825_));
 sg13g2_a21oi_1 _21280_ (.A1(net209),
    .A2(_04826_),
    .Y(_04827_),
    .B1(_08361_));
 sg13g2_nand3b_1 _21281_ (.B(net210),
    .C(_08369_),
    .Y(_04828_),
    .A_N(_04825_));
 sg13g2_nand2b_1 _21282_ (.Y(_02730_),
    .B(_04828_),
    .A_N(_04827_));
 sg13g2_a21o_1 _21283_ (.A2(_08365_),
    .A1(_08368_),
    .B1(_04825_),
    .X(_04829_));
 sg13g2_buf_1 _21284_ (.A(_04829_),
    .X(_04830_));
 sg13g2_nor3_1 _21285_ (.A(_08360_),
    .B(\top_ihp.wb_imem.bits_left[1] ),
    .C(_08362_),
    .Y(_04831_));
 sg13g2_nor2b_1 _21286_ (.A(_08369_),
    .B_N(_08362_),
    .Y(_04832_));
 sg13g2_a21oi_1 _21287_ (.A1(net209),
    .A2(_04831_),
    .Y(_04833_),
    .B1(_04832_));
 sg13g2_nand2b_1 _21288_ (.Y(_04834_),
    .B(_08362_),
    .A_N(net209));
 sg13g2_o21ai_1 _21289_ (.B1(_04834_),
    .Y(_02731_),
    .A1(_04830_),
    .A2(_04833_));
 sg13g2_o21ai_1 _21290_ (.B1(_04823_),
    .Y(_04835_),
    .A1(_04830_),
    .A2(_04831_));
 sg13g2_nand2b_1 _21291_ (.Y(_04836_),
    .B(_04831_),
    .A_N(\top_ihp.wb_imem.bits_left[3] ));
 sg13g2_nor2_1 _21292_ (.A(_04830_),
    .B(_04836_),
    .Y(_04837_));
 sg13g2_and2_1 _21293_ (.A(_04820_),
    .B(_04837_),
    .X(_04838_));
 sg13g2_a21o_1 _21294_ (.A2(_04835_),
    .A1(\top_ihp.wb_imem.bits_left[3] ),
    .B1(_04838_),
    .X(_02732_));
 sg13g2_inv_1 _21295_ (.Y(_04839_),
    .A(_04836_));
 sg13g2_o21ai_1 _21296_ (.B1(net209),
    .Y(_04840_),
    .A1(_04830_),
    .A2(_04839_));
 sg13g2_mux2_1 _21297_ (.A0(_04838_),
    .A1(_04840_),
    .S(\top_ihp.wb_imem.bits_left[4] ),
    .X(_02733_));
 sg13g2_nand3b_1 _21298_ (.B(_04820_),
    .C(_04839_),
    .Y(_04841_),
    .A_N(\top_ihp.wb_imem.bits_left[4] ));
 sg13g2_nor2_1 _21299_ (.A(_08372_),
    .B(net896),
    .Y(_04842_));
 sg13g2_a221oi_1 _21300_ (.B2(_04842_),
    .C1(_04818_),
    .B1(_08373_),
    .A1(_08304_),
    .Y(_04843_),
    .A2(_08357_));
 sg13g2_a21o_1 _21301_ (.A2(_04841_),
    .A1(\top_ihp.wb_imem.bits_left[5] ),
    .B1(_04843_),
    .X(_02734_));
 sg13g2_buf_1 _21302_ (.A(_04820_),
    .X(_04844_));
 sg13g2_buf_1 _21303_ (.A(_04815_),
    .X(_04845_));
 sg13g2_a22oi_1 _21304_ (.Y(_04846_),
    .B1(\top_ihp.oisc.wb_adr_o[0] ),
    .B2(_04845_),
    .A2(net3),
    .A1(net992));
 sg13g2_nor2_1 _21305_ (.A(\top_ihp.wb_dati_rom[24] ),
    .B(net210),
    .Y(_04847_));
 sg13g2_a21oi_1 _21306_ (.A1(_04844_),
    .A2(_04846_),
    .Y(_02735_),
    .B1(_04847_));
 sg13g2_buf_1 _21307_ (.A(_04814_),
    .X(_04848_));
 sg13g2_nor2_1 _21308_ (.A(\top_ihp.wb_dati_rom[17] ),
    .B(net895),
    .Y(_04849_));
 sg13g2_a21oi_1 _21309_ (.A1(_04587_),
    .A2(net887),
    .Y(_04850_),
    .B1(_04849_));
 sg13g2_mux2_1 _21310_ (.A0(\top_ihp.wb_dati_rom[18] ),
    .A1(_04850_),
    .S(net208),
    .X(_02736_));
 sg13g2_nor2_1 _21311_ (.A(\top_ihp.wb_dati_rom[18] ),
    .B(net895),
    .Y(_04851_));
 sg13g2_a21oi_1 _21312_ (.A1(_04592_),
    .A2(net887),
    .Y(_04852_),
    .B1(_04851_));
 sg13g2_mux2_1 _21313_ (.A0(\top_ihp.wb_dati_rom[19] ),
    .A1(_04852_),
    .S(net208),
    .X(_02737_));
 sg13g2_nor2_1 _21314_ (.A(\top_ihp.wb_dati_rom[19] ),
    .B(net895),
    .Y(_04853_));
 sg13g2_a21oi_1 _21315_ (.A1(_04598_),
    .A2(net887),
    .Y(_04854_),
    .B1(_04853_));
 sg13g2_mux2_1 _21316_ (.A0(\top_ihp.wb_dati_rom[20] ),
    .A1(_04854_),
    .S(net208),
    .X(_02738_));
 sg13g2_nor2_1 _21317_ (.A(\top_ihp.wb_dati_rom[20] ),
    .B(net895),
    .Y(_04855_));
 sg13g2_a21oi_1 _21318_ (.A1(_04602_),
    .A2(net887),
    .Y(_04856_),
    .B1(_04855_));
 sg13g2_mux2_1 _21319_ (.A0(\top_ihp.wb_dati_rom[21] ),
    .A1(_04856_),
    .S(net208),
    .X(_02739_));
 sg13g2_nor2_1 _21320_ (.A(\top_ihp.wb_dati_rom[21] ),
    .B(net895),
    .Y(_04857_));
 sg13g2_a21oi_1 _21321_ (.A1(_04606_),
    .A2(net887),
    .Y(_04858_),
    .B1(_04857_));
 sg13g2_mux2_1 _21322_ (.A0(\top_ihp.wb_dati_rom[22] ),
    .A1(_04858_),
    .S(net208),
    .X(_02740_));
 sg13g2_nor2_1 _21323_ (.A(\top_ihp.wb_dati_rom[22] ),
    .B(net895),
    .Y(_04859_));
 sg13g2_a21oi_1 _21324_ (.A1(_04608_),
    .A2(net887),
    .Y(_04860_),
    .B1(_04859_));
 sg13g2_mux2_1 _21325_ (.A0(\top_ihp.wb_dati_rom[23] ),
    .A1(_04860_),
    .S(net208),
    .X(_02741_));
 sg13g2_mux2_1 _21326_ (.A0(\top_ihp.wb_dati_rom[23] ),
    .A1(_04613_),
    .S(net895),
    .X(_04861_));
 sg13g2_mux2_1 _21327_ (.A0(\top_ihp.wb_dati_rom[8] ),
    .A1(_04861_),
    .S(net208),
    .X(_02742_));
 sg13g2_buf_1 _21328_ (.A(_04814_),
    .X(_04862_));
 sg13g2_nor2_1 _21329_ (.A(\top_ihp.wb_dati_rom[8] ),
    .B(net894),
    .Y(_04863_));
 sg13g2_a21oi_1 _21330_ (.A1(_04619_),
    .A2(net887),
    .Y(_04864_),
    .B1(_04863_));
 sg13g2_mux2_1 _21331_ (.A0(\top_ihp.wb_dati_rom[9] ),
    .A1(_04864_),
    .S(net208),
    .X(_02743_));
 sg13g2_nor2_1 _21332_ (.A(\top_ihp.wb_dati_rom[9] ),
    .B(_04862_),
    .Y(_04865_));
 sg13g2_a21oi_1 _21333_ (.A1(_04625_),
    .A2(net887),
    .Y(_04866_),
    .B1(_04865_));
 sg13g2_buf_1 _21334_ (.A(_04820_),
    .X(_04867_));
 sg13g2_mux2_1 _21335_ (.A0(\top_ihp.wb_dati_rom[10] ),
    .A1(_04866_),
    .S(_04867_),
    .X(_02744_));
 sg13g2_buf_1 _21336_ (.A(net896),
    .X(_04868_));
 sg13g2_nor2_1 _21337_ (.A(\top_ihp.wb_dati_rom[10] ),
    .B(_04862_),
    .Y(_04869_));
 sg13g2_a21oi_1 _21338_ (.A1(_04630_),
    .A2(net886),
    .Y(_04870_),
    .B1(_04869_));
 sg13g2_mux2_1 _21339_ (.A0(\top_ihp.wb_dati_rom[11] ),
    .A1(_04870_),
    .S(net207),
    .X(_02745_));
 sg13g2_nor2_1 _21340_ (.A(\top_ihp.wb_dati_rom[24] ),
    .B(net894),
    .Y(_04871_));
 sg13g2_a21oi_1 _21341_ (.A1(_08457_),
    .A2(net886),
    .Y(_04872_),
    .B1(_04871_));
 sg13g2_mux2_1 _21342_ (.A0(\top_ihp.wb_dati_rom[25] ),
    .A1(_04872_),
    .S(net207),
    .X(_02746_));
 sg13g2_mux2_1 _21343_ (.A0(\top_ihp.wb_dati_rom[11] ),
    .A1(_04634_),
    .S(net895),
    .X(_04873_));
 sg13g2_mux2_1 _21344_ (.A0(\top_ihp.wb_dati_rom[12] ),
    .A1(_04873_),
    .S(_04867_),
    .X(_02747_));
 sg13g2_inv_1 _21345_ (.Y(_04874_),
    .A(\top_ihp.wb_dati_rom[13] ));
 sg13g2_nor2_1 _21346_ (.A(\top_ihp.wb_dati_rom[12] ),
    .B(net896),
    .Y(_04875_));
 sg13g2_a21oi_1 _21347_ (.A1(_04640_),
    .A2(_04848_),
    .Y(_04876_),
    .B1(_04875_));
 sg13g2_nand2_1 _21348_ (.Y(_04877_),
    .A(net210),
    .B(_04876_));
 sg13g2_o21ai_1 _21349_ (.B1(_04877_),
    .Y(_02748_),
    .A1(_04874_),
    .A2(_04844_));
 sg13g2_nand2_1 _21350_ (.Y(_04878_),
    .A(_04646_),
    .B(_04845_));
 sg13g2_o21ai_1 _21351_ (.B1(_08304_),
    .Y(_04879_),
    .A1(_04874_),
    .A2(net896));
 sg13g2_nor2_1 _21352_ (.A(_08359_),
    .B(_04879_),
    .Y(_04880_));
 sg13g2_nor2_1 _21353_ (.A(_08305_),
    .B(\top_ihp.wb_dati_rom[14] ),
    .Y(_04881_));
 sg13g2_nand2_1 _21354_ (.Y(_04882_),
    .A(\top_ihp.wb_dati_rom[14] ),
    .B(net896));
 sg13g2_o21ai_1 _21355_ (.B1(_04882_),
    .Y(_04883_),
    .A1(_04874_),
    .A2(_04815_));
 sg13g2_nor2_1 _21356_ (.A(_08304_),
    .B(_04883_),
    .Y(_04884_));
 sg13g2_a221oi_1 _21357_ (.B2(_08359_),
    .C1(_04884_),
    .B1(_04881_),
    .A1(_04878_),
    .Y(_02749_),
    .A2(_04880_));
 sg13g2_nor2_1 _21358_ (.A(\top_ihp.wb_dati_rom[14] ),
    .B(net894),
    .Y(_04885_));
 sg13g2_a21oi_1 _21359_ (.A1(_04649_),
    .A2(net886),
    .Y(_04886_),
    .B1(_04885_));
 sg13g2_mux2_1 _21360_ (.A0(\top_ihp.wb_dati_rom[15] ),
    .A1(_04886_),
    .S(net207),
    .X(_02750_));
 sg13g2_inv_1 _21361_ (.Y(_04887_),
    .A(\top_ihp.wb_dati_rom[15] ));
 sg13g2_nor2_1 _21362_ (.A(\top_ihp.wb_dati_rom[0] ),
    .B(net210),
    .Y(_04888_));
 sg13g2_a21oi_1 _21363_ (.A1(_04887_),
    .A2(net64),
    .Y(_02751_),
    .B1(_04888_));
 sg13g2_inv_1 _21364_ (.Y(_04889_),
    .A(\top_ihp.wb_dati_rom[0] ));
 sg13g2_nor2_1 _21365_ (.A(\top_ihp.wb_dati_rom[1] ),
    .B(_04821_),
    .Y(_04890_));
 sg13g2_a21oi_1 _21366_ (.A1(_04889_),
    .A2(net64),
    .Y(_02752_),
    .B1(_04890_));
 sg13g2_nor2b_1 _21367_ (.A(_04821_),
    .B_N(\top_ihp.wb_dati_rom[2] ),
    .Y(_04891_));
 sg13g2_a21o_1 _21368_ (.A2(net64),
    .A1(\top_ihp.wb_dati_rom[1] ),
    .B1(_04891_),
    .X(_02753_));
 sg13g2_nor2b_1 _21369_ (.A(net209),
    .B_N(\top_ihp.wb_dati_rom[3] ),
    .Y(_04892_));
 sg13g2_a21o_1 _21370_ (.A2(net64),
    .A1(\top_ihp.wb_dati_rom[2] ),
    .B1(_04892_),
    .X(_02754_));
 sg13g2_nor2b_1 _21371_ (.A(net209),
    .B_N(\top_ihp.wb_dati_rom[4] ),
    .Y(_04893_));
 sg13g2_a21o_1 _21372_ (.A2(net64),
    .A1(\top_ihp.wb_dati_rom[3] ),
    .B1(_04893_),
    .X(_02755_));
 sg13g2_nor2b_1 _21373_ (.A(net209),
    .B_N(\top_ihp.wb_dati_rom[5] ),
    .Y(_04894_));
 sg13g2_a21o_1 _21374_ (.A2(_04817_),
    .A1(\top_ihp.wb_dati_rom[4] ),
    .B1(_04894_),
    .X(_02756_));
 sg13g2_nor2_1 _21375_ (.A(\top_ihp.wb_dati_rom[25] ),
    .B(net894),
    .Y(_04895_));
 sg13g2_a21oi_1 _21376_ (.A1(_04383_),
    .A2(net886),
    .Y(_04896_),
    .B1(_04895_));
 sg13g2_mux2_1 _21377_ (.A0(\top_ihp.wb_dati_rom[26] ),
    .A1(_04896_),
    .S(net207),
    .X(_02757_));
 sg13g2_nor2b_1 _21378_ (.A(net209),
    .B_N(\top_ihp.wb_dati_rom[6] ),
    .Y(_04897_));
 sg13g2_a21o_1 _21379_ (.A2(net64),
    .A1(\top_ihp.wb_dati_rom[5] ),
    .B1(_04897_),
    .X(_02758_));
 sg13g2_nor2b_1 _21380_ (.A(_04823_),
    .B_N(\top_ihp.wb_dati_rom[7] ),
    .Y(_04898_));
 sg13g2_a21o_1 _21381_ (.A2(net64),
    .A1(\top_ihp.wb_dati_rom[6] ),
    .B1(_04898_),
    .X(_02759_));
 sg13g2_nor2_1 _21382_ (.A(\top_ihp.wb_dati_rom[26] ),
    .B(net894),
    .Y(_04899_));
 sg13g2_a21oi_1 _21383_ (.A1(_04183_),
    .A2(net886),
    .Y(_04900_),
    .B1(_04899_));
 sg13g2_mux2_1 _21384_ (.A0(\top_ihp.wb_dati_rom[27] ),
    .A1(_04900_),
    .S(net207),
    .X(_02760_));
 sg13g2_nor2_1 _21385_ (.A(\top_ihp.wb_dati_rom[27] ),
    .B(net894),
    .Y(_04901_));
 sg13g2_a21oi_1 _21386_ (.A1(_04187_),
    .A2(net886),
    .Y(_04902_),
    .B1(_04901_));
 sg13g2_mux2_1 _21387_ (.A0(\top_ihp.wb_dati_rom[28] ),
    .A1(_04902_),
    .S(net207),
    .X(_02761_));
 sg13g2_nor2_1 _21388_ (.A(\top_ihp.wb_dati_rom[28] ),
    .B(net894),
    .Y(_04903_));
 sg13g2_a21oi_1 _21389_ (.A1(_04558_),
    .A2(_04868_),
    .Y(_04904_),
    .B1(_04903_));
 sg13g2_mux2_1 _21390_ (.A0(\top_ihp.wb_dati_rom[29] ),
    .A1(_04904_),
    .S(net207),
    .X(_02762_));
 sg13g2_mux2_1 _21391_ (.A0(\top_ihp.wb_dati_rom[29] ),
    .A1(_04563_),
    .S(_04848_),
    .X(_04905_));
 sg13g2_mux2_1 _21392_ (.A0(\top_ihp.wb_dati_rom[30] ),
    .A1(_04905_),
    .S(net207),
    .X(_02763_));
 sg13g2_nor2_1 _21393_ (.A(\top_ihp.wb_dati_rom[30] ),
    .B(net894),
    .Y(_04906_));
 sg13g2_a21oi_1 _21394_ (.A1(_04570_),
    .A2(net886),
    .Y(_04907_),
    .B1(_04906_));
 sg13g2_mux2_1 _21395_ (.A0(\top_ihp.wb_dati_rom[31] ),
    .A1(_04907_),
    .S(net210),
    .X(_02764_));
 sg13g2_nor2_1 _21396_ (.A(\top_ihp.wb_dati_rom[31] ),
    .B(net896),
    .Y(_04908_));
 sg13g2_a21oi_1 _21397_ (.A1(_04578_),
    .A2(_04868_),
    .Y(_04909_),
    .B1(_04908_));
 sg13g2_mux2_1 _21398_ (.A0(\top_ihp.wb_dati_rom[16] ),
    .A1(_04909_),
    .S(net210),
    .X(_02765_));
 sg13g2_nor2_1 _21399_ (.A(\top_ihp.wb_dati_rom[16] ),
    .B(net896),
    .Y(_04910_));
 sg13g2_a21oi_1 _21400_ (.A1(_04582_),
    .A2(net886),
    .Y(_04911_),
    .B1(_04910_));
 sg13g2_mux2_1 _21401_ (.A0(\top_ihp.wb_dati_rom[17] ),
    .A1(_04911_),
    .S(net210),
    .X(_02766_));
 sg13g2_inv_1 _21402_ (.Y(_04912_),
    .A(_08359_));
 sg13g2_nor2_1 _21403_ (.A(_08368_),
    .B(_09609_),
    .Y(_04913_));
 sg13g2_nor2_1 _21404_ (.A(net992),
    .B(_08368_),
    .Y(_04914_));
 sg13g2_inv_1 _21405_ (.Y(_04915_),
    .A(_00318_));
 sg13g2_mux2_1 _21406_ (.A0(_04914_),
    .A1(_04915_),
    .S(_08359_),
    .X(_04916_));
 sg13g2_nor2_1 _21407_ (.A(_00318_),
    .B(net900),
    .Y(_04917_));
 sg13g2_o21ai_1 _21408_ (.B1(_08305_),
    .Y(_04918_),
    .A1(_04913_),
    .A2(_04917_));
 sg13g2_nand2_1 _21409_ (.Y(_04919_),
    .A(_09631_),
    .B(_04917_));
 sg13g2_nand2_1 _21410_ (.Y(_04920_),
    .A(_04918_),
    .B(_04919_));
 sg13g2_a221oi_1 _21411_ (.B2(_08304_),
    .C1(_04920_),
    .B1(_04916_),
    .A1(_04912_),
    .Y(_02767_),
    .A2(_04913_));
 sg13g2_nand2b_1 _21412_ (.Y(_04921_),
    .B(\top_ihp.spi_clk_o ),
    .A_N(\top_ihp.wb_spi.spi_clk_cnt[0] ));
 sg13g2_and2_1 _21413_ (.A(_08168_),
    .B(_08171_),
    .X(_04922_));
 sg13g2_nand4_1 _21414_ (.B(_07988_),
    .C(net974),
    .A(net971),
    .Y(_04923_),
    .D(net857));
 sg13g2_nand2_1 _21415_ (.Y(_04924_),
    .A(_07977_),
    .B(_08469_));
 sg13g2_a22oi_1 _21416_ (.Y(_04925_),
    .B1(_04923_),
    .B2(_04924_),
    .A2(_08186_),
    .A1(_04922_));
 sg13g2_nand4_1 _21417_ (.B(_07989_),
    .C(net974),
    .A(net971),
    .Y(_04926_),
    .D(_07976_));
 sg13g2_nand3_1 _21418_ (.B(net1048),
    .C(net857),
    .A(_07988_),
    .Y(_04927_));
 sg13g2_a21oi_1 _21419_ (.A1(_04926_),
    .A2(_04927_),
    .Y(_04928_),
    .B1(_08188_));
 sg13g2_nand2_1 _21420_ (.Y(_04929_),
    .A(net1019),
    .B(net1048));
 sg13g2_o21ai_1 _21421_ (.B1(_00091_),
    .Y(_04930_),
    .A1(net883),
    .A2(_04929_));
 sg13g2_nor3_2 _21422_ (.A(_04925_),
    .B(_04928_),
    .C(_04930_),
    .Y(_04931_));
 sg13g2_a21o_1 _21423_ (.A2(_04921_),
    .A1(_08192_),
    .B1(_04931_),
    .X(_04932_));
 sg13g2_buf_2 _21424_ (.A(_04932_),
    .X(_04933_));
 sg13g2_inv_2 _21425_ (.Y(_04934_),
    .A(_08192_));
 sg13g2_nor2_1 _21426_ (.A(net1059),
    .B(_04934_),
    .Y(_04935_));
 sg13g2_nand2b_1 _21427_ (.Y(_04936_),
    .B(_04935_),
    .A_N(_04933_));
 sg13g2_buf_1 _21428_ (.A(_04933_),
    .X(_04937_));
 sg13g2_nand2_1 _21429_ (.Y(_04938_),
    .A(net1059),
    .B(_04937_));
 sg13g2_nand2_1 _21430_ (.Y(_02768_),
    .A(_04936_),
    .B(_04938_));
 sg13g2_o21ai_1 _21431_ (.B1(_08193_),
    .Y(_04939_),
    .A1(_08197_),
    .A2(_04921_));
 sg13g2_inv_1 _21432_ (.Y(_04940_),
    .A(_04939_));
 sg13g2_o21ai_1 _21433_ (.B1(_08198_),
    .Y(_04941_),
    .A1(_04931_),
    .A2(_04940_));
 sg13g2_o21ai_1 _21434_ (.B1(_04941_),
    .Y(_02769_),
    .A1(_08198_),
    .A2(_04936_));
 sg13g2_nor3_1 _21435_ (.A(net1059),
    .B(_08198_),
    .C(_04921_),
    .Y(_04942_));
 sg13g2_nor2_1 _21436_ (.A(_04934_),
    .B(_04942_),
    .Y(_04943_));
 sg13g2_o21ai_1 _21437_ (.B1(\top_ihp.wb_spi.bits_left[2] ),
    .Y(_04944_),
    .A1(_04931_),
    .A2(_04943_));
 sg13g2_o21ai_1 _21438_ (.B1(_04944_),
    .Y(_02770_),
    .A1(_08200_),
    .A2(_04936_));
 sg13g2_buf_8 _21439_ (.A(_04933_),
    .X(_04945_));
 sg13g2_buf_8 _21440_ (.A(net443),
    .X(_04946_));
 sg13g2_and3_1 _21441_ (.X(_04947_),
    .A(_08476_),
    .B(_08481_),
    .C(_09639_));
 sg13g2_buf_1 _21442_ (.A(_04947_),
    .X(_04948_));
 sg13g2_nor3_1 _21443_ (.A(net1059),
    .B(\top_ihp.wb_spi.bits_left[3] ),
    .C(_08200_),
    .Y(_04949_));
 sg13g2_and2_1 _21444_ (.A(net1018),
    .B(_04949_),
    .X(_04950_));
 sg13g2_a21oi_1 _21445_ (.A1(_04934_),
    .A2(net802),
    .Y(_04951_),
    .B1(_04950_));
 sg13g2_o21ai_1 _21446_ (.B1(_08193_),
    .Y(_04952_),
    .A1(net1059),
    .A2(_08200_));
 sg13g2_a21oi_1 _21447_ (.A1(net1059),
    .A2(_08202_),
    .Y(_04953_),
    .B1(_04952_));
 sg13g2_o21ai_1 _21448_ (.B1(\top_ihp.wb_spi.bits_left[3] ),
    .Y(_04954_),
    .A1(_04945_),
    .A2(_04953_));
 sg13g2_o21ai_1 _21449_ (.B1(_04954_),
    .Y(_02771_),
    .A1(_04946_),
    .A2(_04951_));
 sg13g2_inv_1 _21450_ (.Y(_04955_),
    .A(\top_ihp.wb_spi.bits_left[4] ));
 sg13g2_a21oi_1 _21451_ (.A1(_08203_),
    .A2(_04949_),
    .Y(_04956_),
    .B1(_04934_));
 sg13g2_o21ai_1 _21452_ (.B1(\top_ihp.wb_spi.bits_left[4] ),
    .Y(_04957_),
    .A1(_04931_),
    .A2(_04956_));
 sg13g2_nor2_1 _21453_ (.A(net1059),
    .B(_08201_),
    .Y(_04958_));
 sg13g2_buf_1 _21454_ (.A(_08193_),
    .X(_04959_));
 sg13g2_nor2_1 _21455_ (.A(_04959_),
    .B(_04727_),
    .Y(_04960_));
 sg13g2_a21oi_1 _21456_ (.A1(_08195_),
    .A2(_04958_),
    .Y(_04961_),
    .B1(_04960_));
 sg13g2_a22oi_1 _21457_ (.Y(_02772_),
    .B1(_04957_),
    .B2(_04961_),
    .A2(_04946_),
    .A1(_04955_));
 sg13g2_buf_1 _21458_ (.A(_08483_),
    .X(_04962_));
 sg13g2_a22oi_1 _21459_ (.Y(_04963_),
    .B1(_04935_),
    .B2(_08202_),
    .A2(_04962_),
    .A1(_04934_));
 sg13g2_a21oi_1 _21460_ (.A1(_08203_),
    .A2(_04958_),
    .Y(_04964_),
    .B1(_04934_));
 sg13g2_o21ai_1 _21461_ (.B1(\top_ihp.wb_spi.bits_left[5] ),
    .Y(_04965_),
    .A1(_04931_),
    .A2(_04964_));
 sg13g2_o21ai_1 _21462_ (.B1(_04965_),
    .Y(_02773_),
    .A1(net206),
    .A2(_04963_));
 sg13g2_buf_1 _21463_ (.A(_08193_),
    .X(_04966_));
 sg13g2_buf_1 _21464_ (.A(net779),
    .X(_04967_));
 sg13g2_nor2_1 _21465_ (.A(net1018),
    .B(_00185_),
    .Y(_04968_));
 sg13g2_a22oi_1 _21466_ (.Y(_04969_),
    .B1(net759),
    .B2(_04968_),
    .A2(net5),
    .A1(net979));
 sg13g2_nand2_1 _21467_ (.Y(_04970_),
    .A(\top_ihp.wb_dati_spi[0] ),
    .B(net444));
 sg13g2_o21ai_1 _21468_ (.B1(_04970_),
    .Y(_02774_),
    .A1(net206),
    .A2(_04969_));
 sg13g2_buf_1 _21469_ (.A(_08193_),
    .X(_04971_));
 sg13g2_nor2b_1 _21470_ (.A(net980),
    .B_N(_04113_),
    .Y(_04972_));
 sg13g2_a22oi_1 _21471_ (.Y(_04973_),
    .B1(net759),
    .B2(_04972_),
    .A2(\top_ihp.wb_dati_spi[9] ),
    .A1(_04971_));
 sg13g2_nand2_1 _21472_ (.Y(_04974_),
    .A(\top_ihp.wb_dati_spi[10] ),
    .B(net444));
 sg13g2_o21ai_1 _21473_ (.B1(_04974_),
    .Y(_02775_),
    .A1(net206),
    .A2(_04973_));
 sg13g2_nor2b_1 _21474_ (.A(net980),
    .B_N(_04115_),
    .Y(_04975_));
 sg13g2_a22oi_1 _21475_ (.Y(_04976_),
    .B1(net759),
    .B2(_04975_),
    .A2(\top_ihp.wb_dati_spi[10] ),
    .A1(_04971_));
 sg13g2_nand2_1 _21476_ (.Y(_04977_),
    .A(\top_ihp.wb_dati_spi[11] ),
    .B(net444));
 sg13g2_o21ai_1 _21477_ (.B1(_04977_),
    .Y(_02776_),
    .A1(net206),
    .A2(_04976_));
 sg13g2_nor2b_1 _21478_ (.A(net980),
    .B_N(_04117_),
    .Y(_04978_));
 sg13g2_a22oi_1 _21479_ (.Y(_04979_),
    .B1(net759),
    .B2(_04978_),
    .A2(\top_ihp.wb_dati_spi[11] ),
    .A1(net978));
 sg13g2_nand2_1 _21480_ (.Y(_04980_),
    .A(\top_ihp.wb_dati_spi[12] ),
    .B(net444));
 sg13g2_o21ai_1 _21481_ (.B1(_04980_),
    .Y(_02777_),
    .A1(net206),
    .A2(_04979_));
 sg13g2_nor2b_1 _21482_ (.A(net980),
    .B_N(_04119_),
    .Y(_04981_));
 sg13g2_a22oi_1 _21483_ (.Y(_04982_),
    .B1(net759),
    .B2(_04981_),
    .A2(\top_ihp.wb_dati_spi[12] ),
    .A1(net978));
 sg13g2_buf_1 _21484_ (.A(_04933_),
    .X(_04983_));
 sg13g2_nand2_1 _21485_ (.Y(_04984_),
    .A(\top_ihp.wb_dati_spi[13] ),
    .B(net442));
 sg13g2_o21ai_1 _21486_ (.B1(_04984_),
    .Y(_02778_),
    .A1(net206),
    .A2(_04982_));
 sg13g2_buf_1 _21487_ (.A(_08193_),
    .X(_04985_));
 sg13g2_nor2b_1 _21488_ (.A(net977),
    .B_N(_04121_),
    .Y(_04986_));
 sg13g2_a22oi_1 _21489_ (.Y(_04987_),
    .B1(net759),
    .B2(_04986_),
    .A2(\top_ihp.wb_dati_spi[13] ),
    .A1(net978));
 sg13g2_nand2_1 _21490_ (.Y(_04988_),
    .A(\top_ihp.wb_dati_spi[14] ),
    .B(net442));
 sg13g2_o21ai_1 _21491_ (.B1(_04988_),
    .Y(_02779_),
    .A1(net206),
    .A2(_04987_));
 sg13g2_nor2b_1 _21492_ (.A(net977),
    .B_N(_04124_),
    .Y(_04989_));
 sg13g2_a22oi_1 _21493_ (.Y(_04990_),
    .B1(net759),
    .B2(_04989_),
    .A2(\top_ihp.wb_dati_spi[14] ),
    .A1(net978));
 sg13g2_nand2_1 _21494_ (.Y(_04991_),
    .A(\top_ihp.wb_dati_spi[15] ),
    .B(net442));
 sg13g2_o21ai_1 _21495_ (.B1(_04991_),
    .Y(_02780_),
    .A1(net206),
    .A2(_04990_));
 sg13g2_buf_1 _21496_ (.A(_04933_),
    .X(_04992_));
 sg13g2_buf_1 _21497_ (.A(_08483_),
    .X(_04993_));
 sg13g2_and3_1 _21498_ (.X(_04994_),
    .A(net1023),
    .B(_08478_),
    .C(_08481_));
 sg13g2_buf_2 _21499_ (.A(_04994_),
    .X(_04995_));
 sg13g2_buf_1 _21500_ (.A(_04995_),
    .X(_04996_));
 sg13g2_inv_1 _21501_ (.Y(_04997_),
    .A(_00185_));
 sg13g2_a22oi_1 _21502_ (.Y(_04998_),
    .B1(net777),
    .B2(_04997_),
    .A2(net778),
    .A1(_04126_));
 sg13g2_nor2_1 _21503_ (.A(net977),
    .B(_04998_),
    .Y(_04999_));
 sg13g2_a21oi_1 _21504_ (.A1(net972),
    .A2(\top_ihp.wb_dati_spi[15] ),
    .Y(_05000_),
    .B1(_04999_));
 sg13g2_nand2_1 _21505_ (.Y(_05001_),
    .A(\top_ihp.wb_dati_spi[16] ),
    .B(_04983_));
 sg13g2_o21ai_1 _21506_ (.B1(_05001_),
    .Y(_02781_),
    .A1(net441),
    .A2(_05000_));
 sg13g2_inv_1 _21507_ (.Y(_05002_),
    .A(_00186_));
 sg13g2_a22oi_1 _21508_ (.Y(_05003_),
    .B1(net777),
    .B2(_05002_),
    .A2(net778),
    .A1(_04128_));
 sg13g2_nor2_1 _21509_ (.A(net977),
    .B(_05003_),
    .Y(_05004_));
 sg13g2_a21oi_1 _21510_ (.A1(net972),
    .A2(\top_ihp.wb_dati_spi[16] ),
    .Y(_05005_),
    .B1(_05004_));
 sg13g2_nand2_1 _21511_ (.Y(_05006_),
    .A(\top_ihp.wb_dati_spi[17] ),
    .B(_04983_));
 sg13g2_o21ai_1 _21512_ (.B1(_05006_),
    .Y(_02782_),
    .A1(net441),
    .A2(_05005_));
 sg13g2_inv_1 _21513_ (.Y(_05007_),
    .A(_00187_));
 sg13g2_a22oi_1 _21514_ (.Y(_05008_),
    .B1(net777),
    .B2(_05007_),
    .A2(net778),
    .A1(_04130_));
 sg13g2_nor2_1 _21515_ (.A(net977),
    .B(_05008_),
    .Y(_05009_));
 sg13g2_a21oi_1 _21516_ (.A1(net972),
    .A2(\top_ihp.wb_dati_spi[17] ),
    .Y(_05010_),
    .B1(_05009_));
 sg13g2_nand2_1 _21517_ (.Y(_05011_),
    .A(\top_ihp.wb_dati_spi[18] ),
    .B(net442));
 sg13g2_o21ai_1 _21518_ (.B1(_05011_),
    .Y(_02783_),
    .A1(net441),
    .A2(_05010_));
 sg13g2_inv_1 _21519_ (.Y(_05012_),
    .A(_00188_));
 sg13g2_a22oi_1 _21520_ (.Y(_05013_),
    .B1(net777),
    .B2(_05012_),
    .A2(net778),
    .A1(_04134_));
 sg13g2_nor2_1 _21521_ (.A(net977),
    .B(_05013_),
    .Y(_05014_));
 sg13g2_a21oi_1 _21522_ (.A1(net972),
    .A2(\top_ihp.wb_dati_spi[18] ),
    .Y(_05015_),
    .B1(_05014_));
 sg13g2_nand2_1 _21523_ (.Y(_05016_),
    .A(\top_ihp.wb_dati_spi[19] ),
    .B(net442));
 sg13g2_o21ai_1 _21524_ (.B1(_05016_),
    .Y(_02784_),
    .A1(net441),
    .A2(_05015_));
 sg13g2_nor2_1 _21525_ (.A(net1018),
    .B(_00186_),
    .Y(_05017_));
 sg13g2_a22oi_1 _21526_ (.Y(_05018_),
    .B1(net759),
    .B2(_05017_),
    .A2(\top_ihp.wb_dati_spi[0] ),
    .A1(net978));
 sg13g2_nand2_1 _21527_ (.Y(_05019_),
    .A(\top_ihp.wb_dati_spi[1] ),
    .B(net442));
 sg13g2_o21ai_1 _21528_ (.B1(_05019_),
    .Y(_02785_),
    .A1(net441),
    .A2(_05018_));
 sg13g2_inv_1 _21529_ (.Y(_05020_),
    .A(_00189_));
 sg13g2_a22oi_1 _21530_ (.Y(_05021_),
    .B1(net777),
    .B2(_05020_),
    .A2(_08483_),
    .A1(_04138_));
 sg13g2_nor2_1 _21531_ (.A(net977),
    .B(_05021_),
    .Y(_05022_));
 sg13g2_a21oi_1 _21532_ (.A1(net972),
    .A2(\top_ihp.wb_dati_spi[19] ),
    .Y(_05023_),
    .B1(_05022_));
 sg13g2_nand2_1 _21533_ (.Y(_05024_),
    .A(\top_ihp.wb_dati_spi[20] ),
    .B(net442));
 sg13g2_o21ai_1 _21534_ (.B1(_05024_),
    .Y(_02786_),
    .A1(net441),
    .A2(_05023_));
 sg13g2_inv_1 _21535_ (.Y(_05025_),
    .A(_00190_));
 sg13g2_a22oi_1 _21536_ (.Y(_05026_),
    .B1(net777),
    .B2(_05025_),
    .A2(_08483_),
    .A1(_04140_));
 sg13g2_nor2_1 _21537_ (.A(net977),
    .B(_05026_),
    .Y(_05027_));
 sg13g2_a21oi_1 _21538_ (.A1(net972),
    .A2(\top_ihp.wb_dati_spi[20] ),
    .Y(_05028_),
    .B1(_05027_));
 sg13g2_nand2_1 _21539_ (.Y(_05029_),
    .A(\top_ihp.wb_dati_spi[21] ),
    .B(net442));
 sg13g2_o21ai_1 _21540_ (.B1(_05029_),
    .Y(_02787_),
    .A1(_04992_),
    .A2(_05028_));
 sg13g2_buf_1 _21541_ (.A(_08193_),
    .X(_05030_));
 sg13g2_inv_1 _21542_ (.Y(_05031_),
    .A(_00191_));
 sg13g2_a22oi_1 _21543_ (.Y(_05032_),
    .B1(_04996_),
    .B2(_05031_),
    .A2(_08483_),
    .A1(_04142_));
 sg13g2_nor2_1 _21544_ (.A(net976),
    .B(_05032_),
    .Y(_05033_));
 sg13g2_a21oi_1 _21545_ (.A1(net972),
    .A2(\top_ihp.wb_dati_spi[21] ),
    .Y(_05034_),
    .B1(_05033_));
 sg13g2_buf_1 _21546_ (.A(_04933_),
    .X(_05035_));
 sg13g2_nand2_1 _21547_ (.Y(_05036_),
    .A(\top_ihp.wb_dati_spi[22] ),
    .B(net440));
 sg13g2_o21ai_1 _21548_ (.B1(_05036_),
    .Y(_02788_),
    .A1(net441),
    .A2(_05034_));
 sg13g2_inv_1 _21549_ (.Y(_05037_),
    .A(_00192_));
 sg13g2_a22oi_1 _21550_ (.Y(_05038_),
    .B1(_04996_),
    .B2(_05037_),
    .A2(_08483_),
    .A1(_04144_));
 sg13g2_nor2_1 _21551_ (.A(net976),
    .B(_05038_),
    .Y(_05039_));
 sg13g2_a21oi_1 _21552_ (.A1(net979),
    .A2(\top_ihp.wb_dati_spi[22] ),
    .Y(_05040_),
    .B1(_05039_));
 sg13g2_nand2_1 _21553_ (.Y(_05041_),
    .A(\top_ihp.wb_dati_spi[23] ),
    .B(net440));
 sg13g2_o21ai_1 _21554_ (.B1(_05041_),
    .Y(_02789_),
    .A1(_04992_),
    .A2(_05040_));
 sg13g2_nand2_1 _21555_ (.Y(_05042_),
    .A(_04148_),
    .B(_04962_));
 sg13g2_a22oi_1 _21556_ (.Y(_05043_),
    .B1(net802),
    .B2(net1050),
    .A2(net777),
    .A1(_04173_));
 sg13g2_a21oi_1 _21557_ (.A1(_05042_),
    .A2(_05043_),
    .Y(_05044_),
    .B1(net976));
 sg13g2_a21oi_1 _21558_ (.A1(net979),
    .A2(\top_ihp.wb_dati_spi[23] ),
    .Y(_05045_),
    .B1(_05044_));
 sg13g2_nand2_1 _21559_ (.Y(_05046_),
    .A(\top_ihp.wb_dati_spi[24] ),
    .B(net440));
 sg13g2_o21ai_1 _21560_ (.B1(_05046_),
    .Y(_02790_),
    .A1(net441),
    .A2(_05045_));
 sg13g2_buf_1 _21561_ (.A(_04933_),
    .X(_05047_));
 sg13g2_nand2_1 _21562_ (.Y(_05048_),
    .A(_04150_),
    .B(net779));
 sg13g2_a22oi_1 _21563_ (.Y(_05049_),
    .B1(net802),
    .B2(_04136_),
    .A2(net777),
    .A1(_04175_));
 sg13g2_a21oi_1 _21564_ (.A1(_05048_),
    .A2(_05049_),
    .Y(_05050_),
    .B1(net976));
 sg13g2_a21oi_1 _21565_ (.A1(net979),
    .A2(\top_ihp.wb_dati_spi[24] ),
    .Y(_05051_),
    .B1(_05050_));
 sg13g2_nand2_1 _21566_ (.Y(_05052_),
    .A(\top_ihp.wb_dati_spi[25] ),
    .B(_05035_));
 sg13g2_o21ai_1 _21567_ (.B1(_05052_),
    .Y(_02791_),
    .A1(_05047_),
    .A2(_05051_));
 sg13g2_nand2_1 _21568_ (.Y(_05053_),
    .A(_04151_),
    .B(_04993_));
 sg13g2_a22oi_1 _21569_ (.Y(_05054_),
    .B1(net802),
    .B2(_04158_),
    .A2(_04995_),
    .A1(_04113_));
 sg13g2_a21oi_1 _21570_ (.A1(_05053_),
    .A2(_05054_),
    .Y(_05055_),
    .B1(net976));
 sg13g2_a21oi_1 _21571_ (.A1(net979),
    .A2(\top_ihp.wb_dati_spi[25] ),
    .Y(_05056_),
    .B1(_05055_));
 sg13g2_nand2_1 _21572_ (.Y(_05057_),
    .A(\top_ihp.wb_dati_spi[26] ),
    .B(_05035_));
 sg13g2_o21ai_1 _21573_ (.B1(_05057_),
    .Y(_02792_),
    .A1(net439),
    .A2(_05056_));
 sg13g2_nand2_1 _21574_ (.Y(_05058_),
    .A(_04153_),
    .B(_04993_));
 sg13g2_a22oi_1 _21575_ (.Y(_05059_),
    .B1(net802),
    .B2(_04163_),
    .A2(_04995_),
    .A1(_04115_));
 sg13g2_a21oi_1 _21576_ (.A1(_05058_),
    .A2(_05059_),
    .Y(_05060_),
    .B1(_05030_));
 sg13g2_a21oi_1 _21577_ (.A1(net979),
    .A2(\top_ihp.wb_dati_spi[26] ),
    .Y(_05061_),
    .B1(_05060_));
 sg13g2_nand2_1 _21578_ (.Y(_05062_),
    .A(\top_ihp.wb_dati_spi[27] ),
    .B(net440));
 sg13g2_o21ai_1 _21579_ (.B1(_05062_),
    .Y(_02793_),
    .A1(net439),
    .A2(_05061_));
 sg13g2_nand2_1 _21580_ (.Y(_05063_),
    .A(_04155_),
    .B(net778));
 sg13g2_a22oi_1 _21581_ (.Y(_05064_),
    .B1(net802),
    .B2(_04165_),
    .A2(_04995_),
    .A1(_04117_));
 sg13g2_a21oi_1 _21582_ (.A1(_05063_),
    .A2(_05064_),
    .Y(_05065_),
    .B1(net976));
 sg13g2_a21oi_1 _21583_ (.A1(_04966_),
    .A2(\top_ihp.wb_dati_spi[27] ),
    .Y(_05066_),
    .B1(_05065_));
 sg13g2_nand2_1 _21584_ (.Y(_05067_),
    .A(\top_ihp.wb_dati_spi[28] ),
    .B(net440));
 sg13g2_o21ai_1 _21585_ (.B1(_05067_),
    .Y(_02794_),
    .A1(_05047_),
    .A2(_05066_));
 sg13g2_nand2_1 _21586_ (.Y(_05068_),
    .A(_04156_),
    .B(net778));
 sg13g2_a22oi_1 _21587_ (.Y(_05069_),
    .B1(net802),
    .B2(_04167_),
    .A2(_04995_),
    .A1(_04119_));
 sg13g2_a21oi_1 _21588_ (.A1(_05068_),
    .A2(_05069_),
    .Y(_05070_),
    .B1(net976));
 sg13g2_a21oi_1 _21589_ (.A1(_04966_),
    .A2(\top_ihp.wb_dati_spi[28] ),
    .Y(_05071_),
    .B1(_05070_));
 sg13g2_nand2_1 _21590_ (.Y(_05072_),
    .A(\top_ihp.wb_dati_spi[29] ),
    .B(net440));
 sg13g2_o21ai_1 _21591_ (.B1(_05072_),
    .Y(_02795_),
    .A1(net439),
    .A2(_05071_));
 sg13g2_nor2_1 _21592_ (.A(net1018),
    .B(_00187_),
    .Y(_05073_));
 sg13g2_a22oi_1 _21593_ (.Y(_05074_),
    .B1(_04967_),
    .B2(_05073_),
    .A2(\top_ihp.wb_dati_spi[1] ),
    .A1(net978));
 sg13g2_nand2_1 _21594_ (.Y(_05075_),
    .A(\top_ihp.wb_dati_spi[2] ),
    .B(net440));
 sg13g2_o21ai_1 _21595_ (.B1(_05075_),
    .Y(_02796_),
    .A1(net439),
    .A2(_05074_));
 sg13g2_nand2_1 _21596_ (.Y(_05076_),
    .A(_04160_),
    .B(net778));
 sg13g2_a22oi_1 _21597_ (.Y(_05077_),
    .B1(net802),
    .B2(_04169_),
    .A2(_04995_),
    .A1(_04121_));
 sg13g2_a21oi_1 _21598_ (.A1(_05076_),
    .A2(_05077_),
    .Y(_05078_),
    .B1(_05030_));
 sg13g2_a21oi_1 _21599_ (.A1(net979),
    .A2(\top_ihp.wb_dati_spi[29] ),
    .Y(_05079_),
    .B1(_05078_));
 sg13g2_nand2_1 _21600_ (.Y(_05080_),
    .A(\top_ihp.wb_dati_spi[30] ),
    .B(net440));
 sg13g2_o21ai_1 _21601_ (.B1(_05080_),
    .Y(_02797_),
    .A1(net439),
    .A2(_05079_));
 sg13g2_nand2_1 _21602_ (.Y(_05081_),
    .A(_04162_),
    .B(net778));
 sg13g2_a22oi_1 _21603_ (.Y(_05082_),
    .B1(_04948_),
    .B2(_04171_),
    .A2(_04995_),
    .A1(_04124_));
 sg13g2_a21oi_1 _21604_ (.A1(_05081_),
    .A2(_05082_),
    .Y(_05083_),
    .B1(net976));
 sg13g2_a21oi_1 _21605_ (.A1(net979),
    .A2(\top_ihp.wb_dati_spi[30] ),
    .Y(_05084_),
    .B1(_05083_));
 sg13g2_nand2_1 _21606_ (.Y(_05085_),
    .A(\top_ihp.wb_dati_spi[31] ),
    .B(net443));
 sg13g2_o21ai_1 _21607_ (.B1(_05085_),
    .Y(_02798_),
    .A1(net439),
    .A2(_05084_));
 sg13g2_nor2_1 _21608_ (.A(net1018),
    .B(_00188_),
    .Y(_05086_));
 sg13g2_a22oi_1 _21609_ (.Y(_05087_),
    .B1(_04967_),
    .B2(_05086_),
    .A2(\top_ihp.wb_dati_spi[2] ),
    .A1(net978));
 sg13g2_nand2_1 _21610_ (.Y(_05088_),
    .A(\top_ihp.wb_dati_spi[3] ),
    .B(net443));
 sg13g2_o21ai_1 _21611_ (.B1(_05088_),
    .Y(_02799_),
    .A1(net439),
    .A2(_05087_));
 sg13g2_nor2_1 _21612_ (.A(net1018),
    .B(_00189_),
    .Y(_05089_));
 sg13g2_a22oi_1 _21613_ (.Y(_05090_),
    .B1(net779),
    .B2(_05089_),
    .A2(\top_ihp.wb_dati_spi[3] ),
    .A1(net978));
 sg13g2_nand2_1 _21614_ (.Y(_05091_),
    .A(\top_ihp.wb_dati_spi[4] ),
    .B(net443));
 sg13g2_o21ai_1 _21615_ (.B1(_05091_),
    .Y(_02800_),
    .A1(net439),
    .A2(_05090_));
 sg13g2_nor2_1 _21616_ (.A(net1018),
    .B(_00190_),
    .Y(_05092_));
 sg13g2_a22oi_1 _21617_ (.Y(_05093_),
    .B1(net779),
    .B2(_05092_),
    .A2(\top_ihp.wb_dati_spi[4] ),
    .A1(net980));
 sg13g2_nand2_1 _21618_ (.Y(_05094_),
    .A(\top_ihp.wb_dati_spi[5] ),
    .B(net443));
 sg13g2_o21ai_1 _21619_ (.B1(_05094_),
    .Y(_02801_),
    .A1(net444),
    .A2(_05093_));
 sg13g2_nor2_1 _21620_ (.A(net1018),
    .B(_00191_),
    .Y(_05095_));
 sg13g2_a22oi_1 _21621_ (.Y(_05096_),
    .B1(net779),
    .B2(_05095_),
    .A2(\top_ihp.wb_dati_spi[5] ),
    .A1(net980));
 sg13g2_nand2_1 _21622_ (.Y(_05097_),
    .A(\top_ihp.wb_dati_spi[6] ),
    .B(_04945_));
 sg13g2_o21ai_1 _21623_ (.B1(_05097_),
    .Y(_02802_),
    .A1(_04937_),
    .A2(_05096_));
 sg13g2_nor2_1 _21624_ (.A(_08194_),
    .B(_00192_),
    .Y(_05098_));
 sg13g2_a22oi_1 _21625_ (.Y(_05099_),
    .B1(net779),
    .B2(_05098_),
    .A2(\top_ihp.wb_dati_spi[6] ),
    .A1(net980));
 sg13g2_nand2_1 _21626_ (.Y(_05100_),
    .A(\top_ihp.wb_dati_spi[7] ),
    .B(net443));
 sg13g2_o21ai_1 _21627_ (.B1(_05100_),
    .Y(_02803_),
    .A1(net444),
    .A2(_05099_));
 sg13g2_nor2b_1 _21628_ (.A(_04985_),
    .B_N(_04173_),
    .Y(_05101_));
 sg13g2_a22oi_1 _21629_ (.Y(_05102_),
    .B1(net779),
    .B2(_05101_),
    .A2(\top_ihp.wb_dati_spi[7] ),
    .A1(_04959_));
 sg13g2_nand2_1 _21630_ (.Y(_05103_),
    .A(\top_ihp.wb_dati_spi[8] ),
    .B(net443));
 sg13g2_o21ai_1 _21631_ (.B1(_05103_),
    .Y(_02804_),
    .A1(net444),
    .A2(_05102_));
 sg13g2_nor2b_1 _21632_ (.A(_04985_),
    .B_N(_04175_),
    .Y(_05104_));
 sg13g2_a22oi_1 _21633_ (.Y(_05105_),
    .B1(net779),
    .B2(_05104_),
    .A2(\top_ihp.wb_dati_spi[8] ),
    .A1(net980));
 sg13g2_nand2_1 _21634_ (.Y(_05106_),
    .A(\top_ihp.wb_dati_spi[9] ),
    .B(net443));
 sg13g2_o21ai_1 _21635_ (.B1(_05106_),
    .Y(_02805_),
    .A1(net444),
    .A2(_05105_));
 sg13g2_nor2_1 _21636_ (.A(net971),
    .B(net974),
    .Y(_05107_));
 sg13g2_nor2_1 _21637_ (.A(net1048),
    .B(net808),
    .Y(_05108_));
 sg13g2_nor2_1 _21638_ (.A(net974),
    .B(net808),
    .Y(_05109_));
 sg13g2_mux2_1 _21639_ (.A0(_05108_),
    .A1(_05109_),
    .S(_08189_),
    .X(_05110_));
 sg13g2_and2_1 _21640_ (.A(_00091_),
    .B(net883),
    .X(_05111_));
 sg13g2_buf_1 _21641_ (.A(_05111_),
    .X(_05112_));
 sg13g2_o21ai_1 _21642_ (.B1(_05112_),
    .Y(_05113_),
    .A1(_05107_),
    .A2(_05110_));
 sg13g2_o21ai_1 _21643_ (.B1(_05113_),
    .Y(_05114_),
    .A1(_08205_),
    .A2(_08218_));
 sg13g2_o21ai_1 _21644_ (.B1(_04934_),
    .Y(_05115_),
    .A1(_05107_),
    .A2(_05110_));
 sg13g2_nor3_1 _21645_ (.A(_05115_),
    .B(_04188_),
    .C(_05112_),
    .Y(_05116_));
 sg13g2_a21o_1 _21646_ (.A2(_05114_),
    .A1(_00319_),
    .B1(_05116_),
    .X(_02806_));
 sg13g2_inv_1 _21647_ (.Y(_05117_),
    .A(_04558_));
 sg13g2_nor3_1 _21648_ (.A(_05115_),
    .B(_05117_),
    .C(_05112_),
    .Y(_05118_));
 sg13g2_a21o_1 _21649_ (.A2(_05114_),
    .A1(_00320_),
    .B1(_05118_),
    .X(_02807_));
 sg13g2_nor3_1 _21650_ (.A(_05115_),
    .B(_04563_),
    .C(_05112_),
    .Y(_05119_));
 sg13g2_a21o_1 _21651_ (.A2(_05114_),
    .A1(_00321_),
    .B1(_05119_),
    .X(_02808_));
 sg13g2_buf_1 _21652_ (.A(\top_ihp.wb_uart.state[1] ),
    .X(_05120_));
 sg13g2_buf_1 _21653_ (.A(\top_ihp.wb_uart.rx_ready ),
    .X(_05121_));
 sg13g2_buf_1 _21654_ (.A(\top_ihp.wb_uart.tx_ready ),
    .X(_05122_));
 sg13g2_inv_1 _21655_ (.Y(_05123_),
    .A(\top_ihp.wb_uart.state[0] ));
 sg13g2_nor2_1 _21656_ (.A(_05120_),
    .B(_05123_),
    .Y(_05124_));
 sg13g2_a22oi_1 _21657_ (.Y(_05125_),
    .B1(_05122_),
    .B2(_05124_),
    .A2(_05121_),
    .A1(_05120_));
 sg13g2_nor2_1 _21658_ (.A(_09490_),
    .B(net1028),
    .Y(_05126_));
 sg13g2_a21oi_1 _21659_ (.A1(_09490_),
    .A2(_05125_),
    .Y(_02809_),
    .B1(_05126_));
 sg13g2_nor2_1 _21660_ (.A(_05123_),
    .B(_05122_),
    .Y(_05127_));
 sg13g2_a21oi_1 _21661_ (.A1(_05123_),
    .A2(_08641_),
    .Y(_05128_),
    .B1(_05127_));
 sg13g2_nand3b_1 _21662_ (.B(\top_ihp.wb_uart.state[0] ),
    .C(_05120_),
    .Y(_05129_),
    .A_N(_05121_));
 sg13g2_o21ai_1 _21663_ (.B1(_05129_),
    .Y(_02810_),
    .A1(_05120_),
    .A2(_05128_));
 sg13g2_nand3_1 _21664_ (.B(net883),
    .C(_08488_),
    .A(_05123_),
    .Y(_05130_));
 sg13g2_nand2b_1 _21665_ (.Y(_05131_),
    .B(_05120_),
    .A_N(_05121_));
 sg13g2_o21ai_1 _21666_ (.B1(_05131_),
    .Y(_02811_),
    .A1(_05120_),
    .A2(_05130_));
 sg13g2_nand3_1 _21667_ (.B(_08490_),
    .C(_08462_),
    .A(net1055),
    .Y(_05132_));
 sg13g2_buf_1 _21668_ (.A(_05132_),
    .X(_05133_));
 sg13g2_xnor2_1 _21669_ (.Y(_05134_),
    .A(_08536_),
    .B(_08532_));
 sg13g2_nor2_1 _21670_ (.A(_05133_),
    .B(_05134_),
    .Y(_02812_));
 sg13g2_inv_1 _21671_ (.Y(_05135_),
    .A(_08538_));
 sg13g2_xnor2_1 _21672_ (.Y(_05136_),
    .A(_05135_),
    .B(_08537_));
 sg13g2_nor2_1 _21673_ (.A(_05133_),
    .B(_05136_),
    .Y(_02813_));
 sg13g2_o21ai_1 _21674_ (.B1(_08539_),
    .Y(_05137_),
    .A1(_05135_),
    .A2(_08537_));
 sg13g2_inv_1 _21675_ (.Y(_05138_),
    .A(_08539_));
 sg13g2_nand4_1 _21676_ (.B(_08538_),
    .C(_05138_),
    .A(_08536_),
    .Y(_05139_),
    .D(_08532_));
 sg13g2_a21oi_1 _21677_ (.A1(_05137_),
    .A2(_05139_),
    .Y(_02814_),
    .B1(_05133_));
 sg13g2_nor2_1 _21678_ (.A(_00183_),
    .B(_08540_),
    .Y(_05140_));
 sg13g2_nand2_1 _21679_ (.Y(_05141_),
    .A(_08532_),
    .B(_05140_));
 sg13g2_xor2_1 _21680_ (.B(_05141_),
    .A(\top_ihp.wb_uart.uart_rx.bit_cnt[3] ),
    .X(_05142_));
 sg13g2_nor2_1 _21681_ (.A(_05133_),
    .B(_05142_),
    .Y(_02815_));
 sg13g2_and2_1 _21682_ (.A(_08528_),
    .B(_08527_),
    .X(_05143_));
 sg13g2_inv_1 _21683_ (.Y(_05144_),
    .A(_05133_));
 sg13g2_nor3_1 _21684_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[8] ),
    .B(_08510_),
    .C(_08516_),
    .Y(_05145_));
 sg13g2_inv_1 _21685_ (.Y(_05146_),
    .A(_08519_));
 sg13g2_nand4_1 _21686_ (.B(_08520_),
    .C(_08522_),
    .A(_05146_),
    .Y(_05147_),
    .D(_08523_));
 sg13g2_nor3_1 _21687_ (.A(_08518_),
    .B(_08529_),
    .C(_05147_),
    .Y(_05148_));
 sg13g2_nand4_1 _21688_ (.B(_05144_),
    .C(_05145_),
    .A(_05143_),
    .Y(_05149_),
    .D(_05148_));
 sg13g2_buf_1 _21689_ (.A(_05149_),
    .X(_05150_));
 sg13g2_nor2_1 _21690_ (.A(_08536_),
    .B(_05150_),
    .Y(_05151_));
 sg13g2_nand3_1 _21691_ (.B(_05138_),
    .C(_05151_),
    .A(_05135_),
    .Y(_05152_));
 sg13g2_nand2_1 _21692_ (.Y(_05153_),
    .A(_00183_),
    .B(_08493_));
 sg13g2_nand2_1 _21693_ (.Y(_05154_),
    .A(\top_ihp.wb_dati_uart[0] ),
    .B(_05152_));
 sg13g2_o21ai_1 _21694_ (.B1(_05154_),
    .Y(_02816_),
    .A1(_05152_),
    .A2(_05153_));
 sg13g2_inv_1 _21695_ (.Y(_05155_),
    .A(_05150_));
 sg13g2_nand2_1 _21696_ (.Y(_05156_),
    .A(_08536_),
    .B(_05155_));
 sg13g2_nor3_1 _21697_ (.A(_08538_),
    .B(_08539_),
    .C(_05156_),
    .Y(_05157_));
 sg13g2_mux2_1 _21698_ (.A0(\top_ihp.wb_dati_uart[1] ),
    .A1(net1072),
    .S(_05157_),
    .X(_02817_));
 sg13g2_nor2_1 _21699_ (.A(_05135_),
    .B(_08539_),
    .Y(_05158_));
 sg13g2_nand2_1 _21700_ (.Y(_05159_),
    .A(_05151_),
    .B(_05158_));
 sg13g2_mux2_1 _21701_ (.A0(net1072),
    .A1(\top_ihp.wb_dati_uart[2] ),
    .S(_05159_),
    .X(_02818_));
 sg13g2_nor2b_1 _21702_ (.A(_05156_),
    .B_N(_05158_),
    .Y(_05160_));
 sg13g2_mux2_1 _21703_ (.A0(\top_ihp.wb_dati_uart[3] ),
    .A1(net1072),
    .S(_05160_),
    .X(_02819_));
 sg13g2_nor2_1 _21704_ (.A(_08536_),
    .B(_08538_),
    .Y(_05161_));
 sg13g2_a22oi_1 _21705_ (.Y(_05162_),
    .B1(_05161_),
    .B2(_08539_),
    .A2(_05158_),
    .A1(_08536_));
 sg13g2_nand2b_1 _21706_ (.Y(_05163_),
    .B(_00183_),
    .A_N(_05162_));
 sg13g2_o21ai_1 _21707_ (.B1(\top_ihp.wb_dati_uart[4] ),
    .Y(_05164_),
    .A1(_05150_),
    .A2(_05163_));
 sg13g2_nand4_1 _21708_ (.B(_08539_),
    .C(_08493_),
    .A(_05135_),
    .Y(_05165_),
    .D(_05151_));
 sg13g2_nand2_1 _21709_ (.Y(_02820_),
    .A(_05164_),
    .B(_05165_));
 sg13g2_nor3_1 _21710_ (.A(_08538_),
    .B(_05138_),
    .C(_05156_),
    .Y(_05166_));
 sg13g2_mux2_1 _21711_ (.A0(\top_ihp.wb_dati_uart[5] ),
    .A1(net1072),
    .S(_05166_),
    .X(_02821_));
 sg13g2_nor3_1 _21712_ (.A(_08536_),
    .B(_08540_),
    .C(_05150_),
    .Y(_05167_));
 sg13g2_mux2_1 _21713_ (.A0(\top_ihp.wb_dati_uart[6] ),
    .A1(net1072),
    .S(_05167_),
    .X(_02822_));
 sg13g2_nor2_1 _21714_ (.A(_08540_),
    .B(_05156_),
    .Y(_05168_));
 sg13g2_mux2_1 _21715_ (.A0(\top_ihp.wb_dati_uart[7] ),
    .A1(net1072),
    .S(_05168_),
    .X(_02823_));
 sg13g2_nand2_1 _21716_ (.Y(_05169_),
    .A(_08462_),
    .B(_08491_));
 sg13g2_a21oi_1 _21717_ (.A1(_05146_),
    .A2(_00092_),
    .Y(_05170_),
    .B1(_08569_));
 sg13g2_a21o_1 _21718_ (.A2(_05170_),
    .A1(_08529_),
    .B1(_05148_),
    .X(_05171_));
 sg13g2_a22oi_1 _21719_ (.Y(_05172_),
    .B1(_05171_),
    .B2(_05143_),
    .A2(_05170_),
    .A1(_05147_));
 sg13g2_nand2_1 _21720_ (.Y(_05173_),
    .A(_08494_),
    .B(_08491_));
 sg13g2_a21oi_1 _21721_ (.A1(_05145_),
    .A2(_05172_),
    .Y(_05174_),
    .B1(_05173_));
 sg13g2_a21o_1 _21722_ (.A2(_05169_),
    .A1(_05121_),
    .B1(_05174_),
    .X(_02824_));
 sg13g2_nand2_2 _21723_ (.Y(_05175_),
    .A(_08639_),
    .B(_08638_));
 sg13g2_xnor2_1 _21724_ (.Y(_05176_),
    .A(_08642_),
    .B(_08676_));
 sg13g2_nor2_1 _21725_ (.A(_05175_),
    .B(_05176_),
    .Y(_02825_));
 sg13g2_nand2_1 _21726_ (.Y(_05177_),
    .A(_08642_),
    .B(_08676_));
 sg13g2_xor2_1 _21727_ (.B(_05177_),
    .A(_08643_),
    .X(_05178_));
 sg13g2_nor2_1 _21728_ (.A(_05175_),
    .B(_05178_),
    .Y(_02826_));
 sg13g2_o21ai_1 _21729_ (.B1(\top_ihp.wb_uart.uart_tx.bit_cnt[2] ),
    .Y(_05179_),
    .A1(_08658_),
    .A2(_08674_));
 sg13g2_nand2_1 _21730_ (.Y(_05180_),
    .A(_08642_),
    .B(_08643_));
 sg13g2_xor2_1 _21731_ (.B(_05180_),
    .A(_00184_),
    .X(_05181_));
 sg13g2_nand2_1 _21732_ (.Y(_05182_),
    .A(_08676_),
    .B(_05181_));
 sg13g2_a21oi_1 _21733_ (.A1(_05179_),
    .A2(_05182_),
    .Y(_02827_),
    .B1(_05175_));
 sg13g2_xor2_1 _21734_ (.B(_08677_),
    .A(\top_ihp.wb_uart.uart_tx.bit_cnt[3] ),
    .X(_05183_));
 sg13g2_nor2_1 _21735_ (.A(_05175_),
    .B(_05183_),
    .Y(_02828_));
 sg13g2_mux2_1 _21736_ (.A0(net1050),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[0] ),
    .S(net532),
    .X(_02829_));
 sg13g2_mux2_1 _21737_ (.A0(_04136_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[1] ),
    .S(net532),
    .X(_02830_));
 sg13g2_mux2_1 _21738_ (.A0(_04158_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[2] ),
    .S(net532),
    .X(_02831_));
 sg13g2_mux2_1 _21739_ (.A0(_04163_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[3] ),
    .S(net532),
    .X(_02832_));
 sg13g2_mux2_1 _21740_ (.A0(_04165_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[4] ),
    .S(net532),
    .X(_02833_));
 sg13g2_mux2_1 _21741_ (.A0(_04167_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[5] ),
    .S(net532),
    .X(_02834_));
 sg13g2_mux2_1 _21742_ (.A0(_04169_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[6] ),
    .S(net532),
    .X(_02835_));
 sg13g2_mux2_1 _21743_ (.A0(_04171_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[7] ),
    .S(_08685_),
    .X(_02836_));
 sg13g2_nand3_1 _21744_ (.B(net837),
    .C(_08488_),
    .A(_08638_),
    .Y(_05184_));
 sg13g2_o21ai_1 _21745_ (.B1(_05184_),
    .Y(_05185_),
    .A1(_08638_),
    .A2(_05122_));
 sg13g2_o21ai_1 _21746_ (.B1(_08639_),
    .Y(_05186_),
    .A1(_05122_),
    .A2(_08681_));
 sg13g2_o21ai_1 _21747_ (.B1(_05186_),
    .Y(_02837_),
    .A1(_08639_),
    .A2(_05185_));
 sg13g2_inv_1 _21748_ (.Y(_05187_),
    .A(\top_ihp.oisc.decoder.decoded[0] ));
 sg13g2_buf_1 _21749_ (.A(_09884_),
    .X(_05188_));
 sg13g2_a221oi_1 _21750_ (.B2(_10390_),
    .C1(_10289_),
    .B1(_10383_),
    .A1(net987),
    .Y(_05189_),
    .A2(_10287_));
 sg13g2_buf_2 _21751_ (.A(_05189_),
    .X(_05190_));
 sg13g2_nor2b_1 _21752_ (.A(_09884_),
    .B_N(_09925_),
    .Y(_05191_));
 sg13g2_buf_2 _21753_ (.A(_05191_),
    .X(_05192_));
 sg13g2_o21ai_1 _21754_ (.B1(_05190_),
    .Y(_05193_),
    .A1(_10429_),
    .A2(_05192_));
 sg13g2_a21o_1 _21755_ (.A2(_09955_),
    .A1(_09950_),
    .B1(net944),
    .X(_05194_));
 sg13g2_or2_1 _21756_ (.X(_05195_),
    .B(_10457_),
    .A(_05194_));
 sg13g2_and2_1 _21757_ (.A(_10383_),
    .B(_10390_),
    .X(_05196_));
 sg13g2_buf_1 _21758_ (.A(_05196_),
    .X(_05197_));
 sg13g2_buf_1 _21759_ (.A(_05197_),
    .X(_05198_));
 sg13g2_nand3_1 _21760_ (.B(_10429_),
    .C(_10457_),
    .A(net737),
    .Y(_05199_));
 sg13g2_o21ai_1 _21761_ (.B1(_05199_),
    .Y(_05200_),
    .A1(_05193_),
    .A2(_05195_));
 sg13g2_nand2b_1 _21762_ (.Y(_05201_),
    .B(_05200_),
    .A_N(_10359_));
 sg13g2_buf_1 _21763_ (.A(_05201_),
    .X(_05202_));
 sg13g2_nand2_1 _21764_ (.Y(_05203_),
    .A(_05190_),
    .B(_05202_));
 sg13g2_or3_1 _21765_ (.A(_10359_),
    .B(_05197_),
    .C(_10457_),
    .X(_05204_));
 sg13g2_buf_1 _21766_ (.A(_05204_),
    .X(_05205_));
 sg13g2_nand4_1 _21767_ (.B(_05197_),
    .C(_10429_),
    .A(_10359_),
    .Y(_05206_),
    .D(_10457_));
 sg13g2_a21oi_2 _21768_ (.B1(_10291_),
    .Y(_05207_),
    .A2(_05206_),
    .A1(_05205_));
 sg13g2_buf_8 _21769_ (.A(_05207_),
    .X(_05208_));
 sg13g2_nor2_2 _21770_ (.A(_09958_),
    .B(net555),
    .Y(_05209_));
 sg13g2_nor3_1 _21771_ (.A(net776),
    .B(_05203_),
    .C(_05209_),
    .Y(_05210_));
 sg13g2_a21o_1 _21772_ (.A2(_10287_),
    .A1(_09788_),
    .B1(_10289_),
    .X(_05211_));
 sg13g2_buf_1 _21773_ (.A(_05211_),
    .X(_05212_));
 sg13g2_nor2_1 _21774_ (.A(_09958_),
    .B(net775),
    .Y(_05213_));
 sg13g2_buf_2 _21775_ (.A(_05213_),
    .X(_05214_));
 sg13g2_nand2_1 _21776_ (.Y(_05215_),
    .A(net765),
    .B(_05214_));
 sg13g2_nor2_1 _21777_ (.A(net805),
    .B(_05207_),
    .Y(_05216_));
 sg13g2_buf_2 _21778_ (.A(_05216_),
    .X(_05217_));
 sg13g2_nor2b_1 _21779_ (.A(_10359_),
    .B_N(_05200_),
    .Y(_05218_));
 sg13g2_buf_8 _21780_ (.A(_05218_),
    .X(_05219_));
 sg13g2_a21o_1 _21781_ (.A2(_05217_),
    .A1(net788),
    .B1(_05219_),
    .X(_05220_));
 sg13g2_nor2_1 _21782_ (.A(_05215_),
    .B(_05220_),
    .Y(_05221_));
 sg13g2_nand2_1 _21783_ (.Y(_05222_),
    .A(net787),
    .B(net786));
 sg13g2_nand2_1 _21784_ (.Y(_05223_),
    .A(net776),
    .B(_09958_));
 sg13g2_nor2_2 _21785_ (.A(net787),
    .B(_05223_),
    .Y(_05224_));
 sg13g2_nor2_1 _21786_ (.A(net555),
    .B(_05224_),
    .Y(_05225_));
 sg13g2_nand2_1 _21787_ (.Y(_05226_),
    .A(net737),
    .B(_10429_));
 sg13g2_buf_2 _21788_ (.A(_05226_),
    .X(_05227_));
 sg13g2_nor2_1 _21789_ (.A(_05212_),
    .B(_05227_),
    .Y(_05228_));
 sg13g2_nand2_1 _21790_ (.Y(_05229_),
    .A(_05219_),
    .B(_05228_));
 sg13g2_a21oi_1 _21791_ (.A1(_05222_),
    .A2(_05225_),
    .Y(_05230_),
    .B1(_05229_));
 sg13g2_nor4_1 _21792_ (.A(net789),
    .B(_05210_),
    .C(_05221_),
    .D(_05230_),
    .Y(_05231_));
 sg13g2_a21oi_1 _21793_ (.A1(_05187_),
    .A2(net769),
    .Y(_00325_),
    .B1(_05231_));
 sg13g2_buf_1 _21794_ (.A(_10291_),
    .X(_05232_));
 sg13g2_inv_1 _21795_ (.Y(_05233_),
    .A(_10430_));
 sg13g2_nor2_1 _21796_ (.A(net765),
    .B(_05233_),
    .Y(_05234_));
 sg13g2_nand2_1 _21797_ (.Y(_05235_),
    .A(net758),
    .B(_05234_));
 sg13g2_nor4_1 _21798_ (.A(net789),
    .B(_05209_),
    .C(_05220_),
    .D(_05235_),
    .Y(_05236_));
 sg13g2_a21o_1 _21799_ (.A2(_08808_),
    .A1(_07958_),
    .B1(_05236_),
    .X(_00326_));
 sg13g2_nand2_1 _21800_ (.Y(_05237_),
    .A(_10291_),
    .B(net737));
 sg13g2_nor2_2 _21801_ (.A(net788),
    .B(net786),
    .Y(_05238_));
 sg13g2_nor3_1 _21802_ (.A(net805),
    .B(net555),
    .C(_05238_),
    .Y(_05239_));
 sg13g2_nor4_1 _21803_ (.A(net789),
    .B(net742),
    .C(_05237_),
    .D(_05239_),
    .Y(_05240_));
 sg13g2_a21o_1 _21804_ (.A2(net768),
    .A1(_08208_),
    .B1(_05240_),
    .X(_00327_));
 sg13g2_inv_1 _21805_ (.Y(_05241_),
    .A(_05215_));
 sg13g2_buf_8 _21806_ (.A(_05202_),
    .X(_05242_));
 sg13g2_a21oi_2 _21807_ (.B1(_05242_),
    .Y(_05243_),
    .A2(_05241_),
    .A1(_05192_));
 sg13g2_or2_1 _21808_ (.X(_05244_),
    .B(_05224_),
    .A(net555));
 sg13g2_xnor2_1 _21809_ (.Y(_05245_),
    .A(net775),
    .B(net737));
 sg13g2_nand3_1 _21810_ (.B(_05244_),
    .C(_05245_),
    .A(net742),
    .Y(_05246_));
 sg13g2_o21ai_1 _21811_ (.B1(net758),
    .Y(_05247_),
    .A1(net776),
    .A2(net765));
 sg13g2_nand2_1 _21812_ (.Y(_05248_),
    .A(_05217_),
    .B(_05247_));
 sg13g2_nor2_1 _21813_ (.A(net765),
    .B(net742),
    .Y(_05249_));
 sg13g2_o21ai_1 _21814_ (.B1(net775),
    .Y(_05250_),
    .A1(net788),
    .A2(_05249_));
 sg13g2_a21oi_1 _21815_ (.A1(_09958_),
    .A2(_05250_),
    .Y(_05251_),
    .B1(net555));
 sg13g2_nor2_1 _21816_ (.A(_05228_),
    .B(_05251_),
    .Y(_05252_));
 sg13g2_o21ai_1 _21817_ (.B1(net737),
    .Y(_05253_),
    .A1(net787),
    .A2(net742));
 sg13g2_a221oi_1 _21818_ (.B2(_05214_),
    .C1(_05219_),
    .B1(_05253_),
    .A1(_05248_),
    .Y(_05254_),
    .A2(_05252_));
 sg13g2_a21oi_1 _21819_ (.A1(_05243_),
    .A2(_05246_),
    .Y(_05255_),
    .B1(_05254_));
 sg13g2_buf_1 _21820_ (.A(net782),
    .X(_05256_));
 sg13g2_mux2_1 _21821_ (.A0(_09703_),
    .A1(_05255_),
    .S(net757),
    .X(_00328_));
 sg13g2_nor2_1 _21822_ (.A(net776),
    .B(net737),
    .Y(_05257_));
 sg13g2_nand2_1 _21823_ (.Y(_05258_),
    .A(_05233_),
    .B(_05257_));
 sg13g2_nor2_1 _21824_ (.A(net775),
    .B(_05234_),
    .Y(_05259_));
 sg13g2_a221oi_1 _21825_ (.B2(_05259_),
    .C1(_05217_),
    .B1(_05258_),
    .A1(net775),
    .Y(_05260_),
    .A2(_05205_));
 sg13g2_nor2_1 _21826_ (.A(net758),
    .B(net737),
    .Y(_05261_));
 sg13g2_o21ai_1 _21827_ (.B1(_05261_),
    .Y(_05262_),
    .A1(net805),
    .A2(net555));
 sg13g2_a21oi_1 _21828_ (.A1(_05235_),
    .A2(_05262_),
    .Y(_05263_),
    .B1(net788));
 sg13g2_o21ai_1 _21829_ (.B1(_05242_),
    .Y(_05264_),
    .A1(_05260_),
    .A2(_05263_));
 sg13g2_nand4_1 _21830_ (.B(_05190_),
    .C(_05192_),
    .A(_05233_),
    .Y(_05265_),
    .D(_05209_));
 sg13g2_o21ai_1 _21831_ (.B1(_05265_),
    .Y(_05266_),
    .A1(_05209_),
    .A2(_05264_));
 sg13g2_mux2_1 _21832_ (.A0(_09676_),
    .A1(_05266_),
    .S(net757),
    .X(_00329_));
 sg13g2_nand2_1 _21833_ (.Y(_05267_),
    .A(net758),
    .B(net742));
 sg13g2_nand2_1 _21834_ (.Y(_05268_),
    .A(net765),
    .B(_05192_));
 sg13g2_o21ai_1 _21835_ (.B1(_05268_),
    .Y(_05269_),
    .A1(_05227_),
    .A2(_05202_));
 sg13g2_nor2_1 _21836_ (.A(net737),
    .B(_05238_),
    .Y(_05270_));
 sg13g2_o21ai_1 _21837_ (.B1(_05219_),
    .Y(_05271_),
    .A1(net787),
    .A2(_05270_));
 sg13g2_nand2_1 _21838_ (.Y(_05272_),
    .A(_05198_),
    .B(net205));
 sg13g2_a22oi_1 _21839_ (.Y(_05273_),
    .B1(_05271_),
    .B2(_05272_),
    .A2(_05269_),
    .A1(net786));
 sg13g2_nand2_1 _21840_ (.Y(_05274_),
    .A(_05244_),
    .B(_05261_));
 sg13g2_o21ai_1 _21841_ (.B1(_05274_),
    .Y(_05275_),
    .A1(_05267_),
    .A2(_05273_));
 sg13g2_mux2_1 _21842_ (.A0(_09689_),
    .A1(_05275_),
    .S(net757),
    .X(_00330_));
 sg13g2_nor2_1 _21843_ (.A(net758),
    .B(_05227_),
    .Y(_05276_));
 sg13g2_o21ai_1 _21844_ (.B1(_05276_),
    .Y(_05277_),
    .A1(net555),
    .A2(_05224_));
 sg13g2_and2_1 _21845_ (.A(_05193_),
    .B(_05277_),
    .X(_05278_));
 sg13g2_nand3_1 _21846_ (.B(_05190_),
    .C(_05224_),
    .A(net742),
    .Y(_05279_));
 sg13g2_a22oi_1 _21847_ (.Y(_05280_),
    .B1(_05279_),
    .B2(_05243_),
    .A2(_05278_),
    .A1(net205));
 sg13g2_nand2_1 _21848_ (.Y(_05281_),
    .A(net782),
    .B(_05280_));
 sg13g2_o21ai_1 _21849_ (.B1(_05281_),
    .Y(_00331_),
    .A1(_09699_),
    .A2(_05256_));
 sg13g2_nor2_1 _21850_ (.A(net758),
    .B(net742),
    .Y(_05282_));
 sg13g2_a221oi_1 _21851_ (.B2(_10390_),
    .C1(_05282_),
    .B1(_10383_),
    .A1(net788),
    .Y(_05283_),
    .A2(net758));
 sg13g2_nor3_1 _21852_ (.A(_05217_),
    .B(_05251_),
    .C(_05283_),
    .Y(_05284_));
 sg13g2_a22oi_1 _21853_ (.Y(_05285_),
    .B1(_05253_),
    .B2(net786),
    .A2(_05238_),
    .A1(net787));
 sg13g2_o21ai_1 _21854_ (.B1(net205),
    .Y(_05286_),
    .A1(net775),
    .A2(_05285_));
 sg13g2_nor2_1 _21855_ (.A(_05284_),
    .B(_05286_),
    .Y(_05287_));
 sg13g2_nor2b_1 _21856_ (.A(_05227_),
    .B_N(_05214_),
    .Y(_05288_));
 sg13g2_nor2_1 _21857_ (.A(net776),
    .B(_09958_),
    .Y(_05289_));
 sg13g2_and2_1 _21858_ (.A(_05190_),
    .B(_05289_),
    .X(_05290_));
 sg13g2_nor3_1 _21859_ (.A(_10291_),
    .B(_05227_),
    .C(_05223_),
    .Y(_05291_));
 sg13g2_o21ai_1 _21860_ (.B1(net805),
    .Y(_05292_),
    .A1(_05290_),
    .A2(_05291_));
 sg13g2_o21ai_1 _21861_ (.B1(_05292_),
    .Y(_05293_),
    .A1(net758),
    .A2(_05206_));
 sg13g2_nor3_1 _21862_ (.A(net205),
    .B(_05288_),
    .C(_05293_),
    .Y(_05294_));
 sg13g2_nor3_1 _21863_ (.A(net789),
    .B(_05287_),
    .C(_05294_),
    .Y(_05295_));
 sg13g2_a21o_1 _21864_ (.A2(net768),
    .A1(\top_ihp.oisc.decoder.decoded[1] ),
    .B1(_05295_),
    .X(_00332_));
 sg13g2_inv_1 _21865_ (.Y(_05296_),
    .A(\top_ihp.oisc.decoder.decoded[2] ));
 sg13g2_nand3_1 _21866_ (.B(net775),
    .C(net765),
    .A(net776),
    .Y(_05297_));
 sg13g2_nand2_1 _21867_ (.Y(_05298_),
    .A(_05237_),
    .B(_05297_));
 sg13g2_o21ai_1 _21868_ (.B1(net775),
    .Y(_05299_),
    .A1(net742),
    .A2(_05205_));
 sg13g2_a22oi_1 _21869_ (.Y(_05300_),
    .B1(_05299_),
    .B2(net788),
    .A2(_05298_),
    .A1(_05233_));
 sg13g2_o21ai_1 _21870_ (.B1(_05214_),
    .Y(_05301_),
    .A1(_05249_),
    .A2(_05257_));
 sg13g2_o21ai_1 _21871_ (.B1(_05301_),
    .Y(_05302_),
    .A1(_05209_),
    .A2(_05300_));
 sg13g2_nor2b_1 _21872_ (.A(_05217_),
    .B_N(_05302_),
    .Y(_05303_));
 sg13g2_nand2_1 _21873_ (.Y(_05304_),
    .A(net787),
    .B(_05238_));
 sg13g2_o21ai_1 _21874_ (.B1(net205),
    .Y(_05305_),
    .A1(_05237_),
    .A2(_05304_));
 sg13g2_a21oi_1 _21875_ (.A1(_05198_),
    .A2(_05289_),
    .Y(_05306_),
    .B1(_05224_));
 sg13g2_o21ai_1 _21876_ (.B1(_05219_),
    .Y(_05307_),
    .A1(_05267_),
    .A2(_05306_));
 sg13g2_o21ai_1 _21877_ (.B1(_05307_),
    .Y(_05308_),
    .A1(_05303_),
    .A2(_05305_));
 sg13g2_nor2_1 _21878_ (.A(_05235_),
    .B(_05225_),
    .Y(_05309_));
 sg13g2_nor2_1 _21879_ (.A(net789),
    .B(_05309_),
    .Y(_05310_));
 sg13g2_a22oi_1 _21880_ (.Y(_00333_),
    .B1(_05308_),
    .B2(_05310_),
    .A2(net769),
    .A1(_05296_));
 sg13g2_inv_1 _21881_ (.Y(_05311_),
    .A(\top_ihp.oisc.decoder.decoded[3] ));
 sg13g2_nor3_1 _21882_ (.A(net787),
    .B(net786),
    .C(_05232_),
    .Y(_05312_));
 sg13g2_a21o_1 _21883_ (.A2(_05214_),
    .A1(net787),
    .B1(_05312_),
    .X(_05313_));
 sg13g2_a221oi_1 _21884_ (.B2(_05188_),
    .C1(_05208_),
    .B1(_05313_),
    .A1(_05192_),
    .Y(_05314_),
    .A2(_05214_));
 sg13g2_nor3_1 _21885_ (.A(_05227_),
    .B(net205),
    .C(_05314_),
    .Y(_05315_));
 sg13g2_mux2_1 _21886_ (.A0(_10392_),
    .A1(net788),
    .S(_05217_),
    .X(_05316_));
 sg13g2_o21ai_1 _21887_ (.B1(_05232_),
    .Y(_05317_),
    .A1(_09958_),
    .A2(_05253_));
 sg13g2_nor3_1 _21888_ (.A(_05219_),
    .B(_05316_),
    .C(_05317_),
    .Y(_05318_));
 sg13g2_o21ai_1 _21889_ (.B1(net782),
    .Y(_05319_),
    .A1(_05315_),
    .A2(_05318_));
 sg13g2_o21ai_1 _21890_ (.B1(_05319_),
    .Y(_00334_),
    .A1(_05311_),
    .A2(net757));
 sg13g2_nor2_1 _21891_ (.A(_05214_),
    .B(_05238_),
    .Y(_05320_));
 sg13g2_a21oi_1 _21892_ (.A1(_05188_),
    .A2(_09917_),
    .Y(_05321_),
    .B1(_05320_));
 sg13g2_o21ai_1 _21893_ (.B1(_05234_),
    .Y(_05322_),
    .A1(net555),
    .A2(_05321_));
 sg13g2_a21oi_1 _21894_ (.A1(_05190_),
    .A2(_05217_),
    .Y(_05323_),
    .B1(_05293_));
 sg13g2_a221oi_1 _21895_ (.B2(net205),
    .C1(_08806_),
    .B1(_05323_),
    .A1(_05243_),
    .Y(_05324_),
    .A2(_05322_));
 sg13g2_a21o_1 _21896_ (.A2(net768),
    .A1(\top_ihp.oisc.decoder.decoded[4] ),
    .B1(_05324_),
    .X(_00335_));
 sg13g2_o21ai_1 _21897_ (.B1(_05203_),
    .Y(_05325_),
    .A1(net205),
    .A2(_05215_));
 sg13g2_nor3_1 _21898_ (.A(_09875_),
    .B(_05219_),
    .C(_05215_),
    .Y(_05326_));
 sg13g2_a221oi_1 _21899_ (.B2(_05192_),
    .C1(_05326_),
    .B1(_05325_),
    .A1(_05219_),
    .Y(_05327_),
    .A2(_05309_));
 sg13g2_nand2_1 _21900_ (.Y(_05328_),
    .A(\top_ihp.oisc.decoder.decoded[5] ),
    .B(net768));
 sg13g2_o21ai_1 _21901_ (.B1(_05328_),
    .Y(_00336_),
    .A1(_08807_),
    .A2(_05327_));
 sg13g2_inv_1 _21902_ (.Y(_05329_),
    .A(_05229_));
 sg13g2_o21ai_1 _21903_ (.B1(_05229_),
    .Y(_05330_),
    .A1(_09875_),
    .A2(_05203_));
 sg13g2_nor4_1 _21904_ (.A(net805),
    .B(net786),
    .C(_05203_),
    .D(_05208_),
    .Y(_05331_));
 sg13g2_a221oi_1 _21905_ (.B2(net786),
    .C1(_05331_),
    .B1(_05330_),
    .A1(_05192_),
    .Y(_05332_),
    .A2(_05329_));
 sg13g2_buf_1 _21906_ (.A(_08806_),
    .X(_05333_));
 sg13g2_nand2_1 _21907_ (.Y(_05334_),
    .A(\top_ihp.oisc.decoder.decoded[6] ),
    .B(net756));
 sg13g2_o21ai_1 _21908_ (.B1(_05334_),
    .Y(_00337_),
    .A1(_08807_),
    .A2(_05332_));
 sg13g2_o21ai_1 _21909_ (.B1(net776),
    .Y(_05335_),
    .A1(net805),
    .A2(_09949_));
 sg13g2_nand3_1 _21910_ (.B(_05190_),
    .C(_05335_),
    .A(net782),
    .Y(_05336_));
 sg13g2_nand2_1 _21911_ (.Y(_05337_),
    .A(\top_ihp.oisc.decoder.decoded[7] ),
    .B(_05333_));
 sg13g2_o21ai_1 _21912_ (.B1(_05337_),
    .Y(_00338_),
    .A1(_05243_),
    .A2(_05336_));
 sg13g2_mux2_1 _21913_ (.A0(_09712_),
    .A1(_09805_),
    .S(_05256_),
    .X(_00339_));
 sg13g2_mux2_1 _21914_ (.A0(_09730_),
    .A1(_09833_),
    .S(net757),
    .X(_00340_));
 sg13g2_nand2_1 _21915_ (.Y(_05338_),
    .A(net1023),
    .B(net756));
 sg13g2_o21ai_1 _21916_ (.B1(_05338_),
    .Y(_00341_),
    .A1(net769),
    .A2(net776));
 sg13g2_nand2_1 _21917_ (.Y(_05339_),
    .A(net945),
    .B(net756));
 sg13g2_o21ai_1 _21918_ (.B1(_05339_),
    .Y(_00342_),
    .A1(net769),
    .A2(net805));
 sg13g2_nand2_1 _21919_ (.Y(_05340_),
    .A(_09793_),
    .B(net756));
 sg13g2_o21ai_1 _21920_ (.B1(_05340_),
    .Y(_00343_),
    .A1(net769),
    .A2(_09958_));
 sg13g2_mux2_1 _21921_ (.A0(\top_ihp.oisc.decoder.instruction[16] ),
    .A1(_09651_),
    .S(net757),
    .X(_00344_));
 sg13g2_nand2_1 _21922_ (.Y(_05341_),
    .A(\top_ihp.oisc.decoder.instruction[17] ),
    .B(net756));
 sg13g2_o21ai_1 _21923_ (.B1(_05341_),
    .Y(_00345_),
    .A1(net769),
    .A2(_10029_));
 sg13g2_mux2_1 _21924_ (.A0(\top_ihp.oisc.decoder.instruction[18] ),
    .A1(_10048_),
    .S(net757),
    .X(_00346_));
 sg13g2_inv_1 _21925_ (.Y(_05342_),
    .A(\top_ihp.oisc.decoder.instruction[19] ));
 sg13g2_or2_1 _21926_ (.X(_05343_),
    .B(_10075_),
    .A(_08804_));
 sg13g2_buf_2 _21927_ (.A(_05343_),
    .X(_05344_));
 sg13g2_o21ai_1 _21928_ (.B1(_05344_),
    .Y(_00347_),
    .A1(_05342_),
    .A2(net757));
 sg13g2_buf_1 _21929_ (.A(net782),
    .X(_05345_));
 sg13g2_mux2_1 _21930_ (.A0(_09681_),
    .A1(_10136_),
    .S(_05345_),
    .X(_00348_));
 sg13g2_mux2_1 _21931_ (.A0(_10087_),
    .A1(_10161_),
    .S(net755),
    .X(_00349_));
 sg13g2_mux2_1 _21932_ (.A0(_10183_),
    .A1(_10179_),
    .S(net755),
    .X(_00350_));
 sg13g2_nand2_1 _21933_ (.Y(_05346_),
    .A(_10196_),
    .B(net756));
 sg13g2_o21ai_1 _21934_ (.B1(_05346_),
    .Y(_00351_),
    .A1(net769),
    .A2(_09777_));
 sg13g2_mux2_1 _21935_ (.A0(_10211_),
    .A1(_09628_),
    .S(net755),
    .X(_00352_));
 sg13g2_mux2_1 _21936_ (.A0(_10231_),
    .A1(_10227_),
    .S(net755),
    .X(_00353_));
 sg13g2_mux2_1 _21937_ (.A0(_10243_),
    .A1(_09812_),
    .S(net755),
    .X(_00354_));
 sg13g2_nand2_1 _21938_ (.Y(_05347_),
    .A(\top_ihp.oisc.decoder.instruction[27] ),
    .B(net756));
 sg13g2_o21ai_1 _21939_ (.B1(_05347_),
    .Y(_00355_),
    .A1(net768),
    .A2(_09841_));
 sg13g2_mux2_1 _21940_ (.A0(\top_ihp.oisc.decoder.instruction[28] ),
    .A1(_09882_),
    .S(net755),
    .X(_00356_));
 sg13g2_mux2_1 _21941_ (.A0(\top_ihp.oisc.decoder.instruction[29] ),
    .A1(_09923_),
    .S(net755),
    .X(_00357_));
 sg13g2_nand2_1 _21942_ (.Y(_05348_),
    .A(\top_ihp.oisc.decoder.instruction[30] ),
    .B(net756));
 sg13g2_o21ai_1 _21943_ (.B1(_05348_),
    .Y(_00358_),
    .A1(net768),
    .A2(_05194_));
 sg13g2_mux2_1 _21944_ (.A0(_09851_),
    .A1(_10339_),
    .S(net755),
    .X(_00359_));
 sg13g2_mux2_1 _21945_ (.A0(_09679_),
    .A1(_10473_),
    .S(_05345_),
    .X(_00360_));
 sg13g2_nand2_1 _21946_ (.Y(_05349_),
    .A(_09740_),
    .B(_05333_));
 sg13g2_o21ai_1 _21947_ (.B1(_05349_),
    .Y(_00361_),
    .A1(_08808_),
    .A2(_09636_));
 sg13g2_nand2_1 _21948_ (.Y(_05350_),
    .A(_09715_),
    .B(net789));
 sg13g2_o21ai_1 _21949_ (.B1(_05350_),
    .Y(_00362_),
    .A1(net768),
    .A2(_10110_));
 sg13g2_nand2_1 _21950_ (.Y(_05351_),
    .A(\top_ihp.oisc.micro_state[1] ),
    .B(_07959_));
 sg13g2_nor2_1 _21951_ (.A(net1052),
    .B(_05351_),
    .Y(_05352_));
 sg13g2_buf_1 _21952_ (.A(_05352_),
    .X(_05353_));
 sg13g2_nand3b_1 _21953_ (.B(_09674_),
    .C(_09682_),
    .Y(_05354_),
    .A_N(_09688_));
 sg13g2_buf_2 _21954_ (.A(_05354_),
    .X(_05355_));
 sg13g2_and2_1 _21955_ (.A(_09590_),
    .B(_05355_),
    .X(_05356_));
 sg13g2_buf_1 _21956_ (.A(_05356_),
    .X(_05357_));
 sg13g2_inv_1 _21957_ (.Y(_05358_),
    .A(_00198_));
 sg13g2_a22oi_1 _21958_ (.Y(_05359_),
    .B1(_05357_),
    .B2(_05358_),
    .A2(net941),
    .A1(_09280_));
 sg13g2_buf_1 _21959_ (.A(_05359_),
    .X(_05360_));
 sg13g2_nand2_1 _21960_ (.Y(_05361_),
    .A(_09065_),
    .B(net941));
 sg13g2_nand3_1 _21961_ (.B(_09681_),
    .C(_05355_),
    .A(net1052),
    .Y(_05362_));
 sg13g2_inv_1 _21962_ (.Y(_05363_),
    .A(_09735_));
 sg13g2_buf_1 _21963_ (.A(_05363_),
    .X(_05364_));
 sg13g2_nor2_1 _21964_ (.A(_09723_),
    .B(_00199_),
    .Y(_05365_));
 sg13g2_and2_1 _21965_ (.A(_05355_),
    .B(_05365_),
    .X(_05366_));
 sg13g2_buf_1 _21966_ (.A(_05366_),
    .X(_05367_));
 sg13g2_nand3_1 _21967_ (.B(_05367_),
    .C(net941),
    .A(net975),
    .Y(_05368_));
 sg13g2_buf_1 _21968_ (.A(_05368_),
    .X(_05369_));
 sg13g2_a221oi_1 _21969_ (.B2(_05362_),
    .C1(_05369_),
    .B1(_05361_),
    .A1(net1047),
    .Y(_05370_),
    .A2(_08802_));
 sg13g2_buf_2 _21970_ (.A(_05370_),
    .X(_05371_));
 sg13g2_and2_1 _21971_ (.A(_05360_),
    .B(_05371_),
    .X(_05372_));
 sg13g2_buf_1 _21972_ (.A(_05372_),
    .X(_05373_));
 sg13g2_buf_1 _21973_ (.A(_09735_),
    .X(_05374_));
 sg13g2_inv_1 _21974_ (.Y(_05375_),
    .A(_00197_));
 sg13g2_a22oi_1 _21975_ (.Y(_05376_),
    .B1(_05357_),
    .B2(_05375_),
    .A2(net941),
    .A1(\top_ihp.oisc.micro_op[14] ));
 sg13g2_buf_2 _21976_ (.A(_05376_),
    .X(_05377_));
 sg13g2_o21ai_1 _21977_ (.B1(_05377_),
    .Y(_05378_),
    .A1(net1017),
    .A2(net856));
 sg13g2_o21ai_1 _21978_ (.B1(_05378_),
    .Y(_05379_),
    .A1(_08805_),
    .A2(_10103_));
 sg13g2_buf_8 _21979_ (.A(_05379_),
    .X(_05380_));
 sg13g2_inv_1 _21980_ (.Y(_05381_),
    .A(_00196_));
 sg13g2_a22oi_1 _21981_ (.Y(_05382_),
    .B1(_05357_),
    .B2(_05381_),
    .A2(net941),
    .A1(\top_ihp.oisc.micro_op[13] ));
 sg13g2_buf_1 _21982_ (.A(_05382_),
    .X(_05383_));
 sg13g2_inv_1 _21983_ (.Y(_05384_),
    .A(_05383_));
 sg13g2_mux2_1 _21984_ (.A0(_09651_),
    .A1(_05384_),
    .S(_08804_),
    .X(_05385_));
 sg13g2_buf_1 _21985_ (.A(_05385_),
    .X(_05386_));
 sg13g2_nor3_1 _21986_ (.A(net1020),
    .B(net754),
    .C(_05386_),
    .Y(_05387_));
 sg13g2_buf_8 _21987_ (.A(_05387_),
    .X(_05388_));
 sg13g2_and2_1 _21988_ (.A(_05373_),
    .B(net729),
    .X(_05389_));
 sg13g2_buf_1 _21989_ (.A(_05389_),
    .X(_05390_));
 sg13g2_nand2_1 _21990_ (.Y(_05391_),
    .A(\top_ihp.oisc.regs[21][0] ),
    .B(_05390_));
 sg13g2_a21o_1 _21991_ (.A2(_08802_),
    .A1(net1047),
    .B1(_05377_),
    .X(_05392_));
 sg13g2_o21ai_1 _21992_ (.B1(_05392_),
    .Y(_05393_),
    .A1(net807),
    .A2(_10029_));
 sg13g2_buf_1 _21993_ (.A(_05393_),
    .X(_05394_));
 sg13g2_o21ai_1 _21994_ (.B1(_05383_),
    .Y(_05395_),
    .A1(net1017),
    .A2(net856));
 sg13g2_o21ai_1 _21995_ (.B1(_05395_),
    .Y(_05396_),
    .A1(_08804_),
    .A2(_09651_));
 sg13g2_buf_1 _21996_ (.A(_05396_),
    .X(_05397_));
 sg13g2_buf_8 _21997_ (.A(_05397_),
    .X(_05398_));
 sg13g2_o21ai_1 _21998_ (.B1(_05360_),
    .Y(_05399_),
    .A1(net1017),
    .A2(net856));
 sg13g2_o21ai_1 _21999_ (.B1(_05399_),
    .Y(_05400_),
    .A1(net807),
    .A2(_10048_));
 sg13g2_buf_2 _22000_ (.A(_05400_),
    .X(_05401_));
 sg13g2_nor4_1 _22001_ (.A(_05374_),
    .B(_05394_),
    .C(_05398_),
    .D(_05401_),
    .Y(_05402_));
 sg13g2_buf_2 _22002_ (.A(_05402_),
    .X(_05403_));
 sg13g2_a22oi_1 _22003_ (.Y(_05404_),
    .B1(_05357_),
    .B2(_09681_),
    .A2(net941),
    .A1(_09065_));
 sg13g2_buf_1 _22004_ (.A(_05404_),
    .X(_05405_));
 sg13g2_nand2_1 _22005_ (.Y(_05406_),
    .A(net807),
    .B(_05405_));
 sg13g2_nand2_1 _22006_ (.Y(_05407_),
    .A(_08796_),
    .B(_04092_));
 sg13g2_nand2_2 _22007_ (.Y(_05408_),
    .A(_09732_),
    .B(net1016));
 sg13g2_nand3_1 _22008_ (.B(_05367_),
    .C(_05408_),
    .A(net807),
    .Y(_05409_));
 sg13g2_buf_1 _22009_ (.A(_05409_),
    .X(_05410_));
 sg13g2_a221oi_1 _22010_ (.B2(_05344_),
    .C1(net1020),
    .B1(_05410_),
    .A1(_05406_),
    .Y(_05411_),
    .A2(_05407_));
 sg13g2_buf_2 _22011_ (.A(_05411_),
    .X(_05412_));
 sg13g2_buf_8 _22012_ (.A(_05412_),
    .X(_05413_));
 sg13g2_nand3_1 _22013_ (.B(_05403_),
    .C(net673),
    .A(\top_ihp.oisc.regs[58][0] ),
    .Y(_05414_));
 sg13g2_buf_1 _22014_ (.A(net975),
    .X(_05415_));
 sg13g2_buf_8 _22015_ (.A(_05386_),
    .X(_05416_));
 sg13g2_nand3_1 _22016_ (.B(net753),
    .C(net751),
    .A(net940),
    .Y(_05417_));
 sg13g2_buf_2 _22017_ (.A(_05417_),
    .X(_05418_));
 sg13g2_inv_1 _22018_ (.Y(_05419_),
    .A(_09280_));
 sg13g2_nand3_1 _22019_ (.B(_05358_),
    .C(_05355_),
    .A(net1052),
    .Y(_05420_));
 sg13g2_o21ai_1 _22020_ (.B1(_05420_),
    .Y(_05421_),
    .A1(_05419_),
    .A2(_05408_));
 sg13g2_buf_1 _22021_ (.A(_05421_),
    .X(_05422_));
 sg13g2_nor2_1 _22022_ (.A(_05405_),
    .B(_05422_),
    .Y(_05423_));
 sg13g2_nand2_1 _22023_ (.Y(_05424_),
    .A(_05355_),
    .B(_05365_));
 sg13g2_nand2_1 _22024_ (.Y(_05425_),
    .A(_05424_),
    .B(net941));
 sg13g2_nor2_1 _22025_ (.A(_04092_),
    .B(_05425_),
    .Y(_05426_));
 sg13g2_a21oi_1 _22026_ (.A1(_05423_),
    .A2(_05426_),
    .Y(_05427_),
    .B1(net984));
 sg13g2_nor2_1 _22027_ (.A(_05418_),
    .B(_05427_),
    .Y(_05428_));
 sg13g2_buf_1 _22028_ (.A(_05428_),
    .X(_05429_));
 sg13g2_buf_8 _22029_ (.A(net554),
    .X(_05430_));
 sg13g2_a21oi_2 _22030_ (.B1(_05369_),
    .Y(_05431_),
    .A2(_08802_),
    .A1(net1047));
 sg13g2_and2_1 _22031_ (.A(_09066_),
    .B(_05431_),
    .X(_05432_));
 sg13g2_buf_2 _22032_ (.A(_05432_),
    .X(_05433_));
 sg13g2_mux2_1 _22033_ (.A0(_10048_),
    .A1(_05422_),
    .S(net807),
    .X(_05434_));
 sg13g2_buf_8 _22034_ (.A(_05434_),
    .X(_05435_));
 sg13g2_nor4_2 _22035_ (.A(_04078_),
    .B(_05380_),
    .C(net752),
    .Y(_05436_),
    .D(_05435_));
 sg13g2_and2_1 _22036_ (.A(_05433_),
    .B(_05436_),
    .X(_05437_));
 sg13g2_buf_2 _22037_ (.A(_05437_),
    .X(_05438_));
 sg13g2_buf_8 _22038_ (.A(_05438_),
    .X(_05439_));
 sg13g2_buf_8 _22039_ (.A(net553),
    .X(_05440_));
 sg13g2_a22oi_1 _22040_ (.Y(_05441_),
    .B1(net437),
    .B2(\top_ihp.oisc.regs[22][0] ),
    .A2(net438),
    .A1(\top_ihp.oisc.regs[7][0] ));
 sg13g2_o21ai_1 _22041_ (.B1(_05362_),
    .Y(_05442_),
    .A1(_09066_),
    .A2(_05408_));
 sg13g2_buf_2 _22042_ (.A(_05442_),
    .X(_05443_));
 sg13g2_a21oi_1 _22043_ (.A1(_07984_),
    .A2(_08802_),
    .Y(_05444_),
    .B1(_05443_));
 sg13g2_nor3_1 _22044_ (.A(net1017),
    .B(_09735_),
    .C(net856),
    .Y(_05445_));
 sg13g2_a22oi_1 _22045_ (.Y(_05446_),
    .B1(_05445_),
    .B2(_08796_),
    .A2(_05444_),
    .A1(net975));
 sg13g2_nand2_1 _22046_ (.Y(_05447_),
    .A(_05424_),
    .B(_05408_));
 sg13g2_o21ai_1 _22047_ (.B1(_05447_),
    .Y(_05448_),
    .A1(_08221_),
    .A2(net856));
 sg13g2_o21ai_1 _22048_ (.B1(_05448_),
    .Y(_05449_),
    .A1(net807),
    .A2(_10075_));
 sg13g2_buf_2 _22049_ (.A(_05449_),
    .X(_05450_));
 sg13g2_nor3_2 _22050_ (.A(net1021),
    .B(_05446_),
    .C(_05450_),
    .Y(_05451_));
 sg13g2_buf_1 _22051_ (.A(_05451_),
    .X(_05452_));
 sg13g2_nor4_2 _22052_ (.A(net984),
    .B(net754),
    .C(_05416_),
    .Y(_05453_),
    .D(_05435_));
 sg13g2_and2_1 _22053_ (.A(net728),
    .B(_05453_),
    .X(_05454_));
 sg13g2_buf_2 _22054_ (.A(_05454_),
    .X(_05455_));
 sg13g2_buf_1 _22055_ (.A(_05455_),
    .X(_05456_));
 sg13g2_nor4_1 _22056_ (.A(net1021),
    .B(net754),
    .C(net752),
    .D(_05401_),
    .Y(_05457_));
 sg13g2_buf_2 _22057_ (.A(_05457_),
    .X(_05458_));
 sg13g2_and2_1 _22058_ (.A(_05371_),
    .B(_05458_),
    .X(_05459_));
 sg13g2_buf_2 _22059_ (.A(_05459_),
    .X(_05460_));
 sg13g2_buf_8 _22060_ (.A(_05460_),
    .X(_05461_));
 sg13g2_a22oi_1 _22061_ (.Y(_05462_),
    .B1(net435),
    .B2(\top_ihp.oisc.regs[31][0] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[36][0] ));
 sg13g2_nand4_1 _22062_ (.B(_05414_),
    .C(_05441_),
    .A(_05391_),
    .Y(_05463_),
    .D(_05462_));
 sg13g2_nand2_1 _22063_ (.Y(_05464_),
    .A(net975),
    .B(net753));
 sg13g2_buf_2 _22064_ (.A(_05464_),
    .X(_05465_));
 sg13g2_nor2_1 _22065_ (.A(net1020),
    .B(net752),
    .Y(_05466_));
 sg13g2_buf_2 _22066_ (.A(_05466_),
    .X(_05467_));
 sg13g2_nor2_1 _22067_ (.A(net1020),
    .B(_05401_),
    .Y(_05468_));
 sg13g2_buf_8 _22068_ (.A(_05468_),
    .X(_05469_));
 sg13g2_nand2_1 _22069_ (.Y(_05470_),
    .A(_09066_),
    .B(_05431_));
 sg13g2_nor4_1 _22070_ (.A(_05465_),
    .B(_05467_),
    .C(net727),
    .D(_05470_),
    .Y(_05471_));
 sg13g2_buf_2 _22071_ (.A(_05471_),
    .X(_05472_));
 sg13g2_buf_8 _22072_ (.A(net552),
    .X(_05473_));
 sg13g2_nor2_1 _22073_ (.A(_09735_),
    .B(net754),
    .Y(_05474_));
 sg13g2_buf_8 _22074_ (.A(_05474_),
    .X(_05475_));
 sg13g2_a21o_1 _22075_ (.A2(_04092_),
    .A1(_08796_),
    .B1(_05444_),
    .X(_05476_));
 sg13g2_buf_2 _22076_ (.A(_05476_),
    .X(_05477_));
 sg13g2_and2_1 _22077_ (.A(net975),
    .B(_05477_),
    .X(_05478_));
 sg13g2_buf_8 _22078_ (.A(_05478_),
    .X(_05479_));
 sg13g2_nand4_1 _22079_ (.B(_05431_),
    .C(_05422_),
    .A(_05415_),
    .Y(_05480_),
    .D(_05383_));
 sg13g2_nor3_2 _22080_ (.A(_05475_),
    .B(net726),
    .C(_05480_),
    .Y(_05481_));
 sg13g2_buf_8 _22081_ (.A(_05481_),
    .X(_05482_));
 sg13g2_buf_1 _22082_ (.A(net551),
    .X(_05483_));
 sg13g2_a22oi_1 _22083_ (.Y(_05484_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[25][0] ),
    .A2(net434),
    .A1(\top_ihp.oisc.regs[20][0] ));
 sg13g2_buf_8 _22084_ (.A(_05467_),
    .X(_05485_));
 sg13g2_buf_1 _22085_ (.A(net672),
    .X(_05486_));
 sg13g2_buf_1 _22086_ (.A(_05373_),
    .X(_05487_));
 sg13g2_buf_8 _22087_ (.A(_05475_),
    .X(_05488_));
 sg13g2_buf_1 _22088_ (.A(net671),
    .X(_05489_));
 sg13g2_nand3_1 _22089_ (.B(_05487_),
    .C(net549),
    .A(\top_ihp.oisc.regs[23][0] ),
    .Y(_05490_));
 sg13g2_buf_8 _22090_ (.A(_05465_),
    .X(_05491_));
 sg13g2_buf_8 _22091_ (.A(net670),
    .X(_05492_));
 sg13g2_nand3_1 _22092_ (.B(_05424_),
    .C(net941),
    .A(net975),
    .Y(_05493_));
 sg13g2_nor4_1 _22093_ (.A(_04092_),
    .B(_05443_),
    .C(_05422_),
    .D(_05493_),
    .Y(_05494_));
 sg13g2_buf_1 _22094_ (.A(_05494_),
    .X(_05495_));
 sg13g2_nand3_1 _22095_ (.B(net548),
    .C(_05495_),
    .A(\top_ihp.oisc.regs[2][0] ),
    .Y(_05496_));
 sg13g2_nand2_1 _22096_ (.Y(_05497_),
    .A(_05490_),
    .B(_05496_));
 sg13g2_and2_1 _22097_ (.A(net729),
    .B(net749),
    .X(_05498_));
 sg13g2_buf_2 _22098_ (.A(_05498_),
    .X(_05499_));
 sg13g2_buf_8 _22099_ (.A(_05499_),
    .X(_05500_));
 sg13g2_buf_8 _22100_ (.A(net432),
    .X(_05501_));
 sg13g2_a22oi_1 _22101_ (.Y(_05502_),
    .B1(net204),
    .B2(\top_ihp.oisc.regs[4][0] ),
    .A2(_05497_),
    .A1(net550));
 sg13g2_a21oi_1 _22102_ (.A1(net754),
    .A2(net752),
    .Y(_05503_),
    .B1(net1020));
 sg13g2_nor2_1 _22103_ (.A(_05427_),
    .B(_05503_),
    .Y(_05504_));
 sg13g2_buf_2 _22104_ (.A(_05504_),
    .X(_05505_));
 sg13g2_buf_8 _22105_ (.A(_05505_),
    .X(_05506_));
 sg13g2_buf_8 _22106_ (.A(net547),
    .X(_05507_));
 sg13g2_nand2_1 _22107_ (.Y(_05508_),
    .A(_09280_),
    .B(_05353_));
 sg13g2_a221oi_1 _22108_ (.B2(_05508_),
    .C1(_05493_),
    .B1(_05420_),
    .A1(_07984_),
    .Y(_05509_),
    .A2(_08802_));
 sg13g2_buf_2 _22109_ (.A(_05509_),
    .X(_05510_));
 sg13g2_nand2_1 _22110_ (.Y(_05511_),
    .A(_05405_),
    .B(_05510_));
 sg13g2_buf_2 _22111_ (.A(_05511_),
    .X(_05512_));
 sg13g2_nor2_1 _22112_ (.A(_05418_),
    .B(net774),
    .Y(_05513_));
 sg13g2_buf_1 _22113_ (.A(_05513_),
    .X(_05514_));
 sg13g2_buf_8 _22114_ (.A(net546),
    .X(_05515_));
 sg13g2_a22oi_1 _22115_ (.Y(_05516_),
    .B1(net430),
    .B2(\top_ihp.oisc.regs[14][0] ),
    .A2(net431),
    .A1(\top_ihp.oisc.regs[1][0] ));
 sg13g2_nand2_1 _22116_ (.Y(_05517_),
    .A(net975),
    .B(net751));
 sg13g2_buf_8 _22117_ (.A(_05517_),
    .X(_05518_));
 sg13g2_buf_8 _22118_ (.A(net725),
    .X(_05519_));
 sg13g2_buf_8 _22119_ (.A(net669),
    .X(_05520_));
 sg13g2_a21o_1 _22120_ (.A2(_05426_),
    .A1(_05423_),
    .B1(net1020),
    .X(_05521_));
 sg13g2_buf_1 _22121_ (.A(_05521_),
    .X(_05522_));
 sg13g2_buf_2 _22122_ (.A(_05522_),
    .X(_05523_));
 sg13g2_nand3_1 _22123_ (.B(net671),
    .C(net724),
    .A(\top_ihp.oisc.regs[5][0] ),
    .Y(_05524_));
 sg13g2_and2_1 _22124_ (.A(_05405_),
    .B(_05510_),
    .X(_05525_));
 sg13g2_buf_1 _22125_ (.A(_05525_),
    .X(_05526_));
 sg13g2_nand3_1 _22126_ (.B(net548),
    .C(_05526_),
    .A(\top_ihp.oisc.regs[8][0] ),
    .Y(_05527_));
 sg13g2_nand2_1 _22127_ (.Y(_05528_),
    .A(_05524_),
    .B(_05527_));
 sg13g2_nor3_2 _22128_ (.A(net670),
    .B(_05479_),
    .C(_05480_),
    .Y(_05529_));
 sg13g2_buf_8 _22129_ (.A(_05529_),
    .X(_05530_));
 sg13g2_buf_8 _22130_ (.A(net429),
    .X(_05531_));
 sg13g2_a22oi_1 _22131_ (.Y(_05532_),
    .B1(_05531_),
    .B2(\top_ihp.oisc.regs[29][0] ),
    .A2(_05528_),
    .A1(net545));
 sg13g2_nand4_1 _22132_ (.B(_05502_),
    .C(_05516_),
    .A(_05484_),
    .Y(_05533_),
    .D(_05532_));
 sg13g2_nand2_1 _22133_ (.Y(_05534_),
    .A(net940),
    .B(_05435_));
 sg13g2_buf_1 _22134_ (.A(_05534_),
    .X(_05535_));
 sg13g2_o21ai_1 _22135_ (.B1(_05433_),
    .Y(_05536_),
    .A1(_09735_),
    .A2(_05377_));
 sg13g2_buf_1 _22136_ (.A(_05536_),
    .X(_05537_));
 sg13g2_nor3_2 _22137_ (.A(net672),
    .B(net723),
    .C(net748),
    .Y(_05538_));
 sg13g2_nor2_1 _22138_ (.A(_09065_),
    .B(_05369_),
    .Y(_05539_));
 sg13g2_nand4_1 _22139_ (.B(_08805_),
    .C(_05378_),
    .A(net940),
    .Y(_05540_),
    .D(_05539_));
 sg13g2_nor4_1 _22140_ (.A(net984),
    .B(net751),
    .C(_05401_),
    .D(_05540_),
    .Y(_05541_));
 sg13g2_buf_1 _22141_ (.A(_05541_),
    .X(_05542_));
 sg13g2_buf_1 _22142_ (.A(_05542_),
    .X(_05543_));
 sg13g2_a22oi_1 _22143_ (.Y(_05544_),
    .B1(net668),
    .B2(\top_ihp.oisc.regs[28][0] ),
    .A2(_05538_),
    .A1(\top_ihp.oisc.regs[24][0] ));
 sg13g2_nor3_2 _22144_ (.A(_04078_),
    .B(net752),
    .C(_05435_),
    .Y(_05545_));
 sg13g2_nor2b_1 _22145_ (.A(net748),
    .B_N(_05545_),
    .Y(_05546_));
 sg13g2_buf_2 _22146_ (.A(_05546_),
    .X(_05547_));
 sg13g2_buf_8 _22147_ (.A(_05547_),
    .X(_05548_));
 sg13g2_nand3_1 _22148_ (.B(_05360_),
    .C(_05377_),
    .A(_05431_),
    .Y(_05549_));
 sg13g2_nor3_2 _22149_ (.A(net725),
    .B(net726),
    .C(_05549_),
    .Y(_05550_));
 sg13g2_buf_8 _22150_ (.A(_05550_),
    .X(_05551_));
 sg13g2_a22oi_1 _22151_ (.Y(_05552_),
    .B1(net543),
    .B2(\top_ihp.oisc.regs[19][0] ),
    .A2(_05548_),
    .A1(\top_ihp.oisc.regs[18][0] ));
 sg13g2_nand3_1 _22152_ (.B(net754),
    .C(net751),
    .A(net940),
    .Y(_05553_));
 sg13g2_buf_2 _22153_ (.A(_05553_),
    .X(_05554_));
 sg13g2_nor2_1 _22154_ (.A(_05554_),
    .B(_05427_),
    .Y(_05555_));
 sg13g2_buf_2 _22155_ (.A(_05555_),
    .X(_05556_));
 sg13g2_nand2_1 _22156_ (.Y(_05557_),
    .A(_05383_),
    .B(_05510_));
 sg13g2_nor3_1 _22157_ (.A(_05465_),
    .B(net726),
    .C(_05557_),
    .Y(_05558_));
 sg13g2_buf_2 _22158_ (.A(_05558_),
    .X(_05559_));
 sg13g2_a22oi_1 _22159_ (.Y(_05560_),
    .B1(_05559_),
    .B2(\top_ihp.oisc.regs[13][0] ),
    .A2(_05556_),
    .A1(\top_ihp.oisc.regs[3][0] ));
 sg13g2_nor3_1 _22160_ (.A(_05475_),
    .B(net726),
    .C(_05557_),
    .Y(_05561_));
 sg13g2_buf_2 _22161_ (.A(_05561_),
    .X(_05562_));
 sg13g2_or4_1 _22162_ (.A(_04092_),
    .B(_05443_),
    .C(_05422_),
    .D(_05493_),
    .X(_05563_));
 sg13g2_nor4_1 _22163_ (.A(_04079_),
    .B(net754),
    .C(net752),
    .D(_05563_),
    .Y(_05564_));
 sg13g2_buf_2 _22164_ (.A(_05564_),
    .X(_05565_));
 sg13g2_a22oi_1 _22165_ (.Y(_05566_),
    .B1(_05565_),
    .B2(\top_ihp.oisc.regs[6][0] ),
    .A2(_05562_),
    .A1(\top_ihp.oisc.regs[9][0] ));
 sg13g2_nand4_1 _22166_ (.B(_05552_),
    .C(_05560_),
    .A(_05544_),
    .Y(_05567_),
    .D(_05566_));
 sg13g2_nand2_1 _22167_ (.Y(_05568_),
    .A(_05443_),
    .B(_05510_));
 sg13g2_nor2_1 _22168_ (.A(_05418_),
    .B(_05568_),
    .Y(_05569_));
 sg13g2_buf_2 _22169_ (.A(_05569_),
    .X(_05570_));
 sg13g2_buf_8 _22170_ (.A(_05570_),
    .X(_05571_));
 sg13g2_nor3_1 _22171_ (.A(_05467_),
    .B(net726),
    .C(_05549_),
    .Y(_05572_));
 sg13g2_buf_2 _22172_ (.A(_05572_),
    .X(_05573_));
 sg13g2_buf_8 _22173_ (.A(_05573_),
    .X(_05574_));
 sg13g2_a22oi_1 _22174_ (.Y(_05575_),
    .B1(net427),
    .B2(\top_ihp.oisc.regs[17][0] ),
    .A2(net428),
    .A1(\top_ihp.oisc.regs[15][0] ));
 sg13g2_nand2_1 _22175_ (.Y(_05576_),
    .A(_08082_),
    .B(_04086_));
 sg13g2_nor2_1 _22176_ (.A(_05554_),
    .B(_05568_),
    .Y(_05577_));
 sg13g2_buf_2 _22177_ (.A(_05577_),
    .X(_05578_));
 sg13g2_nand2_1 _22178_ (.Y(_05579_),
    .A(\top_ihp.oisc.regs[11][0] ),
    .B(_05578_));
 sg13g2_nand3_1 _22179_ (.B(_05576_),
    .C(_05579_),
    .A(_05575_),
    .Y(_05580_));
 sg13g2_o21ai_1 _22180_ (.B1(_05415_),
    .Y(_05581_),
    .A1(net751),
    .A2(_05435_));
 sg13g2_buf_2 _22181_ (.A(_05581_),
    .X(_05582_));
 sg13g2_nor2_1 _22182_ (.A(net669),
    .B(net723),
    .Y(_05583_));
 sg13g2_a22oi_1 _22183_ (.Y(_05584_),
    .B1(_05583_),
    .B2(\top_ihp.oisc.regs[26][0] ),
    .A2(_05582_),
    .A1(\top_ihp.oisc.regs[16][0] ));
 sg13g2_nor3_1 _22184_ (.A(_05374_),
    .B(net751),
    .C(_05401_),
    .Y(_05585_));
 sg13g2_buf_2 _22185_ (.A(_05585_),
    .X(_05586_));
 sg13g2_and3_1 _22186_ (.X(_05587_),
    .A(net671),
    .B(net673),
    .C(net722));
 sg13g2_buf_1 _22187_ (.A(_05587_),
    .X(_05588_));
 sg13g2_nand2_1 _22188_ (.Y(_05589_),
    .A(\top_ihp.oisc.regs[60][0] ),
    .B(_05588_));
 sg13g2_o21ai_1 _22189_ (.B1(_05589_),
    .Y(_05590_),
    .A1(_05537_),
    .A2(_05584_));
 sg13g2_or3_1 _22190_ (.A(_05567_),
    .B(_05580_),
    .C(_05590_),
    .X(_05591_));
 sg13g2_nor3_1 _22191_ (.A(net1021),
    .B(_05477_),
    .C(_05450_),
    .Y(_05592_));
 sg13g2_buf_2 _22192_ (.A(_05592_),
    .X(_05593_));
 sg13g2_and2_1 _22193_ (.A(_05453_),
    .B(_05593_),
    .X(_05594_));
 sg13g2_buf_2 _22194_ (.A(_05594_),
    .X(_05595_));
 sg13g2_buf_1 _22195_ (.A(_05595_),
    .X(_05596_));
 sg13g2_nor3_1 _22196_ (.A(net1020),
    .B(net754),
    .C(_05397_),
    .Y(_05597_));
 sg13g2_buf_8 _22197_ (.A(_05597_),
    .X(_05598_));
 sg13g2_nor4_2 _22198_ (.A(net984),
    .B(_05401_),
    .C(_05477_),
    .Y(_05599_),
    .D(_05450_));
 sg13g2_and2_1 _22199_ (.A(_05598_),
    .B(_05599_),
    .X(_05600_));
 sg13g2_buf_2 _22200_ (.A(_05600_),
    .X(_05601_));
 sg13g2_buf_2 _22201_ (.A(_05601_),
    .X(_05602_));
 sg13g2_a22oi_1 _22202_ (.Y(_05603_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[47][0] ),
    .A2(net426),
    .A1(\top_ihp.oisc.regs[37][0] ));
 sg13g2_and2_1 _22203_ (.A(_05436_),
    .B(_05593_),
    .X(_05604_));
 sg13g2_buf_2 _22204_ (.A(_05604_),
    .X(_05605_));
 sg13g2_buf_2 _22205_ (.A(_05605_),
    .X(_05606_));
 sg13g2_and2_1 _22206_ (.A(_05371_),
    .B(_05403_),
    .X(_05607_));
 sg13g2_buf_2 _22207_ (.A(_05607_),
    .X(_05608_));
 sg13g2_buf_2 _22208_ (.A(_05608_),
    .X(_05609_));
 sg13g2_a22oi_1 _22209_ (.Y(_05610_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[27][0] ),
    .A2(net424),
    .A1(\top_ihp.oisc.regs[39][0] ));
 sg13g2_nand4_1 _22210_ (.B(_05344_),
    .C(_05477_),
    .A(net975),
    .Y(_05611_),
    .D(_05448_));
 sg13g2_buf_2 _22211_ (.A(_05611_),
    .X(_05612_));
 sg13g2_nor3_1 _22212_ (.A(_05468_),
    .B(_05612_),
    .C(_05503_),
    .Y(_05613_));
 sg13g2_buf_2 _22213_ (.A(_05613_),
    .X(_05614_));
 sg13g2_buf_2 _22214_ (.A(_05614_),
    .X(_05615_));
 sg13g2_nor4_1 _22215_ (.A(_05475_),
    .B(net725),
    .C(net727),
    .D(_05612_),
    .Y(_05616_));
 sg13g2_buf_1 _22216_ (.A(_05616_),
    .X(_05617_));
 sg13g2_buf_8 _22217_ (.A(net542),
    .X(_05618_));
 sg13g2_a22oi_1 _22218_ (.Y(_05619_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[34][0] ),
    .A2(net422),
    .A1(\top_ihp.oisc.regs[32][0] ));
 sg13g2_or2_1 _22219_ (.X(_05620_),
    .B(_05444_),
    .A(net1020));
 sg13g2_a221oi_1 _22220_ (.B2(_05410_),
    .C1(_05620_),
    .B1(_05344_),
    .A1(_08796_),
    .Y(_05621_),
    .A2(net782));
 sg13g2_buf_2 _22221_ (.A(_05621_),
    .X(_05622_));
 sg13g2_nor4_2 _22222_ (.A(net984),
    .B(net753),
    .C(net752),
    .Y(_05623_),
    .D(_05435_));
 sg13g2_and2_1 _22223_ (.A(_05622_),
    .B(_05623_),
    .X(_05624_));
 sg13g2_buf_2 _22224_ (.A(_05624_),
    .X(_05625_));
 sg13g2_buf_1 _22225_ (.A(_05625_),
    .X(_05626_));
 sg13g2_nor4_2 _22226_ (.A(net670),
    .B(_05485_),
    .C(net723),
    .Y(_05627_),
    .D(_05612_));
 sg13g2_buf_8 _22227_ (.A(_05627_),
    .X(_05628_));
 sg13g2_buf_8 _22228_ (.A(_05628_),
    .X(_05629_));
 sg13g2_a22oi_1 _22229_ (.Y(_05630_),
    .B1(net202),
    .B2(\top_ihp.oisc.regs[44][0] ),
    .A2(net420),
    .A1(\top_ihp.oisc.regs[51][0] ));
 sg13g2_nand4_1 _22230_ (.B(_05610_),
    .C(_05619_),
    .A(_05603_),
    .Y(_05631_),
    .D(_05630_));
 sg13g2_nor4_1 _22231_ (.A(_05463_),
    .B(_05533_),
    .C(_05591_),
    .D(_05631_),
    .Y(_05632_));
 sg13g2_nor4_2 _22232_ (.A(net984),
    .B(net753),
    .C(net751),
    .Y(_05633_),
    .D(_05401_));
 sg13g2_and2_1 _22233_ (.A(net728),
    .B(_05633_),
    .X(_05634_));
 sg13g2_buf_1 _22234_ (.A(_05634_),
    .X(_05635_));
 sg13g2_buf_1 _22235_ (.A(_05635_),
    .X(_05636_));
 sg13g2_nand2_1 _22236_ (.Y(_05637_),
    .A(_05344_),
    .B(_05410_));
 sg13g2_nor3_1 _22237_ (.A(net984),
    .B(net753),
    .C(_05477_),
    .Y(_05638_));
 sg13g2_and3_1 _22238_ (.X(_05639_),
    .A(_05637_),
    .B(_05586_),
    .C(_05638_));
 sg13g2_buf_1 _22239_ (.A(_05639_),
    .X(_05640_));
 sg13g2_buf_1 _22240_ (.A(_05640_),
    .X(_05641_));
 sg13g2_a22oi_1 _22241_ (.Y(_05642_),
    .B1(net417),
    .B2(\top_ihp.oisc.regs[57][0] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[40][0] ));
 sg13g2_and2_1 _22242_ (.A(_05403_),
    .B(_05452_),
    .X(_05643_));
 sg13g2_buf_1 _22243_ (.A(_05643_),
    .X(_05644_));
 sg13g2_buf_1 _22244_ (.A(_05644_),
    .X(_05645_));
 sg13g2_and2_1 _22245_ (.A(_05453_),
    .B(_05622_),
    .X(_05646_));
 sg13g2_buf_2 _22246_ (.A(_05646_),
    .X(_05647_));
 sg13g2_buf_1 _22247_ (.A(_05647_),
    .X(_05648_));
 sg13g2_a22oi_1 _22248_ (.Y(_05649_),
    .B1(net415),
    .B2(\top_ihp.oisc.regs[53][0] ),
    .A2(net416),
    .A1(\top_ihp.oisc.regs[42][0] ));
 sg13g2_and2_1 _22249_ (.A(net673),
    .B(_05436_),
    .X(_05650_));
 sg13g2_buf_1 _22250_ (.A(_05650_),
    .X(_05651_));
 sg13g2_buf_1 _22251_ (.A(_05651_),
    .X(_05652_));
 sg13g2_and2_1 _22252_ (.A(_05412_),
    .B(_05633_),
    .X(_05653_));
 sg13g2_buf_4 _22253_ (.X(_05654_),
    .A(_05653_));
 sg13g2_a22oi_1 _22254_ (.Y(_05655_),
    .B1(_05654_),
    .B2(\top_ihp.oisc.regs[56][0] ),
    .A2(net201),
    .A1(\top_ihp.oisc.regs[54][0] ));
 sg13g2_and2_1 _22255_ (.A(net673),
    .B(_05458_),
    .X(_05656_));
 sg13g2_buf_2 _22256_ (.A(_05656_),
    .X(_05657_));
 sg13g2_and2_1 _22257_ (.A(_05433_),
    .B(_05458_),
    .X(_05658_));
 sg13g2_buf_2 _22258_ (.A(_05658_),
    .X(_05659_));
 sg13g2_buf_8 _22259_ (.A(_05659_),
    .X(_05660_));
 sg13g2_a22oi_1 _22260_ (.Y(_05661_),
    .B1(net414),
    .B2(\top_ihp.oisc.regs[30][0] ),
    .A2(_05657_),
    .A1(\top_ihp.oisc.regs[62][0] ));
 sg13g2_nand4_1 _22261_ (.B(_05649_),
    .C(_05655_),
    .A(_05642_),
    .Y(_05662_),
    .D(_05661_));
 sg13g2_and2_1 _22262_ (.A(_05458_),
    .B(_05622_),
    .X(_05663_));
 sg13g2_buf_2 _22263_ (.A(_05663_),
    .X(_05664_));
 sg13g2_buf_8 _22264_ (.A(_05664_),
    .X(_05665_));
 sg13g2_nor3_1 _22265_ (.A(net1021),
    .B(net753),
    .C(net752),
    .Y(_05666_));
 sg13g2_buf_2 _22266_ (.A(_05666_),
    .X(_05667_));
 sg13g2_and2_1 _22267_ (.A(_05667_),
    .B(_05599_),
    .X(_05668_));
 sg13g2_buf_2 _22268_ (.A(_05668_),
    .X(_05669_));
 sg13g2_buf_2 _22269_ (.A(_05669_),
    .X(_05670_));
 sg13g2_a22oi_1 _22270_ (.Y(_05671_),
    .B1(net412),
    .B2(\top_ihp.oisc.regs[43][0] ),
    .A2(net413),
    .A1(\top_ihp.oisc.regs[63][0] ));
 sg13g2_and3_1 _22271_ (.X(_05672_),
    .A(net671),
    .B(net722),
    .C(_05622_));
 sg13g2_buf_1 _22272_ (.A(_05672_),
    .X(_05673_));
 sg13g2_buf_1 _22273_ (.A(_05673_),
    .X(_05674_));
 sg13g2_and2_1 _22274_ (.A(_05413_),
    .B(_05623_),
    .X(_05675_));
 sg13g2_buf_1 _22275_ (.A(_05675_),
    .X(_05676_));
 sg13g2_buf_1 _22276_ (.A(_05676_),
    .X(_05677_));
 sg13g2_a22oi_1 _22277_ (.Y(_05678_),
    .B1(net199),
    .B2(\top_ihp.oisc.regs[50][0] ),
    .A2(net200),
    .A1(\top_ihp.oisc.regs[61][0] ));
 sg13g2_and2_1 _22278_ (.A(net729),
    .B(_05599_),
    .X(_05679_));
 sg13g2_buf_2 _22279_ (.A(_05679_),
    .X(_05680_));
 sg13g2_buf_1 _22280_ (.A(_05680_),
    .X(_05681_));
 sg13g2_and4_1 _22281_ (.A(net672),
    .B(net727),
    .C(_05637_),
    .D(_05638_),
    .X(_05682_));
 sg13g2_buf_2 _22282_ (.A(_05682_),
    .X(_05683_));
 sg13g2_buf_1 _22283_ (.A(_05683_),
    .X(_05684_));
 sg13g2_a22oi_1 _22284_ (.Y(_05685_),
    .B1(_05684_),
    .B2(\top_ihp.oisc.regs[59][0] ),
    .A2(net411),
    .A1(\top_ihp.oisc.regs[45][0] ));
 sg13g2_and2_1 _22285_ (.A(_05436_),
    .B(net728),
    .X(_05686_));
 sg13g2_buf_1 _22286_ (.A(_05686_),
    .X(_05687_));
 sg13g2_a22oi_1 _22287_ (.Y(_05688_),
    .B1(_05667_),
    .B2(\top_ihp.oisc.regs[10][0] ),
    .A2(net729),
    .A1(\top_ihp.oisc.regs[12][0] ));
 sg13g2_nor2_1 _22288_ (.A(net774),
    .B(_05688_),
    .Y(_05689_));
 sg13g2_a21oi_1 _22289_ (.A1(\top_ihp.oisc.regs[38][0] ),
    .A2(_05687_),
    .Y(_05690_),
    .B1(_05689_));
 sg13g2_nand4_1 _22290_ (.B(_05678_),
    .C(_05685_),
    .A(_05671_),
    .Y(_05691_),
    .D(_05690_));
 sg13g2_o21ai_1 _22291_ (.B1(net940),
    .Y(_05692_),
    .A1(net782),
    .A2(_05425_));
 sg13g2_a21oi_1 _22292_ (.A1(_05517_),
    .A2(net726),
    .Y(_05693_),
    .B1(net721));
 sg13g2_nand2_1 _22293_ (.Y(_05694_),
    .A(net807),
    .B(_05367_));
 sg13g2_a21oi_1 _22294_ (.A1(net940),
    .A2(net753),
    .Y(_05695_),
    .B1(_05408_));
 sg13g2_o21ai_1 _22295_ (.B1(_05344_),
    .Y(_05696_),
    .A1(_05694_),
    .A2(_05695_));
 sg13g2_a221oi_1 _22296_ (.B2(net940),
    .C1(net727),
    .B1(_05696_),
    .A1(_05692_),
    .Y(_05697_),
    .A2(_05693_));
 sg13g2_nor2_1 _22297_ (.A(net984),
    .B(_05450_),
    .Y(_05698_));
 sg13g2_mux2_1 _22298_ (.A0(_05433_),
    .A1(_05692_),
    .S(_05475_),
    .X(_05699_));
 sg13g2_o21ai_1 _22299_ (.B1(_05364_),
    .Y(_05700_),
    .A1(net753),
    .A2(_05386_));
 sg13g2_buf_2 _22300_ (.A(_05700_),
    .X(_05701_));
 sg13g2_nand3_1 _22301_ (.B(_05470_),
    .C(_05701_),
    .A(net726),
    .Y(_05702_));
 sg13g2_o21ai_1 _22302_ (.B1(_05702_),
    .Y(_05703_),
    .A1(_05698_),
    .A2(_05699_));
 sg13g2_a21oi_1 _22303_ (.A1(_05582_),
    .A2(_05451_),
    .Y(_05704_),
    .B1(_05373_));
 sg13g2_or2_1 _22304_ (.X(_05705_),
    .B(_05704_),
    .A(net671));
 sg13g2_and3_1 _22305_ (.X(_05706_),
    .A(_05697_),
    .B(_05703_),
    .C(_05705_));
 sg13g2_buf_8 _22306_ (.A(_05706_),
    .X(_05707_));
 sg13g2_buf_8 _22307_ (.A(_05707_),
    .X(_05708_));
 sg13g2_and2_1 _22308_ (.A(_05633_),
    .B(_05593_),
    .X(_05709_));
 sg13g2_buf_2 _22309_ (.A(_05709_),
    .X(_05710_));
 sg13g2_buf_1 _22310_ (.A(_05710_),
    .X(_05711_));
 sg13g2_and3_1 _22311_ (.X(_05712_),
    .A(_05465_),
    .B(_05412_),
    .C(_05582_));
 sg13g2_buf_2 _22312_ (.A(_05712_),
    .X(_05713_));
 sg13g2_buf_8 _22313_ (.A(_05713_),
    .X(_05714_));
 sg13g2_buf_8 _22314_ (.A(net409),
    .X(_05715_));
 sg13g2_a22oi_1 _22315_ (.Y(_05716_),
    .B1(net197),
    .B2(\top_ihp.oisc.regs[48][0] ),
    .A2(net410),
    .A1(\top_ihp.oisc.regs[41][0] ));
 sg13g2_and2_1 _22316_ (.A(_05593_),
    .B(_05623_),
    .X(_05717_));
 sg13g2_buf_1 _22317_ (.A(_05717_),
    .X(_05718_));
 sg13g2_buf_2 _22318_ (.A(_05718_),
    .X(_05719_));
 sg13g2_and3_1 _22319_ (.X(_05720_),
    .A(net723),
    .B(_05701_),
    .C(_05593_));
 sg13g2_buf_2 _22320_ (.A(_05720_),
    .X(_05721_));
 sg13g2_buf_1 _22321_ (.A(_05721_),
    .X(_05722_));
 sg13g2_a22oi_1 _22322_ (.Y(_05723_),
    .B1(net407),
    .B2(\top_ihp.oisc.regs[33][0] ),
    .A2(net408),
    .A1(\top_ihp.oisc.regs[35][0] ));
 sg13g2_and2_1 _22323_ (.A(net728),
    .B(_05458_),
    .X(_05724_));
 sg13g2_buf_1 _22324_ (.A(_05724_),
    .X(_05725_));
 sg13g2_buf_2 _22325_ (.A(_05725_),
    .X(_05726_));
 sg13g2_and3_1 _22326_ (.X(_05727_),
    .A(_05475_),
    .B(_05412_),
    .C(_05582_));
 sg13g2_buf_2 _22327_ (.A(_05727_),
    .X(_05728_));
 sg13g2_buf_2 _22328_ (.A(_05728_),
    .X(_05729_));
 sg13g2_a22oi_1 _22329_ (.Y(_05730_),
    .B1(_05729_),
    .B2(\top_ihp.oisc.regs[52][0] ),
    .A2(net406),
    .A1(\top_ihp.oisc.regs[46][0] ));
 sg13g2_and3_1 _22330_ (.X(_05731_),
    .A(net723),
    .B(_05701_),
    .C(_05622_));
 sg13g2_buf_1 _22331_ (.A(_05731_),
    .X(_05732_));
 sg13g2_buf_2 _22332_ (.A(_05732_),
    .X(_05733_));
 sg13g2_and4_1 _22333_ (.A(_05475_),
    .B(_05446_),
    .C(_05637_),
    .D(_05545_),
    .X(_05734_));
 sg13g2_buf_2 _22334_ (.A(_05734_),
    .X(_05735_));
 sg13g2_buf_1 _22335_ (.A(_05735_),
    .X(_05736_));
 sg13g2_a22oi_1 _22336_ (.Y(_05737_),
    .B1(net403),
    .B2(\top_ihp.oisc.regs[55][0] ),
    .A2(net404),
    .A1(\top_ihp.oisc.regs[49][0] ));
 sg13g2_nand4_1 _22337_ (.B(_05723_),
    .C(_05730_),
    .A(_05716_),
    .Y(_05738_),
    .D(_05737_));
 sg13g2_nor4_2 _22338_ (.A(_05662_),
    .B(_05691_),
    .C(net63),
    .Y(_05739_),
    .D(_05738_));
 sg13g2_nand3_1 _22339_ (.B(_05703_),
    .C(_05705_),
    .A(_05697_),
    .Y(_05740_));
 sg13g2_buf_8 _22340_ (.A(_05740_),
    .X(_05741_));
 sg13g2_buf_8 _22341_ (.A(_05741_),
    .X(_05742_));
 sg13g2_or3_1 _22342_ (.A(net835),
    .B(_05431_),
    .C(_05614_),
    .X(_05743_));
 sg13g2_buf_8 _22343_ (.A(_05743_),
    .X(_05744_));
 sg13g2_inv_2 _22344_ (.Y(_05745_),
    .A(_05744_));
 sg13g2_buf_1 _22345_ (.A(_05745_),
    .X(_05746_));
 sg13g2_o21ai_1 _22346_ (.B1(net27),
    .Y(_05747_),
    .A1(\top_ihp.oisc.regs[0][0] ),
    .A2(net62));
 sg13g2_a22oi_1 _22347_ (.Y(_00388_),
    .B1(_05747_),
    .B2(_05576_),
    .A2(_05739_),
    .A1(_05632_));
 sg13g2_nor3_2 _22348_ (.A(net1021),
    .B(_05398_),
    .C(_05563_),
    .Y(_05748_));
 sg13g2_and2_1 _22349_ (.A(_05465_),
    .B(_05748_),
    .X(_05749_));
 sg13g2_buf_2 _22350_ (.A(_05749_),
    .X(_05750_));
 sg13g2_a22oi_1 _22351_ (.Y(_05751_),
    .B1(_05750_),
    .B2(\top_ihp.oisc.regs[2][10] ),
    .A2(_05562_),
    .A1(\top_ihp.oisc.regs[9][10] ));
 sg13g2_a22oi_1 _22352_ (.Y(_05752_),
    .B1(net543),
    .B2(\top_ihp.oisc.regs[19][10] ),
    .A2(_05499_),
    .A1(\top_ihp.oisc.regs[4][10] ));
 sg13g2_and2_1 _22353_ (.A(net729),
    .B(_05526_),
    .X(_05753_));
 sg13g2_buf_1 _22354_ (.A(_05753_),
    .X(_05754_));
 sg13g2_a22oi_1 _22355_ (.Y(_05755_),
    .B1(_05754_),
    .B2(\top_ihp.oisc.regs[12][10] ),
    .A2(_05573_),
    .A1(\top_ihp.oisc.regs[17][10] ));
 sg13g2_a22oi_1 _22356_ (.Y(_05756_),
    .B1(_05570_),
    .B2(\top_ihp.oisc.regs[15][10] ),
    .A2(_05529_),
    .A1(\top_ihp.oisc.regs[29][10] ));
 sg13g2_nand4_1 _22357_ (.B(_05752_),
    .C(_05755_),
    .A(_05751_),
    .Y(_05757_),
    .D(_05756_));
 sg13g2_nor3_1 _22358_ (.A(_05467_),
    .B(net727),
    .C(net748),
    .Y(_05758_));
 sg13g2_buf_8 _22359_ (.A(_05758_),
    .X(_05759_));
 sg13g2_and2_1 _22360_ (.A(net729),
    .B(_05522_),
    .X(_05760_));
 sg13g2_buf_4 _22361_ (.X(_05761_),
    .A(_05760_));
 sg13g2_a22oi_1 _22362_ (.Y(_05762_),
    .B1(_05761_),
    .B2(\top_ihp.oisc.regs[5][10] ),
    .A2(_05759_),
    .A1(\top_ihp.oisc.regs[16][10] ));
 sg13g2_a22oi_1 _22363_ (.Y(_05763_),
    .B1(_05578_),
    .B2(\top_ihp.oisc.regs[11][10] ),
    .A2(_05542_),
    .A1(\top_ihp.oisc.regs[28][10] ));
 sg13g2_nor3_1 _22364_ (.A(net725),
    .B(_05534_),
    .C(net748),
    .Y(_05764_));
 sg13g2_buf_4 _22365_ (.X(_05765_),
    .A(_05764_));
 sg13g2_a22oi_1 _22366_ (.Y(_05766_),
    .B1(_05765_),
    .B2(\top_ihp.oisc.regs[26][10] ),
    .A2(_05547_),
    .A1(\top_ihp.oisc.regs[18][10] ));
 sg13g2_a22oi_1 _22367_ (.Y(_05767_),
    .B1(_05481_),
    .B2(\top_ihp.oisc.regs[25][10] ),
    .A2(_05438_),
    .A1(\top_ihp.oisc.regs[22][10] ));
 sg13g2_nand4_1 _22368_ (.B(_05763_),
    .C(_05766_),
    .A(_05762_),
    .Y(_05768_),
    .D(_05767_));
 sg13g2_mux2_1 _22369_ (.A0(\top_ihp.oisc.regs[10][10] ),
    .A1(\top_ihp.oisc.regs[8][10] ),
    .S(net725),
    .X(_05769_));
 sg13g2_buf_8 _22370_ (.A(net670),
    .X(_05770_));
 sg13g2_a22oi_1 _22371_ (.Y(_05771_),
    .B1(_05769_),
    .B2(net541),
    .A2(net721),
    .A1(\top_ihp.oisc.regs[14][10] ));
 sg13g2_nor2_1 _22372_ (.A(net774),
    .B(_05771_),
    .Y(_05772_));
 sg13g2_a22oi_1 _22373_ (.Y(_05773_),
    .B1(_05718_),
    .B2(\top_ihp.oisc.regs[35][10] ),
    .A2(_05625_),
    .A1(\top_ihp.oisc.regs[51][10] ));
 sg13g2_nor3_1 _22374_ (.A(_05467_),
    .B(_05534_),
    .C(net748),
    .Y(_05774_));
 sg13g2_buf_2 _22375_ (.A(_05774_),
    .X(_05775_));
 sg13g2_buf_8 _22376_ (.A(_05775_),
    .X(_05776_));
 sg13g2_nand2_1 _22377_ (.Y(_05777_),
    .A(\top_ihp.oisc.regs[24][10] ),
    .B(net402));
 sg13g2_buf_8 _22378_ (.A(_05556_),
    .X(_05778_));
 sg13g2_a22oi_1 _22379_ (.Y(_05779_),
    .B1(net401),
    .B2(\top_ihp.oisc.regs[3][10] ),
    .A2(net547),
    .A1(\top_ihp.oisc.regs[1][10] ));
 sg13g2_nand3_1 _22380_ (.B(_05777_),
    .C(_05779_),
    .A(_05773_),
    .Y(_05780_));
 sg13g2_or4_1 _22381_ (.A(_05757_),
    .B(_05768_),
    .C(_05772_),
    .D(_05780_),
    .X(_05781_));
 sg13g2_buf_2 _22382_ (.A(_05471_),
    .X(_05782_));
 sg13g2_buf_8 _22383_ (.A(_05664_),
    .X(_05783_));
 sg13g2_buf_8 _22384_ (.A(_05565_),
    .X(_05784_));
 sg13g2_and2_1 _22385_ (.A(\top_ihp.oisc.regs[6][10] ),
    .B(net667),
    .X(_05785_));
 sg13g2_a221oi_1 _22386_ (.B2(\top_ihp.oisc.regs[63][10] ),
    .C1(_05785_),
    .B1(net400),
    .A1(\top_ihp.oisc.regs[20][10] ),
    .Y(_05786_),
    .A2(_05782_));
 sg13g2_buf_1 _22387_ (.A(_05651_),
    .X(_05787_));
 sg13g2_and2_1 _22388_ (.A(_05403_),
    .B(_05412_),
    .X(_05788_));
 sg13g2_buf_1 _22389_ (.A(_05788_),
    .X(_05789_));
 sg13g2_buf_8 _22390_ (.A(_05789_),
    .X(_05790_));
 sg13g2_buf_8 _22391_ (.A(_05790_),
    .X(_05791_));
 sg13g2_a22oi_1 _22392_ (.Y(_05792_),
    .B1(net195),
    .B2(\top_ihp.oisc.regs[58][10] ),
    .A2(net196),
    .A1(\top_ihp.oisc.regs[54][10] ));
 sg13g2_buf_1 _22393_ (.A(_05735_),
    .X(_05793_));
 sg13g2_a22oi_1 _22394_ (.Y(_05794_),
    .B1(net398),
    .B2(\top_ihp.oisc.regs[55][10] ),
    .A2(net424),
    .A1(\top_ihp.oisc.regs[39][10] ));
 sg13g2_buf_2 _22395_ (.A(_05595_),
    .X(_05795_));
 sg13g2_buf_2 _22396_ (.A(_05725_),
    .X(_05796_));
 sg13g2_a22oi_1 _22397_ (.Y(_05797_),
    .B1(_05796_),
    .B2(\top_ihp.oisc.regs[46][10] ),
    .A2(net397),
    .A1(\top_ihp.oisc.regs[37][10] ));
 sg13g2_nand4_1 _22398_ (.B(_05792_),
    .C(_05794_),
    .A(_05786_),
    .Y(_05798_),
    .D(_05797_));
 sg13g2_buf_2 _22399_ (.A(_05676_),
    .X(_05799_));
 sg13g2_buf_2 _22400_ (.A(_05710_),
    .X(_05800_));
 sg13g2_a22oi_1 _22401_ (.Y(_05801_),
    .B1(net395),
    .B2(\top_ihp.oisc.regs[41][10] ),
    .A2(net194),
    .A1(\top_ihp.oisc.regs[50][10] ));
 sg13g2_buf_2 _22402_ (.A(_05680_),
    .X(_05802_));
 sg13g2_and3_1 _22403_ (.X(_05803_),
    .A(net670),
    .B(net673),
    .C(net722));
 sg13g2_buf_2 _22404_ (.A(_05803_),
    .X(_05804_));
 sg13g2_buf_8 _22405_ (.A(_05804_),
    .X(_05805_));
 sg13g2_a22oi_1 _22406_ (.Y(_05806_),
    .B1(net193),
    .B2(\top_ihp.oisc.regs[56][10] ),
    .A2(net394),
    .A1(\top_ihp.oisc.regs[45][10] ));
 sg13g2_nand3_1 _22407_ (.B(_05801_),
    .C(_05806_),
    .A(net62),
    .Y(_05807_));
 sg13g2_nor3_1 _22408_ (.A(_05781_),
    .B(_05798_),
    .C(_05807_),
    .Y(_05808_));
 sg13g2_buf_1 _22409_ (.A(_05644_),
    .X(_05809_));
 sg13g2_buf_2 _22410_ (.A(_05728_),
    .X(_05810_));
 sg13g2_a22oi_1 _22411_ (.Y(_05811_),
    .B1(net392),
    .B2(\top_ihp.oisc.regs[52][10] ),
    .A2(net393),
    .A1(\top_ihp.oisc.regs[42][10] ));
 sg13g2_buf_8 _22412_ (.A(_05657_),
    .X(_05812_));
 sg13g2_a22oi_1 _22413_ (.Y(_05813_),
    .B1(net192),
    .B2(\top_ihp.oisc.regs[62][10] ),
    .A2(_05456_),
    .A1(\top_ihp.oisc.regs[36][10] ));
 sg13g2_buf_8 _22414_ (.A(_05721_),
    .X(_05814_));
 sg13g2_a22oi_1 _22415_ (.Y(_05815_),
    .B1(net391),
    .B2(\top_ihp.oisc.regs[33][10] ),
    .A2(net419),
    .A1(\top_ihp.oisc.regs[44][10] ));
 sg13g2_a22oi_1 _22416_ (.Y(_05816_),
    .B1(net409),
    .B2(\top_ihp.oisc.regs[48][10] ),
    .A2(_05608_),
    .A1(\top_ihp.oisc.regs[27][10] ));
 sg13g2_nand4_1 _22417_ (.B(_05813_),
    .C(_05815_),
    .A(_05811_),
    .Y(_05817_),
    .D(_05816_));
 sg13g2_nand2_1 _22418_ (.Y(_05818_),
    .A(_05360_),
    .B(_05371_));
 sg13g2_nor4_1 _22419_ (.A(net1021),
    .B(_05818_),
    .C(_05377_),
    .D(net751),
    .Y(_05819_));
 sg13g2_buf_2 _22420_ (.A(_05819_),
    .X(_05820_));
 sg13g2_buf_2 _22421_ (.A(_05820_),
    .X(_05821_));
 sg13g2_or4_1 _22422_ (.A(_05369_),
    .B(_05405_),
    .C(_05422_),
    .D(_05377_),
    .X(_05822_));
 sg13g2_nor4_1 _22423_ (.A(net1021),
    .B(net782),
    .C(_05383_),
    .D(_05822_),
    .Y(_05823_));
 sg13g2_buf_2 _22424_ (.A(_05823_),
    .X(_05824_));
 sg13g2_buf_1 _22425_ (.A(_05824_),
    .X(_05825_));
 sg13g2_a22oi_1 _22426_ (.Y(_05826_),
    .B1(net720),
    .B2(\top_ihp.oisc.regs[23][10] ),
    .A2(net666),
    .A1(\top_ihp.oisc.regs[21][10] ));
 sg13g2_nand2_1 _22427_ (.Y(_05827_),
    .A(_08029_),
    .B(net803));
 sg13g2_buf_1 _22428_ (.A(_05559_),
    .X(_05828_));
 sg13g2_a22oi_1 _22429_ (.Y(_05829_),
    .B1(net390),
    .B2(\top_ihp.oisc.regs[13][10] ),
    .A2(net438),
    .A1(\top_ihp.oisc.regs[7][10] ));
 sg13g2_buf_8 _22430_ (.A(_05460_),
    .X(_05830_));
 sg13g2_a22oi_1 _22431_ (.Y(_05831_),
    .B1(net415),
    .B2(\top_ihp.oisc.regs[53][10] ),
    .A2(net389),
    .A1(\top_ihp.oisc.regs[31][10] ));
 sg13g2_nand4_1 _22432_ (.B(_05827_),
    .C(_05829_),
    .A(_05826_),
    .Y(_05832_),
    .D(_05831_));
 sg13g2_buf_2 _22433_ (.A(_05683_),
    .X(_05833_));
 sg13g2_a22oi_1 _22434_ (.Y(_05834_),
    .B1(net191),
    .B2(\top_ihp.oisc.regs[59][10] ),
    .A2(net412),
    .A1(\top_ihp.oisc.regs[43][10] ));
 sg13g2_buf_8 _22435_ (.A(_05659_),
    .X(_05835_));
 sg13g2_buf_1 _22436_ (.A(_05673_),
    .X(_05836_));
 sg13g2_a22oi_1 _22437_ (.Y(_05837_),
    .B1(net190),
    .B2(\top_ihp.oisc.regs[61][10] ),
    .A2(net388),
    .A1(\top_ihp.oisc.regs[30][10] ));
 sg13g2_nand2_1 _22438_ (.Y(_05838_),
    .A(_05834_),
    .B(_05837_));
 sg13g2_buf_2 _22439_ (.A(_05601_),
    .X(_05839_));
 sg13g2_a22oi_1 _22440_ (.Y(_05840_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[34][10] ),
    .A2(net387),
    .A1(\top_ihp.oisc.regs[47][10] ));
 sg13g2_buf_2 _22441_ (.A(_05732_),
    .X(_05841_));
 sg13g2_a22oi_1 _22442_ (.Y(_05842_),
    .B1(net386),
    .B2(\top_ihp.oisc.regs[49][10] ),
    .A2(net422),
    .A1(\top_ihp.oisc.regs[32][10] ));
 sg13g2_buf_1 _22443_ (.A(_05635_),
    .X(_05843_));
 sg13g2_buf_1 _22444_ (.A(_05687_),
    .X(_05844_));
 sg13g2_a22oi_1 _22445_ (.Y(_05845_),
    .B1(net384),
    .B2(\top_ihp.oisc.regs[38][10] ),
    .A2(net385),
    .A1(\top_ihp.oisc.regs[40][10] ));
 sg13g2_and3_1 _22446_ (.X(_05846_),
    .A(net671),
    .B(_05413_),
    .C(net722));
 sg13g2_buf_8 _22447_ (.A(_05846_),
    .X(_05847_));
 sg13g2_buf_1 _22448_ (.A(net383),
    .X(_05848_));
 sg13g2_a22oi_1 _22449_ (.Y(_05849_),
    .B1(net189),
    .B2(\top_ihp.oisc.regs[60][10] ),
    .A2(net417),
    .A1(\top_ihp.oisc.regs[57][10] ));
 sg13g2_nand4_1 _22450_ (.B(_05842_),
    .C(_05845_),
    .A(_05840_),
    .Y(_05850_),
    .D(_05849_));
 sg13g2_nor4_2 _22451_ (.A(_05817_),
    .B(_05832_),
    .C(_05838_),
    .Y(_05851_),
    .D(_05850_));
 sg13g2_inv_1 _22452_ (.Y(_05852_),
    .A(_00214_));
 sg13g2_o21ai_1 _22453_ (.B1(net27),
    .Y(_05853_),
    .A1(_05852_),
    .A2(net62));
 sg13g2_a22oi_1 _22454_ (.Y(_00389_),
    .B1(_05853_),
    .B2(_05827_),
    .A2(_05851_),
    .A1(_05808_));
 sg13g2_buf_2 _22455_ (.A(_05608_),
    .X(_05854_));
 sg13g2_buf_2 _22456_ (.A(_05713_),
    .X(_05855_));
 sg13g2_a22oi_1 _22457_ (.Y(_05856_),
    .B1(net381),
    .B2(\top_ihp.oisc.regs[48][11] ),
    .A2(_05854_),
    .A1(\top_ihp.oisc.regs[27][11] ));
 sg13g2_buf_8 _22458_ (.A(_05578_),
    .X(_05857_));
 sg13g2_a22oi_1 _22459_ (.Y(_05858_),
    .B1(net380),
    .B2(\top_ihp.oisc.regs[11][11] ),
    .A2(_05573_),
    .A1(\top_ihp.oisc.regs[17][11] ));
 sg13g2_a22oi_1 _22460_ (.Y(_05859_),
    .B1(_05500_),
    .B2(\top_ihp.oisc.regs[4][11] ),
    .A2(net803),
    .A1(_08036_));
 sg13g2_and2_1 _22461_ (.A(_05858_),
    .B(_05859_),
    .X(_05860_));
 sg13g2_buf_2 _22462_ (.A(_05680_),
    .X(_05861_));
 sg13g2_a22oi_1 _22463_ (.Y(_05862_),
    .B1(net379),
    .B2(\top_ihp.oisc.regs[45][11] ),
    .A2(net414),
    .A1(\top_ihp.oisc.regs[30][11] ));
 sg13g2_buf_1 _22464_ (.A(_05676_),
    .X(_05863_));
 sg13g2_buf_1 _22465_ (.A(_05687_),
    .X(_05864_));
 sg13g2_a22oi_1 _22466_ (.Y(_05865_),
    .B1(net378),
    .B2(\top_ihp.oisc.regs[38][11] ),
    .A2(net188),
    .A1(\top_ihp.oisc.regs[50][11] ));
 sg13g2_nand4_1 _22467_ (.B(_05860_),
    .C(_05862_),
    .A(_05856_),
    .Y(_05866_),
    .D(_05865_));
 sg13g2_buf_8 _22468_ (.A(_05804_),
    .X(_05867_));
 sg13g2_a22oi_1 _22469_ (.Y(_05868_),
    .B1(net189),
    .B2(\top_ihp.oisc.regs[60][11] ),
    .A2(net187),
    .A1(\top_ihp.oisc.regs[56][11] ));
 sg13g2_buf_1 _22470_ (.A(_05647_),
    .X(_05869_));
 sg13g2_buf_2 _22471_ (.A(_05625_),
    .X(_05870_));
 sg13g2_a22oi_1 _22472_ (.Y(_05871_),
    .B1(net376),
    .B2(\top_ihp.oisc.regs[51][11] ),
    .A2(net377),
    .A1(\top_ihp.oisc.regs[53][11] ));
 sg13g2_buf_1 _22473_ (.A(_05455_),
    .X(_05872_));
 sg13g2_buf_2 _22474_ (.A(_05616_),
    .X(_05873_));
 sg13g2_a22oi_1 _22475_ (.Y(_05874_),
    .B1(net539),
    .B2(\top_ihp.oisc.regs[34][11] ),
    .A2(net375),
    .A1(\top_ihp.oisc.regs[36][11] ));
 sg13g2_buf_1 _22476_ (.A(_05683_),
    .X(_05875_));
 sg13g2_a22oi_1 _22477_ (.Y(_05876_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[39][11] ),
    .A2(net186),
    .A1(\top_ihp.oisc.regs[59][11] ));
 sg13g2_nand4_1 _22478_ (.B(_05871_),
    .C(_05874_),
    .A(_05868_),
    .Y(_05877_),
    .D(_05876_));
 sg13g2_a22oi_1 _22479_ (.Y(_05878_),
    .B1(net401),
    .B2(\top_ihp.oisc.regs[3][11] ),
    .A2(net668),
    .A1(\top_ihp.oisc.regs[28][11] ));
 sg13g2_a22oi_1 _22480_ (.Y(_05879_),
    .B1(net543),
    .B2(\top_ihp.oisc.regs[19][11] ),
    .A2(net554),
    .A1(\top_ihp.oisc.regs[7][11] ));
 sg13g2_a22oi_1 _22481_ (.Y(_05880_),
    .B1(net402),
    .B2(\top_ihp.oisc.regs[24][11] ),
    .A2(net552),
    .A1(\top_ihp.oisc.regs[20][11] ));
 sg13g2_a22oi_1 _22482_ (.Y(_05881_),
    .B1(net544),
    .B2(\top_ihp.oisc.regs[18][11] ),
    .A2(net553),
    .A1(\top_ihp.oisc.regs[22][11] ));
 sg13g2_and4_1 _22483_ (.A(_05878_),
    .B(_05879_),
    .C(_05880_),
    .D(_05881_),
    .X(_05882_));
 sg13g2_buf_8 _22484_ (.A(_05562_),
    .X(_05883_));
 sg13g2_buf_8 _22485_ (.A(net374),
    .X(_05884_));
 sg13g2_buf_2 _22486_ (.A(net667),
    .X(_05885_));
 sg13g2_a22oi_1 _22487_ (.Y(_05886_),
    .B1(net538),
    .B2(\top_ihp.oisc.regs[6][11] ),
    .A2(net185),
    .A1(\top_ihp.oisc.regs[9][11] ));
 sg13g2_buf_1 _22488_ (.A(net547),
    .X(_05887_));
 sg13g2_buf_8 _22489_ (.A(_05754_),
    .X(_05888_));
 sg13g2_buf_8 _22490_ (.A(net372),
    .X(_05889_));
 sg13g2_a22oi_1 _22491_ (.Y(_05890_),
    .B1(net184),
    .B2(\top_ihp.oisc.regs[12][11] ),
    .A2(net373),
    .A1(\top_ihp.oisc.regs[1][11] ));
 sg13g2_nand3_1 _22492_ (.B(_05886_),
    .C(_05890_),
    .A(_05882_),
    .Y(_05891_));
 sg13g2_buf_8 _22493_ (.A(_05759_),
    .X(_05892_));
 sg13g2_buf_8 _22494_ (.A(net371),
    .X(_05893_));
 sg13g2_a22oi_1 _22495_ (.Y(_05894_),
    .B1(net666),
    .B2(\top_ihp.oisc.regs[21][11] ),
    .A2(net183),
    .A1(\top_ihp.oisc.regs[16][11] ));
 sg13g2_buf_8 _22496_ (.A(net429),
    .X(_05895_));
 sg13g2_buf_1 _22497_ (.A(_05571_),
    .X(_05896_));
 sg13g2_a22oi_1 _22498_ (.Y(_05897_),
    .B1(net181),
    .B2(\top_ihp.oisc.regs[15][11] ),
    .A2(net182),
    .A1(\top_ihp.oisc.regs[29][11] ));
 sg13g2_buf_8 _22499_ (.A(_05559_),
    .X(_05898_));
 sg13g2_buf_1 _22500_ (.A(net370),
    .X(_05899_));
 sg13g2_buf_8 _22501_ (.A(_05750_),
    .X(_05900_));
 sg13g2_buf_8 _22502_ (.A(net369),
    .X(_05901_));
 sg13g2_a22oi_1 _22503_ (.Y(_05902_),
    .B1(net179),
    .B2(\top_ihp.oisc.regs[2][11] ),
    .A2(_05899_),
    .A1(\top_ihp.oisc.regs[13][11] ));
 sg13g2_buf_8 _22504_ (.A(net551),
    .X(_05903_));
 sg13g2_nor3_1 _22505_ (.A(_05475_),
    .B(net725),
    .C(_05511_),
    .Y(_05904_));
 sg13g2_buf_1 _22506_ (.A(_05904_),
    .X(_05905_));
 sg13g2_and2_1 _22507_ (.A(\top_ihp.oisc.regs[5][11] ),
    .B(_05761_),
    .X(_05906_));
 sg13g2_a221oi_1 _22508_ (.B2(\top_ihp.oisc.regs[10][11] ),
    .C1(_05906_),
    .B1(net537),
    .A1(\top_ihp.oisc.regs[25][11] ),
    .Y(_05907_),
    .A2(net368));
 sg13g2_nand4_1 _22509_ (.B(_05897_),
    .C(_05902_),
    .A(_05894_),
    .Y(_05908_),
    .D(_05907_));
 sg13g2_nor4_1 _22510_ (.A(_05866_),
    .B(_05877_),
    .C(_05891_),
    .D(_05908_),
    .Y(_05909_));
 sg13g2_nand2_1 _22511_ (.Y(_05910_),
    .A(\top_ihp.oisc.regs[37][11] ),
    .B(net426));
 sg13g2_buf_8 _22512_ (.A(_05765_),
    .X(_05911_));
 sg13g2_nor2_1 _22513_ (.A(_05503_),
    .B(_05511_),
    .Y(_05912_));
 sg13g2_buf_1 _22514_ (.A(_05912_),
    .X(_05913_));
 sg13g2_buf_2 _22515_ (.A(_05913_),
    .X(_05914_));
 sg13g2_a22oi_1 _22516_ (.Y(_05915_),
    .B1(net536),
    .B2(\top_ihp.oisc.regs[8][11] ),
    .A2(net367),
    .A1(\top_ihp.oisc.regs[26][11] ));
 sg13g2_a22oi_1 _22517_ (.Y(_05916_),
    .B1(net720),
    .B2(\top_ihp.oisc.regs[23][11] ),
    .A2(net430),
    .A1(\top_ihp.oisc.regs[14][11] ));
 sg13g2_nand3_1 _22518_ (.B(_05915_),
    .C(_05916_),
    .A(_05910_),
    .Y(_05917_));
 sg13g2_buf_8 _22519_ (.A(_05741_),
    .X(_05918_));
 sg13g2_buf_1 _22520_ (.A(_05732_),
    .X(_05919_));
 sg13g2_a22oi_1 _22521_ (.Y(_05920_),
    .B1(net366),
    .B2(\top_ihp.oisc.regs[49][11] ),
    .A2(net435),
    .A1(\top_ihp.oisc.regs[31][11] ));
 sg13g2_a22oi_1 _22522_ (.Y(_05921_),
    .B1(net387),
    .B2(\top_ihp.oisc.regs[47][11] ),
    .A2(net393),
    .A1(\top_ihp.oisc.regs[42][11] ));
 sg13g2_nand3_1 _22523_ (.B(_05920_),
    .C(_05921_),
    .A(net61),
    .Y(_05922_));
 sg13g2_buf_1 _22524_ (.A(_05651_),
    .X(_05923_));
 sg13g2_buf_8 _22525_ (.A(_05790_),
    .X(_05924_));
 sg13g2_a22oi_1 _22526_ (.Y(_05925_),
    .B1(net177),
    .B2(\top_ihp.oisc.regs[58][11] ),
    .A2(net178),
    .A1(\top_ihp.oisc.regs[54][11] ));
 sg13g2_a22oi_1 _22527_ (.Y(_05926_),
    .B1(net410),
    .B2(\top_ihp.oisc.regs[41][11] ),
    .A2(net417),
    .A1(\top_ihp.oisc.regs[57][11] ));
 sg13g2_buf_1 _22528_ (.A(_05664_),
    .X(_05927_));
 sg13g2_a22oi_1 _22529_ (.Y(_05928_),
    .B1(net365),
    .B2(\top_ihp.oisc.regs[63][11] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[40][11] ));
 sg13g2_buf_2 _22530_ (.A(_05728_),
    .X(_05929_));
 sg13g2_a22oi_1 _22531_ (.Y(_05930_),
    .B1(net364),
    .B2(\top_ihp.oisc.regs[52][11] ),
    .A2(net200),
    .A1(\top_ihp.oisc.regs[61][11] ));
 sg13g2_nand4_1 _22532_ (.B(_05926_),
    .C(_05928_),
    .A(_05925_),
    .Y(_05931_),
    .D(_05930_));
 sg13g2_buf_2 _22533_ (.A(_05614_),
    .X(_05932_));
 sg13g2_a22oi_1 _22534_ (.Y(_05933_),
    .B1(net396),
    .B2(\top_ihp.oisc.regs[46][11] ),
    .A2(net363),
    .A1(\top_ihp.oisc.regs[32][11] ));
 sg13g2_buf_2 _22535_ (.A(_05669_),
    .X(_05934_));
 sg13g2_buf_2 _22536_ (.A(_05718_),
    .X(_05935_));
 sg13g2_a22oi_1 _22537_ (.Y(_05936_),
    .B1(net361),
    .B2(\top_ihp.oisc.regs[35][11] ),
    .A2(_05934_),
    .A1(\top_ihp.oisc.regs[43][11] ));
 sg13g2_buf_2 _22538_ (.A(_05721_),
    .X(_05937_));
 sg13g2_a22oi_1 _22539_ (.Y(_05938_),
    .B1(net403),
    .B2(\top_ihp.oisc.regs[55][11] ),
    .A2(net360),
    .A1(\top_ihp.oisc.regs[33][11] ));
 sg13g2_buf_1 _22540_ (.A(_05657_),
    .X(_05939_));
 sg13g2_a22oi_1 _22541_ (.Y(_05940_),
    .B1(net202),
    .B2(\top_ihp.oisc.regs[44][11] ),
    .A2(net176),
    .A1(\top_ihp.oisc.regs[62][11] ));
 sg13g2_nand4_1 _22542_ (.B(_05936_),
    .C(_05938_),
    .A(_05933_),
    .Y(_05941_),
    .D(_05940_));
 sg13g2_nor4_2 _22543_ (.A(_05917_),
    .B(_05922_),
    .C(_05931_),
    .Y(_05942_),
    .D(_05941_));
 sg13g2_buf_1 _22544_ (.A(net27),
    .X(_05943_));
 sg13g2_buf_8 _22545_ (.A(_05707_),
    .X(_05944_));
 sg13g2_nand2_1 _22546_ (.Y(_05945_),
    .A(_00215_),
    .B(net60));
 sg13g2_a22oi_1 _22547_ (.Y(_05946_),
    .B1(net26),
    .B2(_05945_),
    .A2(net760),
    .A1(_08036_));
 sg13g2_a21oi_1 _22548_ (.A1(_05909_),
    .A2(_05942_),
    .Y(_00390_),
    .B1(_05946_));
 sg13g2_nand2_1 _22549_ (.Y(_05947_),
    .A(\top_ihp.oisc.regs[41][12] ),
    .B(net395));
 sg13g2_a22oi_1 _22550_ (.Y(_05948_),
    .B1(net397),
    .B2(\top_ihp.oisc.regs[37][12] ),
    .A2(net411),
    .A1(\top_ihp.oisc.regs[45][12] ));
 sg13g2_buf_1 _22551_ (.A(_05735_),
    .X(_05949_));
 sg13g2_a22oi_1 _22552_ (.Y(_05950_),
    .B1(net359),
    .B2(\top_ihp.oisc.regs[55][12] ),
    .A2(net406),
    .A1(\top_ihp.oisc.regs[46][12] ));
 sg13g2_buf_2 _22553_ (.A(_05601_),
    .X(_05951_));
 sg13g2_a22oi_1 _22554_ (.Y(_05952_),
    .B1(net358),
    .B2(\top_ihp.oisc.regs[47][12] ),
    .A2(net413),
    .A1(\top_ihp.oisc.regs[63][12] ));
 sg13g2_nand4_1 _22555_ (.B(_05948_),
    .C(_05950_),
    .A(_05947_),
    .Y(_05953_),
    .D(_05952_));
 sg13g2_buf_1 _22556_ (.A(_05455_),
    .X(_05954_));
 sg13g2_a22oi_1 _22557_ (.Y(_05955_),
    .B1(net388),
    .B2(\top_ihp.oisc.regs[30][12] ),
    .A2(net357),
    .A1(\top_ihp.oisc.regs[36][12] ));
 sg13g2_a22oi_1 _22558_ (.Y(_05956_),
    .B1(net197),
    .B2(\top_ihp.oisc.regs[48][12] ),
    .A2(net422),
    .A1(\top_ihp.oisc.regs[32][12] ));
 sg13g2_a22oi_1 _22559_ (.Y(_05957_),
    .B1(net193),
    .B2(\top_ihp.oisc.regs[56][12] ),
    .A2(net198),
    .A1(\top_ihp.oisc.regs[59][12] ));
 sg13g2_a22oi_1 _22560_ (.Y(_05958_),
    .B1(net194),
    .B2(\top_ihp.oisc.regs[50][12] ),
    .A2(net377),
    .A1(\top_ihp.oisc.regs[53][12] ));
 sg13g2_nand4_1 _22561_ (.B(_05956_),
    .C(_05957_),
    .A(_05955_),
    .Y(_05959_),
    .D(_05958_));
 sg13g2_buf_8 _22562_ (.A(_05460_),
    .X(_05960_));
 sg13g2_buf_2 _22563_ (.A(_05625_),
    .X(_05961_));
 sg13g2_a22oi_1 _22564_ (.Y(_05962_),
    .B1(net355),
    .B2(\top_ihp.oisc.regs[51][12] ),
    .A2(net356),
    .A1(\top_ihp.oisc.regs[31][12] ));
 sg13g2_a22oi_1 _22565_ (.Y(_05963_),
    .B1(net189),
    .B2(\top_ihp.oisc.regs[60][12] ),
    .A2(net539),
    .A1(\top_ihp.oisc.regs[34][12] ));
 sg13g2_a22oi_1 _22566_ (.Y(_05964_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[27][12] ),
    .A2(net178),
    .A1(\top_ihp.oisc.regs[54][12] ));
 sg13g2_buf_1 _22567_ (.A(_05673_),
    .X(_05965_));
 sg13g2_buf_2 _22568_ (.A(_05605_),
    .X(_05966_));
 sg13g2_a22oi_1 _22569_ (.Y(_05967_),
    .B1(net354),
    .B2(\top_ihp.oisc.regs[39][12] ),
    .A2(net175),
    .A1(\top_ihp.oisc.regs[61][12] ));
 sg13g2_nand4_1 _22570_ (.B(_05963_),
    .C(_05964_),
    .A(_05962_),
    .Y(_05968_),
    .D(_05967_));
 sg13g2_nor4_1 _22571_ (.A(_05708_),
    .B(_05953_),
    .C(_05959_),
    .D(_05968_),
    .Y(_05969_));
 sg13g2_buf_2 _22572_ (.A(_05824_),
    .X(_05970_));
 sg13g2_and2_1 _22573_ (.A(_08033_),
    .B(net835),
    .X(_05971_));
 sg13g2_a221oi_1 _22574_ (.B2(\top_ihp.oisc.regs[23][12] ),
    .C1(_05971_),
    .B1(net719),
    .A1(\top_ihp.oisc.regs[3][12] ),
    .Y(_05972_),
    .A2(_05556_));
 sg13g2_a22oi_1 _22575_ (.Y(_05973_),
    .B1(net544),
    .B2(\top_ihp.oisc.regs[18][12] ),
    .A2(net553),
    .A1(\top_ihp.oisc.regs[22][12] ));
 sg13g2_a22oi_1 _22576_ (.Y(_05974_),
    .B1(_05482_),
    .B2(\top_ihp.oisc.regs[25][12] ),
    .A2(net554),
    .A1(\top_ihp.oisc.regs[7][12] ));
 sg13g2_a22oi_1 _22577_ (.Y(_05975_),
    .B1(_05754_),
    .B2(\top_ihp.oisc.regs[12][12] ),
    .A2(_05505_),
    .A1(\top_ihp.oisc.regs[1][12] ));
 sg13g2_and4_1 _22578_ (.A(_05972_),
    .B(_05973_),
    .C(_05974_),
    .D(_05975_),
    .X(_05976_));
 sg13g2_a22oi_1 _22579_ (.Y(_05977_),
    .B1(net177),
    .B2(\top_ihp.oisc.regs[58][12] ),
    .A2(net417),
    .A1(\top_ihp.oisc.regs[57][12] ));
 sg13g2_buf_1 _22580_ (.A(_05718_),
    .X(_05978_));
 sg13g2_a22oi_1 _22581_ (.Y(_05979_),
    .B1(net392),
    .B2(\top_ihp.oisc.regs[52][12] ),
    .A2(net353),
    .A1(\top_ihp.oisc.regs[35][12] ));
 sg13g2_nand3_1 _22582_ (.B(_05977_),
    .C(_05979_),
    .A(_05976_),
    .Y(_05980_));
 sg13g2_buf_1 _22583_ (.A(_05669_),
    .X(_05981_));
 sg13g2_a22oi_1 _22584_ (.Y(_05982_),
    .B1(net366),
    .B2(\top_ihp.oisc.regs[49][12] ),
    .A2(net352),
    .A1(\top_ihp.oisc.regs[43][12] ));
 sg13g2_buf_8 _22585_ (.A(_05657_),
    .X(_05983_));
 sg13g2_a22oi_1 _22586_ (.Y(_05984_),
    .B1(net378),
    .B2(\top_ihp.oisc.regs[38][12] ),
    .A2(net174),
    .A1(\top_ihp.oisc.regs[62][12] ));
 sg13g2_a22oi_1 _22587_ (.Y(_05985_),
    .B1(net391),
    .B2(\top_ihp.oisc.regs[33][12] ),
    .A2(net419),
    .A1(\top_ihp.oisc.regs[44][12] ));
 sg13g2_buf_1 _22588_ (.A(_05635_),
    .X(_05986_));
 sg13g2_a22oi_1 _22589_ (.Y(_05987_),
    .B1(net393),
    .B2(\top_ihp.oisc.regs[42][12] ),
    .A2(net351),
    .A1(\top_ihp.oisc.regs[40][12] ));
 sg13g2_nand4_1 _22590_ (.B(_05984_),
    .C(_05985_),
    .A(_05982_),
    .Y(_05988_),
    .D(_05987_));
 sg13g2_a22oi_1 _22591_ (.Y(_05989_),
    .B1(net370),
    .B2(\top_ihp.oisc.regs[13][12] ),
    .A2(_05530_),
    .A1(\top_ihp.oisc.regs[29][12] ));
 sg13g2_a22oi_1 _22592_ (.Y(_05990_),
    .B1(net665),
    .B2(\top_ihp.oisc.regs[8][12] ),
    .A2(net546),
    .A1(\top_ihp.oisc.regs[14][12] ));
 sg13g2_nand2_1 _22593_ (.Y(_05991_),
    .A(\top_ihp.oisc.regs[24][12] ),
    .B(net402));
 sg13g2_a22oi_1 _22594_ (.Y(_05992_),
    .B1(net537),
    .B2(\top_ihp.oisc.regs[10][12] ),
    .A2(_05562_),
    .A1(\top_ihp.oisc.regs[9][12] ));
 sg13g2_and4_1 _22595_ (.A(_05989_),
    .B(_05990_),
    .C(_05991_),
    .D(_05992_),
    .X(_05993_));
 sg13g2_buf_8 _22596_ (.A(net380),
    .X(_05994_));
 sg13g2_a22oi_1 _22597_ (.Y(_05995_),
    .B1(net183),
    .B2(\top_ihp.oisc.regs[16][12] ),
    .A2(net173),
    .A1(\top_ihp.oisc.regs[11][12] ));
 sg13g2_a22oi_1 _22598_ (.Y(_05996_),
    .B1(net538),
    .B2(\top_ihp.oisc.regs[6][12] ),
    .A2(net204),
    .A1(\top_ihp.oisc.regs[4][12] ));
 sg13g2_nand3_1 _22599_ (.B(_05995_),
    .C(_05996_),
    .A(_05993_),
    .Y(_05997_));
 sg13g2_a22oi_1 _22600_ (.Y(_05998_),
    .B1(_05821_),
    .B2(\top_ihp.oisc.regs[21][12] ),
    .A2(net181),
    .A1(\top_ihp.oisc.regs[15][12] ));
 sg13g2_buf_8 _22601_ (.A(net427),
    .X(_05999_));
 sg13g2_a22oi_1 _22602_ (.Y(_06000_),
    .B1(net172),
    .B2(\top_ihp.oisc.regs[17][12] ),
    .A2(net434),
    .A1(\top_ihp.oisc.regs[20][12] ));
 sg13g2_buf_2 _22603_ (.A(net668),
    .X(_06001_));
 sg13g2_buf_2 _22604_ (.A(net543),
    .X(_06002_));
 sg13g2_a22oi_1 _22605_ (.Y(_06003_),
    .B1(net350),
    .B2(\top_ihp.oisc.regs[19][12] ),
    .A2(_06001_),
    .A1(\top_ihp.oisc.regs[28][12] ));
 sg13g2_and2_1 _22606_ (.A(\top_ihp.oisc.regs[5][12] ),
    .B(_05761_),
    .X(_06004_));
 sg13g2_a221oi_1 _22607_ (.B2(\top_ihp.oisc.regs[26][12] ),
    .C1(_06004_),
    .B1(_05911_),
    .A1(\top_ihp.oisc.regs[2][12] ),
    .Y(_06005_),
    .A2(_05900_));
 sg13g2_nand4_1 _22608_ (.B(_06000_),
    .C(_06003_),
    .A(_05998_),
    .Y(_06006_),
    .D(_06005_));
 sg13g2_nor4_1 _22609_ (.A(_05980_),
    .B(_05988_),
    .C(_05997_),
    .D(_06006_),
    .Y(_06007_));
 sg13g2_buf_8 _22610_ (.A(_05707_),
    .X(_06008_));
 sg13g2_buf_2 _22611_ (.A(_05744_),
    .X(_06009_));
 sg13g2_a21oi_1 _22612_ (.A1(_00216_),
    .A2(net59),
    .Y(_06010_),
    .B1(_06009_));
 sg13g2_nor2_1 _22613_ (.A(_05971_),
    .B(_06010_),
    .Y(_06011_));
 sg13g2_a21oi_1 _22614_ (.A1(_05969_),
    .A2(_06007_),
    .Y(_00391_),
    .B1(_06011_));
 sg13g2_nand2_1 _22615_ (.Y(_06012_),
    .A(\top_ihp.oisc.regs[62][13] ),
    .B(net176));
 sg13g2_a22oi_1 _22616_ (.Y(_06013_),
    .B1(net381),
    .B2(\top_ihp.oisc.regs[48][13] ),
    .A2(net186),
    .A1(\top_ihp.oisc.regs[59][13] ));
 sg13g2_a22oi_1 _22617_ (.Y(_06014_),
    .B1(net382),
    .B2(\top_ihp.oisc.regs[27][13] ),
    .A2(net413),
    .A1(\top_ihp.oisc.regs[63][13] ));
 sg13g2_a22oi_1 _22618_ (.Y(_06015_),
    .B1(_05929_),
    .B2(\top_ihp.oisc.regs[52][13] ),
    .A2(_05710_),
    .A1(\top_ihp.oisc.regs[41][13] ));
 sg13g2_nand4_1 _22619_ (.B(_06013_),
    .C(_06014_),
    .A(_06012_),
    .Y(_06016_),
    .D(_06015_));
 sg13g2_buf_8 _22620_ (.A(_05741_),
    .X(_06017_));
 sg13g2_buf_1 _22621_ (.A(_05725_),
    .X(_06018_));
 sg13g2_a22oi_1 _22622_ (.Y(_06019_),
    .B1(net349),
    .B2(\top_ihp.oisc.regs[46][13] ),
    .A2(_05615_),
    .A1(\top_ihp.oisc.regs[32][13] ));
 sg13g2_buf_1 _22623_ (.A(_05640_),
    .X(_06020_));
 sg13g2_a22oi_1 _22624_ (.Y(_06021_),
    .B1(net348),
    .B2(\top_ihp.oisc.regs[57][13] ),
    .A2(net435),
    .A1(\top_ihp.oisc.regs[31][13] ));
 sg13g2_nand3_1 _22625_ (.B(_06019_),
    .C(_06021_),
    .A(net57),
    .Y(_06022_));
 sg13g2_buf_1 _22626_ (.A(net835),
    .X(_06023_));
 sg13g2_nand2_1 _22627_ (.Y(_06024_),
    .A(_08046_),
    .B(net801));
 sg13g2_a22oi_1 _22628_ (.Y(_06025_),
    .B1(net719),
    .B2(\top_ihp.oisc.regs[23][13] ),
    .A2(_05820_),
    .A1(\top_ihp.oisc.regs[21][13] ));
 sg13g2_nand2_1 _22629_ (.Y(_06026_),
    .A(_06024_),
    .B(_06025_));
 sg13g2_a221oi_1 _22630_ (.B2(\top_ihp.oisc.regs[15][13] ),
    .C1(_06026_),
    .B1(net428),
    .A1(\top_ihp.oisc.regs[9][13] ),
    .Y(_06027_),
    .A2(net374));
 sg13g2_a22oi_1 _22631_ (.Y(_06028_),
    .B1(_05937_),
    .B2(\top_ihp.oisc.regs[33][13] ),
    .A2(net200),
    .A1(\top_ihp.oisc.regs[61][13] ));
 sg13g2_buf_2 _22632_ (.A(_05847_),
    .X(_06029_));
 sg13g2_a22oi_1 _22633_ (.Y(_06030_),
    .B1(net171),
    .B2(\top_ihp.oisc.regs[60][13] ),
    .A2(net352),
    .A1(\top_ihp.oisc.regs[43][13] ));
 sg13g2_a22oi_1 _22634_ (.Y(_06031_),
    .B1(_05839_),
    .B2(\top_ihp.oisc.regs[47][13] ),
    .A2(_05863_),
    .A1(\top_ihp.oisc.regs[50][13] ));
 sg13g2_nand4_1 _22635_ (.B(_06028_),
    .C(_06030_),
    .A(_06027_),
    .Y(_06032_),
    .D(_06031_));
 sg13g2_a22oi_1 _22636_ (.Y(_06033_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[34][13] ),
    .A2(net196),
    .A1(\top_ihp.oisc.regs[54][13] ));
 sg13g2_a22oi_1 _22637_ (.Y(_06034_),
    .B1(net202),
    .B2(\top_ihp.oisc.regs[44][13] ),
    .A2(net424),
    .A1(\top_ihp.oisc.regs[39][13] ));
 sg13g2_a22oi_1 _22638_ (.Y(_06035_),
    .B1(net386),
    .B2(\top_ihp.oisc.regs[49][13] ),
    .A2(net408),
    .A1(\top_ihp.oisc.regs[35][13] ));
 sg13g2_a22oi_1 _22639_ (.Y(_06036_),
    .B1(net177),
    .B2(\top_ihp.oisc.regs[58][13] ),
    .A2(net378),
    .A1(\top_ihp.oisc.regs[38][13] ));
 sg13g2_nand4_1 _22640_ (.B(_06034_),
    .C(_06035_),
    .A(_06033_),
    .Y(_06037_),
    .D(_06036_));
 sg13g2_nor4_2 _22641_ (.A(_06016_),
    .B(_06022_),
    .C(_06032_),
    .Y(_06038_),
    .D(_06037_));
 sg13g2_a22oi_1 _22642_ (.Y(_06039_),
    .B1(net420),
    .B2(\top_ihp.oisc.regs[51][13] ),
    .A2(_05654_),
    .A1(\top_ihp.oisc.regs[56][13] ));
 sg13g2_buf_1 _22643_ (.A(_05595_),
    .X(_06040_));
 sg13g2_a22oi_1 _22644_ (.Y(_06041_),
    .B1(net347),
    .B2(\top_ihp.oisc.regs[37][13] ),
    .A2(net351),
    .A1(\top_ihp.oisc.regs[40][13] ));
 sg13g2_buf_8 _22645_ (.A(_05659_),
    .X(_06042_));
 sg13g2_a22oi_1 _22646_ (.Y(_06043_),
    .B1(net346),
    .B2(\top_ihp.oisc.regs[30][13] ),
    .A2(net416),
    .A1(\top_ihp.oisc.regs[42][13] ));
 sg13g2_a22oi_1 _22647_ (.Y(_06044_),
    .B1(net411),
    .B2(\top_ihp.oisc.regs[45][13] ),
    .A2(_05455_),
    .A1(\top_ihp.oisc.regs[36][13] ));
 sg13g2_nand4_1 _22648_ (.B(_06041_),
    .C(_06043_),
    .A(_06039_),
    .Y(_06045_),
    .D(_06044_));
 sg13g2_buf_8 _22649_ (.A(_05761_),
    .X(_06046_));
 sg13g2_a22oi_1 _22650_ (.Y(_06047_),
    .B1(net345),
    .B2(\top_ihp.oisc.regs[5][13] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[29][13] ));
 sg13g2_a22oi_1 _22651_ (.Y(_06048_),
    .B1(net537),
    .B2(\top_ihp.oisc.regs[10][13] ),
    .A2(net546),
    .A1(\top_ihp.oisc.regs[14][13] ));
 sg13g2_a22oi_1 _22652_ (.Y(_06049_),
    .B1(net402),
    .B2(\top_ihp.oisc.regs[24][13] ),
    .A2(net372),
    .A1(\top_ihp.oisc.regs[12][13] ));
 sg13g2_a22oi_1 _22653_ (.Y(_06050_),
    .B1(net371),
    .B2(\top_ihp.oisc.regs[16][13] ),
    .A2(net553),
    .A1(\top_ihp.oisc.regs[22][13] ));
 sg13g2_nand4_1 _22654_ (.B(_06048_),
    .C(_06049_),
    .A(_06047_),
    .Y(_06051_),
    .D(_06050_));
 sg13g2_buf_1 _22655_ (.A(_05647_),
    .X(_06052_));
 sg13g2_a22oi_1 _22656_ (.Y(_06053_),
    .B1(net398),
    .B2(\top_ihp.oisc.regs[55][13] ),
    .A2(net344),
    .A1(\top_ihp.oisc.regs[53][13] ));
 sg13g2_nand2b_1 _22657_ (.Y(_06054_),
    .B(_06053_),
    .A_N(_06051_));
 sg13g2_a22oi_1 _22658_ (.Y(_06055_),
    .B1(net373),
    .B2(\top_ihp.oisc.regs[1][13] ),
    .A2(net434),
    .A1(\top_ihp.oisc.regs[20][13] ));
 sg13g2_a22oi_1 _22659_ (.Y(_06056_),
    .B1(net179),
    .B2(\top_ihp.oisc.regs[2][13] ),
    .A2(_05903_),
    .A1(\top_ihp.oisc.regs[25][13] ));
 sg13g2_buf_2 _22660_ (.A(_05542_),
    .X(_06057_));
 sg13g2_a22oi_1 _22661_ (.Y(_06058_),
    .B1(net180),
    .B2(\top_ihp.oisc.regs[13][13] ),
    .A2(net664),
    .A1(\top_ihp.oisc.regs[28][13] ));
 sg13g2_buf_8 _22662_ (.A(net401),
    .X(_06059_));
 sg13g2_a22oi_1 _22663_ (.Y(_06060_),
    .B1(net667),
    .B2(\top_ihp.oisc.regs[6][13] ),
    .A2(net170),
    .A1(\top_ihp.oisc.regs[3][13] ));
 sg13g2_nand4_1 _22664_ (.B(_06056_),
    .C(_06058_),
    .A(_06055_),
    .Y(_06061_),
    .D(_06060_));
 sg13g2_buf_8 _22665_ (.A(_05547_),
    .X(_06062_));
 sg13g2_buf_8 _22666_ (.A(net534),
    .X(_06063_));
 sg13g2_a22oi_1 _22667_ (.Y(_06064_),
    .B1(net350),
    .B2(\top_ihp.oisc.regs[19][13] ),
    .A2(net343),
    .A1(\top_ihp.oisc.regs[18][13] ));
 sg13g2_buf_2 _22668_ (.A(net554),
    .X(_06065_));
 sg13g2_buf_1 _22669_ (.A(_05857_),
    .X(_06066_));
 sg13g2_a22oi_1 _22670_ (.Y(_06067_),
    .B1(net169),
    .B2(\top_ihp.oisc.regs[11][13] ),
    .A2(net342),
    .A1(\top_ihp.oisc.regs[7][13] ));
 sg13g2_buf_8 _22671_ (.A(net367),
    .X(_06068_));
 sg13g2_a22oi_1 _22672_ (.Y(_06069_),
    .B1(net536),
    .B2(\top_ihp.oisc.regs[8][13] ),
    .A2(net168),
    .A1(\top_ihp.oisc.regs[26][13] ));
 sg13g2_a22oi_1 _22673_ (.Y(_06070_),
    .B1(net172),
    .B2(\top_ihp.oisc.regs[17][13] ),
    .A2(net204),
    .A1(\top_ihp.oisc.regs[4][13] ));
 sg13g2_nand4_1 _22674_ (.B(_06067_),
    .C(_06069_),
    .A(_06064_),
    .Y(_06071_),
    .D(_06070_));
 sg13g2_nor4_1 _22675_ (.A(_06045_),
    .B(_06054_),
    .C(_06061_),
    .D(_06071_),
    .Y(_06072_));
 sg13g2_a21o_1 _22676_ (.A2(net63),
    .A1(_00217_),
    .B1(net58),
    .X(_06073_));
 sg13g2_a22oi_1 _22677_ (.Y(_00392_),
    .B1(_06073_),
    .B2(_06024_),
    .A2(_06072_),
    .A1(_06038_));
 sg13g2_a22oi_1 _22678_ (.Y(_06074_),
    .B1(_05713_),
    .B2(\top_ihp.oisc.regs[48][14] ),
    .A2(_05605_),
    .A1(\top_ihp.oisc.regs[39][14] ));
 sg13g2_a22oi_1 _22679_ (.Y(_06075_),
    .B1(_05728_),
    .B2(\top_ihp.oisc.regs[52][14] ),
    .A2(_05680_),
    .A1(\top_ihp.oisc.regs[45][14] ));
 sg13g2_a22oi_1 _22680_ (.Y(_06076_),
    .B1(_05654_),
    .B2(\top_ihp.oisc.regs[56][14] ),
    .A2(_05640_),
    .A1(\top_ihp.oisc.regs[57][14] ));
 sg13g2_a22oi_1 _22681_ (.Y(_06077_),
    .B1(_05735_),
    .B2(\top_ihp.oisc.regs[55][14] ),
    .A2(_05614_),
    .A1(\top_ihp.oisc.regs[32][14] ));
 sg13g2_and4_1 _22682_ (.A(_06074_),
    .B(_06075_),
    .C(_06076_),
    .D(_06077_),
    .X(_06078_));
 sg13g2_a22oi_1 _22683_ (.Y(_06079_),
    .B1(net346),
    .B2(\top_ihp.oisc.regs[30][14] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[36][14] ));
 sg13g2_buf_1 _22684_ (.A(_05608_),
    .X(_06080_));
 sg13g2_a22oi_1 _22685_ (.Y(_06081_),
    .B1(_05545_),
    .B2(\top_ihp.oisc.regs[38][14] ),
    .A2(net722),
    .A1(\top_ihp.oisc.regs[44][14] ));
 sg13g2_nor3_1 _22686_ (.A(_05770_),
    .B(_05612_),
    .C(_06081_),
    .Y(_06082_));
 sg13g2_a21oi_1 _22687_ (.A1(\top_ihp.oisc.regs[27][14] ),
    .A2(net341),
    .Y(_06083_),
    .B1(_06082_));
 sg13g2_nand4_1 _22688_ (.B(_06078_),
    .C(_06079_),
    .A(net61),
    .Y(_06084_),
    .D(_06083_));
 sg13g2_a22oi_1 _22689_ (.Y(_06085_),
    .B1(net171),
    .B2(\top_ihp.oisc.regs[60][14] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[53][14] ));
 sg13g2_buf_2 _22690_ (.A(_05710_),
    .X(_06086_));
 sg13g2_a22oi_1 _22691_ (.Y(_06087_),
    .B1(net340),
    .B2(\top_ihp.oisc.regs[41][14] ),
    .A2(net188),
    .A1(\top_ihp.oisc.regs[50][14] ));
 sg13g2_nand3_1 _22692_ (.B(net728),
    .C(_05633_),
    .A(\top_ihp.oisc.regs[40][14] ),
    .Y(_06088_));
 sg13g2_nand2_1 _22693_ (.Y(_06089_),
    .A(\top_ihp.oisc.regs[19][14] ),
    .B(net543));
 sg13g2_nand2_1 _22694_ (.Y(_06090_),
    .A(_08014_),
    .B(net801));
 sg13g2_buf_2 _22695_ (.A(_05820_),
    .X(_06091_));
 sg13g2_a22oi_1 _22696_ (.Y(_06092_),
    .B1(_05970_),
    .B2(\top_ihp.oisc.regs[23][14] ),
    .A2(_06091_),
    .A1(\top_ihp.oisc.regs[21][14] ));
 sg13g2_and4_1 _22697_ (.A(_06088_),
    .B(_06089_),
    .C(_06090_),
    .D(_06092_),
    .X(_06093_));
 sg13g2_buf_1 _22698_ (.A(_05535_),
    .X(_06094_));
 sg13g2_nand3_1 _22699_ (.B(net671),
    .C(net662),
    .A(\top_ihp.oisc.regs[54][14] ),
    .Y(_06095_));
 sg13g2_nand3_1 _22700_ (.B(net548),
    .C(net727),
    .A(\top_ihp.oisc.regs[58][14] ),
    .Y(_06096_));
 sg13g2_nand2_1 _22701_ (.Y(_06097_),
    .A(_05485_),
    .B(net673));
 sg13g2_a21oi_1 _22702_ (.A1(_06095_),
    .A2(_06096_),
    .Y(_06098_),
    .B1(_06097_));
 sg13g2_a21oi_1 _22703_ (.A1(\top_ihp.oisc.regs[31][14] ),
    .A2(net389),
    .Y(_06099_),
    .B1(_06098_));
 sg13g2_nand4_1 _22704_ (.B(_06087_),
    .C(_06093_),
    .A(_06085_),
    .Y(_06100_),
    .D(_06099_));
 sg13g2_a22oi_1 _22705_ (.Y(_06101_),
    .B1(_05841_),
    .B2(\top_ihp.oisc.regs[49][14] ),
    .A2(net365),
    .A1(\top_ihp.oisc.regs[63][14] ));
 sg13g2_buf_8 _22706_ (.A(net402),
    .X(_06102_));
 sg13g2_nand2_1 _22707_ (.Y(_06103_),
    .A(\top_ihp.oisc.regs[24][14] ),
    .B(net167));
 sg13g2_a22oi_1 _22708_ (.Y(_06104_),
    .B1(net373),
    .B2(\top_ihp.oisc.regs[1][14] ),
    .A2(net342),
    .A1(\top_ihp.oisc.regs[7][14] ));
 sg13g2_nand3_1 _22709_ (.B(_06103_),
    .C(_06104_),
    .A(_06101_),
    .Y(_06105_));
 sg13g2_buf_8 _22710_ (.A(_05778_),
    .X(_06106_));
 sg13g2_a22oi_1 _22711_ (.Y(_06107_),
    .B1(net166),
    .B2(\top_ihp.oisc.regs[3][14] ),
    .A2(net204),
    .A1(\top_ihp.oisc.regs[4][14] ));
 sg13g2_a22oi_1 _22712_ (.Y(_06108_),
    .B1(net184),
    .B2(\top_ihp.oisc.regs[12][14] ),
    .A2(net173),
    .A1(\top_ihp.oisc.regs[11][14] ));
 sg13g2_a22oi_1 _22713_ (.Y(_06109_),
    .B1(net168),
    .B2(\top_ihp.oisc.regs[26][14] ),
    .A2(net538),
    .A1(\top_ihp.oisc.regs[6][14] ));
 sg13g2_nor2_1 _22714_ (.A(_05554_),
    .B(_05612_),
    .Y(_06110_));
 sg13g2_mux2_1 _22715_ (.A0(\top_ihp.oisc.regs[42][14] ),
    .A1(\top_ihp.oisc.regs[34][14] ),
    .S(net662),
    .X(_06111_));
 sg13g2_a22oi_1 _22716_ (.Y(_06112_),
    .B1(_06110_),
    .B2(_06111_),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[22][14] ));
 sg13g2_nand4_1 _22717_ (.B(_06108_),
    .C(_06109_),
    .A(_06107_),
    .Y(_06113_),
    .D(_06112_));
 sg13g2_nor4_1 _22718_ (.A(_06084_),
    .B(_06100_),
    .C(_06105_),
    .D(_06113_),
    .Y(_06114_));
 sg13g2_buf_8 _22719_ (.A(net345),
    .X(_06115_));
 sg13g2_a22oi_1 _22720_ (.Y(_06116_),
    .B1(net165),
    .B2(\top_ihp.oisc.regs[5][14] ),
    .A2(net371),
    .A1(\top_ihp.oisc.regs[16][14] ));
 sg13g2_a22oi_1 _22721_ (.Y(_06117_),
    .B1(net181),
    .B2(\top_ihp.oisc.regs[15][14] ),
    .A2(_05899_),
    .A1(\top_ihp.oisc.regs[13][14] ));
 sg13g2_mux2_1 _22722_ (.A0(\top_ihp.oisc.regs[10][14] ),
    .A1(\top_ihp.oisc.regs[8][14] ),
    .S(net545),
    .X(_06118_));
 sg13g2_nor2_2 _22723_ (.A(net671),
    .B(_05512_),
    .Y(_06119_));
 sg13g2_a22oi_1 _22724_ (.Y(_06120_),
    .B1(_06118_),
    .B2(_06119_),
    .A2(net535),
    .A1(\top_ihp.oisc.regs[28][14] ));
 sg13g2_a22oi_1 _22725_ (.Y(_06121_),
    .B1(_05999_),
    .B2(\top_ihp.oisc.regs[17][14] ),
    .A2(net434),
    .A1(\top_ihp.oisc.regs[20][14] ));
 sg13g2_nand4_1 _22726_ (.B(_06117_),
    .C(_06120_),
    .A(_06116_),
    .Y(_06122_),
    .D(_06121_));
 sg13g2_and2_1 _22727_ (.A(\top_ihp.oisc.regs[46][14] ),
    .B(net728),
    .X(_06123_));
 sg13g2_a22oi_1 _22728_ (.Y(_06124_),
    .B1(_06123_),
    .B2(_05458_),
    .A2(net185),
    .A1(\top_ihp.oisc.regs[9][14] ));
 sg13g2_a22oi_1 _22729_ (.Y(_06125_),
    .B1(net182),
    .B2(\top_ihp.oisc.regs[29][14] ),
    .A2(_05483_),
    .A1(\top_ihp.oisc.regs[25][14] ));
 sg13g2_and2_1 _22730_ (.A(\top_ihp.oisc.regs[43][14] ),
    .B(_05593_),
    .X(_06126_));
 sg13g2_a22oi_1 _22731_ (.Y(_06127_),
    .B1(_06126_),
    .B2(_05403_),
    .A2(net430),
    .A1(\top_ihp.oisc.regs[14][14] ));
 sg13g2_a22oi_1 _22732_ (.Y(_06128_),
    .B1(net179),
    .B2(\top_ihp.oisc.regs[2][14] ),
    .A2(_06062_),
    .A1(\top_ihp.oisc.regs[18][14] ));
 sg13g2_nand4_1 _22733_ (.B(_06125_),
    .C(_06127_),
    .A(_06124_),
    .Y(_06129_),
    .D(_06128_));
 sg13g2_a22oi_1 _22734_ (.Y(_06130_),
    .B1(net407),
    .B2(\top_ihp.oisc.regs[33][14] ),
    .A2(net190),
    .A1(\top_ihp.oisc.regs[61][14] ));
 sg13g2_a22oi_1 _22735_ (.Y(_06131_),
    .B1(net361),
    .B2(\top_ihp.oisc.regs[35][14] ),
    .A2(net191),
    .A1(\top_ihp.oisc.regs[59][14] ));
 sg13g2_a22oi_1 _22736_ (.Y(_06132_),
    .B1(net355),
    .B2(\top_ihp.oisc.regs[51][14] ),
    .A2(net176),
    .A1(\top_ihp.oisc.regs[62][14] ));
 sg13g2_a22oi_1 _22737_ (.Y(_06133_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[47][14] ),
    .A2(net426),
    .A1(\top_ihp.oisc.regs[37][14] ));
 sg13g2_nand4_1 _22738_ (.B(_06131_),
    .C(_06132_),
    .A(_06130_),
    .Y(_06134_),
    .D(_06133_));
 sg13g2_nor3_1 _22739_ (.A(_06122_),
    .B(_06129_),
    .C(_06134_),
    .Y(_06135_));
 sg13g2_inv_1 _22740_ (.Y(_06136_),
    .A(_00218_));
 sg13g2_o21ai_1 _22741_ (.B1(net27),
    .Y(_06137_),
    .A1(_06136_),
    .A2(net62));
 sg13g2_a22oi_1 _22742_ (.Y(_00393_),
    .B1(_06137_),
    .B2(_06090_),
    .A2(_06135_),
    .A1(_06114_));
 sg13g2_a22oi_1 _22743_ (.Y(_06138_),
    .B1(net349),
    .B2(\top_ihp.oisc.regs[46][15] ),
    .A2(net435),
    .A1(\top_ihp.oisc.regs[31][15] ));
 sg13g2_buf_1 _22744_ (.A(_05687_),
    .X(_06139_));
 sg13g2_a22oi_1 _22745_ (.Y(_06140_),
    .B1(net339),
    .B2(\top_ihp.oisc.regs[38][15] ),
    .A2(net188),
    .A1(\top_ihp.oisc.regs[50][15] ));
 sg13g2_buf_2 _22746_ (.A(_05614_),
    .X(_06141_));
 sg13g2_a22oi_1 _22747_ (.Y(_06142_),
    .B1(net381),
    .B2(\top_ihp.oisc.regs[48][15] ),
    .A2(net338),
    .A1(\top_ihp.oisc.regs[32][15] ));
 sg13g2_buf_2 _22748_ (.A(_05605_),
    .X(_06143_));
 sg13g2_a22oi_1 _22749_ (.Y(_06144_),
    .B1(net420),
    .B2(\top_ihp.oisc.regs[51][15] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[39][15] ));
 sg13g2_nand4_1 _22750_ (.B(_06140_),
    .C(_06142_),
    .A(_06138_),
    .Y(_06145_),
    .D(_06144_));
 sg13g2_buf_8 _22751_ (.A(_05438_),
    .X(_06146_));
 sg13g2_and2_1 _22752_ (.A(\top_ihp.oisc.regs[26][15] ),
    .B(_05765_),
    .X(_06147_));
 sg13g2_a221oi_1 _22753_ (.B2(\top_ihp.oisc.regs[13][15] ),
    .C1(_06147_),
    .B1(net390),
    .A1(\top_ihp.oisc.regs[22][15] ),
    .Y(_06148_),
    .A2(_06146_));
 sg13g2_buf_8 _22754_ (.A(net374),
    .X(_06149_));
 sg13g2_a22oi_1 _22755_ (.Y(_06150_),
    .B1(net173),
    .B2(\top_ihp.oisc.regs[11][15] ),
    .A2(net164),
    .A1(\top_ihp.oisc.regs[9][15] ));
 sg13g2_a22oi_1 _22756_ (.Y(_06151_),
    .B1(net167),
    .B2(\top_ihp.oisc.regs[24][15] ),
    .A2(net667),
    .A1(\top_ihp.oisc.regs[6][15] ));
 sg13g2_a22oi_1 _22757_ (.Y(_06152_),
    .B1(net383),
    .B2(\top_ihp.oisc.regs[60][15] ),
    .A2(net201),
    .A1(\top_ihp.oisc.regs[54][15] ));
 sg13g2_nand4_1 _22758_ (.B(_06150_),
    .C(_06151_),
    .A(_06148_),
    .Y(_06153_),
    .D(_06152_));
 sg13g2_a22oi_1 _22759_ (.Y(_06154_),
    .B1(net183),
    .B2(\top_ihp.oisc.regs[16][15] ),
    .A2(net373),
    .A1(\top_ihp.oisc.regs[1][15] ));
 sg13g2_a22oi_1 _22760_ (.Y(_06155_),
    .B1(net350),
    .B2(\top_ihp.oisc.regs[19][15] ),
    .A2(net430),
    .A1(\top_ihp.oisc.regs[14][15] ));
 sg13g2_buf_8 _22761_ (.A(_05500_),
    .X(_06156_));
 sg13g2_a22oi_1 _22762_ (.Y(_06157_),
    .B1(net179),
    .B2(\top_ihp.oisc.regs[2][15] ),
    .A2(net163),
    .A1(\top_ihp.oisc.regs[4][15] ));
 sg13g2_a22oi_1 _22763_ (.Y(_06158_),
    .B1(net343),
    .B2(\top_ihp.oisc.regs[18][15] ),
    .A2(net535),
    .A1(\top_ihp.oisc.regs[28][15] ));
 sg13g2_nand4_1 _22764_ (.B(_06155_),
    .C(_06157_),
    .A(_06154_),
    .Y(_06159_),
    .D(_06158_));
 sg13g2_a22oi_1 _22765_ (.Y(_06160_),
    .B1(net166),
    .B2(\top_ihp.oisc.regs[3][15] ),
    .A2(net434),
    .A1(\top_ihp.oisc.regs[20][15] ));
 sg13g2_a22oi_1 _22766_ (.Y(_06161_),
    .B1(net165),
    .B2(\top_ihp.oisc.regs[5][15] ),
    .A2(net184),
    .A1(\top_ihp.oisc.regs[12][15] ));
 sg13g2_a22oi_1 _22767_ (.Y(_06162_),
    .B1(net182),
    .B2(\top_ihp.oisc.regs[29][15] ),
    .A2(_05483_),
    .A1(\top_ihp.oisc.regs[25][15] ));
 sg13g2_buf_2 _22768_ (.A(net428),
    .X(_06163_));
 sg13g2_a22oi_1 _22769_ (.Y(_06164_),
    .B1(net172),
    .B2(\top_ihp.oisc.regs[17][15] ),
    .A2(net162),
    .A1(\top_ihp.oisc.regs[15][15] ));
 sg13g2_nand4_1 _22770_ (.B(_06161_),
    .C(_06162_),
    .A(_06160_),
    .Y(_06165_),
    .D(_06164_));
 sg13g2_nor4_1 _22771_ (.A(_06145_),
    .B(_06153_),
    .C(_06159_),
    .D(_06165_),
    .Y(_06166_));
 sg13g2_a22oi_1 _22772_ (.Y(_06167_),
    .B1(net408),
    .B2(\top_ihp.oisc.regs[35][15] ),
    .A2(net417),
    .A1(\top_ihp.oisc.regs[57][15] ));
 sg13g2_a22oi_1 _22773_ (.Y(_06168_),
    .B1(net379),
    .B2(\top_ihp.oisc.regs[45][15] ),
    .A2(_05659_),
    .A1(\top_ihp.oisc.regs[30][15] ));
 sg13g2_a22oi_1 _22774_ (.Y(_06169_),
    .B1(net359),
    .B2(\top_ihp.oisc.regs[55][15] ),
    .A2(net542),
    .A1(\top_ihp.oisc.regs[34][15] ));
 sg13g2_a22oi_1 _22775_ (.Y(_06170_),
    .B1(net186),
    .B2(\top_ihp.oisc.regs[59][15] ),
    .A2(_05647_),
    .A1(\top_ihp.oisc.regs[53][15] ));
 sg13g2_nand4_1 _22776_ (.B(_06168_),
    .C(_06169_),
    .A(_06167_),
    .Y(_06171_),
    .D(_06170_));
 sg13g2_buf_1 _22777_ (.A(_05644_),
    .X(_06172_));
 sg13g2_nand2_1 _22778_ (.Y(_06173_),
    .A(\top_ihp.oisc.regs[42][15] ),
    .B(net336));
 sg13g2_nand3_1 _22779_ (.B(net750),
    .C(net549),
    .A(\top_ihp.oisc.regs[23][15] ),
    .Y(_06174_));
 sg13g2_buf_1 _22780_ (.A(_05526_),
    .X(_06175_));
 sg13g2_nand3_1 _22781_ (.B(net548),
    .C(net747),
    .A(\top_ihp.oisc.regs[10][15] ),
    .Y(_06176_));
 sg13g2_nand3_1 _22782_ (.B(_06174_),
    .C(_06176_),
    .A(net550),
    .Y(_06177_));
 sg13g2_nand3_1 _22783_ (.B(net750),
    .C(net549),
    .A(\top_ihp.oisc.regs[21][15] ),
    .Y(_06178_));
 sg13g2_nand3_1 _22784_ (.B(net548),
    .C(net747),
    .A(\top_ihp.oisc.regs[8][15] ),
    .Y(_06179_));
 sg13g2_nand3_1 _22785_ (.B(_06178_),
    .C(_06179_),
    .A(net545),
    .Y(_06180_));
 sg13g2_a22oi_1 _22786_ (.Y(_06181_),
    .B1(_06177_),
    .B2(_06180_),
    .A2(net404),
    .A1(\top_ihp.oisc.regs[49][15] ));
 sg13g2_nand3_1 _22787_ (.B(_06173_),
    .C(_06181_),
    .A(net61),
    .Y(_06182_));
 sg13g2_nor2_2 _22788_ (.A(_04123_),
    .B(net804),
    .Y(_06183_));
 sg13g2_a221oi_1 _22789_ (.B2(\top_ihp.oisc.regs[41][15] ),
    .C1(_06183_),
    .B1(net340),
    .A1(\top_ihp.oisc.regs[7][15] ),
    .Y(_06184_),
    .A2(_05430_));
 sg13g2_a22oi_1 _22790_ (.Y(_06185_),
    .B1(net387),
    .B2(\top_ihp.oisc.regs[47][15] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[40][15] ));
 sg13g2_a22oi_1 _22791_ (.Y(_06186_),
    .B1(net365),
    .B2(\top_ihp.oisc.regs[63][15] ),
    .A2(net375),
    .A1(\top_ihp.oisc.regs[36][15] ));
 sg13g2_a22oi_1 _22792_ (.Y(_06187_),
    .B1(net382),
    .B2(\top_ihp.oisc.regs[27][15] ),
    .A2(net200),
    .A1(\top_ihp.oisc.regs[61][15] ));
 sg13g2_nand4_1 _22793_ (.B(_06185_),
    .C(_06186_),
    .A(_06184_),
    .Y(_06188_),
    .D(_06187_));
 sg13g2_buf_8 _22794_ (.A(net419),
    .X(_06189_));
 sg13g2_a22oi_1 _22795_ (.Y(_06190_),
    .B1(net193),
    .B2(\top_ihp.oisc.regs[56][15] ),
    .A2(net161),
    .A1(\top_ihp.oisc.regs[44][15] ));
 sg13g2_a22oi_1 _22796_ (.Y(_06191_),
    .B1(net195),
    .B2(\top_ihp.oisc.regs[58][15] ),
    .A2(net397),
    .A1(\top_ihp.oisc.regs[37][15] ));
 sg13g2_a22oi_1 _22797_ (.Y(_06192_),
    .B1(net405),
    .B2(\top_ihp.oisc.regs[52][15] ),
    .A2(net391),
    .A1(\top_ihp.oisc.regs[33][15] ));
 sg13g2_a22oi_1 _22798_ (.Y(_06193_),
    .B1(net412),
    .B2(\top_ihp.oisc.regs[43][15] ),
    .A2(net192),
    .A1(\top_ihp.oisc.regs[62][15] ));
 sg13g2_nand4_1 _22799_ (.B(_06191_),
    .C(_06192_),
    .A(_06190_),
    .Y(_06194_),
    .D(_06193_));
 sg13g2_nor4_2 _22800_ (.A(_06171_),
    .B(_06182_),
    .C(_06188_),
    .Y(_06195_),
    .D(_06194_));
 sg13g2_a21oi_1 _22801_ (.A1(_00219_),
    .A2(net59),
    .Y(_06196_),
    .B1(net58));
 sg13g2_nor2_1 _22802_ (.A(_06183_),
    .B(_06196_),
    .Y(_06197_));
 sg13g2_a21oi_1 _22803_ (.A1(_06166_),
    .A2(_06195_),
    .Y(_00394_),
    .B1(_06197_));
 sg13g2_a22oi_1 _22804_ (.Y(_06198_),
    .B1(net348),
    .B2(\top_ihp.oisc.regs[57][16] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[40][16] ));
 sg13g2_a22oi_1 _22805_ (.Y(_06199_),
    .B1(net161),
    .B2(\top_ihp.oisc.regs[44][16] ),
    .A2(net347),
    .A1(\top_ihp.oisc.regs[37][16] ));
 sg13g2_a22oi_1 _22806_ (.Y(_06200_),
    .B1(net338),
    .B2(\top_ihp.oisc.regs[32][16] ),
    .A2(net186),
    .A1(\top_ihp.oisc.regs[59][16] ));
 sg13g2_a22oi_1 _22807_ (.Y(_06201_),
    .B1(net383),
    .B2(\top_ihp.oisc.regs[60][16] ),
    .A2(net406),
    .A1(\top_ihp.oisc.regs[46][16] ));
 sg13g2_nand4_1 _22808_ (.B(_06199_),
    .C(_06200_),
    .A(_06198_),
    .Y(_06202_),
    .D(_06201_));
 sg13g2_a22oi_1 _22809_ (.Y(_06203_),
    .B1(net407),
    .B2(\top_ihp.oisc.regs[33][16] ),
    .A2(_05951_),
    .A1(\top_ihp.oisc.regs[47][16] ));
 sg13g2_a22oi_1 _22810_ (.Y(_06204_),
    .B1(net177),
    .B2(\top_ihp.oisc.regs[58][16] ),
    .A2(net362),
    .A1(\top_ihp.oisc.regs[43][16] ));
 sg13g2_nand3_1 _22811_ (.B(_06203_),
    .C(_06204_),
    .A(net61),
    .Y(_06205_));
 sg13g2_a22oi_1 _22812_ (.Y(_06206_),
    .B1(net405),
    .B2(\top_ihp.oisc.regs[52][16] ),
    .A2(net340),
    .A1(\top_ihp.oisc.regs[41][16] ));
 sg13g2_a22oi_1 _22813_ (.Y(_06207_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[34][16] ),
    .A2(net346),
    .A1(\top_ihp.oisc.regs[30][16] ));
 sg13g2_a22oi_1 _22814_ (.Y(_06208_),
    .B1(net187),
    .B2(\top_ihp.oisc.regs[56][16] ),
    .A2(net435),
    .A1(\top_ihp.oisc.regs[31][16] ));
 sg13g2_a22oi_1 _22815_ (.Y(_06209_),
    .B1(net175),
    .B2(\top_ihp.oisc.regs[61][16] ),
    .A2(net174),
    .A1(\top_ihp.oisc.regs[62][16] ));
 sg13g2_nand4_1 _22816_ (.B(_06207_),
    .C(_06208_),
    .A(_06206_),
    .Y(_06210_),
    .D(_06209_));
 sg13g2_a22oi_1 _22817_ (.Y(_06211_),
    .B1(net398),
    .B2(\top_ihp.oisc.regs[55][16] ),
    .A2(net366),
    .A1(\top_ihp.oisc.regs[49][16] ));
 sg13g2_a22oi_1 _22818_ (.Y(_06212_),
    .B1(net355),
    .B2(\top_ihp.oisc.regs[51][16] ),
    .A2(net196),
    .A1(\top_ihp.oisc.regs[54][16] ));
 sg13g2_a22oi_1 _22819_ (.Y(_06213_),
    .B1(net354),
    .B2(\top_ihp.oisc.regs[39][16] ),
    .A2(net336),
    .A1(\top_ihp.oisc.regs[42][16] ));
 sg13g2_a22oi_1 _22820_ (.Y(_06214_),
    .B1(net365),
    .B2(\top_ihp.oisc.regs[63][16] ),
    .A2(net344),
    .A1(\top_ihp.oisc.regs[53][16] ));
 sg13g2_nand4_1 _22821_ (.B(_06212_),
    .C(_06213_),
    .A(_06211_),
    .Y(_06215_),
    .D(_06214_));
 sg13g2_nor4_2 _22822_ (.A(_06202_),
    .B(_06205_),
    .C(_06210_),
    .Y(_06216_),
    .D(_06215_));
 sg13g2_a22oi_1 _22823_ (.Y(_06217_),
    .B1(net749),
    .B2(\top_ihp.oisc.regs[6][16] ),
    .A2(net724),
    .A1(\top_ihp.oisc.regs[7][16] ));
 sg13g2_nand2_1 _22824_ (.Y(_06218_),
    .A(_08010_),
    .B(_04085_));
 sg13g2_o21ai_1 _22825_ (.B1(_06218_),
    .Y(_06219_),
    .A1(_05418_),
    .A2(_06217_));
 sg13g2_a221oi_1 _22826_ (.B2(\top_ihp.oisc.regs[48][16] ),
    .C1(_06219_),
    .B1(net409),
    .A1(\top_ihp.oisc.regs[20][16] ),
    .Y(_06220_),
    .A2(net540));
 sg13g2_a22oi_1 _22827_ (.Y(_06221_),
    .B1(_05775_),
    .B2(\top_ihp.oisc.regs[24][16] ),
    .A2(_05505_),
    .A1(\top_ihp.oisc.regs[1][16] ));
 sg13g2_a22oi_1 _22828_ (.Y(_06222_),
    .B1(_05888_),
    .B2(\top_ihp.oisc.regs[12][16] ),
    .A2(_05543_),
    .A1(\top_ihp.oisc.regs[28][16] ));
 sg13g2_and2_1 _22829_ (.A(_06221_),
    .B(_06222_),
    .X(_06223_));
 sg13g2_a22oi_1 _22830_ (.Y(_06224_),
    .B1(net353),
    .B2(\top_ihp.oisc.regs[35][16] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[36][16] ));
 sg13g2_a22oi_1 _22831_ (.Y(_06225_),
    .B1(net341),
    .B2(\top_ihp.oisc.regs[27][16] ),
    .A2(_05676_),
    .A1(\top_ihp.oisc.regs[50][16] ));
 sg13g2_nand4_1 _22832_ (.B(_06223_),
    .C(_06224_),
    .A(_06220_),
    .Y(_06226_),
    .D(_06225_));
 sg13g2_a22oi_1 _22833_ (.Y(_06227_),
    .B1(net168),
    .B2(\top_ihp.oisc.regs[26][16] ),
    .A2(net430),
    .A1(\top_ihp.oisc.regs[14][16] ));
 sg13g2_nand3_1 _22834_ (.B(_05487_),
    .C(_05486_),
    .A(\top_ihp.oisc.regs[23][16] ),
    .Y(_06228_));
 sg13g2_nand3_1 _22835_ (.B(net669),
    .C(net724),
    .A(\top_ihp.oisc.regs[5][16] ),
    .Y(_06229_));
 sg13g2_nand3_1 _22836_ (.B(_05371_),
    .C(net722),
    .A(\top_ihp.oisc.regs[29][16] ),
    .Y(_06230_));
 sg13g2_nand3_1 _22837_ (.B(_06229_),
    .C(_06230_),
    .A(_06228_),
    .Y(_06231_));
 sg13g2_nand2_1 _22838_ (.Y(_06232_),
    .A(net549),
    .B(_06231_));
 sg13g2_a22oi_1 _22839_ (.Y(_06233_),
    .B1(net162),
    .B2(\top_ihp.oisc.regs[15][16] ),
    .A2(net170),
    .A1(\top_ihp.oisc.regs[3][16] ));
 sg13g2_a22oi_1 _22840_ (.Y(_06234_),
    .B1(net369),
    .B2(\top_ihp.oisc.regs[2][16] ),
    .A2(net390),
    .A1(\top_ihp.oisc.regs[13][16] ));
 sg13g2_nand4_1 _22841_ (.B(_06232_),
    .C(_06233_),
    .A(_06227_),
    .Y(_06235_),
    .D(_06234_));
 sg13g2_a22oi_1 _22842_ (.Y(_06236_),
    .B1(_05844_),
    .B2(\top_ihp.oisc.regs[38][16] ),
    .A2(net379),
    .A1(\top_ihp.oisc.regs[45][16] ));
 sg13g2_a22oi_1 _22843_ (.Y(_06237_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[25][16] ),
    .A2(_05390_),
    .A1(\top_ihp.oisc.regs[21][16] ));
 sg13g2_buf_8 _22844_ (.A(net427),
    .X(_06238_));
 sg13g2_a22oi_1 _22845_ (.Y(_06239_),
    .B1(_06238_),
    .B2(\top_ihp.oisc.regs[17][16] ),
    .A2(_06062_),
    .A1(\top_ihp.oisc.regs[18][16] ));
 sg13g2_mux2_1 _22846_ (.A0(\top_ihp.oisc.regs[10][16] ),
    .A1(\top_ihp.oisc.regs[8][16] ),
    .S(_05518_),
    .X(_06240_));
 sg13g2_a22oi_1 _22847_ (.Y(_06241_),
    .B1(_06119_),
    .B2(_06240_),
    .A2(_05759_),
    .A1(\top_ihp.oisc.regs[16][16] ));
 sg13g2_a22oi_1 _22848_ (.Y(_06242_),
    .B1(net374),
    .B2(\top_ihp.oisc.regs[9][16] ),
    .A2(_05499_),
    .A1(\top_ihp.oisc.regs[4][16] ));
 sg13g2_and2_1 _22849_ (.A(_06241_),
    .B(_06242_),
    .X(_06243_));
 sg13g2_nand4_1 _22850_ (.B(_06237_),
    .C(_06239_),
    .A(_06236_),
    .Y(_06244_),
    .D(_06243_));
 sg13g2_nand2_1 _22851_ (.Y(_06245_),
    .A(\top_ihp.oisc.regs[11][16] ),
    .B(net169));
 sg13g2_nor2_2 _22852_ (.A(_05818_),
    .B(_05554_),
    .Y(_06246_));
 sg13g2_a22oi_1 _22853_ (.Y(_06247_),
    .B1(_06246_),
    .B2(\top_ihp.oisc.regs[19][16] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[22][16] ));
 sg13g2_nand2_1 _22854_ (.Y(_06248_),
    .A(_06245_),
    .B(_06247_));
 sg13g2_nor4_1 _22855_ (.A(_06226_),
    .B(_06235_),
    .C(_06244_),
    .D(_06248_),
    .Y(_06249_));
 sg13g2_inv_1 _22856_ (.Y(_06250_),
    .A(_00220_));
 sg13g2_o21ai_1 _22857_ (.B1(_05746_),
    .Y(_06251_),
    .A1(_06250_),
    .A2(net62));
 sg13g2_a22oi_1 _22858_ (.Y(_00395_),
    .B1(_06251_),
    .B2(_06218_),
    .A2(_06249_),
    .A1(_06216_));
 sg13g2_a22oi_1 _22859_ (.Y(_06252_),
    .B1(_05750_),
    .B2(\top_ihp.oisc.regs[2][17] ),
    .A2(_05529_),
    .A1(\top_ihp.oisc.regs[29][17] ));
 sg13g2_a22oi_1 _22860_ (.Y(_06253_),
    .B1(_05761_),
    .B2(\top_ihp.oisc.regs[5][17] ),
    .A2(net370),
    .A1(\top_ihp.oisc.regs[13][17] ));
 sg13g2_a22oi_1 _22861_ (.Y(_06254_),
    .B1(net552),
    .B2(\top_ihp.oisc.regs[20][17] ),
    .A2(net553),
    .A1(\top_ihp.oisc.regs[22][17] ));
 sg13g2_nand2_1 _22862_ (.Y(_06255_),
    .A(\top_ihp.oisc.regs[12][17] ),
    .B(_05526_));
 sg13g2_nand4_1 _22863_ (.B(\top_ihp.oisc.regs[23][17] ),
    .C(_05373_),
    .A(net940),
    .Y(_06256_),
    .D(_05416_));
 sg13g2_o21ai_1 _22864_ (.B1(_06256_),
    .Y(_06257_),
    .A1(net672),
    .A2(_06255_));
 sg13g2_a22oi_1 _22865_ (.Y(_06258_),
    .B1(_06257_),
    .B2(_05489_),
    .A2(net544),
    .A1(\top_ihp.oisc.regs[18][17] ));
 sg13g2_and4_1 _22866_ (.A(_06252_),
    .B(_06253_),
    .C(_06254_),
    .D(_06258_),
    .X(_06259_));
 sg13g2_a22oi_1 _22867_ (.Y(_06260_),
    .B1(net749),
    .B2(\top_ihp.oisc.regs[6][17] ),
    .A2(net724),
    .A1(\top_ihp.oisc.regs[7][17] ));
 sg13g2_a22oi_1 _22868_ (.Y(_06261_),
    .B1(_06091_),
    .B2(\top_ihp.oisc.regs[21][17] ),
    .A2(net801),
    .A1(_08005_));
 sg13g2_o21ai_1 _22869_ (.B1(_06261_),
    .Y(_06262_),
    .A1(_05418_),
    .A2(_06260_));
 sg13g2_a21oi_1 _22870_ (.A1(\top_ihp.oisc.regs[61][17] ),
    .A2(net175),
    .Y(_06263_),
    .B1(_06262_));
 sg13g2_a22oi_1 _22871_ (.Y(_06264_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[27][17] ),
    .A2(net192),
    .A1(\top_ihp.oisc.regs[62][17] ));
 sg13g2_nand3_1 _22872_ (.B(_06263_),
    .C(_06264_),
    .A(_06259_),
    .Y(_06265_));
 sg13g2_a22oi_1 _22873_ (.Y(_06266_),
    .B1(net172),
    .B2(\top_ihp.oisc.regs[17][17] ),
    .A2(net430),
    .A1(\top_ihp.oisc.regs[14][17] ));
 sg13g2_a22oi_1 _22874_ (.Y(_06267_),
    .B1(net535),
    .B2(\top_ihp.oisc.regs[28][17] ),
    .A2(net163),
    .A1(\top_ihp.oisc.regs[4][17] ));
 sg13g2_nor2_1 _22875_ (.A(_05535_),
    .B(net748),
    .Y(_06268_));
 sg13g2_mux2_1 _22876_ (.A0(\top_ihp.oisc.regs[26][17] ),
    .A1(\top_ihp.oisc.regs[24][17] ),
    .S(net669),
    .X(_06269_));
 sg13g2_a22oi_1 _22877_ (.Y(_06270_),
    .B1(_06268_),
    .B2(_06269_),
    .A2(net380),
    .A1(\top_ihp.oisc.regs[11][17] ));
 sg13g2_buf_1 _22878_ (.A(net543),
    .X(_06271_));
 sg13g2_a22oi_1 _22879_ (.Y(_06272_),
    .B1(net164),
    .B2(\top_ihp.oisc.regs[9][17] ),
    .A2(net335),
    .A1(\top_ihp.oisc.regs[19][17] ));
 sg13g2_nand4_1 _22880_ (.B(_06267_),
    .C(_06270_),
    .A(_06266_),
    .Y(_06273_),
    .D(_06272_));
 sg13g2_a22oi_1 _22881_ (.Y(_06274_),
    .B1(net536),
    .B2(\top_ihp.oisc.regs[8][17] ),
    .A2(net373),
    .A1(\top_ihp.oisc.regs[1][17] ));
 sg13g2_a22oi_1 _22882_ (.Y(_06275_),
    .B1(net181),
    .B2(\top_ihp.oisc.regs[15][17] ),
    .A2(net166),
    .A1(\top_ihp.oisc.regs[3][17] ));
 sg13g2_buf_1 _22883_ (.A(net537),
    .X(_06276_));
 sg13g2_nor2_2 _22884_ (.A(net672),
    .B(net748),
    .Y(_06277_));
 sg13g2_and3_1 _22885_ (.X(_06278_),
    .A(\top_ihp.oisc.regs[16][17] ),
    .B(net662),
    .C(_06277_));
 sg13g2_a221oi_1 _22886_ (.B2(\top_ihp.oisc.regs[10][17] ),
    .C1(_06278_),
    .B1(net334),
    .A1(\top_ihp.oisc.regs[39][17] ),
    .Y(_06279_),
    .A2(_06143_));
 sg13g2_nand3_1 _22887_ (.B(_06275_),
    .C(_06279_),
    .A(_06274_),
    .Y(_06280_));
 sg13g2_a22oi_1 _22888_ (.Y(_06281_),
    .B1(net386),
    .B2(\top_ihp.oisc.regs[49][17] ),
    .A2(_05618_),
    .A1(\top_ihp.oisc.regs[34][17] ));
 sg13g2_a22oi_1 _22889_ (.Y(_06282_),
    .B1(_05800_),
    .B2(\top_ihp.oisc.regs[41][17] ),
    .A2(_05839_),
    .A1(\top_ihp.oisc.regs[47][17] ));
 sg13g2_a22oi_1 _22890_ (.Y(_06283_),
    .B1(_05935_),
    .B2(\top_ihp.oisc.regs[35][17] ),
    .A2(net348),
    .A1(\top_ihp.oisc.regs[57][17] ));
 sg13g2_a22oi_1 _22891_ (.Y(_06284_),
    .B1(net197),
    .B2(\top_ihp.oisc.regs[48][17] ),
    .A2(net178),
    .A1(\top_ihp.oisc.regs[54][17] ));
 sg13g2_nand4_1 _22892_ (.B(_06282_),
    .C(_06283_),
    .A(_06281_),
    .Y(_06285_),
    .D(_06284_));
 sg13g2_nor4_1 _22893_ (.A(_06265_),
    .B(_06273_),
    .C(_06280_),
    .D(_06285_),
    .Y(_06286_));
 sg13g2_a22oi_1 _22894_ (.Y(_06287_),
    .B1(_05670_),
    .B2(\top_ihp.oisc.regs[43][17] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[40][17] ));
 sg13g2_a22oi_1 _22895_ (.Y(_06288_),
    .B1(_05864_),
    .B2(\top_ihp.oisc.regs[38][17] ),
    .A2(net186),
    .A1(\top_ihp.oisc.regs[59][17] ));
 sg13g2_a22oi_1 _22896_ (.Y(_06289_),
    .B1(net391),
    .B2(\top_ihp.oisc.regs[33][17] ),
    .A2(net389),
    .A1(\top_ihp.oisc.regs[31][17] ));
 sg13g2_a22oi_1 _22897_ (.Y(_06290_),
    .B1(net347),
    .B2(\top_ihp.oisc.regs[37][17] ),
    .A2(net416),
    .A1(\top_ihp.oisc.regs[42][17] ));
 sg13g2_nand4_1 _22898_ (.B(_06288_),
    .C(_06289_),
    .A(_06287_),
    .Y(_06291_),
    .D(_06290_));
 sg13g2_a22oi_1 _22899_ (.Y(_06292_),
    .B1(net189),
    .B2(\top_ihp.oisc.regs[60][17] ),
    .A2(_05949_),
    .A1(\top_ihp.oisc.regs[55][17] ));
 sg13g2_a22oi_1 _22900_ (.Y(_06293_),
    .B1(_05867_),
    .B2(\top_ihp.oisc.regs[56][17] ),
    .A2(net400),
    .A1(\top_ihp.oisc.regs[63][17] ));
 sg13g2_a22oi_1 _22901_ (.Y(_06294_),
    .B1(net392),
    .B2(\top_ihp.oisc.regs[52][17] ),
    .A2(_05625_),
    .A1(\top_ihp.oisc.regs[51][17] ));
 sg13g2_a22oi_1 _22902_ (.Y(_06295_),
    .B1(net379),
    .B2(\top_ihp.oisc.regs[45][17] ),
    .A2(_05872_),
    .A1(\top_ihp.oisc.regs[36][17] ));
 sg13g2_nand4_1 _22903_ (.B(_06293_),
    .C(_06294_),
    .A(_06292_),
    .Y(_06296_),
    .D(_06295_));
 sg13g2_and3_1 _22904_ (.X(_06297_),
    .A(_05371_),
    .B(_05492_),
    .C(net722));
 sg13g2_a22oi_1 _22905_ (.Y(_06298_),
    .B1(_06297_),
    .B2(\top_ihp.oisc.regs[25][17] ),
    .A2(_06018_),
    .A1(\top_ihp.oisc.regs[46][17] ));
 sg13g2_a22oi_1 _22906_ (.Y(_06299_),
    .B1(net202),
    .B2(\top_ihp.oisc.regs[44][17] ),
    .A2(net199),
    .A1(\top_ihp.oisc.regs[50][17] ));
 sg13g2_a22oi_1 _22907_ (.Y(_06300_),
    .B1(net177),
    .B2(\top_ihp.oisc.regs[58][17] ),
    .A2(_05615_),
    .A1(\top_ihp.oisc.regs[32][17] ));
 sg13g2_a22oi_1 _22908_ (.Y(_06301_),
    .B1(net388),
    .B2(\top_ihp.oisc.regs[30][17] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[53][17] ));
 sg13g2_nand4_1 _22909_ (.B(_06299_),
    .C(_06300_),
    .A(_06298_),
    .Y(_06302_),
    .D(_06301_));
 sg13g2_nor4_2 _22910_ (.A(_05708_),
    .B(_06291_),
    .C(_06296_),
    .Y(_06303_),
    .D(_06302_));
 sg13g2_buf_1 _22911_ (.A(net783),
    .X(_06304_));
 sg13g2_nand2_1 _22912_ (.Y(_06305_),
    .A(_00221_),
    .B(net60));
 sg13g2_a22oi_1 _22913_ (.Y(_06306_),
    .B1(net26),
    .B2(_06305_),
    .A2(net746),
    .A1(_08005_));
 sg13g2_a21oi_1 _22914_ (.A1(_06286_),
    .A2(_06303_),
    .Y(_00396_),
    .B1(_06306_));
 sg13g2_a22oi_1 _22915_ (.Y(_06307_),
    .B1(_06018_),
    .B2(\top_ihp.oisc.regs[46][18] ),
    .A2(net539),
    .A1(\top_ihp.oisc.regs[34][18] ));
 sg13g2_a22oi_1 _22916_ (.Y(_06308_),
    .B1(net392),
    .B2(\top_ihp.oisc.regs[52][18] ),
    .A2(net174),
    .A1(\top_ihp.oisc.regs[62][18] ));
 sg13g2_a22oi_1 _22917_ (.Y(_06309_),
    .B1(_05733_),
    .B2(\top_ihp.oisc.regs[49][18] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[39][18] ));
 sg13g2_buf_1 _22918_ (.A(_05640_),
    .X(_06310_));
 sg13g2_a22oi_1 _22919_ (.Y(_06311_),
    .B1(net178),
    .B2(\top_ihp.oisc.regs[54][18] ),
    .A2(net333),
    .A1(\top_ihp.oisc.regs[57][18] ));
 sg13g2_nand4_1 _22920_ (.B(_06308_),
    .C(_06309_),
    .A(_06307_),
    .Y(_06312_),
    .D(_06311_));
 sg13g2_a22oi_1 _22921_ (.Y(_06313_),
    .B1(net376),
    .B2(\top_ihp.oisc.regs[51][18] ),
    .A2(net357),
    .A1(\top_ihp.oisc.regs[36][18] ));
 sg13g2_a22oi_1 _22922_ (.Y(_06314_),
    .B1(_05861_),
    .B2(\top_ihp.oisc.regs[45][18] ),
    .A2(net393),
    .A1(\top_ihp.oisc.regs[42][18] ));
 sg13g2_a22oi_1 _22923_ (.Y(_06315_),
    .B1(net383),
    .B2(\top_ihp.oisc.regs[60][18] ),
    .A2(net341),
    .A1(\top_ihp.oisc.regs[27][18] ));
 sg13g2_nand2_1 _22924_ (.Y(_06316_),
    .A(\top_ihp.oisc.regs[28][18] ),
    .B(_05543_));
 sg13g2_a22oi_1 _22925_ (.Y(_06317_),
    .B1(_05970_),
    .B2(\top_ihp.oisc.regs[23][18] ),
    .A2(net801),
    .A1(net1070));
 sg13g2_nand2_1 _22926_ (.Y(_06318_),
    .A(_06316_),
    .B(_06317_));
 sg13g2_a21oi_1 _22927_ (.A1(\top_ihp.oisc.regs[48][18] ),
    .A2(net409),
    .Y(_06319_),
    .B1(_06318_));
 sg13g2_nand4_1 _22928_ (.B(_06314_),
    .C(_06315_),
    .A(_06313_),
    .Y(_06320_),
    .D(_06319_));
 sg13g2_a22oi_1 _22929_ (.Y(_06321_),
    .B1(_05526_),
    .B2(\top_ihp.oisc.regs[12][18] ),
    .A2(_05373_),
    .A1(\top_ihp.oisc.regs[21][18] ));
 sg13g2_or2_1 _22930_ (.X(_06322_),
    .B(_06321_),
    .A(net672));
 sg13g2_nand3_1 _22931_ (.B(net550),
    .C(net747),
    .A(\top_ihp.oisc.regs[14][18] ),
    .Y(_06323_));
 sg13g2_a21oi_1 _22932_ (.A1(_06322_),
    .A2(_06323_),
    .Y(_06324_),
    .B1(net541));
 sg13g2_a221oi_1 _22933_ (.B2(\top_ihp.oisc.regs[5][18] ),
    .C1(_06324_),
    .B1(net345),
    .A1(\top_ihp.oisc.regs[11][18] ),
    .Y(_06325_),
    .A2(net380));
 sg13g2_a22oi_1 _22934_ (.Y(_06326_),
    .B1(net432),
    .B2(\top_ihp.oisc.regs[4][18] ),
    .A2(net553),
    .A1(\top_ihp.oisc.regs[22][18] ));
 sg13g2_a22oi_1 _22935_ (.Y(_06327_),
    .B1(_05750_),
    .B2(\top_ihp.oisc.regs[2][18] ),
    .A2(net544),
    .A1(\top_ihp.oisc.regs[18][18] ));
 sg13g2_and2_1 _22936_ (.A(_06326_),
    .B(_06327_),
    .X(_06328_));
 sg13g2_a22oi_1 _22937_ (.Y(_06329_),
    .B1(net193),
    .B2(\top_ihp.oisc.regs[56][18] ),
    .A2(net359),
    .A1(\top_ihp.oisc.regs[55][18] ));
 sg13g2_a22oi_1 _22938_ (.Y(_06330_),
    .B1(_06139_),
    .B2(\top_ihp.oisc.regs[38][18] ),
    .A2(net346),
    .A1(\top_ihp.oisc.regs[30][18] ));
 sg13g2_nand4_1 _22939_ (.B(_06328_),
    .C(_06329_),
    .A(_06325_),
    .Y(_06331_),
    .D(_06330_));
 sg13g2_a22oi_1 _22940_ (.Y(_06332_),
    .B1(_05935_),
    .B2(\top_ihp.oisc.regs[35][18] ),
    .A2(net191),
    .A1(\top_ihp.oisc.regs[59][18] ));
 sg13g2_a22oi_1 _22941_ (.Y(_06333_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[47][18] ),
    .A2(net190),
    .A1(\top_ihp.oisc.regs[61][18] ));
 sg13g2_a22oi_1 _22942_ (.Y(_06334_),
    .B1(net426),
    .B2(\top_ihp.oisc.regs[37][18] ),
    .A2(net194),
    .A1(\top_ihp.oisc.regs[50][18] ));
 sg13g2_a22oi_1 _22943_ (.Y(_06335_),
    .B1(net177),
    .B2(\top_ihp.oisc.regs[58][18] ),
    .A2(_06189_),
    .A1(\top_ihp.oisc.regs[44][18] ));
 sg13g2_nand4_1 _22944_ (.B(_06333_),
    .C(_06334_),
    .A(_06332_),
    .Y(_06336_),
    .D(_06335_));
 sg13g2_nor4_2 _22945_ (.A(_06312_),
    .B(_06320_),
    .C(_06331_),
    .Y(_06337_),
    .D(_06336_));
 sg13g2_a22oi_1 _22946_ (.Y(_06338_),
    .B1(net182),
    .B2(\top_ihp.oisc.regs[29][18] ),
    .A2(net438),
    .A1(\top_ihp.oisc.regs[7][18] ));
 sg13g2_a22oi_1 _22947_ (.Y(_06339_),
    .B1(net185),
    .B2(\top_ihp.oisc.regs[9][18] ),
    .A2(net170),
    .A1(\top_ihp.oisc.regs[3][18] ));
 sg13g2_mux2_1 _22948_ (.A0(\top_ihp.oisc.regs[24][18] ),
    .A1(\top_ihp.oisc.regs[16][18] ),
    .S(net662),
    .X(_06340_));
 sg13g2_a22oi_1 _22949_ (.Y(_06341_),
    .B1(_06340_),
    .B2(_06277_),
    .A2(net367),
    .A1(\top_ihp.oisc.regs[26][18] ));
 sg13g2_a22oi_1 _22950_ (.Y(_06342_),
    .B1(net334),
    .B2(\top_ihp.oisc.regs[10][18] ),
    .A2(net431),
    .A1(\top_ihp.oisc.regs[1][18] ));
 sg13g2_nand4_1 _22951_ (.B(_06339_),
    .C(_06341_),
    .A(_06338_),
    .Y(_06343_),
    .D(_06342_));
 sg13g2_a22oi_1 _22952_ (.Y(_06344_),
    .B1(net536),
    .B2(\top_ihp.oisc.regs[8][18] ),
    .A2(net667),
    .A1(\top_ihp.oisc.regs[6][18] ));
 sg13g2_a22oi_1 _22953_ (.Y(_06345_),
    .B1(_06246_),
    .B2(\top_ihp.oisc.regs[19][18] ),
    .A2(net160),
    .A1(\top_ihp.oisc.regs[17][18] ));
 sg13g2_a22oi_1 _22954_ (.Y(_06346_),
    .B1(net181),
    .B2(\top_ihp.oisc.regs[15][18] ),
    .A2(net540),
    .A1(\top_ihp.oisc.regs[20][18] ));
 sg13g2_and2_1 _22955_ (.A(\top_ihp.oisc.regs[13][18] ),
    .B(_05426_),
    .X(_06347_));
 sg13g2_nor4_1 _22956_ (.A(net541),
    .B(net550),
    .C(net662),
    .D(net726),
    .Y(_06348_));
 sg13g2_a22oi_1 _22957_ (.Y(_06349_),
    .B1(_06347_),
    .B2(_06348_),
    .A2(net368),
    .A1(\top_ihp.oisc.regs[25][18] ));
 sg13g2_nand4_1 _22958_ (.B(_06345_),
    .C(_06346_),
    .A(_06344_),
    .Y(_06350_),
    .D(_06349_));
 sg13g2_a22oi_1 _22959_ (.Y(_06351_),
    .B1(net407),
    .B2(\top_ihp.oisc.regs[33][18] ),
    .A2(net365),
    .A1(\top_ihp.oisc.regs[63][18] ));
 sg13g2_a22oi_1 _22960_ (.Y(_06352_),
    .B1(_05670_),
    .B2(\top_ihp.oisc.regs[43][18] ),
    .A2(_05960_),
    .A1(\top_ihp.oisc.regs[31][18] ));
 sg13g2_a22oi_1 _22961_ (.Y(_06353_),
    .B1(_05800_),
    .B2(\top_ihp.oisc.regs[41][18] ),
    .A2(net385),
    .A1(\top_ihp.oisc.regs[40][18] ));
 sg13g2_a22oi_1 _22962_ (.Y(_06354_),
    .B1(net363),
    .B2(\top_ihp.oisc.regs[32][18] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[53][18] ));
 sg13g2_nand4_1 _22963_ (.B(_06352_),
    .C(_06353_),
    .A(_06351_),
    .Y(_06355_),
    .D(_06354_));
 sg13g2_nor4_1 _22964_ (.A(net63),
    .B(_06343_),
    .C(_06350_),
    .D(_06355_),
    .Y(_06356_));
 sg13g2_nand2_1 _22965_ (.Y(_06357_),
    .A(_00222_),
    .B(net60));
 sg13g2_a22oi_1 _22966_ (.Y(_06358_),
    .B1(net26),
    .B2(_06357_),
    .A2(net746),
    .A1(_07995_));
 sg13g2_a21oi_1 _22967_ (.A1(_06337_),
    .A2(_06356_),
    .Y(_00397_),
    .B1(_06358_));
 sg13g2_nand2_1 _22968_ (.Y(_06359_),
    .A(\top_ihp.oisc.regs[58][19] ),
    .B(_05791_));
 sg13g2_a22oi_1 _22969_ (.Y(_06360_),
    .B1(_05861_),
    .B2(\top_ihp.oisc.regs[45][19] ),
    .A2(net389),
    .A1(\top_ihp.oisc.regs[31][19] ));
 sg13g2_a22oi_1 _22970_ (.Y(_06361_),
    .B1(_05795_),
    .B2(\top_ihp.oisc.regs[37][19] ),
    .A2(net352),
    .A1(\top_ihp.oisc.regs[43][19] ));
 sg13g2_a22oi_1 _22971_ (.Y(_06362_),
    .B1(net542),
    .B2(\top_ihp.oisc.regs[34][19] ),
    .A2(_05659_),
    .A1(\top_ihp.oisc.regs[30][19] ));
 sg13g2_nand4_1 _22972_ (.B(_06360_),
    .C(_06361_),
    .A(_06359_),
    .Y(_06363_),
    .D(_06362_));
 sg13g2_a22oi_1 _22973_ (.Y(_06364_),
    .B1(net189),
    .B2(\top_ihp.oisc.regs[60][19] ),
    .A2(net393),
    .A1(\top_ihp.oisc.regs[42][19] ));
 sg13g2_a22oi_1 _22974_ (.Y(_06365_),
    .B1(_05719_),
    .B2(\top_ihp.oisc.regs[35][19] ),
    .A2(net382),
    .A1(\top_ihp.oisc.regs[27][19] ));
 sg13g2_nand3_1 _22975_ (.B(_06364_),
    .C(_06365_),
    .A(net61),
    .Y(_06366_));
 sg13g2_nand2_1 _22976_ (.Y(_06367_),
    .A(_07999_),
    .B(net835));
 sg13g2_a22oi_1 _22977_ (.Y(_06368_),
    .B1(net719),
    .B2(\top_ihp.oisc.regs[23][19] ),
    .A2(_05820_),
    .A1(\top_ihp.oisc.regs[21][19] ));
 sg13g2_nand2_1 _22978_ (.Y(_06369_),
    .A(_06367_),
    .B(_06368_));
 sg13g2_a221oi_1 _22979_ (.B2(\top_ihp.oisc.regs[17][19] ),
    .C1(_06369_),
    .B1(net427),
    .A1(\top_ihp.oisc.regs[6][19] ),
    .Y(_06370_),
    .A2(net667));
 sg13g2_a22oi_1 _22980_ (.Y(_06371_),
    .B1(net197),
    .B2(\top_ihp.oisc.regs[48][19] ),
    .A2(net200),
    .A1(\top_ihp.oisc.regs[61][19] ));
 sg13g2_a22oi_1 _22981_ (.Y(_06372_),
    .B1(net376),
    .B2(\top_ihp.oisc.regs[51][19] ),
    .A2(_05864_),
    .A1(\top_ihp.oisc.regs[38][19] ));
 sg13g2_a22oi_1 _22982_ (.Y(_06373_),
    .B1(net340),
    .B2(\top_ihp.oisc.regs[41][19] ),
    .A2(_05875_),
    .A1(\top_ihp.oisc.regs[59][19] ));
 sg13g2_nand4_1 _22983_ (.B(_06371_),
    .C(_06372_),
    .A(_06370_),
    .Y(_06374_),
    .D(_06373_));
 sg13g2_a22oi_1 _22984_ (.Y(_06375_),
    .B1(net202),
    .B2(\top_ihp.oisc.regs[44][19] ),
    .A2(net357),
    .A1(\top_ihp.oisc.regs[36][19] ));
 sg13g2_a22oi_1 _22985_ (.Y(_06376_),
    .B1(net396),
    .B2(\top_ihp.oisc.regs[46][19] ),
    .A2(net348),
    .A1(\top_ihp.oisc.regs[57][19] ));
 sg13g2_a22oi_1 _22986_ (.Y(_06377_),
    .B1(net407),
    .B2(\top_ihp.oisc.regs[33][19] ),
    .A2(_05606_),
    .A1(\top_ihp.oisc.regs[39][19] ));
 sg13g2_a22oi_1 _22987_ (.Y(_06378_),
    .B1(net405),
    .B2(\top_ihp.oisc.regs[52][19] ),
    .A2(_05951_),
    .A1(\top_ihp.oisc.regs[47][19] ));
 sg13g2_nand4_1 _22988_ (.B(_06376_),
    .C(_06377_),
    .A(_06375_),
    .Y(_06379_),
    .D(_06378_));
 sg13g2_nor4_2 _22989_ (.A(_06363_),
    .B(_06366_),
    .C(_06374_),
    .Y(_06380_),
    .D(_06379_));
 sg13g2_a22oi_1 _22990_ (.Y(_06381_),
    .B1(net403),
    .B2(\top_ihp.oisc.regs[55][19] ),
    .A2(net351),
    .A1(\top_ihp.oisc.regs[40][19] ));
 sg13g2_a22oi_1 _22991_ (.Y(_06382_),
    .B1(_05863_),
    .B2(\top_ihp.oisc.regs[50][19] ),
    .A2(net377),
    .A1(\top_ihp.oisc.regs[53][19] ));
 sg13g2_a22oi_1 _22992_ (.Y(_06383_),
    .B1(net338),
    .B2(\top_ihp.oisc.regs[32][19] ),
    .A2(net174),
    .A1(\top_ihp.oisc.regs[62][19] ));
 sg13g2_a22oi_1 _22993_ (.Y(_06384_),
    .B1(_05804_),
    .B2(\top_ihp.oisc.regs[56][19] ),
    .A2(_05732_),
    .A1(\top_ihp.oisc.regs[49][19] ));
 sg13g2_nand4_1 _22994_ (.B(_06382_),
    .C(_06383_),
    .A(_06381_),
    .Y(_06385_),
    .D(_06384_));
 sg13g2_a22oi_1 _22995_ (.Y(_06386_),
    .B1(net371),
    .B2(\top_ihp.oisc.regs[16][19] ),
    .A2(net533),
    .A1(\top_ihp.oisc.regs[22][19] ));
 sg13g2_a22oi_1 _22996_ (.Y(_06387_),
    .B1(net374),
    .B2(\top_ihp.oisc.regs[9][19] ),
    .A2(net668),
    .A1(\top_ihp.oisc.regs[28][19] ));
 sg13g2_a22oi_1 _22997_ (.Y(_06388_),
    .B1(net428),
    .B2(\top_ihp.oisc.regs[15][19] ),
    .A2(net401),
    .A1(\top_ihp.oisc.regs[3][19] ));
 sg13g2_a22oi_1 _22998_ (.Y(_06389_),
    .B1(net665),
    .B2(\top_ihp.oisc.regs[8][19] ),
    .A2(_05765_),
    .A1(\top_ihp.oisc.regs[26][19] ));
 sg13g2_nand4_1 _22999_ (.B(_06387_),
    .C(_06388_),
    .A(_06386_),
    .Y(_06390_),
    .D(_06389_));
 sg13g2_a22oi_1 _23000_ (.Y(_06391_),
    .B1(net365),
    .B2(\top_ihp.oisc.regs[63][19] ),
    .A2(net196),
    .A1(\top_ihp.oisc.regs[54][19] ));
 sg13g2_nand2b_1 _23001_ (.Y(_06392_),
    .B(_06391_),
    .A_N(_06390_));
 sg13g2_a22oi_1 _23002_ (.Y(_06393_),
    .B1(net180),
    .B2(\top_ihp.oisc.regs[13][19] ),
    .A2(net335),
    .A1(\top_ihp.oisc.regs[19][19] ));
 sg13g2_a22oi_1 _23003_ (.Y(_06394_),
    .B1(net173),
    .B2(\top_ihp.oisc.regs[11][19] ),
    .A2(net203),
    .A1(\top_ihp.oisc.regs[29][19] ));
 sg13g2_a22oi_1 _23004_ (.Y(_06395_),
    .B1(net334),
    .B2(\top_ihp.oisc.regs[10][19] ),
    .A2(net540),
    .A1(\top_ihp.oisc.regs[20][19] ));
 sg13g2_a22oi_1 _23005_ (.Y(_06396_),
    .B1(net369),
    .B2(\top_ihp.oisc.regs[2][19] ),
    .A2(net368),
    .A1(\top_ihp.oisc.regs[25][19] ));
 sg13g2_nand4_1 _23006_ (.B(_06394_),
    .C(_06395_),
    .A(_06393_),
    .Y(_06397_),
    .D(_06396_));
 sg13g2_a22oi_1 _23007_ (.Y(_06398_),
    .B1(net167),
    .B2(\top_ihp.oisc.regs[24][19] ),
    .A2(net184),
    .A1(\top_ihp.oisc.regs[12][19] ));
 sg13g2_a22oi_1 _23008_ (.Y(_06399_),
    .B1(net373),
    .B2(\top_ihp.oisc.regs[1][19] ),
    .A2(net204),
    .A1(\top_ihp.oisc.regs[4][19] ));
 sg13g2_a22oi_1 _23009_ (.Y(_06400_),
    .B1(net165),
    .B2(\top_ihp.oisc.regs[5][19] ),
    .A2(net430),
    .A1(\top_ihp.oisc.regs[14][19] ));
 sg13g2_a22oi_1 _23010_ (.Y(_06401_),
    .B1(net343),
    .B2(\top_ihp.oisc.regs[18][19] ),
    .A2(net342),
    .A1(\top_ihp.oisc.regs[7][19] ));
 sg13g2_nand4_1 _23011_ (.B(_06399_),
    .C(_06400_),
    .A(_06398_),
    .Y(_06402_),
    .D(_06401_));
 sg13g2_nor4_1 _23012_ (.A(_06385_),
    .B(_06392_),
    .C(_06397_),
    .D(_06402_),
    .Y(_06403_));
 sg13g2_a21o_1 _23013_ (.A2(net63),
    .A1(_00223_),
    .B1(net58),
    .X(_06404_));
 sg13g2_a22oi_1 _23014_ (.Y(_00398_),
    .B1(_06404_),
    .B2(_06367_),
    .A2(_06403_),
    .A1(_06380_));
 sg13g2_a22oi_1 _23015_ (.Y(_06405_),
    .B1(net360),
    .B2(\top_ihp.oisc.regs[33][1] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[39][1] ));
 sg13g2_a22oi_1 _23016_ (.Y(_06406_),
    .B1(net340),
    .B2(\top_ihp.oisc.regs[41][1] ),
    .A2(net186),
    .A1(\top_ihp.oisc.regs[59][1] ));
 sg13g2_a22oi_1 _23017_ (.Y(_06407_),
    .B1(net187),
    .B2(\top_ihp.oisc.regs[56][1] ),
    .A2(net411),
    .A1(\top_ihp.oisc.regs[45][1] ));
 sg13g2_a22oi_1 _23018_ (.Y(_06408_),
    .B1(net353),
    .B2(\top_ihp.oisc.regs[35][1] ),
    .A2(_05608_),
    .A1(\top_ihp.oisc.regs[27][1] ));
 sg13g2_nand4_1 _23019_ (.B(_06406_),
    .C(_06407_),
    .A(_06405_),
    .Y(_06409_),
    .D(_06408_));
 sg13g2_a22oi_1 _23020_ (.Y(_06410_),
    .B1(net355),
    .B2(\top_ihp.oisc.regs[51][1] ),
    .A2(net358),
    .A1(\top_ihp.oisc.regs[47][1] ));
 sg13g2_a22oi_1 _23021_ (.Y(_06411_),
    .B1(net392),
    .B2(\top_ihp.oisc.regs[52][1] ),
    .A2(net338),
    .A1(\top_ihp.oisc.regs[32][1] ));
 sg13g2_nand3_1 _23022_ (.B(_06410_),
    .C(_06411_),
    .A(net61),
    .Y(_06412_));
 sg13g2_a22oi_1 _23023_ (.Y(_06413_),
    .B1(net396),
    .B2(\top_ihp.oisc.regs[46][1] ),
    .A2(net199),
    .A1(\top_ihp.oisc.regs[50][1] ));
 sg13g2_a22oi_1 _23024_ (.Y(_06414_),
    .B1(net176),
    .B2(\top_ihp.oisc.regs[62][1] ),
    .A2(net178),
    .A1(\top_ihp.oisc.regs[54][1] ));
 sg13g2_a22oi_1 _23025_ (.Y(_06415_),
    .B1(net161),
    .B2(\top_ihp.oisc.regs[44][1] ),
    .A2(net413),
    .A1(\top_ihp.oisc.regs[63][1] ));
 sg13g2_a22oi_1 _23026_ (.Y(_06416_),
    .B1(net339),
    .B2(\top_ihp.oisc.regs[38][1] ),
    .A2(net414),
    .A1(\top_ihp.oisc.regs[30][1] ));
 sg13g2_nand4_1 _23027_ (.B(_06414_),
    .C(_06415_),
    .A(_06413_),
    .Y(_06417_),
    .D(_06416_));
 sg13g2_a22oi_1 _23028_ (.Y(_06418_),
    .B1(net412),
    .B2(\top_ihp.oisc.regs[43][1] ),
    .A2(net344),
    .A1(\top_ihp.oisc.regs[53][1] ));
 sg13g2_a22oi_1 _23029_ (.Y(_06419_),
    .B1(net398),
    .B2(\top_ihp.oisc.regs[55][1] ),
    .A2(net190),
    .A1(\top_ihp.oisc.regs[61][1] ));
 sg13g2_a22oi_1 _23030_ (.Y(_06420_),
    .B1(net197),
    .B2(\top_ihp.oisc.regs[48][1] ),
    .A2(net356),
    .A1(\top_ihp.oisc.regs[31][1] ));
 sg13g2_a22oi_1 _23031_ (.Y(_06421_),
    .B1(net177),
    .B2(\top_ihp.oisc.regs[58][1] ),
    .A2(net417),
    .A1(\top_ihp.oisc.regs[57][1] ));
 sg13g2_nand4_1 _23032_ (.B(_06419_),
    .C(_06420_),
    .A(_06418_),
    .Y(_06422_),
    .D(_06421_));
 sg13g2_nor4_2 _23033_ (.A(_06409_),
    .B(_06412_),
    .C(_06417_),
    .Y(_06423_),
    .D(_06422_));
 sg13g2_nand2_1 _23034_ (.Y(_06424_),
    .A(\top_ihp.oisc.regs[8][1] ),
    .B(net536));
 sg13g2_a22oi_1 _23035_ (.Y(_06425_),
    .B1(net184),
    .B2(\top_ihp.oisc.regs[12][1] ),
    .A2(net534),
    .A1(\top_ihp.oisc.regs[18][1] ));
 sg13g2_nor2_2 _23036_ (.A(_05554_),
    .B(net774),
    .Y(_06426_));
 sg13g2_a22oi_1 _23037_ (.Y(_06427_),
    .B1(_06426_),
    .B2(\top_ihp.oisc.regs[10][1] ),
    .A2(_05428_),
    .A1(\top_ihp.oisc.regs[7][1] ));
 sg13g2_a22oi_1 _23038_ (.Y(_06428_),
    .B1(_05578_),
    .B2(\top_ihp.oisc.regs[11][1] ),
    .A2(_05538_),
    .A1(\top_ihp.oisc.regs[24][1] ));
 sg13g2_a22oi_1 _23039_ (.Y(_06429_),
    .B1(_05765_),
    .B2(\top_ihp.oisc.regs[26][1] ),
    .A2(_05761_),
    .A1(\top_ihp.oisc.regs[5][1] ));
 sg13g2_a22oi_1 _23040_ (.Y(_06430_),
    .B1(_05759_),
    .B2(\top_ihp.oisc.regs[16][1] ),
    .A2(_05559_),
    .A1(\top_ihp.oisc.regs[13][1] ));
 sg13g2_and4_1 _23041_ (.A(_06427_),
    .B(_06428_),
    .C(_06429_),
    .D(_06430_),
    .X(_06431_));
 sg13g2_nand3_1 _23042_ (.B(_06425_),
    .C(_06431_),
    .A(_06424_),
    .Y(_06432_));
 sg13g2_a22oi_1 _23043_ (.Y(_06433_),
    .B1(net366),
    .B2(\top_ihp.oisc.regs[49][1] ),
    .A2(net542),
    .A1(\top_ihp.oisc.regs[34][1] ));
 sg13g2_and2_1 _23044_ (.A(\top_ihp.oisc.regs[28][1] ),
    .B(net668),
    .X(_06434_));
 sg13g2_a221oi_1 _23045_ (.B2(\top_ihp.oisc.regs[14][1] ),
    .C1(_06434_),
    .B1(net546),
    .A1(\top_ihp.oisc.regs[20][1] ),
    .Y(_06435_),
    .A2(net540));
 sg13g2_a22oi_1 _23046_ (.Y(_06436_),
    .B1(net418),
    .B2(\top_ihp.oisc.regs[40][1] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[36][1] ));
 sg13g2_a22oi_1 _23047_ (.Y(_06437_),
    .B1(net393),
    .B2(\top_ihp.oisc.regs[42][1] ),
    .A2(_05588_),
    .A1(\top_ihp.oisc.regs[60][1] ));
 sg13g2_nand4_1 _23048_ (.B(_06435_),
    .C(_06436_),
    .A(_06433_),
    .Y(_06438_),
    .D(_06437_));
 sg13g2_a22oi_1 _23049_ (.Y(_06439_),
    .B1(net179),
    .B2(\top_ihp.oisc.regs[2][1] ),
    .A2(net162),
    .A1(\top_ihp.oisc.regs[15][1] ));
 sg13g2_a22oi_1 _23050_ (.Y(_06440_),
    .B1(net538),
    .B2(\top_ihp.oisc.regs[6][1] ),
    .A2(net163),
    .A1(\top_ihp.oisc.regs[4][1] ));
 sg13g2_a22oi_1 _23051_ (.Y(_06441_),
    .B1(net160),
    .B2(\top_ihp.oisc.regs[17][1] ),
    .A2(net368),
    .A1(\top_ihp.oisc.regs[25][1] ));
 sg13g2_a22oi_1 _23052_ (.Y(_06442_),
    .B1(net335),
    .B2(\top_ihp.oisc.regs[19][1] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[29][1] ));
 sg13g2_nand4_1 _23053_ (.B(_06440_),
    .C(_06441_),
    .A(_06439_),
    .Y(_06443_),
    .D(_06442_));
 sg13g2_a22oi_1 _23054_ (.Y(_06444_),
    .B1(net166),
    .B2(\top_ihp.oisc.regs[3][1] ),
    .A2(net373),
    .A1(\top_ihp.oisc.regs[1][1] ));
 sg13g2_a22oi_1 _23055_ (.Y(_06445_),
    .B1(net185),
    .B2(\top_ihp.oisc.regs[9][1] ),
    .A2(_05440_),
    .A1(\top_ihp.oisc.regs[22][1] ));
 sg13g2_nand2_1 _23056_ (.Y(_06446_),
    .A(_08078_),
    .B(_06023_));
 sg13g2_a22oi_1 _23057_ (.Y(_06447_),
    .B1(net719),
    .B2(\top_ihp.oisc.regs[23][1] ),
    .A2(net663),
    .A1(\top_ihp.oisc.regs[21][1] ));
 sg13g2_nand2_1 _23058_ (.Y(_06448_),
    .A(_06446_),
    .B(_06447_));
 sg13g2_a21oi_1 _23059_ (.A1(\top_ihp.oisc.regs[37][1] ),
    .A2(net426),
    .Y(_06449_),
    .B1(_06448_));
 sg13g2_nand3_1 _23060_ (.B(_06445_),
    .C(_06449_),
    .A(_06444_),
    .Y(_06450_));
 sg13g2_nor4_1 _23061_ (.A(_06432_),
    .B(_06438_),
    .C(_06443_),
    .D(_06450_),
    .Y(_06451_));
 sg13g2_inv_1 _23062_ (.Y(_06452_),
    .A(_00205_));
 sg13g2_o21ai_1 _23063_ (.B1(net27),
    .Y(_06453_),
    .A1(_06452_),
    .A2(net62));
 sg13g2_a22oi_1 _23064_ (.Y(_00399_),
    .B1(_06453_),
    .B2(_06446_),
    .A2(_06451_),
    .A1(_06423_));
 sg13g2_a22oi_1 _23065_ (.Y(_06454_),
    .B1(net363),
    .B2(\top_ihp.oisc.regs[32][20] ),
    .A2(net201),
    .A1(\top_ihp.oisc.regs[54][20] ));
 sg13g2_a22oi_1 _23066_ (.Y(_06455_),
    .B1(net344),
    .B2(\top_ihp.oisc.regs[53][20] ),
    .A2(net389),
    .A1(\top_ihp.oisc.regs[31][20] ));
 sg13g2_a22oi_1 _23067_ (.Y(_06456_),
    .B1(_05867_),
    .B2(\top_ihp.oisc.regs[56][20] ),
    .A2(_05735_),
    .A1(\top_ihp.oisc.regs[55][20] ));
 sg13g2_a22oi_1 _23068_ (.Y(_06457_),
    .B1(_05929_),
    .B2(\top_ihp.oisc.regs[52][20] ),
    .A2(_05681_),
    .A1(\top_ihp.oisc.regs[45][20] ));
 sg13g2_nand4_1 _23069_ (.B(_06455_),
    .C(_06456_),
    .A(_06454_),
    .Y(_06458_),
    .D(_06457_));
 sg13g2_a22oi_1 _23070_ (.Y(_06459_),
    .B1(net376),
    .B2(\top_ihp.oisc.regs[51][20] ),
    .A2(_05677_),
    .A1(\top_ihp.oisc.regs[50][20] ));
 sg13g2_a22oi_1 _23071_ (.Y(_06460_),
    .B1(_05606_),
    .B2(\top_ihp.oisc.regs[39][20] ),
    .A2(net192),
    .A1(\top_ihp.oisc.regs[62][20] ));
 sg13g2_a22oi_1 _23072_ (.Y(_06461_),
    .B1(_05795_),
    .B2(\top_ihp.oisc.regs[37][20] ),
    .A2(_05645_),
    .A1(\top_ihp.oisc.regs[42][20] ));
 sg13g2_nand2_1 _23073_ (.Y(_06462_),
    .A(net723),
    .B(_05433_));
 sg13g2_a22oi_1 _23074_ (.Y(_06463_),
    .B1(_05701_),
    .B2(\top_ihp.oisc.regs[16][20] ),
    .A2(net721),
    .A1(\top_ihp.oisc.regs[22][20] ));
 sg13g2_nor2_1 _23075_ (.A(_06462_),
    .B(_06463_),
    .Y(_06464_));
 sg13g2_a21oi_1 _23076_ (.A1(\top_ihp.oisc.regs[33][20] ),
    .A2(_05814_),
    .Y(_06465_),
    .B1(_06464_));
 sg13g2_nand4_1 _23077_ (.B(_06460_),
    .C(_06461_),
    .A(_06459_),
    .Y(_06466_),
    .D(_06465_));
 sg13g2_a22oi_1 _23078_ (.Y(_06467_),
    .B1(_05629_),
    .B2(\top_ihp.oisc.regs[44][20] ),
    .A2(_06139_),
    .A1(\top_ihp.oisc.regs[38][20] ));
 sg13g2_a22oi_1 _23079_ (.Y(_06468_),
    .B1(net412),
    .B2(\top_ihp.oisc.regs[43][20] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[40][20] ));
 sg13g2_a22oi_1 _23080_ (.Y(_06469_),
    .B1(net410),
    .B2(\top_ihp.oisc.regs[41][20] ),
    .A2(_05684_),
    .A1(\top_ihp.oisc.regs[59][20] ));
 sg13g2_a22oi_1 _23081_ (.Y(_06470_),
    .B1(net171),
    .B2(\top_ihp.oisc.regs[60][20] ),
    .A2(_05714_),
    .A1(\top_ihp.oisc.regs[48][20] ));
 sg13g2_nand4_1 _23082_ (.B(_06468_),
    .C(_06469_),
    .A(_06467_),
    .Y(_06471_),
    .D(_06470_));
 sg13g2_nand2_1 _23083_ (.Y(_06472_),
    .A(\top_ihp.oisc.regs[49][20] ),
    .B(net386));
 sg13g2_a22oi_1 _23084_ (.Y(_06473_),
    .B1(_05796_),
    .B2(\top_ihp.oisc.regs[46][20] ),
    .A2(_05602_),
    .A1(\top_ihp.oisc.regs[47][20] ));
 sg13g2_nand3_1 _23085_ (.B(_06472_),
    .C(_06473_),
    .A(_05742_),
    .Y(_06474_));
 sg13g2_nor4_2 _23086_ (.A(_06458_),
    .B(_06466_),
    .C(_06471_),
    .Y(_06475_),
    .D(_06474_));
 sg13g2_a22oi_1 _23087_ (.Y(_06476_),
    .B1(_05924_),
    .B2(\top_ihp.oisc.regs[58][20] ),
    .A2(net375),
    .A1(\top_ihp.oisc.regs[36][20] ));
 sg13g2_a22oi_1 _23088_ (.Y(_06477_),
    .B1(net353),
    .B2(\top_ihp.oisc.regs[35][20] ),
    .A2(net413),
    .A1(\top_ihp.oisc.regs[63][20] ));
 sg13g2_a22oi_1 _23089_ (.Y(_06478_),
    .B1(net539),
    .B2(\top_ihp.oisc.regs[34][20] ),
    .A2(net341),
    .A1(\top_ihp.oisc.regs[27][20] ));
 sg13g2_a22oi_1 _23090_ (.Y(_06479_),
    .B1(_06042_),
    .B2(\top_ihp.oisc.regs[30][20] ),
    .A2(net333),
    .A1(\top_ihp.oisc.regs[57][20] ));
 sg13g2_nand4_1 _23091_ (.B(_06477_),
    .C(_06478_),
    .A(_06476_),
    .Y(_06480_),
    .D(_06479_));
 sg13g2_a22oi_1 _23092_ (.Y(_06481_),
    .B1(net536),
    .B2(\top_ihp.oisc.regs[8][20] ),
    .A2(net334),
    .A1(\top_ihp.oisc.regs[10][20] ));
 sg13g2_a22oi_1 _23093_ (.Y(_06482_),
    .B1(_06102_),
    .B2(\top_ihp.oisc.regs[24][20] ),
    .A2(net431),
    .A1(\top_ihp.oisc.regs[1][20] ));
 sg13g2_mux2_1 _23094_ (.A0(\top_ihp.oisc.regs[14][20] ),
    .A1(\top_ihp.oisc.regs[12][20] ),
    .S(net669),
    .X(_06483_));
 sg13g2_nor2_2 _23095_ (.A(net670),
    .B(net774),
    .Y(_06484_));
 sg13g2_a22oi_1 _23096_ (.Y(_06485_),
    .B1(_06483_),
    .B2(_06484_),
    .A2(net368),
    .A1(\top_ihp.oisc.regs[25][20] ));
 sg13g2_a22oi_1 _23097_ (.Y(_06486_),
    .B1(_06149_),
    .B2(\top_ihp.oisc.regs[9][20] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[29][20] ));
 sg13g2_nand4_1 _23098_ (.B(_06482_),
    .C(_06485_),
    .A(_06481_),
    .Y(_06487_),
    .D(_06486_));
 sg13g2_a22oi_1 _23099_ (.Y(_06488_),
    .B1(_06106_),
    .B2(\top_ihp.oisc.regs[3][20] ),
    .A2(net350),
    .A1(\top_ihp.oisc.regs[19][20] ));
 sg13g2_a22oi_1 _23100_ (.Y(_06489_),
    .B1(_06068_),
    .B2(\top_ihp.oisc.regs[26][20] ),
    .A2(net369),
    .A1(\top_ihp.oisc.regs[2][20] ));
 sg13g2_nand2_1 _23101_ (.Y(_06490_),
    .A(\top_ihp.oisc.regs[61][20] ),
    .B(net190));
 sg13g2_and2_1 _23102_ (.A(_07990_),
    .B(net803),
    .X(_06491_));
 sg13g2_a221oi_1 _23103_ (.B2(\top_ihp.oisc.regs[23][20] ),
    .C1(_06491_),
    .B1(net720),
    .A1(\top_ihp.oisc.regs[21][20] ),
    .Y(_06492_),
    .A2(net666));
 sg13g2_nand4_1 _23104_ (.B(_06489_),
    .C(_06490_),
    .A(_06488_),
    .Y(_06493_),
    .D(_06492_));
 sg13g2_a22oi_1 _23105_ (.Y(_06494_),
    .B1(net428),
    .B2(\top_ihp.oisc.regs[15][20] ),
    .A2(_06057_),
    .A1(\top_ihp.oisc.regs[28][20] ));
 sg13g2_a22oi_1 _23106_ (.Y(_06495_),
    .B1(_06046_),
    .B2(\top_ihp.oisc.regs[5][20] ),
    .A2(net427),
    .A1(\top_ihp.oisc.regs[17][20] ));
 sg13g2_a22oi_1 _23107_ (.Y(_06496_),
    .B1(net370),
    .B2(\top_ihp.oisc.regs[13][20] ),
    .A2(net544),
    .A1(\top_ihp.oisc.regs[18][20] ));
 sg13g2_a22oi_1 _23108_ (.Y(_06497_),
    .B1(net667),
    .B2(\top_ihp.oisc.regs[6][20] ),
    .A2(_05429_),
    .A1(\top_ihp.oisc.regs[7][20] ));
 sg13g2_and4_1 _23109_ (.A(_06494_),
    .B(_06495_),
    .C(_06496_),
    .D(_06497_),
    .X(_06498_));
 sg13g2_nand2_1 _23110_ (.Y(_06499_),
    .A(\top_ihp.oisc.regs[20][20] ),
    .B(_05473_));
 sg13g2_a22oi_1 _23111_ (.Y(_06500_),
    .B1(_06066_),
    .B2(\top_ihp.oisc.regs[11][20] ),
    .A2(_05501_),
    .A1(\top_ihp.oisc.regs[4][20] ));
 sg13g2_nand3_1 _23112_ (.B(_06499_),
    .C(_06500_),
    .A(_06498_),
    .Y(_06501_));
 sg13g2_nor4_1 _23113_ (.A(_06480_),
    .B(_06487_),
    .C(_06493_),
    .D(_06501_),
    .Y(_06502_));
 sg13g2_a21oi_1 _23114_ (.A1(_00224_),
    .A2(net59),
    .Y(_06503_),
    .B1(_06009_));
 sg13g2_nor2_1 _23115_ (.A(_06491_),
    .B(_06503_),
    .Y(_06504_));
 sg13g2_a21oi_1 _23116_ (.A1(_06475_),
    .A2(_06502_),
    .Y(_00400_),
    .B1(_06504_));
 sg13g2_nand2_1 _23117_ (.Y(_06505_),
    .A(_08169_),
    .B(net801));
 sg13g2_a21o_1 _23118_ (.A2(net63),
    .A1(_00225_),
    .B1(net58),
    .X(_06506_));
 sg13g2_a22oi_1 _23119_ (.Y(_06507_),
    .B1(_05602_),
    .B2(\top_ihp.oisc.regs[47][21] ),
    .A2(net175),
    .A1(\top_ihp.oisc.regs[61][21] ));
 sg13g2_a22oi_1 _23120_ (.Y(_06508_),
    .B1(net187),
    .B2(\top_ihp.oisc.regs[56][21] ),
    .A2(_06040_),
    .A1(\top_ihp.oisc.regs[37][21] ));
 sg13g2_a22oi_1 _23121_ (.Y(_06509_),
    .B1(net406),
    .B2(\top_ihp.oisc.regs[46][21] ),
    .A2(net353),
    .A1(\top_ihp.oisc.regs[35][21] ));
 sg13g2_a22oi_1 _23122_ (.Y(_06510_),
    .B1(net399),
    .B2(\top_ihp.oisc.regs[58][21] ),
    .A2(_05665_),
    .A1(\top_ihp.oisc.regs[63][21] ));
 sg13g2_nand4_1 _23123_ (.B(_06508_),
    .C(_06509_),
    .A(_06507_),
    .Y(_06511_),
    .D(_06510_));
 sg13g2_a22oi_1 _23124_ (.Y(_06512_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[27][21] ),
    .A2(net385),
    .A1(\top_ihp.oisc.regs[40][21] ));
 sg13g2_a22oi_1 _23125_ (.Y(_06513_),
    .B1(net176),
    .B2(\top_ihp.oisc.regs[62][21] ),
    .A2(net348),
    .A1(\top_ihp.oisc.regs[57][21] ));
 sg13g2_nand3_1 _23126_ (.B(_06512_),
    .C(_06513_),
    .A(net57),
    .Y(_06514_));
 sg13g2_a22oi_1 _23127_ (.Y(_06515_),
    .B1(_05618_),
    .B2(\top_ihp.oisc.regs[34][21] ),
    .A2(net344),
    .A1(\top_ihp.oisc.regs[53][21] ));
 sg13g2_a22oi_1 _23128_ (.Y(_06516_),
    .B1(net355),
    .B2(\top_ihp.oisc.regs[51][21] ),
    .A2(net435),
    .A1(\top_ihp.oisc.regs[31][21] ));
 sg13g2_a22oi_1 _23129_ (.Y(_06517_),
    .B1(net412),
    .B2(\top_ihp.oisc.regs[43][21] ),
    .A2(net357),
    .A1(\top_ihp.oisc.regs[36][21] ));
 sg13g2_a22oi_1 _23130_ (.Y(_06518_),
    .B1(net392),
    .B2(\top_ihp.oisc.regs[52][21] ),
    .A2(net393),
    .A1(\top_ihp.oisc.regs[42][21] ));
 sg13g2_nand4_1 _23131_ (.B(_06516_),
    .C(_06517_),
    .A(_06515_),
    .Y(_06519_),
    .D(_06518_));
 sg13g2_a22oi_1 _23132_ (.Y(_06520_),
    .B1(net189),
    .B2(\top_ihp.oisc.regs[60][21] ),
    .A2(net394),
    .A1(\top_ihp.oisc.regs[45][21] ));
 sg13g2_a22oi_1 _23133_ (.Y(_06521_),
    .B1(net398),
    .B2(\top_ihp.oisc.regs[55][21] ),
    .A2(net407),
    .A1(\top_ihp.oisc.regs[33][21] ));
 sg13g2_a22oi_1 _23134_ (.Y(_06522_),
    .B1(_05844_),
    .B2(\top_ihp.oisc.regs[38][21] ),
    .A2(net194),
    .A1(\top_ihp.oisc.regs[50][21] ));
 sg13g2_a22oi_1 _23135_ (.Y(_06523_),
    .B1(net395),
    .B2(\top_ihp.oisc.regs[41][21] ),
    .A2(_06189_),
    .A1(\top_ihp.oisc.regs[44][21] ));
 sg13g2_nand4_1 _23136_ (.B(_06521_),
    .C(_06522_),
    .A(_06520_),
    .Y(_06524_),
    .D(_06523_));
 sg13g2_nor4_2 _23137_ (.A(_06511_),
    .B(_06514_),
    .C(_06519_),
    .Y(_06525_),
    .D(_06524_));
 sg13g2_a22oi_1 _23138_ (.Y(_06526_),
    .B1(net197),
    .B2(\top_ihp.oisc.regs[48][21] ),
    .A2(net178),
    .A1(\top_ihp.oisc.regs[54][21] ));
 sg13g2_a22oi_1 _23139_ (.Y(_06527_),
    .B1(net363),
    .B2(\top_ihp.oisc.regs[32][21] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[39][21] ));
 sg13g2_a22oi_1 _23140_ (.Y(_06528_),
    .B1(net366),
    .B2(\top_ihp.oisc.regs[49][21] ),
    .A2(net198),
    .A1(\top_ihp.oisc.regs[59][21] ));
 sg13g2_a22oi_1 _23141_ (.Y(_06529_),
    .B1(net719),
    .B2(\top_ihp.oisc.regs[23][21] ),
    .A2(net663),
    .A1(\top_ihp.oisc.regs[21][21] ));
 sg13g2_nand2_1 _23142_ (.Y(_06530_),
    .A(_06505_),
    .B(_06529_));
 sg13g2_a21oi_1 _23143_ (.A1(\top_ihp.oisc.regs[30][21] ),
    .A2(net346),
    .Y(_06531_),
    .B1(_06530_));
 sg13g2_nand4_1 _23144_ (.B(_06527_),
    .C(_06528_),
    .A(_06526_),
    .Y(_06532_),
    .D(_06531_));
 sg13g2_mux2_1 _23145_ (.A0(\top_ihp.oisc.regs[6][21] ),
    .A1(\top_ihp.oisc.regs[2][21] ),
    .S(net541),
    .X(_06533_));
 sg13g2_a22oi_1 _23146_ (.Y(_06534_),
    .B1(_06533_),
    .B2(_05748_),
    .A2(net536),
    .A1(\top_ihp.oisc.regs[8][21] ));
 sg13g2_a22oi_1 _23147_ (.Y(_06535_),
    .B1(net165),
    .B2(\top_ihp.oisc.regs[5][21] ),
    .A2(net335),
    .A1(\top_ihp.oisc.regs[19][21] ));
 sg13g2_a22oi_1 _23148_ (.Y(_06536_),
    .B1(net172),
    .B2(\top_ihp.oisc.regs[17][21] ),
    .A2(net533),
    .A1(\top_ihp.oisc.regs[22][21] ));
 sg13g2_a22oi_1 _23149_ (.Y(_06537_),
    .B1(net371),
    .B2(\top_ihp.oisc.regs[16][21] ),
    .A2(net170),
    .A1(\top_ihp.oisc.regs[3][21] ));
 sg13g2_nand4_1 _23150_ (.B(_06535_),
    .C(_06536_),
    .A(_06534_),
    .Y(_06538_),
    .D(_06537_));
 sg13g2_mux2_1 _23151_ (.A0(\top_ihp.oisc.regs[26][21] ),
    .A1(\top_ihp.oisc.regs[24][21] ),
    .S(net545),
    .X(_06539_));
 sg13g2_a22oi_1 _23152_ (.Y(_06540_),
    .B1(_06539_),
    .B2(net727),
    .A2(_05545_),
    .A1(\top_ihp.oisc.regs[18][21] ));
 sg13g2_and2_1 _23153_ (.A(\top_ihp.oisc.regs[10][21] ),
    .B(net537),
    .X(_06541_));
 sg13g2_a221oi_1 _23154_ (.B2(\top_ihp.oisc.regs[12][21] ),
    .C1(_06541_),
    .B1(net184),
    .A1(\top_ihp.oisc.regs[14][21] ),
    .Y(_06542_),
    .A2(net430));
 sg13g2_o21ai_1 _23155_ (.B1(_06542_),
    .Y(_06543_),
    .A1(net748),
    .A2(_06540_));
 sg13g2_nand2_1 _23156_ (.Y(_06544_),
    .A(\top_ihp.oisc.regs[15][21] ),
    .B(_05896_));
 sg13g2_a22oi_1 _23157_ (.Y(_06545_),
    .B1(net182),
    .B2(\top_ihp.oisc.regs[29][21] ),
    .A2(net342),
    .A1(\top_ihp.oisc.regs[7][21] ));
 sg13g2_a22oi_1 _23158_ (.Y(_06546_),
    .B1(net380),
    .B2(\top_ihp.oisc.regs[11][21] ),
    .A2(net540),
    .A1(\top_ihp.oisc.regs[20][21] ));
 sg13g2_a22oi_1 _23159_ (.Y(_06547_),
    .B1(net370),
    .B2(\top_ihp.oisc.regs[13][21] ),
    .A2(net664),
    .A1(\top_ihp.oisc.regs[28][21] ));
 sg13g2_a22oi_1 _23160_ (.Y(_06548_),
    .B1(_05883_),
    .B2(\top_ihp.oisc.regs[9][21] ),
    .A2(net432),
    .A1(\top_ihp.oisc.regs[4][21] ));
 sg13g2_a22oi_1 _23161_ (.Y(_06549_),
    .B1(net547),
    .B2(\top_ihp.oisc.regs[1][21] ),
    .A2(net551),
    .A1(\top_ihp.oisc.regs[25][21] ));
 sg13g2_and4_1 _23162_ (.A(_06546_),
    .B(_06547_),
    .C(_06548_),
    .D(_06549_),
    .X(_06550_));
 sg13g2_nand3_1 _23163_ (.B(_06545_),
    .C(_06550_),
    .A(_06544_),
    .Y(_06551_));
 sg13g2_nor4_1 _23164_ (.A(_06532_),
    .B(_06538_),
    .C(_06543_),
    .D(_06551_),
    .Y(_06552_));
 sg13g2_a22oi_1 _23165_ (.Y(_00401_),
    .B1(_06525_),
    .B2(_06552_),
    .A2(_06506_),
    .A1(_06505_));
 sg13g2_nand2_1 _23166_ (.Y(_06553_),
    .A(\top_ihp.oisc.regs[39][22] ),
    .B(net354));
 sg13g2_a22oi_1 _23167_ (.Y(_06554_),
    .B1(net406),
    .B2(\top_ihp.oisc.regs[46][22] ),
    .A2(net352),
    .A1(\top_ihp.oisc.regs[43][22] ));
 sg13g2_a22oi_1 _23168_ (.Y(_06555_),
    .B1(net187),
    .B2(\top_ihp.oisc.regs[56][22] ),
    .A2(_05595_),
    .A1(\top_ihp.oisc.regs[37][22] ));
 sg13g2_a22oi_1 _23169_ (.Y(_06556_),
    .B1(net353),
    .B2(\top_ihp.oisc.regs[35][22] ),
    .A2(net174),
    .A1(\top_ihp.oisc.regs[62][22] ));
 sg13g2_nand4_1 _23170_ (.B(_06554_),
    .C(_06555_),
    .A(_06553_),
    .Y(_06557_),
    .D(_06556_));
 sg13g2_and2_1 _23171_ (.A(\top_ihp.oisc.regs[6][22] ),
    .B(net667),
    .X(_06558_));
 sg13g2_a221oi_1 _23172_ (.B2(\top_ihp.oisc.regs[59][22] ),
    .C1(_06558_),
    .B1(_05683_),
    .A1(\top_ihp.oisc.regs[9][22] ),
    .Y(_06559_),
    .A2(net374));
 sg13g2_a22oi_1 _23173_ (.Y(_06560_),
    .B1(net387),
    .B2(\top_ihp.oisc.regs[47][22] ),
    .A2(net200),
    .A1(\top_ihp.oisc.regs[61][22] ));
 sg13g2_a22oi_1 _23174_ (.Y(_06561_),
    .B1(net391),
    .B2(\top_ihp.oisc.regs[33][22] ),
    .A2(net389),
    .A1(\top_ihp.oisc.regs[31][22] ));
 sg13g2_a22oi_1 _23175_ (.Y(_06562_),
    .B1(net539),
    .B2(\top_ihp.oisc.regs[34][22] ),
    .A2(net411),
    .A1(\top_ihp.oisc.regs[45][22] ));
 sg13g2_nand4_1 _23176_ (.B(_06560_),
    .C(_06561_),
    .A(_06559_),
    .Y(_06563_),
    .D(_06562_));
 sg13g2_a22oi_1 _23177_ (.Y(_06564_),
    .B1(_06046_),
    .B2(\top_ihp.oisc.regs[5][22] ),
    .A2(_05892_),
    .A1(\top_ihp.oisc.regs[16][22] ));
 sg13g2_a22oi_1 _23178_ (.Y(_06565_),
    .B1(_05574_),
    .B2(\top_ihp.oisc.regs[17][22] ),
    .A2(_05530_),
    .A1(\top_ihp.oisc.regs[29][22] ));
 sg13g2_a22oi_1 _23179_ (.Y(_06566_),
    .B1(_05898_),
    .B2(\top_ihp.oisc.regs[13][22] ),
    .A2(_05551_),
    .A1(\top_ihp.oisc.regs[19][22] ));
 sg13g2_a22oi_1 _23180_ (.Y(_06567_),
    .B1(net380),
    .B2(\top_ihp.oisc.regs[11][22] ),
    .A2(net554),
    .A1(\top_ihp.oisc.regs[7][22] ));
 sg13g2_nand4_1 _23181_ (.B(_06565_),
    .C(_06566_),
    .A(_06564_),
    .Y(_06568_),
    .D(_06567_));
 sg13g2_nand2b_1 _23182_ (.Y(_06569_),
    .B(net57),
    .A_N(_06568_));
 sg13g2_a22oi_1 _23183_ (.Y(_06570_),
    .B1(net195),
    .B2(\top_ihp.oisc.regs[58][22] ),
    .A2(net423),
    .A1(\top_ihp.oisc.regs[27][22] ));
 sg13g2_a22oi_1 _23184_ (.Y(_06571_),
    .B1(net398),
    .B2(\top_ihp.oisc.regs[55][22] ),
    .A2(net384),
    .A1(\top_ihp.oisc.regs[38][22] ));
 sg13g2_a22oi_1 _23185_ (.Y(_06572_),
    .B1(net388),
    .B2(\top_ihp.oisc.regs[30][22] ),
    .A2(net385),
    .A1(\top_ihp.oisc.regs[40][22] ));
 sg13g2_a22oi_1 _23186_ (.Y(_06573_),
    .B1(net196),
    .B2(\top_ihp.oisc.regs[54][22] ),
    .A2(net344),
    .A1(\top_ihp.oisc.regs[53][22] ));
 sg13g2_nand4_1 _23187_ (.B(_06571_),
    .C(_06572_),
    .A(_06570_),
    .Y(_06574_),
    .D(_06573_));
 sg13g2_nor4_1 _23188_ (.A(_06557_),
    .B(_06563_),
    .C(_06569_),
    .D(_06574_),
    .Y(_06575_));
 sg13g2_nor2_1 _23189_ (.A(_08180_),
    .B(net804),
    .Y(_06576_));
 sg13g2_a221oi_1 _23190_ (.B2(\top_ihp.oisc.regs[2][22] ),
    .C1(_06576_),
    .B1(net369),
    .A1(\top_ihp.oisc.regs[41][22] ),
    .Y(_06577_),
    .A2(_05710_));
 sg13g2_a22oi_1 _23191_ (.Y(_06578_),
    .B1(net419),
    .B2(\top_ihp.oisc.regs[44][22] ),
    .A2(net416),
    .A1(\top_ihp.oisc.regs[42][22] ));
 sg13g2_a22oi_1 _23192_ (.Y(_06579_),
    .B1(net404),
    .B2(\top_ihp.oisc.regs[49][22] ),
    .A2(net409),
    .A1(\top_ihp.oisc.regs[48][22] ));
 sg13g2_a22oi_1 _23193_ (.Y(_06580_),
    .B1(_06297_),
    .B2(\top_ihp.oisc.regs[25][22] ),
    .A2(_05640_),
    .A1(\top_ihp.oisc.regs[57][22] ));
 sg13g2_nand4_1 _23194_ (.B(_06578_),
    .C(_06579_),
    .A(_06577_),
    .Y(_06581_),
    .D(_06580_));
 sg13g2_a22oi_1 _23195_ (.Y(_06582_),
    .B1(net392),
    .B2(\top_ihp.oisc.regs[52][22] ),
    .A2(net420),
    .A1(\top_ihp.oisc.regs[51][22] ));
 sg13g2_a22oi_1 _23196_ (.Y(_06583_),
    .B1(_05847_),
    .B2(\top_ihp.oisc.regs[60][22] ),
    .A2(net188),
    .A1(\top_ihp.oisc.regs[50][22] ));
 sg13g2_a22oi_1 _23197_ (.Y(_06584_),
    .B1(net338),
    .B2(\top_ihp.oisc.regs[32][22] ),
    .A2(net413),
    .A1(\top_ihp.oisc.regs[63][22] ));
 sg13g2_a22oi_1 _23198_ (.Y(_06585_),
    .B1(_05667_),
    .B2(\top_ihp.oisc.regs[18][22] ),
    .A2(net729),
    .A1(\top_ihp.oisc.regs[20][22] ));
 sg13g2_nor2_1 _23199_ (.A(_06462_),
    .B(_06585_),
    .Y(_06586_));
 sg13g2_a21oi_1 _23200_ (.A1(\top_ihp.oisc.regs[36][22] ),
    .A2(net436),
    .Y(_06587_),
    .B1(_06586_));
 sg13g2_nand4_1 _23201_ (.B(_06583_),
    .C(_06584_),
    .A(_06582_),
    .Y(_06588_),
    .D(_06587_));
 sg13g2_nor2_1 _23202_ (.A(_04093_),
    .B(_05822_),
    .Y(_06589_));
 sg13g2_mux2_1 _23203_ (.A0(\top_ihp.oisc.regs[23][22] ),
    .A1(\top_ihp.oisc.regs[21][22] ),
    .S(net545),
    .X(_06590_));
 sg13g2_a22oi_1 _23204_ (.Y(_06591_),
    .B1(_06589_),
    .B2(_06590_),
    .A2(net167),
    .A1(\top_ihp.oisc.regs[24][22] ));
 sg13g2_a22oi_1 _23205_ (.Y(_06592_),
    .B1(net166),
    .B2(\top_ihp.oisc.regs[3][22] ),
    .A2(net535),
    .A1(\top_ihp.oisc.regs[28][22] ));
 sg13g2_mux2_1 _23206_ (.A0(\top_ihp.oisc.regs[10][22] ),
    .A1(\top_ihp.oisc.regs[8][22] ),
    .S(net669),
    .X(_06593_));
 sg13g2_a22oi_1 _23207_ (.Y(_06594_),
    .B1(_06119_),
    .B2(_06593_),
    .A2(net162),
    .A1(\top_ihp.oisc.regs[15][22] ));
 sg13g2_a22oi_1 _23208_ (.Y(_06595_),
    .B1(net431),
    .B2(\top_ihp.oisc.regs[1][22] ),
    .A2(net163),
    .A1(\top_ihp.oisc.regs[4][22] ));
 sg13g2_nand4_1 _23209_ (.B(_06592_),
    .C(_06594_),
    .A(_06591_),
    .Y(_06596_),
    .D(_06595_));
 sg13g2_nand2_1 _23210_ (.Y(_06597_),
    .A(\top_ihp.oisc.regs[22][22] ),
    .B(_05440_));
 sg13g2_mux2_1 _23211_ (.A0(\top_ihp.oisc.regs[14][22] ),
    .A1(\top_ihp.oisc.regs[12][22] ),
    .S(net545),
    .X(_06598_));
 sg13g2_a22oi_1 _23212_ (.Y(_06599_),
    .B1(_06484_),
    .B2(_06598_),
    .A2(net168),
    .A1(\top_ihp.oisc.regs[26][22] ));
 sg13g2_nand2_1 _23213_ (.Y(_06600_),
    .A(_06597_),
    .B(_06599_));
 sg13g2_nor4_1 _23214_ (.A(_06581_),
    .B(_06588_),
    .C(_06596_),
    .D(_06600_),
    .Y(_06601_));
 sg13g2_a21oi_1 _23215_ (.A1(_00226_),
    .A2(_05707_),
    .Y(_06602_),
    .B1(net58));
 sg13g2_nor2_1 _23216_ (.A(_06576_),
    .B(_06602_),
    .Y(_06603_));
 sg13g2_a21oi_1 _23217_ (.A1(_06575_),
    .A2(_06601_),
    .Y(_00402_),
    .B1(_06603_));
 sg13g2_a22oi_1 _23218_ (.Y(_06604_),
    .B1(net191),
    .B2(\top_ihp.oisc.regs[59][23] ),
    .A2(_05654_),
    .A1(\top_ihp.oisc.regs[56][23] ));
 sg13g2_a22oi_1 _23219_ (.Y(_06605_),
    .B1(_05677_),
    .B2(\top_ihp.oisc.regs[50][23] ),
    .A2(net352),
    .A1(\top_ihp.oisc.regs[43][23] ));
 sg13g2_a22oi_1 _23220_ (.Y(_06606_),
    .B1(net364),
    .B2(\top_ihp.oisc.regs[52][23] ),
    .A2(_05721_),
    .A1(\top_ihp.oisc.regs[33][23] ));
 sg13g2_a22oi_1 _23221_ (.Y(_06607_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[32][23] ),
    .A2(net389),
    .A1(\top_ihp.oisc.regs[31][23] ));
 sg13g2_nand4_1 _23222_ (.B(_06605_),
    .C(_06606_),
    .A(_06604_),
    .Y(_06608_),
    .D(_06607_));
 sg13g2_a22oi_1 _23223_ (.Y(_06609_),
    .B1(_05775_),
    .B2(\top_ihp.oisc.regs[24][23] ),
    .A2(net552),
    .A1(\top_ihp.oisc.regs[20][23] ));
 sg13g2_a22oi_1 _23224_ (.Y(_06610_),
    .B1(_05573_),
    .B2(\top_ihp.oisc.regs[17][23] ),
    .A2(_05570_),
    .A1(\top_ihp.oisc.regs[15][23] ));
 sg13g2_mux2_1 _23225_ (.A0(\top_ihp.oisc.regs[12][23] ),
    .A1(\top_ihp.oisc.regs[8][23] ),
    .S(net670),
    .X(_06611_));
 sg13g2_nor2_1 _23226_ (.A(net672),
    .B(net774),
    .Y(_06612_));
 sg13g2_a22oi_1 _23227_ (.Y(_06613_),
    .B1(_06611_),
    .B2(_06612_),
    .A2(_05765_),
    .A1(\top_ihp.oisc.regs[26][23] ));
 sg13g2_a22oi_1 _23228_ (.Y(_06614_),
    .B1(_05513_),
    .B2(\top_ihp.oisc.regs[14][23] ),
    .A2(_05439_),
    .A1(\top_ihp.oisc.regs[22][23] ));
 sg13g2_and4_1 _23229_ (.A(_06609_),
    .B(_06610_),
    .C(_06613_),
    .D(_06614_),
    .X(_06615_));
 sg13g2_nand3_1 _23230_ (.B(_05469_),
    .C(net673),
    .A(\top_ihp.oisc.regs[58][23] ),
    .Y(_06616_));
 sg13g2_nand3_1 _23231_ (.B(_06094_),
    .C(net728),
    .A(\top_ihp.oisc.regs[34][23] ),
    .Y(_06617_));
 sg13g2_a21o_1 _23232_ (.A2(_06617_),
    .A1(_06616_),
    .B1(_05554_),
    .X(_06618_));
 sg13g2_a22oi_1 _23233_ (.Y(_06619_),
    .B1(net345),
    .B2(\top_ihp.oisc.regs[5][23] ),
    .A2(_05903_),
    .A1(\top_ihp.oisc.regs[25][23] ));
 sg13g2_a22oi_1 _23234_ (.Y(_06620_),
    .B1(net164),
    .B2(\top_ihp.oisc.regs[9][23] ),
    .A2(net170),
    .A1(\top_ihp.oisc.regs[3][23] ));
 sg13g2_nand4_1 _23235_ (.B(_06618_),
    .C(_06619_),
    .A(_06615_),
    .Y(_06621_),
    .D(_06620_));
 sg13g2_nand3_1 _23236_ (.B(_05667_),
    .C(net747),
    .A(\top_ihp.oisc.regs[10][23] ),
    .Y(_06622_));
 sg13g2_nand3_1 _23237_ (.B(net721),
    .C(net749),
    .A(\top_ihp.oisc.regs[6][23] ),
    .Y(_06623_));
 sg13g2_nand2_1 _23238_ (.Y(_06624_),
    .A(_06622_),
    .B(_06623_));
 sg13g2_a221oi_1 _23239_ (.B2(\top_ihp.oisc.regs[21][23] ),
    .C1(_06624_),
    .B1(net666),
    .A1(\top_ihp.oisc.regs[35][23] ),
    .Y(_06625_),
    .A2(net353));
 sg13g2_nand2_1 _23240_ (.Y(_06626_),
    .A(\top_ihp.oisc.regs[11][23] ),
    .B(net169));
 sg13g2_a22oi_1 _23241_ (.Y(_06627_),
    .B1(_05825_),
    .B2(\top_ihp.oisc.regs[23][23] ),
    .A2(net783),
    .A1(net1061));
 sg13g2_a22oi_1 _23242_ (.Y(_06628_),
    .B1(net350),
    .B2(\top_ihp.oisc.regs[19][23] ),
    .A2(net438),
    .A1(\top_ihp.oisc.regs[7][23] ));
 sg13g2_nand4_1 _23243_ (.B(_06626_),
    .C(_06627_),
    .A(_06625_),
    .Y(_06629_),
    .D(_06628_));
 sg13g2_a22oi_1 _23244_ (.Y(_06630_),
    .B1(net179),
    .B2(\top_ihp.oisc.regs[2][23] ),
    .A2(net180),
    .A1(\top_ihp.oisc.regs[13][23] ));
 sg13g2_a22oi_1 _23245_ (.Y(_06631_),
    .B1(net183),
    .B2(\top_ihp.oisc.regs[16][23] ),
    .A2(net182),
    .A1(\top_ihp.oisc.regs[29][23] ));
 sg13g2_a22oi_1 _23246_ (.Y(_06632_),
    .B1(net535),
    .B2(\top_ihp.oisc.regs[28][23] ),
    .A2(_05887_),
    .A1(\top_ihp.oisc.regs[1][23] ));
 sg13g2_a22oi_1 _23247_ (.Y(_06633_),
    .B1(net343),
    .B2(\top_ihp.oisc.regs[18][23] ),
    .A2(net204),
    .A1(\top_ihp.oisc.regs[4][23] ));
 sg13g2_nand4_1 _23248_ (.B(_06631_),
    .C(_06632_),
    .A(_06630_),
    .Y(_06634_),
    .D(_06633_));
 sg13g2_nor4_1 _23249_ (.A(_06608_),
    .B(_06621_),
    .C(_06629_),
    .D(_06634_),
    .Y(_06635_));
 sg13g2_nand2_1 _23250_ (.Y(_06636_),
    .A(_05488_),
    .B(_05518_));
 sg13g2_nor3_2 _23251_ (.A(_06636_),
    .B(_06094_),
    .C(_05612_),
    .Y(_06637_));
 sg13g2_a22oi_1 _23252_ (.Y(_06638_),
    .B1(_06637_),
    .B2(\top_ihp.oisc.regs[44][23] ),
    .A2(net404),
    .A1(\top_ihp.oisc.regs[49][23] ));
 sg13g2_a22oi_1 _23253_ (.Y(_06639_),
    .B1(net379),
    .B2(\top_ihp.oisc.regs[45][23] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[36][23] ));
 sg13g2_a22oi_1 _23254_ (.Y(_06640_),
    .B1(_05949_),
    .B2(\top_ihp.oisc.regs[55][23] ),
    .A2(net341),
    .A1(\top_ihp.oisc.regs[27][23] ));
 sg13g2_a22oi_1 _23255_ (.Y(_06641_),
    .B1(_05626_),
    .B2(\top_ihp.oisc.regs[51][23] ),
    .A2(net377),
    .A1(\top_ihp.oisc.regs[53][23] ));
 sg13g2_nand4_1 _23256_ (.B(_06639_),
    .C(_06640_),
    .A(_06638_),
    .Y(_06642_),
    .D(_06641_));
 sg13g2_a22oi_1 _23257_ (.Y(_06643_),
    .B1(net176),
    .B2(\top_ihp.oisc.regs[62][23] ),
    .A2(net385),
    .A1(\top_ihp.oisc.regs[40][23] ));
 sg13g2_a22oi_1 _23258_ (.Y(_06644_),
    .B1(_06029_),
    .B2(\top_ihp.oisc.regs[60][23] ),
    .A2(_06042_),
    .A1(\top_ihp.oisc.regs[30][23] ));
 sg13g2_a22oi_1 _23259_ (.Y(_06645_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[39][23] ),
    .A2(net358),
    .A1(\top_ihp.oisc.regs[47][23] ));
 sg13g2_a22oi_1 _23260_ (.Y(_06646_),
    .B1(net175),
    .B2(\top_ihp.oisc.regs[61][23] ),
    .A2(_05809_),
    .A1(\top_ihp.oisc.regs[42][23] ));
 sg13g2_nand4_1 _23261_ (.B(_06644_),
    .C(_06645_),
    .A(_06643_),
    .Y(_06647_),
    .D(_06646_));
 sg13g2_a22oi_1 _23262_ (.Y(_06648_),
    .B1(net426),
    .B2(\top_ihp.oisc.regs[37][23] ),
    .A2(_05927_),
    .A1(\top_ihp.oisc.regs[63][23] ));
 sg13g2_a22oi_1 _23263_ (.Y(_06649_),
    .B1(net197),
    .B2(\top_ihp.oisc.regs[48][23] ),
    .A2(net348),
    .A1(\top_ihp.oisc.regs[57][23] ));
 sg13g2_a22oi_1 _23264_ (.Y(_06650_),
    .B1(net384),
    .B2(\top_ihp.oisc.regs[38][23] ),
    .A2(net178),
    .A1(\top_ihp.oisc.regs[54][23] ));
 sg13g2_a22oi_1 _23265_ (.Y(_06651_),
    .B1(net349),
    .B2(\top_ihp.oisc.regs[46][23] ),
    .A2(_06086_),
    .A1(\top_ihp.oisc.regs[41][23] ));
 sg13g2_nand4_1 _23266_ (.B(_06649_),
    .C(_06650_),
    .A(_06648_),
    .Y(_06652_),
    .D(_06651_));
 sg13g2_nor4_2 _23267_ (.A(_05944_),
    .B(_06642_),
    .C(_06647_),
    .Y(_06653_),
    .D(_06652_));
 sg13g2_nand2_1 _23268_ (.Y(_06654_),
    .A(_00227_),
    .B(net60));
 sg13g2_a22oi_1 _23269_ (.Y(_06655_),
    .B1(net26),
    .B2(_06654_),
    .A2(net746),
    .A1(_08163_));
 sg13g2_a21oi_1 _23270_ (.A1(_06635_),
    .A2(_06653_),
    .Y(_00403_),
    .B1(_06655_));
 sg13g2_a22oi_1 _23271_ (.Y(_06656_),
    .B1(_05848_),
    .B2(\top_ihp.oisc.regs[60][24] ),
    .A2(_06080_),
    .A1(\top_ihp.oisc.regs[27][24] ));
 sg13g2_a22oi_1 _23272_ (.Y(_06657_),
    .B1(net404),
    .B2(\top_ihp.oisc.regs[49][24] ),
    .A2(net419),
    .A1(\top_ihp.oisc.regs[44][24] ));
 sg13g2_a22oi_1 _23273_ (.Y(_06658_),
    .B1(net397),
    .B2(\top_ihp.oisc.regs[37][24] ),
    .A2(net351),
    .A1(\top_ihp.oisc.regs[40][24] ));
 sg13g2_a22oi_1 _23274_ (.Y(_06659_),
    .B1(net379),
    .B2(\top_ihp.oisc.regs[45][24] ),
    .A2(_05665_),
    .A1(\top_ihp.oisc.regs[63][24] ));
 sg13g2_nand4_1 _23275_ (.B(_06657_),
    .C(_06658_),
    .A(_06656_),
    .Y(_06660_),
    .D(_06659_));
 sg13g2_a22oi_1 _23276_ (.Y(_06661_),
    .B1(_05924_),
    .B2(\top_ihp.oisc.regs[58][24] ),
    .A2(net178),
    .A1(\top_ihp.oisc.regs[54][24] ));
 sg13g2_a22oi_1 _23277_ (.Y(_06662_),
    .B1(_05726_),
    .B2(\top_ihp.oisc.regs[46][24] ),
    .A2(_05981_),
    .A1(\top_ihp.oisc.regs[43][24] ));
 sg13g2_a22oi_1 _23278_ (.Y(_06663_),
    .B1(net420),
    .B2(\top_ihp.oisc.regs[51][24] ),
    .A2(net333),
    .A1(\top_ihp.oisc.regs[57][24] ));
 sg13g2_a22oi_1 _23279_ (.Y(_06664_),
    .B1(_05701_),
    .B2(\top_ihp.oisc.regs[8][24] ),
    .A2(net721),
    .A1(\top_ihp.oisc.regs[14][24] ));
 sg13g2_nor2_1 _23280_ (.A(net774),
    .B(_06664_),
    .Y(_06665_));
 sg13g2_a21oi_1 _23281_ (.A1(\top_ihp.oisc.regs[31][24] ),
    .A2(net389),
    .Y(_06666_),
    .B1(_06665_));
 sg13g2_nand4_1 _23282_ (.B(_06662_),
    .C(_06663_),
    .A(_06661_),
    .Y(_06667_),
    .D(_06666_));
 sg13g2_a22oi_1 _23283_ (.Y(_06668_),
    .B1(_06106_),
    .B2(\top_ihp.oisc.regs[3][24] ),
    .A2(_06001_),
    .A1(\top_ihp.oisc.regs[28][24] ));
 sg13g2_a22oi_1 _23284_ (.Y(_06669_),
    .B1(net168),
    .B2(\top_ihp.oisc.regs[26][24] ),
    .A2(_05473_),
    .A1(\top_ihp.oisc.regs[20][24] ));
 sg13g2_a22oi_1 _23285_ (.Y(_06670_),
    .B1(net173),
    .B2(\top_ihp.oisc.regs[11][24] ),
    .A2(_05828_),
    .A1(\top_ihp.oisc.regs[13][24] ));
 sg13g2_a22oi_1 _23286_ (.Y(_06671_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[25][24] ),
    .A2(net533),
    .A1(\top_ihp.oisc.regs[22][24] ));
 sg13g2_nand4_1 _23287_ (.B(_06669_),
    .C(_06670_),
    .A(_06668_),
    .Y(_06672_),
    .D(_06671_));
 sg13g2_mux2_1 _23288_ (.A0(\top_ihp.oisc.regs[6][24] ),
    .A1(\top_ihp.oisc.regs[2][24] ),
    .S(_05770_),
    .X(_06673_));
 sg13g2_a22oi_1 _23289_ (.Y(_06674_),
    .B1(_05748_),
    .B2(_06673_),
    .A2(net182),
    .A1(\top_ihp.oisc.regs[29][24] ));
 sg13g2_a22oi_1 _23290_ (.Y(_06675_),
    .B1(_05893_),
    .B2(\top_ihp.oisc.regs[16][24] ),
    .A2(_06065_),
    .A1(\top_ihp.oisc.regs[7][24] ));
 sg13g2_a22oi_1 _23291_ (.Y(_06676_),
    .B1(net666),
    .B2(\top_ihp.oisc.regs[21][24] ),
    .A2(net803),
    .A1(_08154_));
 sg13g2_inv_1 _23292_ (.Y(_06677_),
    .A(_06676_));
 sg13g2_a221oi_1 _23293_ (.B2(\top_ihp.oisc.regs[38][24] ),
    .C1(_06677_),
    .B1(net378),
    .A1(\top_ihp.oisc.regs[17][24] ),
    .Y(_06678_),
    .A2(net427));
 sg13g2_nand3_1 _23294_ (.B(_06675_),
    .C(_06678_),
    .A(_06674_),
    .Y(_06679_));
 sg13g2_nor4_1 _23295_ (.A(_06660_),
    .B(_06667_),
    .C(_06672_),
    .D(_06679_),
    .Y(_06680_));
 sg13g2_a22oi_1 _23296_ (.Y(_06681_),
    .B1(_05605_),
    .B2(\top_ihp.oisc.regs[39][24] ),
    .A2(_05683_),
    .A1(\top_ihp.oisc.regs[59][24] ));
 sg13g2_a22oi_1 _23297_ (.Y(_06682_),
    .B1(net542),
    .B2(\top_ihp.oisc.regs[34][24] ),
    .A2(_05614_),
    .A1(\top_ihp.oisc.regs[32][24] ));
 sg13g2_and2_1 _23298_ (.A(_06681_),
    .B(_06682_),
    .X(_06683_));
 sg13g2_a22oi_1 _23299_ (.Y(_06684_),
    .B1(_05761_),
    .B2(\top_ihp.oisc.regs[5][24] ),
    .A2(_05538_),
    .A1(\top_ihp.oisc.regs[24][24] ));
 sg13g2_a22oi_1 _23300_ (.Y(_06685_),
    .B1(_05548_),
    .B2(\top_ihp.oisc.regs[18][24] ),
    .A2(_05499_),
    .A1(\top_ihp.oisc.regs[4][24] ));
 sg13g2_and2_1 _23301_ (.A(_06684_),
    .B(_06685_),
    .X(_06686_));
 sg13g2_a22oi_1 _23302_ (.Y(_06687_),
    .B1(net372),
    .B2(\top_ihp.oisc.regs[12][24] ),
    .A2(net431),
    .A1(\top_ihp.oisc.regs[1][24] ));
 sg13g2_nand3_1 _23303_ (.B(net750),
    .C(_05489_),
    .A(\top_ihp.oisc.regs[23][24] ),
    .Y(_06688_));
 sg13g2_nand3_1 _23304_ (.B(net548),
    .C(_06175_),
    .A(\top_ihp.oisc.regs[10][24] ),
    .Y(_06689_));
 sg13g2_nand2_1 _23305_ (.Y(_06690_),
    .A(_06688_),
    .B(_06689_));
 sg13g2_a22oi_1 _23306_ (.Y(_06691_),
    .B1(_06690_),
    .B2(net550),
    .A2(_06271_),
    .A1(\top_ihp.oisc.regs[19][24] ));
 sg13g2_nand4_1 _23307_ (.B(_06686_),
    .C(_06687_),
    .A(_06683_),
    .Y(_06692_),
    .D(_06691_));
 sg13g2_a22oi_1 _23308_ (.Y(_06693_),
    .B1(net405),
    .B2(\top_ihp.oisc.regs[52][24] ),
    .A2(net388),
    .A1(\top_ihp.oisc.regs[30][24] ));
 sg13g2_a22oi_1 _23309_ (.Y(_06694_),
    .B1(net360),
    .B2(\top_ihp.oisc.regs[33][24] ),
    .A2(_05812_),
    .A1(\top_ihp.oisc.regs[62][24] ));
 sg13g2_a22oi_1 _23310_ (.Y(_06695_),
    .B1(net403),
    .B2(\top_ihp.oisc.regs[55][24] ),
    .A2(net188),
    .A1(\top_ihp.oisc.regs[50][24] ));
 sg13g2_a22oi_1 _23311_ (.Y(_06696_),
    .B1(_05855_),
    .B2(\top_ihp.oisc.regs[48][24] ),
    .A2(net377),
    .A1(\top_ihp.oisc.regs[53][24] ));
 sg13g2_nand4_1 _23312_ (.B(_06694_),
    .C(_06695_),
    .A(_06693_),
    .Y(_06697_),
    .D(_06696_));
 sg13g2_a22oi_1 _23313_ (.Y(_06698_),
    .B1(net395),
    .B2(\top_ihp.oisc.regs[41][24] ),
    .A2(_05954_),
    .A1(\top_ihp.oisc.regs[36][24] ));
 sg13g2_a22oi_1 _23314_ (.Y(_06699_),
    .B1(net193),
    .B2(\top_ihp.oisc.regs[56][24] ),
    .A2(_06172_),
    .A1(\top_ihp.oisc.regs[42][24] ));
 sg13g2_and2_1 _23315_ (.A(\top_ihp.oisc.regs[35][24] ),
    .B(_05718_),
    .X(_06700_));
 sg13g2_a221oi_1 _23316_ (.B2(\top_ihp.oisc.regs[15][24] ),
    .C1(_06700_),
    .B1(net428),
    .A1(\top_ihp.oisc.regs[9][24] ),
    .Y(_06701_),
    .A2(net374));
 sg13g2_a22oi_1 _23317_ (.Y(_06702_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[47][24] ),
    .A2(net175),
    .A1(\top_ihp.oisc.regs[61][24] ));
 sg13g2_nand4_1 _23318_ (.B(_06699_),
    .C(_06701_),
    .A(_06698_),
    .Y(_06703_),
    .D(_06702_));
 sg13g2_nor4_1 _23319_ (.A(net60),
    .B(_06692_),
    .C(_06697_),
    .D(_06703_),
    .Y(_06704_));
 sg13g2_nand2_1 _23320_ (.Y(_06705_),
    .A(_00228_),
    .B(net60));
 sg13g2_a22oi_1 _23321_ (.Y(_06706_),
    .B1(_05943_),
    .B2(_06705_),
    .A2(_06304_),
    .A1(_08154_));
 sg13g2_a21oi_1 _23322_ (.A1(_06680_),
    .A2(_06704_),
    .Y(_00404_),
    .B1(_06706_));
 sg13g2_a22oi_1 _23323_ (.Y(_06707_),
    .B1(net426),
    .B2(\top_ihp.oisc.regs[37][25] ),
    .A2(net198),
    .A1(\top_ihp.oisc.regs[59][25] ));
 sg13g2_a22oi_1 _23324_ (.Y(_06708_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[32][25] ),
    .A2(net351),
    .A1(\top_ihp.oisc.regs[40][25] ));
 sg13g2_a22oi_1 _23325_ (.Y(_06709_),
    .B1(net340),
    .B2(\top_ihp.oisc.regs[41][25] ),
    .A2(net341),
    .A1(\top_ihp.oisc.regs[27][25] ));
 sg13g2_a22oi_1 _23326_ (.Y(_06710_),
    .B1(net399),
    .B2(\top_ihp.oisc.regs[58][25] ),
    .A2(net542),
    .A1(\top_ihp.oisc.regs[34][25] ));
 sg13g2_nand4_1 _23327_ (.B(_06708_),
    .C(_06709_),
    .A(_06707_),
    .Y(_06711_),
    .D(_06710_));
 sg13g2_a22oi_1 _23328_ (.Y(_06712_),
    .B1(net167),
    .B2(\top_ihp.oisc.regs[24][25] ),
    .A2(net367),
    .A1(\top_ihp.oisc.regs[26][25] ));
 sg13g2_a22oi_1 _23329_ (.Y(_06713_),
    .B1(net180),
    .B2(\top_ihp.oisc.regs[13][25] ),
    .A2(net203),
    .A1(\top_ihp.oisc.regs[29][25] ));
 sg13g2_a22oi_1 _23330_ (.Y(_06714_),
    .B1(net535),
    .B2(\top_ihp.oisc.regs[28][25] ),
    .A2(net438),
    .A1(\top_ihp.oisc.regs[7][25] ));
 sg13g2_a22oi_1 _23331_ (.Y(_06715_),
    .B1(net534),
    .B2(\top_ihp.oisc.regs[18][25] ),
    .A2(net368),
    .A1(\top_ihp.oisc.regs[25][25] ));
 sg13g2_nand4_1 _23332_ (.B(_06713_),
    .C(_06714_),
    .A(_06712_),
    .Y(_06716_),
    .D(_06715_));
 sg13g2_a22oi_1 _23333_ (.Y(_06717_),
    .B1(net169),
    .B2(\top_ihp.oisc.regs[11][25] ),
    .A2(net434),
    .A1(\top_ihp.oisc.regs[20][25] ));
 sg13g2_a22oi_1 _23334_ (.Y(_06718_),
    .B1(net334),
    .B2(\top_ihp.oisc.regs[10][25] ),
    .A2(net164),
    .A1(\top_ihp.oisc.regs[9][25] ));
 sg13g2_a22oi_1 _23335_ (.Y(_06719_),
    .B1(net181),
    .B2(\top_ihp.oisc.regs[15][25] ),
    .A2(net163),
    .A1(\top_ihp.oisc.regs[4][25] ));
 sg13g2_a22oi_1 _23336_ (.Y(_06720_),
    .B1(net165),
    .B2(\top_ihp.oisc.regs[5][25] ),
    .A2(_05784_),
    .A1(\top_ihp.oisc.regs[6][25] ));
 sg13g2_nand4_1 _23337_ (.B(_06718_),
    .C(_06719_),
    .A(_06717_),
    .Y(_06721_),
    .D(_06720_));
 sg13g2_mux2_1 _23338_ (.A0(\top_ihp.oisc.regs[12][25] ),
    .A1(\top_ihp.oisc.regs[8][25] ),
    .S(net541),
    .X(_06722_));
 sg13g2_a22oi_1 _23339_ (.Y(_06723_),
    .B1(_06722_),
    .B2(net545),
    .A2(net721),
    .A1(\top_ihp.oisc.regs[14][25] ));
 sg13g2_a22oi_1 _23340_ (.Y(_06724_),
    .B1(net427),
    .B2(\top_ihp.oisc.regs[17][25] ),
    .A2(net401),
    .A1(\top_ihp.oisc.regs[3][25] ));
 sg13g2_a22oi_1 _23341_ (.Y(_06725_),
    .B1(_05824_),
    .B2(\top_ihp.oisc.regs[23][25] ),
    .A2(net835),
    .A1(_08157_));
 sg13g2_inv_1 _23342_ (.Y(_06726_),
    .A(_06725_));
 sg13g2_a221oi_1 _23343_ (.B2(\top_ihp.oisc.regs[21][25] ),
    .C1(_06726_),
    .B1(net663),
    .A1(\top_ihp.oisc.regs[22][25] ),
    .Y(_06727_),
    .A2(_05439_));
 sg13g2_a22oi_1 _23344_ (.Y(_06728_),
    .B1(net371),
    .B2(\top_ihp.oisc.regs[16][25] ),
    .A2(net547),
    .A1(\top_ihp.oisc.regs[1][25] ));
 sg13g2_a22oi_1 _23345_ (.Y(_06729_),
    .B1(_05750_),
    .B2(\top_ihp.oisc.regs[2][25] ),
    .A2(net543),
    .A1(\top_ihp.oisc.regs[19][25] ));
 sg13g2_and4_1 _23346_ (.A(_06724_),
    .B(_06727_),
    .C(_06728_),
    .D(_06729_),
    .X(_06730_));
 sg13g2_o21ai_1 _23347_ (.B1(_06730_),
    .Y(_06731_),
    .A1(net774),
    .A2(_06723_));
 sg13g2_nor4_1 _23348_ (.A(_06711_),
    .B(_06716_),
    .C(_06721_),
    .D(_06731_),
    .Y(_06732_));
 sg13g2_nand2_1 _23349_ (.Y(_06733_),
    .A(\top_ihp.oisc.regs[54][25] ),
    .B(net196));
 sg13g2_a22oi_1 _23350_ (.Y(_06734_),
    .B1(net364),
    .B2(\top_ihp.oisc.regs[52][25] ),
    .A2(net419),
    .A1(\top_ihp.oisc.regs[44][25] ));
 sg13g2_a22oi_1 _23351_ (.Y(_06735_),
    .B1(net352),
    .B2(\top_ihp.oisc.regs[43][25] ),
    .A2(net333),
    .A1(\top_ihp.oisc.regs[57][25] ));
 sg13g2_a22oi_1 _23352_ (.Y(_06736_),
    .B1(net409),
    .B2(\top_ihp.oisc.regs[48][25] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[36][25] ));
 sg13g2_nand4_1 _23353_ (.B(_06734_),
    .C(_06735_),
    .A(_06733_),
    .Y(_06737_),
    .D(_06736_));
 sg13g2_a22oi_1 _23354_ (.Y(_06738_),
    .B1(net360),
    .B2(\top_ihp.oisc.regs[33][25] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[53][25] ));
 sg13g2_a22oi_1 _23355_ (.Y(_06739_),
    .B1(net349),
    .B2(\top_ihp.oisc.regs[46][25] ),
    .A2(net358),
    .A1(\top_ihp.oisc.regs[47][25] ));
 sg13g2_nand3_1 _23356_ (.B(_06738_),
    .C(_06739_),
    .A(net61),
    .Y(_06740_));
 sg13g2_a22oi_1 _23357_ (.Y(_06741_),
    .B1(net394),
    .B2(\top_ihp.oisc.regs[45][25] ),
    .A2(net199),
    .A1(\top_ihp.oisc.regs[50][25] ));
 sg13g2_a22oi_1 _23358_ (.Y(_06742_),
    .B1(net384),
    .B2(\top_ihp.oisc.regs[38][25] ),
    .A2(net400),
    .A1(\top_ihp.oisc.regs[63][25] ));
 sg13g2_a22oi_1 _23359_ (.Y(_06743_),
    .B1(net408),
    .B2(\top_ihp.oisc.regs[35][25] ),
    .A2(net393),
    .A1(\top_ihp.oisc.regs[42][25] ));
 sg13g2_a22oi_1 _23360_ (.Y(_06744_),
    .B1(net187),
    .B2(\top_ihp.oisc.regs[56][25] ),
    .A2(net174),
    .A1(\top_ihp.oisc.regs[62][25] ));
 sg13g2_nand4_1 _23361_ (.B(_06742_),
    .C(_06743_),
    .A(_06741_),
    .Y(_06745_),
    .D(_06744_));
 sg13g2_a22oi_1 _23362_ (.Y(_06746_),
    .B1(net189),
    .B2(\top_ihp.oisc.regs[60][25] ),
    .A2(net354),
    .A1(\top_ihp.oisc.regs[39][25] ));
 sg13g2_a22oi_1 _23363_ (.Y(_06747_),
    .B1(net386),
    .B2(\top_ihp.oisc.regs[49][25] ),
    .A2(net376),
    .A1(\top_ihp.oisc.regs[51][25] ));
 sg13g2_a22oi_1 _23364_ (.Y(_06748_),
    .B1(net190),
    .B2(\top_ihp.oisc.regs[61][25] ),
    .A2(net388),
    .A1(\top_ihp.oisc.regs[30][25] ));
 sg13g2_a22oi_1 _23365_ (.Y(_06749_),
    .B1(net403),
    .B2(\top_ihp.oisc.regs[55][25] ),
    .A2(net435),
    .A1(\top_ihp.oisc.regs[31][25] ));
 sg13g2_nand4_1 _23366_ (.B(_06747_),
    .C(_06748_),
    .A(_06746_),
    .Y(_06750_),
    .D(_06749_));
 sg13g2_nor4_2 _23367_ (.A(_06737_),
    .B(_06740_),
    .C(_06745_),
    .Y(_06751_),
    .D(_06750_));
 sg13g2_nand2_1 _23368_ (.Y(_06752_),
    .A(_00229_),
    .B(net59));
 sg13g2_a22oi_1 _23369_ (.Y(_06753_),
    .B1(net26),
    .B2(_06752_),
    .A2(net746),
    .A1(_08157_));
 sg13g2_a21oi_1 _23370_ (.A1(_06732_),
    .A2(_06751_),
    .Y(_00405_),
    .B1(_06753_));
 sg13g2_a22oi_1 _23371_ (.Y(_06754_),
    .B1(net376),
    .B2(\top_ihp.oisc.regs[51][26] ),
    .A2(net400),
    .A1(\top_ihp.oisc.regs[63][26] ));
 sg13g2_a22oi_1 _23372_ (.Y(_06755_),
    .B1(_05810_),
    .B2(\top_ihp.oisc.regs[52][26] ),
    .A2(net414),
    .A1(\top_ihp.oisc.regs[30][26] ));
 sg13g2_a22oi_1 _23373_ (.Y(_06756_),
    .B1(net383),
    .B2(\top_ihp.oisc.regs[60][26] ),
    .A2(_05617_),
    .A1(\top_ihp.oisc.regs[34][26] ));
 sg13g2_a22oi_1 _23374_ (.Y(_06757_),
    .B1(_05978_),
    .B2(\top_ihp.oisc.regs[35][26] ),
    .A2(net416),
    .A1(\top_ihp.oisc.regs[42][26] ));
 sg13g2_nand4_1 _23375_ (.B(_06755_),
    .C(_06756_),
    .A(_06754_),
    .Y(_06758_),
    .D(_06757_));
 sg13g2_a22oi_1 _23376_ (.Y(_06759_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[39][26] ),
    .A2(net199),
    .A1(\top_ihp.oisc.regs[50][26] ));
 sg13g2_a22oi_1 _23377_ (.Y(_06760_),
    .B1(net161),
    .B2(\top_ihp.oisc.regs[44][26] ),
    .A2(net192),
    .A1(\top_ihp.oisc.regs[62][26] ));
 sg13g2_a22oi_1 _23378_ (.Y(_06761_),
    .B1(net191),
    .B2(\top_ihp.oisc.regs[59][26] ),
    .A2(net377),
    .A1(\top_ihp.oisc.regs[53][26] ));
 sg13g2_a22oi_1 _23379_ (.Y(_06762_),
    .B1(net404),
    .B2(\top_ihp.oisc.regs[49][26] ),
    .A2(_05986_),
    .A1(\top_ihp.oisc.regs[40][26] ));
 sg13g2_nand4_1 _23380_ (.B(_06760_),
    .C(_06761_),
    .A(_06759_),
    .Y(_06763_),
    .D(_06762_));
 sg13g2_nand2_1 _23381_ (.Y(_06764_),
    .A(\top_ihp.oisc.regs[33][26] ),
    .B(net407));
 sg13g2_a22oi_1 _23382_ (.Y(_06765_),
    .B1(net395),
    .B2(\top_ihp.oisc.regs[41][26] ),
    .A2(net339),
    .A1(\top_ihp.oisc.regs[38][26] ));
 sg13g2_nand3_1 _23383_ (.B(_06764_),
    .C(_06765_),
    .A(net57),
    .Y(_06766_));
 sg13g2_a22oi_1 _23384_ (.Y(_06767_),
    .B1(net363),
    .B2(\top_ihp.oisc.regs[32][26] ),
    .A2(net190),
    .A1(\top_ihp.oisc.regs[61][26] ));
 sg13g2_a22oi_1 _23385_ (.Y(_06768_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[27][26] ),
    .A2(net387),
    .A1(\top_ihp.oisc.regs[47][26] ));
 sg13g2_a22oi_1 _23386_ (.Y(_06769_),
    .B1(net398),
    .B2(\top_ihp.oisc.regs[55][26] ),
    .A2(net362),
    .A1(\top_ihp.oisc.regs[43][26] ));
 sg13g2_a22oi_1 _23387_ (.Y(_06770_),
    .B1(net396),
    .B2(\top_ihp.oisc.regs[46][26] ),
    .A2(net417),
    .A1(\top_ihp.oisc.regs[57][26] ));
 sg13g2_nand4_1 _23388_ (.B(_06768_),
    .C(_06769_),
    .A(_06767_),
    .Y(_06771_),
    .D(_06770_));
 sg13g2_nor4_2 _23389_ (.A(_06758_),
    .B(_06763_),
    .C(_06766_),
    .Y(_06772_),
    .D(_06771_));
 sg13g2_mux2_1 _23390_ (.A0(\top_ihp.oisc.regs[6][26] ),
    .A1(\top_ihp.oisc.regs[2][26] ),
    .S(net541),
    .X(_06773_));
 sg13g2_a22oi_1 _23391_ (.Y(_06774_),
    .B1(_05748_),
    .B2(_06773_),
    .A2(net390),
    .A1(\top_ihp.oisc.regs[13][26] ));
 sg13g2_a22oi_1 _23392_ (.Y(_06775_),
    .B1(net535),
    .B2(\top_ihp.oisc.regs[28][26] ),
    .A2(net533),
    .A1(\top_ihp.oisc.regs[22][26] ));
 sg13g2_a22oi_1 _23393_ (.Y(_06776_),
    .B1(net163),
    .B2(\top_ihp.oisc.regs[4][26] ),
    .A2(net368),
    .A1(\top_ihp.oisc.regs[25][26] ));
 sg13g2_a22oi_1 _23394_ (.Y(_06777_),
    .B1(_05531_),
    .B2(\top_ihp.oisc.regs[29][26] ),
    .A2(net547),
    .A1(\top_ihp.oisc.regs[1][26] ));
 sg13g2_nand4_1 _23395_ (.B(_06775_),
    .C(_06776_),
    .A(_06774_),
    .Y(_06778_),
    .D(_06777_));
 sg13g2_nand2_1 _23396_ (.Y(_06779_),
    .A(\top_ihp.oisc.regs[45][26] ),
    .B(net394));
 sg13g2_a22oi_1 _23397_ (.Y(_06780_),
    .B1(net160),
    .B2(\top_ihp.oisc.regs[17][26] ),
    .A2(net783),
    .A1(_07980_));
 sg13g2_a22oi_1 _23398_ (.Y(_06781_),
    .B1(_06426_),
    .B2(\top_ihp.oisc.regs[10][26] ),
    .A2(net374),
    .A1(\top_ihp.oisc.regs[9][26] ));
 sg13g2_nand3_1 _23399_ (.B(net750),
    .C(net549),
    .A(\top_ihp.oisc.regs[21][26] ),
    .Y(_06782_));
 sg13g2_nand3_1 _23400_ (.B(net548),
    .C(net747),
    .A(\top_ihp.oisc.regs[8][26] ),
    .Y(_06783_));
 sg13g2_nand2_1 _23401_ (.Y(_06784_),
    .A(_06782_),
    .B(_06783_));
 sg13g2_a22oi_1 _23402_ (.Y(_06785_),
    .B1(_06784_),
    .B2(_05520_),
    .A2(_06271_),
    .A1(\top_ihp.oisc.regs[19][26] ));
 sg13g2_nand4_1 _23403_ (.B(_06780_),
    .C(_06781_),
    .A(_06779_),
    .Y(_06786_),
    .D(_06785_));
 sg13g2_a22oi_1 _23404_ (.Y(_06787_),
    .B1(net181),
    .B2(\top_ihp.oisc.regs[15][26] ),
    .A2(net170),
    .A1(\top_ihp.oisc.regs[3][26] ));
 sg13g2_nand2_1 _23405_ (.Y(_06788_),
    .A(\top_ihp.oisc.regs[7][26] ),
    .B(net342));
 sg13g2_a22oi_1 _23406_ (.Y(_06789_),
    .B1(net173),
    .B2(\top_ihp.oisc.regs[11][26] ),
    .A2(net534),
    .A1(\top_ihp.oisc.regs[18][26] ));
 sg13g2_nand3_1 _23407_ (.B(net750),
    .C(net672),
    .A(\top_ihp.oisc.regs[23][26] ),
    .Y(_06790_));
 sg13g2_nand3_1 _23408_ (.B(_05519_),
    .C(net724),
    .A(\top_ihp.oisc.regs[5][26] ),
    .Y(_06791_));
 sg13g2_nand2_1 _23409_ (.Y(_06792_),
    .A(_06790_),
    .B(_06791_));
 sg13g2_mux2_1 _23410_ (.A0(\top_ihp.oisc.regs[14][26] ),
    .A1(\top_ihp.oisc.regs[12][26] ),
    .S(net669),
    .X(_06793_));
 sg13g2_a22oi_1 _23411_ (.Y(_06794_),
    .B1(_06793_),
    .B2(_06484_),
    .A2(_06792_),
    .A1(net549));
 sg13g2_nand4_1 _23412_ (.B(_06788_),
    .C(_06789_),
    .A(_06787_),
    .Y(_06795_),
    .D(_06794_));
 sg13g2_mux2_1 _23413_ (.A0(\top_ihp.oisc.regs[26][26] ),
    .A1(\top_ihp.oisc.regs[24][26] ),
    .S(net545),
    .X(_06796_));
 sg13g2_a22oi_1 _23414_ (.Y(_06797_),
    .B1(_06796_),
    .B2(net727),
    .A2(_05582_),
    .A1(\top_ihp.oisc.regs[16][26] ));
 sg13g2_a22oi_1 _23415_ (.Y(_06798_),
    .B1(_05804_),
    .B2(\top_ihp.oisc.regs[56][26] ),
    .A2(_05460_),
    .A1(\top_ihp.oisc.regs[31][26] ));
 sg13g2_a22oi_1 _23416_ (.Y(_06799_),
    .B1(_05651_),
    .B2(\top_ihp.oisc.regs[54][26] ),
    .A2(_05472_),
    .A1(\top_ihp.oisc.regs[20][26] ));
 sg13g2_a22oi_1 _23417_ (.Y(_06800_),
    .B1(_05789_),
    .B2(\top_ihp.oisc.regs[58][26] ),
    .A2(_05713_),
    .A1(\top_ihp.oisc.regs[48][26] ));
 sg13g2_a22oi_1 _23418_ (.Y(_06801_),
    .B1(_05595_),
    .B2(\top_ihp.oisc.regs[37][26] ),
    .A2(_05455_),
    .A1(\top_ihp.oisc.regs[36][26] ));
 sg13g2_and4_1 _23419_ (.A(_06798_),
    .B(_06799_),
    .C(_06800_),
    .D(_06801_),
    .X(_06802_));
 sg13g2_o21ai_1 _23420_ (.B1(_06802_),
    .Y(_06803_),
    .A1(_05537_),
    .A2(_06797_));
 sg13g2_nor4_1 _23421_ (.A(_06778_),
    .B(_06786_),
    .C(_06795_),
    .D(_06803_),
    .Y(_06804_));
 sg13g2_nand2_1 _23422_ (.Y(_06805_),
    .A(_00230_),
    .B(_06008_));
 sg13g2_a22oi_1 _23423_ (.Y(_06806_),
    .B1(_05943_),
    .B2(_06805_),
    .A2(_06304_),
    .A1(_07980_));
 sg13g2_a21oi_1 _23424_ (.A1(_06772_),
    .A2(_06804_),
    .Y(_00406_),
    .B1(_06806_));
 sg13g2_a22oi_1 _23425_ (.Y(_06807_),
    .B1(net193),
    .B2(\top_ihp.oisc.regs[56][27] ),
    .A2(net403),
    .A1(\top_ihp.oisc.regs[55][27] ));
 sg13g2_a22oi_1 _23426_ (.Y(_06808_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[47][27] ),
    .A2(net175),
    .A1(\top_ihp.oisc.regs[61][27] ));
 sg13g2_a22oi_1 _23427_ (.Y(_06809_),
    .B1(net370),
    .B2(\top_ihp.oisc.regs[13][27] ),
    .A2(net544),
    .A1(\top_ihp.oisc.regs[18][27] ));
 sg13g2_a22oi_1 _23428_ (.Y(_06810_),
    .B1(_05562_),
    .B2(\top_ihp.oisc.regs[9][27] ),
    .A2(_05481_),
    .A1(\top_ihp.oisc.regs[25][27] ));
 sg13g2_a22oi_1 _23429_ (.Y(_06811_),
    .B1(_05750_),
    .B2(\top_ihp.oisc.regs[2][27] ),
    .A2(net668),
    .A1(\top_ihp.oisc.regs[28][27] ));
 sg13g2_a22oi_1 _23430_ (.Y(_06812_),
    .B1(net552),
    .B2(\top_ihp.oisc.regs[20][27] ),
    .A2(net553),
    .A1(\top_ihp.oisc.regs[22][27] ));
 sg13g2_and4_1 _23431_ (.A(_06809_),
    .B(_06810_),
    .C(_06811_),
    .D(_06812_),
    .X(_06813_));
 sg13g2_nand3_1 _23432_ (.B(_06808_),
    .C(_06813_),
    .A(_06807_),
    .Y(_06814_));
 sg13g2_a22oi_1 _23433_ (.Y(_06815_),
    .B1(_06276_),
    .B2(\top_ihp.oisc.regs[10][27] ),
    .A2(net367),
    .A1(\top_ihp.oisc.regs[26][27] ));
 sg13g2_a22oi_1 _23434_ (.Y(_06816_),
    .B1(_05914_),
    .B2(\top_ihp.oisc.regs[8][27] ),
    .A2(net720),
    .A1(\top_ihp.oisc.regs[23][27] ));
 sg13g2_nand2_1 _23435_ (.Y(_06817_),
    .A(\top_ihp.oisc.regs[60][27] ),
    .B(net171));
 sg13g2_nand4_1 _23436_ (.B(_06815_),
    .C(_06816_),
    .A(net61),
    .Y(_06818_),
    .D(_06817_));
 sg13g2_a22oi_1 _23437_ (.Y(_06819_),
    .B1(_05596_),
    .B2(\top_ihp.oisc.regs[37][27] ),
    .A2(_05787_),
    .A1(\top_ihp.oisc.regs[54][27] ));
 sg13g2_a22oi_1 _23438_ (.Y(_06820_),
    .B1(net412),
    .B2(\top_ihp.oisc.regs[43][27] ),
    .A2(_05648_),
    .A1(\top_ihp.oisc.regs[53][27] ));
 sg13g2_a22oi_1 _23439_ (.Y(_06821_),
    .B1(net177),
    .B2(\top_ihp.oisc.regs[58][27] ),
    .A2(net378),
    .A1(\top_ihp.oisc.regs[38][27] ));
 sg13g2_a22oi_1 _23440_ (.Y(_06822_),
    .B1(net366),
    .B2(\top_ihp.oisc.regs[49][27] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[40][27] ));
 sg13g2_nand4_1 _23441_ (.B(_06820_),
    .C(_06821_),
    .A(_06819_),
    .Y(_06823_),
    .D(_06822_));
 sg13g2_a22oi_1 _23442_ (.Y(_06824_),
    .B1(net394),
    .B2(\top_ihp.oisc.regs[45][27] ),
    .A2(_05799_),
    .A1(\top_ihp.oisc.regs[50][27] ));
 sg13g2_a22oi_1 _23443_ (.Y(_06825_),
    .B1(net405),
    .B2(\top_ihp.oisc.regs[52][27] ),
    .A2(net360),
    .A1(\top_ihp.oisc.regs[33][27] ));
 sg13g2_a22oi_1 _23444_ (.Y(_06826_),
    .B1(net395),
    .B2(\top_ihp.oisc.regs[41][27] ),
    .A2(net539),
    .A1(\top_ihp.oisc.regs[34][27] ));
 sg13g2_a22oi_1 _23445_ (.Y(_06827_),
    .B1(_05629_),
    .B2(\top_ihp.oisc.regs[44][27] ),
    .A2(net356),
    .A1(\top_ihp.oisc.regs[31][27] ));
 sg13g2_nand4_1 _23446_ (.B(_06825_),
    .C(_06826_),
    .A(_06824_),
    .Y(_06828_),
    .D(_06827_));
 sg13g2_nor4_2 _23447_ (.A(_06814_),
    .B(_06818_),
    .C(_06823_),
    .Y(_06829_),
    .D(_06828_));
 sg13g2_a22oi_1 _23448_ (.Y(_06830_),
    .B1(_05761_),
    .B2(\top_ihp.oisc.regs[5][27] ),
    .A2(_05505_),
    .A1(\top_ihp.oisc.regs[1][27] ));
 sg13g2_a22oi_1 _23449_ (.Y(_06831_),
    .B1(_05759_),
    .B2(\top_ihp.oisc.regs[16][27] ),
    .A2(_05570_),
    .A1(\top_ihp.oisc.regs[15][27] ));
 sg13g2_a22oi_1 _23450_ (.Y(_06832_),
    .B1(_05565_),
    .B2(\top_ihp.oisc.regs[6][27] ),
    .A2(net554),
    .A1(\top_ihp.oisc.regs[7][27] ));
 sg13g2_a22oi_1 _23451_ (.Y(_06833_),
    .B1(_05556_),
    .B2(\top_ihp.oisc.regs[3][27] ),
    .A2(_05550_),
    .A1(\top_ihp.oisc.regs[19][27] ));
 sg13g2_and4_1 _23452_ (.A(_06830_),
    .B(_06831_),
    .C(_06832_),
    .D(_06833_),
    .X(_06834_));
 sg13g2_a22oi_1 _23453_ (.Y(_06835_),
    .B1(net182),
    .B2(\top_ihp.oisc.regs[29][27] ),
    .A2(_05515_),
    .A1(\top_ihp.oisc.regs[14][27] ));
 sg13g2_a22oi_1 _23454_ (.Y(_06836_),
    .B1(net167),
    .B2(\top_ihp.oisc.regs[24][27] ),
    .A2(net372),
    .A1(\top_ihp.oisc.regs[12][27] ));
 sg13g2_nand3_1 _23455_ (.B(_06835_),
    .C(_06836_),
    .A(_06834_),
    .Y(_06837_));
 sg13g2_nand2_1 _23456_ (.Y(_06838_),
    .A(\top_ihp.oisc.regs[11][27] ),
    .B(net169));
 sg13g2_a22oi_1 _23457_ (.Y(_06839_),
    .B1(_05821_),
    .B2(\top_ihp.oisc.regs[21][27] ),
    .A2(net803),
    .A1(_08290_));
 sg13g2_a22oi_1 _23458_ (.Y(_06840_),
    .B1(net160),
    .B2(\top_ihp.oisc.regs[17][27] ),
    .A2(net432),
    .A1(\top_ihp.oisc.regs[4][27] ));
 sg13g2_a22oi_1 _23459_ (.Y(_06841_),
    .B1(net381),
    .B2(\top_ihp.oisc.regs[48][27] ),
    .A2(net186),
    .A1(\top_ihp.oisc.regs[59][27] ));
 sg13g2_nand4_1 _23460_ (.B(_06839_),
    .C(_06840_),
    .A(_06838_),
    .Y(_06842_),
    .D(_06841_));
 sg13g2_a22oi_1 _23461_ (.Y(_06843_),
    .B1(net361),
    .B2(\top_ihp.oisc.regs[35][27] ),
    .A2(_05939_),
    .A1(\top_ihp.oisc.regs[62][27] ));
 sg13g2_a22oi_1 _23462_ (.Y(_06844_),
    .B1(net396),
    .B2(\top_ihp.oisc.regs[46][27] ),
    .A2(net365),
    .A1(\top_ihp.oisc.regs[63][27] ));
 sg13g2_nand2_1 _23463_ (.Y(_06845_),
    .A(_06843_),
    .B(_06844_));
 sg13g2_a22oi_1 _23464_ (.Y(_06846_),
    .B1(net354),
    .B2(\top_ihp.oisc.regs[39][27] ),
    .A2(_05954_),
    .A1(\top_ihp.oisc.regs[36][27] ));
 sg13g2_a22oi_1 _23465_ (.Y(_06847_),
    .B1(net355),
    .B2(\top_ihp.oisc.regs[51][27] ),
    .A2(net422),
    .A1(\top_ihp.oisc.regs[32][27] ));
 sg13g2_a22oi_1 _23466_ (.Y(_06848_),
    .B1(_05835_),
    .B2(\top_ihp.oisc.regs[30][27] ),
    .A2(net336),
    .A1(\top_ihp.oisc.regs[42][27] ));
 sg13g2_a22oi_1 _23467_ (.Y(_06849_),
    .B1(_05609_),
    .B2(\top_ihp.oisc.regs[27][27] ),
    .A2(net417),
    .A1(\top_ihp.oisc.regs[57][27] ));
 sg13g2_nand4_1 _23468_ (.B(_06847_),
    .C(_06848_),
    .A(_06846_),
    .Y(_06850_),
    .D(_06849_));
 sg13g2_nor4_1 _23469_ (.A(_06837_),
    .B(_06842_),
    .C(_06845_),
    .D(_06850_),
    .Y(_06851_));
 sg13g2_nand2_1 _23470_ (.Y(_06852_),
    .A(_00231_),
    .B(net59));
 sg13g2_a22oi_1 _23471_ (.Y(_06853_),
    .B1(net26),
    .B2(_06852_),
    .A2(net746),
    .A1(_08290_));
 sg13g2_a21oi_1 _23472_ (.A1(_06829_),
    .A2(_06851_),
    .Y(_00407_),
    .B1(_06853_));
 sg13g2_a22oi_1 _23473_ (.Y(_06854_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[32][28] ),
    .A2(net346),
    .A1(\top_ihp.oisc.regs[30][28] ));
 sg13g2_a22oi_1 _23474_ (.Y(_06855_),
    .B1(net364),
    .B2(\top_ihp.oisc.regs[52][28] ),
    .A2(_05456_),
    .A1(\top_ihp.oisc.regs[36][28] ));
 sg13g2_a22oi_1 _23475_ (.Y(_06856_),
    .B1(net198),
    .B2(\top_ihp.oisc.regs[59][28] ),
    .A2(net351),
    .A1(\top_ihp.oisc.regs[40][28] ));
 sg13g2_a22oi_1 _23476_ (.Y(_06857_),
    .B1(net391),
    .B2(\top_ihp.oisc.regs[33][28] ),
    .A2(_05978_),
    .A1(\top_ihp.oisc.regs[35][28] ));
 sg13g2_nand4_1 _23477_ (.B(_06855_),
    .C(_06856_),
    .A(_06854_),
    .Y(_06858_),
    .D(_06857_));
 sg13g2_a22oi_1 _23478_ (.Y(_06859_),
    .B1(net410),
    .B2(\top_ihp.oisc.regs[41][28] ),
    .A2(net419),
    .A1(\top_ihp.oisc.regs[44][28] ));
 sg13g2_a22oi_1 _23479_ (.Y(_06860_),
    .B1(net383),
    .B2(\top_ihp.oisc.regs[60][28] ),
    .A2(net201),
    .A1(\top_ihp.oisc.regs[54][28] ));
 sg13g2_a22oi_1 _23480_ (.Y(_06861_),
    .B1(net404),
    .B2(\top_ihp.oisc.regs[49][28] ),
    .A2(net377),
    .A1(\top_ihp.oisc.regs[53][28] ));
 sg13g2_a22oi_1 _23481_ (.Y(_06862_),
    .B1(net400),
    .B2(\top_ihp.oisc.regs[63][28] ),
    .A2(net333),
    .A1(\top_ihp.oisc.regs[57][28] ));
 sg13g2_nand4_1 _23482_ (.B(_06860_),
    .C(_06861_),
    .A(_06859_),
    .Y(_06863_),
    .D(_06862_));
 sg13g2_nand2_1 _23483_ (.Y(_06864_),
    .A(\top_ihp.oisc.regs[61][28] ),
    .B(_05836_));
 sg13g2_a22oi_1 _23484_ (.Y(_06865_),
    .B1(net355),
    .B2(\top_ihp.oisc.regs[51][28] ),
    .A2(net397),
    .A1(\top_ihp.oisc.regs[37][28] ));
 sg13g2_nand3_1 _23485_ (.B(_06864_),
    .C(_06865_),
    .A(net57),
    .Y(_06866_));
 sg13g2_a22oi_1 _23486_ (.Y(_06867_),
    .B1(net719),
    .B2(\top_ihp.oisc.regs[23][28] ),
    .A2(net663),
    .A1(\top_ihp.oisc.regs[21][28] ));
 sg13g2_nand2_1 _23487_ (.Y(_06868_),
    .A(_08276_),
    .B(net801));
 sg13g2_nand2_1 _23488_ (.Y(_06869_),
    .A(_06867_),
    .B(_06868_));
 sg13g2_a221oi_1 _23489_ (.B2(\top_ihp.oisc.regs[5][28] ),
    .C1(_06869_),
    .B1(net345),
    .A1(\top_ihp.oisc.regs[1][28] ),
    .Y(_06870_),
    .A2(_05507_));
 sg13g2_a22oi_1 _23490_ (.Y(_06871_),
    .B1(net354),
    .B2(\top_ihp.oisc.regs[39][28] ),
    .A2(net387),
    .A1(\top_ihp.oisc.regs[47][28] ));
 sg13g2_a22oi_1 _23491_ (.Y(_06872_),
    .B1(net194),
    .B2(\top_ihp.oisc.regs[50][28] ),
    .A2(net362),
    .A1(\top_ihp.oisc.regs[43][28] ));
 sg13g2_a22oi_1 _23492_ (.Y(_06873_),
    .B1(net349),
    .B2(\top_ihp.oisc.regs[46][28] ),
    .A2(net336),
    .A1(\top_ihp.oisc.regs[42][28] ));
 sg13g2_nand4_1 _23493_ (.B(_06871_),
    .C(_06872_),
    .A(_06870_),
    .Y(_06874_),
    .D(_06873_));
 sg13g2_nor4_2 _23494_ (.A(_06858_),
    .B(_06863_),
    .C(_06866_),
    .Y(_06875_),
    .D(_06874_));
 sg13g2_a22oi_1 _23495_ (.Y(_06876_),
    .B1(net339),
    .B2(\top_ihp.oisc.regs[38][28] ),
    .A2(_05654_),
    .A1(\top_ihp.oisc.regs[56][28] ));
 sg13g2_a22oi_1 _23496_ (.Y(_06877_),
    .B1(net359),
    .B2(\top_ihp.oisc.regs[55][28] ),
    .A2(net411),
    .A1(\top_ihp.oisc.regs[45][28] ));
 sg13g2_a22oi_1 _23497_ (.Y(_06878_),
    .B1(net341),
    .B2(\top_ihp.oisc.regs[27][28] ),
    .A2(net174),
    .A1(\top_ihp.oisc.regs[62][28] ));
 sg13g2_a22oi_1 _23498_ (.Y(_06879_),
    .B1(net399),
    .B2(\top_ihp.oisc.regs[58][28] ),
    .A2(_05460_),
    .A1(\top_ihp.oisc.regs[31][28] ));
 sg13g2_nand4_1 _23499_ (.B(_06877_),
    .C(_06878_),
    .A(_06876_),
    .Y(_06880_),
    .D(_06879_));
 sg13g2_a22oi_1 _23500_ (.Y(_06881_),
    .B1(net381),
    .B2(\top_ihp.oisc.regs[48][28] ),
    .A2(net542),
    .A1(\top_ihp.oisc.regs[34][28] ));
 sg13g2_a22oi_1 _23501_ (.Y(_06882_),
    .B1(_05514_),
    .B2(\top_ihp.oisc.regs[14][28] ),
    .A2(net553),
    .A1(\top_ihp.oisc.regs[22][28] ));
 sg13g2_a22oi_1 _23502_ (.Y(_06883_),
    .B1(_05775_),
    .B2(\top_ihp.oisc.regs[24][28] ),
    .A2(net668),
    .A1(\top_ihp.oisc.regs[28][28] ));
 sg13g2_and2_1 _23503_ (.A(_06882_),
    .B(_06883_),
    .X(_06884_));
 sg13g2_a22oi_1 _23504_ (.Y(_06885_),
    .B1(net371),
    .B2(\top_ihp.oisc.regs[16][28] ),
    .A2(net401),
    .A1(\top_ihp.oisc.regs[3][28] ));
 sg13g2_a22oi_1 _23505_ (.Y(_06886_),
    .B1(net665),
    .B2(\top_ihp.oisc.regs[8][28] ),
    .A2(net368),
    .A1(\top_ihp.oisc.regs[25][28] ));
 sg13g2_nand4_1 _23506_ (.B(_06884_),
    .C(_06885_),
    .A(_06881_),
    .Y(_06887_),
    .D(_06886_));
 sg13g2_a22oi_1 _23507_ (.Y(_06888_),
    .B1(net343),
    .B2(\top_ihp.oisc.regs[18][28] ),
    .A2(net342),
    .A1(\top_ihp.oisc.regs[7][28] ));
 sg13g2_a22oi_1 _23508_ (.Y(_06889_),
    .B1(net350),
    .B2(\top_ihp.oisc.regs[19][28] ),
    .A2(net163),
    .A1(\top_ihp.oisc.regs[4][28] ));
 sg13g2_a22oi_1 _23509_ (.Y(_06890_),
    .B1(net334),
    .B2(\top_ihp.oisc.regs[10][28] ),
    .A2(net203),
    .A1(\top_ihp.oisc.regs[29][28] ));
 sg13g2_a22oi_1 _23510_ (.Y(_06891_),
    .B1(net184),
    .B2(\top_ihp.oisc.regs[12][28] ),
    .A2(net540),
    .A1(\top_ihp.oisc.regs[20][28] ));
 sg13g2_nand4_1 _23511_ (.B(_06889_),
    .C(_06890_),
    .A(_06888_),
    .Y(_06892_),
    .D(_06891_));
 sg13g2_a22oi_1 _23512_ (.Y(_06893_),
    .B1(net179),
    .B2(\top_ihp.oisc.regs[2][28] ),
    .A2(_05999_),
    .A1(\top_ihp.oisc.regs[17][28] ));
 sg13g2_a22oi_1 _23513_ (.Y(_06894_),
    .B1(net538),
    .B2(\top_ihp.oisc.regs[6][28] ),
    .A2(net180),
    .A1(\top_ihp.oisc.regs[13][28] ));
 sg13g2_a22oi_1 _23514_ (.Y(_06895_),
    .B1(net173),
    .B2(\top_ihp.oisc.regs[11][28] ),
    .A2(net164),
    .A1(\top_ihp.oisc.regs[9][28] ));
 sg13g2_a22oi_1 _23515_ (.Y(_06896_),
    .B1(net168),
    .B2(\top_ihp.oisc.regs[26][28] ),
    .A2(net162),
    .A1(\top_ihp.oisc.regs[15][28] ));
 sg13g2_nand4_1 _23516_ (.B(_06894_),
    .C(_06895_),
    .A(_06893_),
    .Y(_06897_),
    .D(_06896_));
 sg13g2_nor4_1 _23517_ (.A(_06880_),
    .B(_06887_),
    .C(_06892_),
    .D(_06897_),
    .Y(_06898_));
 sg13g2_a21o_1 _23518_ (.A2(net63),
    .A1(_00069_),
    .B1(net58),
    .X(_06899_));
 sg13g2_a22oi_1 _23519_ (.Y(_00408_),
    .B1(_06899_),
    .B2(_06868_),
    .A2(_06898_),
    .A1(_06875_));
 sg13g2_a22oi_1 _23520_ (.Y(_06900_),
    .B1(net349),
    .B2(\top_ihp.oisc.regs[46][29] ),
    .A2(_06141_),
    .A1(\top_ihp.oisc.regs[32][29] ));
 sg13g2_a22oi_1 _23521_ (.Y(_06901_),
    .B1(net161),
    .B2(\top_ihp.oisc.regs[44][29] ),
    .A2(net414),
    .A1(\top_ihp.oisc.regs[30][29] ));
 sg13g2_a22oi_1 _23522_ (.Y(_06902_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[39][29] ),
    .A2(net201),
    .A1(\top_ihp.oisc.regs[54][29] ));
 sg13g2_a22oi_1 _23523_ (.Y(_06903_),
    .B1(net382),
    .B2(\top_ihp.oisc.regs[27][29] ),
    .A2(_05983_),
    .A1(\top_ihp.oisc.regs[62][29] ));
 sg13g2_nand4_1 _23524_ (.B(_06901_),
    .C(_06902_),
    .A(_06900_),
    .Y(_06904_),
    .D(_06903_));
 sg13g2_a22oi_1 _23525_ (.Y(_06905_),
    .B1(_05848_),
    .B2(\top_ihp.oisc.regs[60][29] ),
    .A2(_05733_),
    .A1(\top_ihp.oisc.regs[49][29] ));
 sg13g2_a22oi_1 _23526_ (.Y(_06906_),
    .B1(net336),
    .B2(\top_ihp.oisc.regs[42][29] ),
    .A2(_05636_),
    .A1(\top_ihp.oisc.regs[40][29] ));
 sg13g2_a22oi_1 _23527_ (.Y(_06907_),
    .B1(_05855_),
    .B2(\top_ihp.oisc.regs[48][29] ),
    .A2(net347),
    .A1(\top_ihp.oisc.regs[37][29] ));
 sg13g2_a22oi_1 _23528_ (.Y(_06908_),
    .B1(_06086_),
    .B2(\top_ihp.oisc.regs[41][29] ),
    .A2(_05601_),
    .A1(\top_ihp.oisc.regs[47][29] ));
 sg13g2_nand4_1 _23529_ (.B(_06906_),
    .C(_06907_),
    .A(_06905_),
    .Y(_06909_),
    .D(_06908_));
 sg13g2_nand2_1 _23530_ (.Y(_06910_),
    .A(\top_ihp.oisc.regs[35][29] ),
    .B(net361));
 sg13g2_a22oi_1 _23531_ (.Y(_06911_),
    .B1(net384),
    .B2(\top_ihp.oisc.regs[38][29] ),
    .A2(net356),
    .A1(\top_ihp.oisc.regs[31][29] ));
 sg13g2_nand3_1 _23532_ (.B(_06910_),
    .C(_06911_),
    .A(net57),
    .Y(_06912_));
 sg13g2_a22oi_1 _23533_ (.Y(_06913_),
    .B1(net719),
    .B2(\top_ihp.oisc.regs[23][29] ),
    .A2(net663),
    .A1(\top_ihp.oisc.regs[21][29] ));
 sg13g2_o21ai_1 _23534_ (.B1(_06913_),
    .Y(_06914_),
    .A1(_08332_),
    .A2(net804));
 sg13g2_a221oi_1 _23535_ (.B2(\top_ihp.oisc.regs[5][29] ),
    .C1(_06914_),
    .B1(net345),
    .A1(\top_ihp.oisc.regs[20][29] ),
    .Y(_06915_),
    .A2(_05782_));
 sg13g2_a22oi_1 _23536_ (.Y(_06916_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[34][29] ),
    .A2(_06020_),
    .A1(\top_ihp.oisc.regs[57][29] ));
 sg13g2_a22oi_1 _23537_ (.Y(_06917_),
    .B1(net194),
    .B2(\top_ihp.oisc.regs[50][29] ),
    .A2(_05965_),
    .A1(\top_ihp.oisc.regs[61][29] ));
 sg13g2_a22oi_1 _23538_ (.Y(_06918_),
    .B1(net394),
    .B2(\top_ihp.oisc.regs[45][29] ),
    .A2(net365),
    .A1(\top_ihp.oisc.regs[63][29] ));
 sg13g2_nand4_1 _23539_ (.B(_06916_),
    .C(_06917_),
    .A(_06915_),
    .Y(_06919_),
    .D(_06918_));
 sg13g2_nor4_1 _23540_ (.A(_06904_),
    .B(_06909_),
    .C(_06912_),
    .D(_06919_),
    .Y(_06920_));
 sg13g2_a22oi_1 _23541_ (.Y(_06921_),
    .B1(net399),
    .B2(\top_ihp.oisc.regs[58][29] ),
    .A2(net420),
    .A1(\top_ihp.oisc.regs[51][29] ));
 sg13g2_a22oi_1 _23542_ (.Y(_06922_),
    .B1(net402),
    .B2(\top_ihp.oisc.regs[24][29] ),
    .A2(net390),
    .A1(\top_ihp.oisc.regs[13][29] ));
 sg13g2_a22oi_1 _23543_ (.Y(_06923_),
    .B1(_05857_),
    .B2(\top_ihp.oisc.regs[11][29] ),
    .A2(net431),
    .A1(\top_ihp.oisc.regs[1][29] ));
 sg13g2_mux2_1 _23544_ (.A0(\top_ihp.oisc.regs[12][29] ),
    .A1(\top_ihp.oisc.regs[8][29] ),
    .S(net670),
    .X(_06924_));
 sg13g2_a22oi_1 _23545_ (.Y(_06925_),
    .B1(_06924_),
    .B2(_05520_),
    .A2(net721),
    .A1(\top_ihp.oisc.regs[14][29] ));
 sg13g2_nand2b_1 _23546_ (.Y(_06926_),
    .B(net747),
    .A_N(_06925_));
 sg13g2_nand4_1 _23547_ (.B(_06922_),
    .C(_06923_),
    .A(_06921_),
    .Y(_06927_),
    .D(_06926_));
 sg13g2_a22oi_1 _23548_ (.Y(_06928_),
    .B1(net191),
    .B2(\top_ihp.oisc.regs[59][29] ),
    .A2(net375),
    .A1(\top_ihp.oisc.regs[36][29] ));
 sg13g2_a22oi_1 _23549_ (.Y(_06929_),
    .B1(net391),
    .B2(\top_ihp.oisc.regs[33][29] ),
    .A2(_05869_),
    .A1(\top_ihp.oisc.regs[53][29] ));
 sg13g2_a22oi_1 _23550_ (.Y(_06930_),
    .B1(net359),
    .B2(\top_ihp.oisc.regs[55][29] ),
    .A2(_05728_),
    .A1(\top_ihp.oisc.regs[52][29] ));
 sg13g2_a22oi_1 _23551_ (.Y(_06931_),
    .B1(_05804_),
    .B2(\top_ihp.oisc.regs[56][29] ),
    .A2(_05669_),
    .A1(\top_ihp.oisc.regs[43][29] ));
 sg13g2_nand4_1 _23552_ (.B(_06929_),
    .C(_06930_),
    .A(_06928_),
    .Y(_06932_),
    .D(_06931_));
 sg13g2_a22oi_1 _23553_ (.Y(_06933_),
    .B1(net334),
    .B2(\top_ihp.oisc.regs[10][29] ),
    .A2(net342),
    .A1(\top_ihp.oisc.regs[7][29] ));
 sg13g2_a22oi_1 _23554_ (.Y(_06934_),
    .B1(net168),
    .B2(\top_ihp.oisc.regs[26][29] ),
    .A2(net369),
    .A1(\top_ihp.oisc.regs[2][29] ));
 sg13g2_a22oi_1 _23555_ (.Y(_06935_),
    .B1(net160),
    .B2(\top_ihp.oisc.regs[17][29] ),
    .A2(net335),
    .A1(\top_ihp.oisc.regs[19][29] ));
 sg13g2_a22oi_1 _23556_ (.Y(_06936_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[25][29] ),
    .A2(net533),
    .A1(\top_ihp.oisc.regs[22][29] ));
 sg13g2_nand4_1 _23557_ (.B(_06934_),
    .C(_06935_),
    .A(_06933_),
    .Y(_06937_),
    .D(_06936_));
 sg13g2_a22oi_1 _23558_ (.Y(_06938_),
    .B1(net538),
    .B2(\top_ihp.oisc.regs[6][29] ),
    .A2(net535),
    .A1(\top_ihp.oisc.regs[28][29] ));
 sg13g2_a22oi_1 _23559_ (.Y(_06939_),
    .B1(net183),
    .B2(\top_ihp.oisc.regs[16][29] ),
    .A2(_06063_),
    .A1(\top_ihp.oisc.regs[18][29] ));
 sg13g2_a22oi_1 _23560_ (.Y(_06940_),
    .B1(_05895_),
    .B2(\top_ihp.oisc.regs[29][29] ),
    .A2(net204),
    .A1(\top_ihp.oisc.regs[4][29] ));
 sg13g2_nand3_1 _23561_ (.B(_05443_),
    .C(_05510_),
    .A(\top_ihp.oisc.regs[15][29] ),
    .Y(_06941_));
 sg13g2_nand3_1 _23562_ (.B(net548),
    .C(_05523_),
    .A(\top_ihp.oisc.regs[3][29] ),
    .Y(_06942_));
 sg13g2_o21ai_1 _23563_ (.B1(_06942_),
    .Y(_06943_),
    .A1(net541),
    .A2(_06941_));
 sg13g2_a22oi_1 _23564_ (.Y(_06944_),
    .B1(_06943_),
    .B2(_05486_),
    .A2(net164),
    .A1(\top_ihp.oisc.regs[9][29] ));
 sg13g2_nand4_1 _23565_ (.B(_06939_),
    .C(_06940_),
    .A(_06938_),
    .Y(_06945_),
    .D(_06944_));
 sg13g2_nor4_1 _23566_ (.A(_06927_),
    .B(_06932_),
    .C(_06937_),
    .D(_06945_),
    .Y(_06946_));
 sg13g2_nand2_1 _23567_ (.Y(_06947_),
    .A(_00070_),
    .B(_06008_));
 sg13g2_a22oi_1 _23568_ (.Y(_06948_),
    .B1(net26),
    .B2(_06947_),
    .A2(net746),
    .A1(_08320_));
 sg13g2_a21oi_1 _23569_ (.A1(_06920_),
    .A2(_06946_),
    .Y(_00409_),
    .B1(_06948_));
 sg13g2_a22oi_1 _23570_ (.Y(_06949_),
    .B1(net350),
    .B2(\top_ihp.oisc.regs[19][2] ),
    .A2(net434),
    .A1(\top_ihp.oisc.regs[20][2] ));
 sg13g2_nand2_1 _23571_ (.Y(_06950_),
    .A(\top_ihp.oisc.regs[9][2] ),
    .B(_05884_));
 sg13g2_a22oi_1 _23572_ (.Y(_06951_),
    .B1(net170),
    .B2(\top_ihp.oisc.regs[3][2] ),
    .A2(_06057_),
    .A1(\top_ihp.oisc.regs[28][2] ));
 sg13g2_nand3_1 _23573_ (.B(net669),
    .C(net724),
    .A(\top_ihp.oisc.regs[5][2] ),
    .Y(_06952_));
 sg13g2_nand3_1 _23574_ (.B(net550),
    .C(net747),
    .A(\top_ihp.oisc.regs[14][2] ),
    .Y(_06953_));
 sg13g2_nand2_1 _23575_ (.Y(_06954_),
    .A(_06952_),
    .B(_06953_));
 sg13g2_a22oi_1 _23576_ (.Y(_06955_),
    .B1(_06954_),
    .B2(net549),
    .A2(net432),
    .A1(\top_ihp.oisc.regs[4][2] ));
 sg13g2_nand4_1 _23577_ (.B(_06950_),
    .C(_06951_),
    .A(_06949_),
    .Y(_06956_),
    .D(_06955_));
 sg13g2_mux2_1 _23578_ (.A0(\top_ihp.oisc.regs[24][2] ),
    .A1(\top_ihp.oisc.regs[16][2] ),
    .S(net662),
    .X(_06957_));
 sg13g2_a22oi_1 _23579_ (.Y(_06958_),
    .B1(_06957_),
    .B2(_06277_),
    .A2(_06276_),
    .A1(\top_ihp.oisc.regs[10][2] ));
 sg13g2_a22oi_1 _23580_ (.Y(_06959_),
    .B1(net160),
    .B2(\top_ihp.oisc.regs[17][2] ),
    .A2(net203),
    .A1(\top_ihp.oisc.regs[29][2] ));
 sg13g2_a22oi_1 _23581_ (.Y(_06960_),
    .B1(net173),
    .B2(\top_ihp.oisc.regs[11][2] ),
    .A2(net390),
    .A1(\top_ihp.oisc.regs[13][2] ));
 sg13g2_nand3_1 _23582_ (.B(net550),
    .C(net749),
    .A(\top_ihp.oisc.regs[6][2] ),
    .Y(_06961_));
 sg13g2_nand3_1 _23583_ (.B(_05519_),
    .C(net747),
    .A(\top_ihp.oisc.regs[12][2] ),
    .Y(_06962_));
 sg13g2_nand2_1 _23584_ (.Y(_06963_),
    .A(_06961_),
    .B(_06962_));
 sg13g2_a22oi_1 _23585_ (.Y(_06964_),
    .B1(_06963_),
    .B2(net549),
    .A2(net534),
    .A1(\top_ihp.oisc.regs[18][2] ));
 sg13g2_nand4_1 _23586_ (.B(_06959_),
    .C(_06960_),
    .A(_06958_),
    .Y(_06965_),
    .D(_06964_));
 sg13g2_a22oi_1 _23587_ (.Y(_06966_),
    .B1(net363),
    .B2(\top_ihp.oisc.regs[32][2] ),
    .A2(net424),
    .A1(\top_ihp.oisc.regs[39][2] ));
 sg13g2_a22oi_1 _23588_ (.Y(_06967_),
    .B1(net394),
    .B2(\top_ihp.oisc.regs[45][2] ),
    .A2(net346),
    .A1(\top_ihp.oisc.regs[30][2] ));
 sg13g2_a22oi_1 _23589_ (.Y(_06968_),
    .B1(net428),
    .B2(\top_ihp.oisc.regs[15][2] ),
    .A2(_05482_),
    .A1(\top_ihp.oisc.regs[25][2] ));
 sg13g2_a22oi_1 _23590_ (.Y(_06969_),
    .B1(net367),
    .B2(\top_ihp.oisc.regs[26][2] ),
    .A2(net547),
    .A1(\top_ihp.oisc.regs[1][2] ));
 sg13g2_and2_1 _23591_ (.A(_06968_),
    .B(_06969_),
    .X(_06970_));
 sg13g2_a22oi_1 _23592_ (.Y(_06971_),
    .B1(net663),
    .B2(\top_ihp.oisc.regs[21][2] ),
    .A2(_06023_),
    .A1(_08090_));
 sg13g2_inv_1 _23593_ (.Y(_06972_),
    .A(_06971_));
 sg13g2_a221oi_1 _23594_ (.B2(\top_ihp.oisc.regs[8][2] ),
    .C1(_06972_),
    .B1(_05913_),
    .A1(\top_ihp.oisc.regs[63][2] ),
    .Y(_06973_),
    .A2(_05664_));
 sg13g2_nand4_1 _23595_ (.B(_06967_),
    .C(_06970_),
    .A(_06966_),
    .Y(_06974_),
    .D(_06973_));
 sg13g2_and2_1 _23596_ (.A(\top_ihp.oisc.regs[23][2] ),
    .B(_05825_),
    .X(_06975_));
 sg13g2_a221oi_1 _23597_ (.B2(\top_ihp.oisc.regs[40][2] ),
    .C1(_06975_),
    .B1(net385),
    .A1(\top_ihp.oisc.regs[7][2] ),
    .Y(_06976_),
    .A2(net438));
 sg13g2_a22oi_1 _23598_ (.Y(_06977_),
    .B1(net195),
    .B2(\top_ihp.oisc.regs[58][2] ),
    .A2(net357),
    .A1(\top_ihp.oisc.regs[36][2] ));
 sg13g2_a22oi_1 _23599_ (.Y(_06978_),
    .B1(net202),
    .B2(\top_ihp.oisc.regs[44][2] ),
    .A2(_05923_),
    .A1(\top_ihp.oisc.regs[54][2] ));
 sg13g2_a22oi_1 _23600_ (.Y(_06979_),
    .B1(net405),
    .B2(\top_ihp.oisc.regs[52][2] ),
    .A2(net339),
    .A1(\top_ihp.oisc.regs[38][2] ));
 sg13g2_nand4_1 _23601_ (.B(_06977_),
    .C(_06978_),
    .A(_06976_),
    .Y(_06980_),
    .D(_06979_));
 sg13g2_nor4_1 _23602_ (.A(_06956_),
    .B(_06965_),
    .C(_06974_),
    .D(_06980_),
    .Y(_06981_));
 sg13g2_a22oi_1 _23603_ (.Y(_06982_),
    .B1(net403),
    .B2(\top_ihp.oisc.regs[55][2] ),
    .A2(net347),
    .A1(\top_ihp.oisc.regs[37][2] ));
 sg13g2_a22oi_1 _23604_ (.Y(_06983_),
    .B1(_05719_),
    .B2(\top_ihp.oisc.regs[35][2] ),
    .A2(net416),
    .A1(\top_ihp.oisc.regs[42][2] ));
 sg13g2_a22oi_1 _23605_ (.Y(_06984_),
    .B1(net358),
    .B2(\top_ihp.oisc.regs[47][2] ),
    .A2(_05875_),
    .A1(\top_ihp.oisc.regs[59][2] ));
 sg13g2_a22oi_1 _23606_ (.Y(_06985_),
    .B1(net192),
    .B2(\top_ihp.oisc.regs[62][2] ),
    .A2(net377),
    .A1(\top_ihp.oisc.regs[53][2] ));
 sg13g2_nand4_1 _23607_ (.B(_06983_),
    .C(_06984_),
    .A(_06982_),
    .Y(_06986_),
    .D(_06985_));
 sg13g2_a22oi_1 _23608_ (.Y(_06987_),
    .B1(_05805_),
    .B2(\top_ihp.oisc.regs[56][2] ),
    .A2(_05934_),
    .A1(\top_ihp.oisc.regs[43][2] ));
 sg13g2_a22oi_1 _23609_ (.Y(_06988_),
    .B1(_05726_),
    .B2(\top_ihp.oisc.regs[46][2] ),
    .A2(net188),
    .A1(\top_ihp.oisc.regs[50][2] ));
 sg13g2_a22oi_1 _23610_ (.Y(_06989_),
    .B1(net410),
    .B2(\top_ihp.oisc.regs[41][2] ),
    .A2(_05617_),
    .A1(\top_ihp.oisc.regs[34][2] ));
 sg13g2_a22oi_1 _23611_ (.Y(_06990_),
    .B1(net383),
    .B2(\top_ihp.oisc.regs[60][2] ),
    .A2(net333),
    .A1(\top_ihp.oisc.regs[57][2] ));
 sg13g2_nand4_1 _23612_ (.B(_06988_),
    .C(_06989_),
    .A(_06987_),
    .Y(_06991_),
    .D(_06990_));
 sg13g2_and2_1 _23613_ (.A(\top_ihp.oisc.regs[22][2] ),
    .B(_06146_),
    .X(_06992_));
 sg13g2_a221oi_1 _23614_ (.B2(\top_ihp.oisc.regs[2][2] ),
    .C1(_06992_),
    .B1(_05900_),
    .A1(\top_ihp.oisc.regs[27][2] ),
    .Y(_06993_),
    .A2(net341));
 sg13g2_a22oi_1 _23615_ (.Y(_06994_),
    .B1(_05961_),
    .B2(\top_ihp.oisc.regs[51][2] ),
    .A2(net356),
    .A1(\top_ihp.oisc.regs[31][2] ));
 sg13g2_a22oi_1 _23616_ (.Y(_06995_),
    .B1(net366),
    .B2(\top_ihp.oisc.regs[49][2] ),
    .A2(_05814_),
    .A1(\top_ihp.oisc.regs[33][2] ));
 sg13g2_a22oi_1 _23617_ (.Y(_06996_),
    .B1(_05715_),
    .B2(\top_ihp.oisc.regs[48][2] ),
    .A2(net200),
    .A1(\top_ihp.oisc.regs[61][2] ));
 sg13g2_nand4_1 _23618_ (.B(_06994_),
    .C(_06995_),
    .A(_06993_),
    .Y(_06997_),
    .D(_06996_));
 sg13g2_nor4_2 _23619_ (.A(_05944_),
    .B(_06986_),
    .C(_06991_),
    .Y(_06998_),
    .D(_06997_));
 sg13g2_nand2_1 _23620_ (.Y(_06999_),
    .A(_00206_),
    .B(net59));
 sg13g2_a22oi_1 _23621_ (.Y(_07000_),
    .B1(net26),
    .B2(_06999_),
    .A2(net746),
    .A1(_08090_));
 sg13g2_a21oi_1 _23622_ (.A1(_06981_),
    .A2(_06998_),
    .Y(_00410_),
    .B1(_07000_));
 sg13g2_nand2_1 _23623_ (.Y(_07001_),
    .A(_08307_),
    .B(net801));
 sg13g2_inv_1 _23624_ (.Y(_07002_),
    .A(_00071_));
 sg13g2_o21ai_1 _23625_ (.B1(net27),
    .Y(_07003_),
    .A1(_07002_),
    .A2(net62));
 sg13g2_a22oi_1 _23626_ (.Y(_07004_),
    .B1(net349),
    .B2(\top_ihp.oisc.regs[46][30] ),
    .A2(net379),
    .A1(\top_ihp.oisc.regs[45][30] ));
 sg13g2_a22oi_1 _23627_ (.Y(_07005_),
    .B1(net161),
    .B2(\top_ihp.oisc.regs[44][30] ),
    .A2(net192),
    .A1(\top_ihp.oisc.regs[62][30] ));
 sg13g2_a22oi_1 _23628_ (.Y(_07006_),
    .B1(_05873_),
    .B2(\top_ihp.oisc.regs[34][30] ),
    .A2(_06040_),
    .A1(\top_ihp.oisc.regs[37][30] ));
 sg13g2_a22oi_1 _23629_ (.Y(_07007_),
    .B1(net358),
    .B2(\top_ihp.oisc.regs[47][30] ),
    .A2(_05645_),
    .A1(\top_ihp.oisc.regs[42][30] ));
 sg13g2_nand4_1 _23630_ (.B(_07005_),
    .C(_07006_),
    .A(_07004_),
    .Y(_07008_),
    .D(_07007_));
 sg13g2_a22oi_1 _23631_ (.Y(_07009_),
    .B1(net343),
    .B2(\top_ihp.oisc.regs[18][30] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[22][30] ));
 sg13g2_a22oi_1 _23632_ (.Y(_07010_),
    .B1(net538),
    .B2(\top_ihp.oisc.regs[6][30] ),
    .A2(_05515_),
    .A1(\top_ihp.oisc.regs[14][30] ));
 sg13g2_a22oi_1 _23633_ (.Y(_07011_),
    .B1(net185),
    .B2(\top_ihp.oisc.regs[9][30] ),
    .A2(net664),
    .A1(\top_ihp.oisc.regs[28][30] ));
 sg13g2_a22oi_1 _23634_ (.Y(_07012_),
    .B1(_05501_),
    .B2(\top_ihp.oisc.regs[4][30] ),
    .A2(net438),
    .A1(\top_ihp.oisc.regs[7][30] ));
 sg13g2_nand4_1 _23635_ (.B(_07010_),
    .C(_07011_),
    .A(_07009_),
    .Y(_07013_),
    .D(_07012_));
 sg13g2_a22oi_1 _23636_ (.Y(_07014_),
    .B1(net373),
    .B2(\top_ihp.oisc.regs[1][30] ),
    .A2(net433),
    .A1(\top_ihp.oisc.regs[25][30] ));
 sg13g2_a22oi_1 _23637_ (.Y(_07015_),
    .B1(net183),
    .B2(\top_ihp.oisc.regs[16][30] ),
    .A2(net166),
    .A1(\top_ihp.oisc.regs[3][30] ));
 sg13g2_a22oi_1 _23638_ (.Y(_07016_),
    .B1(net165),
    .B2(\top_ihp.oisc.regs[5][30] ),
    .A2(_05994_),
    .A1(\top_ihp.oisc.regs[11][30] ));
 sg13g2_a22oi_1 _23639_ (.Y(_07017_),
    .B1(net172),
    .B2(\top_ihp.oisc.regs[17][30] ),
    .A2(net335),
    .A1(\top_ihp.oisc.regs[19][30] ));
 sg13g2_nand4_1 _23640_ (.B(_07015_),
    .C(_07016_),
    .A(_07014_),
    .Y(_07018_),
    .D(_07017_));
 sg13g2_a22oi_1 _23641_ (.Y(_07019_),
    .B1(_05453_),
    .B2(\top_ihp.oisc.regs[20][30] ),
    .A2(_05403_),
    .A1(\top_ihp.oisc.regs[26][30] ));
 sg13g2_a22oi_1 _23642_ (.Y(_07020_),
    .B1(net372),
    .B2(\top_ihp.oisc.regs[12][30] ),
    .A2(net370),
    .A1(\top_ihp.oisc.regs[13][30] ));
 sg13g2_a22oi_1 _23643_ (.Y(_07021_),
    .B1(_05571_),
    .B2(\top_ihp.oisc.regs[15][30] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[29][30] ));
 sg13g2_a22oi_1 _23644_ (.Y(_07022_),
    .B1(_05776_),
    .B2(\top_ihp.oisc.regs[24][30] ),
    .A2(_05750_),
    .A1(\top_ihp.oisc.regs[2][30] ));
 sg13g2_a22oi_1 _23645_ (.Y(_07023_),
    .B1(net665),
    .B2(\top_ihp.oisc.regs[8][30] ),
    .A2(net537),
    .A1(\top_ihp.oisc.regs[10][30] ));
 sg13g2_and4_1 _23646_ (.A(_07020_),
    .B(_07021_),
    .C(_07022_),
    .D(_07023_),
    .X(_07024_));
 sg13g2_o21ai_1 _23647_ (.B1(_07024_),
    .Y(_07025_),
    .A1(_05470_),
    .A2(_07019_));
 sg13g2_nor4_1 _23648_ (.A(_07008_),
    .B(_07013_),
    .C(_07018_),
    .D(_07025_),
    .Y(_07026_));
 sg13g2_a22oi_1 _23649_ (.Y(_07027_),
    .B1(net361),
    .B2(\top_ihp.oisc.regs[35][30] ),
    .A2(_05960_),
    .A1(\top_ihp.oisc.regs[31][30] ));
 sg13g2_a22oi_1 _23650_ (.Y(_07028_),
    .B1(_05810_),
    .B2(\top_ihp.oisc.regs[52][30] ),
    .A2(_05648_),
    .A1(\top_ihp.oisc.regs[53][30] ));
 sg13g2_a22oi_1 _23651_ (.Y(_07029_),
    .B1(net403),
    .B2(\top_ihp.oisc.regs[55][30] ),
    .A2(net198),
    .A1(\top_ihp.oisc.regs[59][30] ));
 sg13g2_a22oi_1 _23652_ (.Y(_07030_),
    .B1(net376),
    .B2(\top_ihp.oisc.regs[51][30] ),
    .A2(net414),
    .A1(\top_ihp.oisc.regs[30][30] ));
 sg13g2_nand4_1 _23653_ (.B(_07028_),
    .C(_07029_),
    .A(_07027_),
    .Y(_07031_),
    .D(_07030_));
 sg13g2_a22oi_1 _23654_ (.Y(_07032_),
    .B1(net407),
    .B2(\top_ihp.oisc.regs[33][30] ),
    .A2(net196),
    .A1(\top_ihp.oisc.regs[54][30] ));
 sg13g2_a22oi_1 _23655_ (.Y(_07033_),
    .B1(_05836_),
    .B2(\top_ihp.oisc.regs[61][30] ),
    .A2(net400),
    .A1(\top_ihp.oisc.regs[63][30] ));
 sg13g2_a22oi_1 _23656_ (.Y(_07034_),
    .B1(net194),
    .B2(\top_ihp.oisc.regs[50][30] ),
    .A2(_05641_),
    .A1(\top_ihp.oisc.regs[57][30] ));
 sg13g2_a22oi_1 _23657_ (.Y(_07035_),
    .B1(net719),
    .B2(\top_ihp.oisc.regs[23][30] ),
    .A2(net663),
    .A1(\top_ihp.oisc.regs[21][30] ));
 sg13g2_nand2_1 _23658_ (.Y(_07036_),
    .A(_07001_),
    .B(_07035_));
 sg13g2_a21oi_1 _23659_ (.A1(\top_ihp.oisc.regs[56][30] ),
    .A2(_05804_),
    .Y(_07037_),
    .B1(_07036_));
 sg13g2_nand4_1 _23660_ (.B(_07033_),
    .C(_07034_),
    .A(_07032_),
    .Y(_07038_),
    .D(_07037_));
 sg13g2_a22oi_1 _23661_ (.Y(_07039_),
    .B1(net189),
    .B2(\top_ihp.oisc.regs[60][30] ),
    .A2(net384),
    .A1(\top_ihp.oisc.regs[38][30] ));
 sg13g2_a22oi_1 _23662_ (.Y(_07040_),
    .B1(net195),
    .B2(\top_ihp.oisc.regs[58][30] ),
    .A2(_05711_),
    .A1(\top_ihp.oisc.regs[41][30] ));
 sg13g2_a22oi_1 _23663_ (.Y(_07041_),
    .B1(_05932_),
    .B2(\top_ihp.oisc.regs[32][30] ),
    .A2(net357),
    .A1(\top_ihp.oisc.regs[36][30] ));
 sg13g2_a22oi_1 _23664_ (.Y(_07042_),
    .B1(_05966_),
    .B2(\top_ihp.oisc.regs[39][30] ),
    .A2(net362),
    .A1(\top_ihp.oisc.regs[43][30] ));
 sg13g2_nand4_1 _23665_ (.B(_07040_),
    .C(_07041_),
    .A(_07039_),
    .Y(_07043_),
    .D(_07042_));
 sg13g2_a22oi_1 _23666_ (.Y(_07044_),
    .B1(_05841_),
    .B2(\top_ihp.oisc.regs[49][30] ),
    .A2(_05715_),
    .A1(\top_ihp.oisc.regs[48][30] ));
 sg13g2_a22oi_1 _23667_ (.Y(_07045_),
    .B1(_05609_),
    .B2(\top_ihp.oisc.regs[27][30] ),
    .A2(_05843_),
    .A1(\top_ihp.oisc.regs[40][30] ));
 sg13g2_nand3_1 _23668_ (.B(_07044_),
    .C(_07045_),
    .A(_05742_),
    .Y(_07046_));
 sg13g2_nor4_2 _23669_ (.A(_07031_),
    .B(_07038_),
    .C(_07043_),
    .Y(_07047_),
    .D(_07046_));
 sg13g2_a22oi_1 _23670_ (.Y(_00411_),
    .B1(_07026_),
    .B2(_07047_),
    .A2(_07003_),
    .A1(_07001_));
 sg13g2_nand2_1 _23671_ (.Y(_07048_),
    .A(\top_ihp.oisc.regs[32][31] ),
    .B(net363));
 sg13g2_a22oi_1 _23672_ (.Y(_07049_),
    .B1(net408),
    .B2(\top_ihp.oisc.regs[35][31] ),
    .A2(net413),
    .A1(\top_ihp.oisc.regs[63][31] ));
 sg13g2_a22oi_1 _23673_ (.Y(_07050_),
    .B1(net362),
    .B2(\top_ihp.oisc.regs[43][31] ),
    .A2(net351),
    .A1(\top_ihp.oisc.regs[40][31] ));
 sg13g2_a22oi_1 _23674_ (.Y(_07051_),
    .B1(net364),
    .B2(\top_ihp.oisc.regs[52][31] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[39][31] ));
 sg13g2_nand4_1 _23675_ (.B(_07049_),
    .C(_07050_),
    .A(_07048_),
    .Y(_07052_),
    .D(_07051_));
 sg13g2_a22oi_1 _23676_ (.Y(_07053_),
    .B1(_05870_),
    .B2(\top_ihp.oisc.regs[51][31] ),
    .A2(net358),
    .A1(\top_ihp.oisc.regs[47][31] ));
 sg13g2_a22oi_1 _23677_ (.Y(_07054_),
    .B1(_05937_),
    .B2(\top_ihp.oisc.regs[33][31] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[53][31] ));
 sg13g2_nand3_1 _23678_ (.B(_07053_),
    .C(_07054_),
    .A(_05918_),
    .Y(_07055_));
 sg13g2_a22oi_1 _23679_ (.Y(_07056_),
    .B1(_05596_),
    .B2(\top_ihp.oisc.regs[37][31] ),
    .A2(net199),
    .A1(\top_ihp.oisc.regs[50][31] ));
 sg13g2_nand2_1 _23680_ (.Y(_07057_),
    .A(_09497_),
    .B(net835));
 sg13g2_a22oi_1 _23681_ (.Y(_07058_),
    .B1(_05824_),
    .B2(\top_ihp.oisc.regs[23][31] ),
    .A2(_05820_),
    .A1(\top_ihp.oisc.regs[21][31] ));
 sg13g2_nand2_1 _23682_ (.Y(_07059_),
    .A(_07057_),
    .B(_07058_));
 sg13g2_a221oi_1 _23683_ (.B2(\top_ihp.oisc.regs[13][31] ),
    .C1(_07059_),
    .B1(_05828_),
    .A1(\top_ihp.oisc.regs[7][31] ),
    .Y(_07060_),
    .A2(net554));
 sg13g2_a22oi_1 _23684_ (.Y(_07061_),
    .B1(_05711_),
    .B2(\top_ihp.oisc.regs[41][31] ),
    .A2(_05654_),
    .A1(\top_ihp.oisc.regs[56][31] ));
 sg13g2_a22oi_1 _23685_ (.Y(_07062_),
    .B1(net339),
    .B2(\top_ihp.oisc.regs[38][31] ),
    .A2(net186),
    .A1(\top_ihp.oisc.regs[59][31] ));
 sg13g2_nand4_1 _23686_ (.B(_07060_),
    .C(_07061_),
    .A(_07056_),
    .Y(_07063_),
    .D(_07062_));
 sg13g2_a22oi_1 _23687_ (.Y(_07064_),
    .B1(net190),
    .B2(\top_ihp.oisc.regs[61][31] ),
    .A2(net357),
    .A1(\top_ihp.oisc.regs[36][31] ));
 sg13g2_a22oi_1 _23688_ (.Y(_07065_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[27][31] ),
    .A2(_05802_),
    .A1(\top_ihp.oisc.regs[45][31] ));
 sg13g2_a22oi_1 _23689_ (.Y(_07066_),
    .B1(_05736_),
    .B2(\top_ihp.oisc.regs[55][31] ),
    .A2(_05923_),
    .A1(\top_ihp.oisc.regs[54][31] ));
 sg13g2_a22oi_1 _23690_ (.Y(_07067_),
    .B1(_05919_),
    .B2(\top_ihp.oisc.regs[49][31] ),
    .A2(net346),
    .A1(\top_ihp.oisc.regs[30][31] ));
 sg13g2_nand4_1 _23691_ (.B(_07065_),
    .C(_07066_),
    .A(_07064_),
    .Y(_07068_),
    .D(_07067_));
 sg13g2_nor4_2 _23692_ (.A(_07052_),
    .B(_07055_),
    .C(_07063_),
    .Y(_07069_),
    .D(_07068_));
 sg13g2_a22oi_1 _23693_ (.Y(_07070_),
    .B1(net399),
    .B2(\top_ihp.oisc.regs[58][31] ),
    .A2(_06637_),
    .A1(\top_ihp.oisc.regs[44][31] ));
 sg13g2_a22oi_1 _23694_ (.Y(_07071_),
    .B1(net383),
    .B2(\top_ihp.oisc.regs[60][31] ),
    .A2(net174),
    .A1(\top_ihp.oisc.regs[62][31] ));
 sg13g2_a22oi_1 _23695_ (.Y(_07072_),
    .B1(net406),
    .B2(\top_ihp.oisc.regs[46][31] ),
    .A2(net333),
    .A1(\top_ihp.oisc.regs[57][31] ));
 sg13g2_a22oi_1 _23696_ (.Y(_07073_),
    .B1(net409),
    .B2(\top_ihp.oisc.regs[48][31] ),
    .A2(_05644_),
    .A1(\top_ihp.oisc.regs[42][31] ));
 sg13g2_nand4_1 _23697_ (.B(_07071_),
    .C(_07072_),
    .A(_07070_),
    .Y(_07074_),
    .D(_07073_));
 sg13g2_a22oi_1 _23698_ (.Y(_07075_),
    .B1(net537),
    .B2(\top_ihp.oisc.regs[10][31] ),
    .A2(_05776_),
    .A1(\top_ihp.oisc.regs[24][31] ));
 sg13g2_a22oi_1 _23699_ (.Y(_07076_),
    .B1(net372),
    .B2(\top_ihp.oisc.regs[12][31] ),
    .A2(net551),
    .A1(\top_ihp.oisc.regs[25][31] ));
 sg13g2_a22oi_1 _23700_ (.Y(_07077_),
    .B1(net665),
    .B2(\top_ihp.oisc.regs[8][31] ),
    .A2(net432),
    .A1(\top_ihp.oisc.regs[4][31] ));
 sg13g2_a22oi_1 _23701_ (.Y(_07078_),
    .B1(net380),
    .B2(\top_ihp.oisc.regs[11][31] ),
    .A2(net552),
    .A1(\top_ihp.oisc.regs[20][31] ));
 sg13g2_nand4_1 _23702_ (.B(_07076_),
    .C(_07077_),
    .A(_07075_),
    .Y(_07079_),
    .D(_07078_));
 sg13g2_a22oi_1 _23703_ (.Y(_07080_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[34][31] ),
    .A2(net356),
    .A1(\top_ihp.oisc.regs[31][31] ));
 sg13g2_nand2b_1 _23704_ (.Y(_07081_),
    .B(_07080_),
    .A_N(_07079_));
 sg13g2_a22oi_1 _23705_ (.Y(_07082_),
    .B1(net165),
    .B2(\top_ihp.oisc.regs[5][31] ),
    .A2(_05507_),
    .A1(\top_ihp.oisc.regs[1][31] ));
 sg13g2_a22oi_1 _23706_ (.Y(_07083_),
    .B1(net172),
    .B2(\top_ihp.oisc.regs[17][31] ),
    .A2(net534),
    .A1(\top_ihp.oisc.regs[18][31] ));
 sg13g2_a22oi_1 _23707_ (.Y(_07084_),
    .B1(net185),
    .B2(\top_ihp.oisc.regs[9][31] ),
    .A2(net664),
    .A1(\top_ihp.oisc.regs[28][31] ));
 sg13g2_a22oi_1 _23708_ (.Y(_07085_),
    .B1(net335),
    .B2(\top_ihp.oisc.regs[19][31] ),
    .A2(net546),
    .A1(\top_ihp.oisc.regs[14][31] ));
 sg13g2_nand4_1 _23709_ (.B(_07083_),
    .C(_07084_),
    .A(_07082_),
    .Y(_07086_),
    .D(_07085_));
 sg13g2_a22oi_1 _23710_ (.Y(_07087_),
    .B1(net538),
    .B2(\top_ihp.oisc.regs[6][31] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[22][31] ));
 sg13g2_a22oi_1 _23711_ (.Y(_07088_),
    .B1(net166),
    .B2(\top_ihp.oisc.regs[3][31] ),
    .A2(_05895_),
    .A1(\top_ihp.oisc.regs[29][31] ));
 sg13g2_a22oi_1 _23712_ (.Y(_07089_),
    .B1(net183),
    .B2(\top_ihp.oisc.regs[16][31] ),
    .A2(net369),
    .A1(\top_ihp.oisc.regs[2][31] ));
 sg13g2_a22oi_1 _23713_ (.Y(_07090_),
    .B1(net168),
    .B2(\top_ihp.oisc.regs[26][31] ),
    .A2(net162),
    .A1(\top_ihp.oisc.regs[15][31] ));
 sg13g2_nand4_1 _23714_ (.B(_07088_),
    .C(_07089_),
    .A(_07087_),
    .Y(_07091_),
    .D(_07090_));
 sg13g2_nor4_1 _23715_ (.A(_07074_),
    .B(_07081_),
    .C(_07086_),
    .D(_07091_),
    .Y(_07092_));
 sg13g2_a21o_1 _23716_ (.A2(net63),
    .A1(_00072_),
    .B1(net58),
    .X(_07093_));
 sg13g2_a22oi_1 _23717_ (.Y(_00412_),
    .B1(_07093_),
    .B2(_07057_),
    .A2(_07092_),
    .A1(_07069_));
 sg13g2_and2_1 _23718_ (.A(_08086_),
    .B(net803),
    .X(_07094_));
 sg13g2_a221oi_1 _23719_ (.B2(\top_ihp.oisc.regs[23][3] ),
    .C1(_07094_),
    .B1(net720),
    .A1(\top_ihp.oisc.regs[21][3] ),
    .Y(_07095_),
    .A2(net666));
 sg13g2_a22oi_1 _23720_ (.Y(_07096_),
    .B1(net165),
    .B2(\top_ihp.oisc.regs[5][3] ),
    .A2(_06156_),
    .A1(\top_ihp.oisc.regs[4][3] ));
 sg13g2_a22oi_1 _23721_ (.Y(_07097_),
    .B1(net164),
    .B2(\top_ihp.oisc.regs[9][3] ),
    .A2(net390),
    .A1(\top_ihp.oisc.regs[13][3] ));
 sg13g2_a22oi_1 _23722_ (.Y(_07098_),
    .B1(net162),
    .B2(\top_ihp.oisc.regs[15][3] ),
    .A2(_06059_),
    .A1(\top_ihp.oisc.regs[3][3] ));
 sg13g2_nand4_1 _23723_ (.B(_07096_),
    .C(_07097_),
    .A(_07095_),
    .Y(_07099_),
    .D(_07098_));
 sg13g2_a22oi_1 _23724_ (.Y(_07100_),
    .B1(net167),
    .B2(\top_ihp.oisc.regs[24][3] ),
    .A2(net184),
    .A1(\top_ihp.oisc.regs[12][3] ));
 sg13g2_a22oi_1 _23725_ (.Y(_07101_),
    .B1(_05887_),
    .B2(\top_ihp.oisc.regs[1][3] ),
    .A2(net540),
    .A1(\top_ihp.oisc.regs[20][3] ));
 sg13g2_mux2_1 _23726_ (.A0(\top_ihp.oisc.regs[6][3] ),
    .A1(\top_ihp.oisc.regs[2][3] ),
    .S(net541),
    .X(_07102_));
 sg13g2_a22oi_1 _23727_ (.Y(_07103_),
    .B1(_05748_),
    .B2(_07102_),
    .A2(net664),
    .A1(\top_ihp.oisc.regs[28][3] ));
 sg13g2_a22oi_1 _23728_ (.Y(_07104_),
    .B1(net160),
    .B2(\top_ihp.oisc.regs[17][3] ),
    .A2(net438),
    .A1(\top_ihp.oisc.regs[7][3] ));
 sg13g2_nand4_1 _23729_ (.B(_07101_),
    .C(_07103_),
    .A(_07100_),
    .Y(_07105_),
    .D(_07104_));
 sg13g2_a22oi_1 _23730_ (.Y(_07106_),
    .B1(_05905_),
    .B2(\top_ihp.oisc.regs[10][3] ),
    .A2(net546),
    .A1(\top_ihp.oisc.regs[14][3] ));
 sg13g2_a22oi_1 _23731_ (.Y(_07107_),
    .B1(_05765_),
    .B2(\top_ihp.oisc.regs[26][3] ),
    .A2(net544),
    .A1(\top_ihp.oisc.regs[18][3] ));
 sg13g2_a22oi_1 _23732_ (.Y(_07108_),
    .B1(net371),
    .B2(\top_ihp.oisc.regs[16][3] ),
    .A2(net543),
    .A1(\top_ihp.oisc.regs[19][3] ));
 sg13g2_a22oi_1 _23733_ (.Y(_07109_),
    .B1(net665),
    .B2(\top_ihp.oisc.regs[8][3] ),
    .A2(_05529_),
    .A1(\top_ihp.oisc.regs[29][3] ));
 sg13g2_and4_1 _23734_ (.A(_07106_),
    .B(_07107_),
    .C(_07108_),
    .D(_07109_),
    .X(_07110_));
 sg13g2_a22oi_1 _23735_ (.Y(_07111_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[34][3] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[53][3] ));
 sg13g2_nand2_1 _23736_ (.Y(_07112_),
    .A(\top_ihp.oisc.regs[11][3] ),
    .B(net169));
 sg13g2_a22oi_1 _23737_ (.Y(_07113_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[25][3] ),
    .A2(net533),
    .A1(\top_ihp.oisc.regs[22][3] ));
 sg13g2_nand4_1 _23738_ (.B(_07111_),
    .C(_07112_),
    .A(_07110_),
    .Y(_07114_),
    .D(_07113_));
 sg13g2_a22oi_1 _23739_ (.Y(_07115_),
    .B1(net396),
    .B2(\top_ihp.oisc.regs[46][3] ),
    .A2(net426),
    .A1(\top_ihp.oisc.regs[37][3] ));
 sg13g2_a22oi_1 _23740_ (.Y(_07116_),
    .B1(net195),
    .B2(\top_ihp.oisc.regs[58][3] ),
    .A2(net363),
    .A1(\top_ihp.oisc.regs[32][3] ));
 sg13g2_a22oi_1 _23741_ (.Y(_07117_),
    .B1(_05793_),
    .B2(\top_ihp.oisc.regs[55][3] ),
    .A2(net387),
    .A1(\top_ihp.oisc.regs[47][3] ));
 sg13g2_a22oi_1 _23742_ (.Y(_07118_),
    .B1(net202),
    .B2(\top_ihp.oisc.regs[44][3] ),
    .A2(net357),
    .A1(\top_ihp.oisc.regs[36][3] ));
 sg13g2_nand4_1 _23743_ (.B(_07116_),
    .C(_07117_),
    .A(_07115_),
    .Y(_07119_),
    .D(_07118_));
 sg13g2_nor4_1 _23744_ (.A(_07099_),
    .B(_07105_),
    .C(_07114_),
    .D(_07119_),
    .Y(_07120_));
 sg13g2_a22oi_1 _23745_ (.Y(_07121_),
    .B1(_05787_),
    .B2(\top_ihp.oisc.regs[54][3] ),
    .A2(_05636_),
    .A1(\top_ihp.oisc.regs[40][3] ));
 sg13g2_a22oi_1 _23746_ (.Y(_07122_),
    .B1(net362),
    .B2(\top_ihp.oisc.regs[43][3] ),
    .A2(_05660_),
    .A1(\top_ihp.oisc.regs[30][3] ));
 sg13g2_a22oi_1 _23747_ (.Y(_07123_),
    .B1(net364),
    .B2(\top_ihp.oisc.regs[52][3] ),
    .A2(net378),
    .A1(\top_ihp.oisc.regs[38][3] ));
 sg13g2_a22oi_1 _23748_ (.Y(_07124_),
    .B1(_05681_),
    .B2(\top_ihp.oisc.regs[45][3] ),
    .A2(net188),
    .A1(\top_ihp.oisc.regs[50][3] ));
 sg13g2_nand4_1 _23749_ (.B(_07122_),
    .C(_07123_),
    .A(_07121_),
    .Y(_07125_),
    .D(_07124_));
 sg13g2_a22oi_1 _23750_ (.Y(_07126_),
    .B1(net395),
    .B2(\top_ihp.oisc.regs[41][3] ),
    .A2(net191),
    .A1(\top_ihp.oisc.regs[59][3] ));
 sg13g2_a22oi_1 _23751_ (.Y(_07127_),
    .B1(net382),
    .B2(\top_ihp.oisc.regs[27][3] ),
    .A2(_05812_),
    .A1(\top_ihp.oisc.regs[62][3] ));
 sg13g2_a22oi_1 _23752_ (.Y(_07128_),
    .B1(net171),
    .B2(\top_ihp.oisc.regs[60][3] ),
    .A2(_06310_),
    .A1(\top_ihp.oisc.regs[57][3] ));
 sg13g2_nand2_1 _23753_ (.Y(_07129_),
    .A(_05492_),
    .B(net673));
 sg13g2_a22oi_1 _23754_ (.Y(_07130_),
    .B1(_05586_),
    .B2(\top_ihp.oisc.regs[56][3] ),
    .A2(_05582_),
    .A1(\top_ihp.oisc.regs[48][3] ));
 sg13g2_nor2_1 _23755_ (.A(_07129_),
    .B(_07130_),
    .Y(_07131_));
 sg13g2_a21oi_1 _23756_ (.A1(\top_ihp.oisc.regs[61][3] ),
    .A2(_05674_),
    .Y(_07132_),
    .B1(_07131_));
 sg13g2_nand4_1 _23757_ (.B(_07127_),
    .C(_07128_),
    .A(_07126_),
    .Y(_07133_),
    .D(_07132_));
 sg13g2_a22oi_1 _23758_ (.Y(_07134_),
    .B1(net361),
    .B2(\top_ihp.oisc.regs[35][3] ),
    .A2(net354),
    .A1(\top_ihp.oisc.regs[39][3] ));
 sg13g2_a22oi_1 _23759_ (.Y(_07135_),
    .B1(_06172_),
    .B2(\top_ihp.oisc.regs[42][3] ),
    .A2(net356),
    .A1(\top_ihp.oisc.regs[31][3] ));
 sg13g2_a22oi_1 _23760_ (.Y(_07136_),
    .B1(_05919_),
    .B2(\top_ihp.oisc.regs[49][3] ),
    .A2(_05783_),
    .A1(\top_ihp.oisc.regs[63][3] ));
 sg13g2_a22oi_1 _23761_ (.Y(_07137_),
    .B1(_05722_),
    .B2(\top_ihp.oisc.regs[33][3] ),
    .A2(net420),
    .A1(\top_ihp.oisc.regs[51][3] ));
 sg13g2_nand4_1 _23762_ (.B(_07135_),
    .C(_07136_),
    .A(_07134_),
    .Y(_07138_),
    .D(_07137_));
 sg13g2_nor4_2 _23763_ (.A(net60),
    .B(_07125_),
    .C(_07133_),
    .Y(_07139_),
    .D(_07138_));
 sg13g2_a21oi_1 _23764_ (.A1(_00207_),
    .A2(_05707_),
    .Y(_07140_),
    .B1(_05744_));
 sg13g2_nor2_1 _23765_ (.A(_07094_),
    .B(_07140_),
    .Y(_07141_));
 sg13g2_a21oi_1 _23766_ (.A1(_07120_),
    .A2(_07139_),
    .Y(_00413_),
    .B1(_07141_));
 sg13g2_a22oi_1 _23767_ (.Y(_07142_),
    .B1(net360),
    .B2(\top_ihp.oisc.regs[33][4] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[39][4] ));
 sg13g2_a22oi_1 _23768_ (.Y(_07143_),
    .B1(_06052_),
    .B2(\top_ihp.oisc.regs[53][4] ),
    .A2(net351),
    .A1(\top_ihp.oisc.regs[40][4] ));
 sg13g2_a22oi_1 _23769_ (.Y(_07144_),
    .B1(net379),
    .B2(\top_ihp.oisc.regs[45][4] ),
    .A2(net201),
    .A1(\top_ihp.oisc.regs[54][4] ));
 sg13g2_a22oi_1 _23770_ (.Y(_07145_),
    .B1(net198),
    .B2(\top_ihp.oisc.regs[59][4] ),
    .A2(net352),
    .A1(\top_ihp.oisc.regs[43][4] ));
 sg13g2_nand4_1 _23771_ (.B(_07143_),
    .C(_07144_),
    .A(_07142_),
    .Y(_07146_),
    .D(_07145_));
 sg13g2_a22oi_1 _23772_ (.Y(_07147_),
    .B1(net665),
    .B2(\top_ihp.oisc.regs[8][4] ),
    .A2(net401),
    .A1(\top_ihp.oisc.regs[3][4] ));
 sg13g2_a22oi_1 _23773_ (.Y(_07148_),
    .B1(net668),
    .B2(\top_ihp.oisc.regs[28][4] ),
    .A2(_05514_),
    .A1(\top_ihp.oisc.regs[14][4] ));
 sg13g2_and4_1 _23774_ (.A(\top_ihp.oisc.regs[34][4] ),
    .B(net723),
    .C(_05667_),
    .D(net728),
    .X(_07149_));
 sg13g2_a21oi_1 _23775_ (.A1(\top_ihp.oisc.regs[16][4] ),
    .A2(_05759_),
    .Y(_07150_),
    .B1(_07149_));
 sg13g2_a22oi_1 _23776_ (.Y(_07151_),
    .B1(_05765_),
    .B2(\top_ihp.oisc.regs[26][4] ),
    .A2(_05505_),
    .A1(\top_ihp.oisc.regs[1][4] ));
 sg13g2_and4_1 _23777_ (.A(_07147_),
    .B(_07148_),
    .C(_07150_),
    .D(_07151_),
    .X(_07152_));
 sg13g2_a22oi_1 _23778_ (.Y(_07153_),
    .B1(_06115_),
    .B2(\top_ihp.oisc.regs[5][4] ),
    .A2(net534),
    .A1(\top_ihp.oisc.regs[18][4] ));
 sg13g2_a22oi_1 _23779_ (.Y(_07154_),
    .B1(_05885_),
    .B2(\top_ihp.oisc.regs[6][4] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[22][4] ));
 sg13g2_nand3_1 _23780_ (.B(_07153_),
    .C(_07154_),
    .A(_07152_),
    .Y(_07155_));
 sg13g2_and2_1 _23781_ (.A(_08109_),
    .B(net803),
    .X(_07156_));
 sg13g2_a221oi_1 _23782_ (.B2(\top_ihp.oisc.regs[23][4] ),
    .C1(_07156_),
    .B1(net720),
    .A1(\top_ihp.oisc.regs[24][4] ),
    .Y(_07157_),
    .A2(net402));
 sg13g2_nand2_1 _23783_ (.Y(_07158_),
    .A(\top_ihp.oisc.regs[21][4] ),
    .B(net666));
 sg13g2_nand3_1 _23784_ (.B(_05667_),
    .C(net749),
    .A(\top_ihp.oisc.regs[2][4] ),
    .Y(_07159_));
 sg13g2_nand4_1 _23785_ (.B(net729),
    .C(net662),
    .A(\top_ihp.oisc.regs[20][4] ),
    .Y(_07160_),
    .D(_05433_));
 sg13g2_and3_1 _23786_ (.X(_07161_),
    .A(_07158_),
    .B(_07159_),
    .C(_07160_));
 sg13g2_a22oi_1 _23787_ (.Y(_07162_),
    .B1(_05994_),
    .B2(\top_ihp.oisc.regs[11][4] ),
    .A2(net203),
    .A1(\top_ihp.oisc.regs[29][4] ));
 sg13g2_a22oi_1 _23788_ (.Y(_07163_),
    .B1(net180),
    .B2(\top_ihp.oisc.regs[13][4] ),
    .A2(net163),
    .A1(\top_ihp.oisc.regs[4][4] ));
 sg13g2_nand4_1 _23789_ (.B(_07161_),
    .C(_07162_),
    .A(_07157_),
    .Y(_07164_),
    .D(_07163_));
 sg13g2_a22oi_1 _23790_ (.Y(_07165_),
    .B1(_05889_),
    .B2(\top_ihp.oisc.regs[12][4] ),
    .A2(_06002_),
    .A1(\top_ihp.oisc.regs[19][4] ));
 sg13g2_a22oi_1 _23791_ (.Y(_07166_),
    .B1(net172),
    .B2(\top_ihp.oisc.regs[17][4] ),
    .A2(_05884_),
    .A1(\top_ihp.oisc.regs[9][4] ));
 sg13g2_a22oi_1 _23792_ (.Y(_07167_),
    .B1(net334),
    .B2(\top_ihp.oisc.regs[10][4] ),
    .A2(_05896_),
    .A1(\top_ihp.oisc.regs[15][4] ));
 sg13g2_a22oi_1 _23793_ (.Y(_07168_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[25][4] ),
    .A2(_06065_),
    .A1(\top_ihp.oisc.regs[7][4] ));
 sg13g2_nand4_1 _23794_ (.B(_07166_),
    .C(_07167_),
    .A(_07165_),
    .Y(_07169_),
    .D(_07168_));
 sg13g2_nor4_1 _23795_ (.A(_07146_),
    .B(_07155_),
    .C(_07164_),
    .D(_07169_),
    .Y(_07170_));
 sg13g2_a22oi_1 _23796_ (.Y(_07171_),
    .B1(net382),
    .B2(\top_ihp.oisc.regs[27][4] ),
    .A2(net375),
    .A1(\top_ihp.oisc.regs[36][4] ));
 sg13g2_a22oi_1 _23797_ (.Y(_07172_),
    .B1(_05593_),
    .B2(\top_ihp.oisc.regs[47][4] ),
    .A2(_05452_),
    .A1(\top_ihp.oisc.regs[46][4] ));
 sg13g2_inv_1 _23798_ (.Y(_07173_),
    .A(_07172_));
 sg13g2_a22oi_1 _23799_ (.Y(_07174_),
    .B1(_07173_),
    .B2(_05458_),
    .A2(_05588_),
    .A1(\top_ihp.oisc.regs[60][4] ));
 sg13g2_a22oi_1 _23800_ (.Y(_07175_),
    .B1(net338),
    .B2(\top_ihp.oisc.regs[32][4] ),
    .A2(_05673_),
    .A1(\top_ihp.oisc.regs[61][4] ));
 sg13g2_nand3_1 _23801_ (.B(_05488_),
    .C(_05469_),
    .A(\top_ihp.oisc.regs[62][4] ),
    .Y(_07176_));
 sg13g2_nand3_1 _23802_ (.B(_05491_),
    .C(net723),
    .A(\top_ihp.oisc.regs[50][4] ),
    .Y(_07177_));
 sg13g2_a21oi_1 _23803_ (.A1(_07176_),
    .A2(_07177_),
    .Y(_07178_),
    .B1(_06097_));
 sg13g2_a21oi_1 _23804_ (.A1(\top_ihp.oisc.regs[44][4] ),
    .A2(_06637_),
    .Y(_07179_),
    .B1(_07178_));
 sg13g2_nand4_1 _23805_ (.B(_07174_),
    .C(_07175_),
    .A(_07171_),
    .Y(_07180_),
    .D(_07179_));
 sg13g2_a22oi_1 _23806_ (.Y(_07181_),
    .B1(net361),
    .B2(\top_ihp.oisc.regs[35][4] ),
    .A2(net397),
    .A1(\top_ihp.oisc.regs[37][4] ));
 sg13g2_a22oi_1 _23807_ (.Y(_07182_),
    .B1(net339),
    .B2(\top_ihp.oisc.regs[38][4] ),
    .A2(net400),
    .A1(\top_ihp.oisc.regs[63][4] ));
 sg13g2_a22oi_1 _23808_ (.Y(_07183_),
    .B1(net366),
    .B2(\top_ihp.oisc.regs[49][4] ),
    .A2(_06310_),
    .A1(\top_ihp.oisc.regs[57][4] ));
 sg13g2_a22oi_1 _23809_ (.Y(_07184_),
    .B1(net359),
    .B2(\top_ihp.oisc.regs[55][4] ),
    .A2(net409),
    .A1(\top_ihp.oisc.regs[48][4] ));
 sg13g2_nand4_1 _23810_ (.B(_07182_),
    .C(_07183_),
    .A(_07181_),
    .Y(_07185_),
    .D(_07184_));
 sg13g2_a22oi_1 _23811_ (.Y(_07186_),
    .B1(_05729_),
    .B2(\top_ihp.oisc.regs[52][4] ),
    .A2(net410),
    .A1(\top_ihp.oisc.regs[41][4] ));
 sg13g2_a22oi_1 _23812_ (.Y(_07187_),
    .B1(net195),
    .B2(\top_ihp.oisc.regs[58][4] ),
    .A2(_05870_),
    .A1(\top_ihp.oisc.regs[51][4] ));
 sg13g2_a22oi_1 _23813_ (.Y(_07188_),
    .B1(_05835_),
    .B2(\top_ihp.oisc.regs[30][4] ),
    .A2(net336),
    .A1(\top_ihp.oisc.regs[42][4] ));
 sg13g2_a22oi_1 _23814_ (.Y(_07189_),
    .B1(_05654_),
    .B2(\top_ihp.oisc.regs[56][4] ),
    .A2(_05461_),
    .A1(\top_ihp.oisc.regs[31][4] ));
 sg13g2_nand4_1 _23815_ (.B(_07187_),
    .C(_07188_),
    .A(_07186_),
    .Y(_07190_),
    .D(_07189_));
 sg13g2_nor4_2 _23816_ (.A(net60),
    .B(_07180_),
    .C(_07185_),
    .Y(_07191_),
    .D(_07190_));
 sg13g2_a21oi_1 _23817_ (.A1(_00208_),
    .A2(_05707_),
    .Y(_07192_),
    .B1(_05744_));
 sg13g2_nor2_1 _23818_ (.A(_07156_),
    .B(_07192_),
    .Y(_07193_));
 sg13g2_a21oi_1 _23819_ (.A1(_07170_),
    .A2(_07191_),
    .Y(_00414_),
    .B1(_07193_));
 sg13g2_a22oi_1 _23820_ (.Y(_07194_),
    .B1(_05927_),
    .B2(\top_ihp.oisc.regs[63][5] ),
    .A2(_05652_),
    .A1(\top_ihp.oisc.regs[54][5] ));
 sg13g2_a22oi_1 _23821_ (.Y(_07195_),
    .B1(net171),
    .B2(\top_ihp.oisc.regs[60][5] ),
    .A2(net364),
    .A1(\top_ihp.oisc.regs[52][5] ));
 sg13g2_a22oi_1 _23822_ (.Y(_07196_),
    .B1(net382),
    .B2(\top_ihp.oisc.regs[27][5] ),
    .A2(_05660_),
    .A1(\top_ihp.oisc.regs[30][5] ));
 sg13g2_a22oi_1 _23823_ (.Y(_07197_),
    .B1(net539),
    .B2(\top_ihp.oisc.regs[34][5] ),
    .A2(_05981_),
    .A1(\top_ihp.oisc.regs[43][5] ));
 sg13g2_nand4_1 _23824_ (.B(_07195_),
    .C(_07196_),
    .A(_07194_),
    .Y(_07198_),
    .D(_07197_));
 sg13g2_a22oi_1 _23825_ (.Y(_07199_),
    .B1(net161),
    .B2(\top_ihp.oisc.regs[44][5] ),
    .A2(_05626_),
    .A1(\top_ihp.oisc.regs[51][5] ));
 sg13g2_a22oi_1 _23826_ (.Y(_07200_),
    .B1(net387),
    .B2(\top_ihp.oisc.regs[47][5] ),
    .A2(_05809_),
    .A1(\top_ihp.oisc.regs[42][5] ));
 sg13g2_a22oi_1 _23827_ (.Y(_07201_),
    .B1(net187),
    .B2(\top_ihp.oisc.regs[56][5] ),
    .A2(net347),
    .A1(\top_ihp.oisc.regs[37][5] ));
 sg13g2_a22oi_1 _23828_ (.Y(_07202_),
    .B1(_05833_),
    .B2(\top_ihp.oisc.regs[59][5] ),
    .A2(_05830_),
    .A1(\top_ihp.oisc.regs[31][5] ));
 sg13g2_nand4_1 _23829_ (.B(_07200_),
    .C(_07201_),
    .A(_07199_),
    .Y(_07203_),
    .D(_07202_));
 sg13g2_nand2_1 _23830_ (.Y(_07204_),
    .A(\top_ihp.oisc.regs[58][5] ),
    .B(_05791_));
 sg13g2_a22oi_1 _23831_ (.Y(_07205_),
    .B1(net354),
    .B2(\top_ihp.oisc.regs[39][5] ),
    .A2(net339),
    .A1(\top_ihp.oisc.regs[38][5] ));
 sg13g2_nand3_1 _23832_ (.B(_07204_),
    .C(_07205_),
    .A(_06017_),
    .Y(_07206_));
 sg13g2_a22oi_1 _23833_ (.Y(_07207_),
    .B1(net361),
    .B2(\top_ihp.oisc.regs[35][5] ),
    .A2(_06052_),
    .A1(\top_ihp.oisc.regs[53][5] ));
 sg13g2_a22oi_1 _23834_ (.Y(_07208_),
    .B1(_05932_),
    .B2(\top_ihp.oisc.regs[32][5] ),
    .A2(net385),
    .A1(\top_ihp.oisc.regs[40][5] ));
 sg13g2_a22oi_1 _23835_ (.Y(_07209_),
    .B1(net194),
    .B2(\top_ihp.oisc.regs[50][5] ),
    .A2(net176),
    .A1(\top_ihp.oisc.regs[62][5] ));
 sg13g2_a22oi_1 _23836_ (.Y(_07210_),
    .B1(net396),
    .B2(\top_ihp.oisc.regs[46][5] ),
    .A2(_05641_),
    .A1(\top_ihp.oisc.regs[57][5] ));
 sg13g2_nand4_1 _23837_ (.B(_07208_),
    .C(_07209_),
    .A(_07207_),
    .Y(_07211_),
    .D(_07210_));
 sg13g2_nor4_2 _23838_ (.A(_07198_),
    .B(_07203_),
    .C(_07206_),
    .Y(_07212_),
    .D(_07211_));
 sg13g2_a22oi_1 _23839_ (.Y(_07213_),
    .B1(net381),
    .B2(\top_ihp.oisc.regs[48][5] ),
    .A2(_05674_),
    .A1(\top_ihp.oisc.regs[61][5] ));
 sg13g2_a22oi_1 _23840_ (.Y(_07214_),
    .B1(net359),
    .B2(\top_ihp.oisc.regs[55][5] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[36][5] ));
 sg13g2_a22oi_1 _23841_ (.Y(_07215_),
    .B1(net404),
    .B2(\top_ihp.oisc.regs[49][5] ),
    .A2(_05721_),
    .A1(\top_ihp.oisc.regs[33][5] ));
 sg13g2_a22oi_1 _23842_ (.Y(_07216_),
    .B1(net340),
    .B2(\top_ihp.oisc.regs[41][5] ),
    .A2(_05680_),
    .A1(\top_ihp.oisc.regs[45][5] ));
 sg13g2_nand4_1 _23843_ (.B(_07214_),
    .C(_07215_),
    .A(_07213_),
    .Y(_07217_),
    .D(_07216_));
 sg13g2_mux2_1 _23844_ (.A0(\top_ihp.oisc.regs[14][5] ),
    .A1(\top_ihp.oisc.regs[12][5] ),
    .S(net725),
    .X(_07218_));
 sg13g2_a22oi_1 _23845_ (.Y(_07219_),
    .B1(_06484_),
    .B2(_07218_),
    .A2(net547),
    .A1(\top_ihp.oisc.regs[1][5] ));
 sg13g2_a22oi_1 _23846_ (.Y(_07220_),
    .B1(net551),
    .B2(\top_ihp.oisc.regs[25][5] ),
    .A2(net552),
    .A1(\top_ihp.oisc.regs[20][5] ));
 sg13g2_and2_1 _23847_ (.A(_07219_),
    .B(_07220_),
    .X(_07221_));
 sg13g2_and2_1 _23848_ (.A(\top_ihp.oisc.regs[21][5] ),
    .B(_05390_),
    .X(_07222_));
 sg13g2_a221oi_1 _23849_ (.B2(\top_ihp.oisc.regs[10][5] ),
    .C1(_07222_),
    .B1(_05905_),
    .A1(\top_ihp.oisc.regs[26][5] ),
    .Y(_07223_),
    .A2(net367));
 sg13g2_a22oi_1 _23850_ (.Y(_07224_),
    .B1(net160),
    .B2(\top_ihp.oisc.regs[17][5] ),
    .A2(_05883_),
    .A1(\top_ihp.oisc.regs[9][5] ));
 sg13g2_a22oi_1 _23851_ (.Y(_07225_),
    .B1(net345),
    .B2(\top_ihp.oisc.regs[5][5] ),
    .A2(net664),
    .A1(\top_ihp.oisc.regs[28][5] ));
 sg13g2_nand4_1 _23852_ (.B(_07223_),
    .C(_07224_),
    .A(_07221_),
    .Y(_07226_),
    .D(_07225_));
 sg13g2_nor2_1 _23853_ (.A(_08140_),
    .B(net804),
    .Y(_07227_));
 sg13g2_a221oi_1 _23854_ (.B2(\top_ihp.oisc.regs[8][5] ),
    .C1(_07227_),
    .B1(net665),
    .A1(\top_ihp.oisc.regs[23][5] ),
    .Y(_07228_),
    .A2(net720));
 sg13g2_a22oi_1 _23855_ (.Y(_07229_),
    .B1(net343),
    .B2(\top_ihp.oisc.regs[18][5] ),
    .A2(net342),
    .A1(\top_ihp.oisc.regs[7][5] ));
 sg13g2_a22oi_1 _23856_ (.Y(_07230_),
    .B1(net167),
    .B2(\top_ihp.oisc.regs[24][5] ),
    .A2(_06163_),
    .A1(\top_ihp.oisc.regs[15][5] ));
 sg13g2_a22oi_1 _23857_ (.Y(_07231_),
    .B1(_06002_),
    .B2(\top_ihp.oisc.regs[19][5] ),
    .A2(_06156_),
    .A1(\top_ihp.oisc.regs[4][5] ));
 sg13g2_nand4_1 _23858_ (.B(_07229_),
    .C(_07230_),
    .A(_07228_),
    .Y(_07232_),
    .D(_07231_));
 sg13g2_a22oi_1 _23859_ (.Y(_07233_),
    .B1(_05885_),
    .B2(\top_ihp.oisc.regs[6][5] ),
    .A2(net166),
    .A1(\top_ihp.oisc.regs[3][5] ));
 sg13g2_a22oi_1 _23860_ (.Y(_07234_),
    .B1(net183),
    .B2(\top_ihp.oisc.regs[16][5] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[22][5] ));
 sg13g2_a22oi_1 _23861_ (.Y(_07235_),
    .B1(net180),
    .B2(\top_ihp.oisc.regs[13][5] ),
    .A2(net203),
    .A1(\top_ihp.oisc.regs[29][5] ));
 sg13g2_a22oi_1 _23862_ (.Y(_07236_),
    .B1(net179),
    .B2(\top_ihp.oisc.regs[2][5] ),
    .A2(net380),
    .A1(\top_ihp.oisc.regs[11][5] ));
 sg13g2_nand4_1 _23863_ (.B(_07234_),
    .C(_07235_),
    .A(_07233_),
    .Y(_07237_),
    .D(_07236_));
 sg13g2_nor4_1 _23864_ (.A(_07217_),
    .B(_07226_),
    .C(_07232_),
    .D(_07237_),
    .Y(_07238_));
 sg13g2_a21oi_1 _23865_ (.A1(_00209_),
    .A2(_05707_),
    .Y(_07239_),
    .B1(_05744_));
 sg13g2_nor2_1 _23866_ (.A(_07227_),
    .B(_07239_),
    .Y(_07240_));
 sg13g2_a21oi_1 _23867_ (.A1(_07212_),
    .A2(_07238_),
    .Y(_00415_),
    .B1(_07240_));
 sg13g2_a22oi_1 _23868_ (.Y(_07241_),
    .B1(net408),
    .B2(\top_ihp.oisc.regs[35][6] ),
    .A2(net539),
    .A1(\top_ihp.oisc.regs[34][6] ));
 sg13g2_a22oi_1 _23869_ (.Y(_07242_),
    .B1(net171),
    .B2(\top_ihp.oisc.regs[60][6] ),
    .A2(_05732_),
    .A1(\top_ihp.oisc.regs[49][6] ));
 sg13g2_a22oi_1 _23870_ (.Y(_07243_),
    .B1(net391),
    .B2(\top_ihp.oisc.regs[33][6] ),
    .A2(_05652_),
    .A1(\top_ihp.oisc.regs[54][6] ));
 sg13g2_a22oi_1 _23871_ (.Y(_07244_),
    .B1(net419),
    .B2(\top_ihp.oisc.regs[44][6] ),
    .A2(_05673_),
    .A1(\top_ihp.oisc.regs[61][6] ));
 sg13g2_nand4_1 _23872_ (.B(_07242_),
    .C(_07243_),
    .A(_07241_),
    .Y(_07245_),
    .D(_07244_));
 sg13g2_a22oi_1 _23873_ (.Y(_07246_),
    .B1(net349),
    .B2(\top_ihp.oisc.regs[46][6] ),
    .A2(net192),
    .A1(\top_ihp.oisc.regs[62][6] ));
 sg13g2_a22oi_1 _23874_ (.Y(_07247_),
    .B1(net392),
    .B2(\top_ihp.oisc.regs[52][6] ),
    .A2(net375),
    .A1(\top_ihp.oisc.regs[36][6] ));
 sg13g2_a22oi_1 _23875_ (.Y(_07248_),
    .B1(net397),
    .B2(\top_ihp.oisc.regs[37][6] ),
    .A2(net411),
    .A1(\top_ihp.oisc.regs[45][6] ));
 sg13g2_a22oi_1 _23876_ (.Y(_07249_),
    .B1(_05701_),
    .B2(\top_ihp.oisc.regs[8][6] ),
    .A2(net721),
    .A1(\top_ihp.oisc.regs[14][6] ));
 sg13g2_nor2_1 _23877_ (.A(_05512_),
    .B(_07249_),
    .Y(_07250_));
 sg13g2_a21oi_1 _23878_ (.A1(\top_ihp.oisc.regs[32][6] ),
    .A2(net338),
    .Y(_07251_),
    .B1(_07250_));
 sg13g2_nand4_1 _23879_ (.B(_07247_),
    .C(_07248_),
    .A(_07246_),
    .Y(_07252_),
    .D(_07251_));
 sg13g2_mux2_1 _23880_ (.A0(\top_ihp.oisc.regs[24][6] ),
    .A1(\top_ihp.oisc.regs[16][6] ),
    .S(net662),
    .X(_07253_));
 sg13g2_a22oi_1 _23881_ (.Y(_07254_),
    .B1(_07253_),
    .B2(_06277_),
    .A2(net343),
    .A1(\top_ihp.oisc.regs[18][6] ));
 sg13g2_a22oi_1 _23882_ (.Y(_07255_),
    .B1(_05889_),
    .B2(\top_ihp.oisc.regs[12][6] ),
    .A2(net434),
    .A1(\top_ihp.oisc.regs[20][6] ));
 sg13g2_a22oi_1 _23883_ (.Y(_07256_),
    .B1(net749),
    .B2(\top_ihp.oisc.regs[6][6] ),
    .A2(net724),
    .A1(\top_ihp.oisc.regs[7][6] ));
 sg13g2_nand3_1 _23884_ (.B(net750),
    .C(_05701_),
    .A(\top_ihp.oisc.regs[17][6] ),
    .Y(_07257_));
 sg13g2_o21ai_1 _23885_ (.B1(_07257_),
    .Y(_07258_),
    .A1(_05418_),
    .A2(_07256_));
 sg13g2_a21oi_1 _23886_ (.A1(\top_ihp.oisc.regs[10][6] ),
    .A2(_06426_),
    .Y(_07259_),
    .B1(_07258_));
 sg13g2_a22oi_1 _23887_ (.Y(_07260_),
    .B1(net185),
    .B2(\top_ihp.oisc.regs[9][6] ),
    .A2(net203),
    .A1(\top_ihp.oisc.regs[29][6] ));
 sg13g2_nand4_1 _23888_ (.B(_07255_),
    .C(_07259_),
    .A(_07254_),
    .Y(_07261_),
    .D(_07260_));
 sg13g2_a22oi_1 _23889_ (.Y(_07262_),
    .B1(_06068_),
    .B2(\top_ihp.oisc.regs[26][6] ),
    .A2(_05901_),
    .A1(\top_ihp.oisc.regs[2][6] ));
 sg13g2_a22oi_1 _23890_ (.Y(_07263_),
    .B1(net181),
    .B2(\top_ihp.oisc.regs[15][6] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[22][6] ));
 sg13g2_a22oi_1 _23891_ (.Y(_07264_),
    .B1(_05523_),
    .B2(\top_ihp.oisc.regs[5][6] ),
    .A2(net750),
    .A1(\top_ihp.oisc.regs[21][6] ));
 sg13g2_nand3_1 _23892_ (.B(net750),
    .C(_05598_),
    .A(\top_ihp.oisc.regs[23][6] ),
    .Y(_07265_));
 sg13g2_o21ai_1 _23893_ (.B1(_07265_),
    .Y(_07266_),
    .A1(_06636_),
    .A2(_07264_));
 sg13g2_a221oi_1 _23894_ (.B2(\top_ihp.oisc.regs[43][6] ),
    .C1(_07266_),
    .B1(net362),
    .A1(_08122_),
    .Y(_07267_),
    .A2(_04087_));
 sg13g2_nand3_1 _23895_ (.B(_07263_),
    .C(_07267_),
    .A(_07262_),
    .Y(_07268_));
 sg13g2_nor4_1 _23896_ (.A(_07245_),
    .B(_07252_),
    .C(_07261_),
    .D(_07268_),
    .Y(_07269_));
 sg13g2_a22oi_1 _23897_ (.Y(_07270_),
    .B1(_05833_),
    .B2(\top_ihp.oisc.regs[59][6] ),
    .A2(net356),
    .A1(\top_ihp.oisc.regs[31][6] ));
 sg13g2_a22oi_1 _23898_ (.Y(_07271_),
    .B1(net395),
    .B2(\top_ihp.oisc.regs[41][6] ),
    .A2(_05854_),
    .A1(\top_ihp.oisc.regs[27][6] ));
 sg13g2_a22oi_1 _23899_ (.Y(_07272_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[47][6] ),
    .A2(_05843_),
    .A1(\top_ihp.oisc.regs[40][6] ));
 sg13g2_a22oi_1 _23900_ (.Y(_07273_),
    .B1(net384),
    .B2(\top_ihp.oisc.regs[38][6] ),
    .A2(_05783_),
    .A1(\top_ihp.oisc.regs[63][6] ));
 sg13g2_nand4_1 _23901_ (.B(_07271_),
    .C(_07272_),
    .A(_07270_),
    .Y(_07274_),
    .D(_07273_));
 sg13g2_a22oi_1 _23902_ (.Y(_07275_),
    .B1(net398),
    .B2(\top_ihp.oisc.regs[55][6] ),
    .A2(net355),
    .A1(\top_ihp.oisc.regs[51][6] ));
 sg13g2_a22oi_1 _23903_ (.Y(_07276_),
    .B1(_05799_),
    .B2(\top_ihp.oisc.regs[50][6] ),
    .A2(net348),
    .A1(\top_ihp.oisc.regs[57][6] ));
 sg13g2_a22oi_1 _23904_ (.Y(_07277_),
    .B1(net195),
    .B2(\top_ihp.oisc.regs[58][6] ),
    .A2(net344),
    .A1(\top_ihp.oisc.regs[53][6] ));
 sg13g2_a22oi_1 _23905_ (.Y(_07278_),
    .B1(net197),
    .B2(\top_ihp.oisc.regs[48][6] ),
    .A2(net336),
    .A1(\top_ihp.oisc.regs[42][6] ));
 sg13g2_nand4_1 _23906_ (.B(_07276_),
    .C(_07277_),
    .A(_07275_),
    .Y(_07279_),
    .D(_07278_));
 sg13g2_a22oi_1 _23907_ (.Y(_07280_),
    .B1(_05898_),
    .B2(\top_ihp.oisc.regs[13][6] ),
    .A2(_05506_),
    .A1(\top_ihp.oisc.regs[1][6] ));
 sg13g2_a22oi_1 _23908_ (.Y(_07281_),
    .B1(_06246_),
    .B2(\top_ihp.oisc.regs[19][6] ),
    .A2(_05578_),
    .A1(\top_ihp.oisc.regs[11][6] ));
 sg13g2_a22oi_1 _23909_ (.Y(_07282_),
    .B1(net664),
    .B2(\top_ihp.oisc.regs[28][6] ),
    .A2(net551),
    .A1(\top_ihp.oisc.regs[25][6] ));
 sg13g2_a22oi_1 _23910_ (.Y(_07283_),
    .B1(net401),
    .B2(\top_ihp.oisc.regs[3][6] ),
    .A2(_05499_),
    .A1(\top_ihp.oisc.regs[4][6] ));
 sg13g2_and4_1 _23911_ (.A(_07280_),
    .B(_07281_),
    .C(_07282_),
    .D(_07283_),
    .X(_07284_));
 sg13g2_nand2_1 _23912_ (.Y(_07285_),
    .A(\top_ihp.oisc.regs[39][6] ),
    .B(_05966_));
 sg13g2_a22oi_1 _23913_ (.Y(_07286_),
    .B1(_05805_),
    .B2(\top_ihp.oisc.regs[56][6] ),
    .A2(net388),
    .A1(\top_ihp.oisc.regs[30][6] ));
 sg13g2_nand4_1 _23914_ (.B(_07284_),
    .C(_07285_),
    .A(_06017_),
    .Y(_07287_),
    .D(_07286_));
 sg13g2_nor3_1 _23915_ (.A(_07274_),
    .B(_07279_),
    .C(_07287_),
    .Y(_07288_));
 sg13g2_nand2_1 _23916_ (.Y(_07289_),
    .A(_00210_),
    .B(net59));
 sg13g2_a22oi_1 _23917_ (.Y(_07290_),
    .B1(net27),
    .B2(_07289_),
    .A2(net746),
    .A1(_08122_));
 sg13g2_a21oi_1 _23918_ (.A1(_07269_),
    .A2(_07288_),
    .Y(_00416_),
    .B1(_07290_));
 sg13g2_a22oi_1 _23919_ (.Y(_07291_),
    .B1(net171),
    .B2(\top_ihp.oisc.regs[60][7] ),
    .A2(net198),
    .A1(\top_ihp.oisc.regs[59][7] ));
 sg13g2_a22oi_1 _23920_ (.Y(_07292_),
    .B1(net362),
    .B2(\top_ihp.oisc.regs[43][7] ),
    .A2(_05830_),
    .A1(\top_ihp.oisc.regs[31][7] ));
 sg13g2_a22oi_1 _23921_ (.Y(_07293_),
    .B1(net399),
    .B2(\top_ihp.oisc.regs[58][7] ),
    .A2(_05714_),
    .A1(\top_ihp.oisc.regs[48][7] ));
 sg13g2_a22oi_1 _23922_ (.Y(_07294_),
    .B1(net364),
    .B2(\top_ihp.oisc.regs[52][7] ),
    .A2(_05635_),
    .A1(\top_ihp.oisc.regs[40][7] ));
 sg13g2_nand4_1 _23923_ (.B(_07292_),
    .C(_07293_),
    .A(_07291_),
    .Y(_07295_),
    .D(_07294_));
 sg13g2_a22oi_1 _23924_ (.Y(_07296_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[47][7] ),
    .A2(net175),
    .A1(\top_ihp.oisc.regs[61][7] ));
 sg13g2_a22oi_1 _23925_ (.Y(_07297_),
    .B1(_06020_),
    .B2(\top_ihp.oisc.regs[57][7] ),
    .A2(net375),
    .A1(\top_ihp.oisc.regs[36][7] ));
 sg13g2_nand3_1 _23926_ (.B(_07296_),
    .C(_07297_),
    .A(_05918_),
    .Y(_07298_));
 sg13g2_nand2_1 _23927_ (.Y(_07299_),
    .A(_08116_),
    .B(net835));
 sg13g2_a22oi_1 _23928_ (.Y(_07300_),
    .B1(_05824_),
    .B2(\top_ihp.oisc.regs[23][7] ),
    .A2(_05820_),
    .A1(\top_ihp.oisc.regs[21][7] ));
 sg13g2_a22oi_1 _23929_ (.Y(_07301_),
    .B1(_05565_),
    .B2(\top_ihp.oisc.regs[6][7] ),
    .A2(_05542_),
    .A1(\top_ihp.oisc.regs[28][7] ));
 sg13g2_nand3_1 _23930_ (.B(_07300_),
    .C(_07301_),
    .A(_07299_),
    .Y(_07302_));
 sg13g2_a221oi_1 _23931_ (.B2(\top_ihp.oisc.regs[37][7] ),
    .C1(_07302_),
    .B1(net347),
    .A1(\top_ihp.oisc.regs[42][7] ),
    .Y(_07303_),
    .A2(net416));
 sg13g2_a22oi_1 _23932_ (.Y(_07304_),
    .B1(_05793_),
    .B2(\top_ihp.oisc.regs[55][7] ),
    .A2(net422),
    .A1(\top_ihp.oisc.regs[32][7] ));
 sg13g2_a22oi_1 _23933_ (.Y(_07305_),
    .B1(net386),
    .B2(\top_ihp.oisc.regs[49][7] ),
    .A2(net199),
    .A1(\top_ihp.oisc.regs[50][7] ));
 sg13g2_nand3_1 _23934_ (.B(_07304_),
    .C(_07305_),
    .A(_07303_),
    .Y(_07306_));
 sg13g2_a22oi_1 _23935_ (.Y(_07307_),
    .B1(_05722_),
    .B2(\top_ihp.oisc.regs[33][7] ),
    .A2(_05961_),
    .A1(\top_ihp.oisc.regs[51][7] ));
 sg13g2_a22oi_1 _23936_ (.Y(_07308_),
    .B1(net202),
    .B2(\top_ihp.oisc.regs[44][7] ),
    .A2(_05873_),
    .A1(\top_ihp.oisc.regs[34][7] ));
 sg13g2_a22oi_1 _23937_ (.Y(_07309_),
    .B1(_05802_),
    .B2(\top_ihp.oisc.regs[45][7] ),
    .A2(net176),
    .A1(\top_ihp.oisc.regs[62][7] ));
 sg13g2_a22oi_1 _23938_ (.Y(_07310_),
    .B1(net410),
    .B2(\top_ihp.oisc.regs[41][7] ),
    .A2(net378),
    .A1(\top_ihp.oisc.regs[38][7] ));
 sg13g2_nand4_1 _23939_ (.B(_07308_),
    .C(_07309_),
    .A(_07307_),
    .Y(_07311_),
    .D(_07310_));
 sg13g2_nor4_2 _23940_ (.A(_07295_),
    .B(_07298_),
    .C(_07306_),
    .Y(_07312_),
    .D(_07311_));
 sg13g2_a22oi_1 _23941_ (.Y(_07313_),
    .B1(net187),
    .B2(\top_ihp.oisc.regs[56][7] ),
    .A2(net414),
    .A1(\top_ihp.oisc.regs[30][7] ));
 sg13g2_a22oi_1 _23942_ (.Y(_07314_),
    .B1(net382),
    .B2(\top_ihp.oisc.regs[27][7] ),
    .A2(net540),
    .A1(\top_ihp.oisc.regs[20][7] ));
 sg13g2_a22oi_1 _23943_ (.Y(_07315_),
    .B1(net337),
    .B2(\top_ihp.oisc.regs[39][7] ),
    .A2(_05647_),
    .A1(\top_ihp.oisc.regs[53][7] ));
 sg13g2_a22oi_1 _23944_ (.Y(_07316_),
    .B1(net406),
    .B2(\top_ihp.oisc.regs[46][7] ),
    .A2(_05664_),
    .A1(\top_ihp.oisc.regs[63][7] ));
 sg13g2_nand4_1 _23945_ (.B(_07314_),
    .C(_07315_),
    .A(_07313_),
    .Y(_07317_),
    .D(_07316_));
 sg13g2_and2_1 _23946_ (.A(\top_ihp.oisc.regs[29][7] ),
    .B(net429),
    .X(_07318_));
 sg13g2_a221oi_1 _23947_ (.B2(\top_ihp.oisc.regs[12][7] ),
    .C1(_07318_),
    .B1(net372),
    .A1(\top_ihp.oisc.regs[25][7] ),
    .Y(_07319_),
    .A2(net551));
 sg13g2_a22oi_1 _23948_ (.Y(_07320_),
    .B1(net402),
    .B2(\top_ihp.oisc.regs[24][7] ),
    .A2(_05430_),
    .A1(\top_ihp.oisc.regs[7][7] ));
 sg13g2_a22oi_1 _23949_ (.Y(_07321_),
    .B1(net164),
    .B2(\top_ihp.oisc.regs[9][7] ),
    .A2(net432),
    .A1(\top_ihp.oisc.regs[4][7] ));
 sg13g2_a22oi_1 _23950_ (.Y(_07322_),
    .B1(net353),
    .B2(\top_ihp.oisc.regs[35][7] ),
    .A2(net201),
    .A1(\top_ihp.oisc.regs[54][7] ));
 sg13g2_nand4_1 _23951_ (.B(_07320_),
    .C(_07321_),
    .A(_07319_),
    .Y(_07323_),
    .D(_07322_));
 sg13g2_a22oi_1 _23952_ (.Y(_07324_),
    .B1(net169),
    .B2(\top_ihp.oisc.regs[11][7] ),
    .A2(_06238_),
    .A1(\top_ihp.oisc.regs[17][7] ));
 sg13g2_a22oi_1 _23953_ (.Y(_07325_),
    .B1(net350),
    .B2(\top_ihp.oisc.regs[19][7] ),
    .A2(net431),
    .A1(\top_ihp.oisc.regs[1][7] ));
 sg13g2_a22oi_1 _23954_ (.Y(_07326_),
    .B1(_06115_),
    .B2(\top_ihp.oisc.regs[5][7] ),
    .A2(net546),
    .A1(\top_ihp.oisc.regs[14][7] ));
 sg13g2_a22oi_1 _23955_ (.Y(_07327_),
    .B1(net180),
    .B2(\top_ihp.oisc.regs[13][7] ),
    .A2(net533),
    .A1(\top_ihp.oisc.regs[22][7] ));
 sg13g2_nand4_1 _23956_ (.B(_07325_),
    .C(_07326_),
    .A(_07324_),
    .Y(_07328_),
    .D(_07327_));
 sg13g2_a22oi_1 _23957_ (.Y(_07329_),
    .B1(_05901_),
    .B2(\top_ihp.oisc.regs[2][7] ),
    .A2(_06063_),
    .A1(\top_ihp.oisc.regs[18][7] ));
 sg13g2_a22oi_1 _23958_ (.Y(_07330_),
    .B1(_05893_),
    .B2(\top_ihp.oisc.regs[16][7] ),
    .A2(net162),
    .A1(\top_ihp.oisc.regs[15][7] ));
 sg13g2_a22oi_1 _23959_ (.Y(_07331_),
    .B1(net536),
    .B2(\top_ihp.oisc.regs[8][7] ),
    .A2(_05911_),
    .A1(\top_ihp.oisc.regs[26][7] ));
 sg13g2_a22oi_1 _23960_ (.Y(_07332_),
    .B1(_06426_),
    .B2(\top_ihp.oisc.regs[10][7] ),
    .A2(_06059_),
    .A1(\top_ihp.oisc.regs[3][7] ));
 sg13g2_nand4_1 _23961_ (.B(_07330_),
    .C(_07331_),
    .A(_07329_),
    .Y(_07333_),
    .D(_07332_));
 sg13g2_nor4_1 _23962_ (.A(_07317_),
    .B(_07323_),
    .C(_07328_),
    .D(_07333_),
    .Y(_07334_));
 sg13g2_inv_1 _23963_ (.Y(_07335_),
    .A(_00211_));
 sg13g2_o21ai_1 _23964_ (.B1(net27),
    .Y(_07336_),
    .A1(_07335_),
    .A2(net62));
 sg13g2_a22oi_1 _23965_ (.Y(_00417_),
    .B1(_07336_),
    .B2(_07299_),
    .A2(_07334_),
    .A1(_07312_));
 sg13g2_a22oi_1 _23966_ (.Y(_07337_),
    .B1(_06029_),
    .B2(\top_ihp.oisc.regs[60][8] ),
    .A2(net406),
    .A1(\top_ihp.oisc.regs[46][8] ));
 sg13g2_a22oi_1 _23967_ (.Y(_07338_),
    .B1(net340),
    .B2(\top_ihp.oisc.regs[41][8] ),
    .A2(_05983_),
    .A1(\top_ihp.oisc.regs[62][8] ));
 sg13g2_a22oi_1 _23968_ (.Y(_07339_),
    .B1(net381),
    .B2(\top_ihp.oisc.regs[48][8] ),
    .A2(_06141_),
    .A1(\top_ihp.oisc.regs[32][8] ));
 sg13g2_a22oi_1 _23969_ (.Y(_07340_),
    .B1(_05545_),
    .B2(\top_ihp.oisc.regs[22][8] ),
    .A2(net722),
    .A1(\top_ihp.oisc.regs[28][8] ));
 sg13g2_nor2_1 _23970_ (.A(_05540_),
    .B(_07340_),
    .Y(_07341_));
 sg13g2_a21oi_1 _23971_ (.A1(\top_ihp.oisc.regs[63][8] ),
    .A2(net413),
    .Y(_07342_),
    .B1(_07341_));
 sg13g2_nand4_1 _23972_ (.B(_07338_),
    .C(_07339_),
    .A(_07337_),
    .Y(_07343_),
    .D(_07342_));
 sg13g2_a22oi_1 _23973_ (.Y(_07344_),
    .B1(net193),
    .B2(\top_ihp.oisc.regs[56][8] ),
    .A2(net411),
    .A1(\top_ihp.oisc.regs[45][8] ));
 sg13g2_a22oi_1 _23974_ (.Y(_07345_),
    .B1(net399),
    .B2(\top_ihp.oisc.regs[58][8] ),
    .A2(_06080_),
    .A1(\top_ihp.oisc.regs[27][8] ));
 sg13g2_a22oi_1 _23975_ (.Y(_07346_),
    .B1(_06143_),
    .B2(\top_ihp.oisc.regs[39][8] ),
    .A2(net414),
    .A1(\top_ihp.oisc.regs[30][8] ));
 sg13g2_a22oi_1 _23976_ (.Y(_07347_),
    .B1(net188),
    .B2(\top_ihp.oisc.regs[50][8] ),
    .A2(_05986_),
    .A1(\top_ihp.oisc.regs[40][8] ));
 sg13g2_nand4_1 _23977_ (.B(_07345_),
    .C(_07346_),
    .A(_07344_),
    .Y(_07348_),
    .D(_07347_));
 sg13g2_a22oi_1 _23978_ (.Y(_07349_),
    .B1(net369),
    .B2(\top_ihp.oisc.regs[2][8] ),
    .A2(net370),
    .A1(\top_ihp.oisc.regs[13][8] ));
 sg13g2_a22oi_1 _23979_ (.Y(_07350_),
    .B1(net427),
    .B2(\top_ihp.oisc.regs[17][8] ),
    .A2(net551),
    .A1(\top_ihp.oisc.regs[25][8] ));
 sg13g2_a22oi_1 _23980_ (.Y(_07351_),
    .B1(_05784_),
    .B2(\top_ihp.oisc.regs[6][8] ),
    .A2(net554),
    .A1(\top_ihp.oisc.regs[7][8] ));
 sg13g2_a22oi_1 _23981_ (.Y(_07352_),
    .B1(net432),
    .B2(\top_ihp.oisc.regs[4][8] ),
    .A2(_05472_),
    .A1(\top_ihp.oisc.regs[20][8] ));
 sg13g2_nand4_1 _23982_ (.B(_07350_),
    .C(_07351_),
    .A(_07349_),
    .Y(_07353_),
    .D(_07352_));
 sg13g2_nand2b_1 _23983_ (.Y(_07354_),
    .B(net57),
    .A_N(_07353_));
 sg13g2_a22oi_1 _23984_ (.Y(_07355_),
    .B1(net386),
    .B2(\top_ihp.oisc.regs[49][8] ),
    .A2(net412),
    .A1(\top_ihp.oisc.regs[43][8] ));
 sg13g2_a22oi_1 _23985_ (.Y(_07356_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[47][8] ),
    .A2(net397),
    .A1(\top_ihp.oisc.regs[37][8] ));
 sg13g2_a22oi_1 _23986_ (.Y(_07357_),
    .B1(_05736_),
    .B2(\top_ihp.oisc.regs[55][8] ),
    .A2(net336),
    .A1(\top_ihp.oisc.regs[42][8] ));
 sg13g2_a22oi_1 _23987_ (.Y(_07358_),
    .B1(net384),
    .B2(\top_ihp.oisc.regs[38][8] ),
    .A2(net344),
    .A1(\top_ihp.oisc.regs[53][8] ));
 sg13g2_nand4_1 _23988_ (.B(_07356_),
    .C(_07357_),
    .A(_07355_),
    .Y(_07359_),
    .D(_07358_));
 sg13g2_nor4_1 _23989_ (.A(_07343_),
    .B(_07348_),
    .C(_07354_),
    .D(_07359_),
    .Y(_07360_));
 sg13g2_a22oi_1 _23990_ (.Y(_07361_),
    .B1(_06163_),
    .B2(\top_ihp.oisc.regs[15][8] ),
    .A2(_06149_),
    .A1(\top_ihp.oisc.regs[9][8] ));
 sg13g2_a22oi_1 _23991_ (.Y(_07362_),
    .B1(net345),
    .B2(\top_ihp.oisc.regs[5][8] ),
    .A2(net372),
    .A1(\top_ihp.oisc.regs[12][8] ));
 sg13g2_a22oi_1 _23992_ (.Y(_07363_),
    .B1(net335),
    .B2(\top_ihp.oisc.regs[19][8] ),
    .A2(net534),
    .A1(\top_ihp.oisc.regs[18][8] ));
 sg13g2_a22oi_1 _23993_ (.Y(_07364_),
    .B1(_05892_),
    .B2(\top_ihp.oisc.regs[16][8] ),
    .A2(_05778_),
    .A1(\top_ihp.oisc.regs[3][8] ));
 sg13g2_nand4_1 _23994_ (.B(_07362_),
    .C(_07363_),
    .A(_07361_),
    .Y(_07365_),
    .D(_07364_));
 sg13g2_a22oi_1 _23995_ (.Y(_07366_),
    .B1(net360),
    .B2(\top_ihp.oisc.regs[33][8] ),
    .A2(net542),
    .A1(\top_ihp.oisc.regs[34][8] ));
 sg13g2_nand2_1 _23996_ (.Y(_07367_),
    .A(_08100_),
    .B(net803));
 sg13g2_a22oi_1 _23997_ (.Y(_07368_),
    .B1(net720),
    .B2(\top_ihp.oisc.regs[23][8] ),
    .A2(net666),
    .A1(\top_ihp.oisc.regs[21][8] ));
 sg13g2_a22oi_1 _23998_ (.Y(_07369_),
    .B1(net367),
    .B2(\top_ihp.oisc.regs[26][8] ),
    .A2(_05506_),
    .A1(\top_ihp.oisc.regs[1][8] ));
 sg13g2_nand4_1 _23999_ (.B(_07367_),
    .C(_07368_),
    .A(_07366_),
    .Y(_07370_),
    .D(_07369_));
 sg13g2_a22oi_1 _24000_ (.Y(_07371_),
    .B1(net196),
    .B2(\top_ihp.oisc.regs[54][8] ),
    .A2(net435),
    .A1(\top_ihp.oisc.regs[31][8] ));
 sg13g2_a22oi_1 _24001_ (.Y(_07372_),
    .B1(net408),
    .B2(\top_ihp.oisc.regs[35][8] ),
    .A2(net420),
    .A1(\top_ihp.oisc.regs[51][8] ));
 sg13g2_a22oi_1 _24002_ (.Y(_07373_),
    .B1(net191),
    .B2(\top_ihp.oisc.regs[59][8] ),
    .A2(net375),
    .A1(\top_ihp.oisc.regs[36][8] ));
 sg13g2_a22oi_1 _24003_ (.Y(_07374_),
    .B1(net161),
    .B2(\top_ihp.oisc.regs[44][8] ),
    .A2(net333),
    .A1(\top_ihp.oisc.regs[57][8] ));
 sg13g2_nand4_1 _24004_ (.B(_07372_),
    .C(_07373_),
    .A(_07371_),
    .Y(_07375_),
    .D(_07374_));
 sg13g2_nand2_1 _24005_ (.Y(_07376_),
    .A(\top_ihp.oisc.regs[11][8] ),
    .B(net169));
 sg13g2_a22oi_1 _24006_ (.Y(_07377_),
    .B1(_06102_),
    .B2(\top_ihp.oisc.regs[24][8] ),
    .A2(net203),
    .A1(\top_ihp.oisc.regs[29][8] ));
 sg13g2_a22oi_1 _24007_ (.Y(_07378_),
    .B1(net405),
    .B2(\top_ihp.oisc.regs[52][8] ),
    .A2(_05965_),
    .A1(\top_ihp.oisc.regs[61][8] ));
 sg13g2_mux2_1 _24008_ (.A0(\top_ihp.oisc.regs[14][8] ),
    .A1(\top_ihp.oisc.regs[10][8] ),
    .S(_05491_),
    .X(_07379_));
 sg13g2_a22oi_1 _24009_ (.Y(_07380_),
    .B1(_07379_),
    .B2(net550),
    .A2(_05701_),
    .A1(\top_ihp.oisc.regs[8][8] ));
 sg13g2_nand2b_1 _24010_ (.Y(_07381_),
    .B(_06175_),
    .A_N(_07380_));
 sg13g2_nand4_1 _24011_ (.B(_07377_),
    .C(_07378_),
    .A(_07376_),
    .Y(_07382_),
    .D(_07381_));
 sg13g2_nor4_1 _24012_ (.A(_07365_),
    .B(_07370_),
    .C(_07375_),
    .D(_07382_),
    .Y(_07383_));
 sg13g2_a21o_1 _24013_ (.A2(net63),
    .A1(_00212_),
    .B1(net58),
    .X(_07384_));
 sg13g2_a22oi_1 _24014_ (.Y(_00418_),
    .B1(_07384_),
    .B2(_07367_),
    .A2(_07383_),
    .A1(_07360_));
 sg13g2_a22oi_1 _24015_ (.Y(_07385_),
    .B1(net410),
    .B2(\top_ihp.oisc.regs[41][9] ),
    .A2(_05461_),
    .A1(\top_ihp.oisc.regs[31][9] ));
 sg13g2_a22oi_1 _24016_ (.Y(_07386_),
    .B1(net378),
    .B2(\top_ihp.oisc.regs[38][9] ),
    .A2(_05872_),
    .A1(\top_ihp.oisc.regs[36][9] ));
 sg13g2_a22oi_1 _24017_ (.Y(_07387_),
    .B1(net199),
    .B2(\top_ihp.oisc.regs[50][9] ),
    .A2(net352),
    .A1(\top_ihp.oisc.regs[43][9] ));
 sg13g2_a22oi_1 _24018_ (.Y(_07388_),
    .B1(net358),
    .B2(\top_ihp.oisc.regs[47][9] ),
    .A2(_05869_),
    .A1(\top_ihp.oisc.regs[53][9] ));
 sg13g2_nand4_1 _24019_ (.B(_07386_),
    .C(_07387_),
    .A(_07385_),
    .Y(_07389_),
    .D(_07388_));
 sg13g2_a22oi_1 _24020_ (.Y(_07390_),
    .B1(_05939_),
    .B2(\top_ihp.oisc.regs[62][9] ),
    .A2(_05588_),
    .A1(\top_ihp.oisc.regs[60][9] ));
 sg13g2_a22oi_1 _24021_ (.Y(_07391_),
    .B1(net376),
    .B2(\top_ihp.oisc.regs[51][9] ),
    .A2(net200),
    .A1(\top_ihp.oisc.regs[61][9] ));
 sg13g2_a22oi_1 _24022_ (.Y(_07392_),
    .B1(net359),
    .B2(\top_ihp.oisc.regs[55][9] ),
    .A2(net416),
    .A1(\top_ihp.oisc.regs[42][9] ));
 sg13g2_a22oi_1 _24023_ (.Y(_07393_),
    .B1(net399),
    .B2(\top_ihp.oisc.regs[58][9] ),
    .A2(net201),
    .A1(\top_ihp.oisc.regs[54][9] ));
 sg13g2_nand4_1 _24024_ (.B(_07391_),
    .C(_07392_),
    .A(_07390_),
    .Y(_07394_),
    .D(_07393_));
 sg13g2_a22oi_1 _24025_ (.Y(_07395_),
    .B1(net386),
    .B2(\top_ihp.oisc.regs[49][9] ),
    .A2(net385),
    .A1(\top_ihp.oisc.regs[40][9] ));
 sg13g2_a22oi_1 _24026_ (.Y(_07396_),
    .B1(net193),
    .B2(\top_ihp.oisc.regs[56][9] ),
    .A2(net198),
    .A1(\top_ihp.oisc.regs[59][9] ));
 sg13g2_a22oi_1 _24027_ (.Y(_07397_),
    .B1(net381),
    .B2(\top_ihp.oisc.regs[48][9] ),
    .A2(net338),
    .A1(\top_ihp.oisc.regs[32][9] ));
 sg13g2_a22oi_1 _24028_ (.Y(_07398_),
    .B1(net360),
    .B2(\top_ihp.oisc.regs[33][9] ),
    .A2(net400),
    .A1(\top_ihp.oisc.regs[63][9] ));
 sg13g2_nand4_1 _24029_ (.B(_07396_),
    .C(_07397_),
    .A(_07395_),
    .Y(_07399_),
    .D(_07398_));
 sg13g2_nand2_1 _24030_ (.Y(_07400_),
    .A(\top_ihp.oisc.regs[30][9] ),
    .B(net388));
 sg13g2_a22oi_1 _24031_ (.Y(_07401_),
    .B1(net396),
    .B2(\top_ihp.oisc.regs[46][9] ),
    .A2(net348),
    .A1(\top_ihp.oisc.regs[57][9] ));
 sg13g2_nand3_1 _24032_ (.B(_07400_),
    .C(_07401_),
    .A(net57),
    .Y(_07402_));
 sg13g2_nor4_1 _24033_ (.A(_07389_),
    .B(_07394_),
    .C(_07399_),
    .D(_07402_),
    .Y(_07403_));
 sg13g2_a22oi_1 _24034_ (.Y(_07404_),
    .B1(_06066_),
    .B2(\top_ihp.oisc.regs[11][9] ),
    .A2(net185),
    .A1(\top_ihp.oisc.regs[9][9] ));
 sg13g2_nand2_1 _24035_ (.Y(_07405_),
    .A(\top_ihp.oisc.regs[25][9] ),
    .B(net433));
 sg13g2_nand2_1 _24036_ (.Y(_07406_),
    .A(_07404_),
    .B(_07405_));
 sg13g2_a22oi_1 _24037_ (.Y(_07407_),
    .B1(net204),
    .B2(\top_ihp.oisc.regs[4][9] ),
    .A2(net533),
    .A1(\top_ihp.oisc.regs[22][9] ));
 sg13g2_a22oi_1 _24038_ (.Y(_07408_),
    .B1(_05914_),
    .B2(\top_ihp.oisc.regs[8][9] ),
    .A2(net428),
    .A1(\top_ihp.oisc.regs[15][9] ));
 sg13g2_a22oi_1 _24039_ (.Y(_07409_),
    .B1(net170),
    .B2(\top_ihp.oisc.regs[3][9] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[29][9] ));
 sg13g2_a22oi_1 _24040_ (.Y(_07410_),
    .B1(_05888_),
    .B2(\top_ihp.oisc.regs[12][9] ),
    .A2(net431),
    .A1(\top_ihp.oisc.regs[1][9] ));
 sg13g2_nand4_1 _24041_ (.B(_07408_),
    .C(_07409_),
    .A(_07407_),
    .Y(_07411_),
    .D(_07410_));
 sg13g2_and2_1 _24042_ (.A(\top_ihp.oisc.regs[19][9] ),
    .B(_05551_),
    .X(_07412_));
 sg13g2_a221oi_1 _24043_ (.B2(\top_ihp.oisc.regs[17][9] ),
    .C1(_07412_),
    .B1(_05574_),
    .A1(\top_ihp.oisc.regs[13][9] ),
    .Y(_07413_),
    .A2(net390));
 sg13g2_a22oi_1 _24044_ (.Y(_07414_),
    .B1(_05759_),
    .B2(\top_ihp.oisc.regs[16][9] ),
    .A2(_05565_),
    .A1(\top_ihp.oisc.regs[6][9] ));
 sg13g2_nand3_1 _24045_ (.B(_05388_),
    .C(net724),
    .A(\top_ihp.oisc.regs[5][9] ),
    .Y(_07415_));
 sg13g2_nand3_1 _24046_ (.B(_05667_),
    .C(net749),
    .A(\top_ihp.oisc.regs[2][9] ),
    .Y(_07416_));
 sg13g2_nand2_1 _24047_ (.Y(_07417_),
    .A(\top_ihp.oisc.regs[18][9] ),
    .B(net544));
 sg13g2_and4_1 _24048_ (.A(_07414_),
    .B(_07415_),
    .C(_07416_),
    .D(_07417_),
    .X(_07418_));
 sg13g2_a22oi_1 _24049_ (.Y(_07419_),
    .B1(net408),
    .B2(\top_ihp.oisc.regs[35][9] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[39][9] ));
 sg13g2_a22oi_1 _24050_ (.Y(_07420_),
    .B1(_06637_),
    .B2(\top_ihp.oisc.regs[44][9] ),
    .A2(net347),
    .A1(\top_ihp.oisc.regs[37][9] ));
 sg13g2_nand4_1 _24051_ (.B(_07418_),
    .C(_07419_),
    .A(_07413_),
    .Y(_07421_),
    .D(_07420_));
 sg13g2_and2_1 _24052_ (.A(\top_ihp.oisc.regs[23][9] ),
    .B(_05824_),
    .X(_07422_));
 sg13g2_a221oi_1 _24053_ (.B2(\top_ihp.oisc.regs[21][9] ),
    .C1(_07422_),
    .B1(net663),
    .A1(_08103_),
    .Y(_07423_),
    .A2(net801));
 sg13g2_a22oi_1 _24054_ (.Y(_07424_),
    .B1(net664),
    .B2(\top_ihp.oisc.regs[28][9] ),
    .A2(net546),
    .A1(\top_ihp.oisc.regs[14][9] ));
 sg13g2_mux2_1 _24055_ (.A0(\top_ihp.oisc.regs[26][9] ),
    .A1(\top_ihp.oisc.regs[24][9] ),
    .S(net725),
    .X(_07425_));
 sg13g2_a22oi_1 _24056_ (.Y(_07426_),
    .B1(_06268_),
    .B2(_07425_),
    .A2(net552),
    .A1(\top_ihp.oisc.regs[20][9] ));
 sg13g2_a22oi_1 _24057_ (.Y(_07427_),
    .B1(net537),
    .B2(\top_ihp.oisc.regs[10][9] ),
    .A2(_05429_),
    .A1(\top_ihp.oisc.regs[7][9] ));
 sg13g2_and4_1 _24058_ (.A(_07423_),
    .B(_07424_),
    .C(_07426_),
    .D(_07427_),
    .X(_07428_));
 sg13g2_a22oi_1 _24059_ (.Y(_07429_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[27][9] ),
    .A2(net394),
    .A1(\top_ihp.oisc.regs[45][9] ));
 sg13g2_a22oi_1 _24060_ (.Y(_07430_),
    .B1(net405),
    .B2(\top_ihp.oisc.regs[52][9] ),
    .A2(net421),
    .A1(\top_ihp.oisc.regs[34][9] ));
 sg13g2_nand3_1 _24061_ (.B(_07429_),
    .C(_07430_),
    .A(_07428_),
    .Y(_07431_));
 sg13g2_nor4_1 _24062_ (.A(_07406_),
    .B(_07411_),
    .C(_07421_),
    .D(_07431_),
    .Y(_07432_));
 sg13g2_nand2_1 _24063_ (.Y(_07433_),
    .A(_00213_),
    .B(net59));
 sg13g2_a22oi_1 _24064_ (.Y(_07434_),
    .B1(_05746_),
    .B2(_07433_),
    .A2(net783),
    .A1(_08103_));
 sg13g2_a21oi_1 _24065_ (.A1(_07403_),
    .A2(_07432_),
    .Y(_00419_),
    .B1(_07434_));
 sg13g2_buf_1 _24066_ (.A(net783),
    .X(_07435_));
 sg13g2_nand2_1 _24067_ (.Y(_07436_),
    .A(_07973_),
    .B(_05351_));
 sg13g2_buf_2 _24068_ (.A(_07436_),
    .X(_07437_));
 sg13g2_buf_1 _24069_ (.A(_07437_),
    .X(_07438_));
 sg13g2_or2_1 _24070_ (.X(_07439_),
    .B(_08815_),
    .A(_08810_));
 sg13g2_buf_1 _24071_ (.A(_07439_),
    .X(_07440_));
 sg13g2_nand2_1 _24072_ (.Y(_07441_),
    .A(_08817_),
    .B(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_nor2_1 _24073_ (.A(_07440_),
    .B(_07441_),
    .Y(_07442_));
 sg13g2_buf_1 _24074_ (.A(_07442_),
    .X(_07443_));
 sg13g2_buf_1 _24075_ (.A(_07443_),
    .X(_07444_));
 sg13g2_nand2_1 _24076_ (.Y(_07445_),
    .A(_08813_),
    .B(_08815_));
 sg13g2_nor3_1 _24077_ (.A(_08818_),
    .B(_08817_),
    .C(_07445_),
    .Y(_07446_));
 sg13g2_buf_1 _24078_ (.A(_07446_),
    .X(_07447_));
 sg13g2_buf_1 _24079_ (.A(_07447_),
    .X(_07448_));
 sg13g2_buf_1 _24080_ (.A(net863),
    .X(_07449_));
 sg13g2_nand2_1 _24081_ (.Y(_07450_),
    .A(_08818_),
    .B(\top_ihp.oisc.reg_rb[3] ));
 sg13g2_nand2_2 _24082_ (.Y(_07451_),
    .A(_08810_),
    .B(\top_ihp.oisc.reg_rb[0] ));
 sg13g2_nor2_1 _24083_ (.A(_07450_),
    .B(_07451_),
    .Y(_07452_));
 sg13g2_buf_1 _24084_ (.A(_07452_),
    .X(_07453_));
 sg13g2_buf_2 _24085_ (.A(_07453_),
    .X(_07454_));
 sg13g2_buf_2 _24086_ (.A(net831),
    .X(_07455_));
 sg13g2_a22oi_1 _24087_ (.Y(_07456_),
    .B1(_07455_),
    .B2(\top_ihp.oisc.regs[15][0] ),
    .A2(net846),
    .A1(\top_ihp.oisc.regs[8][0] ));
 sg13g2_or2_1 _24088_ (.X(_07457_),
    .B(_08813_),
    .A(_08814_));
 sg13g2_buf_1 _24089_ (.A(_07457_),
    .X(_07458_));
 sg13g2_nor3_1 _24090_ (.A(_08818_),
    .B(_08817_),
    .C(_07458_),
    .Y(_07459_));
 sg13g2_buf_1 _24091_ (.A(_07459_),
    .X(_07460_));
 sg13g2_buf_1 _24092_ (.A(_07460_),
    .X(_07461_));
 sg13g2_buf_1 _24093_ (.A(net845),
    .X(_07462_));
 sg13g2_nor2_1 _24094_ (.A(_07450_),
    .B(_07458_),
    .Y(_07463_));
 sg13g2_buf_1 _24095_ (.A(_07463_),
    .X(_07464_));
 sg13g2_buf_1 _24096_ (.A(_07464_),
    .X(_07465_));
 sg13g2_a22oi_1 _24097_ (.Y(_07466_),
    .B1(net829),
    .B2(\top_ihp.oisc.regs[14][0] ),
    .A2(net830),
    .A1(\top_ihp.oisc.regs[10][0] ));
 sg13g2_nand2_1 _24098_ (.Y(_07467_),
    .A(_07456_),
    .B(_07466_));
 sg13g2_a21oi_1 _24099_ (.A1(\top_ihp.oisc.regs[5][0] ),
    .A2(net800),
    .Y(_07468_),
    .B1(_07467_));
 sg13g2_nor3_1 _24100_ (.A(\top_ihp.oisc.reg_rb[3] ),
    .B(\top_ihp.oisc.reg_rb[2] ),
    .C(_07440_),
    .Y(_07469_));
 sg13g2_buf_1 _24101_ (.A(_07469_),
    .X(_07470_));
 sg13g2_buf_1 _24102_ (.A(_07470_),
    .X(_07471_));
 sg13g2_nor2_1 _24103_ (.A(_07441_),
    .B(_07451_),
    .Y(_07472_));
 sg13g2_buf_1 _24104_ (.A(_07472_),
    .X(_07473_));
 sg13g2_buf_1 _24105_ (.A(_07473_),
    .X(_07474_));
 sg13g2_buf_1 _24106_ (.A(net798),
    .X(_07475_));
 sg13g2_nor2_1 _24107_ (.A(_07440_),
    .B(_07450_),
    .Y(_07476_));
 sg13g2_buf_2 _24108_ (.A(_07476_),
    .X(_07477_));
 sg13g2_buf_1 _24109_ (.A(_07477_),
    .X(_07478_));
 sg13g2_nor2_1 _24110_ (.A(_07445_),
    .B(_07450_),
    .Y(_07479_));
 sg13g2_buf_1 _24111_ (.A(_07479_),
    .X(_07480_));
 sg13g2_buf_1 _24112_ (.A(_07480_),
    .X(_07481_));
 sg13g2_a22oi_1 _24113_ (.Y(_07482_),
    .B1(net826),
    .B2(\top_ihp.oisc.regs[12][0] ),
    .A2(net827),
    .A1(\top_ihp.oisc.regs[13][0] ));
 sg13g2_nor2_1 _24114_ (.A(net922),
    .B(net1016),
    .Y(_07483_));
 sg13g2_buf_1 _24115_ (.A(_07483_),
    .X(_07484_));
 sg13g2_buf_1 _24116_ (.A(_07484_),
    .X(_07485_));
 sg13g2_nor3_1 _24117_ (.A(_08818_),
    .B(_08817_),
    .C(_07440_),
    .Y(_07486_));
 sg13g2_buf_1 _24118_ (.A(_07486_),
    .X(_07487_));
 sg13g2_buf_1 _24119_ (.A(_07487_),
    .X(_07488_));
 sg13g2_a22oi_1 _24120_ (.Y(_07489_),
    .B1(net844),
    .B2(\top_ihp.oisc.regs[9][0] ),
    .A2(net862),
    .A1(\top_ihp.oisc.regs[32][0] ));
 sg13g2_nor3_1 _24121_ (.A(_08818_),
    .B(_08817_),
    .C(_07451_),
    .Y(_07490_));
 sg13g2_buf_2 _24122_ (.A(_07490_),
    .X(_07491_));
 sg13g2_buf_1 _24123_ (.A(_07491_),
    .X(_07492_));
 sg13g2_buf_2 _24124_ (.A(net843),
    .X(_07493_));
 sg13g2_nor4_1 _24125_ (.A(_08818_),
    .B(\top_ihp.oisc.micro_op[11] ),
    .C(_08814_),
    .D(_08810_),
    .Y(_07494_));
 sg13g2_and2_1 _24126_ (.A(net1016),
    .B(_07494_),
    .X(_07495_));
 sg13g2_buf_1 _24127_ (.A(_07495_),
    .X(_07496_));
 sg13g2_buf_1 _24128_ (.A(_07496_),
    .X(_07497_));
 sg13g2_buf_1 _24129_ (.A(net893),
    .X(_07498_));
 sg13g2_a22oi_1 _24130_ (.Y(_07499_),
    .B1(net885),
    .B2(\top_ihp.oisc.regs[0][0] ),
    .A2(net825),
    .A1(\top_ihp.oisc.regs[11][0] ));
 sg13g2_nand3_1 _24131_ (.B(_07489_),
    .C(_07499_),
    .A(_07482_),
    .Y(_07500_));
 sg13g2_a221oi_1 _24132_ (.B2(\top_ihp.oisc.regs[7][0] ),
    .C1(_07500_),
    .B1(net773),
    .A1(\top_ihp.oisc.regs[1][0] ),
    .Y(_07501_),
    .A2(net828));
 sg13g2_nor2_1 _24133_ (.A(_07441_),
    .B(_07458_),
    .Y(_07502_));
 sg13g2_buf_2 _24134_ (.A(_07502_),
    .X(_07503_));
 sg13g2_buf_1 _24135_ (.A(_07503_),
    .X(_07504_));
 sg13g2_buf_1 _24136_ (.A(net797),
    .X(_07505_));
 sg13g2_nor3_1 _24137_ (.A(\top_ihp.oisc.reg_rb[3] ),
    .B(\top_ihp.oisc.reg_rb[2] ),
    .C(_07451_),
    .Y(_07506_));
 sg13g2_buf_2 _24138_ (.A(_07506_),
    .X(_07507_));
 sg13g2_buf_1 _24139_ (.A(_07507_),
    .X(_07508_));
 sg13g2_a22oi_1 _24140_ (.Y(_07509_),
    .B1(net824),
    .B2(\top_ihp.oisc.regs[3][0] ),
    .A2(net772),
    .A1(\top_ihp.oisc.regs[6][0] ));
 sg13g2_nor3_1 _24141_ (.A(\top_ihp.oisc.reg_rb[3] ),
    .B(\top_ihp.oisc.reg_rb[2] ),
    .C(_07458_),
    .Y(_07510_));
 sg13g2_buf_1 _24142_ (.A(_07510_),
    .X(_07511_));
 sg13g2_buf_1 _24143_ (.A(_07511_),
    .X(_07512_));
 sg13g2_nor2_1 _24144_ (.A(_07441_),
    .B(_07445_),
    .Y(_07513_));
 sg13g2_buf_1 _24145_ (.A(_07513_),
    .X(_07514_));
 sg13g2_buf_1 _24146_ (.A(_07514_),
    .X(_07515_));
 sg13g2_a22oi_1 _24147_ (.Y(_07516_),
    .B1(net796),
    .B2(\top_ihp.oisc.regs[4][0] ),
    .A2(net823),
    .A1(\top_ihp.oisc.regs[2][0] ));
 sg13g2_nand4_1 _24148_ (.B(_07501_),
    .C(_07509_),
    .A(_07468_),
    .Y(_07517_),
    .D(_07516_));
 sg13g2_buf_1 _24149_ (.A(net783),
    .X(_07518_));
 sg13g2_a21oi_1 _24150_ (.A1(net864),
    .A2(_07517_),
    .Y(_07519_),
    .B1(net744));
 sg13g2_a21oi_1 _24151_ (.A1(_08459_),
    .A2(net745),
    .Y(_00420_),
    .B1(_07519_));
 sg13g2_buf_1 _24152_ (.A(_07487_),
    .X(_07520_));
 sg13g2_a22oi_1 _24153_ (.Y(_07521_),
    .B1(net842),
    .B2(\top_ihp.oisc.regs[9][10] ),
    .A2(net846),
    .A1(\top_ihp.oisc.regs[8][10] ));
 sg13g2_a22oi_1 _24154_ (.Y(_07522_),
    .B1(net830),
    .B2(\top_ihp.oisc.regs[10][10] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[15][10] ));
 sg13g2_nand2_1 _24155_ (.Y(_07523_),
    .A(_07521_),
    .B(_07522_));
 sg13g2_a21oi_1 _24156_ (.A1(\top_ihp.oisc.regs[7][10] ),
    .A2(net773),
    .Y(_07524_),
    .B1(_07523_));
 sg13g2_buf_1 _24157_ (.A(_07464_),
    .X(_07525_));
 sg13g2_a22oi_1 _24158_ (.Y(_07526_),
    .B1(net826),
    .B2(\top_ihp.oisc.regs[12][10] ),
    .A2(net822),
    .A1(\top_ihp.oisc.regs[14][10] ));
 sg13g2_a22oi_1 _24159_ (.Y(_07527_),
    .B1(net825),
    .B2(\top_ihp.oisc.regs[11][10] ),
    .A2(net862),
    .A1(\top_ihp.oisc.regs[32][10] ));
 sg13g2_a22oi_1 _24160_ (.Y(_07528_),
    .B1(net885),
    .B2(_05852_),
    .A2(_07477_),
    .A1(\top_ihp.oisc.regs[13][10] ));
 sg13g2_nand3_1 _24161_ (.B(_07527_),
    .C(_07528_),
    .A(_07526_),
    .Y(_07529_));
 sg13g2_a221oi_1 _24162_ (.B2(\top_ihp.oisc.regs[3][10] ),
    .C1(_07529_),
    .B1(net824),
    .A1(\top_ihp.oisc.regs[1][10] ),
    .Y(_07530_),
    .A2(net828));
 sg13g2_buf_1 _24163_ (.A(_07504_),
    .X(_07531_));
 sg13g2_buf_1 _24164_ (.A(_07511_),
    .X(_07532_));
 sg13g2_a22oi_1 _24165_ (.Y(_07533_),
    .B1(net821),
    .B2(\top_ihp.oisc.regs[2][10] ),
    .A2(net771),
    .A1(\top_ihp.oisc.regs[6][10] ));
 sg13g2_buf_1 _24166_ (.A(_07443_),
    .X(_07534_));
 sg13g2_a22oi_1 _24167_ (.Y(_07535_),
    .B1(net796),
    .B2(\top_ihp.oisc.regs[4][10] ),
    .A2(net795),
    .A1(\top_ihp.oisc.regs[5][10] ));
 sg13g2_nand4_1 _24168_ (.B(_07530_),
    .C(_07533_),
    .A(_07524_),
    .Y(_07536_),
    .D(_07535_));
 sg13g2_buf_1 _24169_ (.A(net783),
    .X(_07537_));
 sg13g2_a21oi_1 _24170_ (.A1(net864),
    .A2(_07536_),
    .Y(_07538_),
    .B1(net743));
 sg13g2_a21oi_1 _24171_ (.A1(_08414_),
    .A2(net745),
    .Y(_00421_),
    .B1(_07538_));
 sg13g2_buf_1 _24172_ (.A(net885),
    .X(_07539_));
 sg13g2_buf_1 _24173_ (.A(_07443_),
    .X(_07540_));
 sg13g2_buf_1 _24174_ (.A(_07514_),
    .X(_07541_));
 sg13g2_buf_1 _24175_ (.A(_07470_),
    .X(_07542_));
 sg13g2_and2_1 _24176_ (.A(\top_ihp.oisc.regs[1][11] ),
    .B(net820),
    .X(_07543_));
 sg13g2_a221oi_1 _24177_ (.B2(\top_ihp.oisc.regs[4][11] ),
    .C1(_07543_),
    .B1(net793),
    .A1(\top_ihp.oisc.regs[5][11] ),
    .Y(_07544_),
    .A2(net794));
 sg13g2_nor3_1 _24178_ (.A(\top_ihp.oisc.reg_rb[3] ),
    .B(\top_ihp.oisc.reg_rb[2] ),
    .C(_07451_),
    .Y(_07545_));
 sg13g2_buf_2 _24179_ (.A(_07545_),
    .X(_07546_));
 sg13g2_buf_1 _24180_ (.A(_07546_),
    .X(_07547_));
 sg13g2_buf_1 _24181_ (.A(_07480_),
    .X(_07548_));
 sg13g2_buf_1 _24182_ (.A(_07487_),
    .X(_07549_));
 sg13g2_buf_1 _24183_ (.A(_07453_),
    .X(_07550_));
 sg13g2_a21oi_1 _24184_ (.A1(\top_ihp.oisc.regs[15][11] ),
    .A2(net817),
    .Y(_07551_),
    .B1(net893));
 sg13g2_a22oi_1 _24185_ (.Y(_07552_),
    .B1(net843),
    .B2(\top_ihp.oisc.regs[11][11] ),
    .A2(net845),
    .A1(\top_ihp.oisc.regs[10][11] ));
 sg13g2_nand2_1 _24186_ (.Y(_07553_),
    .A(_07551_),
    .B(_07552_));
 sg13g2_a221oi_1 _24187_ (.B2(\top_ihp.oisc.regs[9][11] ),
    .C1(_07553_),
    .B1(net841),
    .A1(\top_ihp.oisc.regs[12][11] ),
    .Y(_07554_),
    .A2(net818));
 sg13g2_buf_1 _24188_ (.A(_07484_),
    .X(_07555_));
 sg13g2_buf_1 _24189_ (.A(_07477_),
    .X(_07556_));
 sg13g2_a22oi_1 _24190_ (.Y(_07557_),
    .B1(net816),
    .B2(\top_ihp.oisc.regs[13][11] ),
    .A2(net860),
    .A1(\top_ihp.oisc.regs[32][11] ));
 sg13g2_a22oi_1 _24191_ (.Y(_07558_),
    .B1(net829),
    .B2(\top_ihp.oisc.regs[14][11] ),
    .A2(net846),
    .A1(\top_ihp.oisc.regs[8][11] ));
 sg13g2_buf_1 _24192_ (.A(_07473_),
    .X(_07559_));
 sg13g2_a22oi_1 _24193_ (.Y(_07560_),
    .B1(net797),
    .B2(\top_ihp.oisc.regs[6][11] ),
    .A2(net792),
    .A1(\top_ihp.oisc.regs[7][11] ));
 sg13g2_nand4_1 _24194_ (.B(_07557_),
    .C(_07558_),
    .A(_07554_),
    .Y(_07561_),
    .D(_07560_));
 sg13g2_a221oi_1 _24195_ (.B2(\top_ihp.oisc.regs[3][11] ),
    .C1(_07561_),
    .B1(net819),
    .A1(\top_ihp.oisc.regs[2][11] ),
    .Y(_07562_),
    .A2(net821));
 sg13g2_buf_1 _24196_ (.A(_07555_),
    .X(_07563_));
 sg13g2_a221oi_1 _24197_ (.B2(_07562_),
    .C1(net840),
    .B1(_07544_),
    .A1(_00215_),
    .Y(_07564_),
    .A2(net861));
 sg13g2_buf_1 _24198_ (.A(net804),
    .X(_07565_));
 sg13g2_mux2_1 _24199_ (.A0(_08028_),
    .A1(_07564_),
    .S(net770),
    .X(_00422_));
 sg13g2_a22oi_1 _24200_ (.Y(_07566_),
    .B1(net816),
    .B2(\top_ihp.oisc.regs[13][12] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[15][12] ));
 sg13g2_a22oi_1 _24201_ (.Y(_07567_),
    .B1(net842),
    .B2(\top_ihp.oisc.regs[9][12] ),
    .A2(net830),
    .A1(\top_ihp.oisc.regs[10][12] ));
 sg13g2_nand2_1 _24202_ (.Y(_07568_),
    .A(_07566_),
    .B(_07567_));
 sg13g2_a21oi_1 _24203_ (.A1(\top_ihp.oisc.regs[7][12] ),
    .A2(net773),
    .Y(_07569_),
    .B1(_07568_));
 sg13g2_buf_1 _24204_ (.A(_07511_),
    .X(_07570_));
 sg13g2_a22oi_1 _24205_ (.Y(_07571_),
    .B1(net826),
    .B2(\top_ihp.oisc.regs[12][12] ),
    .A2(net862),
    .A1(\top_ihp.oisc.regs[32][12] ));
 sg13g2_a22oi_1 _24206_ (.Y(_07572_),
    .B1(net825),
    .B2(\top_ihp.oisc.regs[11][12] ),
    .A2(_07448_),
    .A1(\top_ihp.oisc.regs[8][12] ));
 sg13g2_inv_1 _24207_ (.Y(_07573_),
    .A(_00216_));
 sg13g2_a22oi_1 _24208_ (.Y(_07574_),
    .B1(net885),
    .B2(_07573_),
    .A2(net822),
    .A1(\top_ihp.oisc.regs[14][12] ));
 sg13g2_nand3_1 _24209_ (.B(_07572_),
    .C(_07574_),
    .A(_07571_),
    .Y(_07575_));
 sg13g2_a221oi_1 _24210_ (.B2(\top_ihp.oisc.regs[2][12] ),
    .C1(_07575_),
    .B1(net815),
    .A1(\top_ihp.oisc.regs[3][12] ),
    .Y(_07576_),
    .A2(_07507_));
 sg13g2_buf_1 _24211_ (.A(_07470_),
    .X(_07577_));
 sg13g2_a22oi_1 _24212_ (.Y(_07578_),
    .B1(net772),
    .B2(\top_ihp.oisc.regs[6][12] ),
    .A2(net814),
    .A1(\top_ihp.oisc.regs[1][12] ));
 sg13g2_a22oi_1 _24213_ (.Y(_07579_),
    .B1(net796),
    .B2(\top_ihp.oisc.regs[4][12] ),
    .A2(net795),
    .A1(\top_ihp.oisc.regs[5][12] ));
 sg13g2_nand4_1 _24214_ (.B(_07576_),
    .C(_07578_),
    .A(_07569_),
    .Y(_07580_),
    .D(_07579_));
 sg13g2_a21oi_1 _24215_ (.A1(net864),
    .A2(_07580_),
    .Y(_07581_),
    .B1(net743));
 sg13g2_a21oi_1 _24216_ (.A1(_04594_),
    .A2(net745),
    .Y(_00423_),
    .B1(_07581_));
 sg13g2_and2_1 _24217_ (.A(\top_ihp.oisc.regs[1][13] ),
    .B(net820),
    .X(_07582_));
 sg13g2_a221oi_1 _24218_ (.B2(\top_ihp.oisc.regs[4][13] ),
    .C1(_07582_),
    .B1(net793),
    .A1(\top_ihp.oisc.regs[5][13] ),
    .Y(_07583_),
    .A2(net794));
 sg13g2_a21oi_1 _24219_ (.A1(\top_ihp.oisc.regs[15][13] ),
    .A2(net817),
    .Y(_07584_),
    .B1(net893));
 sg13g2_a22oi_1 _24220_ (.Y(_07585_),
    .B1(net843),
    .B2(\top_ihp.oisc.regs[11][13] ),
    .A2(net845),
    .A1(\top_ihp.oisc.regs[10][13] ));
 sg13g2_nand2_1 _24221_ (.Y(_07586_),
    .A(_07584_),
    .B(_07585_));
 sg13g2_a221oi_1 _24222_ (.B2(\top_ihp.oisc.regs[9][13] ),
    .C1(_07586_),
    .B1(net841),
    .A1(\top_ihp.oisc.regs[12][13] ),
    .Y(_07587_),
    .A2(net818));
 sg13g2_a22oi_1 _24223_ (.Y(_07588_),
    .B1(net816),
    .B2(\top_ihp.oisc.regs[13][13] ),
    .A2(net860),
    .A1(\top_ihp.oisc.regs[32][13] ));
 sg13g2_a22oi_1 _24224_ (.Y(_07589_),
    .B1(net829),
    .B2(\top_ihp.oisc.regs[14][13] ),
    .A2(net846),
    .A1(\top_ihp.oisc.regs[8][13] ));
 sg13g2_a22oi_1 _24225_ (.Y(_07590_),
    .B1(net797),
    .B2(\top_ihp.oisc.regs[6][13] ),
    .A2(net792),
    .A1(\top_ihp.oisc.regs[7][13] ));
 sg13g2_nand4_1 _24226_ (.B(_07588_),
    .C(_07589_),
    .A(_07587_),
    .Y(_07591_),
    .D(_07590_));
 sg13g2_a221oi_1 _24227_ (.B2(\top_ihp.oisc.regs[3][13] ),
    .C1(_07591_),
    .B1(net819),
    .A1(\top_ihp.oisc.regs[2][13] ),
    .Y(_07592_),
    .A2(net821));
 sg13g2_a221oi_1 _24228_ (.B2(_07592_),
    .C1(net840),
    .B1(_07583_),
    .A1(_00217_),
    .Y(_07593_),
    .A2(net861));
 sg13g2_mux2_1 _24229_ (.A0(_08050_),
    .A1(_07593_),
    .S(net770),
    .X(_00424_));
 sg13g2_a22oi_1 _24230_ (.Y(_07594_),
    .B1(net826),
    .B2(\top_ihp.oisc.regs[12][14] ),
    .A2(net846),
    .A1(\top_ihp.oisc.regs[8][14] ));
 sg13g2_buf_1 _24231_ (.A(_07477_),
    .X(_07595_));
 sg13g2_a22oi_1 _24232_ (.Y(_07596_),
    .B1(net842),
    .B2(\top_ihp.oisc.regs[9][14] ),
    .A2(net813),
    .A1(\top_ihp.oisc.regs[13][14] ));
 sg13g2_nand2_1 _24233_ (.Y(_07597_),
    .A(_07594_),
    .B(_07596_));
 sg13g2_a21oi_1 _24234_ (.A1(\top_ihp.oisc.regs[5][14] ),
    .A2(net800),
    .Y(_07598_),
    .B1(_07597_));
 sg13g2_buf_2 _24235_ (.A(net843),
    .X(_07599_));
 sg13g2_a22oi_1 _24236_ (.Y(_07600_),
    .B1(net812),
    .B2(\top_ihp.oisc.regs[11][14] ),
    .A2(net822),
    .A1(\top_ihp.oisc.regs[14][14] ));
 sg13g2_a22oi_1 _24237_ (.Y(_07601_),
    .B1(net799),
    .B2(\top_ihp.oisc.regs[15][14] ),
    .A2(net862),
    .A1(\top_ihp.oisc.regs[32][14] ));
 sg13g2_buf_1 _24238_ (.A(_07460_),
    .X(_07602_));
 sg13g2_buf_1 _24239_ (.A(_07497_),
    .X(_07603_));
 sg13g2_a22oi_1 _24240_ (.Y(_07604_),
    .B1(net884),
    .B2(_06136_),
    .A2(net839),
    .A1(\top_ihp.oisc.regs[10][14] ));
 sg13g2_nand3_1 _24241_ (.B(_07601_),
    .C(_07604_),
    .A(_07600_),
    .Y(_07605_));
 sg13g2_a221oi_1 _24242_ (.B2(\top_ihp.oisc.regs[7][14] ),
    .C1(_07605_),
    .B1(net773),
    .A1(\top_ihp.oisc.regs[1][14] ),
    .Y(_07606_),
    .A2(net828));
 sg13g2_a22oi_1 _24243_ (.Y(_07607_),
    .B1(net824),
    .B2(\top_ihp.oisc.regs[3][14] ),
    .A2(net771),
    .A1(\top_ihp.oisc.regs[6][14] ));
 sg13g2_a22oi_1 _24244_ (.Y(_07608_),
    .B1(net796),
    .B2(\top_ihp.oisc.regs[4][14] ),
    .A2(net823),
    .A1(\top_ihp.oisc.regs[2][14] ));
 sg13g2_nand4_1 _24245_ (.B(_07606_),
    .C(_07607_),
    .A(_07598_),
    .Y(_07609_),
    .D(_07608_));
 sg13g2_a21oi_1 _24246_ (.A1(net864),
    .A2(_07609_),
    .Y(_07610_),
    .B1(net743));
 sg13g2_a21oi_1 _24247_ (.A1(_08231_),
    .A2(net745),
    .Y(_00425_),
    .B1(_07610_));
 sg13g2_and2_1 _24248_ (.A(\top_ihp.oisc.regs[1][15] ),
    .B(net820),
    .X(_07611_));
 sg13g2_a221oi_1 _24249_ (.B2(\top_ihp.oisc.regs[4][15] ),
    .C1(_07611_),
    .B1(net793),
    .A1(\top_ihp.oisc.regs[5][15] ),
    .Y(_07612_),
    .A2(net794));
 sg13g2_a21oi_1 _24250_ (.A1(\top_ihp.oisc.regs[14][15] ),
    .A2(_07464_),
    .Y(_07613_),
    .B1(net893));
 sg13g2_a22oi_1 _24251_ (.Y(_07614_),
    .B1(_07480_),
    .B2(\top_ihp.oisc.regs[12][15] ),
    .A2(net845),
    .A1(\top_ihp.oisc.regs[10][15] ));
 sg13g2_nand2_1 _24252_ (.Y(_07615_),
    .A(_07613_),
    .B(_07614_));
 sg13g2_a221oi_1 _24253_ (.B2(\top_ihp.oisc.regs[9][15] ),
    .C1(_07615_),
    .B1(net841),
    .A1(\top_ihp.oisc.regs[15][15] ),
    .Y(_07616_),
    .A2(net831));
 sg13g2_a22oi_1 _24254_ (.Y(_07617_),
    .B1(net816),
    .B2(\top_ihp.oisc.regs[13][15] ),
    .A2(net860),
    .A1(\top_ihp.oisc.regs[32][15] ));
 sg13g2_a22oi_1 _24255_ (.Y(_07618_),
    .B1(net812),
    .B2(\top_ihp.oisc.regs[11][15] ),
    .A2(net846),
    .A1(\top_ihp.oisc.regs[8][15] ));
 sg13g2_a22oi_1 _24256_ (.Y(_07619_),
    .B1(net797),
    .B2(\top_ihp.oisc.regs[6][15] ),
    .A2(net792),
    .A1(\top_ihp.oisc.regs[7][15] ));
 sg13g2_nand4_1 _24257_ (.B(_07617_),
    .C(_07618_),
    .A(_07616_),
    .Y(_07620_),
    .D(_07619_));
 sg13g2_a221oi_1 _24258_ (.B2(\top_ihp.oisc.regs[3][15] ),
    .C1(_07620_),
    .B1(net819),
    .A1(\top_ihp.oisc.regs[2][15] ),
    .Y(_07621_),
    .A2(net821));
 sg13g2_a221oi_1 _24259_ (.B2(_07621_),
    .C1(net840),
    .B1(_07612_),
    .A1(_00219_),
    .Y(_07622_),
    .A2(net861));
 sg13g2_mux2_1 _24260_ (.A0(_08009_),
    .A1(_07622_),
    .S(net770),
    .X(_00426_));
 sg13g2_a22oi_1 _24261_ (.Y(_07623_),
    .B1(_07556_),
    .B2(\top_ihp.oisc.regs[13][16] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[15][16] ));
 sg13g2_a22oi_1 _24262_ (.Y(_07624_),
    .B1(net829),
    .B2(\top_ihp.oisc.regs[14][16] ),
    .A2(net846),
    .A1(\top_ihp.oisc.regs[8][16] ));
 sg13g2_nand2_1 _24263_ (.Y(_07625_),
    .A(_07623_),
    .B(_07624_));
 sg13g2_a21oi_1 _24264_ (.A1(\top_ihp.oisc.regs[5][16] ),
    .A2(net800),
    .Y(_07626_),
    .B1(_07625_));
 sg13g2_a22oi_1 _24265_ (.Y(_07627_),
    .B1(net826),
    .B2(\top_ihp.oisc.regs[12][16] ),
    .A2(net839),
    .A1(\top_ihp.oisc.regs[10][16] ));
 sg13g2_buf_1 _24266_ (.A(_07484_),
    .X(_07628_));
 sg13g2_a22oi_1 _24267_ (.Y(_07629_),
    .B1(net844),
    .B2(\top_ihp.oisc.regs[9][16] ),
    .A2(net859),
    .A1(\top_ihp.oisc.regs[32][16] ));
 sg13g2_a22oi_1 _24268_ (.Y(_07630_),
    .B1(net884),
    .B2(_06250_),
    .A2(net825),
    .A1(\top_ihp.oisc.regs[11][16] ));
 sg13g2_nand3_1 _24269_ (.B(_07629_),
    .C(_07630_),
    .A(_07627_),
    .Y(_07631_));
 sg13g2_a221oi_1 _24270_ (.B2(\top_ihp.oisc.regs[7][16] ),
    .C1(_07631_),
    .B1(net773),
    .A1(\top_ihp.oisc.regs[1][16] ),
    .Y(_07632_),
    .A2(net828));
 sg13g2_a22oi_1 _24271_ (.Y(_07633_),
    .B1(net824),
    .B2(\top_ihp.oisc.regs[3][16] ),
    .A2(net771),
    .A1(\top_ihp.oisc.regs[6][16] ));
 sg13g2_buf_1 _24272_ (.A(_07514_),
    .X(_07634_));
 sg13g2_a22oi_1 _24273_ (.Y(_07635_),
    .B1(net791),
    .B2(\top_ihp.oisc.regs[4][16] ),
    .A2(net815),
    .A1(\top_ihp.oisc.regs[2][16] ));
 sg13g2_nand4_1 _24274_ (.B(_07632_),
    .C(_07633_),
    .A(_07626_),
    .Y(_07636_),
    .D(_07635_));
 sg13g2_a21oi_1 _24275_ (.A1(net864),
    .A2(_07636_),
    .Y(_07637_),
    .B1(net743));
 sg13g2_a21oi_1 _24276_ (.A1(_08022_),
    .A2(net745),
    .Y(_00427_),
    .B1(_07637_));
 sg13g2_and2_1 _24277_ (.A(\top_ihp.oisc.regs[1][17] ),
    .B(net820),
    .X(_07638_));
 sg13g2_a221oi_1 _24278_ (.B2(\top_ihp.oisc.regs[4][17] ),
    .C1(_07638_),
    .B1(net793),
    .A1(\top_ihp.oisc.regs[5][17] ),
    .Y(_07639_),
    .A2(net794));
 sg13g2_a21oi_1 _24279_ (.A1(\top_ihp.oisc.regs[9][17] ),
    .A2(_07487_),
    .Y(_07640_),
    .B1(net893));
 sg13g2_a22oi_1 _24280_ (.Y(_07641_),
    .B1(net845),
    .B2(\top_ihp.oisc.regs[10][17] ),
    .A2(_07453_),
    .A1(\top_ihp.oisc.regs[15][17] ));
 sg13g2_nand2_1 _24281_ (.Y(_07642_),
    .A(_07640_),
    .B(_07641_));
 sg13g2_a221oi_1 _24282_ (.B2(\top_ihp.oisc.regs[12][17] ),
    .C1(_07642_),
    .B1(net826),
    .A1(\top_ihp.oisc.regs[8][17] ),
    .Y(_07643_),
    .A2(net863));
 sg13g2_buf_1 _24283_ (.A(net859),
    .X(_07644_));
 sg13g2_a22oi_1 _24284_ (.Y(_07645_),
    .B1(net813),
    .B2(\top_ihp.oisc.regs[13][17] ),
    .A2(net838),
    .A1(\top_ihp.oisc.regs[32][17] ));
 sg13g2_a22oi_1 _24285_ (.Y(_07646_),
    .B1(net812),
    .B2(\top_ihp.oisc.regs[11][17] ),
    .A2(net822),
    .A1(\top_ihp.oisc.regs[14][17] ));
 sg13g2_a22oi_1 _24286_ (.Y(_07647_),
    .B1(net797),
    .B2(\top_ihp.oisc.regs[6][17] ),
    .A2(net792),
    .A1(\top_ihp.oisc.regs[7][17] ));
 sg13g2_nand4_1 _24287_ (.B(_07645_),
    .C(_07646_),
    .A(_07643_),
    .Y(_07648_),
    .D(_07647_));
 sg13g2_a221oi_1 _24288_ (.B2(\top_ihp.oisc.regs[3][17] ),
    .C1(_07648_),
    .B1(net819),
    .A1(\top_ihp.oisc.regs[2][17] ),
    .Y(_07649_),
    .A2(net821));
 sg13g2_a221oi_1 _24289_ (.B2(_07649_),
    .C1(net840),
    .B1(_07639_),
    .A1(_00221_),
    .Y(_07650_),
    .A2(net861));
 sg13g2_mux2_1 _24290_ (.A0(_08006_),
    .A1(_07650_),
    .S(net770),
    .X(_00428_));
 sg13g2_a22oi_1 _24291_ (.Y(_07651_),
    .B1(net816),
    .B2(\top_ihp.oisc.regs[13][18] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[15][18] ));
 sg13g2_a22oi_1 _24292_ (.Y(_07652_),
    .B1(net829),
    .B2(\top_ihp.oisc.regs[14][18] ),
    .A2(net830),
    .A1(\top_ihp.oisc.regs[10][18] ));
 sg13g2_nand2_1 _24293_ (.Y(_07653_),
    .A(_07651_),
    .B(_07652_));
 sg13g2_a21oi_1 _24294_ (.A1(\top_ihp.oisc.regs[7][18] ),
    .A2(net773),
    .Y(_07654_),
    .B1(_07653_));
 sg13g2_a22oi_1 _24295_ (.Y(_07655_),
    .B1(net818),
    .B2(\top_ihp.oisc.regs[12][18] ),
    .A2(net863),
    .A1(\top_ihp.oisc.regs[8][18] ));
 sg13g2_a22oi_1 _24296_ (.Y(_07656_),
    .B1(net844),
    .B2(\top_ihp.oisc.regs[9][18] ),
    .A2(net859),
    .A1(\top_ihp.oisc.regs[32][18] ));
 sg13g2_inv_1 _24297_ (.Y(_07657_),
    .A(_00222_));
 sg13g2_a22oi_1 _24298_ (.Y(_07658_),
    .B1(net884),
    .B2(_07657_),
    .A2(net825),
    .A1(\top_ihp.oisc.regs[11][18] ));
 sg13g2_nand3_1 _24299_ (.B(_07656_),
    .C(_07658_),
    .A(_07655_),
    .Y(_07659_));
 sg13g2_a221oi_1 _24300_ (.B2(\top_ihp.oisc.regs[3][18] ),
    .C1(_07659_),
    .B1(_07507_),
    .A1(\top_ihp.oisc.regs[1][18] ),
    .Y(_07660_),
    .A2(net828));
 sg13g2_a22oi_1 _24301_ (.Y(_07661_),
    .B1(net821),
    .B2(\top_ihp.oisc.regs[2][18] ),
    .A2(net771),
    .A1(\top_ihp.oisc.regs[6][18] ));
 sg13g2_a22oi_1 _24302_ (.Y(_07662_),
    .B1(net791),
    .B2(\top_ihp.oisc.regs[4][18] ),
    .A2(net795),
    .A1(\top_ihp.oisc.regs[5][18] ));
 sg13g2_nand4_1 _24303_ (.B(_07660_),
    .C(_07661_),
    .A(_07654_),
    .Y(_07663_),
    .D(_07662_));
 sg13g2_a21oi_1 _24304_ (.A1(net864),
    .A2(_07663_),
    .Y(_07664_),
    .B1(net743));
 sg13g2_a21oi_1 _24305_ (.A1(_08258_),
    .A2(net745),
    .Y(_00429_),
    .B1(_07664_));
 sg13g2_and2_1 _24306_ (.A(\top_ihp.oisc.regs[1][19] ),
    .B(net820),
    .X(_07665_));
 sg13g2_a221oi_1 _24307_ (.B2(\top_ihp.oisc.regs[4][19] ),
    .C1(_07665_),
    .B1(net793),
    .A1(\top_ihp.oisc.regs[5][19] ),
    .Y(_07666_),
    .A2(net794));
 sg13g2_a21oi_1 _24308_ (.A1(\top_ihp.oisc.regs[8][19] ),
    .A2(_07447_),
    .Y(_07667_),
    .B1(net893));
 sg13g2_a22oi_1 _24309_ (.Y(_07668_),
    .B1(_07480_),
    .B2(\top_ihp.oisc.regs[12][19] ),
    .A2(_07453_),
    .A1(\top_ihp.oisc.regs[15][19] ));
 sg13g2_nand2_1 _24310_ (.Y(_07669_),
    .A(_07667_),
    .B(_07668_));
 sg13g2_a221oi_1 _24311_ (.B2(\top_ihp.oisc.regs[9][19] ),
    .C1(_07669_),
    .B1(net841),
    .A1(\top_ihp.oisc.regs[13][19] ),
    .Y(_07670_),
    .A2(net827));
 sg13g2_a22oi_1 _24312_ (.Y(_07671_),
    .B1(net829),
    .B2(\top_ihp.oisc.regs[14][19] ),
    .A2(net838),
    .A1(\top_ihp.oisc.regs[32][19] ));
 sg13g2_a22oi_1 _24313_ (.Y(_07672_),
    .B1(net812),
    .B2(\top_ihp.oisc.regs[11][19] ),
    .A2(net830),
    .A1(\top_ihp.oisc.regs[10][19] ));
 sg13g2_a22oi_1 _24314_ (.Y(_07673_),
    .B1(net797),
    .B2(\top_ihp.oisc.regs[6][19] ),
    .A2(net792),
    .A1(\top_ihp.oisc.regs[7][19] ));
 sg13g2_nand4_1 _24315_ (.B(_07671_),
    .C(_07672_),
    .A(_07670_),
    .Y(_07674_),
    .D(_07673_));
 sg13g2_a221oi_1 _24316_ (.B2(\top_ihp.oisc.regs[3][19] ),
    .C1(_07674_),
    .B1(net819),
    .A1(\top_ihp.oisc.regs[2][19] ),
    .Y(_07675_),
    .A2(net821));
 sg13g2_a221oi_1 _24317_ (.B2(_07675_),
    .C1(net840),
    .B1(_07666_),
    .A1(_00223_),
    .Y(_07676_),
    .A2(net861));
 sg13g2_mux2_1 _24318_ (.A0(net1071),
    .A1(_07676_),
    .S(net770),
    .X(_00430_));
 sg13g2_buf_1 _24319_ (.A(_07464_),
    .X(_07677_));
 sg13g2_a22oi_1 _24320_ (.Y(_07678_),
    .B1(net812),
    .B2(\top_ihp.oisc.regs[11][1] ),
    .A2(_07677_),
    .A1(\top_ihp.oisc.regs[14][1] ));
 sg13g2_a22oi_1 _24321_ (.Y(_07679_),
    .B1(net842),
    .B2(\top_ihp.oisc.regs[9][1] ),
    .A2(net813),
    .A1(\top_ihp.oisc.regs[13][1] ));
 sg13g2_nand2_1 _24322_ (.Y(_07680_),
    .A(_07678_),
    .B(_07679_));
 sg13g2_a21oi_1 _24323_ (.A1(\top_ihp.oisc.regs[7][1] ),
    .A2(net773),
    .Y(_07681_),
    .B1(_07680_));
 sg13g2_buf_1 _24324_ (.A(_07447_),
    .X(_07682_));
 sg13g2_a22oi_1 _24325_ (.Y(_07683_),
    .B1(net858),
    .B2(\top_ihp.oisc.regs[8][1] ),
    .A2(net862),
    .A1(\top_ihp.oisc.regs[32][1] ));
 sg13g2_a22oi_1 _24326_ (.Y(_07684_),
    .B1(net818),
    .B2(\top_ihp.oisc.regs[12][1] ),
    .A2(net831),
    .A1(\top_ihp.oisc.regs[15][1] ));
 sg13g2_a22oi_1 _24327_ (.Y(_07685_),
    .B1(net884),
    .B2(_06452_),
    .A2(net839),
    .A1(\top_ihp.oisc.regs[10][1] ));
 sg13g2_nand3_1 _24328_ (.B(_07684_),
    .C(_07685_),
    .A(_07683_),
    .Y(_07686_));
 sg13g2_a221oi_1 _24329_ (.B2(\top_ihp.oisc.regs[2][1] ),
    .C1(_07686_),
    .B1(net815),
    .A1(\top_ihp.oisc.regs[3][1] ),
    .Y(_07687_),
    .A2(_07507_));
 sg13g2_a22oi_1 _24330_ (.Y(_07688_),
    .B1(net772),
    .B2(\top_ihp.oisc.regs[6][1] ),
    .A2(net814),
    .A1(\top_ihp.oisc.regs[1][1] ));
 sg13g2_a22oi_1 _24331_ (.Y(_07689_),
    .B1(net791),
    .B2(\top_ihp.oisc.regs[4][1] ),
    .A2(net795),
    .A1(\top_ihp.oisc.regs[5][1] ));
 sg13g2_nand4_1 _24332_ (.B(_07687_),
    .C(_07688_),
    .A(_07681_),
    .Y(_07690_),
    .D(_07689_));
 sg13g2_a21oi_1 _24333_ (.A1(net864),
    .A2(_07690_),
    .Y(_07691_),
    .B1(net743));
 sg13g2_a21oi_1 _24334_ (.A1(_08452_),
    .A2(_07435_),
    .Y(_00431_),
    .B1(_07691_));
 sg13g2_a22oi_1 _24335_ (.Y(_07692_),
    .B1(_07599_),
    .B2(\top_ihp.oisc.regs[11][20] ),
    .A2(_07520_),
    .A1(\top_ihp.oisc.regs[9][20] ));
 sg13g2_a22oi_1 _24336_ (.Y(_07693_),
    .B1(_07556_),
    .B2(\top_ihp.oisc.regs[13][20] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[15][20] ));
 sg13g2_nand2_1 _24337_ (.Y(_07694_),
    .A(_07692_),
    .B(_07693_));
 sg13g2_a21oi_1 _24338_ (.A1(\top_ihp.oisc.regs[7][20] ),
    .A2(_07475_),
    .Y(_07695_),
    .B1(_07694_));
 sg13g2_a22oi_1 _24339_ (.Y(_07696_),
    .B1(_07548_),
    .B2(\top_ihp.oisc.regs[12][20] ),
    .A2(_07485_),
    .A1(\top_ihp.oisc.regs[32][20] ));
 sg13g2_a22oi_1 _24340_ (.Y(_07697_),
    .B1(net839),
    .B2(\top_ihp.oisc.regs[10][20] ),
    .A2(net863),
    .A1(\top_ihp.oisc.regs[8][20] ));
 sg13g2_inv_1 _24341_ (.Y(_07698_),
    .A(_00224_));
 sg13g2_a22oi_1 _24342_ (.Y(_07699_),
    .B1(net884),
    .B2(_07698_),
    .A2(_07525_),
    .A1(\top_ihp.oisc.regs[14][20] ));
 sg13g2_nand3_1 _24343_ (.B(_07697_),
    .C(_07699_),
    .A(_07696_),
    .Y(_07700_));
 sg13g2_a221oi_1 _24344_ (.B2(\top_ihp.oisc.regs[2][20] ),
    .C1(_07700_),
    .B1(net815),
    .A1(\top_ihp.oisc.regs[3][20] ),
    .Y(_07701_),
    .A2(_07507_));
 sg13g2_a22oi_1 _24345_ (.Y(_07702_),
    .B1(net772),
    .B2(\top_ihp.oisc.regs[6][20] ),
    .A2(net814),
    .A1(\top_ihp.oisc.regs[1][20] ));
 sg13g2_a22oi_1 _24346_ (.Y(_07703_),
    .B1(net791),
    .B2(\top_ihp.oisc.regs[4][20] ),
    .A2(net795),
    .A1(\top_ihp.oisc.regs[5][20] ));
 sg13g2_nand4_1 _24347_ (.B(_07701_),
    .C(_07702_),
    .A(_07695_),
    .Y(_07704_),
    .D(_07703_));
 sg13g2_a21oi_1 _24348_ (.A1(net864),
    .A2(_07704_),
    .Y(_07705_),
    .B1(_07537_));
 sg13g2_a21oi_1 _24349_ (.A1(_07991_),
    .A2(net745),
    .Y(_00432_),
    .B1(_07705_));
 sg13g2_and2_1 _24350_ (.A(\top_ihp.oisc.regs[2][21] ),
    .B(_07511_),
    .X(_07706_));
 sg13g2_a221oi_1 _24351_ (.B2(\top_ihp.oisc.regs[4][21] ),
    .C1(_07706_),
    .B1(net793),
    .A1(\top_ihp.oisc.regs[6][21] ),
    .Y(_07707_),
    .A2(net772));
 sg13g2_buf_1 _24352_ (.A(_07496_),
    .X(_07708_));
 sg13g2_a21oi_1 _24353_ (.A1(\top_ihp.oisc.regs[9][21] ),
    .A2(_07487_),
    .Y(_07709_),
    .B1(net892));
 sg13g2_a22oi_1 _24354_ (.Y(_07710_),
    .B1(_07454_),
    .B2(\top_ihp.oisc.regs[15][21] ),
    .A2(_07447_),
    .A1(\top_ihp.oisc.regs[8][21] ));
 sg13g2_nand2_1 _24355_ (.Y(_07711_),
    .A(_07709_),
    .B(_07710_));
 sg13g2_a221oi_1 _24356_ (.B2(\top_ihp.oisc.regs[11][21] ),
    .C1(_07711_),
    .B1(_07599_),
    .A1(\top_ihp.oisc.regs[12][21] ),
    .Y(_07712_),
    .A2(_07548_));
 sg13g2_a22oi_1 _24357_ (.Y(_07713_),
    .B1(net813),
    .B2(\top_ihp.oisc.regs[13][21] ),
    .A2(net838),
    .A1(\top_ihp.oisc.regs[32][21] ));
 sg13g2_a22oi_1 _24358_ (.Y(_07714_),
    .B1(net829),
    .B2(\top_ihp.oisc.regs[14][21] ),
    .A2(_07462_),
    .A1(\top_ihp.oisc.regs[10][21] ));
 sg13g2_a22oi_1 _24359_ (.Y(_07715_),
    .B1(net792),
    .B2(\top_ihp.oisc.regs[7][21] ),
    .A2(_07443_),
    .A1(\top_ihp.oisc.regs[5][21] ));
 sg13g2_nand4_1 _24360_ (.B(_07713_),
    .C(_07714_),
    .A(_07712_),
    .Y(_07716_),
    .D(_07715_));
 sg13g2_a221oi_1 _24361_ (.B2(\top_ihp.oisc.regs[3][21] ),
    .C1(_07716_),
    .B1(net819),
    .A1(\top_ihp.oisc.regs[1][21] ),
    .Y(_07717_),
    .A2(net814));
 sg13g2_a221oi_1 _24362_ (.B2(_07717_),
    .C1(net840),
    .B1(_07707_),
    .A1(_00225_),
    .Y(_07718_),
    .A2(net861));
 sg13g2_mux2_1 _24363_ (.A0(_08153_),
    .A1(_07718_),
    .S(net770),
    .X(_00433_));
 sg13g2_a22oi_1 _24364_ (.Y(_07719_),
    .B1(net796),
    .B2(\top_ihp.oisc.regs[4][22] ),
    .A2(net814),
    .A1(\top_ihp.oisc.regs[1][22] ));
 sg13g2_nand2_1 _24365_ (.Y(_07720_),
    .A(\top_ihp.oisc.regs[5][22] ),
    .B(net794));
 sg13g2_buf_1 _24366_ (.A(_07480_),
    .X(_07721_));
 sg13g2_a22oi_1 _24367_ (.Y(_07722_),
    .B1(net844),
    .B2(\top_ihp.oisc.regs[9][22] ),
    .A2(_07721_),
    .A1(\top_ihp.oisc.regs[12][22] ));
 sg13g2_a21o_1 _24368_ (.A2(net817),
    .A1(\top_ihp.oisc.regs[15][22] ),
    .B1(_07708_),
    .X(_07723_));
 sg13g2_a221oi_1 _24369_ (.B2(\top_ihp.oisc.regs[11][22] ),
    .C1(_07723_),
    .B1(net843),
    .A1(\top_ihp.oisc.regs[10][22] ),
    .Y(_07724_),
    .A2(net839));
 sg13g2_a22oi_1 _24370_ (.Y(_07725_),
    .B1(net827),
    .B2(\top_ihp.oisc.regs[13][22] ),
    .A2(net859),
    .A1(\top_ihp.oisc.regs[32][22] ));
 sg13g2_a22oi_1 _24371_ (.Y(_07726_),
    .B1(net822),
    .B2(\top_ihp.oisc.regs[14][22] ),
    .A2(_07448_),
    .A1(\top_ihp.oisc.regs[8][22] ));
 sg13g2_nand4_1 _24372_ (.B(_07724_),
    .C(_07725_),
    .A(_07722_),
    .Y(_07727_),
    .D(_07726_));
 sg13g2_a221oi_1 _24373_ (.B2(\top_ihp.oisc.regs[6][22] ),
    .C1(_07727_),
    .B1(net771),
    .A1(\top_ihp.oisc.regs[7][22] ),
    .Y(_07728_),
    .A2(net798));
 sg13g2_a22oi_1 _24374_ (.Y(_07729_),
    .B1(_07546_),
    .B2(\top_ihp.oisc.regs[3][22] ),
    .A2(net823),
    .A1(\top_ihp.oisc.regs[2][22] ));
 sg13g2_nand4_1 _24375_ (.B(_07720_),
    .C(_07728_),
    .A(_07719_),
    .Y(_07730_),
    .D(_07729_));
 sg13g2_a21oi_1 _24376_ (.A1(_00226_),
    .A2(net885),
    .Y(_07731_),
    .B1(net860));
 sg13g2_a21oi_1 _24377_ (.A1(_07730_),
    .A2(_07731_),
    .Y(_07732_),
    .B1(net743));
 sg13g2_a21oi_1 _24378_ (.A1(_08393_),
    .A2(net745),
    .Y(_00434_),
    .B1(_07732_));
 sg13g2_a22oi_1 _24379_ (.Y(_07733_),
    .B1(net816),
    .B2(\top_ihp.oisc.regs[13][23] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[15][23] ));
 sg13g2_a22oi_1 _24380_ (.Y(_07734_),
    .B1(net829),
    .B2(\top_ihp.oisc.regs[14][23] ),
    .A2(_07449_),
    .A1(\top_ihp.oisc.regs[8][23] ));
 sg13g2_nand2_1 _24381_ (.Y(_07735_),
    .A(_07733_),
    .B(_07734_));
 sg13g2_a21oi_1 _24382_ (.A1(\top_ihp.oisc.regs[5][23] ),
    .A2(net800),
    .Y(_07736_),
    .B1(_07735_));
 sg13g2_a22oi_1 _24383_ (.Y(_07737_),
    .B1(net818),
    .B2(\top_ihp.oisc.regs[12][23] ),
    .A2(net839),
    .A1(\top_ihp.oisc.regs[10][23] ));
 sg13g2_a22oi_1 _24384_ (.Y(_07738_),
    .B1(net844),
    .B2(\top_ihp.oisc.regs[9][23] ),
    .A2(net859),
    .A1(\top_ihp.oisc.regs[32][23] ));
 sg13g2_inv_1 _24385_ (.Y(_07739_),
    .A(_00227_));
 sg13g2_a22oi_1 _24386_ (.Y(_07740_),
    .B1(net884),
    .B2(_07739_),
    .A2(net825),
    .A1(\top_ihp.oisc.regs[11][23] ));
 sg13g2_nand3_1 _24387_ (.B(_07738_),
    .C(_07740_),
    .A(_07737_),
    .Y(_07741_));
 sg13g2_a221oi_1 _24388_ (.B2(\top_ihp.oisc.regs[7][23] ),
    .C1(_07741_),
    .B1(net798),
    .A1(\top_ihp.oisc.regs[1][23] ),
    .Y(_07742_),
    .A2(net828));
 sg13g2_a22oi_1 _24389_ (.Y(_07743_),
    .B1(net824),
    .B2(\top_ihp.oisc.regs[3][23] ),
    .A2(net771),
    .A1(\top_ihp.oisc.regs[6][23] ));
 sg13g2_a22oi_1 _24390_ (.Y(_07744_),
    .B1(net791),
    .B2(\top_ihp.oisc.regs[4][23] ),
    .A2(net815),
    .A1(\top_ihp.oisc.regs[2][23] ));
 sg13g2_nand4_1 _24391_ (.B(_07742_),
    .C(_07743_),
    .A(_07736_),
    .Y(_07745_),
    .D(_07744_));
 sg13g2_a21oi_1 _24392_ (.A1(_07438_),
    .A2(_07745_),
    .Y(_07746_),
    .B1(_07537_));
 sg13g2_a21oi_1 _24393_ (.A1(_10220_),
    .A2(_07435_),
    .Y(_00435_),
    .B1(_07746_));
 sg13g2_and2_1 _24394_ (.A(\top_ihp.oisc.regs[1][24] ),
    .B(_07542_),
    .X(_07747_));
 sg13g2_a221oi_1 _24395_ (.B2(\top_ihp.oisc.regs[4][24] ),
    .C1(_07747_),
    .B1(_07541_),
    .A1(\top_ihp.oisc.regs[5][24] ),
    .Y(_07748_),
    .A2(_07540_));
 sg13g2_a21oi_1 _24396_ (.A1(\top_ihp.oisc.regs[15][24] ),
    .A2(net817),
    .Y(_07749_),
    .B1(net892));
 sg13g2_a22oi_1 _24397_ (.Y(_07750_),
    .B1(net843),
    .B2(\top_ihp.oisc.regs[11][24] ),
    .A2(net845),
    .A1(\top_ihp.oisc.regs[10][24] ));
 sg13g2_nand2_1 _24398_ (.Y(_07751_),
    .A(_07749_),
    .B(_07750_));
 sg13g2_a221oi_1 _24399_ (.B2(\top_ihp.oisc.regs[9][24] ),
    .C1(_07751_),
    .B1(_07549_),
    .A1(\top_ihp.oisc.regs[12][24] ),
    .Y(_07752_),
    .A2(net810));
 sg13g2_a22oi_1 _24400_ (.Y(_07753_),
    .B1(net813),
    .B2(\top_ihp.oisc.regs[13][24] ),
    .A2(net838),
    .A1(\top_ihp.oisc.regs[32][24] ));
 sg13g2_a22oi_1 _24401_ (.Y(_07754_),
    .B1(_07677_),
    .B2(\top_ihp.oisc.regs[14][24] ),
    .A2(net858),
    .A1(\top_ihp.oisc.regs[8][24] ));
 sg13g2_a22oi_1 _24402_ (.Y(_07755_),
    .B1(_07504_),
    .B2(\top_ihp.oisc.regs[6][24] ),
    .A2(net792),
    .A1(\top_ihp.oisc.regs[7][24] ));
 sg13g2_nand4_1 _24403_ (.B(_07753_),
    .C(_07754_),
    .A(_07752_),
    .Y(_07756_),
    .D(_07755_));
 sg13g2_a221oi_1 _24404_ (.B2(\top_ihp.oisc.regs[3][24] ),
    .C1(_07756_),
    .B1(net819),
    .A1(\top_ihp.oisc.regs[2][24] ),
    .Y(_07757_),
    .A2(_07532_));
 sg13g2_a221oi_1 _24405_ (.B2(_07757_),
    .C1(net840),
    .B1(_07748_),
    .A1(_00228_),
    .Y(_07758_),
    .A2(net861));
 sg13g2_mux2_1 _24406_ (.A0(_08155_),
    .A1(_07758_),
    .S(net770),
    .X(_00436_));
 sg13g2_a22oi_1 _24407_ (.Y(_07759_),
    .B1(net830),
    .B2(\top_ihp.oisc.regs[10][25] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[15][25] ));
 sg13g2_a22oi_1 _24408_ (.Y(_07760_),
    .B1(net816),
    .B2(\top_ihp.oisc.regs[13][25] ),
    .A2(net822),
    .A1(\top_ihp.oisc.regs[14][25] ));
 sg13g2_nand2_1 _24409_ (.Y(_07761_),
    .A(_07759_),
    .B(_07760_));
 sg13g2_a21oi_1 _24410_ (.A1(\top_ihp.oisc.regs[5][25] ),
    .A2(net800),
    .Y(_07762_),
    .B1(_07761_));
 sg13g2_a22oi_1 _24411_ (.Y(_07763_),
    .B1(net818),
    .B2(\top_ihp.oisc.regs[12][25] ),
    .A2(net863),
    .A1(\top_ihp.oisc.regs[8][25] ));
 sg13g2_a22oi_1 _24412_ (.Y(_07764_),
    .B1(net844),
    .B2(\top_ihp.oisc.regs[9][25] ),
    .A2(net859),
    .A1(\top_ihp.oisc.regs[32][25] ));
 sg13g2_inv_1 _24413_ (.Y(_07765_),
    .A(_00229_));
 sg13g2_a22oi_1 _24414_ (.Y(_07766_),
    .B1(net884),
    .B2(_07765_),
    .A2(net825),
    .A1(\top_ihp.oisc.regs[11][25] ));
 sg13g2_nand3_1 _24415_ (.B(_07764_),
    .C(_07766_),
    .A(_07763_),
    .Y(_07767_));
 sg13g2_a221oi_1 _24416_ (.B2(\top_ihp.oisc.regs[7][25] ),
    .C1(_07767_),
    .B1(net798),
    .A1(\top_ihp.oisc.regs[1][25] ),
    .Y(_07768_),
    .A2(net828));
 sg13g2_a22oi_1 _24417_ (.Y(_07769_),
    .B1(net824),
    .B2(\top_ihp.oisc.regs[3][25] ),
    .A2(net771),
    .A1(\top_ihp.oisc.regs[6][25] ));
 sg13g2_a22oi_1 _24418_ (.Y(_07770_),
    .B1(net791),
    .B2(\top_ihp.oisc.regs[4][25] ),
    .A2(net815),
    .A1(\top_ihp.oisc.regs[2][25] ));
 sg13g2_nand4_1 _24419_ (.B(_07768_),
    .C(_07769_),
    .A(_07762_),
    .Y(_07771_),
    .D(_07770_));
 sg13g2_a21oi_1 _24420_ (.A1(_07438_),
    .A2(_07771_),
    .Y(_07772_),
    .B1(net743));
 sg13g2_a21oi_1 _24421_ (.A1(_08437_),
    .A2(net744),
    .Y(_00437_),
    .B1(_07772_));
 sg13g2_a22oi_1 _24422_ (.Y(_07773_),
    .B1(net796),
    .B2(\top_ihp.oisc.regs[4][26] ),
    .A2(net814),
    .A1(\top_ihp.oisc.regs[1][26] ));
 sg13g2_nand2_1 _24423_ (.Y(_07774_),
    .A(\top_ihp.oisc.regs[5][26] ),
    .B(net794));
 sg13g2_a22oi_1 _24424_ (.Y(_07775_),
    .B1(net844),
    .B2(\top_ihp.oisc.regs[9][26] ),
    .A2(net831),
    .A1(\top_ihp.oisc.regs[15][26] ));
 sg13g2_a21o_1 _24425_ (.A2(_07464_),
    .A1(\top_ihp.oisc.regs[14][26] ),
    .B1(_07708_),
    .X(_07776_));
 sg13g2_a221oi_1 _24426_ (.B2(\top_ihp.oisc.regs[12][26] ),
    .C1(_07776_),
    .B1(net810),
    .A1(\top_ihp.oisc.regs[10][26] ),
    .Y(_07777_),
    .A2(net845));
 sg13g2_a22oi_1 _24427_ (.Y(_07778_),
    .B1(net827),
    .B2(\top_ihp.oisc.regs[13][26] ),
    .A2(net859),
    .A1(\top_ihp.oisc.regs[32][26] ));
 sg13g2_a22oi_1 _24428_ (.Y(_07779_),
    .B1(_07493_),
    .B2(\top_ihp.oisc.regs[11][26] ),
    .A2(net863),
    .A1(\top_ihp.oisc.regs[8][26] ));
 sg13g2_nand4_1 _24429_ (.B(_07777_),
    .C(_07778_),
    .A(_07775_),
    .Y(_07780_),
    .D(_07779_));
 sg13g2_a221oi_1 _24430_ (.B2(\top_ihp.oisc.regs[6][26] ),
    .C1(_07780_),
    .B1(_07531_),
    .A1(\top_ihp.oisc.regs[7][26] ),
    .Y(_07781_),
    .A2(net798));
 sg13g2_a22oi_1 _24431_ (.Y(_07782_),
    .B1(_07546_),
    .B2(\top_ihp.oisc.regs[3][26] ),
    .A2(net823),
    .A1(\top_ihp.oisc.regs[2][26] ));
 sg13g2_nand4_1 _24432_ (.B(_07774_),
    .C(_07781_),
    .A(_07773_),
    .Y(_07783_),
    .D(_07782_));
 sg13g2_a21oi_1 _24433_ (.A1(_00230_),
    .A2(net885),
    .Y(_07784_),
    .B1(net860));
 sg13g2_a21oi_1 _24434_ (.A1(_07783_),
    .A2(_07784_),
    .Y(_07785_),
    .B1(_04088_));
 sg13g2_a21oi_1 _24435_ (.A1(_07989_),
    .A2(net744),
    .Y(_00438_),
    .B1(_07785_));
 sg13g2_and2_1 _24436_ (.A(\top_ihp.oisc.regs[1][27] ),
    .B(net820),
    .X(_07786_));
 sg13g2_a221oi_1 _24437_ (.B2(\top_ihp.oisc.regs[4][27] ),
    .C1(_07786_),
    .B1(net793),
    .A1(\top_ihp.oisc.regs[5][27] ),
    .Y(_07787_),
    .A2(_07540_));
 sg13g2_a21oi_1 _24438_ (.A1(\top_ihp.oisc.regs[15][27] ),
    .A2(net817),
    .Y(_07788_),
    .B1(net892));
 sg13g2_a22oi_1 _24439_ (.Y(_07789_),
    .B1(net843),
    .B2(\top_ihp.oisc.regs[11][27] ),
    .A2(_07447_),
    .A1(\top_ihp.oisc.regs[8][27] ));
 sg13g2_nand2_1 _24440_ (.Y(_07790_),
    .A(_07788_),
    .B(_07789_));
 sg13g2_a221oi_1 _24441_ (.B2(\top_ihp.oisc.regs[13][27] ),
    .C1(_07790_),
    .B1(_07478_),
    .A1(\top_ihp.oisc.regs[14][27] ),
    .Y(_07791_),
    .A2(_07525_));
 sg13g2_a22oi_1 _24442_ (.Y(_07792_),
    .B1(_07481_),
    .B2(\top_ihp.oisc.regs[12][27] ),
    .A2(net838),
    .A1(\top_ihp.oisc.regs[32][27] ));
 sg13g2_a22oi_1 _24443_ (.Y(_07793_),
    .B1(net842),
    .B2(\top_ihp.oisc.regs[9][27] ),
    .A2(_07602_),
    .A1(\top_ihp.oisc.regs[10][27] ));
 sg13g2_a22oi_1 _24444_ (.Y(_07794_),
    .B1(net797),
    .B2(\top_ihp.oisc.regs[6][27] ),
    .A2(net792),
    .A1(\top_ihp.oisc.regs[7][27] ));
 sg13g2_nand4_1 _24445_ (.B(_07792_),
    .C(_07793_),
    .A(_07791_),
    .Y(_07795_),
    .D(_07794_));
 sg13g2_a221oi_1 _24446_ (.B2(\top_ihp.oisc.regs[3][27] ),
    .C1(_07795_),
    .B1(net819),
    .A1(\top_ihp.oisc.regs[2][27] ),
    .Y(_07796_),
    .A2(net821));
 sg13g2_a221oi_1 _24447_ (.B2(_07796_),
    .C1(net840),
    .B1(_07787_),
    .A1(_00231_),
    .Y(_07797_),
    .A2(net861));
 sg13g2_mux2_1 _24448_ (.A0(_08284_),
    .A1(_07797_),
    .S(net770),
    .X(_00439_));
 sg13g2_and2_1 _24449_ (.A(\top_ihp.oisc.regs[1][28] ),
    .B(net820),
    .X(_07798_));
 sg13g2_a221oi_1 _24450_ (.B2(\top_ihp.oisc.regs[4][28] ),
    .C1(_07798_),
    .B1(_07541_),
    .A1(\top_ihp.oisc.regs[5][28] ),
    .Y(_07799_),
    .A2(_07444_));
 sg13g2_a21oi_1 _24451_ (.A1(\top_ihp.oisc.regs[15][28] ),
    .A2(net817),
    .Y(_07800_),
    .B1(net892));
 sg13g2_a22oi_1 _24452_ (.Y(_07801_),
    .B1(net843),
    .B2(\top_ihp.oisc.regs[11][28] ),
    .A2(net845),
    .A1(\top_ihp.oisc.regs[10][28] ));
 sg13g2_nand2_1 _24453_ (.Y(_07802_),
    .A(_07800_),
    .B(_07801_));
 sg13g2_a221oi_1 _24454_ (.B2(\top_ihp.oisc.regs[9][28] ),
    .C1(_07802_),
    .B1(net841),
    .A1(\top_ihp.oisc.regs[12][28] ),
    .Y(_07803_),
    .A2(_07721_));
 sg13g2_a22oi_1 _24455_ (.Y(_07804_),
    .B1(net813),
    .B2(\top_ihp.oisc.regs[13][28] ),
    .A2(net838),
    .A1(\top_ihp.oisc.regs[32][28] ));
 sg13g2_a22oi_1 _24456_ (.Y(_07805_),
    .B1(net811),
    .B2(\top_ihp.oisc.regs[14][28] ),
    .A2(net858),
    .A1(\top_ihp.oisc.regs[8][28] ));
 sg13g2_a22oi_1 _24457_ (.Y(_07806_),
    .B1(_07503_),
    .B2(\top_ihp.oisc.regs[6][28] ),
    .A2(_07559_),
    .A1(\top_ihp.oisc.regs[7][28] ));
 sg13g2_nand4_1 _24458_ (.B(_07804_),
    .C(_07805_),
    .A(_07803_),
    .Y(_07807_),
    .D(_07806_));
 sg13g2_a221oi_1 _24459_ (.B2(\top_ihp.oisc.regs[3][28] ),
    .C1(_07807_),
    .B1(_07547_),
    .A1(\top_ihp.oisc.regs[2][28] ),
    .Y(_07808_),
    .A2(_07532_));
 sg13g2_a221oi_1 _24460_ (.B2(_07808_),
    .C1(_07563_),
    .B1(_07799_),
    .A1(_00069_),
    .Y(_07809_),
    .A2(_07539_));
 sg13g2_mux2_1 _24461_ (.A0(_08277_),
    .A1(_07809_),
    .S(_07565_),
    .X(_00440_));
 sg13g2_a22oi_1 _24462_ (.Y(_07810_),
    .B1(net842),
    .B2(\top_ihp.oisc.regs[9][29] ),
    .A2(net811),
    .A1(\top_ihp.oisc.regs[14][29] ));
 sg13g2_a22oi_1 _24463_ (.Y(_07811_),
    .B1(net826),
    .B2(\top_ihp.oisc.regs[12][29] ),
    .A2(net830),
    .A1(\top_ihp.oisc.regs[10][29] ));
 sg13g2_nand2_1 _24464_ (.Y(_07812_),
    .A(_07810_),
    .B(_07811_));
 sg13g2_a21oi_1 _24465_ (.A1(\top_ihp.oisc.regs[2][29] ),
    .A2(net823),
    .Y(_07813_),
    .B1(_07812_));
 sg13g2_a22oi_1 _24466_ (.Y(_07814_),
    .B1(net858),
    .B2(\top_ihp.oisc.regs[8][29] ),
    .A2(net862),
    .A1(\top_ihp.oisc.regs[32][29] ));
 sg13g2_a22oi_1 _24467_ (.Y(_07815_),
    .B1(net827),
    .B2(\top_ihp.oisc.regs[13][29] ),
    .A2(net831),
    .A1(\top_ihp.oisc.regs[15][29] ));
 sg13g2_inv_1 _24468_ (.Y(_07816_),
    .A(_00070_));
 sg13g2_a22oi_1 _24469_ (.Y(_07817_),
    .B1(_07603_),
    .B2(_07816_),
    .A2(net825),
    .A1(\top_ihp.oisc.regs[11][29] ));
 sg13g2_nand3_1 _24470_ (.B(_07815_),
    .C(_07817_),
    .A(_07814_),
    .Y(_07818_));
 sg13g2_a221oi_1 _24471_ (.B2(\top_ihp.oisc.regs[4][29] ),
    .C1(_07818_),
    .B1(_07514_),
    .A1(\top_ihp.oisc.regs[7][29] ),
    .Y(_07819_),
    .A2(net798));
 sg13g2_a22oi_1 _24472_ (.Y(_07820_),
    .B1(net824),
    .B2(\top_ihp.oisc.regs[3][29] ),
    .A2(net814),
    .A1(\top_ihp.oisc.regs[1][29] ));
 sg13g2_a22oi_1 _24473_ (.Y(_07821_),
    .B1(net772),
    .B2(\top_ihp.oisc.regs[6][29] ),
    .A2(net795),
    .A1(\top_ihp.oisc.regs[5][29] ));
 sg13g2_nand4_1 _24474_ (.B(_07819_),
    .C(_07820_),
    .A(_07813_),
    .Y(_07822_),
    .D(_07821_));
 sg13g2_a21oi_1 _24475_ (.A1(_07437_),
    .A2(_07822_),
    .Y(_07823_),
    .B1(net760));
 sg13g2_a21oi_1 _24476_ (.A1(_08344_),
    .A2(net744),
    .Y(_00441_),
    .B1(_07823_));
 sg13g2_and2_1 _24477_ (.A(\top_ihp.oisc.regs[1][2] ),
    .B(_07542_),
    .X(_07824_));
 sg13g2_a221oi_1 _24478_ (.B2(\top_ihp.oisc.regs[4][2] ),
    .C1(_07824_),
    .B1(net793),
    .A1(\top_ihp.oisc.regs[5][2] ),
    .Y(_07825_),
    .A2(net800));
 sg13g2_a21oi_1 _24479_ (.A1(\top_ihp.oisc.regs[15][2] ),
    .A2(net817),
    .Y(_07826_),
    .B1(net892));
 sg13g2_a22oi_1 _24480_ (.Y(_07827_),
    .B1(_07491_),
    .B2(\top_ihp.oisc.regs[11][2] ),
    .A2(_07461_),
    .A1(\top_ihp.oisc.regs[10][2] ));
 sg13g2_nand2_1 _24481_ (.Y(_07828_),
    .A(_07826_),
    .B(_07827_));
 sg13g2_a221oi_1 _24482_ (.B2(\top_ihp.oisc.regs[9][2] ),
    .C1(_07828_),
    .B1(net841),
    .A1(\top_ihp.oisc.regs[12][2] ),
    .Y(_07829_),
    .A2(net810));
 sg13g2_a22oi_1 _24483_ (.Y(_07830_),
    .B1(net813),
    .B2(\top_ihp.oisc.regs[13][2] ),
    .A2(net838),
    .A1(\top_ihp.oisc.regs[32][2] ));
 sg13g2_a22oi_1 _24484_ (.Y(_07831_),
    .B1(net811),
    .B2(\top_ihp.oisc.regs[14][2] ),
    .A2(_07682_),
    .A1(\top_ihp.oisc.regs[8][2] ));
 sg13g2_a22oi_1 _24485_ (.Y(_07832_),
    .B1(_07503_),
    .B2(\top_ihp.oisc.regs[6][2] ),
    .A2(_07559_),
    .A1(\top_ihp.oisc.regs[7][2] ));
 sg13g2_nand4_1 _24486_ (.B(_07830_),
    .C(_07831_),
    .A(_07829_),
    .Y(_07833_),
    .D(_07832_));
 sg13g2_a221oi_1 _24487_ (.B2(\top_ihp.oisc.regs[3][2] ),
    .C1(_07833_),
    .B1(_07547_),
    .A1(\top_ihp.oisc.regs[2][2] ),
    .Y(_07834_),
    .A2(_07512_));
 sg13g2_a221oi_1 _24488_ (.B2(_07834_),
    .C1(_07563_),
    .B1(_07825_),
    .A1(_00206_),
    .Y(_07835_),
    .A2(_07539_));
 sg13g2_mux2_1 _24489_ (.A0(_08091_),
    .A1(_07835_),
    .S(_07565_),
    .X(_00442_));
 sg13g2_a22oi_1 _24490_ (.Y(_07836_),
    .B1(net812),
    .B2(\top_ihp.oisc.regs[11][30] ),
    .A2(net811),
    .A1(\top_ihp.oisc.regs[14][30] ));
 sg13g2_a22oi_1 _24491_ (.Y(_07837_),
    .B1(_07520_),
    .B2(\top_ihp.oisc.regs[9][30] ),
    .A2(net827),
    .A1(\top_ihp.oisc.regs[13][30] ));
 sg13g2_nand2_1 _24492_ (.Y(_07838_),
    .A(_07836_),
    .B(_07837_));
 sg13g2_a21oi_1 _24493_ (.A1(\top_ihp.oisc.regs[7][30] ),
    .A2(_07475_),
    .Y(_07839_),
    .B1(_07838_));
 sg13g2_a22oi_1 _24494_ (.Y(_07840_),
    .B1(net858),
    .B2(\top_ihp.oisc.regs[8][30] ),
    .A2(_07485_),
    .A1(\top_ihp.oisc.regs[32][30] ));
 sg13g2_a22oi_1 _24495_ (.Y(_07841_),
    .B1(net818),
    .B2(\top_ihp.oisc.regs[12][30] ),
    .A2(net831),
    .A1(\top_ihp.oisc.regs[15][30] ));
 sg13g2_a22oi_1 _24496_ (.Y(_07842_),
    .B1(_07603_),
    .B2(_07002_),
    .A2(_07602_),
    .A1(\top_ihp.oisc.regs[10][30] ));
 sg13g2_nand3_1 _24497_ (.B(_07841_),
    .C(_07842_),
    .A(_07840_),
    .Y(_07843_));
 sg13g2_a221oi_1 _24498_ (.B2(\top_ihp.oisc.regs[2][30] ),
    .C1(_07843_),
    .B1(net815),
    .A1(\top_ihp.oisc.regs[3][30] ),
    .Y(_07844_),
    .A2(_07507_));
 sg13g2_a22oi_1 _24499_ (.Y(_07845_),
    .B1(net772),
    .B2(\top_ihp.oisc.regs[6][30] ),
    .A2(net814),
    .A1(\top_ihp.oisc.regs[1][30] ));
 sg13g2_a22oi_1 _24500_ (.Y(_07846_),
    .B1(_07634_),
    .B2(\top_ihp.oisc.regs[4][30] ),
    .A2(net795),
    .A1(\top_ihp.oisc.regs[5][30] ));
 sg13g2_nand4_1 _24501_ (.B(_07844_),
    .C(_07845_),
    .A(_07839_),
    .Y(_07847_),
    .D(_07846_));
 sg13g2_a21oi_1 _24502_ (.A1(_07437_),
    .A2(_07847_),
    .Y(_07848_),
    .B1(net760));
 sg13g2_a21oi_1 _24503_ (.A1(_08315_),
    .A2(net744),
    .Y(_00443_),
    .B1(_07848_));
 sg13g2_and2_1 _24504_ (.A(\top_ihp.oisc.regs[2][31] ),
    .B(_07511_),
    .X(_07849_));
 sg13g2_a221oi_1 _24505_ (.B2(\top_ihp.oisc.regs[6][31] ),
    .C1(_07849_),
    .B1(_07505_),
    .A1(\top_ihp.oisc.regs[5][31] ),
    .Y(_07850_),
    .A2(net800));
 sg13g2_a21oi_1 _24506_ (.A1(\top_ihp.oisc.regs[15][31] ),
    .A2(_07550_),
    .Y(_07851_),
    .B1(net892));
 sg13g2_a22oi_1 _24507_ (.Y(_07852_),
    .B1(_07491_),
    .B2(\top_ihp.oisc.regs[11][31] ),
    .A2(_07460_),
    .A1(\top_ihp.oisc.regs[10][31] ));
 sg13g2_nand2_1 _24508_ (.Y(_07853_),
    .A(_07851_),
    .B(_07852_));
 sg13g2_a221oi_1 _24509_ (.B2(\top_ihp.oisc.regs[9][31] ),
    .C1(_07853_),
    .B1(net841),
    .A1(\top_ihp.oisc.regs[12][31] ),
    .Y(_07854_),
    .A2(net810));
 sg13g2_a22oi_1 _24510_ (.Y(_07855_),
    .B1(_07595_),
    .B2(\top_ihp.oisc.regs[13][31] ),
    .A2(_07644_),
    .A1(\top_ihp.oisc.regs[32][31] ));
 sg13g2_a22oi_1 _24511_ (.Y(_07856_),
    .B1(net811),
    .B2(\top_ihp.oisc.regs[14][31] ),
    .A2(net858),
    .A1(\top_ihp.oisc.regs[8][31] ));
 sg13g2_a22oi_1 _24512_ (.Y(_07857_),
    .B1(_07546_),
    .B2(\top_ihp.oisc.regs[3][31] ),
    .A2(_07473_),
    .A1(\top_ihp.oisc.regs[7][31] ));
 sg13g2_nand4_1 _24513_ (.B(_07855_),
    .C(_07856_),
    .A(_07854_),
    .Y(_07858_),
    .D(_07857_));
 sg13g2_a221oi_1 _24514_ (.B2(\top_ihp.oisc.regs[4][31] ),
    .C1(_07858_),
    .B1(net796),
    .A1(\top_ihp.oisc.regs[1][31] ),
    .Y(_07859_),
    .A2(_07577_));
 sg13g2_a221oi_1 _24515_ (.B2(_07859_),
    .C1(net860),
    .B1(_07850_),
    .A1(_00072_),
    .Y(_07860_),
    .A2(_07498_));
 sg13g2_mux2_1 _24516_ (.A0(_09498_),
    .A1(_07860_),
    .S(net804),
    .X(_00444_));
 sg13g2_a22oi_1 _24517_ (.Y(_07861_),
    .B1(net816),
    .B2(\top_ihp.oisc.regs[13][3] ),
    .A2(net846),
    .A1(\top_ihp.oisc.regs[8][3] ));
 sg13g2_a22oi_1 _24518_ (.Y(_07862_),
    .B1(_07465_),
    .B2(\top_ihp.oisc.regs[14][3] ),
    .A2(_07462_),
    .A1(\top_ihp.oisc.regs[10][3] ));
 sg13g2_nand2_1 _24519_ (.Y(_07863_),
    .A(_07861_),
    .B(_07862_));
 sg13g2_a21oi_1 _24520_ (.A1(\top_ihp.oisc.regs[5][3] ),
    .A2(net795),
    .Y(_07864_),
    .B1(_07863_));
 sg13g2_a22oi_1 _24521_ (.Y(_07865_),
    .B1(_07493_),
    .B2(\top_ihp.oisc.regs[11][3] ),
    .A2(net810),
    .A1(\top_ihp.oisc.regs[12][3] ));
 sg13g2_a22oi_1 _24522_ (.Y(_07866_),
    .B1(net844),
    .B2(\top_ihp.oisc.regs[9][3] ),
    .A2(net859),
    .A1(\top_ihp.oisc.regs[32][3] ));
 sg13g2_inv_1 _24523_ (.Y(_07867_),
    .A(_00207_));
 sg13g2_a22oi_1 _24524_ (.Y(_07868_),
    .B1(net884),
    .B2(_07867_),
    .A2(net831),
    .A1(\top_ihp.oisc.regs[15][3] ));
 sg13g2_nand3_1 _24525_ (.B(_07866_),
    .C(_07868_),
    .A(_07865_),
    .Y(_07869_));
 sg13g2_a221oi_1 _24526_ (.B2(\top_ihp.oisc.regs[7][3] ),
    .C1(_07869_),
    .B1(_07474_),
    .A1(\top_ihp.oisc.regs[1][3] ),
    .Y(_07870_),
    .A2(_07471_));
 sg13g2_a22oi_1 _24527_ (.Y(_07871_),
    .B1(net824),
    .B2(\top_ihp.oisc.regs[3][3] ),
    .A2(net771),
    .A1(\top_ihp.oisc.regs[6][3] ));
 sg13g2_a22oi_1 _24528_ (.Y(_07872_),
    .B1(net791),
    .B2(\top_ihp.oisc.regs[4][3] ),
    .A2(_07570_),
    .A1(\top_ihp.oisc.regs[2][3] ));
 sg13g2_nand4_1 _24529_ (.B(_07870_),
    .C(_07871_),
    .A(_07864_),
    .Y(_07873_),
    .D(_07872_));
 sg13g2_a21oi_1 _24530_ (.A1(_07437_),
    .A2(_07873_),
    .Y(_07874_),
    .B1(net760));
 sg13g2_a21oi_1 _24531_ (.A1(_04178_),
    .A2(net744),
    .Y(_00445_),
    .B1(_07874_));
 sg13g2_and2_1 _24532_ (.A(\top_ihp.oisc.regs[1][4] ),
    .B(_07470_),
    .X(_07875_));
 sg13g2_a221oi_1 _24533_ (.B2(\top_ihp.oisc.regs[4][4] ),
    .C1(_07875_),
    .B1(net796),
    .A1(\top_ihp.oisc.regs[5][4] ),
    .Y(_07876_),
    .A2(net800));
 sg13g2_a21oi_1 _24534_ (.A1(\top_ihp.oisc.regs[15][4] ),
    .A2(_07550_),
    .Y(_07877_),
    .B1(net892));
 sg13g2_a22oi_1 _24535_ (.Y(_07878_),
    .B1(_07491_),
    .B2(\top_ihp.oisc.regs[11][4] ),
    .A2(_07460_),
    .A1(\top_ihp.oisc.regs[10][4] ));
 sg13g2_nand2_1 _24536_ (.Y(_07879_),
    .A(_07877_),
    .B(_07878_));
 sg13g2_a221oi_1 _24537_ (.B2(\top_ihp.oisc.regs[9][4] ),
    .C1(_07879_),
    .B1(_07549_),
    .A1(\top_ihp.oisc.regs[12][4] ),
    .Y(_07880_),
    .A2(net810));
 sg13g2_a22oi_1 _24538_ (.Y(_07881_),
    .B1(_07595_),
    .B2(\top_ihp.oisc.regs[13][4] ),
    .A2(net838),
    .A1(\top_ihp.oisc.regs[32][4] ));
 sg13g2_a22oi_1 _24539_ (.Y(_07882_),
    .B1(net811),
    .B2(\top_ihp.oisc.regs[14][4] ),
    .A2(net858),
    .A1(\top_ihp.oisc.regs[8][4] ));
 sg13g2_a22oi_1 _24540_ (.Y(_07883_),
    .B1(_07503_),
    .B2(\top_ihp.oisc.regs[6][4] ),
    .A2(_07473_),
    .A1(\top_ihp.oisc.regs[7][4] ));
 sg13g2_nand4_1 _24541_ (.B(_07881_),
    .C(_07882_),
    .A(_07880_),
    .Y(_07884_),
    .D(_07883_));
 sg13g2_a221oi_1 _24542_ (.B2(\top_ihp.oisc.regs[3][4] ),
    .C1(_07884_),
    .B1(_07546_),
    .A1(\top_ihp.oisc.regs[2][4] ),
    .Y(_07885_),
    .A2(net823));
 sg13g2_a221oi_1 _24543_ (.B2(_07885_),
    .C1(_07555_),
    .B1(_07876_),
    .A1(_00208_),
    .Y(_07886_),
    .A2(_07498_));
 sg13g2_mux2_1 _24544_ (.A0(_08110_),
    .A1(_07886_),
    .S(net804),
    .X(_00446_));
 sg13g2_inv_1 _24545_ (.Y(_07887_),
    .A(_08127_));
 sg13g2_a22oi_1 _24546_ (.Y(_07888_),
    .B1(_07465_),
    .B2(\top_ihp.oisc.regs[14][5] ),
    .A2(_07449_),
    .A1(\top_ihp.oisc.regs[8][5] ));
 sg13g2_a22oi_1 _24547_ (.Y(_07889_),
    .B1(net812),
    .B2(\top_ihp.oisc.regs[11][5] ),
    .A2(net841),
    .A1(\top_ihp.oisc.regs[9][5] ));
 sg13g2_nand2_1 _24548_ (.Y(_07890_),
    .A(_07888_),
    .B(_07889_));
 sg13g2_a21oi_1 _24549_ (.A1(\top_ihp.oisc.regs[5][5] ),
    .A2(_07534_),
    .Y(_07891_),
    .B1(_07890_));
 sg13g2_a22oi_1 _24550_ (.Y(_07892_),
    .B1(net818),
    .B2(\top_ihp.oisc.regs[12][5] ),
    .A2(_07478_),
    .A1(\top_ihp.oisc.regs[13][5] ));
 sg13g2_a22oi_1 _24551_ (.Y(_07893_),
    .B1(net831),
    .B2(\top_ihp.oisc.regs[15][5] ),
    .A2(_07628_),
    .A1(\top_ihp.oisc.regs[32][5] ));
 sg13g2_inv_1 _24552_ (.Y(_07894_),
    .A(_00209_));
 sg13g2_a22oi_1 _24553_ (.Y(_07895_),
    .B1(net893),
    .B2(_07894_),
    .A2(net839),
    .A1(\top_ihp.oisc.regs[10][5] ));
 sg13g2_nand3_1 _24554_ (.B(_07893_),
    .C(_07895_),
    .A(_07892_),
    .Y(_07896_));
 sg13g2_a221oi_1 _24555_ (.B2(\top_ihp.oisc.regs[7][5] ),
    .C1(_07896_),
    .B1(_07474_),
    .A1(\top_ihp.oisc.regs[1][5] ),
    .Y(_07897_),
    .A2(net820));
 sg13g2_a22oi_1 _24556_ (.Y(_07898_),
    .B1(_07508_),
    .B2(\top_ihp.oisc.regs[3][5] ),
    .A2(_07531_),
    .A1(\top_ihp.oisc.regs[6][5] ));
 sg13g2_a22oi_1 _24557_ (.Y(_07899_),
    .B1(_07634_),
    .B2(\top_ihp.oisc.regs[4][5] ),
    .A2(_07570_),
    .A1(\top_ihp.oisc.regs[2][5] ));
 sg13g2_nand4_1 _24558_ (.B(_07897_),
    .C(_07898_),
    .A(_07891_),
    .Y(_07900_),
    .D(_07899_));
 sg13g2_a21oi_1 _24559_ (.A1(_07437_),
    .A2(_07900_),
    .Y(_07901_),
    .B1(net760));
 sg13g2_a21oi_1 _24560_ (.A1(_07887_),
    .A2(_07518_),
    .Y(_00447_),
    .B1(_07901_));
 sg13g2_a22oi_1 _24561_ (.Y(_07902_),
    .B1(_07515_),
    .B2(\top_ihp.oisc.regs[4][6] ),
    .A2(_07577_),
    .A1(\top_ihp.oisc.regs[1][6] ));
 sg13g2_nand2_1 _24562_ (.Y(_07903_),
    .A(\top_ihp.oisc.regs[5][6] ),
    .B(net794));
 sg13g2_a22oi_1 _24563_ (.Y(_07904_),
    .B1(_07488_),
    .B2(\top_ihp.oisc.regs[9][6] ),
    .A2(net810),
    .A1(\top_ihp.oisc.regs[12][6] ));
 sg13g2_a21o_1 _24564_ (.A2(_07453_),
    .A1(\top_ihp.oisc.regs[15][6] ),
    .B1(_07496_),
    .X(_07905_));
 sg13g2_a221oi_1 _24565_ (.B2(\top_ihp.oisc.regs[11][6] ),
    .C1(_07905_),
    .B1(_07492_),
    .A1(\top_ihp.oisc.regs[10][6] ),
    .Y(_07906_),
    .A2(_07461_));
 sg13g2_a22oi_1 _24566_ (.Y(_07907_),
    .B1(net827),
    .B2(\top_ihp.oisc.regs[13][6] ),
    .A2(_07628_),
    .A1(\top_ihp.oisc.regs[32][6] ));
 sg13g2_a22oi_1 _24567_ (.Y(_07908_),
    .B1(net822),
    .B2(\top_ihp.oisc.regs[14][6] ),
    .A2(net863),
    .A1(\top_ihp.oisc.regs[8][6] ));
 sg13g2_nand4_1 _24568_ (.B(_07906_),
    .C(_07907_),
    .A(_07904_),
    .Y(_07909_),
    .D(_07908_));
 sg13g2_a221oi_1 _24569_ (.B2(\top_ihp.oisc.regs[6][6] ),
    .C1(_07909_),
    .B1(net797),
    .A1(\top_ihp.oisc.regs[7][6] ),
    .Y(_07910_),
    .A2(net798));
 sg13g2_a22oi_1 _24570_ (.Y(_07911_),
    .B1(_07546_),
    .B2(\top_ihp.oisc.regs[3][6] ),
    .A2(_07512_),
    .A1(\top_ihp.oisc.regs[2][6] ));
 sg13g2_nand4_1 _24571_ (.B(_07903_),
    .C(_07910_),
    .A(_07902_),
    .Y(_07912_),
    .D(_07911_));
 sg13g2_a21oi_1 _24572_ (.A1(_00210_),
    .A2(net885),
    .Y(_07913_),
    .B1(net860));
 sg13g2_a21oi_1 _24573_ (.A1(_07912_),
    .A2(_07913_),
    .Y(_07914_),
    .B1(_04088_));
 sg13g2_a21oi_1 _24574_ (.A1(_08399_),
    .A2(net744),
    .Y(_00448_),
    .B1(_07914_));
 sg13g2_a22oi_1 _24575_ (.Y(_07915_),
    .B1(net842),
    .B2(\top_ihp.oisc.regs[9][7] ),
    .A2(net811),
    .A1(\top_ihp.oisc.regs[14][7] ));
 sg13g2_a22oi_1 _24576_ (.Y(_07916_),
    .B1(net826),
    .B2(\top_ihp.oisc.regs[12][7] ),
    .A2(net830),
    .A1(\top_ihp.oisc.regs[10][7] ));
 sg13g2_nand2_1 _24577_ (.Y(_07917_),
    .A(_07915_),
    .B(_07916_));
 sg13g2_a21oi_1 _24578_ (.A1(\top_ihp.oisc.regs[2][7] ),
    .A2(net823),
    .Y(_07918_),
    .B1(_07917_));
 sg13g2_a22oi_1 _24579_ (.Y(_07919_),
    .B1(net858),
    .B2(\top_ihp.oisc.regs[8][7] ),
    .A2(net862),
    .A1(\top_ihp.oisc.regs[32][7] ));
 sg13g2_a22oi_1 _24580_ (.Y(_07920_),
    .B1(net827),
    .B2(\top_ihp.oisc.regs[13][7] ),
    .A2(_07454_),
    .A1(\top_ihp.oisc.regs[15][7] ));
 sg13g2_a22oi_1 _24581_ (.Y(_07921_),
    .B1(net893),
    .B2(_07335_),
    .A2(_07492_),
    .A1(\top_ihp.oisc.regs[11][7] ));
 sg13g2_nand3_1 _24582_ (.B(_07920_),
    .C(_07921_),
    .A(_07919_),
    .Y(_07922_));
 sg13g2_a221oi_1 _24583_ (.B2(\top_ihp.oisc.regs[4][7] ),
    .C1(_07922_),
    .B1(_07514_),
    .A1(\top_ihp.oisc.regs[7][7] ),
    .Y(_07923_),
    .A2(net798));
 sg13g2_a22oi_1 _24584_ (.Y(_07924_),
    .B1(_07508_),
    .B2(\top_ihp.oisc.regs[3][7] ),
    .A2(_07471_),
    .A1(\top_ihp.oisc.regs[1][7] ));
 sg13g2_a22oi_1 _24585_ (.Y(_07925_),
    .B1(_07505_),
    .B2(\top_ihp.oisc.regs[6][7] ),
    .A2(_07534_),
    .A1(\top_ihp.oisc.regs[5][7] ));
 sg13g2_nand4_1 _24586_ (.B(_07923_),
    .C(_07924_),
    .A(_07918_),
    .Y(_07926_),
    .D(_07925_));
 sg13g2_a21oi_1 _24587_ (.A1(_07437_),
    .A2(_07926_),
    .Y(_07927_),
    .B1(net760));
 sg13g2_a21oi_1 _24588_ (.A1(_08406_),
    .A2(_07518_),
    .Y(_00449_),
    .B1(_07927_));
 sg13g2_and2_1 _24589_ (.A(\top_ihp.oisc.regs[1][8] ),
    .B(_07470_),
    .X(_07928_));
 sg13g2_a221oi_1 _24590_ (.B2(\top_ihp.oisc.regs[4][8] ),
    .C1(_07928_),
    .B1(_07515_),
    .A1(\top_ihp.oisc.regs[5][8] ),
    .Y(_07929_),
    .A2(_07444_));
 sg13g2_a21oi_1 _24591_ (.A1(\top_ihp.oisc.regs[15][8] ),
    .A2(net817),
    .Y(_07930_),
    .B1(net892));
 sg13g2_a22oi_1 _24592_ (.Y(_07931_),
    .B1(_07491_),
    .B2(\top_ihp.oisc.regs[11][8] ),
    .A2(_07460_),
    .A1(\top_ihp.oisc.regs[10][8] ));
 sg13g2_nand2_1 _24593_ (.Y(_07932_),
    .A(_07930_),
    .B(_07931_));
 sg13g2_a221oi_1 _24594_ (.B2(\top_ihp.oisc.regs[9][8] ),
    .C1(_07932_),
    .B1(_07488_),
    .A1(\top_ihp.oisc.regs[12][8] ),
    .Y(_07933_),
    .A2(net810));
 sg13g2_a22oi_1 _24595_ (.Y(_07934_),
    .B1(net813),
    .B2(\top_ihp.oisc.regs[13][8] ),
    .A2(_07644_),
    .A1(\top_ihp.oisc.regs[32][8] ));
 sg13g2_a22oi_1 _24596_ (.Y(_07935_),
    .B1(net811),
    .B2(\top_ihp.oisc.regs[14][8] ),
    .A2(_07682_),
    .A1(\top_ihp.oisc.regs[8][8] ));
 sg13g2_a22oi_1 _24597_ (.Y(_07936_),
    .B1(_07503_),
    .B2(\top_ihp.oisc.regs[6][8] ),
    .A2(_07473_),
    .A1(\top_ihp.oisc.regs[7][8] ));
 sg13g2_nand4_1 _24598_ (.B(_07934_),
    .C(_07935_),
    .A(_07933_),
    .Y(_07937_),
    .D(_07936_));
 sg13g2_a221oi_1 _24599_ (.B2(\top_ihp.oisc.regs[3][8] ),
    .C1(_07937_),
    .B1(_07546_),
    .A1(\top_ihp.oisc.regs[2][8] ),
    .Y(_07938_),
    .A2(net823));
 sg13g2_a221oi_1 _24600_ (.B2(_07938_),
    .C1(net860),
    .B1(_07929_),
    .A1(_00212_),
    .Y(_07939_),
    .A2(net885));
 sg13g2_mux2_1 _24601_ (.A0(_08101_),
    .A1(_07939_),
    .S(net804),
    .X(_00450_));
 sg13g2_a22oi_1 _24602_ (.Y(_07940_),
    .B1(net842),
    .B2(\top_ihp.oisc.regs[9][9] ),
    .A2(_07481_),
    .A1(\top_ihp.oisc.regs[12][9] ));
 sg13g2_a22oi_1 _24603_ (.Y(_07941_),
    .B1(net812),
    .B2(\top_ihp.oisc.regs[11][9] ),
    .A2(_07455_),
    .A1(\top_ihp.oisc.regs[15][9] ));
 sg13g2_nand2_1 _24604_ (.Y(_07942_),
    .A(_07940_),
    .B(_07941_));
 sg13g2_a21oi_1 _24605_ (.A1(\top_ihp.oisc.regs[7][9] ),
    .A2(net773),
    .Y(_07943_),
    .B1(_07942_));
 sg13g2_a22oi_1 _24606_ (.Y(_07944_),
    .B1(net863),
    .B2(\top_ihp.oisc.regs[8][9] ),
    .A2(net862),
    .A1(\top_ihp.oisc.regs[32][9] ));
 sg13g2_a22oi_1 _24607_ (.Y(_07945_),
    .B1(net822),
    .B2(\top_ihp.oisc.regs[14][9] ),
    .A2(net839),
    .A1(\top_ihp.oisc.regs[10][9] ));
 sg13g2_inv_1 _24608_ (.Y(_07946_),
    .A(_00213_));
 sg13g2_a22oi_1 _24609_ (.Y(_07947_),
    .B1(_07497_),
    .B2(_07946_),
    .A2(_07477_),
    .A1(\top_ihp.oisc.regs[13][9] ));
 sg13g2_nand3_1 _24610_ (.B(_07945_),
    .C(_07947_),
    .A(_07944_),
    .Y(_07948_));
 sg13g2_a221oi_1 _24611_ (.B2(\top_ihp.oisc.regs[2][9] ),
    .C1(_07948_),
    .B1(net815),
    .A1(\top_ihp.oisc.regs[3][9] ),
    .Y(_07949_),
    .A2(_07507_));
 sg13g2_a22oi_1 _24612_ (.Y(_07950_),
    .B1(net772),
    .B2(\top_ihp.oisc.regs[6][9] ),
    .A2(net828),
    .A1(\top_ihp.oisc.regs[1][9] ));
 sg13g2_a22oi_1 _24613_ (.Y(_07951_),
    .B1(net791),
    .B2(\top_ihp.oisc.regs[4][9] ),
    .A2(_07443_),
    .A1(\top_ihp.oisc.regs[5][9] ));
 sg13g2_nand4_1 _24614_ (.B(_07949_),
    .C(_07950_),
    .A(_07943_),
    .Y(_07952_),
    .D(_07951_));
 sg13g2_a21oi_1 _24615_ (.A1(_07437_),
    .A2(_07952_),
    .Y(_07953_),
    .B1(net760));
 sg13g2_a21oi_1 _24616_ (.A1(_10506_),
    .A2(net744),
    .Y(_00451_),
    .B1(_07953_));
 sg13g2_a21oi_1 _24617_ (.A1(_08304_),
    .A2(_08359_),
    .Y(_00323_),
    .B1(_09605_));
 sg13g2_mux4_1 _24618_ (.S0(_08642_),
    .A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[0] ),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[1] ),
    .A2(\top_ihp.wb_uart.uart_tx.tx_data_latch[2] ),
    .A3(\top_ihp.wb_uart.uart_tx.tx_data_latch[3] ),
    .S1(_08643_),
    .X(_07954_));
 sg13g2_mux4_1 _24619_ (.S0(_08642_),
    .A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[4] ),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[5] ),
    .A2(\top_ihp.wb_uart.uart_tx.tx_data_latch[6] ),
    .A3(\top_ihp.wb_uart.uart_tx.tx_data_latch[7] ),
    .S1(_08643_),
    .X(_07955_));
 sg13g2_mux2_1 _24620_ (.A0(_07954_),
    .A1(_07955_),
    .S(\top_ihp.wb_uart.uart_tx.bit_cnt[2] ),
    .X(_07956_));
 sg13g2_nand2b_1 _24621_ (.Y(_07957_),
    .B(_08637_),
    .A_N(_08639_));
 sg13g2_o21ai_1 _24622_ (.B1(_07957_),
    .Y(_00324_),
    .A1(_05175_),
    .A2(_07956_));
 sg13g2_nor2_1 _24623_ (.A(net982),
    .B(net2133),
    .Y(\top_ihp.ram_clk_o ));
 sg13g2_and2_1 _24624_ (.A(net943),
    .B(\top_ihp.wb_emem.cmd[63] ),
    .X(\top_ihp.ram_data_o ));
 sg13g2_nor2_1 _24625_ (.A(net2132),
    .B(\top_ihp.rom_cs_o ),
    .Y(\top_ihp.rom_clk_o ));
 sg13g2_and2_1 _24626_ (.A(_08366_),
    .B(\top_ihp.wb_dati_rom[7] ),
    .X(\top_ihp.rom_data_o ));
 sg13g2_and2_1 _24627_ (.A(_08195_),
    .B(\top_ihp.wb_dati_spi[31] ),
    .X(\top_ihp.spi_data_o ));
 sg13g2_inv_1 _14561__1 (.Y(net2016),
    .A(clknet_leaf_18_clk));
 sg13g2_buf_1 _24629_ (.A(net1431),
    .X(uio_oe[0]));
 sg13g2_buf_1 _24630_ (.A(net1432),
    .X(uio_oe[1]));
 sg13g2_buf_1 _24631_ (.A(net1433),
    .X(uio_oe[2]));
 sg13g2_buf_1 _24632_ (.A(net1434),
    .X(uio_oe[3]));
 sg13g2_buf_1 _24633_ (.A(net1435),
    .X(uio_oe[4]));
 sg13g2_buf_1 _24634_ (.A(net1436),
    .X(uio_oe[5]));
 sg13g2_buf_1 _24635_ (.A(net1437),
    .X(uio_oe[6]));
 sg13g2_buf_1 _24636_ (.A(net1438),
    .X(uio_oe[7]));
 sg13g2_buf_1 _24637_ (.A(\top_ihp.spi_data_o ),
    .X(net10));
 sg13g2_buf_1 _24638_ (.A(\top_ihp.spi_cs_o_1 ),
    .X(net11));
 sg13g2_buf_1 _24639_ (.A(\top_ihp.spi_cs_o_2 ),
    .X(net12));
 sg13g2_buf_1 _24640_ (.A(\top_ihp.spi_cs_o_3 ),
    .X(net13));
 sg13g2_buf_1 _24641_ (.A(\top_ihp.gpio_o_1 ),
    .X(net14));
 sg13g2_buf_1 _24642_ (.A(\top_ihp.gpio_o_2 ),
    .X(net15));
 sg13g2_buf_1 _24643_ (.A(\top_ihp.gpio_o_3 ),
    .X(net16));
 sg13g2_buf_1 _24644_ (.A(\top_ihp.gpio_o_4 ),
    .X(net17));
 sg13g2_buf_1 _24645_ (.A(\top_ihp.tx ),
    .X(net18));
 sg13g2_buf_1 _24646_ (.A(\top_ihp.rom_clk_o ),
    .X(net19));
 sg13g2_buf_1 _24647_ (.A(\top_ihp.rom_data_o ),
    .X(net20));
 sg13g2_buf_1 _24648_ (.A(\top_ihp.rom_cs_o ),
    .X(net21));
 sg13g2_buf_1 _24649_ (.A(\top_ihp.ram_clk_o ),
    .X(net22));
 sg13g2_buf_1 _24650_ (.A(\top_ihp.ram_data_o ),
    .X(net23));
 sg13g2_buf_1 _24651_ (.A(\top_ihp.ram_cs_o ),
    .X(net24));
 sg13g2_buf_1 _24652_ (.A(\top_ihp.spi_clk_o ),
    .X(net25));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1141),
    .D(_00325_),
    .Q_N(_13522_),
    .Q(\top_ihp.oisc.decoder.decoded[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1145),
    .D(_00326_),
    .Q_N(_13521_),
    .Q(\top_ihp.oisc.decoder.decoded[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1145),
    .D(_00327_),
    .Q_N(_13520_),
    .Q(\top_ihp.oisc.decoder.decoded[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1146),
    .D(_00328_),
    .Q_N(_13519_),
    .Q(\top_ihp.oisc.decoder.decoded[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1146),
    .D(_00329_),
    .Q_N(_13518_),
    .Q(\top_ihp.oisc.decoder.decoded[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1146),
    .D(_00330_),
    .Q_N(_13517_),
    .Q(\top_ihp.oisc.decoder.decoded[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1146),
    .D(_00331_),
    .Q_N(_00085_),
    .Q(\top_ihp.oisc.decoder.decoded[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1141),
    .D(_00332_),
    .Q_N(_13516_),
    .Q(\top_ihp.oisc.decoder.decoded[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1141),
    .D(_00333_),
    .Q_N(_13515_),
    .Q(\top_ihp.oisc.decoder.decoded[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1145),
    .D(_00334_),
    .Q_N(_13514_),
    .Q(\top_ihp.oisc.decoder.decoded[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1141),
    .D(_00335_),
    .Q_N(_13513_),
    .Q(\top_ihp.oisc.decoder.decoded[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1141),
    .D(_00336_),
    .Q_N(_13512_),
    .Q(\top_ihp.oisc.decoder.decoded[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1145),
    .D(_00337_),
    .Q_N(_13511_),
    .Q(\top_ihp.oisc.decoder.decoded[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1145),
    .D(_00338_),
    .Q_N(_13510_),
    .Q(\top_ihp.oisc.decoder.decoded[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1144),
    .D(_00339_),
    .Q_N(_13509_),
    .Q(\top_ihp.oisc.decoder.instruction[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1144),
    .D(_00340_),
    .Q_N(_13508_),
    .Q(\top_ihp.oisc.decoder.instruction[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1144),
    .D(_00341_),
    .Q_N(_13507_),
    .Q(\top_ihp.oisc.decoder.instruction[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1143),
    .D(_00342_),
    .Q_N(_13506_),
    .Q(\top_ihp.oisc.decoder.instruction[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1143),
    .D(_00343_),
    .Q_N(_00074_),
    .Q(\top_ihp.oisc.decoder.instruction[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1143),
    .D(_00204_),
    .Q_N(_13505_),
    .Q(\top_ihp.oisc.decoder.instruction[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[16]$_DFFE_PN0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1143),
    .D(_00344_),
    .Q_N(_00200_),
    .Q(\top_ihp.oisc.decoder.instruction[16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[17]$_DFFE_PN0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1143),
    .D(_00345_),
    .Q_N(_00201_),
    .Q(\top_ihp.oisc.decoder.instruction[17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[18]$_DFFE_PN0N_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1131),
    .D(_00346_),
    .Q_N(_00202_),
    .Q(\top_ihp.oisc.decoder.instruction[18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[19]$_DFFE_PN0N_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1132),
    .D(_00347_),
    .Q_N(_00203_),
    .Q(\top_ihp.oisc.decoder.instruction[19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[20]$_DFFE_PN0N_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1144),
    .D(_00348_),
    .Q_N(_13504_),
    .Q(\top_ihp.oisc.decoder.instruction[20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[21]$_DFFE_PN0N_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1147),
    .D(_00349_),
    .Q_N(_00196_),
    .Q(\top_ihp.oisc.decoder.instruction[21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[22]$_DFFE_PN0N_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1144),
    .D(_00350_),
    .Q_N(_00197_),
    .Q(\top_ihp.oisc.decoder.instruction[22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[23]$_DFFE_PN0N_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1144),
    .D(_00351_),
    .Q_N(_00198_),
    .Q(\top_ihp.oisc.decoder.instruction[23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[24]$_DFFE_PN0N_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1143),
    .D(_00352_),
    .Q_N(_00199_),
    .Q(\top_ihp.oisc.decoder.instruction[24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[25]$_DFFE_PN0N_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1143),
    .D(_00353_),
    .Q_N(_13503_),
    .Q(\top_ihp.oisc.decoder.instruction[25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[26]$_DFFE_PN0N_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1145),
    .D(_00354_),
    .Q_N(_13502_),
    .Q(\top_ihp.oisc.decoder.instruction[26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[27]$_DFFE_PN0N_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1143),
    .D(_00355_),
    .Q_N(_13501_),
    .Q(\top_ihp.oisc.decoder.instruction[27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[28]$_DFFE_PN0N_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1148),
    .D(_00356_),
    .Q_N(_13500_),
    .Q(\top_ihp.oisc.decoder.instruction[28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[29]$_DFFE_PN0N_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1148),
    .D(_00357_),
    .Q_N(_13499_),
    .Q(\top_ihp.oisc.decoder.instruction[29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[30]$_DFFE_PN0N_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1144),
    .D(_00358_),
    .Q_N(_13498_),
    .Q(\top_ihp.oisc.decoder.instruction[30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[31]$_DFFE_PN0N_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1146),
    .D(_00359_),
    .Q_N(_13497_),
    .Q(\top_ihp.oisc.decoder.instruction[31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1145),
    .D(_00360_),
    .Q_N(_13496_),
    .Q(\top_ihp.oisc.decoder.instruction[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1148),
    .D(_00361_),
    .Q_N(_13495_),
    .Q(\top_ihp.oisc.decoder.instruction[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1144),
    .D(_00362_),
    .Q_N(_13523_),
    .Q(\top_ihp.oisc.decoder.instruction[9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.mem_addr_lowbits[0]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1439),
    .D(\top_ihp.oisc.wb_adr_o[0] ),
    .Q_N(_13524_),
    .Q(\top_ihp.oisc.mem_addr_lowbits[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.mem_addr_lowbits[1]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1440),
    .D(\top_ihp.oisc.wb_adr_o[1] ),
    .Q_N(_13494_),
    .Q(\top_ihp.oisc.mem_addr_lowbits[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1108),
    .D(_00363_),
    .Q_N(_13493_),
    .Q(\top_ihp.oisc.micro_op[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1108),
    .D(_00364_),
    .Q_N(_13492_),
    .Q(\top_ihp.oisc.micro_op[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1109),
    .D(_00365_),
    .Q_N(_13491_),
    .Q(\top_ihp.oisc.micro_op[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1159),
    .D(_00366_),
    .Q_N(_13490_),
    .Q(\top_ihp.oisc.micro_op[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1109),
    .D(_00367_),
    .Q_N(_13489_),
    .Q(\top_ihp.oisc.micro_op[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1108),
    .D(_00368_),
    .Q_N(_13488_),
    .Q(\top_ihp.oisc.micro_op[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1108),
    .D(_00369_),
    .Q_N(_13487_),
    .Q(\top_ihp.oisc.micro_op[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1108),
    .D(_00370_),
    .Q_N(_13486_),
    .Q(\top_ihp.oisc.micro_op[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1109),
    .D(_00371_),
    .Q_N(_13485_),
    .Q(\top_ihp.oisc.micro_op[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1109),
    .D(_00372_),
    .Q_N(_13484_),
    .Q(\top_ihp.oisc.micro_op[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1109),
    .D(_00373_),
    .Q_N(_13483_),
    .Q(\top_ihp.oisc.micro_op[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1109),
    .D(_00374_),
    .Q_N(_13482_),
    .Q(\top_ihp.oisc.micro_op[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1108),
    .D(_00375_),
    .Q_N(_13481_),
    .Q(\top_ihp.oisc.micro_op[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1108),
    .D(_00376_),
    .Q_N(_13480_),
    .Q(\top_ihp.oisc.micro_op[9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[0]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1441),
    .D(_00377_),
    .Q_N(_00181_),
    .Q(\top_ihp.oisc.micro_pc[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[1]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1442),
    .D(_00378_),
    .Q_N(_00182_),
    .Q(\top_ihp.oisc.micro_pc[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[2]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1443),
    .D(_00379_),
    .Q_N(_00180_),
    .Q(\top_ihp.oisc.micro_pc[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[3]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1444),
    .D(_00380_),
    .Q_N(_00179_),
    .Q(\top_ihp.oisc.micro_pc[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[4]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1445),
    .D(_00381_),
    .Q_N(_00178_),
    .Q(\top_ihp.oisc.micro_pc[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[5]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1446),
    .D(_00382_),
    .Q_N(_00177_),
    .Q(\top_ihp.oisc.micro_pc[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[6]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1447),
    .D(_00383_),
    .Q_N(_00176_),
    .Q(\top_ihp.oisc.micro_pc[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[7]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1448),
    .D(_00384_),
    .Q_N(_00175_),
    .Q(\top_ihp.oisc.micro_pc[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_res_addr[0]$_DFF_PN0_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1157),
    .D(\top_ihp.oisc.reg_rb[0] ),
    .Q_N(_13525_),
    .Q(\top_ihp.oisc.micro_res_addr[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_res_addr[1]$_DFF_PN0_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1158),
    .D(\top_ihp.oisc.reg_rb[1] ),
    .Q_N(_13526_),
    .Q(\top_ihp.oisc.micro_res_addr[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_res_addr[2]$_DFF_PN0_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1147),
    .D(\top_ihp.oisc.reg_rb[2] ),
    .Q_N(_13527_),
    .Q(\top_ihp.oisc.micro_res_addr[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_res_addr[3]$_DFF_PN0_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1158),
    .D(\top_ihp.oisc.reg_rb[3] ),
    .Q_N(_13479_),
    .Q(\top_ihp.oisc.micro_res_addr[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_state[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1146),
    .D(_00385_),
    .Q_N(\top_ihp.oisc.micro_state[0] ),
    .Q(_13599_));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_state[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1146),
    .D(_00386_),
    .Q_N(_13478_),
    .Q(\top_ihp.oisc.micro_state[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_state[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1146),
    .D(_00387_),
    .Q_N(_13477_),
    .Q(\top_ihp.oisc.micro_state[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1219),
    .D(_00388_),
    .Q_N(_13476_),
    .Q(\top_ihp.oisc.op_a[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1248),
    .D(_00389_),
    .Q_N(_13475_),
    .Q(\top_ihp.oisc.op_a[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1219),
    .D(_00390_),
    .Q_N(_13474_),
    .Q(\top_ihp.oisc.op_a[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1219),
    .D(_00391_),
    .Q_N(_13473_),
    .Q(\top_ihp.oisc.op_a[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1153),
    .D(_00392_),
    .Q_N(_13472_),
    .Q(\top_ihp.oisc.op_a[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1222),
    .D(_00393_),
    .Q_N(_13471_),
    .Q(\top_ihp.oisc.op_a[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1152),
    .D(_00394_),
    .Q_N(_13470_),
    .Q(\top_ihp.oisc.op_a[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[16]$_DFFE_PN0N_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1219),
    .D(_00395_),
    .Q_N(_13469_),
    .Q(\top_ihp.oisc.op_a[16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[17]$_DFFE_PN0N_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1225),
    .D(_00396_),
    .Q_N(_13468_),
    .Q(\top_ihp.oisc.op_a[17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[18]$_DFFE_PN0N_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1225),
    .D(_00397_),
    .Q_N(_13467_),
    .Q(\top_ihp.oisc.op_a[18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[19]$_DFFE_PN0N_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1155),
    .D(_00398_),
    .Q_N(_13466_),
    .Q(\top_ihp.oisc.op_a[19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1182),
    .D(_00399_),
    .Q_N(_13465_),
    .Q(\top_ihp.oisc.op_a[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[20]$_DFFE_PN0N_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1240),
    .D(_00400_),
    .Q_N(_13464_),
    .Q(\top_ihp.oisc.op_a[20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[21]$_DFFE_PN0N_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1173),
    .D(_00401_),
    .Q_N(_13463_),
    .Q(\top_ihp.oisc.op_a[21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[22]$_DFFE_PN0N_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1226),
    .D(_00402_),
    .Q_N(_13462_),
    .Q(\top_ihp.oisc.op_a[22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[23]$_DFFE_PN0N_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1223),
    .D(_00403_),
    .Q_N(_13461_),
    .Q(\top_ihp.oisc.op_a[23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[24]$_DFFE_PN0N_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1240),
    .D(_00404_),
    .Q_N(_13460_),
    .Q(\top_ihp.oisc.op_a[24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[25]$_DFFE_PN0N_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1182),
    .D(_00405_),
    .Q_N(_13459_),
    .Q(\top_ihp.oisc.op_a[25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[26]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1150),
    .D(_00406_),
    .Q_N(_13458_),
    .Q(\top_ihp.oisc.op_a[26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[27]$_DFFE_PN0N_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1240),
    .D(_00407_),
    .Q_N(_13457_),
    .Q(\top_ihp.oisc.op_a[27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[28]$_DFFE_PN0N_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1162),
    .D(_00408_),
    .Q_N(_13456_),
    .Q(\top_ihp.oisc.op_a[28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[29]$_DFFE_PN0N_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1235),
    .D(_00409_),
    .Q_N(_13455_),
    .Q(\top_ihp.oisc.op_a[29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1245),
    .D(_00410_),
    .Q_N(_13454_),
    .Q(\top_ihp.oisc.op_a[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[30]$_DFFE_PN0N_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1157),
    .D(_00411_),
    .Q_N(_13453_),
    .Q(\top_ihp.oisc.op_a[30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[31]$_DFFE_PN0N_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1158),
    .D(_00412_),
    .Q_N(_13452_),
    .Q(\top_ihp.oisc.op_a[31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1162),
    .D(_00413_),
    .Q_N(_13451_),
    .Q(\top_ihp.oisc.op_a[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1162),
    .D(_00414_),
    .Q_N(_13450_),
    .Q(\top_ihp.oisc.op_a[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1158),
    .D(_00415_),
    .Q_N(_13449_),
    .Q(\top_ihp.oisc.op_a[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1244),
    .D(_00416_),
    .Q_N(_13448_),
    .Q(\top_ihp.oisc.op_a[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1163),
    .D(_00417_),
    .Q_N(_13447_),
    .Q(\top_ihp.oisc.op_a[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1240),
    .D(_00418_),
    .Q_N(_13446_),
    .Q(\top_ihp.oisc.op_a[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1240),
    .D(_00419_),
    .Q_N(_13445_),
    .Q(\top_ihp.oisc.op_a[9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1159),
    .D(_00420_),
    .Q_N(_13444_),
    .Q(\top_ihp.oisc.op_b[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1152),
    .D(_00421_),
    .Q_N(_13443_),
    .Q(\top_ihp.oisc.op_b[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1152),
    .D(_00422_),
    .Q_N(_13442_),
    .Q(\top_ihp.oisc.op_b[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1152),
    .D(_00423_),
    .Q_N(_13441_),
    .Q(\top_ihp.oisc.op_b[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1152),
    .D(_00424_),
    .Q_N(_13440_),
    .Q(\top_ihp.oisc.op_b[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1152),
    .D(_00425_),
    .Q_N(_13439_),
    .Q(\top_ihp.oisc.op_b[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1152),
    .D(_00426_),
    .Q_N(_13438_),
    .Q(\top_ihp.oisc.op_b[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[16]$_DFFE_PN0N_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1152),
    .D(_00427_),
    .Q_N(_13437_),
    .Q(\top_ihp.oisc.op_b[16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[17]$_DFFE_PN0N_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1150),
    .D(_00428_),
    .Q_N(_13436_),
    .Q(\top_ihp.oisc.op_b[17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[18]$_DFFE_PN0N_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1151),
    .D(_00429_),
    .Q_N(_13435_),
    .Q(\top_ihp.oisc.op_b[18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[19]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1151),
    .D(_00430_),
    .Q_N(_13434_),
    .Q(\top_ihp.oisc.op_b[19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1159),
    .D(_00431_),
    .Q_N(_13433_),
    .Q(\top_ihp.oisc.op_b[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[20]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1150),
    .D(_00432_),
    .Q_N(_13432_),
    .Q(\top_ihp.oisc.op_b[20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[21]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1150),
    .D(_00433_),
    .Q_N(_13431_),
    .Q(\top_ihp.oisc.op_b[21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[22]$_DFFE_PN0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1150),
    .D(_00434_),
    .Q_N(_13430_),
    .Q(\top_ihp.oisc.op_b[22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[23]$_DFFE_PN0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1150),
    .D(_00435_),
    .Q_N(_13429_),
    .Q(\top_ihp.oisc.op_b[23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[24]$_DFFE_PN0N_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1150),
    .D(_00436_),
    .Q_N(_13428_),
    .Q(\top_ihp.oisc.op_b[24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[25]$_DFFE_PN0N_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1150),
    .D(_00437_),
    .Q_N(_13427_),
    .Q(\top_ihp.oisc.op_b[25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[26]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1151),
    .D(_00438_),
    .Q_N(_13426_),
    .Q(\top_ihp.oisc.op_b[26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[27]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1151),
    .D(_00439_),
    .Q_N(_13425_),
    .Q(\top_ihp.oisc.op_b[27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[28]$_DFFE_PN0N_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1159),
    .D(_00440_),
    .Q_N(_13424_),
    .Q(\top_ihp.oisc.op_b[28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[29]$_DFFE_PN0N_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1159),
    .D(_00441_),
    .Q_N(_13423_),
    .Q(\top_ihp.oisc.op_b[29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1159),
    .D(_00442_),
    .Q_N(_13422_),
    .Q(\top_ihp.oisc.op_b[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[30]$_DFFE_PN0N_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1157),
    .D(_00443_),
    .Q_N(_13421_),
    .Q(\top_ihp.oisc.op_b[30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[31]$_DFFE_PN0N_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1157),
    .D(_00444_),
    .Q_N(_13420_),
    .Q(\top_ihp.oisc.op_b[31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1159),
    .D(_00445_),
    .Q_N(_13419_),
    .Q(\top_ihp.oisc.op_b[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1158),
    .D(_00446_),
    .Q_N(_13418_),
    .Q(\top_ihp.oisc.op_b[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1164),
    .D(_00447_),
    .Q_N(_13417_),
    .Q(\top_ihp.oisc.op_b[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1164),
    .D(_00448_),
    .Q_N(_13416_),
    .Q(\top_ihp.oisc.op_b[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1157),
    .D(_00449_),
    .Q_N(_13415_),
    .Q(\top_ihp.oisc.op_b[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1159),
    .D(_00450_),
    .Q_N(_13414_),
    .Q(\top_ihp.oisc.op_b[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1151),
    .D(_00451_),
    .Q_N(_13413_),
    .Q(\top_ihp.oisc.op_b[9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1219),
    .D(_00452_),
    .Q_N(_13412_),
    .Q(\top_ihp.oisc.regs[0][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1221),
    .D(_00453_),
    .Q_N(_00214_),
    .Q(\top_ihp.oisc.regs[0][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1219),
    .D(_00454_),
    .Q_N(_00215_),
    .Q(\top_ihp.oisc.regs[0][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1221),
    .D(_00455_),
    .Q_N(_00216_),
    .Q(\top_ihp.oisc.regs[0][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1219),
    .D(_00456_),
    .Q_N(_00217_),
    .Q(\top_ihp.oisc.regs[0][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1221),
    .D(_00457_),
    .Q_N(_00218_),
    .Q(\top_ihp.oisc.regs[0][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1222),
    .D(_00458_),
    .Q_N(_00219_),
    .Q(\top_ihp.oisc.regs[0][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1220),
    .D(_00459_),
    .Q_N(_00220_),
    .Q(\top_ihp.oisc.regs[0][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1223),
    .D(_00460_),
    .Q_N(_00221_),
    .Q(\top_ihp.oisc.regs[0][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1223),
    .D(_00461_),
    .Q_N(_00222_),
    .Q(\top_ihp.oisc.regs[0][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1172),
    .D(_00462_),
    .Q_N(_00223_),
    .Q(\top_ihp.oisc.regs[0][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1223),
    .D(_00463_),
    .Q_N(_00205_),
    .Q(\top_ihp.oisc.regs[0][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1239),
    .D(_00464_),
    .Q_N(_00224_),
    .Q(\top_ihp.oisc.regs[0][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1173),
    .D(_00465_),
    .Q_N(_00225_),
    .Q(\top_ihp.oisc.regs[0][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1224),
    .D(_00466_),
    .Q_N(_00226_),
    .Q(\top_ihp.oisc.regs[0][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1224),
    .D(_00467_),
    .Q_N(_00227_),
    .Q(\top_ihp.oisc.regs[0][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1239),
    .D(_00468_),
    .Q_N(_00228_),
    .Q(\top_ihp.oisc.regs[0][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1179),
    .D(_00469_),
    .Q_N(_00229_),
    .Q(\top_ihp.oisc.regs[0][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1199),
    .D(_00470_),
    .Q_N(_00230_),
    .Q(\top_ihp.oisc.regs[0][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1239),
    .D(_00471_),
    .Q_N(_00231_),
    .Q(\top_ihp.oisc.regs[0][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1200),
    .D(_00472_),
    .Q_N(_00069_),
    .Q(\top_ihp.oisc.regs[0][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1203),
    .D(_00473_),
    .Q_N(_00070_),
    .Q(\top_ihp.oisc.regs[0][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1243),
    .D(_00474_),
    .Q_N(_00206_),
    .Q(\top_ihp.oisc.regs[0][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1194),
    .D(_00475_),
    .Q_N(_00071_),
    .Q(\top_ihp.oisc.regs[0][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1200),
    .D(_00476_),
    .Q_N(_00072_),
    .Q(\top_ihp.oisc.regs[0][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1192),
    .D(_00477_),
    .Q_N(_00207_),
    .Q(\top_ihp.oisc.regs[0][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1161),
    .D(_00478_),
    .Q_N(_00208_),
    .Q(\top_ihp.oisc.regs[0][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1192),
    .D(_00479_),
    .Q_N(_00209_),
    .Q(\top_ihp.oisc.regs[0][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1243),
    .D(_00480_),
    .Q_N(_00210_),
    .Q(\top_ihp.oisc.regs[0][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1243),
    .D(_00481_),
    .Q_N(_00211_),
    .Q(\top_ihp.oisc.regs[0][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1239),
    .D(_00482_),
    .Q_N(_00212_),
    .Q(\top_ihp.oisc.regs[0][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1226),
    .D(_00483_),
    .Q_N(_00213_),
    .Q(\top_ihp.oisc.regs[0][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][0]$_DFFE_PN1P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1213),
    .D(_00484_),
    .Q_N(\top_ihp.oisc.regs[10][0] ),
    .Q(_00235_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1165),
    .D(_00485_),
    .Q_N(_13411_),
    .Q(\top_ihp.oisc.regs[10][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1175),
    .D(_00486_),
    .Q_N(_13410_),
    .Q(\top_ihp.oisc.regs[10][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1176),
    .D(_00487_),
    .Q_N(_13409_),
    .Q(\top_ihp.oisc.regs[10][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1165),
    .D(_00488_),
    .Q_N(_13408_),
    .Q(\top_ihp.oisc.regs[10][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1209),
    .D(_00489_),
    .Q_N(_13407_),
    .Q(\top_ihp.oisc.regs[10][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1177),
    .D(_00490_),
    .Q_N(_13406_),
    .Q(\top_ihp.oisc.regs[10][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1209),
    .D(_00491_),
    .Q_N(_13405_),
    .Q(\top_ihp.oisc.regs[10][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1213),
    .D(_00492_),
    .Q_N(_13404_),
    .Q(\top_ihp.oisc.regs[10][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1179),
    .D(_00493_),
    .Q_N(_13403_),
    .Q(\top_ihp.oisc.regs[10][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1170),
    .D(_00494_),
    .Q_N(_13402_),
    .Q(\top_ihp.oisc.regs[10][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1182),
    .D(_00495_),
    .Q_N(_13401_),
    .Q(\top_ihp.oisc.regs[10][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1198),
    .D(_00496_),
    .Q_N(_13400_),
    .Q(\top_ihp.oisc.regs[10][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1173),
    .D(_00497_),
    .Q_N(_13399_),
    .Q(\top_ihp.oisc.regs[10][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1213),
    .D(_00498_),
    .Q_N(_13398_),
    .Q(\top_ihp.oisc.regs[10][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1180),
    .D(_00499_),
    .Q_N(_13397_),
    .Q(\top_ihp.oisc.regs[10][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1229),
    .D(_00500_),
    .Q_N(_13396_),
    .Q(\top_ihp.oisc.regs[10][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1180),
    .D(_00501_),
    .Q_N(_13395_),
    .Q(\top_ihp.oisc.regs[10][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1198),
    .D(_00502_),
    .Q_N(_13394_),
    .Q(\top_ihp.oisc.regs[10][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1196),
    .D(_00503_),
    .Q_N(_13393_),
    .Q(\top_ihp.oisc.regs[10][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1203),
    .D(_00504_),
    .Q_N(_13392_),
    .Q(\top_ihp.oisc.regs[10][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1204),
    .D(_00505_),
    .Q_N(_13391_),
    .Q(\top_ihp.oisc.regs[10][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1235),
    .D(_00506_),
    .Q_N(_13390_),
    .Q(\top_ihp.oisc.regs[10][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1192),
    .D(_00507_),
    .Q_N(_13389_),
    .Q(\top_ihp.oisc.regs[10][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1191),
    .D(_00508_),
    .Q_N(_13388_),
    .Q(\top_ihp.oisc.regs[10][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1186),
    .D(_00509_),
    .Q_N(_13387_),
    .Q(\top_ihp.oisc.regs[10][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1191),
    .D(_00510_),
    .Q_N(_13386_),
    .Q(\top_ihp.oisc.regs[10][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1161),
    .D(_00511_),
    .Q_N(_13385_),
    .Q(\top_ihp.oisc.regs[10][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1234),
    .D(_00512_),
    .Q_N(_13384_),
    .Q(\top_ihp.oisc.regs[10][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1234),
    .D(_00513_),
    .Q_N(_13383_),
    .Q(\top_ihp.oisc.regs[10][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1230),
    .D(_00514_),
    .Q_N(_13382_),
    .Q(\top_ihp.oisc.regs[10][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1214),
    .D(_00515_),
    .Q_N(_13381_),
    .Q(\top_ihp.oisc.regs[10][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][0]$_DFFE_PN1P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1213),
    .D(_00516_),
    .Q_N(\top_ihp.oisc.regs[11][0] ),
    .Q(_00236_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1153),
    .D(_00517_),
    .Q_N(_13380_),
    .Q(\top_ihp.oisc.regs[11][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1167),
    .D(_00518_),
    .Q_N(_13379_),
    .Q(\top_ihp.oisc.regs[11][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1175),
    .D(_00519_),
    .Q_N(_13378_),
    .Q(\top_ihp.oisc.regs[11][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1153),
    .D(_00520_),
    .Q_N(_13377_),
    .Q(\top_ihp.oisc.regs[11][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1208),
    .D(_00521_),
    .Q_N(_13376_),
    .Q(\top_ihp.oisc.regs[11][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1209),
    .D(_00522_),
    .Q_N(_13375_),
    .Q(\top_ihp.oisc.regs[11][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1209),
    .D(_00523_),
    .Q_N(_13374_),
    .Q(\top_ihp.oisc.regs[11][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1153),
    .D(_00524_),
    .Q_N(_13373_),
    .Q(\top_ihp.oisc.regs[11][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1179),
    .D(_00525_),
    .Q_N(_13372_),
    .Q(\top_ihp.oisc.regs[11][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1154),
    .D(_00526_),
    .Q_N(_13371_),
    .Q(\top_ihp.oisc.regs[11][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][1]$_DFFE_PN1P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1180),
    .D(_00527_),
    .Q_N(\top_ihp.oisc.regs[11][1] ),
    .Q(_00237_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1229),
    .D(_00528_),
    .Q_N(_13370_),
    .Q(\top_ihp.oisc.regs[11][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1186),
    .D(_00529_),
    .Q_N(_13369_),
    .Q(\top_ihp.oisc.regs[11][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1214),
    .D(_00530_),
    .Q_N(_13368_),
    .Q(\top_ihp.oisc.regs[11][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1214),
    .D(_00531_),
    .Q_N(_13367_),
    .Q(\top_ihp.oisc.regs[11][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1229),
    .D(_00532_),
    .Q_N(_13366_),
    .Q(\top_ihp.oisc.regs[11][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1180),
    .D(_00533_),
    .Q_N(_13365_),
    .Q(\top_ihp.oisc.regs[11][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1198),
    .D(_00534_),
    .Q_N(_13364_),
    .Q(\top_ihp.oisc.regs[11][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1196),
    .D(_00535_),
    .Q_N(_13363_),
    .Q(\top_ihp.oisc.regs[11][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1203),
    .D(_00536_),
    .Q_N(_13362_),
    .Q(\top_ihp.oisc.regs[11][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1204),
    .D(_00537_),
    .Q_N(_13361_),
    .Q(\top_ihp.oisc.regs[11][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][2]$_DFFE_PN1P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1237),
    .D(_00538_),
    .Q_N(\top_ihp.oisc.regs[11][2] ),
    .Q(_00238_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1193),
    .D(_00539_),
    .Q_N(_13360_),
    .Q(\top_ihp.oisc.regs[11][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1191),
    .D(_00540_),
    .Q_N(_13359_),
    .Q(\top_ihp.oisc.regs[11][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][3]$_DFFE_PN1P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1189),
    .D(_00541_),
    .Q_N(\top_ihp.oisc.regs[11][3] ),
    .Q(_00239_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][4]$_DFFE_PN1P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1161),
    .D(_00542_),
    .Q_N(\top_ihp.oisc.regs[11][4] ),
    .Q(_00240_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1192),
    .D(_00543_),
    .Q_N(_13358_),
    .Q(\top_ihp.oisc.regs[11][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1230),
    .D(_00544_),
    .Q_N(_13357_),
    .Q(\top_ihp.oisc.regs[11][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1236),
    .D(_00545_),
    .Q_N(_13356_),
    .Q(\top_ihp.oisc.regs[11][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1232),
    .D(_00546_),
    .Q_N(_13355_),
    .Q(\top_ihp.oisc.regs[11][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1232),
    .D(_00547_),
    .Q_N(_13354_),
    .Q(\top_ihp.oisc.regs[11][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][0]$_DFFE_PN1P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1213),
    .D(_00548_),
    .Q_N(\top_ihp.oisc.regs[12][0] ),
    .Q(_00241_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][10]$_DFFE_PN1P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1166),
    .D(_00549_),
    .Q_N(\top_ihp.oisc.regs[12][10] ),
    .Q(_00242_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][11]$_DFFE_PN1P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1168),
    .D(_00550_),
    .Q_N(\top_ihp.oisc.regs[12][11] ),
    .Q(_00243_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][12]$_DFFE_PN1P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1153),
    .D(_00551_),
    .Q_N(\top_ihp.oisc.regs[12][12] ),
    .Q(_00244_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][13]$_DFFE_PN1P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1153),
    .D(_00552_),
    .Q_N(\top_ihp.oisc.regs[12][13] ),
    .Q(_00245_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][14]$_DFFE_PN1P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1208),
    .D(_00553_),
    .Q_N(\top_ihp.oisc.regs[12][14] ),
    .Q(_00246_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][15]$_DFFE_PN1P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1178),
    .D(_00554_),
    .Q_N(\top_ihp.oisc.regs[12][15] ),
    .Q(_00247_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][16]$_DFFE_PN1P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1178),
    .D(_00555_),
    .Q_N(\top_ihp.oisc.regs[12][16] ),
    .Q(_00248_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][17]$_DFFE_PN1P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1154),
    .D(_00556_),
    .Q_N(\top_ihp.oisc.regs[12][17] ),
    .Q(_00249_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][18]$_DFFE_PN1P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1154),
    .D(_00557_),
    .Q_N(\top_ihp.oisc.regs[12][18] ),
    .Q(_00250_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][19]$_DFFE_PN1P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1154),
    .D(_00558_),
    .Q_N(\top_ihp.oisc.regs[12][19] ),
    .Q(_00251_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][1]$_DFFE_PN1P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1179),
    .D(_00559_),
    .Q_N(\top_ihp.oisc.regs[12][1] ),
    .Q(_00252_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][20]$_DFFE_PN1P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1197),
    .D(_00560_),
    .Q_N(\top_ihp.oisc.regs[12][20] ),
    .Q(_00253_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][21]$_DFFE_PN1P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1154),
    .D(_00561_),
    .Q_N(\top_ihp.oisc.regs[12][21] ),
    .Q(_00254_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][22]$_DFFE_PN1P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1214),
    .D(_00562_),
    .Q_N(\top_ihp.oisc.regs[12][22] ),
    .Q(_00255_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][23]$_DFFE_PN1P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1155),
    .D(_00563_),
    .Q_N(\top_ihp.oisc.regs[12][23] ),
    .Q(_00256_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][24]$_DFFE_PN1P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1229),
    .D(_00564_),
    .Q_N(\top_ihp.oisc.regs[12][24] ),
    .Q(_00257_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][25]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1155),
    .D(_00565_),
    .Q_N(\top_ihp.oisc.regs[12][25] ),
    .Q(_00258_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][26]$_DFFE_PN1P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1197),
    .D(_00566_),
    .Q_N(\top_ihp.oisc.regs[12][26] ),
    .Q(_00259_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][27]$_DFFE_PN1P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1188),
    .D(_00567_),
    .Q_N(\top_ihp.oisc.regs[12][27] ),
    .Q(_00260_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][28]$_DFFE_PN1P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1201),
    .D(_00568_),
    .Q_N(\top_ihp.oisc.regs[12][28] ),
    .Q(_00261_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][29]$_DFFE_PN1P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1203),
    .D(_00569_),
    .Q_N(\top_ihp.oisc.regs[12][29] ),
    .Q(_00262_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][2]$_DFFE_PN1P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1235),
    .D(_00570_),
    .Q_N(\top_ihp.oisc.regs[12][2] ),
    .Q(_00263_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][30]$_DFFE_PN1P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1162),
    .D(_00571_),
    .Q_N(\top_ihp.oisc.regs[12][30] ),
    .Q(_00264_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][31]$_DFFE_PN1P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1160),
    .D(_00572_),
    .Q_N(\top_ihp.oisc.regs[12][31] ),
    .Q(_00265_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][3]$_DFFE_PN1P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1187),
    .D(_00573_),
    .Q_N(\top_ihp.oisc.regs[12][3] ),
    .Q(_00266_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][4]$_DFFE_PN1P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1160),
    .D(_00574_),
    .Q_N(\top_ihp.oisc.regs[12][4] ),
    .Q(_00267_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][5]$_DFFE_PN1P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1162),
    .D(_00575_),
    .Q_N(\top_ihp.oisc.regs[12][5] ),
    .Q(_00268_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][6]$_DFFE_PN1P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1235),
    .D(_00576_),
    .Q_N(\top_ihp.oisc.regs[12][6] ),
    .Q(_00269_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][7]$_DFFE_PN1P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1162),
    .D(_00577_),
    .Q_N(\top_ihp.oisc.regs[12][7] ),
    .Q(_00270_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][8]$_DFFE_PN1P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1232),
    .D(_00578_),
    .Q_N(\top_ihp.oisc.regs[12][8] ),
    .Q(_00271_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][9]$_DFFE_PN1P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1215),
    .D(_00579_),
    .Q_N(\top_ihp.oisc.regs[12][9] ),
    .Q(_00272_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1209),
    .D(_00580_),
    .Q_N(_13353_),
    .Q(\top_ihp.oisc.regs[13][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][10]$_DFFE_PN1P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1167),
    .D(_00581_),
    .Q_N(\top_ihp.oisc.regs[13][10] ),
    .Q(_00273_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][11]$_DFFE_PN1P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1175),
    .D(_00582_),
    .Q_N(\top_ihp.oisc.regs[13][11] ),
    .Q(_00274_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][12]$_DFFE_PN1P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1153),
    .D(_00583_),
    .Q_N(\top_ihp.oisc.regs[13][12] ),
    .Q(_00275_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][13]$_DFFE_PN1P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1153),
    .D(_00584_),
    .Q_N(\top_ihp.oisc.regs[13][13] ),
    .Q(_00276_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][14]$_DFFE_PN1P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1208),
    .D(_00585_),
    .Q_N(\top_ihp.oisc.regs[13][14] ),
    .Q(_00277_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][15]$_DFFE_PN1P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1208),
    .D(_00586_),
    .Q_N(\top_ihp.oisc.regs[13][15] ),
    .Q(_00278_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][16]$_DFFE_PN1P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1211),
    .D(_00587_),
    .Q_N(\top_ihp.oisc.regs[13][16] ),
    .Q(_00279_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][17]$_DFFE_PN1P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1156),
    .D(_00588_),
    .Q_N(\top_ihp.oisc.regs[13][17] ),
    .Q(_00280_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][18]$_DFFE_PN1P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1154),
    .D(_00589_),
    .Q_N(\top_ihp.oisc.regs[13][18] ),
    .Q(_00281_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][19]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1154),
    .D(_00590_),
    .Q_N(\top_ihp.oisc.regs[13][19] ),
    .Q(_00282_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1182),
    .D(_00591_),
    .Q_N(_13352_),
    .Q(\top_ihp.oisc.regs[13][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][20]$_DFFE_PN1P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1229),
    .D(_00592_),
    .Q_N(\top_ihp.oisc.regs[13][20] ),
    .Q(_00283_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][21]$_DFFE_PN1P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1155),
    .D(_00593_),
    .Q_N(\top_ihp.oisc.regs[13][21] ),
    .Q(_00284_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][22]$_DFFE_PN1P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1213),
    .D(_00594_),
    .Q_N(\top_ihp.oisc.regs[13][22] ),
    .Q(_00285_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][23]$_DFFE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1155),
    .D(_00595_),
    .Q_N(\top_ihp.oisc.regs[13][23] ),
    .Q(_00286_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][24]$_DFFE_PN1P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1232),
    .D(_00596_),
    .Q_N(\top_ihp.oisc.regs[13][24] ),
    .Q(_00287_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][25]$_DFFE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1155),
    .D(_00597_),
    .Q_N(\top_ihp.oisc.regs[13][25] ),
    .Q(_00288_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][26]$_DFFE_PN1P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1196),
    .D(_00598_),
    .Q_N(\top_ihp.oisc.regs[13][26] ),
    .Q(_00289_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][27]$_DFFE_PN1P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1186),
    .D(_00599_),
    .Q_N(\top_ihp.oisc.regs[13][27] ),
    .Q(_00290_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][28]$_DFFE_PN1P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1201),
    .D(_00600_),
    .Q_N(\top_ihp.oisc.regs[13][28] ),
    .Q(_00291_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][29]$_DFFE_PN1P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1204),
    .D(_00601_),
    .Q_N(\top_ihp.oisc.regs[13][29] ),
    .Q(_00292_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][2]$_DFFE_PN1P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1237),
    .D(_00602_),
    .Q_N(\top_ihp.oisc.regs[13][2] ),
    .Q(_00293_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][30]$_DFFE_PN1P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1191),
    .D(_00603_),
    .Q_N(\top_ihp.oisc.regs[13][30] ),
    .Q(_00294_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][31]$_DFFE_PN1P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1200),
    .D(_00604_),
    .Q_N(\top_ihp.oisc.regs[13][31] ),
    .Q(_00295_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][3]$_DFFE_PN1P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1187),
    .D(_00605_),
    .Q_N(\top_ihp.oisc.regs[13][3] ),
    .Q(_00296_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][4]$_DFFE_PN1P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1191),
    .D(_00606_),
    .Q_N(\top_ihp.oisc.regs[13][4] ),
    .Q(_00297_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][5]$_DFFE_PN1P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1191),
    .D(_00607_),
    .Q_N(\top_ihp.oisc.regs[13][5] ),
    .Q(_00298_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][6]$_DFFE_PN1P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1236),
    .D(_00608_),
    .Q_N(\top_ihp.oisc.regs[13][6] ),
    .Q(_00299_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][7]$_DFFE_PN1P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1234),
    .D(_00609_),
    .Q_N(\top_ihp.oisc.regs[13][7] ),
    .Q(_00300_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][8]$_DFFE_PN1P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1233),
    .D(_00610_),
    .Q_N(\top_ihp.oisc.regs[13][8] ),
    .Q(_00301_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][9]$_DFFE_PN1P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1215),
    .D(_00611_),
    .Q_N(\top_ihp.oisc.regs[13][9] ),
    .Q(_00302_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1212),
    .D(_00612_),
    .Q_N(_13351_),
    .Q(\top_ihp.oisc.regs[14][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1166),
    .D(_00613_),
    .Q_N(_13350_),
    .Q(\top_ihp.oisc.regs[14][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1211),
    .D(_00614_),
    .Q_N(_13349_),
    .Q(\top_ihp.oisc.regs[14][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1178),
    .D(_00615_),
    .Q_N(_13348_),
    .Q(\top_ihp.oisc.regs[14][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1165),
    .D(_00616_),
    .Q_N(_13347_),
    .Q(\top_ihp.oisc.regs[14][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1211),
    .D(_00617_),
    .Q_N(_13346_),
    .Q(\top_ihp.oisc.regs[14][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1177),
    .D(_00618_),
    .Q_N(_13345_),
    .Q(\top_ihp.oisc.regs[14][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1212),
    .D(_00619_),
    .Q_N(_13344_),
    .Q(\top_ihp.oisc.regs[14][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1166),
    .D(_00620_),
    .Q_N(_13343_),
    .Q(\top_ihp.oisc.regs[14][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1176),
    .D(_00621_),
    .Q_N(_13342_),
    .Q(\top_ihp.oisc.regs[14][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1170),
    .D(_00622_),
    .Q_N(_13341_),
    .Q(\top_ihp.oisc.regs[14][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1183),
    .D(_00623_),
    .Q_N(_13340_),
    .Q(\top_ihp.oisc.regs[14][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1198),
    .D(_00624_),
    .Q_N(_13339_),
    .Q(\top_ihp.oisc.regs[14][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1170),
    .D(_00625_),
    .Q_N(_13338_),
    .Q(\top_ihp.oisc.regs[14][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1214),
    .D(_00626_),
    .Q_N(_13337_),
    .Q(\top_ihp.oisc.regs[14][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1171),
    .D(_00627_),
    .Q_N(_13336_),
    .Q(\top_ihp.oisc.regs[14][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1231),
    .D(_00628_),
    .Q_N(_13335_),
    .Q(\top_ihp.oisc.regs[14][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1173),
    .D(_00629_),
    .Q_N(_13334_),
    .Q(\top_ihp.oisc.regs[14][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1197),
    .D(_00630_),
    .Q_N(_13333_),
    .Q(\top_ihp.oisc.regs[14][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1188),
    .D(_00631_),
    .Q_N(_13332_),
    .Q(\top_ihp.oisc.regs[14][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1187),
    .D(_00632_),
    .Q_N(_13331_),
    .Q(\top_ihp.oisc.regs[14][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1203),
    .D(_00633_),
    .Q_N(_13330_),
    .Q(\top_ihp.oisc.regs[14][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1234),
    .D(_00634_),
    .Q_N(_13329_),
    .Q(\top_ihp.oisc.regs[14][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1194),
    .D(_00635_),
    .Q_N(_13328_),
    .Q(\top_ihp.oisc.regs[14][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1160),
    .D(_00636_),
    .Q_N(_13327_),
    .Q(\top_ihp.oisc.regs[14][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1187),
    .D(_00637_),
    .Q_N(_13326_),
    .Q(\top_ihp.oisc.regs[14][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1187),
    .D(_00638_),
    .Q_N(_13325_),
    .Q(\top_ihp.oisc.regs[14][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1192),
    .D(_00639_),
    .Q_N(_13324_),
    .Q(\top_ihp.oisc.regs[14][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1230),
    .D(_00640_),
    .Q_N(_13323_),
    .Q(\top_ihp.oisc.regs[14][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1234),
    .D(_00641_),
    .Q_N(_13322_),
    .Q(\top_ihp.oisc.regs[14][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1233),
    .D(_00642_),
    .Q_N(_13321_),
    .Q(\top_ihp.oisc.regs[14][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1217),
    .D(_00643_),
    .Q_N(_13320_),
    .Q(\top_ihp.oisc.regs[14][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1216),
    .D(_00644_),
    .Q_N(_13319_),
    .Q(\top_ihp.oisc.regs[15][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1166),
    .D(_00645_),
    .Q_N(_13318_),
    .Q(\top_ihp.oisc.regs[15][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1175),
    .D(_00646_),
    .Q_N(_13317_),
    .Q(\top_ihp.oisc.regs[15][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1211),
    .D(_00647_),
    .Q_N(_13316_),
    .Q(\top_ihp.oisc.regs[15][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1165),
    .D(_00648_),
    .Q_N(_13315_),
    .Q(\top_ihp.oisc.regs[15][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1211),
    .D(_00649_),
    .Q_N(_13314_),
    .Q(\top_ihp.oisc.regs[15][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1177),
    .D(_00650_),
    .Q_N(_13313_),
    .Q(\top_ihp.oisc.regs[15][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1212),
    .D(_00651_),
    .Q_N(_13312_),
    .Q(\top_ihp.oisc.regs[15][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1182),
    .D(_00652_),
    .Q_N(_13311_),
    .Q(\top_ihp.oisc.regs[15][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1170),
    .D(_00653_),
    .Q_N(_13310_),
    .Q(\top_ihp.oisc.regs[15][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1171),
    .D(_00654_),
    .Q_N(_13309_),
    .Q(\top_ihp.oisc.regs[15][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1179),
    .D(_00655_),
    .Q_N(_13308_),
    .Q(\top_ihp.oisc.regs[15][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1229),
    .D(_00656_),
    .Q_N(_13307_),
    .Q(\top_ihp.oisc.regs[15][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1186),
    .D(_00657_),
    .Q_N(_13306_),
    .Q(\top_ihp.oisc.regs[15][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1216),
    .D(_00658_),
    .Q_N(_13305_),
    .Q(\top_ihp.oisc.regs[15][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1171),
    .D(_00659_),
    .Q_N(_13304_),
    .Q(\top_ihp.oisc.regs[15][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1232),
    .D(_00660_),
    .Q_N(_13303_),
    .Q(\top_ihp.oisc.regs[15][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1173),
    .D(_00661_),
    .Q_N(_13302_),
    .Q(\top_ihp.oisc.regs[15][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1198),
    .D(_00662_),
    .Q_N(_13301_),
    .Q(\top_ihp.oisc.regs[15][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1186),
    .D(_00663_),
    .Q_N(_13300_),
    .Q(\top_ihp.oisc.regs[15][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1201),
    .D(_00664_),
    .Q_N(_13299_),
    .Q(\top_ihp.oisc.regs[15][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1203),
    .D(_00665_),
    .Q_N(_13298_),
    .Q(\top_ihp.oisc.regs[15][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1237),
    .D(_00666_),
    .Q_N(_13297_),
    .Q(\top_ihp.oisc.regs[15][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1192),
    .D(_00667_),
    .Q_N(_13296_),
    .Q(\top_ihp.oisc.regs[15][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1193),
    .D(_00668_),
    .Q_N(_13295_),
    .Q(\top_ihp.oisc.regs[15][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1194),
    .D(_00669_),
    .Q_N(_13294_),
    .Q(\top_ihp.oisc.regs[15][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1191),
    .D(_00670_),
    .Q_N(_13293_),
    .Q(\top_ihp.oisc.regs[15][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1191),
    .D(_00671_),
    .Q_N(_13292_),
    .Q(\top_ihp.oisc.regs[15][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1236),
    .D(_00672_),
    .Q_N(_13291_),
    .Q(\top_ihp.oisc.regs[15][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1236),
    .D(_00673_),
    .Q_N(_13290_),
    .Q(\top_ihp.oisc.regs[15][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1231),
    .D(_00674_),
    .Q_N(_13289_),
    .Q(\top_ihp.oisc.regs[15][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1215),
    .D(_00675_),
    .Q_N(_13288_),
    .Q(\top_ihp.oisc.regs[15][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1449),
    .D(_00676_),
    .Q_N(_13287_),
    .Q(\top_ihp.oisc.regs[16][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1450),
    .D(_00677_),
    .Q_N(_13286_),
    .Q(\top_ihp.oisc.regs[16][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1451),
    .D(_00678_),
    .Q_N(_13285_),
    .Q(\top_ihp.oisc.regs[16][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][12]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1452),
    .D(_00679_),
    .Q_N(_13284_),
    .Q(\top_ihp.oisc.regs[16][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][13]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1453),
    .D(_00680_),
    .Q_N(_13283_),
    .Q(\top_ihp.oisc.regs[16][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][14]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1454),
    .D(_00681_),
    .Q_N(_13282_),
    .Q(\top_ihp.oisc.regs[16][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][15]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1455),
    .D(_00682_),
    .Q_N(_13281_),
    .Q(\top_ihp.oisc.regs[16][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][16]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1456),
    .D(_00683_),
    .Q_N(_13280_),
    .Q(\top_ihp.oisc.regs[16][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][17]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1457),
    .D(_00684_),
    .Q_N(_13279_),
    .Q(\top_ihp.oisc.regs[16][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][18]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1458),
    .D(_00685_),
    .Q_N(_13278_),
    .Q(\top_ihp.oisc.regs[16][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][19]$_DFFE_PP_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1459),
    .D(_00686_),
    .Q_N(_13277_),
    .Q(\top_ihp.oisc.regs[16][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1460),
    .D(_00687_),
    .Q_N(_13276_),
    .Q(\top_ihp.oisc.regs[16][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][20]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1461),
    .D(_00688_),
    .Q_N(_13275_),
    .Q(\top_ihp.oisc.regs[16][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][21]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1462),
    .D(_00689_),
    .Q_N(_13274_),
    .Q(\top_ihp.oisc.regs[16][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][22]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1463),
    .D(_00690_),
    .Q_N(_13273_),
    .Q(\top_ihp.oisc.regs[16][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][23]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1464),
    .D(_00691_),
    .Q_N(_13272_),
    .Q(\top_ihp.oisc.regs[16][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][24]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1465),
    .D(_00692_),
    .Q_N(_13271_),
    .Q(\top_ihp.oisc.regs[16][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][25]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1466),
    .D(_00693_),
    .Q_N(_13270_),
    .Q(\top_ihp.oisc.regs[16][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][26]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1467),
    .D(_00694_),
    .Q_N(_13269_),
    .Q(\top_ihp.oisc.regs[16][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][27]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1468),
    .D(_00695_),
    .Q_N(_13268_),
    .Q(\top_ihp.oisc.regs[16][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][28]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1469),
    .D(_00696_),
    .Q_N(_13267_),
    .Q(\top_ihp.oisc.regs[16][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][29]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1470),
    .D(_00697_),
    .Q_N(_13266_),
    .Q(\top_ihp.oisc.regs[16][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1471),
    .D(_00698_),
    .Q_N(_13265_),
    .Q(\top_ihp.oisc.regs[16][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][30]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1472),
    .D(_00699_),
    .Q_N(_13264_),
    .Q(\top_ihp.oisc.regs[16][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][31]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1473),
    .D(_00700_),
    .Q_N(_13263_),
    .Q(\top_ihp.oisc.regs[16][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1474),
    .D(_00701_),
    .Q_N(_13262_),
    .Q(\top_ihp.oisc.regs[16][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1475),
    .D(_00702_),
    .Q_N(_13261_),
    .Q(\top_ihp.oisc.regs[16][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1476),
    .D(_00703_),
    .Q_N(_13260_),
    .Q(\top_ihp.oisc.regs[16][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1477),
    .D(_00704_),
    .Q_N(_13259_),
    .Q(\top_ihp.oisc.regs[16][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1478),
    .D(_00705_),
    .Q_N(_13258_),
    .Q(\top_ihp.oisc.regs[16][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1479),
    .D(_00706_),
    .Q_N(_13257_),
    .Q(\top_ihp.oisc.regs[16][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1480),
    .D(_00707_),
    .Q_N(_13256_),
    .Q(\top_ihp.oisc.regs[16][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1481),
    .D(_00708_),
    .Q_N(_13255_),
    .Q(\top_ihp.oisc.regs[17][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1482),
    .D(_00709_),
    .Q_N(_13254_),
    .Q(\top_ihp.oisc.regs[17][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1483),
    .D(_00710_),
    .Q_N(_13253_),
    .Q(\top_ihp.oisc.regs[17][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][12]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1484),
    .D(_00711_),
    .Q_N(_13252_),
    .Q(\top_ihp.oisc.regs[17][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][13]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1485),
    .D(_00712_),
    .Q_N(_13251_),
    .Q(\top_ihp.oisc.regs[17][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][14]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1486),
    .D(_00713_),
    .Q_N(_13250_),
    .Q(\top_ihp.oisc.regs[17][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][15]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1487),
    .D(_00714_),
    .Q_N(_13249_),
    .Q(\top_ihp.oisc.regs[17][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][16]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1488),
    .D(_00715_),
    .Q_N(_13248_),
    .Q(\top_ihp.oisc.regs[17][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][17]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1489),
    .D(_00716_),
    .Q_N(_13247_),
    .Q(\top_ihp.oisc.regs[17][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][18]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1490),
    .D(_00717_),
    .Q_N(_13246_),
    .Q(\top_ihp.oisc.regs[17][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][19]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1491),
    .D(_00718_),
    .Q_N(_13245_),
    .Q(\top_ihp.oisc.regs[17][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1492),
    .D(_00719_),
    .Q_N(_13244_),
    .Q(\top_ihp.oisc.regs[17][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][20]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1493),
    .D(_00720_),
    .Q_N(_13243_),
    .Q(\top_ihp.oisc.regs[17][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][21]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1494),
    .D(_00721_),
    .Q_N(_13242_),
    .Q(\top_ihp.oisc.regs[17][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][22]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1495),
    .D(_00722_),
    .Q_N(_13241_),
    .Q(\top_ihp.oisc.regs[17][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][23]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1496),
    .D(_00723_),
    .Q_N(_13240_),
    .Q(\top_ihp.oisc.regs[17][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][24]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1497),
    .D(_00724_),
    .Q_N(_13239_),
    .Q(\top_ihp.oisc.regs[17][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][25]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1498),
    .D(_00725_),
    .Q_N(_13238_),
    .Q(\top_ihp.oisc.regs[17][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][26]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1499),
    .D(_00726_),
    .Q_N(_13237_),
    .Q(\top_ihp.oisc.regs[17][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][27]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1500),
    .D(_00727_),
    .Q_N(_13236_),
    .Q(\top_ihp.oisc.regs[17][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][28]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1501),
    .D(_00728_),
    .Q_N(_13235_),
    .Q(\top_ihp.oisc.regs[17][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][29]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1502),
    .D(_00729_),
    .Q_N(_13234_),
    .Q(\top_ihp.oisc.regs[17][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1503),
    .D(_00730_),
    .Q_N(_13233_),
    .Q(\top_ihp.oisc.regs[17][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][30]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1504),
    .D(_00731_),
    .Q_N(_13232_),
    .Q(\top_ihp.oisc.regs[17][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][31]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1505),
    .D(_00732_),
    .Q_N(_13231_),
    .Q(\top_ihp.oisc.regs[17][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1506),
    .D(_00733_),
    .Q_N(_13230_),
    .Q(\top_ihp.oisc.regs[17][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1507),
    .D(_00734_),
    .Q_N(_13229_),
    .Q(\top_ihp.oisc.regs[17][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1508),
    .D(_00735_),
    .Q_N(_13228_),
    .Q(\top_ihp.oisc.regs[17][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1509),
    .D(_00736_),
    .Q_N(_13227_),
    .Q(\top_ihp.oisc.regs[17][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1510),
    .D(_00737_),
    .Q_N(_13226_),
    .Q(\top_ihp.oisc.regs[17][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1511),
    .D(_00738_),
    .Q_N(_13225_),
    .Q(\top_ihp.oisc.regs[17][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1512),
    .D(_00739_),
    .Q_N(_13224_),
    .Q(\top_ihp.oisc.regs[17][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1513),
    .D(_00740_),
    .Q_N(_13223_),
    .Q(\top_ihp.oisc.regs[18][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1514),
    .D(_00741_),
    .Q_N(_13222_),
    .Q(\top_ihp.oisc.regs[18][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1515),
    .D(_00742_),
    .Q_N(_13221_),
    .Q(\top_ihp.oisc.regs[18][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][12]$_DFFE_PP_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1516),
    .D(_00743_),
    .Q_N(_13220_),
    .Q(\top_ihp.oisc.regs[18][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][13]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1517),
    .D(_00744_),
    .Q_N(_13219_),
    .Q(\top_ihp.oisc.regs[18][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][14]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1518),
    .D(_00745_),
    .Q_N(_13218_),
    .Q(\top_ihp.oisc.regs[18][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][15]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1519),
    .D(_00746_),
    .Q_N(_13217_),
    .Q(\top_ihp.oisc.regs[18][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][16]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1520),
    .D(_00747_),
    .Q_N(_13216_),
    .Q(\top_ihp.oisc.regs[18][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][17]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1521),
    .D(_00748_),
    .Q_N(_13215_),
    .Q(\top_ihp.oisc.regs[18][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][18]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1522),
    .D(_00749_),
    .Q_N(_13214_),
    .Q(\top_ihp.oisc.regs[18][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][19]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1523),
    .D(_00750_),
    .Q_N(_13213_),
    .Q(\top_ihp.oisc.regs[18][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1524),
    .D(_00751_),
    .Q_N(_13212_),
    .Q(\top_ihp.oisc.regs[18][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][20]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1525),
    .D(_00752_),
    .Q_N(_13211_),
    .Q(\top_ihp.oisc.regs[18][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][21]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1526),
    .D(_00753_),
    .Q_N(_13210_),
    .Q(\top_ihp.oisc.regs[18][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][22]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1527),
    .D(_00754_),
    .Q_N(_13209_),
    .Q(\top_ihp.oisc.regs[18][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][23]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1528),
    .D(_00755_),
    .Q_N(_13208_),
    .Q(\top_ihp.oisc.regs[18][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][24]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1529),
    .D(_00756_),
    .Q_N(_13207_),
    .Q(\top_ihp.oisc.regs[18][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][25]$_DFFE_PP_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1530),
    .D(_00757_),
    .Q_N(_13206_),
    .Q(\top_ihp.oisc.regs[18][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][26]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1531),
    .D(_00758_),
    .Q_N(_13205_),
    .Q(\top_ihp.oisc.regs[18][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][27]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1532),
    .D(_00759_),
    .Q_N(_13204_),
    .Q(\top_ihp.oisc.regs[18][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][28]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1533),
    .D(_00760_),
    .Q_N(_13203_),
    .Q(\top_ihp.oisc.regs[18][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][29]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1534),
    .D(_00761_),
    .Q_N(_13202_),
    .Q(\top_ihp.oisc.regs[18][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1535),
    .D(_00762_),
    .Q_N(_13201_),
    .Q(\top_ihp.oisc.regs[18][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][30]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1536),
    .D(_00763_),
    .Q_N(_13200_),
    .Q(\top_ihp.oisc.regs[18][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][31]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1537),
    .D(_00764_),
    .Q_N(_13199_),
    .Q(\top_ihp.oisc.regs[18][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1538),
    .D(_00765_),
    .Q_N(_13198_),
    .Q(\top_ihp.oisc.regs[18][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1539),
    .D(_00766_),
    .Q_N(_13197_),
    .Q(\top_ihp.oisc.regs[18][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1540),
    .D(_00767_),
    .Q_N(_13196_),
    .Q(\top_ihp.oisc.regs[18][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1541),
    .D(_00768_),
    .Q_N(_13195_),
    .Q(\top_ihp.oisc.regs[18][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1542),
    .D(_00769_),
    .Q_N(_13194_),
    .Q(\top_ihp.oisc.regs[18][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1543),
    .D(_00770_),
    .Q_N(_13193_),
    .Q(\top_ihp.oisc.regs[18][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1544),
    .D(_00771_),
    .Q_N(_13192_),
    .Q(\top_ihp.oisc.regs[18][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1545),
    .D(_00772_),
    .Q_N(_13191_),
    .Q(\top_ihp.oisc.regs[19][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1546),
    .D(_00773_),
    .Q_N(_13190_),
    .Q(\top_ihp.oisc.regs[19][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1547),
    .D(_00774_),
    .Q_N(_13189_),
    .Q(\top_ihp.oisc.regs[19][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][12]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1548),
    .D(_00775_),
    .Q_N(_13188_),
    .Q(\top_ihp.oisc.regs[19][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][13]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1549),
    .D(_00776_),
    .Q_N(_13187_),
    .Q(\top_ihp.oisc.regs[19][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][14]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1550),
    .D(_00777_),
    .Q_N(_13186_),
    .Q(\top_ihp.oisc.regs[19][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][15]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1551),
    .D(_00778_),
    .Q_N(_13185_),
    .Q(\top_ihp.oisc.regs[19][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][16]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1552),
    .D(_00779_),
    .Q_N(_13184_),
    .Q(\top_ihp.oisc.regs[19][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][17]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1553),
    .D(_00780_),
    .Q_N(_13183_),
    .Q(\top_ihp.oisc.regs[19][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][18]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1554),
    .D(_00781_),
    .Q_N(_13182_),
    .Q(\top_ihp.oisc.regs[19][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][19]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1555),
    .D(_00782_),
    .Q_N(_13181_),
    .Q(\top_ihp.oisc.regs[19][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1556),
    .D(_00783_),
    .Q_N(_13180_),
    .Q(\top_ihp.oisc.regs[19][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][20]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1557),
    .D(_00784_),
    .Q_N(_13179_),
    .Q(\top_ihp.oisc.regs[19][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][21]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1558),
    .D(_00785_),
    .Q_N(_13178_),
    .Q(\top_ihp.oisc.regs[19][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][22]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1559),
    .D(_00786_),
    .Q_N(_13177_),
    .Q(\top_ihp.oisc.regs[19][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][23]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1560),
    .D(_00787_),
    .Q_N(_13176_),
    .Q(\top_ihp.oisc.regs[19][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][24]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1561),
    .D(_00788_),
    .Q_N(_13175_),
    .Q(\top_ihp.oisc.regs[19][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][25]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1562),
    .D(_00789_),
    .Q_N(_13174_),
    .Q(\top_ihp.oisc.regs[19][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][26]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1563),
    .D(_00790_),
    .Q_N(_13173_),
    .Q(\top_ihp.oisc.regs[19][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][27]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1564),
    .D(_00791_),
    .Q_N(_13172_),
    .Q(\top_ihp.oisc.regs[19][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][28]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1565),
    .D(_00792_),
    .Q_N(_13171_),
    .Q(\top_ihp.oisc.regs[19][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][29]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1566),
    .D(_00793_),
    .Q_N(_13170_),
    .Q(\top_ihp.oisc.regs[19][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1567),
    .D(_00794_),
    .Q_N(_13169_),
    .Q(\top_ihp.oisc.regs[19][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][30]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1568),
    .D(_00795_),
    .Q_N(_13168_),
    .Q(\top_ihp.oisc.regs[19][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][31]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1569),
    .D(_00796_),
    .Q_N(_13167_),
    .Q(\top_ihp.oisc.regs[19][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1570),
    .D(_00797_),
    .Q_N(_13166_),
    .Q(\top_ihp.oisc.regs[19][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1571),
    .D(_00798_),
    .Q_N(_13165_),
    .Q(\top_ihp.oisc.regs[19][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1572),
    .D(_00799_),
    .Q_N(_13164_),
    .Q(\top_ihp.oisc.regs[19][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1573),
    .D(_00800_),
    .Q_N(_13163_),
    .Q(\top_ihp.oisc.regs[19][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1574),
    .D(_00801_),
    .Q_N(_13162_),
    .Q(\top_ihp.oisc.regs[19][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1575),
    .D(_00802_),
    .Q_N(_13161_),
    .Q(\top_ihp.oisc.regs[19][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1576),
    .D(_00803_),
    .Q_N(_13160_),
    .Q(\top_ihp.oisc.regs[19][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1212),
    .D(_00804_),
    .Q_N(_13159_),
    .Q(\top_ihp.oisc.regs[1][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1169),
    .D(_00805_),
    .Q_N(_13158_),
    .Q(\top_ihp.oisc.regs[1][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1168),
    .D(_00806_),
    .Q_N(_13157_),
    .Q(\top_ihp.oisc.regs[1][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1176),
    .D(_00807_),
    .Q_N(_13156_),
    .Q(\top_ihp.oisc.regs[1][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1168),
    .D(_00808_),
    .Q_N(_13155_),
    .Q(\top_ihp.oisc.regs[1][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1208),
    .D(_00809_),
    .Q_N(_13154_),
    .Q(\top_ihp.oisc.regs[1][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1177),
    .D(_00810_),
    .Q_N(_13153_),
    .Q(\top_ihp.oisc.regs[1][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1209),
    .D(_00811_),
    .Q_N(_13152_),
    .Q(\top_ihp.oisc.regs[1][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1169),
    .D(_00812_),
    .Q_N(_13151_),
    .Q(\top_ihp.oisc.regs[1][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1179),
    .D(_00813_),
    .Q_N(_13150_),
    .Q(\top_ihp.oisc.regs[1][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1172),
    .D(_00814_),
    .Q_N(_13149_),
    .Q(\top_ihp.oisc.regs[1][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1182),
    .D(_00815_),
    .Q_N(_13148_),
    .Q(\top_ihp.oisc.regs[1][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1198),
    .D(_00816_),
    .Q_N(_13147_),
    .Q(\top_ihp.oisc.regs[1][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1188),
    .D(_00817_),
    .Q_N(_13146_),
    .Q(\top_ihp.oisc.regs[1][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1215),
    .D(_00818_),
    .Q_N(_13145_),
    .Q(\top_ihp.oisc.regs[1][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1181),
    .D(_00819_),
    .Q_N(_13144_),
    .Q(\top_ihp.oisc.regs[1][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1232),
    .D(_00820_),
    .Q_N(_13143_),
    .Q(\top_ihp.oisc.regs[1][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1172),
    .D(_00821_),
    .Q_N(_13142_),
    .Q(\top_ihp.oisc.regs[1][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1196),
    .D(_00822_),
    .Q_N(_13141_),
    .Q(\top_ihp.oisc.regs[1][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1196),
    .D(_00823_),
    .Q_N(_13140_),
    .Q(\top_ihp.oisc.regs[1][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1236),
    .D(_00824_),
    .Q_N(_13139_),
    .Q(\top_ihp.oisc.regs[1][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1234),
    .D(_00825_),
    .Q_N(_13138_),
    .Q(\top_ihp.oisc.regs[1][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1243),
    .D(_00826_),
    .Q_N(_13137_),
    .Q(\top_ihp.oisc.regs[1][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][30]$_DFFE_PN1P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1188),
    .D(_00827_),
    .Q_N(\top_ihp.oisc.regs[1][30] ),
    .Q(_00303_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1200),
    .D(_00828_),
    .Q_N(_13136_),
    .Q(\top_ihp.oisc.regs[1][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1196),
    .D(_00829_),
    .Q_N(_13135_),
    .Q(\top_ihp.oisc.regs[1][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1200),
    .D(_00830_),
    .Q_N(_13134_),
    .Q(\top_ihp.oisc.regs[1][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1200),
    .D(_00831_),
    .Q_N(_13133_),
    .Q(\top_ihp.oisc.regs[1][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1236),
    .D(_00832_),
    .Q_N(_13132_),
    .Q(\top_ihp.oisc.regs[1][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1236),
    .D(_00833_),
    .Q_N(_13131_),
    .Q(\top_ihp.oisc.regs[1][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1239),
    .D(_00834_),
    .Q_N(_13130_),
    .Q(\top_ihp.oisc.regs[1][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1215),
    .D(_00835_),
    .Q_N(_13129_),
    .Q(\top_ihp.oisc.regs[1][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1577),
    .D(_00836_),
    .Q_N(_13128_),
    .Q(\top_ihp.oisc.regs[20][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1578),
    .D(_00837_),
    .Q_N(_13127_),
    .Q(\top_ihp.oisc.regs[20][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1579),
    .D(_00838_),
    .Q_N(_13126_),
    .Q(\top_ihp.oisc.regs[20][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][12]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1580),
    .D(_00839_),
    .Q_N(_13125_),
    .Q(\top_ihp.oisc.regs[20][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][13]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1581),
    .D(_00840_),
    .Q_N(_13124_),
    .Q(\top_ihp.oisc.regs[20][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][14]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1582),
    .D(_00841_),
    .Q_N(_13123_),
    .Q(\top_ihp.oisc.regs[20][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][15]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1583),
    .D(_00842_),
    .Q_N(_13122_),
    .Q(\top_ihp.oisc.regs[20][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][16]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1584),
    .D(_00843_),
    .Q_N(_13121_),
    .Q(\top_ihp.oisc.regs[20][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][17]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1585),
    .D(_00844_),
    .Q_N(_13120_),
    .Q(\top_ihp.oisc.regs[20][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][18]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1586),
    .D(_00845_),
    .Q_N(_13119_),
    .Q(\top_ihp.oisc.regs[20][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][19]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1587),
    .D(_00846_),
    .Q_N(_13118_),
    .Q(\top_ihp.oisc.regs[20][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1588),
    .D(_00847_),
    .Q_N(_13117_),
    .Q(\top_ihp.oisc.regs[20][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][20]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1589),
    .D(_00848_),
    .Q_N(_13116_),
    .Q(\top_ihp.oisc.regs[20][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][21]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1590),
    .D(_00849_),
    .Q_N(_13115_),
    .Q(\top_ihp.oisc.regs[20][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][22]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1591),
    .D(_00850_),
    .Q_N(_13114_),
    .Q(\top_ihp.oisc.regs[20][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][23]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1592),
    .D(_00851_),
    .Q_N(_13113_),
    .Q(\top_ihp.oisc.regs[20][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][24]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1593),
    .D(_00852_),
    .Q_N(_13112_),
    .Q(\top_ihp.oisc.regs[20][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][25]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1594),
    .D(_00853_),
    .Q_N(_13111_),
    .Q(\top_ihp.oisc.regs[20][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][26]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1595),
    .D(_00854_),
    .Q_N(_13110_),
    .Q(\top_ihp.oisc.regs[20][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][27]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1596),
    .D(_00855_),
    .Q_N(_13109_),
    .Q(\top_ihp.oisc.regs[20][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][28]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1597),
    .D(_00856_),
    .Q_N(_13108_),
    .Q(\top_ihp.oisc.regs[20][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][29]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1598),
    .D(_00857_),
    .Q_N(_13107_),
    .Q(\top_ihp.oisc.regs[20][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1599),
    .D(_00858_),
    .Q_N(_13106_),
    .Q(\top_ihp.oisc.regs[20][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][30]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1600),
    .D(_00859_),
    .Q_N(_13105_),
    .Q(\top_ihp.oisc.regs[20][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][31]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1601),
    .D(_00860_),
    .Q_N(_13104_),
    .Q(\top_ihp.oisc.regs[20][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1602),
    .D(_00861_),
    .Q_N(_13103_),
    .Q(\top_ihp.oisc.regs[20][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1603),
    .D(_00862_),
    .Q_N(_13102_),
    .Q(\top_ihp.oisc.regs[20][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1604),
    .D(_00863_),
    .Q_N(_13101_),
    .Q(\top_ihp.oisc.regs[20][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1605),
    .D(_00864_),
    .Q_N(_13100_),
    .Q(\top_ihp.oisc.regs[20][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1606),
    .D(_00865_),
    .Q_N(_13099_),
    .Q(\top_ihp.oisc.regs[20][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1607),
    .D(_00866_),
    .Q_N(_13098_),
    .Q(\top_ihp.oisc.regs[20][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1608),
    .D(_00867_),
    .Q_N(_13097_),
    .Q(\top_ihp.oisc.regs[20][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1609),
    .D(_00868_),
    .Q_N(_13096_),
    .Q(\top_ihp.oisc.regs[21][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1610),
    .D(_00869_),
    .Q_N(_13095_),
    .Q(\top_ihp.oisc.regs[21][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1611),
    .D(_00870_),
    .Q_N(_13094_),
    .Q(\top_ihp.oisc.regs[21][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][12]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1612),
    .D(_00871_),
    .Q_N(_13093_),
    .Q(\top_ihp.oisc.regs[21][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][13]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1613),
    .D(_00872_),
    .Q_N(_13092_),
    .Q(\top_ihp.oisc.regs[21][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][14]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1614),
    .D(_00873_),
    .Q_N(_13091_),
    .Q(\top_ihp.oisc.regs[21][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][15]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1615),
    .D(_00874_),
    .Q_N(_13090_),
    .Q(\top_ihp.oisc.regs[21][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][16]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1616),
    .D(_00875_),
    .Q_N(_13089_),
    .Q(\top_ihp.oisc.regs[21][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][17]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1617),
    .D(_00876_),
    .Q_N(_13088_),
    .Q(\top_ihp.oisc.regs[21][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][18]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1618),
    .D(_00877_),
    .Q_N(_13087_),
    .Q(\top_ihp.oisc.regs[21][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][19]$_DFFE_PP_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1619),
    .D(_00878_),
    .Q_N(_13086_),
    .Q(\top_ihp.oisc.regs[21][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1620),
    .D(_00879_),
    .Q_N(_13085_),
    .Q(\top_ihp.oisc.regs[21][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][20]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1621),
    .D(_00880_),
    .Q_N(_13084_),
    .Q(\top_ihp.oisc.regs[21][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][21]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1622),
    .D(_00881_),
    .Q_N(_13083_),
    .Q(\top_ihp.oisc.regs[21][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][22]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1623),
    .D(_00882_),
    .Q_N(_13082_),
    .Q(\top_ihp.oisc.regs[21][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][23]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1624),
    .D(_00883_),
    .Q_N(_13081_),
    .Q(\top_ihp.oisc.regs[21][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][24]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1625),
    .D(_00884_),
    .Q_N(_13080_),
    .Q(\top_ihp.oisc.regs[21][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][25]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1626),
    .D(_00885_),
    .Q_N(_13079_),
    .Q(\top_ihp.oisc.regs[21][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][26]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1627),
    .D(_00886_),
    .Q_N(_13078_),
    .Q(\top_ihp.oisc.regs[21][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][27]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1628),
    .D(_00887_),
    .Q_N(_13077_),
    .Q(\top_ihp.oisc.regs[21][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][28]$_DFFE_PP_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1629),
    .D(_00888_),
    .Q_N(_13076_),
    .Q(\top_ihp.oisc.regs[21][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][29]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1630),
    .D(_00889_),
    .Q_N(_13075_),
    .Q(\top_ihp.oisc.regs[21][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1631),
    .D(_00890_),
    .Q_N(_13074_),
    .Q(\top_ihp.oisc.regs[21][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][30]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1632),
    .D(_00891_),
    .Q_N(_13073_),
    .Q(\top_ihp.oisc.regs[21][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][31]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1633),
    .D(_00892_),
    .Q_N(_13072_),
    .Q(\top_ihp.oisc.regs[21][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1634),
    .D(_00893_),
    .Q_N(_13071_),
    .Q(\top_ihp.oisc.regs[21][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1635),
    .D(_00894_),
    .Q_N(_13070_),
    .Q(\top_ihp.oisc.regs[21][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1636),
    .D(_00895_),
    .Q_N(_13069_),
    .Q(\top_ihp.oisc.regs[21][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1637),
    .D(_00896_),
    .Q_N(_13068_),
    .Q(\top_ihp.oisc.regs[21][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1638),
    .D(_00897_),
    .Q_N(_13067_),
    .Q(\top_ihp.oisc.regs[21][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1639),
    .D(_00898_),
    .Q_N(_13066_),
    .Q(\top_ihp.oisc.regs[21][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1640),
    .D(_00899_),
    .Q_N(_13065_),
    .Q(\top_ihp.oisc.regs[21][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1641),
    .D(_00900_),
    .Q_N(_13064_),
    .Q(\top_ihp.oisc.regs[22][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1642),
    .D(_00901_),
    .Q_N(_13063_),
    .Q(\top_ihp.oisc.regs[22][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1643),
    .D(_00902_),
    .Q_N(_13062_),
    .Q(\top_ihp.oisc.regs[22][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][12]$_DFFE_PP_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1644),
    .D(_00903_),
    .Q_N(_13061_),
    .Q(\top_ihp.oisc.regs[22][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][13]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1645),
    .D(_00904_),
    .Q_N(_13060_),
    .Q(\top_ihp.oisc.regs[22][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][14]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1646),
    .D(_00905_),
    .Q_N(_13059_),
    .Q(\top_ihp.oisc.regs[22][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][15]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1647),
    .D(_00906_),
    .Q_N(_13058_),
    .Q(\top_ihp.oisc.regs[22][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][16]$_DFFE_PP_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1648),
    .D(_00907_),
    .Q_N(_13057_),
    .Q(\top_ihp.oisc.regs[22][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][17]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1649),
    .D(_00908_),
    .Q_N(_13056_),
    .Q(\top_ihp.oisc.regs[22][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][18]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1650),
    .D(_00909_),
    .Q_N(_13055_),
    .Q(\top_ihp.oisc.regs[22][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][19]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1651),
    .D(_00910_),
    .Q_N(_13054_),
    .Q(\top_ihp.oisc.regs[22][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1652),
    .D(_00911_),
    .Q_N(_13053_),
    .Q(\top_ihp.oisc.regs[22][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][20]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1653),
    .D(_00912_),
    .Q_N(_13052_),
    .Q(\top_ihp.oisc.regs[22][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][21]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1654),
    .D(_00913_),
    .Q_N(_13051_),
    .Q(\top_ihp.oisc.regs[22][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][22]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1655),
    .D(_00914_),
    .Q_N(_13050_),
    .Q(\top_ihp.oisc.regs[22][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][23]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1656),
    .D(_00915_),
    .Q_N(_13049_),
    .Q(\top_ihp.oisc.regs[22][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][24]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1657),
    .D(_00916_),
    .Q_N(_13048_),
    .Q(\top_ihp.oisc.regs[22][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][25]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1658),
    .D(_00917_),
    .Q_N(_13047_),
    .Q(\top_ihp.oisc.regs[22][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][26]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1659),
    .D(_00918_),
    .Q_N(_13046_),
    .Q(\top_ihp.oisc.regs[22][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][27]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1660),
    .D(_00919_),
    .Q_N(_13045_),
    .Q(\top_ihp.oisc.regs[22][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][28]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1661),
    .D(_00920_),
    .Q_N(_13044_),
    .Q(\top_ihp.oisc.regs[22][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][29]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1662),
    .D(_00921_),
    .Q_N(_13043_),
    .Q(\top_ihp.oisc.regs[22][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1663),
    .D(_00922_),
    .Q_N(_13042_),
    .Q(\top_ihp.oisc.regs[22][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][30]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1664),
    .D(_00923_),
    .Q_N(_13041_),
    .Q(\top_ihp.oisc.regs[22][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][31]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1665),
    .D(_00924_),
    .Q_N(_13040_),
    .Q(\top_ihp.oisc.regs[22][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1666),
    .D(_00925_),
    .Q_N(_13039_),
    .Q(\top_ihp.oisc.regs[22][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1667),
    .D(_00926_),
    .Q_N(_13038_),
    .Q(\top_ihp.oisc.regs[22][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1668),
    .D(_00927_),
    .Q_N(_13037_),
    .Q(\top_ihp.oisc.regs[22][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1669),
    .D(_00928_),
    .Q_N(_13036_),
    .Q(\top_ihp.oisc.regs[22][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1670),
    .D(_00929_),
    .Q_N(_13035_),
    .Q(\top_ihp.oisc.regs[22][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1671),
    .D(_00930_),
    .Q_N(_13034_),
    .Q(\top_ihp.oisc.regs[22][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1672),
    .D(_00931_),
    .Q_N(_13033_),
    .Q(\top_ihp.oisc.regs[22][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1673),
    .D(_00932_),
    .Q_N(_13032_),
    .Q(\top_ihp.oisc.regs[23][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1674),
    .D(_00933_),
    .Q_N(_13031_),
    .Q(\top_ihp.oisc.regs[23][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1675),
    .D(_00934_),
    .Q_N(_13030_),
    .Q(\top_ihp.oisc.regs[23][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][12]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1676),
    .D(_00935_),
    .Q_N(_13029_),
    .Q(\top_ihp.oisc.regs[23][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][13]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1677),
    .D(_00936_),
    .Q_N(_13028_),
    .Q(\top_ihp.oisc.regs[23][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][14]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1678),
    .D(_00937_),
    .Q_N(_13027_),
    .Q(\top_ihp.oisc.regs[23][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][15]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1679),
    .D(_00938_),
    .Q_N(_13026_),
    .Q(\top_ihp.oisc.regs[23][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][16]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1680),
    .D(_00939_),
    .Q_N(_13025_),
    .Q(\top_ihp.oisc.regs[23][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][17]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1681),
    .D(_00940_),
    .Q_N(_13024_),
    .Q(\top_ihp.oisc.regs[23][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][18]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1682),
    .D(_00941_),
    .Q_N(_13023_),
    .Q(\top_ihp.oisc.regs[23][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][19]$_DFFE_PP_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1683),
    .D(_00942_),
    .Q_N(_13022_),
    .Q(\top_ihp.oisc.regs[23][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1684),
    .D(_00943_),
    .Q_N(_13021_),
    .Q(\top_ihp.oisc.regs[23][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][20]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1685),
    .D(_00944_),
    .Q_N(_13020_),
    .Q(\top_ihp.oisc.regs[23][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][21]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1686),
    .D(_00945_),
    .Q_N(_13019_),
    .Q(\top_ihp.oisc.regs[23][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][22]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1687),
    .D(_00946_),
    .Q_N(_13018_),
    .Q(\top_ihp.oisc.regs[23][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][23]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1688),
    .D(_00947_),
    .Q_N(_13017_),
    .Q(\top_ihp.oisc.regs[23][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][24]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1689),
    .D(_00948_),
    .Q_N(_13016_),
    .Q(\top_ihp.oisc.regs[23][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][25]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1690),
    .D(_00949_),
    .Q_N(_13015_),
    .Q(\top_ihp.oisc.regs[23][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][26]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1691),
    .D(_00950_),
    .Q_N(_13014_),
    .Q(\top_ihp.oisc.regs[23][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][27]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1692),
    .D(_00951_),
    .Q_N(_13013_),
    .Q(\top_ihp.oisc.regs[23][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][28]$_DFFE_PP_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1693),
    .D(_00952_),
    .Q_N(_13012_),
    .Q(\top_ihp.oisc.regs[23][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][29]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1694),
    .D(_00953_),
    .Q_N(_13011_),
    .Q(\top_ihp.oisc.regs[23][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1695),
    .D(_00954_),
    .Q_N(_13010_),
    .Q(\top_ihp.oisc.regs[23][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][30]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1696),
    .D(_00955_),
    .Q_N(_13009_),
    .Q(\top_ihp.oisc.regs[23][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][31]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1697),
    .D(_00956_),
    .Q_N(_13008_),
    .Q(\top_ihp.oisc.regs[23][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1698),
    .D(_00957_),
    .Q_N(_13007_),
    .Q(\top_ihp.oisc.regs[23][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1699),
    .D(_00958_),
    .Q_N(_13006_),
    .Q(\top_ihp.oisc.regs[23][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1700),
    .D(_00959_),
    .Q_N(_13005_),
    .Q(\top_ihp.oisc.regs[23][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1701),
    .D(_00960_),
    .Q_N(_13004_),
    .Q(\top_ihp.oisc.regs[23][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1702),
    .D(_00961_),
    .Q_N(_13003_),
    .Q(\top_ihp.oisc.regs[23][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1703),
    .D(_00962_),
    .Q_N(_13002_),
    .Q(\top_ihp.oisc.regs[23][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1704),
    .D(_00963_),
    .Q_N(_13001_),
    .Q(\top_ihp.oisc.regs[23][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1705),
    .D(_00964_),
    .Q_N(_13000_),
    .Q(\top_ihp.oisc.regs[24][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1706),
    .D(_00965_),
    .Q_N(_12999_),
    .Q(\top_ihp.oisc.regs[24][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1707),
    .D(_00966_),
    .Q_N(_12998_),
    .Q(\top_ihp.oisc.regs[24][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][12]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1708),
    .D(_00967_),
    .Q_N(_12997_),
    .Q(\top_ihp.oisc.regs[24][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][13]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1709),
    .D(_00968_),
    .Q_N(_12996_),
    .Q(\top_ihp.oisc.regs[24][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][14]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1710),
    .D(_00969_),
    .Q_N(_12995_),
    .Q(\top_ihp.oisc.regs[24][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][15]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1711),
    .D(_00970_),
    .Q_N(_12994_),
    .Q(\top_ihp.oisc.regs[24][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][16]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1712),
    .D(_00971_),
    .Q_N(_12993_),
    .Q(\top_ihp.oisc.regs[24][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][17]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1713),
    .D(_00972_),
    .Q_N(_12992_),
    .Q(\top_ihp.oisc.regs[24][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][18]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1714),
    .D(_00973_),
    .Q_N(_12991_),
    .Q(\top_ihp.oisc.regs[24][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][19]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1715),
    .D(_00974_),
    .Q_N(_12990_),
    .Q(\top_ihp.oisc.regs[24][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1716),
    .D(_00975_),
    .Q_N(_12989_),
    .Q(\top_ihp.oisc.regs[24][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][20]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1717),
    .D(_00976_),
    .Q_N(_12988_),
    .Q(\top_ihp.oisc.regs[24][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][21]$_DFFE_PP_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1718),
    .D(_00977_),
    .Q_N(_12987_),
    .Q(\top_ihp.oisc.regs[24][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][22]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1719),
    .D(_00978_),
    .Q_N(_12986_),
    .Q(\top_ihp.oisc.regs[24][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][23]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1720),
    .D(_00979_),
    .Q_N(_12985_),
    .Q(\top_ihp.oisc.regs[24][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][24]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1721),
    .D(_00980_),
    .Q_N(_12984_),
    .Q(\top_ihp.oisc.regs[24][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][25]$_DFFE_PP_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1722),
    .D(_00981_),
    .Q_N(_12983_),
    .Q(\top_ihp.oisc.regs[24][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][26]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1723),
    .D(_00982_),
    .Q_N(_12982_),
    .Q(\top_ihp.oisc.regs[24][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][27]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1724),
    .D(_00983_),
    .Q_N(_12981_),
    .Q(\top_ihp.oisc.regs[24][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][28]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1725),
    .D(_00984_),
    .Q_N(_12980_),
    .Q(\top_ihp.oisc.regs[24][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][29]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1726),
    .D(_00985_),
    .Q_N(_12979_),
    .Q(\top_ihp.oisc.regs[24][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1727),
    .D(_00986_),
    .Q_N(_12978_),
    .Q(\top_ihp.oisc.regs[24][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][30]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1728),
    .D(_00987_),
    .Q_N(_12977_),
    .Q(\top_ihp.oisc.regs[24][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][31]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1729),
    .D(_00988_),
    .Q_N(_12976_),
    .Q(\top_ihp.oisc.regs[24][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1730),
    .D(_00989_),
    .Q_N(_12975_),
    .Q(\top_ihp.oisc.regs[24][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1731),
    .D(_00990_),
    .Q_N(_12974_),
    .Q(\top_ihp.oisc.regs[24][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1732),
    .D(_00991_),
    .Q_N(_12973_),
    .Q(\top_ihp.oisc.regs[24][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1733),
    .D(_00992_),
    .Q_N(_12972_),
    .Q(\top_ihp.oisc.regs[24][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1734),
    .D(_00993_),
    .Q_N(_12971_),
    .Q(\top_ihp.oisc.regs[24][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1735),
    .D(_00994_),
    .Q_N(_12970_),
    .Q(\top_ihp.oisc.regs[24][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1736),
    .D(_00995_),
    .Q_N(_12969_),
    .Q(\top_ihp.oisc.regs[24][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1737),
    .D(_00996_),
    .Q_N(_12968_),
    .Q(\top_ihp.oisc.regs[25][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1738),
    .D(_00997_),
    .Q_N(_12967_),
    .Q(\top_ihp.oisc.regs[25][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1739),
    .D(_00998_),
    .Q_N(_12966_),
    .Q(\top_ihp.oisc.regs[25][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][12]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1740),
    .D(_00999_),
    .Q_N(_12965_),
    .Q(\top_ihp.oisc.regs[25][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][13]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1741),
    .D(_01000_),
    .Q_N(_12964_),
    .Q(\top_ihp.oisc.regs[25][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][14]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1742),
    .D(_01001_),
    .Q_N(_12963_),
    .Q(\top_ihp.oisc.regs[25][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][15]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1743),
    .D(_01002_),
    .Q_N(_12962_),
    .Q(\top_ihp.oisc.regs[25][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][16]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1744),
    .D(_01003_),
    .Q_N(_12961_),
    .Q(\top_ihp.oisc.regs[25][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][17]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1745),
    .D(_01004_),
    .Q_N(_12960_),
    .Q(\top_ihp.oisc.regs[25][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][18]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1746),
    .D(_01005_),
    .Q_N(_12959_),
    .Q(\top_ihp.oisc.regs[25][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][19]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1747),
    .D(_01006_),
    .Q_N(_12958_),
    .Q(\top_ihp.oisc.regs[25][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1748),
    .D(_01007_),
    .Q_N(_12957_),
    .Q(\top_ihp.oisc.regs[25][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][20]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1749),
    .D(_01008_),
    .Q_N(_12956_),
    .Q(\top_ihp.oisc.regs[25][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][21]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1750),
    .D(_01009_),
    .Q_N(_12955_),
    .Q(\top_ihp.oisc.regs[25][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][22]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1751),
    .D(_01010_),
    .Q_N(_12954_),
    .Q(\top_ihp.oisc.regs[25][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][23]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1752),
    .D(_01011_),
    .Q_N(_12953_),
    .Q(\top_ihp.oisc.regs[25][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][24]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1753),
    .D(_01012_),
    .Q_N(_12952_),
    .Q(\top_ihp.oisc.regs[25][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][25]$_DFFE_PP_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1754),
    .D(_01013_),
    .Q_N(_12951_),
    .Q(\top_ihp.oisc.regs[25][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][26]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1755),
    .D(_01014_),
    .Q_N(_12950_),
    .Q(\top_ihp.oisc.regs[25][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][27]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1756),
    .D(_01015_),
    .Q_N(_12949_),
    .Q(\top_ihp.oisc.regs[25][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][28]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1757),
    .D(_01016_),
    .Q_N(_12948_),
    .Q(\top_ihp.oisc.regs[25][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][29]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1758),
    .D(_01017_),
    .Q_N(_12947_),
    .Q(\top_ihp.oisc.regs[25][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1759),
    .D(_01018_),
    .Q_N(_12946_),
    .Q(\top_ihp.oisc.regs[25][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][30]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1760),
    .D(_01019_),
    .Q_N(_12945_),
    .Q(\top_ihp.oisc.regs[25][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][31]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1761),
    .D(_01020_),
    .Q_N(_12944_),
    .Q(\top_ihp.oisc.regs[25][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1762),
    .D(_01021_),
    .Q_N(_12943_),
    .Q(\top_ihp.oisc.regs[25][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1763),
    .D(_01022_),
    .Q_N(_12942_),
    .Q(\top_ihp.oisc.regs[25][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1764),
    .D(_01023_),
    .Q_N(_12941_),
    .Q(\top_ihp.oisc.regs[25][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1765),
    .D(_01024_),
    .Q_N(_12940_),
    .Q(\top_ihp.oisc.regs[25][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1766),
    .D(_01025_),
    .Q_N(_12939_),
    .Q(\top_ihp.oisc.regs[25][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1767),
    .D(_01026_),
    .Q_N(_12938_),
    .Q(\top_ihp.oisc.regs[25][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1768),
    .D(_01027_),
    .Q_N(_12937_),
    .Q(\top_ihp.oisc.regs[25][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1769),
    .D(_01028_),
    .Q_N(_12936_),
    .Q(\top_ihp.oisc.regs[26][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1770),
    .D(_01029_),
    .Q_N(_12935_),
    .Q(\top_ihp.oisc.regs[26][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1771),
    .D(_01030_),
    .Q_N(_12934_),
    .Q(\top_ihp.oisc.regs[26][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][12]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1772),
    .D(_01031_),
    .Q_N(_12933_),
    .Q(\top_ihp.oisc.regs[26][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][13]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1773),
    .D(_01032_),
    .Q_N(_12932_),
    .Q(\top_ihp.oisc.regs[26][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][14]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1774),
    .D(_01033_),
    .Q_N(_12931_),
    .Q(\top_ihp.oisc.regs[26][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][15]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1775),
    .D(_01034_),
    .Q_N(_12930_),
    .Q(\top_ihp.oisc.regs[26][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][16]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1776),
    .D(_01035_),
    .Q_N(_12929_),
    .Q(\top_ihp.oisc.regs[26][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][17]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1777),
    .D(_01036_),
    .Q_N(_12928_),
    .Q(\top_ihp.oisc.regs[26][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][18]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1778),
    .D(_01037_),
    .Q_N(_12927_),
    .Q(\top_ihp.oisc.regs[26][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][19]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1779),
    .D(_01038_),
    .Q_N(_12926_),
    .Q(\top_ihp.oisc.regs[26][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1780),
    .D(_01039_),
    .Q_N(_12925_),
    .Q(\top_ihp.oisc.regs[26][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][20]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1781),
    .D(_01040_),
    .Q_N(_12924_),
    .Q(\top_ihp.oisc.regs[26][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][21]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1782),
    .D(_01041_),
    .Q_N(_12923_),
    .Q(\top_ihp.oisc.regs[26][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][22]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1783),
    .D(_01042_),
    .Q_N(_12922_),
    .Q(\top_ihp.oisc.regs[26][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][23]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1784),
    .D(_01043_),
    .Q_N(_12921_),
    .Q(\top_ihp.oisc.regs[26][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][24]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1785),
    .D(_01044_),
    .Q_N(_12920_),
    .Q(\top_ihp.oisc.regs[26][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][25]$_DFFE_PP_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1786),
    .D(_01045_),
    .Q_N(_12919_),
    .Q(\top_ihp.oisc.regs[26][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][26]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1787),
    .D(_01046_),
    .Q_N(_12918_),
    .Q(\top_ihp.oisc.regs[26][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][27]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1788),
    .D(_01047_),
    .Q_N(_12917_),
    .Q(\top_ihp.oisc.regs[26][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][28]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1789),
    .D(_01048_),
    .Q_N(_12916_),
    .Q(\top_ihp.oisc.regs[26][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][29]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1790),
    .D(_01049_),
    .Q_N(_12915_),
    .Q(\top_ihp.oisc.regs[26][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1791),
    .D(_01050_),
    .Q_N(_12914_),
    .Q(\top_ihp.oisc.regs[26][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][30]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1792),
    .D(_01051_),
    .Q_N(_12913_),
    .Q(\top_ihp.oisc.regs[26][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][31]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1793),
    .D(_01052_),
    .Q_N(_12912_),
    .Q(\top_ihp.oisc.regs[26][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1794),
    .D(_01053_),
    .Q_N(_12911_),
    .Q(\top_ihp.oisc.regs[26][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1795),
    .D(_01054_),
    .Q_N(_12910_),
    .Q(\top_ihp.oisc.regs[26][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1796),
    .D(_01055_),
    .Q_N(_12909_),
    .Q(\top_ihp.oisc.regs[26][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1797),
    .D(_01056_),
    .Q_N(_12908_),
    .Q(\top_ihp.oisc.regs[26][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1798),
    .D(_01057_),
    .Q_N(_12907_),
    .Q(\top_ihp.oisc.regs[26][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1799),
    .D(_01058_),
    .Q_N(_12906_),
    .Q(\top_ihp.oisc.regs[26][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1800),
    .D(_01059_),
    .Q_N(_12905_),
    .Q(\top_ihp.oisc.regs[26][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1801),
    .D(_01060_),
    .Q_N(_12904_),
    .Q(\top_ihp.oisc.regs[27][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1802),
    .D(_01061_),
    .Q_N(_12903_),
    .Q(\top_ihp.oisc.regs[27][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1803),
    .D(_01062_),
    .Q_N(_12902_),
    .Q(\top_ihp.oisc.regs[27][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][12]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1804),
    .D(_01063_),
    .Q_N(_12901_),
    .Q(\top_ihp.oisc.regs[27][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][13]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1805),
    .D(_01064_),
    .Q_N(_12900_),
    .Q(\top_ihp.oisc.regs[27][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][14]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1806),
    .D(_01065_),
    .Q_N(_12899_),
    .Q(\top_ihp.oisc.regs[27][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][15]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1807),
    .D(_01066_),
    .Q_N(_12898_),
    .Q(\top_ihp.oisc.regs[27][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][16]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1808),
    .D(_01067_),
    .Q_N(_12897_),
    .Q(\top_ihp.oisc.regs[27][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][17]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1809),
    .D(_01068_),
    .Q_N(_12896_),
    .Q(\top_ihp.oisc.regs[27][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][18]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1810),
    .D(_01069_),
    .Q_N(_12895_),
    .Q(\top_ihp.oisc.regs[27][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][19]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1811),
    .D(_01070_),
    .Q_N(_12894_),
    .Q(\top_ihp.oisc.regs[27][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1812),
    .D(_01071_),
    .Q_N(_12893_),
    .Q(\top_ihp.oisc.regs[27][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][20]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1813),
    .D(_01072_),
    .Q_N(_12892_),
    .Q(\top_ihp.oisc.regs[27][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][21]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1814),
    .D(_01073_),
    .Q_N(_12891_),
    .Q(\top_ihp.oisc.regs[27][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][22]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1815),
    .D(_01074_),
    .Q_N(_12890_),
    .Q(\top_ihp.oisc.regs[27][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][23]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1816),
    .D(_01075_),
    .Q_N(_12889_),
    .Q(\top_ihp.oisc.regs[27][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][24]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1817),
    .D(_01076_),
    .Q_N(_12888_),
    .Q(\top_ihp.oisc.regs[27][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][25]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1818),
    .D(_01077_),
    .Q_N(_12887_),
    .Q(\top_ihp.oisc.regs[27][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][26]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1819),
    .D(_01078_),
    .Q_N(_12886_),
    .Q(\top_ihp.oisc.regs[27][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][27]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1820),
    .D(_01079_),
    .Q_N(_12885_),
    .Q(\top_ihp.oisc.regs[27][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][28]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1821),
    .D(_01080_),
    .Q_N(_12884_),
    .Q(\top_ihp.oisc.regs[27][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][29]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1822),
    .D(_01081_),
    .Q_N(_12883_),
    .Q(\top_ihp.oisc.regs[27][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1823),
    .D(_01082_),
    .Q_N(_12882_),
    .Q(\top_ihp.oisc.regs[27][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][30]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1824),
    .D(_01083_),
    .Q_N(_12881_),
    .Q(\top_ihp.oisc.regs[27][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][31]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1825),
    .D(_01084_),
    .Q_N(_12880_),
    .Q(\top_ihp.oisc.regs[27][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1826),
    .D(_01085_),
    .Q_N(_12879_),
    .Q(\top_ihp.oisc.regs[27][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1827),
    .D(_01086_),
    .Q_N(_12878_),
    .Q(\top_ihp.oisc.regs[27][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1828),
    .D(_01087_),
    .Q_N(_12877_),
    .Q(\top_ihp.oisc.regs[27][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1829),
    .D(_01088_),
    .Q_N(_12876_),
    .Q(\top_ihp.oisc.regs[27][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1830),
    .D(_01089_),
    .Q_N(_12875_),
    .Q(\top_ihp.oisc.regs[27][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1831),
    .D(_01090_),
    .Q_N(_12874_),
    .Q(\top_ihp.oisc.regs[27][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1832),
    .D(_01091_),
    .Q_N(_12873_),
    .Q(\top_ihp.oisc.regs[27][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1833),
    .D(_01092_),
    .Q_N(_12872_),
    .Q(\top_ihp.oisc.regs[28][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1834),
    .D(_01093_),
    .Q_N(_12871_),
    .Q(\top_ihp.oisc.regs[28][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1835),
    .D(_01094_),
    .Q_N(_12870_),
    .Q(\top_ihp.oisc.regs[28][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][12]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1836),
    .D(_01095_),
    .Q_N(_12869_),
    .Q(\top_ihp.oisc.regs[28][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][13]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1837),
    .D(_01096_),
    .Q_N(_12868_),
    .Q(\top_ihp.oisc.regs[28][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][14]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1838),
    .D(_01097_),
    .Q_N(_12867_),
    .Q(\top_ihp.oisc.regs[28][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][15]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1839),
    .D(_01098_),
    .Q_N(_12866_),
    .Q(\top_ihp.oisc.regs[28][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][16]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1840),
    .D(_01099_),
    .Q_N(_12865_),
    .Q(\top_ihp.oisc.regs[28][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][17]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1841),
    .D(_01100_),
    .Q_N(_12864_),
    .Q(\top_ihp.oisc.regs[28][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][18]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1842),
    .D(_01101_),
    .Q_N(_12863_),
    .Q(\top_ihp.oisc.regs[28][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][19]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1843),
    .D(_01102_),
    .Q_N(_12862_),
    .Q(\top_ihp.oisc.regs[28][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1844),
    .D(_01103_),
    .Q_N(_12861_),
    .Q(\top_ihp.oisc.regs[28][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][20]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1845),
    .D(_01104_),
    .Q_N(_12860_),
    .Q(\top_ihp.oisc.regs[28][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][21]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1846),
    .D(_01105_),
    .Q_N(_12859_),
    .Q(\top_ihp.oisc.regs[28][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][22]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1847),
    .D(_01106_),
    .Q_N(_12858_),
    .Q(\top_ihp.oisc.regs[28][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][23]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1848),
    .D(_01107_),
    .Q_N(_12857_),
    .Q(\top_ihp.oisc.regs[28][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][24]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1849),
    .D(_01108_),
    .Q_N(_12856_),
    .Q(\top_ihp.oisc.regs[28][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][25]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1850),
    .D(_01109_),
    .Q_N(_12855_),
    .Q(\top_ihp.oisc.regs[28][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][26]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1851),
    .D(_01110_),
    .Q_N(_12854_),
    .Q(\top_ihp.oisc.regs[28][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][27]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1852),
    .D(_01111_),
    .Q_N(_12853_),
    .Q(\top_ihp.oisc.regs[28][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][28]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1853),
    .D(_01112_),
    .Q_N(_12852_),
    .Q(\top_ihp.oisc.regs[28][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][29]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1854),
    .D(_01113_),
    .Q_N(_12851_),
    .Q(\top_ihp.oisc.regs[28][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1855),
    .D(_01114_),
    .Q_N(_12850_),
    .Q(\top_ihp.oisc.regs[28][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][30]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1856),
    .D(_01115_),
    .Q_N(_12849_),
    .Q(\top_ihp.oisc.regs[28][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][31]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1857),
    .D(_01116_),
    .Q_N(_12848_),
    .Q(\top_ihp.oisc.regs[28][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1858),
    .D(_01117_),
    .Q_N(_12847_),
    .Q(\top_ihp.oisc.regs[28][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1859),
    .D(_01118_),
    .Q_N(_12846_),
    .Q(\top_ihp.oisc.regs[28][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1860),
    .D(_01119_),
    .Q_N(_12845_),
    .Q(\top_ihp.oisc.regs[28][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1861),
    .D(_01120_),
    .Q_N(_12844_),
    .Q(\top_ihp.oisc.regs[28][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1862),
    .D(_01121_),
    .Q_N(_12843_),
    .Q(\top_ihp.oisc.regs[28][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1863),
    .D(_01122_),
    .Q_N(_12842_),
    .Q(\top_ihp.oisc.regs[28][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1864),
    .D(_01123_),
    .Q_N(_12841_),
    .Q(\top_ihp.oisc.regs[28][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1865),
    .D(_01124_),
    .Q_N(_12840_),
    .Q(\top_ihp.oisc.regs[29][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1866),
    .D(_01125_),
    .Q_N(_12839_),
    .Q(\top_ihp.oisc.regs[29][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1867),
    .D(_01126_),
    .Q_N(_12838_),
    .Q(\top_ihp.oisc.regs[29][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][12]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1868),
    .D(_01127_),
    .Q_N(_12837_),
    .Q(\top_ihp.oisc.regs[29][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][13]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1869),
    .D(_01128_),
    .Q_N(_12836_),
    .Q(\top_ihp.oisc.regs[29][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][14]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1870),
    .D(_01129_),
    .Q_N(_12835_),
    .Q(\top_ihp.oisc.regs[29][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][15]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1871),
    .D(_01130_),
    .Q_N(_12834_),
    .Q(\top_ihp.oisc.regs[29][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][16]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1872),
    .D(_01131_),
    .Q_N(_12833_),
    .Q(\top_ihp.oisc.regs[29][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][17]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1873),
    .D(_01132_),
    .Q_N(_12832_),
    .Q(\top_ihp.oisc.regs[29][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][18]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1874),
    .D(_01133_),
    .Q_N(_12831_),
    .Q(\top_ihp.oisc.regs[29][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][19]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1875),
    .D(_01134_),
    .Q_N(_12830_),
    .Q(\top_ihp.oisc.regs[29][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1876),
    .D(_01135_),
    .Q_N(_12829_),
    .Q(\top_ihp.oisc.regs[29][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][20]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1877),
    .D(_01136_),
    .Q_N(_12828_),
    .Q(\top_ihp.oisc.regs[29][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][21]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1878),
    .D(_01137_),
    .Q_N(_12827_),
    .Q(\top_ihp.oisc.regs[29][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][22]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1879),
    .D(_01138_),
    .Q_N(_12826_),
    .Q(\top_ihp.oisc.regs[29][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][23]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1880),
    .D(_01139_),
    .Q_N(_12825_),
    .Q(\top_ihp.oisc.regs[29][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][24]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1881),
    .D(_01140_),
    .Q_N(_12824_),
    .Q(\top_ihp.oisc.regs[29][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][25]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1882),
    .D(_01141_),
    .Q_N(_12823_),
    .Q(\top_ihp.oisc.regs[29][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][26]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1883),
    .D(_01142_),
    .Q_N(_12822_),
    .Q(\top_ihp.oisc.regs[29][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][27]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1884),
    .D(_01143_),
    .Q_N(_12821_),
    .Q(\top_ihp.oisc.regs[29][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][28]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1885),
    .D(_01144_),
    .Q_N(_12820_),
    .Q(\top_ihp.oisc.regs[29][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][29]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1886),
    .D(_01145_),
    .Q_N(_12819_),
    .Q(\top_ihp.oisc.regs[29][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1887),
    .D(_01146_),
    .Q_N(_12818_),
    .Q(\top_ihp.oisc.regs[29][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][30]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1888),
    .D(_01147_),
    .Q_N(_12817_),
    .Q(\top_ihp.oisc.regs[29][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][31]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1889),
    .D(_01148_),
    .Q_N(_12816_),
    .Q(\top_ihp.oisc.regs[29][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1890),
    .D(_01149_),
    .Q_N(_12815_),
    .Q(\top_ihp.oisc.regs[29][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1891),
    .D(_01150_),
    .Q_N(_12814_),
    .Q(\top_ihp.oisc.regs[29][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1892),
    .D(_01151_),
    .Q_N(_12813_),
    .Q(\top_ihp.oisc.regs[29][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1893),
    .D(_01152_),
    .Q_N(_12812_),
    .Q(\top_ihp.oisc.regs[29][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1894),
    .D(_01153_),
    .Q_N(_12811_),
    .Q(\top_ihp.oisc.regs[29][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1895),
    .D(_01154_),
    .Q_N(_12810_),
    .Q(\top_ihp.oisc.regs[29][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1896),
    .D(_01155_),
    .Q_N(_12809_),
    .Q(\top_ihp.oisc.regs[29][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1212),
    .D(_01156_),
    .Q_N(_12808_),
    .Q(\top_ihp.oisc.regs[2][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1167),
    .D(_01157_),
    .Q_N(_12807_),
    .Q(\top_ihp.oisc.regs[2][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1175),
    .D(_01158_),
    .Q_N(_12806_),
    .Q(\top_ihp.oisc.regs[2][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1220),
    .D(_01159_),
    .Q_N(_12805_),
    .Q(\top_ihp.oisc.regs[2][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1168),
    .D(_01160_),
    .Q_N(_12804_),
    .Q(\top_ihp.oisc.regs[2][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1211),
    .D(_01161_),
    .Q_N(_12803_),
    .Q(\top_ihp.oisc.regs[2][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1177),
    .D(_01162_),
    .Q_N(_12802_),
    .Q(\top_ihp.oisc.regs[2][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1212),
    .D(_01163_),
    .Q_N(_12801_),
    .Q(\top_ihp.oisc.regs[2][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1166),
    .D(_01164_),
    .Q_N(_12800_),
    .Q(\top_ihp.oisc.regs[2][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1170),
    .D(_01165_),
    .Q_N(_12799_),
    .Q(\top_ihp.oisc.regs[2][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1172),
    .D(_01166_),
    .Q_N(_12798_),
    .Q(\top_ihp.oisc.regs[2][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1179),
    .D(_01167_),
    .Q_N(_12797_),
    .Q(\top_ihp.oisc.regs[2][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1239),
    .D(_01168_),
    .Q_N(_12796_),
    .Q(\top_ihp.oisc.regs[2][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1188),
    .D(_01169_),
    .Q_N(_12795_),
    .Q(\top_ihp.oisc.regs[2][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1223),
    .D(_01170_),
    .Q_N(_12794_),
    .Q(\top_ihp.oisc.regs[2][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1181),
    .D(_01171_),
    .Q_N(_12793_),
    .Q(\top_ihp.oisc.regs[2][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1232),
    .D(_01172_),
    .Q_N(_12792_),
    .Q(\top_ihp.oisc.regs[2][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1172),
    .D(_01173_),
    .Q_N(_12791_),
    .Q(\top_ihp.oisc.regs[2][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1196),
    .D(_01174_),
    .Q_N(_12790_),
    .Q(\top_ihp.oisc.regs[2][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1188),
    .D(_01175_),
    .Q_N(_12789_),
    .Q(\top_ihp.oisc.regs[2][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1203),
    .D(_01176_),
    .Q_N(_12788_),
    .Q(\top_ihp.oisc.regs[2][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1204),
    .D(_01177_),
    .Q_N(_12787_),
    .Q(\top_ihp.oisc.regs[2][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1243),
    .D(_01178_),
    .Q_N(_12786_),
    .Q(\top_ihp.oisc.regs[2][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1194),
    .D(_01179_),
    .Q_N(_12785_),
    .Q(\top_ihp.oisc.regs[2][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1201),
    .D(_01180_),
    .Q_N(_12784_),
    .Q(\top_ihp.oisc.regs[2][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1194),
    .D(_01181_),
    .Q_N(_12783_),
    .Q(\top_ihp.oisc.regs[2][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1194),
    .D(_01182_),
    .Q_N(_12782_),
    .Q(\top_ihp.oisc.regs[2][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1194),
    .D(_01183_),
    .Q_N(_12781_),
    .Q(\top_ihp.oisc.regs[2][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1243),
    .D(_01184_),
    .Q_N(_12780_),
    .Q(\top_ihp.oisc.regs[2][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1237),
    .D(_01185_),
    .Q_N(_12779_),
    .Q(\top_ihp.oisc.regs[2][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1239),
    .D(_01186_),
    .Q_N(_12778_),
    .Q(\top_ihp.oisc.regs[2][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1216),
    .D(_01187_),
    .Q_N(_12777_),
    .Q(\top_ihp.oisc.regs[2][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1897),
    .D(_01188_),
    .Q_N(_12776_),
    .Q(\top_ihp.oisc.regs[30][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1898),
    .D(_01189_),
    .Q_N(_12775_),
    .Q(\top_ihp.oisc.regs[30][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1899),
    .D(_01190_),
    .Q_N(_12774_),
    .Q(\top_ihp.oisc.regs[30][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][12]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1900),
    .D(_01191_),
    .Q_N(_12773_),
    .Q(\top_ihp.oisc.regs[30][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][13]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1901),
    .D(_01192_),
    .Q_N(_12772_),
    .Q(\top_ihp.oisc.regs[30][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][14]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1902),
    .D(_01193_),
    .Q_N(_12771_),
    .Q(\top_ihp.oisc.regs[30][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][15]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1903),
    .D(_01194_),
    .Q_N(_12770_),
    .Q(\top_ihp.oisc.regs[30][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][16]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1904),
    .D(_01195_),
    .Q_N(_12769_),
    .Q(\top_ihp.oisc.regs[30][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][17]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1905),
    .D(_01196_),
    .Q_N(_12768_),
    .Q(\top_ihp.oisc.regs[30][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][18]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1906),
    .D(_01197_),
    .Q_N(_12767_),
    .Q(\top_ihp.oisc.regs[30][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][19]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1907),
    .D(_01198_),
    .Q_N(_12766_),
    .Q(\top_ihp.oisc.regs[30][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1908),
    .D(_01199_),
    .Q_N(_12765_),
    .Q(\top_ihp.oisc.regs[30][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][20]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1909),
    .D(_01200_),
    .Q_N(_12764_),
    .Q(\top_ihp.oisc.regs[30][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][21]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1910),
    .D(_01201_),
    .Q_N(_12763_),
    .Q(\top_ihp.oisc.regs[30][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][22]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1911),
    .D(_01202_),
    .Q_N(_12762_),
    .Q(\top_ihp.oisc.regs[30][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][23]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1912),
    .D(_01203_),
    .Q_N(_12761_),
    .Q(\top_ihp.oisc.regs[30][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][24]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1913),
    .D(_01204_),
    .Q_N(_12760_),
    .Q(\top_ihp.oisc.regs[30][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][25]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1914),
    .D(_01205_),
    .Q_N(_12759_),
    .Q(\top_ihp.oisc.regs[30][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][26]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1915),
    .D(_01206_),
    .Q_N(_12758_),
    .Q(\top_ihp.oisc.regs[30][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][27]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1916),
    .D(_01207_),
    .Q_N(_12757_),
    .Q(\top_ihp.oisc.regs[30][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][28]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1917),
    .D(_01208_),
    .Q_N(_12756_),
    .Q(\top_ihp.oisc.regs[30][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][29]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1918),
    .D(_01209_),
    .Q_N(_12755_),
    .Q(\top_ihp.oisc.regs[30][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1919),
    .D(_01210_),
    .Q_N(_12754_),
    .Q(\top_ihp.oisc.regs[30][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][30]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1920),
    .D(_01211_),
    .Q_N(_12753_),
    .Q(\top_ihp.oisc.regs[30][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][31]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1921),
    .D(_01212_),
    .Q_N(_12752_),
    .Q(\top_ihp.oisc.regs[30][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1922),
    .D(_01213_),
    .Q_N(_12751_),
    .Q(\top_ihp.oisc.regs[30][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1923),
    .D(_01214_),
    .Q_N(_12750_),
    .Q(\top_ihp.oisc.regs[30][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1924),
    .D(_01215_),
    .Q_N(_12749_),
    .Q(\top_ihp.oisc.regs[30][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1925),
    .D(_01216_),
    .Q_N(_12748_),
    .Q(\top_ihp.oisc.regs[30][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1926),
    .D(_01217_),
    .Q_N(_12747_),
    .Q(\top_ihp.oisc.regs[30][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1927),
    .D(_01218_),
    .Q_N(_12746_),
    .Q(\top_ihp.oisc.regs[30][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1928),
    .D(_01219_),
    .Q_N(_12745_),
    .Q(\top_ihp.oisc.regs[30][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1929),
    .D(_01220_),
    .Q_N(_12744_),
    .Q(\top_ihp.oisc.regs[31][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1930),
    .D(_01221_),
    .Q_N(_12743_),
    .Q(\top_ihp.oisc.regs[31][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1931),
    .D(_01222_),
    .Q_N(_12742_),
    .Q(\top_ihp.oisc.regs[31][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][12]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1932),
    .D(_01223_),
    .Q_N(_12741_),
    .Q(\top_ihp.oisc.regs[31][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][13]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1933),
    .D(_01224_),
    .Q_N(_12740_),
    .Q(\top_ihp.oisc.regs[31][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][14]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1934),
    .D(_01225_),
    .Q_N(_12739_),
    .Q(\top_ihp.oisc.regs[31][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][15]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1935),
    .D(_01226_),
    .Q_N(_12738_),
    .Q(\top_ihp.oisc.regs[31][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][16]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1936),
    .D(_01227_),
    .Q_N(_12737_),
    .Q(\top_ihp.oisc.regs[31][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][17]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1937),
    .D(_01228_),
    .Q_N(_12736_),
    .Q(\top_ihp.oisc.regs[31][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][18]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1938),
    .D(_01229_),
    .Q_N(_12735_),
    .Q(\top_ihp.oisc.regs[31][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][19]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1939),
    .D(_01230_),
    .Q_N(_12734_),
    .Q(\top_ihp.oisc.regs[31][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1940),
    .D(_01231_),
    .Q_N(_12733_),
    .Q(\top_ihp.oisc.regs[31][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][20]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1941),
    .D(_01232_),
    .Q_N(_12732_),
    .Q(\top_ihp.oisc.regs[31][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][21]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1942),
    .D(_01233_),
    .Q_N(_12731_),
    .Q(\top_ihp.oisc.regs[31][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][22]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1943),
    .D(_01234_),
    .Q_N(_12730_),
    .Q(\top_ihp.oisc.regs[31][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][23]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1944),
    .D(_01235_),
    .Q_N(_12729_),
    .Q(\top_ihp.oisc.regs[31][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][24]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1945),
    .D(_01236_),
    .Q_N(_12728_),
    .Q(\top_ihp.oisc.regs[31][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][25]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1946),
    .D(_01237_),
    .Q_N(_12727_),
    .Q(\top_ihp.oisc.regs[31][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][26]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1947),
    .D(_01238_),
    .Q_N(_12726_),
    .Q(\top_ihp.oisc.regs[31][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][27]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1948),
    .D(_01239_),
    .Q_N(_12725_),
    .Q(\top_ihp.oisc.regs[31][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][28]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1949),
    .D(_01240_),
    .Q_N(_12724_),
    .Q(\top_ihp.oisc.regs[31][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][29]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1950),
    .D(_01241_),
    .Q_N(_12723_),
    .Q(\top_ihp.oisc.regs[31][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1951),
    .D(_01242_),
    .Q_N(_12722_),
    .Q(\top_ihp.oisc.regs[31][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][30]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1952),
    .D(_01243_),
    .Q_N(_12721_),
    .Q(\top_ihp.oisc.regs[31][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][31]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1953),
    .D(_01244_),
    .Q_N(_12720_),
    .Q(\top_ihp.oisc.regs[31][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1954),
    .D(_01245_),
    .Q_N(_12719_),
    .Q(\top_ihp.oisc.regs[31][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1955),
    .D(_01246_),
    .Q_N(_12718_),
    .Q(\top_ihp.oisc.regs[31][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1956),
    .D(_01247_),
    .Q_N(_12717_),
    .Q(\top_ihp.oisc.regs[31][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1957),
    .D(_01248_),
    .Q_N(_12716_),
    .Q(\top_ihp.oisc.regs[31][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1958),
    .D(_01249_),
    .Q_N(_12715_),
    .Q(\top_ihp.oisc.regs[31][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1959),
    .D(_01250_),
    .Q_N(_12714_),
    .Q(\top_ihp.oisc.regs[31][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1960),
    .D(_01251_),
    .Q_N(_12713_),
    .Q(\top_ihp.oisc.regs[31][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1961),
    .D(_01252_),
    .Q_N(_12712_),
    .Q(\top_ihp.oisc.regs[32][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][10]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1962),
    .D(_01253_),
    .Q_N(_12711_),
    .Q(\top_ihp.oisc.regs[32][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][11]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1963),
    .D(_01254_),
    .Q_N(_12710_),
    .Q(\top_ihp.oisc.regs[32][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][12]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1964),
    .D(_01255_),
    .Q_N(_12709_),
    .Q(\top_ihp.oisc.regs[32][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][13]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1965),
    .D(_01256_),
    .Q_N(_12708_),
    .Q(\top_ihp.oisc.regs[32][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][14]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1966),
    .D(_01257_),
    .Q_N(_12707_),
    .Q(\top_ihp.oisc.regs[32][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][15]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1967),
    .D(_01258_),
    .Q_N(_12706_),
    .Q(\top_ihp.oisc.regs[32][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][16]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1968),
    .D(_01259_),
    .Q_N(_12705_),
    .Q(\top_ihp.oisc.regs[32][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][17]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1969),
    .D(_01260_),
    .Q_N(_12704_),
    .Q(\top_ihp.oisc.regs[32][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][18]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1970),
    .D(_01261_),
    .Q_N(_12703_),
    .Q(\top_ihp.oisc.regs[32][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][19]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1971),
    .D(_01262_),
    .Q_N(_12702_),
    .Q(\top_ihp.oisc.regs[32][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][1]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1972),
    .D(_01263_),
    .Q_N(_12701_),
    .Q(\top_ihp.oisc.regs[32][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][20]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1973),
    .D(_01264_),
    .Q_N(_12700_),
    .Q(\top_ihp.oisc.regs[32][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][21]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1974),
    .D(_01265_),
    .Q_N(_12699_),
    .Q(\top_ihp.oisc.regs[32][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][22]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1975),
    .D(_01266_),
    .Q_N(_12698_),
    .Q(\top_ihp.oisc.regs[32][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][23]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1976),
    .D(_01267_),
    .Q_N(_12697_),
    .Q(\top_ihp.oisc.regs[32][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][24]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1977),
    .D(_01268_),
    .Q_N(_12696_),
    .Q(\top_ihp.oisc.regs[32][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][25]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1978),
    .D(_01269_),
    .Q_N(_12695_),
    .Q(\top_ihp.oisc.regs[32][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][26]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1979),
    .D(_01270_),
    .Q_N(_12694_),
    .Q(\top_ihp.oisc.regs[32][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][27]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1980),
    .D(_01271_),
    .Q_N(_12693_),
    .Q(\top_ihp.oisc.regs[32][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][28]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1981),
    .D(_01272_),
    .Q_N(_12692_),
    .Q(\top_ihp.oisc.regs[32][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][29]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1982),
    .D(_01273_),
    .Q_N(_12691_),
    .Q(\top_ihp.oisc.regs[32][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][2]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1983),
    .D(_01274_),
    .Q_N(_12690_),
    .Q(\top_ihp.oisc.regs[32][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][30]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1984),
    .D(_01275_),
    .Q_N(_12689_),
    .Q(\top_ihp.oisc.regs[32][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][31]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1985),
    .D(_01276_),
    .Q_N(_12688_),
    .Q(\top_ihp.oisc.regs[32][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][3]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1986),
    .D(_01277_),
    .Q_N(_12687_),
    .Q(\top_ihp.oisc.regs[32][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][4]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1987),
    .D(_01278_),
    .Q_N(_12686_),
    .Q(\top_ihp.oisc.regs[32][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][5]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1988),
    .D(_01279_),
    .Q_N(_12685_),
    .Q(\top_ihp.oisc.regs[32][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][6]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1989),
    .D(_01280_),
    .Q_N(_12684_),
    .Q(\top_ihp.oisc.regs[32][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][7]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1990),
    .D(_01281_),
    .Q_N(_12683_),
    .Q(\top_ihp.oisc.regs[32][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][8]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1991),
    .D(_01282_),
    .Q_N(_12682_),
    .Q(\top_ihp.oisc.regs[32][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][9]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1992),
    .D(_01283_),
    .Q_N(_12681_),
    .Q(\top_ihp.oisc.regs[32][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1315),
    .D(_01284_),
    .Q_N(_12680_),
    .Q(\top_ihp.oisc.regs[33][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1364),
    .D(_01285_),
    .Q_N(_12679_),
    .Q(\top_ihp.oisc.regs[33][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1315),
    .D(_01286_),
    .Q_N(_12678_),
    .Q(\top_ihp.oisc.regs[33][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1265),
    .D(_01287_),
    .Q_N(_12677_),
    .Q(\top_ihp.oisc.regs[33][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1317),
    .D(_01288_),
    .Q_N(_12676_),
    .Q(\top_ihp.oisc.regs[33][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1265),
    .D(_01289_),
    .Q_N(_12675_),
    .Q(\top_ihp.oisc.regs[33][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1265),
    .D(_01290_),
    .Q_N(_12674_),
    .Q(\top_ihp.oisc.regs[33][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1364),
    .D(_01291_),
    .Q_N(_12673_),
    .Q(\top_ihp.oisc.regs[33][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1315),
    .D(_01292_),
    .Q_N(_12672_),
    .Q(\top_ihp.oisc.regs[33][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1315),
    .D(_01293_),
    .Q_N(_12671_),
    .Q(\top_ihp.oisc.regs[33][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1372),
    .D(_01294_),
    .Q_N(_12670_),
    .Q(\top_ihp.oisc.regs[33][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1267),
    .D(_01295_),
    .Q_N(_12669_),
    .Q(\top_ihp.oisc.regs[33][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1349),
    .D(_01296_),
    .Q_N(_12668_),
    .Q(\top_ihp.oisc.regs[33][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1372),
    .D(_01297_),
    .Q_N(_12667_),
    .Q(\top_ihp.oisc.regs[33][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1268),
    .D(_01298_),
    .Q_N(_12666_),
    .Q(\top_ihp.oisc.regs[33][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1270),
    .D(_01299_),
    .Q_N(_12665_),
    .Q(\top_ihp.oisc.regs[33][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1329),
    .D(_01300_),
    .Q_N(_12664_),
    .Q(\top_ihp.oisc.regs[33][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1309),
    .D(_01301_),
    .Q_N(_12663_),
    .Q(\top_ihp.oisc.regs[33][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1396),
    .D(_01302_),
    .Q_N(_12662_),
    .Q(\top_ihp.oisc.regs[33][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1396),
    .D(_01303_),
    .Q_N(_12661_),
    .Q(\top_ihp.oisc.regs[33][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1330),
    .D(_01304_),
    .Q_N(_12660_),
    .Q(\top_ihp.oisc.regs[33][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1338),
    .D(_01305_),
    .Q_N(_12659_),
    .Q(\top_ihp.oisc.regs[33][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1355),
    .D(_01306_),
    .Q_N(_12658_),
    .Q(\top_ihp.oisc.regs[33][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1339),
    .D(_01307_),
    .Q_N(_12657_),
    .Q(\top_ihp.oisc.regs[33][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1341),
    .D(_01308_),
    .Q_N(_12656_),
    .Q(\top_ihp.oisc.regs[33][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1341),
    .D(_01309_),
    .Q_N(_12655_),
    .Q(\top_ihp.oisc.regs[33][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1290),
    .D(_01310_),
    .Q_N(_12654_),
    .Q(\top_ihp.oisc.regs[33][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1292),
    .D(_01311_),
    .Q_N(_12653_),
    .Q(\top_ihp.oisc.regs[33][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1281),
    .D(_01312_),
    .Q_N(_12652_),
    .Q(\top_ihp.oisc.regs[33][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1347),
    .D(_01313_),
    .Q_N(_12651_),
    .Q(\top_ihp.oisc.regs[33][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1281),
    .D(_01314_),
    .Q_N(_12650_),
    .Q(\top_ihp.oisc.regs[33][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1277),
    .D(_01315_),
    .Q_N(_12649_),
    .Q(\top_ihp.oisc.regs[33][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1302),
    .D(_01316_),
    .Q_N(_12648_),
    .Q(\top_ihp.oisc.regs[34][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1364),
    .D(_01317_),
    .Q_N(_12647_),
    .Q(\top_ihp.oisc.regs[34][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1364),
    .D(_01318_),
    .Q_N(_12646_),
    .Q(\top_ihp.oisc.regs[34][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1301),
    .D(_01319_),
    .Q_N(_12645_),
    .Q(\top_ihp.oisc.regs[34][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1317),
    .D(_01320_),
    .Q_N(_12644_),
    .Q(\top_ihp.oisc.regs[34][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1299),
    .D(_01321_),
    .Q_N(_12643_),
    .Q(\top_ihp.oisc.regs[34][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][15]$_DFFE_PN1P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1249),
    .D(_01322_),
    .Q_N(\top_ihp.oisc.regs[34][15] ),
    .Q(_00304_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1364),
    .D(_01323_),
    .Q_N(_12642_),
    .Q(\top_ihp.oisc.regs[34][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1307),
    .D(_01324_),
    .Q_N(_12641_),
    .Q(\top_ihp.oisc.regs[34][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1319),
    .D(_01325_),
    .Q_N(_12640_),
    .Q(\top_ihp.oisc.regs[34][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1364),
    .D(_01326_),
    .Q_N(_12639_),
    .Q(\top_ihp.oisc.regs[34][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1270),
    .D(_01327_),
    .Q_N(_12638_),
    .Q(\top_ihp.oisc.regs[34][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1276),
    .D(_01328_),
    .Q_N(_12637_),
    .Q(\top_ihp.oisc.regs[34][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1372),
    .D(_01329_),
    .Q_N(_12636_),
    .Q(\top_ihp.oisc.regs[34][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1268),
    .D(_01330_),
    .Q_N(_12635_),
    .Q(\top_ihp.oisc.regs[34][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1256),
    .D(_01331_),
    .Q_N(_12634_),
    .Q(\top_ihp.oisc.regs[34][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1276),
    .D(_01332_),
    .Q_N(_12633_),
    .Q(\top_ihp.oisc.regs[34][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1256),
    .D(_01333_),
    .Q_N(_12632_),
    .Q(\top_ihp.oisc.regs[34][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1396),
    .D(_01334_),
    .Q_N(_12631_),
    .Q(\top_ihp.oisc.regs[34][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1396),
    .D(_01335_),
    .Q_N(_12630_),
    .Q(\top_ihp.oisc.regs[34][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1277),
    .D(_01336_),
    .Q_N(_12629_),
    .Q(\top_ihp.oisc.regs[34][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1336),
    .D(_01337_),
    .Q_N(_12628_),
    .Q(\top_ihp.oisc.regs[34][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1402),
    .D(_01338_),
    .Q_N(_12627_),
    .Q(\top_ihp.oisc.regs[34][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1402),
    .D(_01339_),
    .Q_N(_12626_),
    .Q(\top_ihp.oisc.regs[34][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][31]$_DFFE_PN1P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1279),
    .D(_01340_),
    .Q_N(\top_ihp.oisc.regs[34][31] ),
    .Q(_00305_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1330),
    .D(_01341_),
    .Q_N(_12625_),
    .Q(\top_ihp.oisc.regs[34][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1280),
    .D(_01342_),
    .Q_N(_12624_),
    .Q(\top_ihp.oisc.regs[34][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1402),
    .D(_01343_),
    .Q_N(_12623_),
    .Q(\top_ihp.oisc.regs[34][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1281),
    .D(_01344_),
    .Q_N(_12622_),
    .Q(\top_ihp.oisc.regs[34][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1347),
    .D(_01345_),
    .Q_N(_12621_),
    .Q(\top_ihp.oisc.regs[34][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1277),
    .D(_01346_),
    .Q_N(_12620_),
    .Q(\top_ihp.oisc.regs[34][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1276),
    .D(_01347_),
    .Q_N(_12619_),
    .Q(\top_ihp.oisc.regs[34][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1315),
    .D(_01348_),
    .Q_N(_12618_),
    .Q(\top_ihp.oisc.regs[35][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1260),
    .D(_01349_),
    .Q_N(_12617_),
    .Q(\top_ihp.oisc.regs[35][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][11]$_DFFE_PN1P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1313),
    .D(_01350_),
    .Q_N(\top_ihp.oisc.regs[35][11] ),
    .Q(_00306_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1259),
    .D(_01351_),
    .Q_N(_12616_),
    .Q(\top_ihp.oisc.regs[35][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1313),
    .D(_01352_),
    .Q_N(_12615_),
    .Q(\top_ihp.oisc.regs[35][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1297),
    .D(_01353_),
    .Q_N(_12614_),
    .Q(\top_ihp.oisc.regs[35][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1297),
    .D(_01354_),
    .Q_N(_12613_),
    .Q(\top_ihp.oisc.regs[35][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1251),
    .D(_01355_),
    .Q_N(_12612_),
    .Q(\top_ihp.oisc.regs[35][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1321),
    .D(_01356_),
    .Q_N(_12611_),
    .Q(\top_ihp.oisc.regs[35][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1371),
    .D(_01357_),
    .Q_N(_12610_),
    .Q(\top_ihp.oisc.regs[35][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1371),
    .D(_01358_),
    .Q_N(_12609_),
    .Q(\top_ihp.oisc.regs[35][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1267),
    .D(_01359_),
    .Q_N(_12608_),
    .Q(\top_ihp.oisc.regs[35][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1276),
    .D(_01360_),
    .Q_N(_12607_),
    .Q(\top_ihp.oisc.regs[35][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1372),
    .D(_01361_),
    .Q_N(_12606_),
    .Q(\top_ihp.oisc.regs[35][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1268),
    .D(_01362_),
    .Q_N(_12605_),
    .Q(\top_ihp.oisc.regs[35][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1254),
    .D(_01363_),
    .Q_N(_12604_),
    .Q(\top_ihp.oisc.regs[35][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1275),
    .D(_01364_),
    .Q_N(_12603_),
    .Q(\top_ihp.oisc.regs[35][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1304),
    .D(_01365_),
    .Q_N(_12602_),
    .Q(\top_ihp.oisc.regs[35][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1395),
    .D(_01366_),
    .Q_N(_12601_),
    .Q(\top_ihp.oisc.regs[35][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1330),
    .D(_01367_),
    .Q_N(_12600_),
    .Q(\top_ihp.oisc.regs[35][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1330),
    .D(_01368_),
    .Q_N(_12599_),
    .Q(\top_ihp.oisc.regs[35][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1282),
    .D(_01369_),
    .Q_N(_12598_),
    .Q(\top_ihp.oisc.regs[35][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1404),
    .D(_01370_),
    .Q_N(_12597_),
    .Q(\top_ihp.oisc.regs[35][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1404),
    .D(_01371_),
    .Q_N(_12596_),
    .Q(\top_ihp.oisc.regs[35][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][31]$_DFFE_PN1P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1281),
    .D(_01372_),
    .Q_N(\top_ihp.oisc.regs[35][31] ),
    .Q(_00307_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1343),
    .D(_01373_),
    .Q_N(_12595_),
    .Q(\top_ihp.oisc.regs[35][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1288),
    .D(_01374_),
    .Q_N(_12594_),
    .Q(\top_ihp.oisc.regs[35][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1402),
    .D(_01375_),
    .Q_N(_12593_),
    .Q(\top_ihp.oisc.regs[35][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1281),
    .D(_01376_),
    .Q_N(_12592_),
    .Q(\top_ihp.oisc.regs[35][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1281),
    .D(_01377_),
    .Q_N(_12591_),
    .Q(\top_ihp.oisc.regs[35][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1284),
    .D(_01378_),
    .Q_N(_12590_),
    .Q(\top_ihp.oisc.regs[35][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1276),
    .D(_01379_),
    .Q_N(_12589_),
    .Q(\top_ihp.oisc.regs[35][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1251),
    .D(_01380_),
    .Q_N(_12588_),
    .Q(\top_ihp.oisc.regs[36][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1319),
    .D(_01381_),
    .Q_N(_12587_),
    .Q(\top_ihp.oisc.regs[36][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1364),
    .D(_01382_),
    .Q_N(_12586_),
    .Q(\top_ihp.oisc.regs[36][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1260),
    .D(_01383_),
    .Q_N(_12585_),
    .Q(\top_ihp.oisc.regs[36][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1379),
    .D(_01384_),
    .Q_N(_12584_),
    .Q(\top_ihp.oisc.regs[36][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1251),
    .D(_01385_),
    .Q_N(_12583_),
    .Q(\top_ihp.oisc.regs[36][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1259),
    .D(_01386_),
    .Q_N(_12582_),
    .Q(\top_ihp.oisc.regs[36][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1251),
    .D(_01387_),
    .Q_N(_12581_),
    .Q(\top_ihp.oisc.regs[36][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1386),
    .D(_01388_),
    .Q_N(_12580_),
    .Q(\top_ihp.oisc.regs[36][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1387),
    .D(_01389_),
    .Q_N(_12579_),
    .Q(\top_ihp.oisc.regs[36][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1388),
    .D(_01390_),
    .Q_N(_12578_),
    .Q(\top_ihp.oisc.regs[36][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1267),
    .D(_01391_),
    .Q_N(_12577_),
    .Q(\top_ihp.oisc.regs[36][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1329),
    .D(_01392_),
    .Q_N(_12576_),
    .Q(\top_ihp.oisc.regs[36][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1388),
    .D(_01393_),
    .Q_N(_12575_),
    .Q(\top_ihp.oisc.regs[36][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1256),
    .D(_01394_),
    .Q_N(_12574_),
    .Q(\top_ihp.oisc.regs[36][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1411),
    .D(_01395_),
    .Q_N(_12573_),
    .Q(\top_ihp.oisc.regs[36][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1413),
    .D(_01396_),
    .Q_N(_12572_),
    .Q(\top_ihp.oisc.regs[36][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1268),
    .D(_01397_),
    .Q_N(_12571_),
    .Q(\top_ihp.oisc.regs[36][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1333),
    .D(_01398_),
    .Q_N(_12570_),
    .Q(\top_ihp.oisc.regs[36][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1413),
    .D(_01399_),
    .Q_N(_12569_),
    .Q(\top_ihp.oisc.regs[36][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1421),
    .D(_01400_),
    .Q_N(_12568_),
    .Q(\top_ihp.oisc.regs[36][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1342),
    .D(_01401_),
    .Q_N(_12567_),
    .Q(\top_ihp.oisc.regs[36][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1339),
    .D(_01402_),
    .Q_N(_12566_),
    .Q(\top_ihp.oisc.regs[36][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1343),
    .D(_01403_),
    .Q_N(_12565_),
    .Q(\top_ihp.oisc.regs[36][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1355),
    .D(_01404_),
    .Q_N(_12564_),
    .Q(\top_ihp.oisc.regs[36][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1336),
    .D(_01405_),
    .Q_N(_12563_),
    .Q(\top_ihp.oisc.regs[36][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1288),
    .D(_01406_),
    .Q_N(_12562_),
    .Q(\top_ihp.oisc.regs[36][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1291),
    .D(_01407_),
    .Q_N(_12561_),
    .Q(\top_ihp.oisc.regs[36][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1284),
    .D(_01408_),
    .Q_N(_12560_),
    .Q(\top_ihp.oisc.regs[36][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1347),
    .D(_01409_),
    .Q_N(_12559_),
    .Q(\top_ihp.oisc.regs[36][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1329),
    .D(_01410_),
    .Q_N(_12558_),
    .Q(\top_ihp.oisc.regs[36][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1412),
    .D(_01411_),
    .Q_N(_12557_),
    .Q(\top_ihp.oisc.regs[36][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1380),
    .D(_01412_),
    .Q_N(_12556_),
    .Q(\top_ihp.oisc.regs[37][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1302),
    .D(_01413_),
    .Q_N(_12555_),
    .Q(\top_ihp.oisc.regs[37][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1301),
    .D(_01414_),
    .Q_N(_12554_),
    .Q(\top_ihp.oisc.regs[37][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1261),
    .D(_01415_),
    .Q_N(_12553_),
    .Q(\top_ihp.oisc.regs[37][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1380),
    .D(_01416_),
    .Q_N(_12552_),
    .Q(\top_ihp.oisc.regs[37][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1263),
    .D(_01417_),
    .Q_N(_12551_),
    .Q(\top_ihp.oisc.regs[37][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1263),
    .D(_01418_),
    .Q_N(_12550_),
    .Q(\top_ihp.oisc.regs[37][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1381),
    .D(_01419_),
    .Q_N(_12549_),
    .Q(\top_ihp.oisc.regs[37][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1390),
    .D(_01420_),
    .Q_N(_12548_),
    .Q(\top_ihp.oisc.regs[37][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1387),
    .D(_01421_),
    .Q_N(_12547_),
    .Q(\top_ihp.oisc.regs[37][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1390),
    .D(_01422_),
    .Q_N(_12546_),
    .Q(\top_ihp.oisc.regs[37][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1253),
    .D(_01423_),
    .Q_N(_12545_),
    .Q(\top_ihp.oisc.regs[37][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1412),
    .D(_01424_),
    .Q_N(_12544_),
    .Q(\top_ihp.oisc.regs[37][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1392),
    .D(_01425_),
    .Q_N(_12543_),
    .Q(\top_ihp.oisc.regs[37][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1256),
    .D(_01426_),
    .Q_N(_12542_),
    .Q(\top_ihp.oisc.regs[37][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1322),
    .D(_01427_),
    .Q_N(_12541_),
    .Q(\top_ihp.oisc.regs[37][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1414),
    .D(_01428_),
    .Q_N(_12540_),
    .Q(\top_ihp.oisc.regs[37][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1255),
    .D(_01429_),
    .Q_N(_12539_),
    .Q(\top_ihp.oisc.regs[37][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1347),
    .D(_01430_),
    .Q_N(_12538_),
    .Q(\top_ihp.oisc.regs[37][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1414),
    .D(_01431_),
    .Q_N(_12537_),
    .Q(\top_ihp.oisc.regs[37][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1404),
    .D(_01432_),
    .Q_N(_12536_),
    .Q(\top_ihp.oisc.regs[37][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1360),
    .D(_01433_),
    .Q_N(_12535_),
    .Q(\top_ihp.oisc.regs[37][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1422),
    .D(_01434_),
    .Q_N(_12534_),
    .Q(\top_ihp.oisc.regs[37][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1421),
    .D(_01435_),
    .Q_N(_12533_),
    .Q(\top_ihp.oisc.regs[37][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1341),
    .D(_01436_),
    .Q_N(_12532_),
    .Q(\top_ihp.oisc.regs[37][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1291),
    .D(_01437_),
    .Q_N(_12531_),
    .Q(\top_ihp.oisc.regs[37][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1293),
    .D(_01438_),
    .Q_N(_12530_),
    .Q(\top_ihp.oisc.regs[37][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1354),
    .D(_01439_),
    .Q_N(_12529_),
    .Q(\top_ihp.oisc.regs[37][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1285),
    .D(_01440_),
    .Q_N(_12528_),
    .Q(\top_ihp.oisc.regs[37][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1333),
    .D(_01441_),
    .Q_N(_12527_),
    .Q(\top_ihp.oisc.regs[37][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1334),
    .D(_01442_),
    .Q_N(_12526_),
    .Q(\top_ihp.oisc.regs[37][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1333),
    .D(_01443_),
    .Q_N(_12525_),
    .Q(\top_ihp.oisc.regs[37][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1383),
    .D(_01444_),
    .Q_N(_12524_),
    .Q(\top_ihp.oisc.regs[38][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1383),
    .D(_01445_),
    .Q_N(_12523_),
    .Q(\top_ihp.oisc.regs[38][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1381),
    .D(_01446_),
    .Q_N(_12522_),
    .Q(\top_ihp.oisc.regs[38][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1263),
    .D(_01447_),
    .Q_N(_12521_),
    .Q(\top_ihp.oisc.regs[38][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1381),
    .D(_01448_),
    .Q_N(_12520_),
    .Q(\top_ihp.oisc.regs[38][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1255),
    .D(_01449_),
    .Q_N(_12519_),
    .Q(\top_ihp.oisc.regs[38][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1250),
    .D(_01450_),
    .Q_N(_12518_),
    .Q(\top_ihp.oisc.regs[38][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1383),
    .D(_01451_),
    .Q_N(_12517_),
    .Q(\top_ihp.oisc.regs[38][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1390),
    .D(_01452_),
    .Q_N(_12516_),
    .Q(\top_ihp.oisc.regs[38][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1390),
    .D(_01453_),
    .Q_N(_12515_),
    .Q(\top_ihp.oisc.regs[38][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1391),
    .D(_01454_),
    .Q_N(_12514_),
    .Q(\top_ihp.oisc.regs[38][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1269),
    .D(_01455_),
    .Q_N(_12513_),
    .Q(\top_ihp.oisc.regs[38][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1416),
    .D(_01456_),
    .Q_N(_12512_),
    .Q(\top_ihp.oisc.regs[38][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1392),
    .D(_01457_),
    .Q_N(_12511_),
    .Q(\top_ihp.oisc.regs[38][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1269),
    .D(_01458_),
    .Q_N(_12510_),
    .Q(\top_ihp.oisc.regs[38][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1349),
    .D(_01459_),
    .Q_N(_12509_),
    .Q(\top_ihp.oisc.regs[38][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1276),
    .D(_01460_),
    .Q_N(_12508_),
    .Q(\top_ihp.oisc.regs[38][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1267),
    .D(_01461_),
    .Q_N(_12507_),
    .Q(\top_ihp.oisc.regs[38][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1418),
    .D(_01462_),
    .Q_N(_12506_),
    .Q(\top_ihp.oisc.regs[38][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1418),
    .D(_01463_),
    .Q_N(_12505_),
    .Q(\top_ihp.oisc.regs[38][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1282),
    .D(_01464_),
    .Q_N(_12504_),
    .Q(\top_ihp.oisc.regs[38][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1282),
    .D(_01465_),
    .Q_N(_12503_),
    .Q(\top_ihp.oisc.regs[38][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1293),
    .D(_01466_),
    .Q_N(_12502_),
    .Q(\top_ihp.oisc.regs[38][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1426),
    .D(_01467_),
    .Q_N(_12501_),
    .Q(\top_ihp.oisc.regs[38][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1342),
    .D(_01468_),
    .Q_N(_12500_),
    .Q(\top_ihp.oisc.regs[38][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1424),
    .D(_01469_),
    .Q_N(_12499_),
    .Q(\top_ihp.oisc.regs[38][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1292),
    .D(_01470_),
    .Q_N(_12498_),
    .Q(\top_ihp.oisc.regs[38][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1407),
    .D(_01471_),
    .Q_N(_12497_),
    .Q(\top_ihp.oisc.regs[38][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1424),
    .D(_01472_),
    .Q_N(_12496_),
    .Q(\top_ihp.oisc.regs[38][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1351),
    .D(_01473_),
    .Q_N(_12495_),
    .Q(\top_ihp.oisc.regs[38][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1332),
    .D(_01474_),
    .Q_N(_12494_),
    .Q(\top_ihp.oisc.regs[38][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1416),
    .D(_01475_),
    .Q_N(_12493_),
    .Q(\top_ihp.oisc.regs[38][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1378),
    .D(_01476_),
    .Q_N(_12492_),
    .Q(\top_ihp.oisc.regs[39][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1302),
    .D(_01477_),
    .Q_N(_12491_),
    .Q(\top_ihp.oisc.regs[39][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1366),
    .D(_01478_),
    .Q_N(_12490_),
    .Q(\top_ihp.oisc.regs[39][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1301),
    .D(_01479_),
    .Q_N(_12489_),
    .Q(\top_ihp.oisc.regs[39][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1378),
    .D(_01480_),
    .Q_N(_12488_),
    .Q(\top_ihp.oisc.regs[39][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1261),
    .D(_01481_),
    .Q_N(_12487_),
    .Q(\top_ihp.oisc.regs[39][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1299),
    .D(_01482_),
    .Q_N(_12486_),
    .Q(\top_ihp.oisc.regs[39][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1378),
    .D(_01483_),
    .Q_N(_12485_),
    .Q(\top_ihp.oisc.regs[39][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1261),
    .D(_01484_),
    .Q_N(_12484_),
    .Q(\top_ihp.oisc.regs[39][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1321),
    .D(_01485_),
    .Q_N(_12483_),
    .Q(\top_ihp.oisc.regs[39][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1376),
    .D(_01486_),
    .Q_N(_12482_),
    .Q(\top_ihp.oisc.regs[39][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1267),
    .D(_01487_),
    .Q_N(_12481_),
    .Q(\top_ihp.oisc.regs[39][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1400),
    .D(_01488_),
    .Q_N(_12480_),
    .Q(\top_ihp.oisc.regs[39][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1256),
    .D(_01489_),
    .Q_N(_12479_),
    .Q(\top_ihp.oisc.regs[39][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1273),
    .D(_01490_),
    .Q_N(_12478_),
    .Q(\top_ihp.oisc.regs[39][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1349),
    .D(_01491_),
    .Q_N(_12477_),
    .Q(\top_ihp.oisc.regs[39][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1276),
    .D(_01492_),
    .Q_N(_12476_),
    .Q(\top_ihp.oisc.regs[39][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1309),
    .D(_01493_),
    .Q_N(_12475_),
    .Q(\top_ihp.oisc.regs[39][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1413),
    .D(_01494_),
    .Q_N(_12474_),
    .Q(\top_ihp.oisc.regs[39][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1413),
    .D(_01495_),
    .Q_N(_12473_),
    .Q(\top_ihp.oisc.regs[39][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1421),
    .D(_01496_),
    .Q_N(_12472_),
    .Q(\top_ihp.oisc.regs[39][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1282),
    .D(_01497_),
    .Q_N(_12471_),
    .Q(\top_ihp.oisc.regs[39][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1282),
    .D(_01498_),
    .Q_N(_12470_),
    .Q(\top_ihp.oisc.regs[39][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1408),
    .D(_01499_),
    .Q_N(_12469_),
    .Q(\top_ihp.oisc.regs[39][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1336),
    .D(_01500_),
    .Q_N(_12468_),
    .Q(\top_ihp.oisc.regs[39][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1343),
    .D(_01501_),
    .Q_N(_12467_),
    .Q(\top_ihp.oisc.regs[39][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1290),
    .D(_01502_),
    .Q_N(_12466_),
    .Q(\top_ihp.oisc.regs[39][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1407),
    .D(_01503_),
    .Q_N(_12465_),
    .Q(\top_ihp.oisc.regs[39][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1354),
    .D(_01504_),
    .Q_N(_12464_),
    .Q(\top_ihp.oisc.regs[39][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1286),
    .D(_01505_),
    .Q_N(_12463_),
    .Q(\top_ihp.oisc.regs[39][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1347),
    .D(_01506_),
    .Q_N(_12462_),
    .Q(\top_ihp.oisc.regs[39][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1277),
    .D(_01507_),
    .Q_N(_12461_),
    .Q(\top_ihp.oisc.regs[39][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1221),
    .D(_01508_),
    .Q_N(_12460_),
    .Q(\top_ihp.oisc.regs[3][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1221),
    .D(_01509_),
    .Q_N(_12459_),
    .Q(\top_ihp.oisc.regs[3][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1222),
    .D(_01510_),
    .Q_N(_12458_),
    .Q(\top_ihp.oisc.regs[3][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1221),
    .D(_01511_),
    .Q_N(_12457_),
    .Q(\top_ihp.oisc.regs[3][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1248),
    .D(_01512_),
    .Q_N(_12456_),
    .Q(\top_ihp.oisc.regs[3][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1222),
    .D(_01513_),
    .Q_N(_12455_),
    .Q(\top_ihp.oisc.regs[3][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1222),
    .D(_01514_),
    .Q_N(_12454_),
    .Q(\top_ihp.oisc.regs[3][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1221),
    .D(_01515_),
    .Q_N(_12453_),
    .Q(\top_ihp.oisc.regs[3][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1225),
    .D(_01516_),
    .Q_N(_12452_),
    .Q(\top_ihp.oisc.regs[3][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1225),
    .D(_01517_),
    .Q_N(_12451_),
    .Q(\top_ihp.oisc.regs[3][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1225),
    .D(_01518_),
    .Q_N(_12450_),
    .Q(\top_ihp.oisc.regs[3][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1225),
    .D(_01519_),
    .Q_N(_12449_),
    .Q(\top_ihp.oisc.regs[3][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1240),
    .D(_01520_),
    .Q_N(_12448_),
    .Q(\top_ihp.oisc.regs[3][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1226),
    .D(_01521_),
    .Q_N(_12447_),
    .Q(\top_ihp.oisc.regs[3][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1226),
    .D(_01522_),
    .Q_N(_12446_),
    .Q(\top_ihp.oisc.regs[3][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1226),
    .D(_01523_),
    .Q_N(_12445_),
    .Q(\top_ihp.oisc.regs[3][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1240),
    .D(_01524_),
    .Q_N(_12444_),
    .Q(\top_ihp.oisc.regs[3][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1225),
    .D(_01525_),
    .Q_N(_12443_),
    .Q(\top_ihp.oisc.regs[3][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1241),
    .D(_01526_),
    .Q_N(_12442_),
    .Q(\top_ihp.oisc.regs[3][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1241),
    .D(_01527_),
    .Q_N(_12441_),
    .Q(\top_ihp.oisc.regs[3][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1244),
    .D(_01528_),
    .Q_N(_12440_),
    .Q(\top_ihp.oisc.regs[3][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1244),
    .D(_01529_),
    .Q_N(_12439_),
    .Q(\top_ihp.oisc.regs[3][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1245),
    .D(_01530_),
    .Q_N(_12438_),
    .Q(\top_ihp.oisc.regs[3][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1200),
    .D(_01531_),
    .Q_N(_12437_),
    .Q(\top_ihp.oisc.regs[3][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1201),
    .D(_01532_),
    .Q_N(_12436_),
    .Q(\top_ihp.oisc.regs[3][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1200),
    .D(_01533_),
    .Q_N(_12435_),
    .Q(\top_ihp.oisc.regs[3][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1202),
    .D(_01534_),
    .Q_N(_12434_),
    .Q(\top_ihp.oisc.regs[3][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1244),
    .D(_01535_),
    .Q_N(_12433_),
    .Q(\top_ihp.oisc.regs[3][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1244),
    .D(_01536_),
    .Q_N(_12432_),
    .Q(\top_ihp.oisc.regs[3][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1244),
    .D(_01537_),
    .Q_N(_12431_),
    .Q(\top_ihp.oisc.regs[3][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1241),
    .D(_01538_),
    .Q_N(_12430_),
    .Q(\top_ihp.oisc.regs[3][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1226),
    .D(_01539_),
    .Q_N(_12429_),
    .Q(\top_ihp.oisc.regs[3][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1382),
    .D(_01540_),
    .Q_N(_12428_),
    .Q(\top_ihp.oisc.regs[40][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1383),
    .D(_01541_),
    .Q_N(_12427_),
    .Q(\top_ihp.oisc.regs[40][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1381),
    .D(_01542_),
    .Q_N(_12426_),
    .Q(\top_ihp.oisc.regs[40][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1259),
    .D(_01543_),
    .Q_N(_12425_),
    .Q(\top_ihp.oisc.regs[40][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1383),
    .D(_01544_),
    .Q_N(_12424_),
    .Q(\top_ihp.oisc.regs[40][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1248),
    .D(_01545_),
    .Q_N(_12423_),
    .Q(\top_ihp.oisc.regs[40][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1259),
    .D(_01546_),
    .Q_N(_12422_),
    .Q(\top_ihp.oisc.regs[40][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1382),
    .D(_01547_),
    .Q_N(_12421_),
    .Q(\top_ihp.oisc.regs[40][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1391),
    .D(_01548_),
    .Q_N(_12420_),
    .Q(\top_ihp.oisc.regs[40][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1384),
    .D(_01549_),
    .Q_N(_12419_),
    .Q(\top_ihp.oisc.regs[40][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1392),
    .D(_01550_),
    .Q_N(_12418_),
    .Q(\top_ihp.oisc.regs[40][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1268),
    .D(_01551_),
    .Q_N(_12417_),
    .Q(\top_ihp.oisc.regs[40][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1416),
    .D(_01552_),
    .Q_N(_12416_),
    .Q(\top_ihp.oisc.regs[40][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1392),
    .D(_01553_),
    .Q_N(_12415_),
    .Q(\top_ihp.oisc.regs[40][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1268),
    .D(_01554_),
    .Q_N(_12414_),
    .Q(\top_ihp.oisc.regs[40][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1349),
    .D(_01555_),
    .Q_N(_12413_),
    .Q(\top_ihp.oisc.regs[40][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1416),
    .D(_01556_),
    .Q_N(_12412_),
    .Q(\top_ihp.oisc.regs[40][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1255),
    .D(_01557_),
    .Q_N(_12411_),
    .Q(\top_ihp.oisc.regs[40][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1418),
    .D(_01558_),
    .Q_N(_12410_),
    .Q(\top_ihp.oisc.regs[40][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1418),
    .D(_01559_),
    .Q_N(_12409_),
    .Q(\top_ihp.oisc.regs[40][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1358),
    .D(_01560_),
    .Q_N(_12408_),
    .Q(\top_ihp.oisc.regs[40][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1424),
    .D(_01561_),
    .Q_N(_12407_),
    .Q(\top_ihp.oisc.regs[40][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1424),
    .D(_01562_),
    .Q_N(_12406_),
    .Q(\top_ihp.oisc.regs[40][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1424),
    .D(_01563_),
    .Q_N(_12405_),
    .Q(\top_ihp.oisc.regs[40][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1336),
    .D(_01564_),
    .Q_N(_12404_),
    .Q(\top_ihp.oisc.regs[40][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1425),
    .D(_01565_),
    .Q_N(_12403_),
    .Q(\top_ihp.oisc.regs[40][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1425),
    .D(_01566_),
    .Q_N(_12402_),
    .Q(\top_ihp.oisc.regs[40][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1423),
    .D(_01567_),
    .Q_N(_12401_),
    .Q(\top_ihp.oisc.regs[40][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1423),
    .D(_01568_),
    .Q_N(_12400_),
    .Q(\top_ihp.oisc.regs[40][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1347),
    .D(_01569_),
    .Q_N(_12399_),
    .Q(\top_ihp.oisc.regs[40][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1346),
    .D(_01570_),
    .Q_N(_12398_),
    .Q(\top_ihp.oisc.regs[40][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1346),
    .D(_01571_),
    .Q_N(_12397_),
    .Q(\top_ihp.oisc.regs[40][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1380),
    .D(_01572_),
    .Q_N(_12396_),
    .Q(\top_ihp.oisc.regs[41][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1384),
    .D(_01573_),
    .Q_N(_12395_),
    .Q(\top_ihp.oisc.regs[41][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1378),
    .D(_01574_),
    .Q_N(_12394_),
    .Q(\top_ihp.oisc.regs[41][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1260),
    .D(_01575_),
    .Q_N(_12393_),
    .Q(\top_ihp.oisc.regs[41][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1381),
    .D(_01576_),
    .Q_N(_12392_),
    .Q(\top_ihp.oisc.regs[41][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1250),
    .D(_01577_),
    .Q_N(_12391_),
    .Q(\top_ihp.oisc.regs[41][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1250),
    .D(_01578_),
    .Q_N(_12390_),
    .Q(\top_ihp.oisc.regs[41][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1381),
    .D(_01579_),
    .Q_N(_12389_),
    .Q(\top_ihp.oisc.regs[41][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1387),
    .D(_01580_),
    .Q_N(_12388_),
    .Q(\top_ihp.oisc.regs[41][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1384),
    .D(_01581_),
    .Q_N(_12387_),
    .Q(\top_ihp.oisc.regs[41][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1390),
    .D(_01582_),
    .Q_N(_12386_),
    .Q(\top_ihp.oisc.regs[41][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1255),
    .D(_01583_),
    .Q_N(_12385_),
    .Q(\top_ihp.oisc.regs[41][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1416),
    .D(_01584_),
    .Q_N(_12384_),
    .Q(\top_ihp.oisc.regs[41][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1392),
    .D(_01585_),
    .Q_N(_12383_),
    .Q(\top_ihp.oisc.regs[41][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1255),
    .D(_01586_),
    .Q_N(_12382_),
    .Q(\top_ihp.oisc.regs[41][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1388),
    .D(_01587_),
    .Q_N(_12381_),
    .Q(\top_ihp.oisc.regs[41][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1418),
    .D(_01588_),
    .Q_N(_12380_),
    .Q(\top_ihp.oisc.regs[41][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1255),
    .D(_01589_),
    .Q_N(_12379_),
    .Q(\top_ihp.oisc.regs[41][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1418),
    .D(_01590_),
    .Q_N(_12378_),
    .Q(\top_ihp.oisc.regs[41][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1418),
    .D(_01591_),
    .Q_N(_12377_),
    .Q(\top_ihp.oisc.regs[41][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1422),
    .D(_01592_),
    .Q_N(_12376_),
    .Q(\top_ihp.oisc.regs[41][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1358),
    .D(_01593_),
    .Q_N(_12375_),
    .Q(\top_ihp.oisc.regs[41][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1404),
    .D(_01594_),
    .Q_N(_12374_),
    .Q(\top_ihp.oisc.regs[41][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1405),
    .D(_01595_),
    .Q_N(_12373_),
    .Q(\top_ihp.oisc.regs[41][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1358),
    .D(_01596_),
    .Q_N(_12372_),
    .Q(\top_ihp.oisc.regs[41][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1360),
    .D(_01597_),
    .Q_N(_12371_),
    .Q(\top_ihp.oisc.regs[41][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1422),
    .D(_01598_),
    .Q_N(_12370_),
    .Q(\top_ihp.oisc.regs[41][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1291),
    .D(_01599_),
    .Q_N(_12369_),
    .Q(\top_ihp.oisc.regs[41][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1423),
    .D(_01600_),
    .Q_N(_12368_),
    .Q(\top_ihp.oisc.regs[41][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1414),
    .D(_01601_),
    .Q_N(_12367_),
    .Q(\top_ihp.oisc.regs[41][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1285),
    .D(_01602_),
    .Q_N(_12366_),
    .Q(\top_ihp.oisc.regs[41][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1412),
    .D(_01603_),
    .Q_N(_12365_),
    .Q(\top_ihp.oisc.regs[41][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1383),
    .D(_01604_),
    .Q_N(_12364_),
    .Q(\top_ihp.oisc.regs[42][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1383),
    .D(_01605_),
    .Q_N(_12363_),
    .Q(\top_ihp.oisc.regs[42][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1382),
    .D(_01606_),
    .Q_N(_12362_),
    .Q(\top_ihp.oisc.regs[42][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1261),
    .D(_01607_),
    .Q_N(_12361_),
    .Q(\top_ihp.oisc.regs[42][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1383),
    .D(_01608_),
    .Q_N(_12360_),
    .Q(\top_ihp.oisc.regs[42][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1260),
    .D(_01609_),
    .Q_N(_12359_),
    .Q(\top_ihp.oisc.regs[42][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1265),
    .D(_01610_),
    .Q_N(_12358_),
    .Q(\top_ihp.oisc.regs[42][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1382),
    .D(_01611_),
    .Q_N(_12357_),
    .Q(\top_ihp.oisc.regs[42][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1391),
    .D(_01612_),
    .Q_N(_12356_),
    .Q(\top_ihp.oisc.regs[42][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1391),
    .D(_01613_),
    .Q_N(_12355_),
    .Q(\top_ihp.oisc.regs[42][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1391),
    .D(_01614_),
    .Q_N(_12354_),
    .Q(\top_ihp.oisc.regs[42][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1305),
    .D(_01615_),
    .Q_N(_12353_),
    .Q(\top_ihp.oisc.regs[42][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1416),
    .D(_01616_),
    .Q_N(_12352_),
    .Q(\top_ihp.oisc.regs[42][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1392),
    .D(_01617_),
    .Q_N(_12351_),
    .Q(\top_ihp.oisc.regs[42][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1270),
    .D(_01618_),
    .Q_N(_12350_),
    .Q(\top_ihp.oisc.regs[42][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1346),
    .D(_01619_),
    .Q_N(_12349_),
    .Q(\top_ihp.oisc.regs[42][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1417),
    .D(_01620_),
    .Q_N(_12348_),
    .Q(\top_ihp.oisc.regs[42][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1304),
    .D(_01621_),
    .Q_N(_12347_),
    .Q(\top_ihp.oisc.regs[42][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1418),
    .D(_01622_),
    .Q_N(_12346_),
    .Q(\top_ihp.oisc.regs[42][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1419),
    .D(_01623_),
    .Q_N(_12345_),
    .Q(\top_ihp.oisc.regs[42][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1424),
    .D(_01624_),
    .Q_N(_12344_),
    .Q(\top_ihp.oisc.regs[42][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1425),
    .D(_01625_),
    .Q_N(_12343_),
    .Q(\top_ihp.oisc.regs[42][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1424),
    .D(_01626_),
    .Q_N(_12342_),
    .Q(\top_ihp.oisc.regs[42][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1425),
    .D(_01627_),
    .Q_N(_12341_),
    .Q(\top_ihp.oisc.regs[42][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1290),
    .D(_01628_),
    .Q_N(_12340_),
    .Q(\top_ihp.oisc.regs[42][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1426),
    .D(_01629_),
    .Q_N(_12339_),
    .Q(\top_ihp.oisc.regs[42][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1425),
    .D(_01630_),
    .Q_N(_12338_),
    .Q(\top_ihp.oisc.regs[42][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1407),
    .D(_01631_),
    .Q_N(_12337_),
    .Q(\top_ihp.oisc.regs[42][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1351),
    .D(_01632_),
    .Q_N(_12336_),
    .Q(\top_ihp.oisc.regs[42][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1333),
    .D(_01633_),
    .Q_N(_12335_),
    .Q(\top_ihp.oisc.regs[42][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1347),
    .D(_01634_),
    .Q_N(_12334_),
    .Q(\top_ihp.oisc.regs[42][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1417),
    .D(_01635_),
    .Q_N(_12333_),
    .Q(\top_ihp.oisc.regs[42][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1313),
    .D(_01636_),
    .Q_N(_12332_),
    .Q(\top_ihp.oisc.regs[43][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1368),
    .D(_01637_),
    .Q_N(_12331_),
    .Q(\top_ihp.oisc.regs[43][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1313),
    .D(_01638_),
    .Q_N(_12330_),
    .Q(\top_ihp.oisc.regs[43][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1263),
    .D(_01639_),
    .Q_N(_12329_),
    .Q(\top_ihp.oisc.regs[43][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1380),
    .D(_01640_),
    .Q_N(_12328_),
    .Q(\top_ihp.oisc.regs[43][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1263),
    .D(_01641_),
    .Q_N(_12327_),
    .Q(\top_ihp.oisc.regs[43][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1297),
    .D(_01642_),
    .Q_N(_12326_),
    .Q(\top_ihp.oisc.regs[43][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1380),
    .D(_01643_),
    .Q_N(_12325_),
    .Q(\top_ihp.oisc.regs[43][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1390),
    .D(_01644_),
    .Q_N(_12324_),
    .Q(\top_ihp.oisc.regs[43][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1384),
    .D(_01645_),
    .Q_N(_12323_),
    .Q(\top_ihp.oisc.regs[43][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1391),
    .D(_01646_),
    .Q_N(_12322_),
    .Q(\top_ihp.oisc.regs[43][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1387),
    .D(_01647_),
    .Q_N(_12321_),
    .Q(\top_ihp.oisc.regs[43][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1393),
    .D(_01648_),
    .Q_N(_12320_),
    .Q(\top_ihp.oisc.regs[43][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1393),
    .D(_01649_),
    .Q_N(_12319_),
    .Q(\top_ihp.oisc.regs[43][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1309),
    .D(_01650_),
    .Q_N(_12318_),
    .Q(\top_ihp.oisc.regs[43][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1389),
    .D(_01651_),
    .Q_N(_12317_),
    .Q(\top_ihp.oisc.regs[43][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1417),
    .D(_01652_),
    .Q_N(_12316_),
    .Q(\top_ihp.oisc.regs[43][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1307),
    .D(_01653_),
    .Q_N(_12315_),
    .Q(\top_ihp.oisc.regs[43][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1419),
    .D(_01654_),
    .Q_N(_12314_),
    .Q(\top_ihp.oisc.regs[43][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1419),
    .D(_01655_),
    .Q_N(_12313_),
    .Q(\top_ihp.oisc.regs[43][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1424),
    .D(_01656_),
    .Q_N(_12312_),
    .Q(\top_ihp.oisc.regs[43][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1426),
    .D(_01657_),
    .Q_N(_12311_),
    .Q(\top_ihp.oisc.regs[43][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1426),
    .D(_01658_),
    .Q_N(_12310_),
    .Q(\top_ihp.oisc.regs[43][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1426),
    .D(_01659_),
    .Q_N(_12309_),
    .Q(\top_ihp.oisc.regs[43][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1291),
    .D(_01660_),
    .Q_N(_12308_),
    .Q(\top_ihp.oisc.regs[43][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1426),
    .D(_01661_),
    .Q_N(_12307_),
    .Q(\top_ihp.oisc.regs[43][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1341),
    .D(_01662_),
    .Q_N(_12306_),
    .Q(\top_ihp.oisc.regs[43][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1402),
    .D(_01663_),
    .Q_N(_12305_),
    .Q(\top_ihp.oisc.regs[43][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1291),
    .D(_01664_),
    .Q_N(_12304_),
    .Q(\top_ihp.oisc.regs[43][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1414),
    .D(_01665_),
    .Q_N(_12303_),
    .Q(\top_ihp.oisc.regs[43][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1333),
    .D(_01666_),
    .Q_N(_12302_),
    .Q(\top_ihp.oisc.regs[43][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1416),
    .D(_01667_),
    .Q_N(_12301_),
    .Q(\top_ihp.oisc.regs[43][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1384),
    .D(_01668_),
    .Q_N(_12300_),
    .Q(\top_ihp.oisc.regs[44][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1384),
    .D(_01669_),
    .Q_N(_12299_),
    .Q(\top_ihp.oisc.regs[44][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1381),
    .D(_01670_),
    .Q_N(_12298_),
    .Q(\top_ihp.oisc.regs[44][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1261),
    .D(_01671_),
    .Q_N(_12297_),
    .Q(\top_ihp.oisc.regs[44][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1381),
    .D(_01672_),
    .Q_N(_12296_),
    .Q(\top_ihp.oisc.regs[44][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1255),
    .D(_01673_),
    .Q_N(_12295_),
    .Q(\top_ihp.oisc.regs[44][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1265),
    .D(_01674_),
    .Q_N(_12294_),
    .Q(\top_ihp.oisc.regs[44][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1384),
    .D(_01675_),
    .Q_N(_12293_),
    .Q(\top_ihp.oisc.regs[44][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1390),
    .D(_01676_),
    .Q_N(_12292_),
    .Q(\top_ihp.oisc.regs[44][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1390),
    .D(_01677_),
    .Q_N(_12291_),
    .Q(\top_ihp.oisc.regs[44][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1392),
    .D(_01678_),
    .Q_N(_12290_),
    .Q(\top_ihp.oisc.regs[44][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1269),
    .D(_01679_),
    .Q_N(_12289_),
    .Q(\top_ihp.oisc.regs[44][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1416),
    .D(_01680_),
    .Q_N(_12288_),
    .Q(\top_ihp.oisc.regs[44][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1392),
    .D(_01681_),
    .Q_N(_12287_),
    .Q(\top_ihp.oisc.regs[44][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1269),
    .D(_01682_),
    .Q_N(_12286_),
    .Q(\top_ihp.oisc.regs[44][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1411),
    .D(_01683_),
    .Q_N(_12285_),
    .Q(\top_ihp.oisc.regs[44][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1417),
    .D(_01684_),
    .Q_N(_12284_),
    .Q(\top_ihp.oisc.regs[44][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1269),
    .D(_01685_),
    .Q_N(_12283_),
    .Q(\top_ihp.oisc.regs[44][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1419),
    .D(_01686_),
    .Q_N(_12282_),
    .Q(\top_ihp.oisc.regs[44][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1419),
    .D(_01687_),
    .Q_N(_12281_),
    .Q(\top_ihp.oisc.regs[44][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1423),
    .D(_01688_),
    .Q_N(_12280_),
    .Q(\top_ihp.oisc.regs[44][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1426),
    .D(_01689_),
    .Q_N(_12279_),
    .Q(\top_ihp.oisc.regs[44][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1426),
    .D(_01690_),
    .Q_N(_12278_),
    .Q(\top_ihp.oisc.regs[44][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1427),
    .D(_01691_),
    .Q_N(_12277_),
    .Q(\top_ihp.oisc.regs[44][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1292),
    .D(_01692_),
    .Q_N(_12276_),
    .Q(\top_ihp.oisc.regs[44][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1336),
    .D(_01693_),
    .Q_N(_12275_),
    .Q(\top_ihp.oisc.regs[44][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1337),
    .D(_01694_),
    .Q_N(_12274_),
    .Q(\top_ihp.oisc.regs[44][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1407),
    .D(_01695_),
    .Q_N(_12273_),
    .Q(\top_ihp.oisc.regs[44][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1337),
    .D(_01696_),
    .Q_N(_12272_),
    .Q(\top_ihp.oisc.regs[44][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1347),
    .D(_01697_),
    .Q_N(_12271_),
    .Q(\top_ihp.oisc.regs[44][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1329),
    .D(_01698_),
    .Q_N(_12270_),
    .Q(\top_ihp.oisc.regs[44][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1332),
    .D(_01699_),
    .Q_N(_12269_),
    .Q(\top_ihp.oisc.regs[44][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1379),
    .D(_01700_),
    .Q_N(_12268_),
    .Q(\top_ihp.oisc.regs[45][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1379),
    .D(_01701_),
    .Q_N(_12267_),
    .Q(\top_ihp.oisc.regs[45][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1380),
    .D(_01702_),
    .Q_N(_12266_),
    .Q(\top_ihp.oisc.regs[45][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1260),
    .D(_01703_),
    .Q_N(_12265_),
    .Q(\top_ihp.oisc.regs[45][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1379),
    .D(_01704_),
    .Q_N(_12264_),
    .Q(\top_ihp.oisc.regs[45][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1260),
    .D(_01705_),
    .Q_N(_12263_),
    .Q(\top_ihp.oisc.regs[45][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1260),
    .D(_01706_),
    .Q_N(_12262_),
    .Q(\top_ihp.oisc.regs[45][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1379),
    .D(_01707_),
    .Q_N(_12261_),
    .Q(\top_ihp.oisc.regs[45][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1386),
    .D(_01708_),
    .Q_N(_12260_),
    .Q(\top_ihp.oisc.regs[45][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1386),
    .D(_01709_),
    .Q_N(_12259_),
    .Q(\top_ihp.oisc.regs[45][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1387),
    .D(_01710_),
    .Q_N(_12258_),
    .Q(\top_ihp.oisc.regs[45][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1267),
    .D(_01711_),
    .Q_N(_12257_),
    .Q(\top_ihp.oisc.regs[45][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1412),
    .D(_01712_),
    .Q_N(_12256_),
    .Q(\top_ihp.oisc.regs[45][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1388),
    .D(_01713_),
    .Q_N(_12255_),
    .Q(\top_ihp.oisc.regs[45][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1273),
    .D(_01714_),
    .Q_N(_12254_),
    .Q(\top_ihp.oisc.regs[45][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1411),
    .D(_01715_),
    .Q_N(_12253_),
    .Q(\top_ihp.oisc.regs[45][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1350),
    .D(_01716_),
    .Q_N(_12252_),
    .Q(\top_ihp.oisc.regs[45][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1268),
    .D(_01717_),
    .Q_N(_12251_),
    .Q(\top_ihp.oisc.regs[45][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1275),
    .D(_01718_),
    .Q_N(_12250_),
    .Q(\top_ihp.oisc.regs[45][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1399),
    .D(_01719_),
    .Q_N(_12249_),
    .Q(\top_ihp.oisc.regs[45][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1289),
    .D(_01720_),
    .Q_N(_12248_),
    .Q(\top_ihp.oisc.regs[45][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1279),
    .D(_01721_),
    .Q_N(_12247_),
    .Q(\top_ihp.oisc.regs[45][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1279),
    .D(_01722_),
    .Q_N(_12246_),
    .Q(\top_ihp.oisc.regs[45][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1423),
    .D(_01723_),
    .Q_N(_12245_),
    .Q(\top_ihp.oisc.regs[45][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1354),
    .D(_01724_),
    .Q_N(_12244_),
    .Q(\top_ihp.oisc.regs[45][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1423),
    .D(_01725_),
    .Q_N(_12243_),
    .Q(\top_ihp.oisc.regs[45][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1338),
    .D(_01726_),
    .Q_N(_12242_),
    .Q(\top_ihp.oisc.regs[45][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1291),
    .D(_01727_),
    .Q_N(_12241_),
    .Q(\top_ihp.oisc.regs[45][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1286),
    .D(_01728_),
    .Q_N(_12240_),
    .Q(\top_ihp.oisc.regs[45][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1413),
    .D(_01729_),
    .Q_N(_12239_),
    .Q(\top_ihp.oisc.regs[45][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1346),
    .D(_01730_),
    .Q_N(_12238_),
    .Q(\top_ihp.oisc.regs[45][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1285),
    .D(_01731_),
    .Q_N(_12237_),
    .Q(\top_ihp.oisc.regs[45][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1319),
    .D(_01732_),
    .Q_N(_12236_),
    .Q(\top_ihp.oisc.regs[46][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1303),
    .D(_01733_),
    .Q_N(_12235_),
    .Q(\top_ihp.oisc.regs[46][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1316),
    .D(_01734_),
    .Q_N(_12234_),
    .Q(\top_ihp.oisc.regs[46][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1261),
    .D(_01735_),
    .Q_N(_12233_),
    .Q(\top_ihp.oisc.regs[46][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1317),
    .D(_01736_),
    .Q_N(_12232_),
    .Q(\top_ihp.oisc.regs[46][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1250),
    .D(_01737_),
    .Q_N(_12231_),
    .Q(\top_ihp.oisc.regs[46][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1250),
    .D(_01738_),
    .Q_N(_12230_),
    .Q(\top_ihp.oisc.regs[46][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1368),
    .D(_01739_),
    .Q_N(_12229_),
    .Q(\top_ihp.oisc.regs[46][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1375),
    .D(_01740_),
    .Q_N(_12228_),
    .Q(\top_ihp.oisc.regs[46][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1319),
    .D(_01741_),
    .Q_N(_12227_),
    .Q(\top_ihp.oisc.regs[46][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1376),
    .D(_01742_),
    .Q_N(_12226_),
    .Q(\top_ihp.oisc.regs[46][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1269),
    .D(_01743_),
    .Q_N(_12225_),
    .Q(\top_ihp.oisc.regs[46][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1376),
    .D(_01744_),
    .Q_N(_12224_),
    .Q(\top_ihp.oisc.regs[46][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1372),
    .D(_01745_),
    .Q_N(_12223_),
    .Q(\top_ihp.oisc.regs[46][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1270),
    .D(_01746_),
    .Q_N(_12222_),
    .Q(\top_ihp.oisc.regs[46][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1376),
    .D(_01747_),
    .Q_N(_12221_),
    .Q(\top_ihp.oisc.regs[46][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1395),
    .D(_01748_),
    .Q_N(_12220_),
    .Q(\top_ihp.oisc.regs[46][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1322),
    .D(_01749_),
    .Q_N(_12219_),
    .Q(\top_ihp.oisc.regs[46][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1396),
    .D(_01750_),
    .Q_N(_12218_),
    .Q(\top_ihp.oisc.regs[46][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1284),
    .D(_01751_),
    .Q_N(_12217_),
    .Q(\top_ihp.oisc.regs[46][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1422),
    .D(_01752_),
    .Q_N(_12216_),
    .Q(\top_ihp.oisc.regs[46][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1288),
    .D(_01753_),
    .Q_N(_12215_),
    .Q(\top_ihp.oisc.regs[46][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1408),
    .D(_01754_),
    .Q_N(_12214_),
    .Q(\top_ihp.oisc.regs[46][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1422),
    .D(_01755_),
    .Q_N(_12213_),
    .Q(\top_ihp.oisc.regs[46][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1338),
    .D(_01756_),
    .Q_N(_12212_),
    .Q(\top_ihp.oisc.regs[46][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1291),
    .D(_01757_),
    .Q_N(_12211_),
    .Q(\top_ihp.oisc.regs[46][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1290),
    .D(_01758_),
    .Q_N(_12210_),
    .Q(\top_ihp.oisc.regs[46][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1402),
    .D(_01759_),
    .Q_N(_12209_),
    .Q(\top_ihp.oisc.regs[46][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1286),
    .D(_01760_),
    .Q_N(_12208_),
    .Q(\top_ihp.oisc.regs[46][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1281),
    .D(_01761_),
    .Q_N(_12207_),
    .Q(\top_ihp.oisc.regs[46][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1285),
    .D(_01762_),
    .Q_N(_12206_),
    .Q(\top_ihp.oisc.regs[46][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1309),
    .D(_01763_),
    .Q_N(_12205_),
    .Q(\top_ihp.oisc.regs[46][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1368),
    .D(_01764_),
    .Q_N(_12204_),
    .Q(\top_ihp.oisc.regs[47][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1368),
    .D(_01765_),
    .Q_N(_12203_),
    .Q(\top_ihp.oisc.regs[47][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1378),
    .D(_01766_),
    .Q_N(_12202_),
    .Q(\top_ihp.oisc.regs[47][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1262),
    .D(_01767_),
    .Q_N(_12201_),
    .Q(\top_ihp.oisc.regs[47][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1378),
    .D(_01768_),
    .Q_N(_12200_),
    .Q(\top_ihp.oisc.regs[47][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1263),
    .D(_01769_),
    .Q_N(_12199_),
    .Q(\top_ihp.oisc.regs[47][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1262),
    .D(_01770_),
    .Q_N(_12198_),
    .Q(\top_ihp.oisc.regs[47][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1379),
    .D(_01771_),
    .Q_N(_12197_),
    .Q(\top_ihp.oisc.regs[47][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1379),
    .D(_01772_),
    .Q_N(_12196_),
    .Q(\top_ihp.oisc.regs[47][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1375),
    .D(_01773_),
    .Q_N(_12195_),
    .Q(\top_ihp.oisc.regs[47][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1386),
    .D(_01774_),
    .Q_N(_12194_),
    .Q(\top_ihp.oisc.regs[47][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1269),
    .D(_01775_),
    .Q_N(_12193_),
    .Q(\top_ihp.oisc.regs[47][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1376),
    .D(_01776_),
    .Q_N(_12192_),
    .Q(\top_ihp.oisc.regs[47][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1372),
    .D(_01777_),
    .Q_N(_12191_),
    .Q(\top_ihp.oisc.regs[47][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1270),
    .D(_01778_),
    .Q_N(_12190_),
    .Q(\top_ihp.oisc.regs[47][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1350),
    .D(_01779_),
    .Q_N(_12189_),
    .Q(\top_ihp.oisc.regs[47][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1350),
    .D(_01780_),
    .Q_N(_12188_),
    .Q(\top_ihp.oisc.regs[47][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1270),
    .D(_01781_),
    .Q_N(_12187_),
    .Q(\top_ihp.oisc.regs[47][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1413),
    .D(_01782_),
    .Q_N(_12186_),
    .Q(\top_ihp.oisc.regs[47][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1351),
    .D(_01783_),
    .Q_N(_12185_),
    .Q(\top_ihp.oisc.regs[47][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1421),
    .D(_01784_),
    .Q_N(_12184_),
    .Q(\top_ihp.oisc.regs[47][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1358),
    .D(_01785_),
    .Q_N(_12183_),
    .Q(\top_ihp.oisc.regs[47][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1407),
    .D(_01786_),
    .Q_N(_12182_),
    .Q(\top_ihp.oisc.regs[47][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1407),
    .D(_01787_),
    .Q_N(_12181_),
    .Q(\top_ihp.oisc.regs[47][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1354),
    .D(_01788_),
    .Q_N(_12180_),
    .Q(\top_ihp.oisc.regs[47][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1337),
    .D(_01789_),
    .Q_N(_12179_),
    .Q(\top_ihp.oisc.regs[47][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1336),
    .D(_01790_),
    .Q_N(_12178_),
    .Q(\top_ihp.oisc.regs[47][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1410),
    .D(_01791_),
    .Q_N(_12177_),
    .Q(\top_ihp.oisc.regs[47][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1399),
    .D(_01792_),
    .Q_N(_12176_),
    .Q(\top_ihp.oisc.regs[47][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1399),
    .D(_01793_),
    .Q_N(_12175_),
    .Q(\top_ihp.oisc.regs[47][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1332),
    .D(_01794_),
    .Q_N(_12174_),
    .Q(\top_ihp.oisc.regs[47][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1400),
    .D(_01795_),
    .Q_N(_12173_),
    .Q(\top_ihp.oisc.regs[47][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1319),
    .D(_01796_),
    .Q_N(_12172_),
    .Q(\top_ihp.oisc.regs[48][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1319),
    .D(_01797_),
    .Q_N(_12171_),
    .Q(\top_ihp.oisc.regs[48][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1365),
    .D(_01798_),
    .Q_N(_12170_),
    .Q(\top_ihp.oisc.regs[48][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1299),
    .D(_01799_),
    .Q_N(_12169_),
    .Q(\top_ihp.oisc.regs[48][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1318),
    .D(_01800_),
    .Q_N(_12168_),
    .Q(\top_ihp.oisc.regs[48][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1251),
    .D(_01801_),
    .Q_N(_12167_),
    .Q(\top_ihp.oisc.regs[48][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1250),
    .D(_01802_),
    .Q_N(_12166_),
    .Q(\top_ihp.oisc.regs[48][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1252),
    .D(_01803_),
    .Q_N(_12165_),
    .Q(\top_ihp.oisc.regs[48][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1307),
    .D(_01804_),
    .Q_N(_12164_),
    .Q(\top_ihp.oisc.regs[48][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1371),
    .D(_01805_),
    .Q_N(_12163_),
    .Q(\top_ihp.oisc.regs[48][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1325),
    .D(_01806_),
    .Q_N(_12162_),
    .Q(\top_ihp.oisc.regs[48][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1372),
    .D(_01807_),
    .Q_N(_12161_),
    .Q(\top_ihp.oisc.regs[48][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1395),
    .D(_01808_),
    .Q_N(_12160_),
    .Q(\top_ihp.oisc.regs[48][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1305),
    .D(_01809_),
    .Q_N(_12159_),
    .Q(\top_ihp.oisc.regs[48][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1272),
    .D(_01810_),
    .Q_N(_12158_),
    .Q(\top_ihp.oisc.regs[48][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1325),
    .D(_01811_),
    .Q_N(_12157_),
    .Q(\top_ihp.oisc.regs[48][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1395),
    .D(_01812_),
    .Q_N(_12156_),
    .Q(\top_ihp.oisc.regs[48][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1305),
    .D(_01813_),
    .Q_N(_12155_),
    .Q(\top_ihp.oisc.regs[48][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1277),
    .D(_01814_),
    .Q_N(_12154_),
    .Q(\top_ihp.oisc.regs[48][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1277),
    .D(_01815_),
    .Q_N(_12153_),
    .Q(\top_ihp.oisc.regs[48][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1281),
    .D(_01816_),
    .Q_N(_12152_),
    .Q(\top_ihp.oisc.regs[48][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1359),
    .D(_01817_),
    .Q_N(_12151_),
    .Q(\top_ihp.oisc.regs[48][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1359),
    .D(_01818_),
    .Q_N(_12150_),
    .Q(\top_ihp.oisc.regs[48][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1358),
    .D(_01819_),
    .Q_N(_12149_),
    .Q(\top_ihp.oisc.regs[48][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1288),
    .D(_01820_),
    .Q_N(_12148_),
    .Q(\top_ihp.oisc.regs[48][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1278),
    .D(_01821_),
    .Q_N(_12147_),
    .Q(\top_ihp.oisc.regs[48][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1292),
    .D(_01822_),
    .Q_N(_12146_),
    .Q(\top_ihp.oisc.regs[48][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1292),
    .D(_01823_),
    .Q_N(_12145_),
    .Q(\top_ihp.oisc.regs[48][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1358),
    .D(_01824_),
    .Q_N(_12144_),
    .Q(\top_ihp.oisc.regs[48][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1334),
    .D(_01825_),
    .Q_N(_12143_),
    .Q(\top_ihp.oisc.regs[48][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1285),
    .D(_01826_),
    .Q_N(_12142_),
    .Q(\top_ihp.oisc.regs[48][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1285),
    .D(_01827_),
    .Q_N(_12141_),
    .Q(\top_ihp.oisc.regs[48][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1319),
    .D(_01828_),
    .Q_N(_12140_),
    .Q(\top_ihp.oisc.regs[49][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1364),
    .D(_01829_),
    .Q_N(_12139_),
    .Q(\top_ihp.oisc.regs[49][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1365),
    .D(_01830_),
    .Q_N(_12138_),
    .Q(\top_ihp.oisc.regs[49][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1264),
    .D(_01831_),
    .Q_N(_12137_),
    .Q(\top_ihp.oisc.regs[49][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1318),
    .D(_01832_),
    .Q_N(_12136_),
    .Q(\top_ihp.oisc.regs[49][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1263),
    .D(_01833_),
    .Q_N(_12135_),
    .Q(\top_ihp.oisc.regs[49][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1266),
    .D(_01834_),
    .Q_N(_12134_),
    .Q(\top_ihp.oisc.regs[49][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1365),
    .D(_01835_),
    .Q_N(_12133_),
    .Q(\top_ihp.oisc.regs[49][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1307),
    .D(_01836_),
    .Q_N(_12132_),
    .Q(\top_ihp.oisc.regs[49][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1321),
    .D(_01837_),
    .Q_N(_12131_),
    .Q(\top_ihp.oisc.regs[49][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1305),
    .D(_01838_),
    .Q_N(_12130_),
    .Q(\top_ihp.oisc.regs[49][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1270),
    .D(_01839_),
    .Q_N(_12129_),
    .Q(\top_ihp.oisc.regs[49][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1376),
    .D(_01840_),
    .Q_N(_12128_),
    .Q(\top_ihp.oisc.regs[49][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1271),
    .D(_01841_),
    .Q_N(_12127_),
    .Q(\top_ihp.oisc.regs[49][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1271),
    .D(_01842_),
    .Q_N(_12126_),
    .Q(\top_ihp.oisc.regs[49][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1400),
    .D(_01843_),
    .Q_N(_12125_),
    .Q(\top_ihp.oisc.regs[49][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1400),
    .D(_01844_),
    .Q_N(_12124_),
    .Q(\top_ihp.oisc.regs[49][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1322),
    .D(_01845_),
    .Q_N(_12123_),
    .Q(\top_ihp.oisc.regs[49][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1399),
    .D(_01846_),
    .Q_N(_12122_),
    .Q(\top_ihp.oisc.regs[49][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1399),
    .D(_01847_),
    .Q_N(_12121_),
    .Q(\top_ihp.oisc.regs[49][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1360),
    .D(_01848_),
    .Q_N(_12120_),
    .Q(\top_ihp.oisc.regs[49][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1359),
    .D(_01849_),
    .Q_N(_12119_),
    .Q(\top_ihp.oisc.regs[49][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1356),
    .D(_01850_),
    .Q_N(_12118_),
    .Q(\top_ihp.oisc.regs[49][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1358),
    .D(_01851_),
    .Q_N(_12117_),
    .Q(\top_ihp.oisc.regs[49][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1355),
    .D(_01852_),
    .Q_N(_12116_),
    .Q(\top_ihp.oisc.regs[49][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1342),
    .D(_01853_),
    .Q_N(_12115_),
    .Q(\top_ihp.oisc.regs[49][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1342),
    .D(_01854_),
    .Q_N(_12114_),
    .Q(\top_ihp.oisc.regs[49][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1338),
    .D(_01855_),
    .Q_N(_12113_),
    .Q(\top_ihp.oisc.regs[49][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1330),
    .D(_01856_),
    .Q_N(_12112_),
    .Q(\top_ihp.oisc.regs[49][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1333),
    .D(_01857_),
    .Q_N(_12111_),
    .Q(\top_ihp.oisc.regs[49][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1332),
    .D(_01858_),
    .Q_N(_12110_),
    .Q(\top_ihp.oisc.regs[49][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1332),
    .D(_01859_),
    .Q_N(_12109_),
    .Q(\top_ihp.oisc.regs[49][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1221),
    .D(_01860_),
    .Q_N(_12108_),
    .Q(\top_ihp.oisc.regs[4][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1249),
    .D(_01861_),
    .Q_N(_12107_),
    .Q(\top_ihp.oisc.regs[4][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1249),
    .D(_01862_),
    .Q_N(_12106_),
    .Q(\top_ihp.oisc.regs[4][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1222),
    .D(_01863_),
    .Q_N(_12105_),
    .Q(\top_ihp.oisc.regs[4][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1248),
    .D(_01864_),
    .Q_N(_12104_),
    .Q(\top_ihp.oisc.regs[4][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1222),
    .D(_01865_),
    .Q_N(_12103_),
    .Q(\top_ihp.oisc.regs[4][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1248),
    .D(_01866_),
    .Q_N(_12102_),
    .Q(\top_ihp.oisc.regs[4][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1249),
    .D(_01867_),
    .Q_N(_12101_),
    .Q(\top_ihp.oisc.regs[4][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1249),
    .D(_01868_),
    .Q_N(_12100_),
    .Q(\top_ihp.oisc.regs[4][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1253),
    .D(_01869_),
    .Q_N(_12099_),
    .Q(\top_ihp.oisc.regs[4][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1253),
    .D(_01870_),
    .Q_N(_12098_),
    .Q(\top_ihp.oisc.regs[4][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1226),
    .D(_01871_),
    .Q_N(_12097_),
    .Q(\top_ihp.oisc.regs[4][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1240),
    .D(_01872_),
    .Q_N(_12096_),
    .Q(\top_ihp.oisc.regs[4][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1275),
    .D(_01873_),
    .Q_N(_12095_),
    .Q(\top_ihp.oisc.regs[4][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1227),
    .D(_01874_),
    .Q_N(_12094_),
    .Q(\top_ihp.oisc.regs[4][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1254),
    .D(_01875_),
    .Q_N(_12093_),
    .Q(\top_ihp.oisc.regs[4][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1275),
    .D(_01876_),
    .Q_N(_12092_),
    .Q(\top_ihp.oisc.regs[4][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1254),
    .D(_01877_),
    .Q_N(_12091_),
    .Q(\top_ihp.oisc.regs[4][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1241),
    .D(_01878_),
    .Q_N(_12090_),
    .Q(\top_ihp.oisc.regs[4][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1241),
    .D(_01879_),
    .Q_N(_12089_),
    .Q(\top_ihp.oisc.regs[4][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1245),
    .D(_01880_),
    .Q_N(_12088_),
    .Q(\top_ihp.oisc.regs[4][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1245),
    .D(_01881_),
    .Q_N(_12087_),
    .Q(\top_ihp.oisc.regs[4][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1245),
    .D(_01882_),
    .Q_N(_12086_),
    .Q(\top_ihp.oisc.regs[4][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1201),
    .D(_01883_),
    .Q_N(_12085_),
    .Q(\top_ihp.oisc.regs[4][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1202),
    .D(_01884_),
    .Q_N(_12084_),
    .Q(\top_ihp.oisc.regs[4][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1196),
    .D(_01885_),
    .Q_N(_12083_),
    .Q(\top_ihp.oisc.regs[4][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1202),
    .D(_01886_),
    .Q_N(_12082_),
    .Q(\top_ihp.oisc.regs[4][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1245),
    .D(_01887_),
    .Q_N(_12081_),
    .Q(\top_ihp.oisc.regs[4][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1244),
    .D(_01888_),
    .Q_N(_12080_),
    .Q(\top_ihp.oisc.regs[4][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1244),
    .D(_01889_),
    .Q_N(_12079_),
    .Q(\top_ihp.oisc.regs[4][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1275),
    .D(_01890_),
    .Q_N(_12078_),
    .Q(\top_ihp.oisc.regs[4][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1254),
    .D(_01891_),
    .Q_N(_12077_),
    .Q(\top_ihp.oisc.regs[4][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1315),
    .D(_01892_),
    .Q_N(_12076_),
    .Q(\top_ihp.oisc.regs[50][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1379),
    .D(_01893_),
    .Q_N(_12075_),
    .Q(\top_ihp.oisc.regs[50][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1378),
    .D(_01894_),
    .Q_N(_12074_),
    .Q(\top_ihp.oisc.regs[50][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1302),
    .D(_01895_),
    .Q_N(_12073_),
    .Q(\top_ihp.oisc.regs[50][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1378),
    .D(_01896_),
    .Q_N(_12072_),
    .Q(\top_ihp.oisc.regs[50][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1250),
    .D(_01897_),
    .Q_N(_12071_),
    .Q(\top_ihp.oisc.regs[50][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1251),
    .D(_01898_),
    .Q_N(_12070_),
    .Q(\top_ihp.oisc.regs[50][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1252),
    .D(_01899_),
    .Q_N(_12069_),
    .Q(\top_ihp.oisc.regs[50][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1386),
    .D(_01900_),
    .Q_N(_12068_),
    .Q(\top_ihp.oisc.regs[50][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1375),
    .D(_01901_),
    .Q_N(_12067_),
    .Q(\top_ihp.oisc.regs[50][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1388),
    .D(_01902_),
    .Q_N(_12066_),
    .Q(\top_ihp.oisc.regs[50][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1308),
    .D(_01903_),
    .Q_N(_12065_),
    .Q(\top_ihp.oisc.regs[50][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1412),
    .D(_01904_),
    .Q_N(_12064_),
    .Q(\top_ihp.oisc.regs[50][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1388),
    .D(_01905_),
    .Q_N(_12063_),
    .Q(\top_ihp.oisc.regs[50][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1322),
    .D(_01906_),
    .Q_N(_12062_),
    .Q(\top_ihp.oisc.regs[50][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1388),
    .D(_01907_),
    .Q_N(_12061_),
    .Q(\top_ihp.oisc.regs[50][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1395),
    .D(_01908_),
    .Q_N(_12060_),
    .Q(\top_ihp.oisc.regs[50][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1321),
    .D(_01909_),
    .Q_N(_12059_),
    .Q(\top_ihp.oisc.regs[50][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1413),
    .D(_01910_),
    .Q_N(_12058_),
    .Q(\top_ihp.oisc.regs[50][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1399),
    .D(_01911_),
    .Q_N(_12057_),
    .Q(\top_ihp.oisc.regs[50][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1421),
    .D(_01912_),
    .Q_N(_12056_),
    .Q(\top_ihp.oisc.regs[50][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1289),
    .D(_01913_),
    .Q_N(_12055_),
    .Q(\top_ihp.oisc.regs[50][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1408),
    .D(_01914_),
    .Q_N(_12054_),
    .Q(\top_ihp.oisc.regs[50][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1339),
    .D(_01915_),
    .Q_N(_12053_),
    .Q(\top_ihp.oisc.regs[50][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1341),
    .D(_01916_),
    .Q_N(_12052_),
    .Q(\top_ihp.oisc.regs[50][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1422),
    .D(_01917_),
    .Q_N(_12051_),
    .Q(\top_ihp.oisc.regs[50][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1290),
    .D(_01918_),
    .Q_N(_12050_),
    .Q(\top_ihp.oisc.regs[50][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1403),
    .D(_01919_),
    .Q_N(_12049_),
    .Q(\top_ihp.oisc.regs[50][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1351),
    .D(_01920_),
    .Q_N(_12048_),
    .Q(\top_ihp.oisc.regs[50][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1341),
    .D(_01921_),
    .Q_N(_12047_),
    .Q(\top_ihp.oisc.regs[50][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1346),
    .D(_01922_),
    .Q_N(_12046_),
    .Q(\top_ihp.oisc.regs[50][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1411),
    .D(_01923_),
    .Q_N(_12045_),
    .Q(\top_ihp.oisc.regs[50][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1368),
    .D(_01924_),
    .Q_N(_12044_),
    .Q(\top_ihp.oisc.regs[51][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1299),
    .D(_01925_),
    .Q_N(_12043_),
    .Q(\top_ihp.oisc.regs[51][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1366),
    .D(_01926_),
    .Q_N(_12042_),
    .Q(\top_ihp.oisc.regs[51][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1301),
    .D(_01927_),
    .Q_N(_12041_),
    .Q(\top_ihp.oisc.regs[51][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1367),
    .D(_01928_),
    .Q_N(_12040_),
    .Q(\top_ihp.oisc.regs[51][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1297),
    .D(_01929_),
    .Q_N(_12039_),
    .Q(\top_ihp.oisc.regs[51][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1299),
    .D(_01930_),
    .Q_N(_12038_),
    .Q(\top_ihp.oisc.regs[51][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1367),
    .D(_01931_),
    .Q_N(_12037_),
    .Q(\top_ihp.oisc.regs[51][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1375),
    .D(_01932_),
    .Q_N(_12036_),
    .Q(\top_ihp.oisc.regs[51][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1386),
    .D(_01933_),
    .Q_N(_12035_),
    .Q(\top_ihp.oisc.regs[51][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1386),
    .D(_01934_),
    .Q_N(_12034_),
    .Q(\top_ihp.oisc.regs[51][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1375),
    .D(_01935_),
    .Q_N(_12033_),
    .Q(\top_ihp.oisc.regs[51][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1411),
    .D(_01936_),
    .Q_N(_12032_),
    .Q(\top_ihp.oisc.regs[51][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1376),
    .D(_01937_),
    .Q_N(_12031_),
    .Q(\top_ihp.oisc.regs[51][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1377),
    .D(_01938_),
    .Q_N(_12030_),
    .Q(\top_ihp.oisc.regs[51][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1411),
    .D(_01939_),
    .Q_N(_12029_),
    .Q(\top_ihp.oisc.regs[51][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1349),
    .D(_01940_),
    .Q_N(_12028_),
    .Q(\top_ihp.oisc.regs[51][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1325),
    .D(_01941_),
    .Q_N(_12027_),
    .Q(\top_ihp.oisc.regs[51][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1396),
    .D(_01942_),
    .Q_N(_12026_),
    .Q(\top_ihp.oisc.regs[51][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1396),
    .D(_01943_),
    .Q_N(_12025_),
    .Q(\top_ihp.oisc.regs[51][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1404),
    .D(_01944_),
    .Q_N(_12024_),
    .Q(\top_ihp.oisc.regs[51][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1355),
    .D(_01945_),
    .Q_N(_12023_),
    .Q(\top_ihp.oisc.regs[51][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1359),
    .D(_01946_),
    .Q_N(_12022_),
    .Q(\top_ihp.oisc.regs[51][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1422),
    .D(_01947_),
    .Q_N(_12021_),
    .Q(\top_ihp.oisc.regs[51][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1354),
    .D(_01948_),
    .Q_N(_12020_),
    .Q(\top_ihp.oisc.regs[51][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1355),
    .D(_01949_),
    .Q_N(_12019_),
    .Q(\top_ihp.oisc.regs[51][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1408),
    .D(_01950_),
    .Q_N(_12018_),
    .Q(\top_ihp.oisc.regs[51][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1410),
    .D(_01951_),
    .Q_N(_12017_),
    .Q(\top_ihp.oisc.regs[51][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1351),
    .D(_01952_),
    .Q_N(_12016_),
    .Q(\top_ihp.oisc.regs[51][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1348),
    .D(_01953_),
    .Q_N(_12015_),
    .Q(\top_ihp.oisc.regs[51][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1329),
    .D(_01954_),
    .Q_N(_12014_),
    .Q(\top_ihp.oisc.regs[51][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1310),
    .D(_01955_),
    .Q_N(_12013_),
    .Q(\top_ihp.oisc.regs[51][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1319),
    .D(_01956_),
    .Q_N(_12012_),
    .Q(\top_ihp.oisc.regs[52][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1369),
    .D(_01957_),
    .Q_N(_12011_),
    .Q(\top_ihp.oisc.regs[52][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1313),
    .D(_01958_),
    .Q_N(_12010_),
    .Q(\top_ihp.oisc.regs[52][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1259),
    .D(_01959_),
    .Q_N(_12009_),
    .Q(\top_ihp.oisc.regs[52][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1318),
    .D(_01960_),
    .Q_N(_12008_),
    .Q(\top_ihp.oisc.regs[52][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1260),
    .D(_01961_),
    .Q_N(_12007_),
    .Q(\top_ihp.oisc.regs[52][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1299),
    .D(_01962_),
    .Q_N(_12006_),
    .Q(\top_ihp.oisc.regs[52][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1367),
    .D(_01963_),
    .Q_N(_12005_),
    .Q(\top_ihp.oisc.regs[52][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1368),
    .D(_01964_),
    .Q_N(_12004_),
    .Q(\top_ihp.oisc.regs[52][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1324),
    .D(_01965_),
    .Q_N(_12003_),
    .Q(\top_ihp.oisc.regs[52][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1386),
    .D(_01966_),
    .Q_N(_12002_),
    .Q(\top_ihp.oisc.regs[52][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1272),
    .D(_01967_),
    .Q_N(_12001_),
    .Q(\top_ihp.oisc.regs[52][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1411),
    .D(_01968_),
    .Q_N(_12000_),
    .Q(\top_ihp.oisc.regs[52][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1388),
    .D(_01969_),
    .Q_N(_11999_),
    .Q(\top_ihp.oisc.regs[52][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1377),
    .D(_01970_),
    .Q_N(_11998_),
    .Q(\top_ihp.oisc.regs[52][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1271),
    .D(_01971_),
    .Q_N(_11997_),
    .Q(\top_ihp.oisc.regs[52][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1400),
    .D(_01972_),
    .Q_N(_11996_),
    .Q(\top_ihp.oisc.regs[52][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1304),
    .D(_01973_),
    .Q_N(_11995_),
    .Q(\top_ihp.oisc.regs[52][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1413),
    .D(_01974_),
    .Q_N(_11994_),
    .Q(\top_ihp.oisc.regs[52][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1397),
    .D(_01975_),
    .Q_N(_11993_),
    .Q(\top_ihp.oisc.regs[52][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1421),
    .D(_01976_),
    .Q_N(_11992_),
    .Q(\top_ihp.oisc.regs[52][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1339),
    .D(_01977_),
    .Q_N(_11991_),
    .Q(\top_ihp.oisc.regs[52][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1293),
    .D(_01978_),
    .Q_N(_11990_),
    .Q(\top_ihp.oisc.regs[52][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1422),
    .D(_01979_),
    .Q_N(_11989_),
    .Q(\top_ihp.oisc.regs[52][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1336),
    .D(_01980_),
    .Q_N(_11988_),
    .Q(\top_ihp.oisc.regs[52][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1421),
    .D(_01981_),
    .Q_N(_11987_),
    .Q(\top_ihp.oisc.regs[52][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1409),
    .D(_01982_),
    .Q_N(_11986_),
    .Q(\top_ihp.oisc.regs[52][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1410),
    .D(_01983_),
    .Q_N(_11985_),
    .Q(\top_ihp.oisc.regs[52][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1286),
    .D(_01984_),
    .Q_N(_11984_),
    .Q(\top_ihp.oisc.regs[52][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1333),
    .D(_01985_),
    .Q_N(_11983_),
    .Q(\top_ihp.oisc.regs[52][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1284),
    .D(_01986_),
    .Q_N(_11982_),
    .Q(\top_ihp.oisc.regs[52][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1284),
    .D(_01987_),
    .Q_N(_11981_),
    .Q(\top_ihp.oisc.regs[52][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1369),
    .D(_01988_),
    .Q_N(_11980_),
    .Q(\top_ihp.oisc.regs[53][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1302),
    .D(_01989_),
    .Q_N(_11979_),
    .Q(\top_ihp.oisc.regs[53][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1367),
    .D(_01990_),
    .Q_N(_11978_),
    .Q(\top_ihp.oisc.regs[53][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1302),
    .D(_01991_),
    .Q_N(_11977_),
    .Q(\top_ihp.oisc.regs[53][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1298),
    .D(_01992_),
    .Q_N(_11976_),
    .Q(\top_ihp.oisc.regs[53][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1298),
    .D(_01993_),
    .Q_N(_11975_),
    .Q(\top_ihp.oisc.regs[53][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1299),
    .D(_01994_),
    .Q_N(_11974_),
    .Q(\top_ihp.oisc.regs[53][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1301),
    .D(_01995_),
    .Q_N(_11973_),
    .Q(\top_ihp.oisc.regs[53][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1377),
    .D(_01996_),
    .Q_N(_11972_),
    .Q(\top_ihp.oisc.regs[53][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1321),
    .D(_01997_),
    .Q_N(_11971_),
    .Q(\top_ihp.oisc.regs[53][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1389),
    .D(_01998_),
    .Q_N(_11970_),
    .Q(\top_ihp.oisc.regs[53][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1387),
    .D(_01999_),
    .Q_N(_11969_),
    .Q(\top_ihp.oisc.regs[53][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1389),
    .D(_02000_),
    .Q_N(_11968_),
    .Q(\top_ihp.oisc.regs[53][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1377),
    .D(_02001_),
    .Q_N(_11967_),
    .Q(\top_ihp.oisc.regs[53][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1324),
    .D(_02002_),
    .Q_N(_11966_),
    .Q(\top_ihp.oisc.regs[53][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1411),
    .D(_02003_),
    .Q_N(_11965_),
    .Q(\top_ihp.oisc.regs[53][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1395),
    .D(_02004_),
    .Q_N(_11964_),
    .Q(\top_ihp.oisc.regs[53][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1325),
    .D(_02005_),
    .Q_N(_11963_),
    .Q(\top_ihp.oisc.regs[53][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1401),
    .D(_02006_),
    .Q_N(_11962_),
    .Q(\top_ihp.oisc.regs[53][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1401),
    .D(_02007_),
    .Q_N(_11961_),
    .Q(\top_ihp.oisc.regs[53][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1404),
    .D(_02008_),
    .Q_N(_11960_),
    .Q(\top_ihp.oisc.regs[53][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1342),
    .D(_02009_),
    .Q_N(_11959_),
    .Q(\top_ihp.oisc.regs[53][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1409),
    .D(_02010_),
    .Q_N(_11958_),
    .Q(\top_ihp.oisc.regs[53][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1409),
    .D(_02011_),
    .Q_N(_11957_),
    .Q(\top_ihp.oisc.regs[53][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1344),
    .D(_02012_),
    .Q_N(_11956_),
    .Q(\top_ihp.oisc.regs[53][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1330),
    .D(_02013_),
    .Q_N(_11955_),
    .Q(\top_ihp.oisc.regs[53][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1421),
    .D(_02014_),
    .Q_N(_11954_),
    .Q(\top_ihp.oisc.regs[53][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1402),
    .D(_02015_),
    .Q_N(_11953_),
    .Q(\top_ihp.oisc.regs[53][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1352),
    .D(_02016_),
    .Q_N(_11952_),
    .Q(\top_ihp.oisc.regs[53][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1333),
    .D(_02017_),
    .Q_N(_11951_),
    .Q(\top_ihp.oisc.regs[53][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1332),
    .D(_02018_),
    .Q_N(_11950_),
    .Q(\top_ihp.oisc.regs[53][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1400),
    .D(_02019_),
    .Q_N(_11949_),
    .Q(\top_ihp.oisc.regs[53][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1315),
    .D(_02020_),
    .Q_N(_11948_),
    .Q(\top_ihp.oisc.regs[54][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1303),
    .D(_02021_),
    .Q_N(_11947_),
    .Q(\top_ihp.oisc.regs[54][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1313),
    .D(_02022_),
    .Q_N(_11946_),
    .Q(\top_ihp.oisc.regs[54][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1301),
    .D(_02023_),
    .Q_N(_11945_),
    .Q(\top_ihp.oisc.regs[54][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1317),
    .D(_02024_),
    .Q_N(_11944_),
    .Q(\top_ihp.oisc.regs[54][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1304),
    .D(_02025_),
    .Q_N(_11943_),
    .Q(\top_ihp.oisc.regs[54][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1297),
    .D(_02026_),
    .Q_N(_11942_),
    .Q(\top_ihp.oisc.regs[54][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1317),
    .D(_02027_),
    .Q_N(_11941_),
    .Q(\top_ihp.oisc.regs[54][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1308),
    .D(_02028_),
    .Q_N(_11940_),
    .Q(\top_ihp.oisc.regs[54][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1324),
    .D(_02029_),
    .Q_N(_11939_),
    .Q(\top_ihp.oisc.regs[54][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1267),
    .D(_02030_),
    .Q_N(_11938_),
    .Q(\top_ihp.oisc.regs[54][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1304),
    .D(_02031_),
    .Q_N(_11937_),
    .Q(\top_ihp.oisc.regs[54][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1322),
    .D(_02032_),
    .Q_N(_11936_),
    .Q(\top_ihp.oisc.regs[54][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1305),
    .D(_02033_),
    .Q_N(_11935_),
    .Q(\top_ihp.oisc.regs[54][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1321),
    .D(_02034_),
    .Q_N(_11934_),
    .Q(\top_ihp.oisc.regs[54][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1325),
    .D(_02035_),
    .Q_N(_11933_),
    .Q(\top_ihp.oisc.regs[54][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1323),
    .D(_02036_),
    .Q_N(_11932_),
    .Q(\top_ihp.oisc.regs[54][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1304),
    .D(_02037_),
    .Q_N(_11931_),
    .Q(\top_ihp.oisc.regs[54][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1287),
    .D(_02038_),
    .Q_N(_11930_),
    .Q(\top_ihp.oisc.regs[54][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1351),
    .D(_02039_),
    .Q_N(_11929_),
    .Q(\top_ihp.oisc.regs[54][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1360),
    .D(_02040_),
    .Q_N(_11928_),
    .Q(\top_ihp.oisc.regs[54][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1282),
    .D(_02041_),
    .Q_N(_11927_),
    .Q(\top_ihp.oisc.regs[54][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1359),
    .D(_02042_),
    .Q_N(_11926_),
    .Q(\top_ihp.oisc.regs[54][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1293),
    .D(_02043_),
    .Q_N(_11925_),
    .Q(\top_ihp.oisc.regs[54][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1355),
    .D(_02044_),
    .Q_N(_11924_),
    .Q(\top_ihp.oisc.regs[54][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1360),
    .D(_02045_),
    .Q_N(_11923_),
    .Q(\top_ihp.oisc.regs[54][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1338),
    .D(_02046_),
    .Q_N(_11922_),
    .Q(\top_ihp.oisc.regs[54][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1356),
    .D(_02047_),
    .Q_N(_11921_),
    .Q(\top_ihp.oisc.regs[54][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1290),
    .D(_02048_),
    .Q_N(_11920_),
    .Q(\top_ihp.oisc.regs[54][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1283),
    .D(_02049_),
    .Q_N(_11919_),
    .Q(\top_ihp.oisc.regs[54][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1330),
    .D(_02050_),
    .Q_N(_11918_),
    .Q(\top_ihp.oisc.regs[54][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1305),
    .D(_02051_),
    .Q_N(_11917_),
    .Q(\top_ihp.oisc.regs[54][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1316),
    .D(_02052_),
    .Q_N(_11916_),
    .Q(\top_ihp.oisc.regs[55][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1302),
    .D(_02053_),
    .Q_N(_11915_),
    .Q(\top_ihp.oisc.regs[55][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1314),
    .D(_02054_),
    .Q_N(_11914_),
    .Q(\top_ihp.oisc.regs[55][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1265),
    .D(_02055_),
    .Q_N(_11913_),
    .Q(\top_ihp.oisc.regs[55][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1298),
    .D(_02056_),
    .Q_N(_11912_),
    .Q(\top_ihp.oisc.regs[55][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1265),
    .D(_02057_),
    .Q_N(_11911_),
    .Q(\top_ihp.oisc.regs[55][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1265),
    .D(_02058_),
    .Q_N(_11910_),
    .Q(\top_ihp.oisc.regs[55][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1365),
    .D(_02059_),
    .Q_N(_11909_),
    .Q(\top_ihp.oisc.regs[55][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1371),
    .D(_02060_),
    .Q_N(_11908_),
    .Q(\top_ihp.oisc.regs[55][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1324),
    .D(_02061_),
    .Q_N(_11907_),
    .Q(\top_ihp.oisc.regs[55][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1372),
    .D(_02062_),
    .Q_N(_11906_),
    .Q(\top_ihp.oisc.regs[55][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1326),
    .D(_02063_),
    .Q_N(_11905_),
    .Q(\top_ihp.oisc.regs[55][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1325),
    .D(_02064_),
    .Q_N(_11904_),
    .Q(\top_ihp.oisc.regs[55][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1373),
    .D(_02065_),
    .Q_N(_11903_),
    .Q(\top_ihp.oisc.regs[55][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1321),
    .D(_02066_),
    .Q_N(_11902_),
    .Q(\top_ihp.oisc.regs[55][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1395),
    .D(_02067_),
    .Q_N(_11901_),
    .Q(\top_ihp.oisc.regs[55][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1398),
    .D(_02068_),
    .Q_N(_11900_),
    .Q(\top_ihp.oisc.regs[55][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1323),
    .D(_02069_),
    .Q_N(_11899_),
    .Q(\top_ihp.oisc.regs[55][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1397),
    .D(_02070_),
    .Q_N(_11898_),
    .Q(\top_ihp.oisc.regs[55][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1352),
    .D(_02071_),
    .Q_N(_11897_),
    .Q(\top_ihp.oisc.regs[55][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1292),
    .D(_02072_),
    .Q_N(_11896_),
    .Q(\top_ihp.oisc.regs[55][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1339),
    .D(_02073_),
    .Q_N(_11895_),
    .Q(\top_ihp.oisc.regs[55][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1408),
    .D(_02074_),
    .Q_N(_11894_),
    .Q(\top_ihp.oisc.regs[55][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1408),
    .D(_02075_),
    .Q_N(_11893_),
    .Q(\top_ihp.oisc.regs[55][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1355),
    .D(_02076_),
    .Q_N(_11892_),
    .Q(\top_ihp.oisc.regs[55][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1337),
    .D(_02077_),
    .Q_N(_11891_),
    .Q(\top_ihp.oisc.regs[55][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1292),
    .D(_02078_),
    .Q_N(_11890_),
    .Q(\top_ihp.oisc.regs[55][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1291),
    .D(_02079_),
    .Q_N(_11889_),
    .Q(\top_ihp.oisc.regs[55][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1358),
    .D(_02080_),
    .Q_N(_11888_),
    .Q(\top_ihp.oisc.regs[55][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1341),
    .D(_02081_),
    .Q_N(_11887_),
    .Q(\top_ihp.oisc.regs[55][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1346),
    .D(_02082_),
    .Q_N(_11886_),
    .Q(\top_ihp.oisc.regs[55][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1335),
    .D(_02083_),
    .Q_N(_11885_),
    .Q(\top_ihp.oisc.regs[55][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1313),
    .D(_02084_),
    .Q_N(_11884_),
    .Q(\top_ihp.oisc.regs[56][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1368),
    .D(_02085_),
    .Q_N(_11883_),
    .Q(\top_ihp.oisc.regs[56][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1366),
    .D(_02086_),
    .Q_N(_11882_),
    .Q(\top_ihp.oisc.regs[56][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1302),
    .D(_02087_),
    .Q_N(_11881_),
    .Q(\top_ihp.oisc.regs[56][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1369),
    .D(_02088_),
    .Q_N(_11880_),
    .Q(\top_ihp.oisc.regs[56][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1306),
    .D(_02089_),
    .Q_N(_11879_),
    .Q(\top_ihp.oisc.regs[56][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1300),
    .D(_02090_),
    .Q_N(_11878_),
    .Q(\top_ihp.oisc.regs[56][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1366),
    .D(_02091_),
    .Q_N(_11877_),
    .Q(\top_ihp.oisc.regs[56][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1324),
    .D(_02092_),
    .Q_N(_11876_),
    .Q(\top_ihp.oisc.regs[56][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1324),
    .D(_02093_),
    .Q_N(_11875_),
    .Q(\top_ihp.oisc.regs[56][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1305),
    .D(_02094_),
    .Q_N(_11874_),
    .Q(\top_ihp.oisc.regs[56][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1267),
    .D(_02095_),
    .Q_N(_11873_),
    .Q(\top_ihp.oisc.regs[56][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1325),
    .D(_02096_),
    .Q_N(_11872_),
    .Q(\top_ihp.oisc.regs[56][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1326),
    .D(_02097_),
    .Q_N(_11871_),
    .Q(\top_ihp.oisc.regs[56][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1273),
    .D(_02098_),
    .Q_N(_11870_),
    .Q(\top_ihp.oisc.regs[56][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1284),
    .D(_02099_),
    .Q_N(_11869_),
    .Q(\top_ihp.oisc.regs[56][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1350),
    .D(_02100_),
    .Q_N(_11868_),
    .Q(\top_ihp.oisc.regs[56][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1307),
    .D(_02101_),
    .Q_N(_11867_),
    .Q(\top_ihp.oisc.regs[56][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1287),
    .D(_02102_),
    .Q_N(_11866_),
    .Q(\top_ihp.oisc.regs[56][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1352),
    .D(_02103_),
    .Q_N(_11865_),
    .Q(\top_ihp.oisc.regs[56][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1283),
    .D(_02104_),
    .Q_N(_11864_),
    .Q(\top_ihp.oisc.regs[56][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1339),
    .D(_02105_),
    .Q_N(_11863_),
    .Q(\top_ihp.oisc.regs[56][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1405),
    .D(_02106_),
    .Q_N(_11862_),
    .Q(\top_ihp.oisc.regs[56][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1288),
    .D(_02107_),
    .Q_N(_11861_),
    .Q(\top_ihp.oisc.regs[56][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1354),
    .D(_02108_),
    .Q_N(_11860_),
    .Q(\top_ihp.oisc.regs[56][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1283),
    .D(_02109_),
    .Q_N(_11859_),
    .Q(\top_ihp.oisc.regs[56][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1405),
    .D(_02110_),
    .Q_N(_11858_),
    .Q(\top_ihp.oisc.regs[56][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1407),
    .D(_02111_),
    .Q_N(_11857_),
    .Q(\top_ihp.oisc.regs[56][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1357),
    .D(_02112_),
    .Q_N(_11856_),
    .Q(\top_ihp.oisc.regs[56][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1294),
    .D(_02113_),
    .Q_N(_11855_),
    .Q(\top_ihp.oisc.regs[56][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1346),
    .D(_02114_),
    .Q_N(_11854_),
    .Q(\top_ihp.oisc.regs[56][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1332),
    .D(_02115_),
    .Q_N(_11853_),
    .Q(\top_ihp.oisc.regs[56][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1314),
    .D(_02116_),
    .Q_N(_11852_),
    .Q(\top_ihp.oisc.regs[57][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1370),
    .D(_02117_),
    .Q_N(_11851_),
    .Q(\top_ihp.oisc.regs[57][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1365),
    .D(_02118_),
    .Q_N(_11850_),
    .Q(\top_ihp.oisc.regs[57][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1298),
    .D(_02119_),
    .Q_N(_11849_),
    .Q(\top_ihp.oisc.regs[57][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1365),
    .D(_02120_),
    .Q_N(_11848_),
    .Q(\top_ihp.oisc.regs[57][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1306),
    .D(_02121_),
    .Q_N(_11847_),
    .Q(\top_ihp.oisc.regs[57][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1298),
    .D(_02122_),
    .Q_N(_11846_),
    .Q(\top_ihp.oisc.regs[57][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1366),
    .D(_02123_),
    .Q_N(_11845_),
    .Q(\top_ihp.oisc.regs[57][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1321),
    .D(_02124_),
    .Q_N(_11844_),
    .Q(\top_ihp.oisc.regs[57][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1324),
    .D(_02125_),
    .Q_N(_11843_),
    .Q(\top_ihp.oisc.regs[57][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1373),
    .D(_02126_),
    .Q_N(_11842_),
    .Q(\top_ihp.oisc.regs[57][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1327),
    .D(_02127_),
    .Q_N(_11841_),
    .Q(\top_ihp.oisc.regs[57][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1322),
    .D(_02128_),
    .Q_N(_11840_),
    .Q(\top_ihp.oisc.regs[57][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1373),
    .D(_02129_),
    .Q_N(_11839_),
    .Q(\top_ihp.oisc.regs[57][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1308),
    .D(_02130_),
    .Q_N(_11838_),
    .Q(\top_ihp.oisc.regs[57][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1326),
    .D(_02131_),
    .Q_N(_11837_),
    .Q(\top_ihp.oisc.regs[57][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1349),
    .D(_02132_),
    .Q_N(_11836_),
    .Q(\top_ihp.oisc.regs[57][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1308),
    .D(_02133_),
    .Q_N(_11835_),
    .Q(\top_ihp.oisc.regs[57][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1397),
    .D(_02134_),
    .Q_N(_11834_),
    .Q(\top_ihp.oisc.regs[57][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1397),
    .D(_02135_),
    .Q_N(_11833_),
    .Q(\top_ihp.oisc.regs[57][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1360),
    .D(_02136_),
    .Q_N(_11832_),
    .Q(\top_ihp.oisc.regs[57][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1338),
    .D(_02137_),
    .Q_N(_11831_),
    .Q(\top_ihp.oisc.regs[57][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1404),
    .D(_02138_),
    .Q_N(_11830_),
    .Q(\top_ihp.oisc.regs[57][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1338),
    .D(_02139_),
    .Q_N(_11829_),
    .Q(\top_ihp.oisc.regs[57][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1338),
    .D(_02140_),
    .Q_N(_11828_),
    .Q(\top_ihp.oisc.regs[57][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1343),
    .D(_02141_),
    .Q_N(_11827_),
    .Q(\top_ihp.oisc.regs[57][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1340),
    .D(_02142_),
    .Q_N(_11826_),
    .Q(\top_ihp.oisc.regs[57][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1402),
    .D(_02143_),
    .Q_N(_11825_),
    .Q(\top_ihp.oisc.regs[57][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1361),
    .D(_02144_),
    .Q_N(_11824_),
    .Q(\top_ihp.oisc.regs[57][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1354),
    .D(_02145_),
    .Q_N(_11823_),
    .Q(\top_ihp.oisc.regs[57][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1329),
    .D(_02146_),
    .Q_N(_11822_),
    .Q(\top_ihp.oisc.regs[57][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1309),
    .D(_02147_),
    .Q_N(_11821_),
    .Q(\top_ihp.oisc.regs[57][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1251),
    .D(_02148_),
    .Q_N(_11820_),
    .Q(\top_ihp.oisc.regs[58][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1303),
    .D(_02149_),
    .Q_N(_11819_),
    .Q(\top_ihp.oisc.regs[58][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1314),
    .D(_02150_),
    .Q_N(_11818_),
    .Q(\top_ihp.oisc.regs[58][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1298),
    .D(_02151_),
    .Q_N(_11817_),
    .Q(\top_ihp.oisc.regs[58][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1365),
    .D(_02152_),
    .Q_N(_11816_),
    .Q(\top_ihp.oisc.regs[58][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1255),
    .D(_02153_),
    .Q_N(_11815_),
    .Q(\top_ihp.oisc.regs[58][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1264),
    .D(_02154_),
    .Q_N(_11814_),
    .Q(\top_ihp.oisc.regs[58][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1365),
    .D(_02155_),
    .Q_N(_11813_),
    .Q(\top_ihp.oisc.regs[58][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1371),
    .D(_02156_),
    .Q_N(_11812_),
    .Q(\top_ihp.oisc.regs[58][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1371),
    .D(_02157_),
    .Q_N(_11811_),
    .Q(\top_ihp.oisc.regs[58][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1371),
    .D(_02158_),
    .Q_N(_11810_),
    .Q(\top_ihp.oisc.regs[58][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1327),
    .D(_02159_),
    .Q_N(_11809_),
    .Q(\top_ihp.oisc.regs[58][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1331),
    .D(_02160_),
    .Q_N(_11808_),
    .Q(\top_ihp.oisc.regs[58][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1322),
    .D(_02161_),
    .Q_N(_11807_),
    .Q(\top_ihp.oisc.regs[58][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1307),
    .D(_02162_),
    .Q_N(_11806_),
    .Q(\top_ihp.oisc.regs[58][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1256),
    .D(_02163_),
    .Q_N(_11805_),
    .Q(\top_ihp.oisc.regs[58][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1348),
    .D(_02164_),
    .Q_N(_11804_),
    .Q(\top_ihp.oisc.regs[58][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1256),
    .D(_02165_),
    .Q_N(_11803_),
    .Q(\top_ihp.oisc.regs[58][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1278),
    .D(_02166_),
    .Q_N(_11802_),
    .Q(\top_ihp.oisc.regs[58][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1397),
    .D(_02167_),
    .Q_N(_11801_),
    .Q(\top_ihp.oisc.regs[58][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1288),
    .D(_02168_),
    .Q_N(_11800_),
    .Q(\top_ihp.oisc.regs[58][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1355),
    .D(_02169_),
    .Q_N(_11799_),
    .Q(\top_ihp.oisc.regs[58][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1339),
    .D(_02170_),
    .Q_N(_11798_),
    .Q(\top_ihp.oisc.regs[58][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1405),
    .D(_02171_),
    .Q_N(_11797_),
    .Q(\top_ihp.oisc.regs[58][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1288),
    .D(_02172_),
    .Q_N(_11796_),
    .Q(\top_ihp.oisc.regs[58][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1289),
    .D(_02173_),
    .Q_N(_11795_),
    .Q(\top_ihp.oisc.regs[58][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1405),
    .D(_02174_),
    .Q_N(_11794_),
    .Q(\top_ihp.oisc.regs[58][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1403),
    .D(_02175_),
    .Q_N(_11793_),
    .Q(\top_ihp.oisc.regs[58][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1352),
    .D(_02176_),
    .Q_N(_11792_),
    .Q(\top_ihp.oisc.regs[58][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1334),
    .D(_02177_),
    .Q_N(_11791_),
    .Q(\top_ihp.oisc.regs[58][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1346),
    .D(_02178_),
    .Q_N(_11790_),
    .Q(\top_ihp.oisc.regs[58][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1309),
    .D(_02179_),
    .Q_N(_11789_),
    .Q(\top_ihp.oisc.regs[58][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1316),
    .D(_02180_),
    .Q_N(_11788_),
    .Q(\top_ihp.oisc.regs[59][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1366),
    .D(_02181_),
    .Q_N(_11787_),
    .Q(\top_ihp.oisc.regs[59][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1366),
    .D(_02182_),
    .Q_N(_11786_),
    .Q(\top_ihp.oisc.regs[59][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1300),
    .D(_02183_),
    .Q_N(_11785_),
    .Q(\top_ihp.oisc.regs[59][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1318),
    .D(_02184_),
    .Q_N(_11784_),
    .Q(\top_ihp.oisc.regs[59][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1297),
    .D(_02185_),
    .Q_N(_11783_),
    .Q(\top_ihp.oisc.regs[59][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1299),
    .D(_02186_),
    .Q_N(_11782_),
    .Q(\top_ihp.oisc.regs[59][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1297),
    .D(_02187_),
    .Q_N(_11781_),
    .Q(\top_ihp.oisc.regs[59][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1375),
    .D(_02188_),
    .Q_N(_11780_),
    .Q(\top_ihp.oisc.regs[59][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1371),
    .D(_02189_),
    .Q_N(_11779_),
    .Q(\top_ihp.oisc.regs[59][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1375),
    .D(_02190_),
    .Q_N(_11778_),
    .Q(\top_ihp.oisc.regs[59][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1257),
    .D(_02191_),
    .Q_N(_11777_),
    .Q(\top_ihp.oisc.regs[59][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1400),
    .D(_02192_),
    .Q_N(_11776_),
    .Q(\top_ihp.oisc.regs[59][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1271),
    .D(_02193_),
    .Q_N(_11775_),
    .Q(\top_ihp.oisc.regs[59][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1257),
    .D(_02194_),
    .Q_N(_11774_),
    .Q(\top_ihp.oisc.regs[59][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1284),
    .D(_02195_),
    .Q_N(_11773_),
    .Q(\top_ihp.oisc.regs[59][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1277),
    .D(_02196_),
    .Q_N(_11772_),
    .Q(\top_ihp.oisc.regs[59][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1257),
    .D(_02197_),
    .Q_N(_11771_),
    .Q(\top_ihp.oisc.regs[59][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1399),
    .D(_02198_),
    .Q_N(_11770_),
    .Q(\top_ihp.oisc.regs[59][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1287),
    .D(_02199_),
    .Q_N(_11769_),
    .Q(\top_ihp.oisc.regs[59][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1359),
    .D(_02200_),
    .Q_N(_11768_),
    .Q(\top_ihp.oisc.regs[59][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1342),
    .D(_02201_),
    .Q_N(_11767_),
    .Q(\top_ihp.oisc.regs[59][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1408),
    .D(_02202_),
    .Q_N(_11766_),
    .Q(\top_ihp.oisc.regs[59][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1408),
    .D(_02203_),
    .Q_N(_11765_),
    .Q(\top_ihp.oisc.regs[59][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1342),
    .D(_02204_),
    .Q_N(_11764_),
    .Q(\top_ihp.oisc.regs[59][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1343),
    .D(_02205_),
    .Q_N(_11763_),
    .Q(\top_ihp.oisc.regs[59][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1341),
    .D(_02206_),
    .Q_N(_11762_),
    .Q(\top_ihp.oisc.regs[59][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1407),
    .D(_02207_),
    .Q_N(_11761_),
    .Q(\top_ihp.oisc.regs[59][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1361),
    .D(_02208_),
    .Q_N(_11760_),
    .Q(\top_ihp.oisc.regs[59][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1344),
    .D(_02209_),
    .Q_N(_11759_),
    .Q(\top_ihp.oisc.regs[59][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1329),
    .D(_02210_),
    .Q_N(_11758_),
    .Q(\top_ihp.oisc.regs[59][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1332),
    .D(_02211_),
    .Q_N(_11757_),
    .Q(\top_ihp.oisc.regs[59][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1223),
    .D(_02212_),
    .Q_N(_11756_),
    .Q(\top_ihp.oisc.regs[5][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1167),
    .D(_02213_),
    .Q_N(_11755_),
    .Q(\top_ihp.oisc.regs[5][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1175),
    .D(_02214_),
    .Q_N(_11754_),
    .Q(\top_ihp.oisc.regs[5][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1220),
    .D(_02215_),
    .Q_N(_11753_),
    .Q(\top_ihp.oisc.regs[5][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1219),
    .D(_02216_),
    .Q_N(_11752_),
    .Q(\top_ihp.oisc.regs[5][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1208),
    .D(_02217_),
    .Q_N(_11751_),
    .Q(\top_ihp.oisc.regs[5][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1177),
    .D(_02218_),
    .Q_N(_11750_),
    .Q(\top_ihp.oisc.regs[5][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1220),
    .D(_02219_),
    .Q_N(_11749_),
    .Q(\top_ihp.oisc.regs[5][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1169),
    .D(_02220_),
    .Q_N(_11748_),
    .Q(\top_ihp.oisc.regs[5][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1172),
    .D(_02221_),
    .Q_N(_11747_),
    .Q(\top_ihp.oisc.regs[5][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1223),
    .D(_02222_),
    .Q_N(_11746_),
    .Q(\top_ihp.oisc.regs[5][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1225),
    .D(_02223_),
    .Q_N(_11745_),
    .Q(\top_ihp.oisc.regs[5][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1183),
    .D(_02224_),
    .Q_N(_11744_),
    .Q(\top_ihp.oisc.regs[5][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1173),
    .D(_02225_),
    .Q_N(_11743_),
    .Q(\top_ihp.oisc.regs[5][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1223),
    .D(_02226_),
    .Q_N(_11742_),
    .Q(\top_ihp.oisc.regs[5][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1227),
    .D(_02227_),
    .Q_N(_11741_),
    .Q(\top_ihp.oisc.regs[5][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1224),
    .D(_02228_),
    .Q_N(_11740_),
    .Q(\top_ihp.oisc.regs[5][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1224),
    .D(_02229_),
    .Q_N(_11739_),
    .Q(\top_ihp.oisc.regs[5][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1239),
    .D(_02230_),
    .Q_N(_11738_),
    .Q(\top_ihp.oisc.regs[5][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1197),
    .D(_02231_),
    .Q_N(_11737_),
    .Q(\top_ihp.oisc.regs[5][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1246),
    .D(_02232_),
    .Q_N(_11736_),
    .Q(\top_ihp.oisc.regs[5][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1246),
    .D(_02233_),
    .Q_N(_11735_),
    .Q(\top_ihp.oisc.regs[5][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1246),
    .D(_02234_),
    .Q_N(_11734_),
    .Q(\top_ihp.oisc.regs[5][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1193),
    .D(_02235_),
    .Q_N(_11733_),
    .Q(\top_ihp.oisc.regs[5][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1201),
    .D(_02236_),
    .Q_N(_11732_),
    .Q(\top_ihp.oisc.regs[5][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1193),
    .D(_02237_),
    .Q_N(_11731_),
    .Q(\top_ihp.oisc.regs[5][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1193),
    .D(_02238_),
    .Q_N(_11730_),
    .Q(\top_ihp.oisc.regs[5][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1193),
    .D(_02239_),
    .Q_N(_11729_),
    .Q(\top_ihp.oisc.regs[5][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1243),
    .D(_02240_),
    .Q_N(_11728_),
    .Q(\top_ihp.oisc.regs[5][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1243),
    .D(_02241_),
    .Q_N(_11727_),
    .Q(\top_ihp.oisc.regs[5][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1242),
    .D(_02242_),
    .Q_N(_11726_),
    .Q(\top_ihp.oisc.regs[5][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1224),
    .D(_02243_),
    .Q_N(_11725_),
    .Q(\top_ihp.oisc.regs[5][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1304),
    .D(_02244_),
    .Q_N(_11724_),
    .Q(\top_ihp.oisc.regs[60][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1368),
    .D(_02245_),
    .Q_N(_11723_),
    .Q(\top_ihp.oisc.regs[60][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1366),
    .D(_02246_),
    .Q_N(_11722_),
    .Q(\top_ihp.oisc.regs[60][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1301),
    .D(_02247_),
    .Q_N(_11721_),
    .Q(\top_ihp.oisc.regs[60][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1318),
    .D(_02248_),
    .Q_N(_11720_),
    .Q(\top_ihp.oisc.regs[60][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1300),
    .D(_02249_),
    .Q_N(_11719_),
    .Q(\top_ihp.oisc.regs[60][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1298),
    .D(_02250_),
    .Q_N(_11718_),
    .Q(\top_ihp.oisc.regs[60][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1370),
    .D(_02251_),
    .Q_N(_11717_),
    .Q(\top_ihp.oisc.regs[60][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1375),
    .D(_02252_),
    .Q_N(_11716_),
    .Q(\top_ihp.oisc.regs[60][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1374),
    .D(_02253_),
    .Q_N(_11715_),
    .Q(\top_ihp.oisc.regs[60][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1373),
    .D(_02254_),
    .Q_N(_11714_),
    .Q(\top_ihp.oisc.regs[60][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1309),
    .D(_02255_),
    .Q_N(_11713_),
    .Q(\top_ihp.oisc.regs[60][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1373),
    .D(_02256_),
    .Q_N(_11712_),
    .Q(\top_ihp.oisc.regs[60][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1376),
    .D(_02257_),
    .Q_N(_11711_),
    .Q(\top_ihp.oisc.regs[60][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1310),
    .D(_02258_),
    .Q_N(_11710_),
    .Q(\top_ihp.oisc.regs[60][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1398),
    .D(_02259_),
    .Q_N(_11709_),
    .Q(\top_ihp.oisc.regs[60][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1398),
    .D(_02260_),
    .Q_N(_11708_),
    .Q(\top_ihp.oisc.regs[60][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1322),
    .D(_02261_),
    .Q_N(_11707_),
    .Q(\top_ihp.oisc.regs[60][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1396),
    .D(_02262_),
    .Q_N(_11706_),
    .Q(\top_ihp.oisc.regs[60][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1331),
    .D(_02263_),
    .Q_N(_11705_),
    .Q(\top_ihp.oisc.regs[60][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1360),
    .D(_02264_),
    .Q_N(_11704_),
    .Q(\top_ihp.oisc.regs[60][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1359),
    .D(_02265_),
    .Q_N(_11703_),
    .Q(\top_ihp.oisc.regs[60][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1404),
    .D(_02266_),
    .Q_N(_11702_),
    .Q(\top_ihp.oisc.regs[60][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1405),
    .D(_02267_),
    .Q_N(_11701_),
    .Q(\top_ihp.oisc.regs[60][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1289),
    .D(_02268_),
    .Q_N(_11700_),
    .Q(\top_ihp.oisc.regs[60][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1343),
    .D(_02269_),
    .Q_N(_11699_),
    .Q(\top_ihp.oisc.regs[60][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1290),
    .D(_02270_),
    .Q_N(_11698_),
    .Q(\top_ihp.oisc.regs[60][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1403),
    .D(_02271_),
    .Q_N(_11697_),
    .Q(\top_ihp.oisc.regs[60][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1336),
    .D(_02272_),
    .Q_N(_11696_),
    .Q(\top_ihp.oisc.regs[60][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1344),
    .D(_02273_),
    .Q_N(_11695_),
    .Q(\top_ihp.oisc.regs[60][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1329),
    .D(_02274_),
    .Q_N(_11694_),
    .Q(\top_ihp.oisc.regs[60][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1309),
    .D(_02275_),
    .Q_N(_11693_),
    .Q(\top_ihp.oisc.regs[60][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1315),
    .D(_02276_),
    .Q_N(_11692_),
    .Q(\top_ihp.oisc.regs[61][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1320),
    .D(_02277_),
    .Q_N(_11691_),
    .Q(\top_ihp.oisc.regs[61][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1313),
    .D(_02278_),
    .Q_N(_11690_),
    .Q(\top_ihp.oisc.regs[61][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1301),
    .D(_02279_),
    .Q_N(_11689_),
    .Q(\top_ihp.oisc.regs[61][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1318),
    .D(_02280_),
    .Q_N(_11688_),
    .Q(\top_ihp.oisc.regs[61][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1264),
    .D(_02281_),
    .Q_N(_11687_),
    .Q(\top_ihp.oisc.regs[61][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1262),
    .D(_02282_),
    .Q_N(_11686_),
    .Q(\top_ihp.oisc.regs[61][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1317),
    .D(_02283_),
    .Q_N(_11685_),
    .Q(\top_ihp.oisc.regs[61][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1269),
    .D(_02284_),
    .Q_N(_11684_),
    .Q(\top_ihp.oisc.regs[61][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1327),
    .D(_02285_),
    .Q_N(_11683_),
    .Q(\top_ihp.oisc.regs[61][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1325),
    .D(_02286_),
    .Q_N(_11682_),
    .Q(\top_ihp.oisc.regs[61][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1326),
    .D(_02287_),
    .Q_N(_11681_),
    .Q(\top_ihp.oisc.regs[61][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1285),
    .D(_02288_),
    .Q_N(_11680_),
    .Q(\top_ihp.oisc.regs[61][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1326),
    .D(_02289_),
    .Q_N(_11679_),
    .Q(\top_ihp.oisc.regs[61][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1270),
    .D(_02290_),
    .Q_N(_11678_),
    .Q(\top_ihp.oisc.regs[61][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1349),
    .D(_02291_),
    .Q_N(_11677_),
    .Q(\top_ihp.oisc.regs[61][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1350),
    .D(_02292_),
    .Q_N(_11676_),
    .Q(\top_ihp.oisc.regs[61][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1323),
    .D(_02293_),
    .Q_N(_11675_),
    .Q(\top_ihp.oisc.regs[61][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1351),
    .D(_02294_),
    .Q_N(_11674_),
    .Q(\top_ihp.oisc.regs[61][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1351),
    .D(_02295_),
    .Q_N(_11673_),
    .Q(\top_ihp.oisc.regs[61][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1359),
    .D(_02296_),
    .Q_N(_11672_),
    .Q(\top_ihp.oisc.regs[61][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1289),
    .D(_02297_),
    .Q_N(_11671_),
    .Q(\top_ihp.oisc.regs[61][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1356),
    .D(_02298_),
    .Q_N(_11670_),
    .Q(\top_ihp.oisc.regs[61][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1293),
    .D(_02299_),
    .Q_N(_11669_),
    .Q(\top_ihp.oisc.regs[61][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1356),
    .D(_02300_),
    .Q_N(_11668_),
    .Q(\top_ihp.oisc.regs[61][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1342),
    .D(_02301_),
    .Q_N(_11667_),
    .Q(\top_ihp.oisc.regs[61][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1289),
    .D(_02302_),
    .Q_N(_11666_),
    .Q(\top_ihp.oisc.regs[61][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1292),
    .D(_02303_),
    .Q_N(_11665_),
    .Q(\top_ihp.oisc.regs[61][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1290),
    .D(_02304_),
    .Q_N(_11664_),
    .Q(\top_ihp.oisc.regs[61][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1354),
    .D(_02305_),
    .Q_N(_11663_),
    .Q(\top_ihp.oisc.regs[61][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1284),
    .D(_02306_),
    .Q_N(_11662_),
    .Q(\top_ihp.oisc.regs[61][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1310),
    .D(_02307_),
    .Q_N(_11661_),
    .Q(\top_ihp.oisc.regs[61][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1303),
    .D(_02308_),
    .Q_N(_11660_),
    .Q(\top_ihp.oisc.regs[62][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1320),
    .D(_02309_),
    .Q_N(_11659_),
    .Q(\top_ihp.oisc.regs[62][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1314),
    .D(_02310_),
    .Q_N(_11658_),
    .Q(\top_ihp.oisc.regs[62][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1263),
    .D(_02311_),
    .Q_N(_11657_),
    .Q(\top_ihp.oisc.regs[62][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1317),
    .D(_02312_),
    .Q_N(_11656_),
    .Q(\top_ihp.oisc.regs[62][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1297),
    .D(_02313_),
    .Q_N(_11655_),
    .Q(\top_ihp.oisc.regs[62][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1264),
    .D(_02314_),
    .Q_N(_11654_),
    .Q(\top_ihp.oisc.regs[62][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1317),
    .D(_02315_),
    .Q_N(_11653_),
    .Q(\top_ihp.oisc.regs[62][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1307),
    .D(_02316_),
    .Q_N(_11652_),
    .Q(\top_ihp.oisc.regs[62][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1324),
    .D(_02317_),
    .Q_N(_11651_),
    .Q(\top_ihp.oisc.regs[62][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1306),
    .D(_02318_),
    .Q_N(_11650_),
    .Q(\top_ihp.oisc.regs[62][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1304),
    .D(_02319_),
    .Q_N(_11649_),
    .Q(\top_ihp.oisc.regs[62][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1400),
    .D(_02320_),
    .Q_N(_11648_),
    .Q(\top_ihp.oisc.regs[62][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1373),
    .D(_02321_),
    .Q_N(_11647_),
    .Q(\top_ihp.oisc.regs[62][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1305),
    .D(_02322_),
    .Q_N(_11646_),
    .Q(\top_ihp.oisc.regs[62][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1349),
    .D(_02323_),
    .Q_N(_11645_),
    .Q(\top_ihp.oisc.regs[62][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1395),
    .D(_02324_),
    .Q_N(_11644_),
    .Q(\top_ihp.oisc.regs[62][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1307),
    .D(_02325_),
    .Q_N(_11643_),
    .Q(\top_ihp.oisc.regs[62][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1399),
    .D(_02326_),
    .Q_N(_11642_),
    .Q(\top_ihp.oisc.regs[62][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1330),
    .D(_02327_),
    .Q_N(_11641_),
    .Q(\top_ihp.oisc.regs[62][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1282),
    .D(_02328_),
    .Q_N(_11640_),
    .Q(\top_ihp.oisc.regs[62][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1282),
    .D(_02329_),
    .Q_N(_11639_),
    .Q(\top_ihp.oisc.regs[62][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1409),
    .D(_02330_),
    .Q_N(_11638_),
    .Q(\top_ihp.oisc.regs[62][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1409),
    .D(_02331_),
    .Q_N(_11637_),
    .Q(\top_ihp.oisc.regs[62][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1288),
    .D(_02332_),
    .Q_N(_11636_),
    .Q(\top_ihp.oisc.regs[62][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1343),
    .D(_02333_),
    .Q_N(_11635_),
    .Q(\top_ihp.oisc.regs[62][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1283),
    .D(_02334_),
    .Q_N(_11634_),
    .Q(\top_ihp.oisc.regs[62][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1403),
    .D(_02335_),
    .Q_N(_11633_),
    .Q(\top_ihp.oisc.regs[62][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1286),
    .D(_02336_),
    .Q_N(_11632_),
    .Q(\top_ihp.oisc.regs[62][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1334),
    .D(_02337_),
    .Q_N(_11631_),
    .Q(\top_ihp.oisc.regs[62][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1285),
    .D(_02338_),
    .Q_N(_11630_),
    .Q(\top_ihp.oisc.regs[62][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1310),
    .D(_02339_),
    .Q_N(_11629_),
    .Q(\top_ihp.oisc.regs[62][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1259),
    .D(_02340_),
    .Q_N(_11628_),
    .Q(\top_ihp.oisc.regs[63][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1249),
    .D(_02341_),
    .Q_N(_11627_),
    .Q(\top_ihp.oisc.regs[63][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1259),
    .D(_02342_),
    .Q_N(_11626_),
    .Q(\top_ihp.oisc.regs[63][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1250),
    .D(_02343_),
    .Q_N(_11625_),
    .Q(\top_ihp.oisc.regs[63][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1248),
    .D(_02344_),
    .Q_N(_11624_),
    .Q(\top_ihp.oisc.regs[63][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1248),
    .D(_02345_),
    .Q_N(_11623_),
    .Q(\top_ihp.oisc.regs[63][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1259),
    .D(_02346_),
    .Q_N(_11622_),
    .Q(\top_ihp.oisc.regs[63][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1248),
    .D(_02347_),
    .Q_N(_11621_),
    .Q(\top_ihp.oisc.regs[63][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1253),
    .D(_02348_),
    .Q_N(_11620_),
    .Q(\top_ihp.oisc.regs[63][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1249),
    .D(_02349_),
    .Q_N(_11619_),
    .Q(\top_ihp.oisc.regs[63][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1253),
    .D(_02350_),
    .Q_N(_11618_),
    .Q(\top_ihp.oisc.regs[63][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1253),
    .D(_02351_),
    .Q_N(_11617_),
    .Q(\top_ihp.oisc.regs[63][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1276),
    .D(_02352_),
    .Q_N(_11616_),
    .Q(\top_ihp.oisc.regs[63][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1256),
    .D(_02353_),
    .Q_N(_11615_),
    .Q(\top_ihp.oisc.regs[63][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1253),
    .D(_02354_),
    .Q_N(_11614_),
    .Q(\top_ihp.oisc.regs[63][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1254),
    .D(_02355_),
    .Q_N(_11613_),
    .Q(\top_ihp.oisc.regs[63][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1275),
    .D(_02356_),
    .Q_N(_11612_),
    .Q(\top_ihp.oisc.regs[63][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1253),
    .D(_02357_),
    .Q_N(_11611_),
    .Q(\top_ihp.oisc.regs[63][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1278),
    .D(_02358_),
    .Q_N(_11610_),
    .Q(\top_ihp.oisc.regs[63][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1278),
    .D(_02359_),
    .Q_N(_11609_),
    .Q(\top_ihp.oisc.regs[63][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1279),
    .D(_02360_),
    .Q_N(_11608_),
    .Q(\top_ihp.oisc.regs[63][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1279),
    .D(_02361_),
    .Q_N(_11607_),
    .Q(\top_ihp.oisc.regs[63][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1279),
    .D(_02362_),
    .Q_N(_11606_),
    .Q(\top_ihp.oisc.regs[63][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1279),
    .D(_02363_),
    .Q_N(_11605_),
    .Q(\top_ihp.oisc.regs[63][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1280),
    .D(_02364_),
    .Q_N(_11604_),
    .Q(\top_ihp.oisc.regs[63][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1280),
    .D(_02365_),
    .Q_N(_11603_),
    .Q(\top_ihp.oisc.regs[63][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1280),
    .D(_02366_),
    .Q_N(_11602_),
    .Q(\top_ihp.oisc.regs[63][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1279),
    .D(_02367_),
    .Q_N(_11601_),
    .Q(\top_ihp.oisc.regs[63][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1280),
    .D(_02368_),
    .Q_N(_11600_),
    .Q(\top_ihp.oisc.regs[63][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1280),
    .D(_02369_),
    .Q_N(_11599_),
    .Q(\top_ihp.oisc.regs[63][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1275),
    .D(_02370_),
    .Q_N(_11598_),
    .Q(\top_ihp.oisc.regs[63][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1275),
    .D(_02371_),
    .Q_N(_11597_),
    .Q(\top_ihp.oisc.regs[63][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1214),
    .D(_02372_),
    .Q_N(_11596_),
    .Q(\top_ihp.oisc.regs[6][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1167),
    .D(_02373_),
    .Q_N(_11595_),
    .Q(\top_ihp.oisc.regs[6][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1168),
    .D(_02374_),
    .Q_N(_11594_),
    .Q(\top_ihp.oisc.regs[6][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1176),
    .D(_02375_),
    .Q_N(_11593_),
    .Q(\top_ihp.oisc.regs[6][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1168),
    .D(_02376_),
    .Q_N(_11592_),
    .Q(\top_ihp.oisc.regs[6][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1210),
    .D(_02377_),
    .Q_N(_11591_),
    .Q(\top_ihp.oisc.regs[6][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1177),
    .D(_02378_),
    .Q_N(_11590_),
    .Q(\top_ihp.oisc.regs[6][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1210),
    .D(_02379_),
    .Q_N(_11589_),
    .Q(\top_ihp.oisc.regs[6][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1176),
    .D(_02380_),
    .Q_N(_11588_),
    .Q(\top_ihp.oisc.regs[6][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1167),
    .D(_02381_),
    .Q_N(_11587_),
    .Q(\top_ihp.oisc.regs[6][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1173),
    .D(_02382_),
    .Q_N(_11586_),
    .Q(\top_ihp.oisc.regs[6][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1180),
    .D(_02383_),
    .Q_N(_11585_),
    .Q(\top_ihp.oisc.regs[6][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1198),
    .D(_02384_),
    .Q_N(_11584_),
    .Q(\top_ihp.oisc.regs[6][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1188),
    .D(_02385_),
    .Q_N(_11583_),
    .Q(\top_ihp.oisc.regs[6][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1183),
    .D(_02386_),
    .Q_N(_11582_),
    .Q(\top_ihp.oisc.regs[6][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1181),
    .D(_02387_),
    .Q_N(_11581_),
    .Q(\top_ihp.oisc.regs[6][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1198),
    .D(_02388_),
    .Q_N(_11580_),
    .Q(\top_ihp.oisc.regs[6][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1173),
    .D(_02389_),
    .Q_N(_11579_),
    .Q(\top_ihp.oisc.regs[6][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1197),
    .D(_02390_),
    .Q_N(_11578_),
    .Q(\top_ihp.oisc.regs[6][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1189),
    .D(_02391_),
    .Q_N(_11577_),
    .Q(\top_ihp.oisc.regs[6][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1204),
    .D(_02392_),
    .Q_N(_11576_),
    .Q(\top_ihp.oisc.regs[6][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1235),
    .D(_02393_),
    .Q_N(_11575_),
    .Q(\top_ihp.oisc.regs[6][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1235),
    .D(_02394_),
    .Q_N(_11574_),
    .Q(\top_ihp.oisc.regs[6][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1193),
    .D(_02395_),
    .Q_N(_11573_),
    .Q(\top_ihp.oisc.regs[6][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1201),
    .D(_02396_),
    .Q_N(_11572_),
    .Q(\top_ihp.oisc.regs[6][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1189),
    .D(_02397_),
    .Q_N(_11571_),
    .Q(\top_ihp.oisc.regs[6][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1193),
    .D(_02398_),
    .Q_N(_11570_),
    .Q(\top_ihp.oisc.regs[6][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1195),
    .D(_02399_),
    .Q_N(_11569_),
    .Q(\top_ihp.oisc.regs[6][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1230),
    .D(_02400_),
    .Q_N(_11568_),
    .Q(\top_ihp.oisc.regs[6][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1199),
    .D(_02401_),
    .Q_N(_11567_),
    .Q(\top_ihp.oisc.regs[6][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1230),
    .D(_02402_),
    .Q_N(_11566_),
    .Q(\top_ihp.oisc.regs[6][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1217),
    .D(_02403_),
    .Q_N(_11565_),
    .Q(\top_ihp.oisc.regs[6][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1209),
    .D(_02404_),
    .Q_N(_11564_),
    .Q(\top_ihp.oisc.regs[7][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1167),
    .D(_02405_),
    .Q_N(_11563_),
    .Q(\top_ihp.oisc.regs[7][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1165),
    .D(_02406_),
    .Q_N(_11562_),
    .Q(\top_ihp.oisc.regs[7][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1175),
    .D(_02407_),
    .Q_N(_11561_),
    .Q(\top_ihp.oisc.regs[7][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1165),
    .D(_02408_),
    .Q_N(_11560_),
    .Q(\top_ihp.oisc.regs[7][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1208),
    .D(_02409_),
    .Q_N(_11559_),
    .Q(\top_ihp.oisc.regs[7][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1208),
    .D(_02410_),
    .Q_N(_11558_),
    .Q(\top_ihp.oisc.regs[7][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1209),
    .D(_02411_),
    .Q_N(_11557_),
    .Q(\top_ihp.oisc.regs[7][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1176),
    .D(_02412_),
    .Q_N(_11556_),
    .Q(\top_ihp.oisc.regs[7][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1167),
    .D(_02413_),
    .Q_N(_11555_),
    .Q(\top_ihp.oisc.regs[7][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1154),
    .D(_02414_),
    .Q_N(_11554_),
    .Q(\top_ihp.oisc.regs[7][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1180),
    .D(_02415_),
    .Q_N(_11553_),
    .Q(\top_ihp.oisc.regs[7][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1217),
    .D(_02416_),
    .Q_N(_11552_),
    .Q(\top_ihp.oisc.regs[7][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1155),
    .D(_02417_),
    .Q_N(_11551_),
    .Q(\top_ihp.oisc.regs[7][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1213),
    .D(_02418_),
    .Q_N(_11550_),
    .Q(\top_ihp.oisc.regs[7][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1181),
    .D(_02419_),
    .Q_N(_11549_),
    .Q(\top_ihp.oisc.regs[7][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1229),
    .D(_02420_),
    .Q_N(_11548_),
    .Q(\top_ihp.oisc.regs[7][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1170),
    .D(_02421_),
    .Q_N(_11547_),
    .Q(\top_ihp.oisc.regs[7][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1199),
    .D(_02422_),
    .Q_N(_11546_),
    .Q(\top_ihp.oisc.regs[7][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1188),
    .D(_02423_),
    .Q_N(_11545_),
    .Q(\top_ihp.oisc.regs[7][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1204),
    .D(_02424_),
    .Q_N(_11544_),
    .Q(\top_ihp.oisc.regs[7][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1204),
    .D(_02425_),
    .Q_N(_11543_),
    .Q(\top_ihp.oisc.regs[7][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1235),
    .D(_02426_),
    .Q_N(_11542_),
    .Q(\top_ihp.oisc.regs[7][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1195),
    .D(_02427_),
    .Q_N(_11541_),
    .Q(\top_ihp.oisc.regs[7][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1202),
    .D(_02428_),
    .Q_N(_11540_),
    .Q(\top_ihp.oisc.regs[7][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1189),
    .D(_02429_),
    .Q_N(_11539_),
    .Q(\top_ihp.oisc.regs[7][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1195),
    .D(_02430_),
    .Q_N(_11538_),
    .Q(\top_ihp.oisc.regs[7][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1192),
    .D(_02431_),
    .Q_N(_11537_),
    .Q(\top_ihp.oisc.regs[7][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1230),
    .D(_02432_),
    .Q_N(_11536_),
    .Q(\top_ihp.oisc.regs[7][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1234),
    .D(_02433_),
    .Q_N(_11535_),
    .Q(\top_ihp.oisc.regs[7][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1230),
    .D(_02434_),
    .Q_N(_11534_),
    .Q(\top_ihp.oisc.regs[7][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1183),
    .D(_02435_),
    .Q_N(_11533_),
    .Q(\top_ihp.oisc.regs[7][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1216),
    .D(_02436_),
    .Q_N(_11532_),
    .Q(\top_ihp.oisc.regs[8][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1166),
    .D(_02437_),
    .Q_N(_11531_),
    .Q(\top_ihp.oisc.regs[8][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1212),
    .D(_02438_),
    .Q_N(_11530_),
    .Q(\top_ihp.oisc.regs[8][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1176),
    .D(_02439_),
    .Q_N(_11529_),
    .Q(\top_ihp.oisc.regs[8][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1165),
    .D(_02440_),
    .Q_N(_11528_),
    .Q(\top_ihp.oisc.regs[8][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1210),
    .D(_02441_),
    .Q_N(_11527_),
    .Q(\top_ihp.oisc.regs[8][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1211),
    .D(_02442_),
    .Q_N(_11526_),
    .Q(\top_ihp.oisc.regs[8][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1218),
    .D(_02443_),
    .Q_N(_11525_),
    .Q(\top_ihp.oisc.regs[8][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1172),
    .D(_02444_),
    .Q_N(_11524_),
    .Q(\top_ihp.oisc.regs[8][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1170),
    .D(_02445_),
    .Q_N(_11523_),
    .Q(\top_ihp.oisc.regs[8][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1171),
    .D(_02446_),
    .Q_N(_11522_),
    .Q(\top_ihp.oisc.regs[8][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1182),
    .D(_02447_),
    .Q_N(_11521_),
    .Q(\top_ihp.oisc.regs[8][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1197),
    .D(_02448_),
    .Q_N(_11520_),
    .Q(\top_ihp.oisc.regs[8][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1186),
    .D(_02449_),
    .Q_N(_11519_),
    .Q(\top_ihp.oisc.regs[8][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1213),
    .D(_02450_),
    .Q_N(_11518_),
    .Q(\top_ihp.oisc.regs[8][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1171),
    .D(_02451_),
    .Q_N(_11517_),
    .Q(\top_ihp.oisc.regs[8][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1229),
    .D(_02452_),
    .Q_N(_11516_),
    .Q(\top_ihp.oisc.regs[8][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1170),
    .D(_02453_),
    .Q_N(_11515_),
    .Q(\top_ihp.oisc.regs[8][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1199),
    .D(_02454_),
    .Q_N(_11514_),
    .Q(\top_ihp.oisc.regs[8][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1189),
    .D(_02455_),
    .Q_N(_11513_),
    .Q(\top_ihp.oisc.regs[8][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1163),
    .D(_02456_),
    .Q_N(_11512_),
    .Q(\top_ihp.oisc.regs[8][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1203),
    .D(_02457_),
    .Q_N(_11511_),
    .Q(\top_ihp.oisc.regs[8][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1237),
    .D(_02458_),
    .Q_N(_11510_),
    .Q(\top_ihp.oisc.regs[8][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1161),
    .D(_02459_),
    .Q_N(_11509_),
    .Q(\top_ihp.oisc.regs[8][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1160),
    .D(_02460_),
    .Q_N(_11508_),
    .Q(\top_ihp.oisc.regs[8][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1163),
    .D(_02461_),
    .Q_N(_11507_),
    .Q(\top_ihp.oisc.regs[8][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1161),
    .D(_02462_),
    .Q_N(_11506_),
    .Q(\top_ihp.oisc.regs[8][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1161),
    .D(_02463_),
    .Q_N(_11505_),
    .Q(\top_ihp.oisc.regs[8][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1230),
    .D(_02464_),
    .Q_N(_11504_),
    .Q(\top_ihp.oisc.regs[8][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1236),
    .D(_02465_),
    .Q_N(_11503_),
    .Q(\top_ihp.oisc.regs[8][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1233),
    .D(_02466_),
    .Q_N(_11502_),
    .Q(\top_ihp.oisc.regs[8][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1215),
    .D(_02467_),
    .Q_N(_11501_),
    .Q(\top_ihp.oisc.regs[8][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1214),
    .D(_02468_),
    .Q_N(_11500_),
    .Q(\top_ihp.oisc.regs[9][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1166),
    .D(_02469_),
    .Q_N(_11499_),
    .Q(\top_ihp.oisc.regs[9][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1168),
    .D(_02470_),
    .Q_N(_11498_),
    .Q(\top_ihp.oisc.regs[9][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1175),
    .D(_02471_),
    .Q_N(_11497_),
    .Q(\top_ihp.oisc.regs[9][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1165),
    .D(_02472_),
    .Q_N(_11496_),
    .Q(\top_ihp.oisc.regs[9][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1211),
    .D(_02473_),
    .Q_N(_11495_),
    .Q(\top_ihp.oisc.regs[9][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1177),
    .D(_02474_),
    .Q_N(_11494_),
    .Q(\top_ihp.oisc.regs[9][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1210),
    .D(_02475_),
    .Q_N(_11493_),
    .Q(\top_ihp.oisc.regs[9][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1172),
    .D(_02476_),
    .Q_N(_11492_),
    .Q(\top_ihp.oisc.regs[9][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1180),
    .D(_02477_),
    .Q_N(_11491_),
    .Q(\top_ihp.oisc.regs[9][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1171),
    .D(_02478_),
    .Q_N(_11490_),
    .Q(\top_ihp.oisc.regs[9][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1182),
    .D(_02479_),
    .Q_N(_11489_),
    .Q(\top_ihp.oisc.regs[9][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1199),
    .D(_02480_),
    .Q_N(_11488_),
    .Q(\top_ihp.oisc.regs[9][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1186),
    .D(_02481_),
    .Q_N(_11487_),
    .Q(\top_ihp.oisc.regs[9][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1215),
    .D(_02482_),
    .Q_N(_11486_),
    .Q(\top_ihp.oisc.regs[9][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1183),
    .D(_02483_),
    .Q_N(_11485_),
    .Q(\top_ihp.oisc.regs[9][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1232),
    .D(_02484_),
    .Q_N(_11484_),
    .Q(\top_ihp.oisc.regs[9][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1179),
    .D(_02485_),
    .Q_N(_11483_),
    .Q(\top_ihp.oisc.regs[9][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1197),
    .D(_02486_),
    .Q_N(_11482_),
    .Q(\top_ihp.oisc.regs[9][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1186),
    .D(_02487_),
    .Q_N(_11481_),
    .Q(\top_ihp.oisc.regs[9][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1160),
    .D(_02488_),
    .Q_N(_11480_),
    .Q(\top_ihp.oisc.regs[9][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1161),
    .D(_02489_),
    .Q_N(_11479_),
    .Q(\top_ihp.oisc.regs[9][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1237),
    .D(_02490_),
    .Q_N(_11478_),
    .Q(\top_ihp.oisc.regs[9][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1160),
    .D(_02491_),
    .Q_N(_11477_),
    .Q(\top_ihp.oisc.regs[9][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1162),
    .D(_02492_),
    .Q_N(_11476_),
    .Q(\top_ihp.oisc.regs[9][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1194),
    .D(_02493_),
    .Q_N(_11475_),
    .Q(\top_ihp.oisc.regs[9][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1160),
    .D(_02494_),
    .Q_N(_11474_),
    .Q(\top_ihp.oisc.regs[9][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1160),
    .D(_02495_),
    .Q_N(_11473_),
    .Q(\top_ihp.oisc.regs[9][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1235),
    .D(_02496_),
    .Q_N(_11472_),
    .Q(\top_ihp.oisc.regs[9][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1234),
    .D(_02497_),
    .Q_N(_11471_),
    .Q(\top_ihp.oisc.regs[9][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1231),
    .D(_02498_),
    .Q_N(_11470_),
    .Q(\top_ihp.oisc.regs[9][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1215),
    .D(_02499_),
    .Q_N(_11469_),
    .Q(\top_ihp.oisc.regs[9][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1147),
    .D(_02500_),
    .Q_N(\top_ihp.oisc.state[0] ),
    .Q(_13600_));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1157),
    .D(_02501_),
    .Q_N(_11468_),
    .Q(\top_ihp.oisc.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1157),
    .D(_02502_),
    .Q_N(_00087_),
    .Q(\top_ihp.oisc.state[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1157),
    .D(_02503_),
    .Q_N(_00086_),
    .Q(\top_ihp.oisc.state[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1158),
    .D(_02504_),
    .Q_N(_00088_),
    .Q(\top_ihp.oisc.state[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[5]$_DFF_PN0_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1158),
    .D(_00002_),
    .Q_N(_00073_),
    .Q(\top_ihp.oisc.state[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1147),
    .D(_02505_),
    .Q_N(_11467_),
    .Q(\top_ihp.oisc.state[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1124),
    .D(_02506_),
    .Q_N(_00185_),
    .Q(\top_ihp.oisc.wb_dat_o[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1126),
    .D(_02507_),
    .Q_N(_11466_),
    .Q(\top_ihp.oisc.wb_dat_o[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1126),
    .D(_02508_),
    .Q_N(_11465_),
    .Q(\top_ihp.oisc.wb_dat_o[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1126),
    .D(_02509_),
    .Q_N(_11464_),
    .Q(\top_ihp.oisc.wb_dat_o[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1128),
    .D(_02510_),
    .Q_N(_11463_),
    .Q(\top_ihp.oisc.wb_dat_o[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1128),
    .D(_02511_),
    .Q_N(_11462_),
    .Q(\top_ihp.oisc.wb_dat_o[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1127),
    .D(_02512_),
    .Q_N(_11461_),
    .Q(\top_ihp.oisc.wb_dat_o[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1127),
    .D(_02513_),
    .Q_N(_11460_),
    .Q(\top_ihp.oisc.wb_dat_o[16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1128),
    .D(_02514_),
    .Q_N(_11459_),
    .Q(\top_ihp.oisc.wb_dat_o[17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1128),
    .D(_02515_),
    .Q_N(_11458_),
    .Q(\top_ihp.oisc.wb_dat_o[18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1128),
    .D(_02516_),
    .Q_N(_11457_),
    .Q(\top_ihp.oisc.wb_dat_o[19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1124),
    .D(_02517_),
    .Q_N(_00186_),
    .Q(\top_ihp.oisc.wb_dat_o[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1132),
    .D(_02518_),
    .Q_N(_11456_),
    .Q(\top_ihp.oisc.wb_dat_o[20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1132),
    .D(_02519_),
    .Q_N(_11455_),
    .Q(\top_ihp.oisc.wb_dat_o[21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1130),
    .D(_02520_),
    .Q_N(_11454_),
    .Q(\top_ihp.oisc.wb_dat_o[22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1128),
    .D(_02521_),
    .Q_N(_11453_),
    .Q(\top_ihp.oisc.wb_dat_o[23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1131),
    .D(_02522_),
    .Q_N(_11452_),
    .Q(\top_ihp.oisc.wb_dat_o[24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1132),
    .D(_02523_),
    .Q_N(_11451_),
    .Q(\top_ihp.oisc.wb_dat_o[25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1130),
    .D(_02524_),
    .Q_N(_11450_),
    .Q(\top_ihp.oisc.wb_dat_o[26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1133),
    .D(_02525_),
    .Q_N(_11449_),
    .Q(\top_ihp.oisc.wb_dat_o[27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1131),
    .D(_02526_),
    .Q_N(_11448_),
    .Q(\top_ihp.oisc.wb_dat_o[28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1130),
    .D(_02527_),
    .Q_N(_11447_),
    .Q(\top_ihp.oisc.wb_dat_o[29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1124),
    .D(_02528_),
    .Q_N(_00187_),
    .Q(\top_ihp.oisc.wb_dat_o[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1131),
    .D(_02529_),
    .Q_N(_11446_),
    .Q(\top_ihp.oisc.wb_dat_o[30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1133),
    .D(_02530_),
    .Q_N(_11445_),
    .Q(\top_ihp.oisc.wb_dat_o[31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1124),
    .D(_02531_),
    .Q_N(_00188_),
    .Q(\top_ihp.oisc.wb_dat_o[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1124),
    .D(_02532_),
    .Q_N(_00189_),
    .Q(\top_ihp.oisc.wb_dat_o[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1124),
    .D(_02533_),
    .Q_N(_00190_),
    .Q(\top_ihp.oisc.wb_dat_o[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1130),
    .D(_02534_),
    .Q_N(_00191_),
    .Q(\top_ihp.oisc.wb_dat_o[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1130),
    .D(_02535_),
    .Q_N(_00192_),
    .Q(\top_ihp.oisc.wb_dat_o[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1131),
    .D(_02536_),
    .Q_N(_11444_),
    .Q(\top_ihp.oisc.wb_dat_o[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1133),
    .D(_02537_),
    .Q_N(_13528_),
    .Q(\top_ihp.oisc.wb_dat_o[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.ack_o$_DFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1131),
    .D(_00003_),
    .Q_N(_11443_),
    .Q(\top_ihp.wb_ack_coproc ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1111),
    .D(_02538_),
    .Q_N(_11442_),
    .Q(\top_ihp.wb_coproc.dat_o[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1090),
    .D(_02539_),
    .Q_N(_11441_),
    .Q(\top_ihp.wb_coproc.dat_o[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1111),
    .D(_02540_),
    .Q_N(_11440_),
    .Q(\top_ihp.wb_coproc.dat_o[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1111),
    .D(_02541_),
    .Q_N(_11439_),
    .Q(\top_ihp.wb_coproc.dat_o[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1111),
    .D(_02542_),
    .Q_N(_11438_),
    .Q(\top_ihp.wb_coproc.dat_o[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1111),
    .D(_02543_),
    .Q_N(_11437_),
    .Q(\top_ihp.wb_coproc.dat_o[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1111),
    .D(_02544_),
    .Q_N(_11436_),
    .Q(\top_ihp.wb_coproc.dat_o[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1111),
    .D(_02545_),
    .Q_N(_11435_),
    .Q(\top_ihp.wb_coproc.dat_o[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1090),
    .D(_02546_),
    .Q_N(_11434_),
    .Q(\top_ihp.wb_coproc.dat_o[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1111),
    .D(_02547_),
    .Q_N(_11433_),
    .Q(\top_ihp.wb_coproc.dat_o[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1123),
    .D(_02548_),
    .Q_N(_11432_),
    .Q(\top_ihp.wb_coproc.dat_o[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1114),
    .D(_02549_),
    .Q_N(_11431_),
    .Q(\top_ihp.wb_coproc.dat_o[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1126),
    .D(_02550_),
    .Q_N(_11430_),
    .Q(\top_ihp.wb_coproc.dat_o[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1129),
    .D(_02551_),
    .Q_N(_11429_),
    .Q(\top_ihp.wb_coproc.dat_o[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1123),
    .D(_02552_),
    .Q_N(_11428_),
    .Q(\top_ihp.wb_coproc.dat_o[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1123),
    .D(_02553_),
    .Q_N(_11427_),
    .Q(\top_ihp.wb_coproc.dat_o[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1125),
    .D(_02554_),
    .Q_N(_11426_),
    .Q(\top_ihp.wb_coproc.dat_o[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1129),
    .D(_02555_),
    .Q_N(_11425_),
    .Q(\top_ihp.wb_coproc.dat_o[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1112),
    .D(_02556_),
    .Q_N(_11424_),
    .Q(\top_ihp.wb_coproc.dat_o[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1112),
    .D(_02557_),
    .Q_N(_11423_),
    .Q(\top_ihp.wb_coproc.dat_o[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1088),
    .D(_02558_),
    .Q_N(_11422_),
    .Q(\top_ihp.wb_coproc.dat_o[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1094),
    .D(_02559_),
    .Q_N(_11421_),
    .Q(\top_ihp.wb_coproc.dat_o[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1088),
    .D(_02560_),
    .Q_N(_11420_),
    .Q(\top_ihp.wb_coproc.dat_o[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1094),
    .D(_02561_),
    .Q_N(_11419_),
    .Q(\top_ihp.wb_coproc.dat_o[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1091),
    .D(_02562_),
    .Q_N(_11418_),
    .Q(\top_ihp.wb_coproc.dat_o[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1088),
    .D(_02563_),
    .Q_N(_11417_),
    .Q(\top_ihp.wb_coproc.dat_o[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1088),
    .D(_02564_),
    .Q_N(_11416_),
    .Q(\top_ihp.wb_coproc.dat_o[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1092),
    .D(_02565_),
    .Q_N(_11415_),
    .Q(\top_ihp.wb_coproc.dat_o[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1092),
    .D(_02566_),
    .Q_N(_11414_),
    .Q(\top_ihp.wb_coproc.dat_o[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1092),
    .D(_02567_),
    .Q_N(_11413_),
    .Q(\top_ihp.wb_coproc.dat_o[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1113),
    .D(_02568_),
    .Q_N(_11412_),
    .Q(\top_ihp.wb_coproc.dat_o[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1113),
    .D(_02569_),
    .Q_N(_11411_),
    .Q(\top_ihp.wb_coproc.dat_o[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1086),
    .D(_02570_),
    .Q_N(_11410_),
    .Q(\top_ihp.wb_coproc.opa[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1086),
    .D(_02571_),
    .Q_N(_11409_),
    .Q(\top_ihp.wb_coproc.opa[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1086),
    .D(_02572_),
    .Q_N(_11408_),
    .Q(\top_ihp.wb_coproc.opa[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1086),
    .D(_02573_),
    .Q_N(_11407_),
    .Q(\top_ihp.wb_coproc.opa[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1090),
    .D(_02574_),
    .Q_N(_11406_),
    .Q(\top_ihp.wb_coproc.opa[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1087),
    .D(_02575_),
    .Q_N(_11405_),
    .Q(\top_ihp.wb_coproc.opa[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1087),
    .D(_02576_),
    .Q_N(_11404_),
    .Q(\top_ihp.wb_coproc.opa[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1087),
    .D(_02577_),
    .Q_N(_11403_),
    .Q(\top_ihp.wb_coproc.opa[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1090),
    .D(_02578_),
    .Q_N(_11402_),
    .Q(\top_ihp.wb_coproc.opa[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1090),
    .D(_02579_),
    .Q_N(_11401_),
    .Q(\top_ihp.wb_coproc.opa[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1123),
    .D(_02580_),
    .Q_N(_11400_),
    .Q(\top_ihp.wb_coproc.opa[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1114),
    .D(_02581_),
    .Q_N(_11399_),
    .Q(\top_ihp.wb_coproc.opa[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1126),
    .D(_02582_),
    .Q_N(_11398_),
    .Q(\top_ihp.wb_coproc.opa[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1126),
    .D(_02583_),
    .Q_N(_11397_),
    .Q(\top_ihp.wb_coproc.opa[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1123),
    .D(_02584_),
    .Q_N(_11396_),
    .Q(\top_ihp.wb_coproc.opa[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1115),
    .D(_02585_),
    .Q_N(_11395_),
    .Q(\top_ihp.wb_coproc.opa[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1125),
    .D(_02586_),
    .Q_N(_11394_),
    .Q(\top_ihp.wb_coproc.opa[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1126),
    .D(_02587_),
    .Q_N(_11393_),
    .Q(\top_ihp.wb_coproc.opa[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1114),
    .D(_02588_),
    .Q_N(_11392_),
    .Q(\top_ihp.wb_coproc.opa[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1125),
    .D(_02589_),
    .Q_N(_11391_),
    .Q(\top_ihp.wb_coproc.opa[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1088),
    .D(_02590_),
    .Q_N(_11390_),
    .Q(\top_ihp.wb_coproc.opa[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1089),
    .D(_02591_),
    .Q_N(_11389_),
    .Q(\top_ihp.wb_coproc.opa[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1077),
    .D(_02592_),
    .Q_N(_11388_),
    .Q(\top_ihp.wb_coproc.opa[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1092),
    .D(_02593_),
    .Q_N(_11387_),
    .Q(\top_ihp.wb_coproc.opa[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1091),
    .D(_02594_),
    .Q_N(_11386_),
    .Q(\top_ihp.wb_coproc.opa[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1088),
    .D(_02595_),
    .Q_N(_11385_),
    .Q(\top_ihp.wb_coproc.opa[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1078),
    .D(_02596_),
    .Q_N(_11384_),
    .Q(\top_ihp.wb_coproc.opa[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1083),
    .D(_02597_),
    .Q_N(_11383_),
    .Q(\top_ihp.wb_coproc.opa[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1092),
    .D(_02598_),
    .Q_N(_11382_),
    .Q(\top_ihp.wb_coproc.opa[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1083),
    .D(_02599_),
    .Q_N(_11381_),
    .Q(\top_ihp.wb_coproc.opa[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1091),
    .D(_02600_),
    .Q_N(_11380_),
    .Q(\top_ihp.wb_coproc.opa[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1091),
    .D(_02601_),
    .Q_N(_11379_),
    .Q(\top_ihp.wb_coproc.opa[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1086),
    .D(_02602_),
    .Q_N(_11378_),
    .Q(\top_ihp.wb_coproc.opb[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1087),
    .D(_02603_),
    .Q_N(_11377_),
    .Q(\top_ihp.wb_coproc.opb[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1086),
    .D(_02604_),
    .Q_N(_11376_),
    .Q(\top_ihp.wb_coproc.opb[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1086),
    .D(_02605_),
    .Q_N(_11375_),
    .Q(\top_ihp.wb_coproc.opb[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1090),
    .D(_02606_),
    .Q_N(_11374_),
    .Q(\top_ihp.wb_coproc.opb[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1086),
    .D(_02607_),
    .Q_N(_11373_),
    .Q(\top_ihp.wb_coproc.opb[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1087),
    .D(_02608_),
    .Q_N(_11372_),
    .Q(\top_ihp.wb_coproc.opb[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1087),
    .D(_02609_),
    .Q_N(_11371_),
    .Q(\top_ihp.wb_coproc.opb[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1090),
    .D(_02610_),
    .Q_N(_11370_),
    .Q(\top_ihp.wb_coproc.opb[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1090),
    .D(_02611_),
    .Q_N(_11369_),
    .Q(\top_ihp.wb_coproc.opb[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1127),
    .D(_02612_),
    .Q_N(_11368_),
    .Q(\top_ihp.wb_coproc.opb[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1112),
    .D(_02613_),
    .Q_N(_11367_),
    .Q(\top_ihp.wb_coproc.opb[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1127),
    .D(_02614_),
    .Q_N(_11366_),
    .Q(\top_ihp.wb_coproc.opb[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1126),
    .D(_02615_),
    .Q_N(_11365_),
    .Q(\top_ihp.wb_coproc.opb[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1123),
    .D(_02616_),
    .Q_N(_11364_),
    .Q(\top_ihp.wb_coproc.opb[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1115),
    .D(_02617_),
    .Q_N(_11363_),
    .Q(\top_ihp.wb_coproc.opb[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1125),
    .D(_02618_),
    .Q_N(_11362_),
    .Q(\top_ihp.wb_coproc.opb[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1127),
    .D(_02619_),
    .Q_N(_11361_),
    .Q(\top_ihp.wb_coproc.opb[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1114),
    .D(_02620_),
    .Q_N(_11360_),
    .Q(\top_ihp.wb_coproc.opb[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1123),
    .D(_02621_),
    .Q_N(_11359_),
    .Q(\top_ihp.wb_coproc.opb[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1089),
    .D(_02622_),
    .Q_N(_11358_),
    .Q(\top_ihp.wb_coproc.opb[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1091),
    .D(_02623_),
    .Q_N(_11357_),
    .Q(\top_ihp.wb_coproc.opb[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1088),
    .D(_02624_),
    .Q_N(_11356_),
    .Q(\top_ihp.wb_coproc.opb[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1092),
    .D(_02625_),
    .Q_N(_11355_),
    .Q(\top_ihp.wb_coproc.opb[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1091),
    .D(_02626_),
    .Q_N(_11354_),
    .Q(\top_ihp.wb_coproc.opb[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1088),
    .D(_02627_),
    .Q_N(_11353_),
    .Q(\top_ihp.wb_coproc.opb[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1078),
    .D(_02628_),
    .Q_N(_11352_),
    .Q(\top_ihp.wb_coproc.opb[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1083),
    .D(_02629_),
    .Q_N(_11351_),
    .Q(\top_ihp.wb_coproc.opb[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1092),
    .D(_02630_),
    .Q_N(_11350_),
    .Q(\top_ihp.wb_coproc.opb[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1084),
    .D(_02631_),
    .Q_N(_11349_),
    .Q(\top_ihp.wb_coproc.opb[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1091),
    .D(_02632_),
    .Q_N(_11348_),
    .Q(\top_ihp.wb_coproc.opb[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1091),
    .D(_02633_),
    .Q_N(_11347_),
    .Q(\top_ihp.wb_coproc.opb[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1993),
    .D(_02634_),
    .Q_N(_00232_),
    .Q(\top_ihp.wb_emem.bit_counter[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1994),
    .D(_02635_),
    .Q_N(_11346_),
    .Q(\top_ihp.wb_emem.bit_counter[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1995),
    .D(_02636_),
    .Q_N(_11345_),
    .Q(\top_ihp.wb_emem.bit_counter[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1996),
    .D(_02637_),
    .Q_N(_11344_),
    .Q(\top_ihp.wb_emem.bit_counter[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1997),
    .D(_02638_),
    .Q_N(_11343_),
    .Q(\top_ihp.wb_emem.bit_counter[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1998),
    .D(_02639_),
    .Q_N(_11342_),
    .Q(\top_ihp.wb_emem.bit_counter[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1999),
    .D(_02640_),
    .Q_N(_11341_),
    .Q(\top_ihp.wb_emem.bit_counter[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2000),
    .D(_02641_),
    .Q_N(_11340_),
    .Q(\top_ihp.wb_emem.bit_counter[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[0]$_DFFE_NN0P_  (.CLK(net2131),
    .RESET_B(net1119),
    .D(_02642_),
    .Q_N(_00155_),
    .Q(\top_ihp.wb_dati_ram[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[10]$_DFFE_NN0P_  (.CLK(net2130),
    .RESET_B(net1119),
    .D(_02643_),
    .Q_N(_00122_),
    .Q(\top_ihp.wb_dati_ram[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[11]$_DFFE_NN0P_  (.CLK(net2129),
    .RESET_B(net1119),
    .D(_02644_),
    .Q_N(_00125_),
    .Q(\top_ihp.wb_dati_ram[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[12]$_DFFE_NN0P_  (.CLK(net2128),
    .RESET_B(net1120),
    .D(_02645_),
    .Q_N(_00143_),
    .Q(\top_ihp.wb_dati_ram[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[13]$_DFFE_NN0P_  (.CLK(net2127),
    .RESET_B(net1120),
    .D(_02646_),
    .Q_N(_00146_),
    .Q(\top_ihp.wb_dati_ram[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[14]$_DFFE_NN0P_  (.CLK(net2126),
    .RESET_B(net1120),
    .D(_02647_),
    .Q_N(_00149_),
    .Q(\top_ihp.wb_dati_ram[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[15]$_DFFE_NN0P_  (.CLK(net2125),
    .RESET_B(net1118),
    .D(_02648_),
    .Q_N(_00152_),
    .Q(\top_ihp.wb_dati_ram[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[16]$_DFFE_NN0P_  (.CLK(net2124),
    .RESET_B(net1118),
    .D(_02649_),
    .Q_N(_00131_),
    .Q(\top_ihp.wb_dati_ram[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[17]$_DFFE_NN0P_  (.CLK(net2123),
    .RESET_B(net1118),
    .D(_02650_),
    .Q_N(_00134_),
    .Q(\top_ihp.wb_dati_ram[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[18]$_DFFE_NN0P_  (.CLK(net2122),
    .RESET_B(net1118),
    .D(_02651_),
    .Q_N(_00137_),
    .Q(\top_ihp.wb_dati_ram[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[19]$_DFFE_NN0P_  (.CLK(net2121),
    .RESET_B(net1118),
    .D(_02652_),
    .Q_N(_00140_),
    .Q(\top_ihp.wb_dati_ram[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[1]$_DFFE_NN0P_  (.CLK(net2120),
    .RESET_B(net1118),
    .D(_02653_),
    .Q_N(_00158_),
    .Q(\top_ihp.wb_dati_ram[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[20]$_DFFE_NN0P_  (.CLK(net2119),
    .RESET_B(net1094),
    .D(_02654_),
    .Q_N(_00077_),
    .Q(\top_ihp.wb_dati_ram[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[21]$_DFFE_NN0P_  (.CLK(net2118),
    .RESET_B(net1094),
    .D(_02655_),
    .Q_N(_00083_),
    .Q(\top_ihp.wb_dati_ram[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[22]$_DFFE_NN0P_  (.CLK(net2117),
    .RESET_B(net1118),
    .D(_02656_),
    .Q_N(_00080_),
    .Q(\top_ihp.wb_dati_ram[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[23]$_DFFE_NN0P_  (.CLK(net2116),
    .RESET_B(net1095),
    .D(_02657_),
    .Q_N(_00113_),
    .Q(\top_ihp.wb_dati_ram[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[24]$_DFFE_NN0P_  (.CLK(net2115),
    .RESET_B(net1119),
    .D(_02658_),
    .Q_N(_11339_),
    .Q(\top_ihp.wb_dati_ram[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[25]$_DFFE_NN0P_  (.CLK(net2114),
    .RESET_B(net1119),
    .D(_02659_),
    .Q_N(_00194_),
    .Q(\top_ihp.wb_dati_ram[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[26]$_DFFE_NN0P_  (.CLK(net2113),
    .RESET_B(net1094),
    .D(_02660_),
    .Q_N(_00095_),
    .Q(\top_ihp.wb_dati_ram[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[27]$_DFFE_NN0P_  (.CLK(net2112),
    .RESET_B(net1094),
    .D(_02661_),
    .Q_N(_00101_),
    .Q(\top_ihp.wb_dati_ram[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[28]$_DFFE_NN0P_  (.CLK(net2111),
    .RESET_B(net1094),
    .D(_02662_),
    .Q_N(_00098_),
    .Q(\top_ihp.wb_dati_ram[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[29]$_DFFE_NN0P_  (.CLK(net2110),
    .RESET_B(net1094),
    .D(_02663_),
    .Q_N(_00104_),
    .Q(\top_ihp.wb_dati_ram[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[2]$_DFFE_NN0P_  (.CLK(net2109),
    .RESET_B(net1095),
    .D(_02664_),
    .Q_N(_00161_),
    .Q(\top_ihp.wb_dati_ram[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[30]$_DFFE_NN0P_  (.CLK(net2108),
    .RESET_B(net1095),
    .D(_02665_),
    .Q_N(_00107_),
    .Q(\top_ihp.wb_dati_ram[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[31]$_DFFE_NN0P_  (.CLK(net2107),
    .RESET_B(net1095),
    .D(_02666_),
    .Q_N(_00128_),
    .Q(\top_ihp.wb_dati_ram[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[32]$_DFFE_NN0P_  (.CLK(net2106),
    .RESET_B(net1104),
    .D(_02667_),
    .Q_N(_11338_),
    .Q(\top_ihp.wb_emem.cmd[32] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[33]$_DFFE_NN0P_  (.CLK(net2105),
    .RESET_B(net1104),
    .D(_02668_),
    .Q_N(_11337_),
    .Q(\top_ihp.wb_emem.cmd[33] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[34]$_DFFE_NN0P_  (.CLK(net2104),
    .RESET_B(net1104),
    .D(_02669_),
    .Q_N(_11336_),
    .Q(\top_ihp.wb_emem.cmd[34] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[35]$_DFFE_NN0P_  (.CLK(net2103),
    .RESET_B(net1104),
    .D(_02670_),
    .Q_N(_11335_),
    .Q(\top_ihp.wb_emem.cmd[35] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[36]$_DFFE_NN0P_  (.CLK(net2102),
    .RESET_B(net1104),
    .D(_02671_),
    .Q_N(_11334_),
    .Q(\top_ihp.wb_emem.cmd[36] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[37]$_DFFE_NN0P_  (.CLK(net2101),
    .RESET_B(net1105),
    .D(_02672_),
    .Q_N(_11333_),
    .Q(\top_ihp.wb_emem.cmd[37] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[38]$_DFFE_NN0P_  (.CLK(net2100),
    .RESET_B(net1105),
    .D(_02673_),
    .Q_N(_11332_),
    .Q(\top_ihp.wb_emem.cmd[38] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[39]$_DFFE_NN0P_  (.CLK(net2099),
    .RESET_B(net1105),
    .D(_02674_),
    .Q_N(_11331_),
    .Q(\top_ihp.wb_emem.cmd[39] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[3]$_DFFE_NN0P_  (.CLK(net2098),
    .RESET_B(net1095),
    .D(_02675_),
    .Q_N(_00164_),
    .Q(\top_ihp.wb_dati_ram[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[40]$_DFFE_NN0P_  (.CLK(net2097),
    .RESET_B(net1105),
    .D(_02676_),
    .Q_N(_11330_),
    .Q(\top_ihp.wb_emem.cmd[40] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[41]$_DFFE_NN0P_  (.CLK(net2096),
    .RESET_B(net1134),
    .D(_02677_),
    .Q_N(_11329_),
    .Q(\top_ihp.wb_emem.cmd[41] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[42]$_DFFE_NN0P_  (.CLK(net2095),
    .RESET_B(net1134),
    .D(_02678_),
    .Q_N(_11328_),
    .Q(\top_ihp.wb_emem.cmd[42] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[43]$_DFFE_NN0P_  (.CLK(net2094),
    .RESET_B(net1136),
    .D(_02679_),
    .Q_N(_11327_),
    .Q(\top_ihp.wb_emem.cmd[43] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[44]$_DFFE_NN0P_  (.CLK(net2093),
    .RESET_B(net1120),
    .D(_02680_),
    .Q_N(_11326_),
    .Q(\top_ihp.wb_emem.cmd[44] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[45]$_DFFE_NN0P_  (.CLK(net2092),
    .RESET_B(net1120),
    .D(_02681_),
    .Q_N(_11325_),
    .Q(\top_ihp.wb_emem.cmd[45] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[46]$_DFFE_NN0P_  (.CLK(net2091),
    .RESET_B(net1120),
    .D(_02682_),
    .Q_N(_11324_),
    .Q(\top_ihp.wb_emem.cmd[46] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[47]$_DFFE_NN0P_  (.CLK(net2090),
    .RESET_B(net1136),
    .D(_02683_),
    .Q_N(_11323_),
    .Q(\top_ihp.wb_emem.cmd[47] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[48]$_DFFE_NN1P_  (.CLK(net2089),
    .RESET_B(net1122),
    .D(_02684_),
    .Q_N(\top_ihp.wb_emem.cmd[48] ),
    .Q(_00308_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[49]$_DFFE_NN0P_  (.CLK(net2088),
    .RESET_B(net1120),
    .D(_02685_),
    .Q_N(_11322_),
    .Q(\top_ihp.wb_emem.cmd[49] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[4]$_DFFE_NN0P_  (.CLK(net2087),
    .RESET_B(net1093),
    .D(_02686_),
    .Q_N(_00167_),
    .Q(\top_ihp.wb_dati_ram[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[50]$_DFFE_NN0P_  (.CLK(net2086),
    .RESET_B(net1120),
    .D(_02687_),
    .Q_N(_11321_),
    .Q(\top_ihp.wb_emem.cmd[50] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[51]$_DFFE_NN1P_  (.CLK(net2085),
    .RESET_B(net1104),
    .D(_02688_),
    .Q_N(\top_ihp.wb_emem.cmd[51] ),
    .Q(_00309_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[52]$_DFFE_NN1P_  (.CLK(net2084),
    .RESET_B(net1106),
    .D(_02689_),
    .Q_N(\top_ihp.wb_emem.cmd[52] ),
    .Q(_00310_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[53]$_DFFE_NN0P_  (.CLK(net2083),
    .RESET_B(net1106),
    .D(_02690_),
    .Q_N(_11320_),
    .Q(\top_ihp.wb_emem.cmd[53] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[54]$_DFFE_NN0P_  (.CLK(net2082),
    .RESET_B(net1106),
    .D(_02691_),
    .Q_N(_11319_),
    .Q(\top_ihp.wb_emem.cmd[54] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[55]$_DFFE_NN1P_  (.CLK(net2081),
    .RESET_B(net1104),
    .D(_02692_),
    .Q_N(\top_ihp.wb_emem.cmd[55] ),
    .Q(_00311_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[56]$_DFFE_NN0P_  (.CLK(net2080),
    .RESET_B(net1104),
    .D(_02693_),
    .Q_N(_11318_),
    .Q(\top_ihp.wb_emem.cmd[56] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[57]$_DFFE_NN1P_  (.CLK(net2079),
    .RESET_B(net1103),
    .D(_02694_),
    .Q_N(\top_ihp.wb_emem.cmd[57] ),
    .Q(_00312_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[58]$_DFFE_NN1P_  (.CLK(net2078),
    .RESET_B(net1103),
    .D(_02695_),
    .Q_N(\top_ihp.wb_emem.cmd[58] ),
    .Q(_00313_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[59]$_DFFE_NN0P_  (.CLK(net2077),
    .RESET_B(net1103),
    .D(_02696_),
    .Q_N(_11317_),
    .Q(\top_ihp.wb_emem.cmd[59] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[5]$_DFFE_NN0P_  (.CLK(net2076),
    .RESET_B(net1092),
    .D(_02697_),
    .Q_N(_00170_),
    .Q(\top_ihp.wb_dati_ram[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[60]$_DFFE_NN0P_  (.CLK(net2075),
    .RESET_B(net1105),
    .D(_02698_),
    .Q_N(_11316_),
    .Q(\top_ihp.wb_emem.cmd[60] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[61]$_DFFE_NN1P_  (.CLK(net2074),
    .RESET_B(net1102),
    .D(_02699_),
    .Q_N(\top_ihp.wb_emem.cmd[61] ),
    .Q(_00314_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[62]$_DFFE_NN1P_  (.CLK(net2073),
    .RESET_B(net1102),
    .D(_02700_),
    .Q_N(\top_ihp.wb_emem.cmd[62] ),
    .Q(_00315_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[63]$_DFFE_NN0P_  (.CLK(net2072),
    .RESET_B(net1102),
    .D(_02701_),
    .Q_N(_11315_),
    .Q(\top_ihp.wb_emem.cmd[63] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[6]$_DFFE_NN0P_  (.CLK(net2071),
    .RESET_B(net1093),
    .D(_02702_),
    .Q_N(_00110_),
    .Q(\top_ihp.wb_dati_ram[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[7]$_DFFE_NN0P_  (.CLK(net2070),
    .RESET_B(net1095),
    .D(_02703_),
    .Q_N(_00173_),
    .Q(\top_ihp.wb_dati_ram[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[8]$_DFFE_NN0P_  (.CLK(net2069),
    .RESET_B(net1095),
    .D(_02704_),
    .Q_N(_00116_),
    .Q(\top_ihp.wb_dati_ram[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[9]$_DFFE_NN0P_  (.CLK(net2068),
    .RESET_B(net1095),
    .D(_02705_),
    .Q_N(_00119_),
    .Q(\top_ihp.wb_dati_ram[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.last_bit$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2001),
    .D(_02706_),
    .Q_N(_11314_),
    .Q(\top_ihp.wb_emem.last_bit ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.last_wait$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2002),
    .D(_02707_),
    .Q_N(_11313_),
    .Q(\top_ihp.wb_emem.last_wait ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.nbits[3]$_SDFFCE_NP1P_  (.CLK(net2067),
    .RESET_B(net2003),
    .D(_02708_),
    .Q_N(_11312_),
    .Q(\top_ihp.wb_emem.nbits[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.nbits[4]$_SDFFCE_NP0P_  (.CLK(net2066),
    .RESET_B(net2004),
    .D(_02709_),
    .Q_N(_11311_),
    .Q(\top_ihp.wb_emem.nbits[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.nbits[5]$_SDFFCE_NP0P_  (.CLK(net2065),
    .RESET_B(net2005),
    .D(_02710_),
    .Q_N(_11310_),
    .Q(\top_ihp.wb_emem.nbits[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.nbits[6]$_SDFFCE_NP0P_  (.CLK(net2064),
    .RESET_B(net2006),
    .D(_02711_),
    .Q_N(_11309_),
    .Q(\top_ihp.wb_emem.nbits[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.state[0]$_DFFE_NN0P_  (.CLK(net2063),
    .RESET_B(net1103),
    .D(_02712_),
    .Q_N(_11308_),
    .Q(\top_ihp.wb_emem.state[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.state[1]$_DFFE_NN0P_  (.CLK(net2062),
    .RESET_B(net1103),
    .D(_02713_),
    .Q_N(_11307_),
    .Q(\top_ihp.wb_emem.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.state[2]$_DFFE_NN0P_  (.CLK(net2061),
    .RESET_B(net1103),
    .D(_02714_),
    .Q_N(_11306_),
    .Q(\top_ihp.wb_emem.state[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.state[3]$_DFFE_NN0P_  (.CLK(net2060),
    .RESET_B(net1103),
    .D(_02715_),
    .Q_N(\top_ihp.ram_cs_o ),
    .Q(\top_ihp.wb_emem.state[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net2007),
    .D(_02716_),
    .Q_N(_00233_),
    .Q(\top_ihp.wb_emem.wait_counter[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2008),
    .D(_02717_),
    .Q_N(_11305_),
    .Q(\top_ihp.wb_emem.wait_counter[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2009),
    .D(_02718_),
    .Q_N(_11304_),
    .Q(\top_ihp.wb_emem.wait_counter[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2010),
    .D(_02719_),
    .Q_N(_11303_),
    .Q(\top_ihp.wb_emem.wait_counter[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2011),
    .D(_02720_),
    .Q_N(_11302_),
    .Q(\top_ihp.wb_emem.wait_counter[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2012),
    .D(_02721_),
    .Q_N(_11301_),
    .Q(\top_ihp.wb_emem.wait_counter[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2013),
    .D(_02722_),
    .Q_N(_11300_),
    .Q(\top_ihp.wb_emem.wait_counter[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net2014),
    .D(_02723_),
    .Q_N(_13529_),
    .Q(\top_ihp.wb_emem.wait_counter[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.ack_o$_DFF_PN0_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1106),
    .D(_00004_),
    .Q_N(_00089_),
    .Q(\top_ihp.wb_ack_gpio ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.dat_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1106),
    .D(_02724_),
    .Q_N(_11299_),
    .Q(\top_ihp.wb_dati_gpio[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1109),
    .D(_02725_),
    .Q_N(_11298_),
    .Q(\top_ihp.gpio_o_1 ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.data_o[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1110),
    .D(_02726_),
    .Q_N(\top_ihp.gpio_o_2 ),
    .Q(_00316_));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1140),
    .D(_02727_),
    .Q_N(_11297_),
    .Q(\top_ihp.gpio_o_3 ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.data_o[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1140),
    .D(_02728_),
    .Q_N(\top_ihp.gpio_o_4 ),
    .Q(_00317_));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[0]$_DFFE_NN0P_  (.CLK(net2059),
    .RESET_B(net1140),
    .D(_02729_),
    .Q_N(_11296_),
    .Q(\top_ihp.wb_imem.bits_left[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[1]$_DFFE_NN0P_  (.CLK(net2058),
    .RESET_B(net1141),
    .D(_02730_),
    .Q_N(_11295_),
    .Q(\top_ihp.wb_imem.bits_left[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[2]$_DFFE_NN0P_  (.CLK(net2057),
    .RESET_B(net1140),
    .D(_02731_),
    .Q_N(_11294_),
    .Q(\top_ihp.wb_imem.bits_left[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[3]$_DFFE_NN0P_  (.CLK(net2056),
    .RESET_B(net1142),
    .D(_02732_),
    .Q_N(_11293_),
    .Q(\top_ihp.wb_imem.bits_left[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[4]$_DFFE_NN0P_  (.CLK(net2055),
    .RESET_B(net1142),
    .D(_02733_),
    .Q_N(_11292_),
    .Q(\top_ihp.wb_imem.bits_left[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[5]$_DFFE_NN0P_  (.CLK(net2054),
    .RESET_B(net1142),
    .D(_02734_),
    .Q_N(_11291_),
    .Q(\top_ihp.wb_imem.bits_left[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[0]$_DFFE_NN0P_  (.CLK(net2053),
    .RESET_B(net1136),
    .D(_02735_),
    .Q_N(_00154_),
    .Q(\top_ihp.wb_dati_rom[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[10]$_DFFE_NN0P_  (.CLK(net2052),
    .RESET_B(net1134),
    .D(_02736_),
    .Q_N(_00121_),
    .Q(\top_ihp.wb_dati_rom[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[11]$_DFFE_NN0P_  (.CLK(net2051),
    .RESET_B(net1136),
    .D(_02737_),
    .Q_N(_00124_),
    .Q(\top_ihp.wb_dati_rom[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[12]$_DFFE_NN0P_  (.CLK(net2050),
    .RESET_B(net1136),
    .D(_02738_),
    .Q_N(_00142_),
    .Q(\top_ihp.wb_dati_rom[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[13]$_DFFE_NN0P_  (.CLK(net2049),
    .RESET_B(net1136),
    .D(_02739_),
    .Q_N(_00145_),
    .Q(\top_ihp.wb_dati_rom[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[14]$_DFFE_NN0P_  (.CLK(net2048),
    .RESET_B(net1136),
    .D(_02740_),
    .Q_N(_00148_),
    .Q(\top_ihp.wb_dati_rom[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[15]$_DFFE_NN0P_  (.CLK(net2047),
    .RESET_B(net1136),
    .D(_02741_),
    .Q_N(_00151_),
    .Q(\top_ihp.wb_dati_rom[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[16]$_DFFE_NN0P_  (.CLK(net2046),
    .RESET_B(net1137),
    .D(_02742_),
    .Q_N(_00130_),
    .Q(\top_ihp.wb_dati_rom[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[17]$_DFFE_NN0P_  (.CLK(net2045),
    .RESET_B(net1137),
    .D(_02743_),
    .Q_N(_00133_),
    .Q(\top_ihp.wb_dati_rom[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[18]$_DFFE_NN0P_  (.CLK(net2044),
    .RESET_B(net1134),
    .D(_02744_),
    .Q_N(_00136_),
    .Q(\top_ihp.wb_dati_rom[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[19]$_DFFE_NN0P_  (.CLK(net2043),
    .RESET_B(net1134),
    .D(_02745_),
    .Q_N(_00139_),
    .Q(\top_ihp.wb_dati_rom[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[1]$_DFFE_NN0P_  (.CLK(net2042),
    .RESET_B(net1137),
    .D(_02746_),
    .Q_N(_00157_),
    .Q(\top_ihp.wb_dati_rom[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[20]$_DFFE_NN0P_  (.CLK(net2041),
    .RESET_B(net1137),
    .D(_02747_),
    .Q_N(_00076_),
    .Q(\top_ihp.wb_dati_rom[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[21]$_DFFE_NN0P_  (.CLK(net2040),
    .RESET_B(net1141),
    .D(_02748_),
    .Q_N(_00082_),
    .Q(\top_ihp.wb_dati_rom[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[22]$_DFFE_NN0P_  (.CLK(net2039),
    .RESET_B(net1139),
    .D(_02749_),
    .Q_N(_00079_),
    .Q(\top_ihp.wb_dati_rom[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[23]$_DFFE_NN0P_  (.CLK(net2038),
    .RESET_B(net1135),
    .D(_02750_),
    .Q_N(_00112_),
    .Q(\top_ihp.wb_dati_rom[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[24]$_DFFE_NN0P_  (.CLK(net2037),
    .RESET_B(net1139),
    .D(_02751_),
    .Q_N(_11290_),
    .Q(\top_ihp.wb_dati_rom[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[25]$_DFFE_NN0P_  (.CLK(net2036),
    .RESET_B(net1139),
    .D(_02752_),
    .Q_N(_00193_),
    .Q(\top_ihp.wb_dati_rom[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[26]$_DFFE_NN0P_  (.CLK(net2035),
    .RESET_B(net1139),
    .D(_02753_),
    .Q_N(_00094_),
    .Q(\top_ihp.wb_dati_rom[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[27]$_DFFE_NN0P_  (.CLK(net2034),
    .RESET_B(net1139),
    .D(_02754_),
    .Q_N(_00100_),
    .Q(\top_ihp.wb_dati_rom[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[28]$_DFFE_NN0P_  (.CLK(net2033),
    .RESET_B(net1139),
    .D(_02755_),
    .Q_N(_00097_),
    .Q(\top_ihp.wb_dati_rom[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[29]$_DFFE_NN0P_  (.CLK(net2032),
    .RESET_B(net1139),
    .D(_02756_),
    .Q_N(_00103_),
    .Q(\top_ihp.wb_dati_rom[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[2]$_DFFE_NN0P_  (.CLK(net2031),
    .RESET_B(net1134),
    .D(_02757_),
    .Q_N(_00160_),
    .Q(\top_ihp.wb_dati_rom[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[30]$_DFFE_NN0P_  (.CLK(net2030),
    .RESET_B(net1139),
    .D(_02758_),
    .Q_N(_00106_),
    .Q(\top_ihp.wb_dati_rom[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[31]$_DFFE_NN0P_  (.CLK(net2029),
    .RESET_B(net1140),
    .D(_02759_),
    .Q_N(_00127_),
    .Q(\top_ihp.wb_dati_rom[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[3]$_DFFE_NN0P_  (.CLK(net2028),
    .RESET_B(net1135),
    .D(_02760_),
    .Q_N(_00163_),
    .Q(\top_ihp.wb_dati_rom[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[4]$_DFFE_NN0P_  (.CLK(net2027),
    .RESET_B(net1135),
    .D(_02761_),
    .Q_N(_00166_),
    .Q(\top_ihp.wb_dati_rom[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[5]$_DFFE_NN0P_  (.CLK(net2026),
    .RESET_B(net1137),
    .D(_02762_),
    .Q_N(_00169_),
    .Q(\top_ihp.wb_dati_rom[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[6]$_DFFE_NN0P_  (.CLK(net2025),
    .RESET_B(net1137),
    .D(_02763_),
    .Q_N(_00109_),
    .Q(\top_ihp.wb_dati_rom[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[7]$_DFFE_NN0P_  (.CLK(net2024),
    .RESET_B(net1135),
    .D(_02764_),
    .Q_N(_00172_),
    .Q(\top_ihp.wb_dati_rom[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[8]$_DFFE_NN0P_  (.CLK(net2023),
    .RESET_B(net1134),
    .D(_02765_),
    .Q_N(_00115_),
    .Q(\top_ihp.wb_dati_rom[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[9]$_DFFE_NN0P_  (.CLK(net2022),
    .RESET_B(net1134),
    .D(_02766_),
    .Q_N(_00118_),
    .Q(\top_ihp.wb_dati_rom[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.spi_cs_o$_DFFE_NN1P_  (.CLK(net2021),
    .RESET_B(net1140),
    .D(_02767_),
    .Q_N(\top_ihp.rom_cs_o ),
    .Q(_00318_));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.state[0]$_DFF_NN1_  (.CLK(net2020),
    .RESET_B(net1140),
    .D(_00323_),
    .Q_N(\top_ihp.wb_imem.state[0] ),
    .Q(_13601_));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.state[1]$_DFF_NN0_  (.CLK(net2019),
    .RESET_B(net1141),
    .D(_00000_),
    .Q_N(_00090_),
    .Q(\top_ihp.wb_imem.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.state[2]$_DFF_NN0_  (.CLK(net2018),
    .RESET_B(net1142),
    .D(_00001_),
    .Q_N(_13530_),
    .Q(\top_ihp.wb_imem.state[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.ack_o$_DFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1131),
    .D(_13604_),
    .Q_N(_11289_),
    .Q(\top_ihp.wb_ack_spi ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1130),
    .D(_02768_),
    .Q_N(_11288_),
    .Q(\top_ihp.wb_spi.bits_left[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1132),
    .D(_02769_),
    .Q_N(_11287_),
    .Q(\top_ihp.wb_spi.bits_left[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1132),
    .D(_02770_),
    .Q_N(_11286_),
    .Q(\top_ihp.wb_spi.bits_left[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1121),
    .D(_02771_),
    .Q_N(_11285_),
    .Q(\top_ihp.wb_spi.bits_left[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1121),
    .D(_02772_),
    .Q_N(_11284_),
    .Q(\top_ihp.wb_spi.bits_left[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1130),
    .D(_02773_),
    .Q_N(_11283_),
    .Q(\top_ihp.wb_spi.bits_left[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1116),
    .D(_02774_),
    .Q_N(_11282_),
    .Q(\top_ihp.wb_dati_spi[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1113),
    .D(_02775_),
    .Q_N(_00138_),
    .Q(\top_ihp.wb_dati_spi[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1113),
    .D(_02776_),
    .Q_N(_00141_),
    .Q(\top_ihp.wb_dati_spi[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1113),
    .D(_02777_),
    .Q_N(_00078_),
    .Q(\top_ihp.wb_dati_spi[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1112),
    .D(_02778_),
    .Q_N(_00084_),
    .Q(\top_ihp.wb_dati_spi[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1112),
    .D(_02779_),
    .Q_N(_00081_),
    .Q(\top_ihp.wb_dati_spi[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1114),
    .D(_02780_),
    .Q_N(_00114_),
    .Q(\top_ihp.wb_dati_spi[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1114),
    .D(_02781_),
    .Q_N(_00117_),
    .Q(\top_ihp.wb_dati_spi[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1114),
    .D(_02782_),
    .Q_N(_00120_),
    .Q(\top_ihp.wb_dati_spi[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1114),
    .D(_02783_),
    .Q_N(_00123_),
    .Q(\top_ihp.wb_dati_spi[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1115),
    .D(_02784_),
    .Q_N(_00126_),
    .Q(\top_ihp.wb_dati_spi[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1116),
    .D(_02785_),
    .Q_N(_00195_),
    .Q(\top_ihp.wb_dati_spi[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1115),
    .D(_02786_),
    .Q_N(_00144_),
    .Q(\top_ihp.wb_dati_spi[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1115),
    .D(_02787_),
    .Q_N(_00147_),
    .Q(\top_ihp.wb_dati_spi[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1124),
    .D(_02788_),
    .Q_N(_00150_),
    .Q(\top_ihp.wb_dati_spi[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1123),
    .D(_02789_),
    .Q_N(_00153_),
    .Q(\top_ihp.wb_dati_spi[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1124),
    .D(_02790_),
    .Q_N(_00156_),
    .Q(\top_ihp.wb_dati_spi[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1116),
    .D(_02791_),
    .Q_N(_00159_),
    .Q(\top_ihp.wb_dati_spi[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1116),
    .D(_02792_),
    .Q_N(_00162_),
    .Q(\top_ihp.wb_dati_spi[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1130),
    .D(_02793_),
    .Q_N(_00165_),
    .Q(\top_ihp.wb_dati_spi[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1116),
    .D(_02794_),
    .Q_N(_00168_),
    .Q(\top_ihp.wb_dati_spi[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1121),
    .D(_02795_),
    .Q_N(_00171_),
    .Q(\top_ihp.wb_dati_spi[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1116),
    .D(_02796_),
    .Q_N(_00096_),
    .Q(\top_ihp.wb_dati_spi[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1121),
    .D(_02797_),
    .Q_N(_00111_),
    .Q(\top_ihp.wb_dati_spi[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1121),
    .D(_02798_),
    .Q_N(_00174_),
    .Q(\top_ihp.wb_dati_spi[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1117),
    .D(_02799_),
    .Q_N(_00102_),
    .Q(\top_ihp.wb_dati_spi[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1117),
    .D(_02800_),
    .Q_N(_00099_),
    .Q(\top_ihp.wb_dati_spi[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1121),
    .D(_02801_),
    .Q_N(_00105_),
    .Q(\top_ihp.wb_dati_spi[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1121),
    .D(_02802_),
    .Q_N(_00108_),
    .Q(\top_ihp.wb_dati_spi[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1118),
    .D(_02803_),
    .Q_N(_00129_),
    .Q(\top_ihp.wb_dati_spi[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1113),
    .D(_02804_),
    .Q_N(_00132_),
    .Q(\top_ihp.wb_dati_spi[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1113),
    .D(_02805_),
    .Q_N(_00135_),
    .Q(\top_ihp.wb_dati_spi[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_clk_cnt[0]$_DFF_NN0_  (.CLK(net2017),
    .RESET_B(net1093),
    .D(_11255_),
    .Q_N(_11255_),
    .Q(\top_ihp.wb_spi.spi_clk_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_clk_cnt[1]$_DFF_NN0_  (.CLK(net2016),
    .RESET_B(net1093),
    .D(_00234_),
    .Q_N(_11281_),
    .Q(\top_ihp.spi_clk_o ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_cs_o_1$_DFFE_PN1P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1105),
    .D(_02806_),
    .Q_N(\top_ihp.spi_cs_o_1 ),
    .Q(_00319_));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_cs_o_2$_DFFE_PN1P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1105),
    .D(_02807_),
    .Q_N(\top_ihp.spi_cs_o_2 ),
    .Q(_00320_));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_cs_o_3$_DFFE_PN1P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1105),
    .D(_02808_),
    .Q_N(\top_ihp.spi_cs_o_3 ),
    .Q(_00321_));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.state$_DFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1132),
    .D(_13605_),
    .Q_N(_00091_),
    .Q(\top_ihp.wb_spi.state ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.ack_o$_SDFFCE_PP0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2015),
    .D(_02809_),
    .Q_N(_00075_),
    .Q(\top_ihp.wb_ack_uart ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.state[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1084),
    .D(_02810_),
    .Q_N(_11280_),
    .Q(\top_ihp.wb_uart.state[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.state[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1084),
    .D(_02811_),
    .Q_N(_11279_),
    .Q(\top_ihp.wb_uart.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.bit_cnt[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1101),
    .D(_02812_),
    .Q_N(_00183_),
    .Q(\top_ihp.wb_uart.uart_rx.bit_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.bit_cnt[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1101),
    .D(_02813_),
    .Q_N(_11278_),
    .Q(\top_ihp.wb_uart.uart_rx.bit_cnt[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.bit_cnt[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1101),
    .D(_02814_),
    .Q_N(_11277_),
    .Q(\top_ihp.wb_uart.uart_rx.bit_cnt[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.bit_cnt[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1101),
    .D(_02815_),
    .Q_N(_13531_),
    .Q(\top_ihp.wb_uart.uart_rx.bit_cnt[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[0]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1080),
    .D(_00005_),
    .Q_N(_13532_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[10]$_DFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1082),
    .D(_00006_),
    .Q_N(_13533_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[11]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1082),
    .D(_00007_),
    .Q_N(_13534_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[12]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1082),
    .D(_00008_),
    .Q_N(_13535_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[13]$_DFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1100),
    .D(_00009_),
    .Q_N(_13536_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[14]$_DFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1100),
    .D(_00010_),
    .Q_N(_13537_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[15]$_DFF_PN0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1100),
    .D(_00011_),
    .Q_N(_13538_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[16]$_DFF_PN0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1100),
    .D(_00012_),
    .Q_N(_13539_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[17]$_DFF_PN0_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1099),
    .D(_00013_),
    .Q_N(_13540_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[18]$_DFF_PN0_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1099),
    .D(_00014_),
    .Q_N(_13541_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[19]$_DFF_PN0_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1099),
    .D(_00015_),
    .Q_N(_13542_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[1]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1080),
    .D(_00016_),
    .Q_N(_13543_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[20]$_DFF_PN0_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1099),
    .D(_00017_),
    .Q_N(_13544_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[21]$_DFF_PN0_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1099),
    .D(_00018_),
    .Q_N(_13545_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[22]$_DFF_PN0_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1101),
    .D(_00019_),
    .Q_N(_13546_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[23]$_DFF_PN0_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1099),
    .D(_00020_),
    .Q_N(_13547_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[24]$_DFF_PN0_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1099),
    .D(_00021_),
    .Q_N(_13548_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[25]$_DFF_PN0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1099),
    .D(_00022_),
    .Q_N(_13549_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[26]$_DFF_PN0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1100),
    .D(_00023_),
    .Q_N(_13550_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[27]$_DFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1100),
    .D(_00024_),
    .Q_N(_13551_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[28]$_DFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1100),
    .D(_00025_),
    .Q_N(_13552_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[29]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1082),
    .D(_00026_),
    .Q_N(_13553_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[2]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1080),
    .D(_00027_),
    .Q_N(_13554_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[30]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1082),
    .D(_00028_),
    .Q_N(_13555_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[31]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1085),
    .D(_00029_),
    .Q_N(_13556_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[3]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1081),
    .D(_00030_),
    .Q_N(_13557_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[4]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1080),
    .D(_00031_),
    .Q_N(_13558_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[5]$_DFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1082),
    .D(_00032_),
    .Q_N(_00092_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[6]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1080),
    .D(_00033_),
    .Q_N(_13559_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[7]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1081),
    .D(_00034_),
    .Q_N(_13560_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[8]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1082),
    .D(_00035_),
    .Q_N(_13561_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[9]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1082),
    .D(_00036_),
    .Q_N(_11276_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1102),
    .D(_02816_),
    .Q_N(_11275_),
    .Q(\top_ihp.wb_dati_uart[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1102),
    .D(_02817_),
    .Q_N(_11274_),
    .Q(\top_ihp.wb_dati_uart[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1102),
    .D(_02818_),
    .Q_N(_11273_),
    .Q(\top_ihp.wb_dati_uart[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1102),
    .D(_02819_),
    .Q_N(_11272_),
    .Q(\top_ihp.wb_dati_uart[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1101),
    .D(_02820_),
    .Q_N(_11271_),
    .Q(\top_ihp.wb_dati_uart[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1102),
    .D(_02821_),
    .Q_N(_11270_),
    .Q(\top_ihp.wb_dati_uart[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1107),
    .D(_02822_),
    .Q_N(_11269_),
    .Q(\top_ihp.wb_dati_uart[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1107),
    .D(_02823_),
    .Q_N(_11268_),
    .Q(\top_ihp.wb_dati_uart[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data_ready$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1084),
    .D(_02824_),
    .Q_N(_13562_),
    .Q(\top_ihp.wb_uart.rx_ready ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.state[0]$_DFF_PN0_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1101),
    .D(\top_ihp.wb_uart.uart_rx.next_state[0] ),
    .Q_N(_13563_),
    .Q(\top_ihp.wb_uart.uart_rx.state[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.state[1]$_DFF_PN0_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1110),
    .D(\top_ihp.wb_uart.uart_rx.next_state[1] ),
    .Q_N(_13564_),
    .Q(\top_ihp.wb_uart.uart_rx.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.state[2]$_DFF_PN0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1110),
    .D(\top_ihp.wb_uart.uart_rx.next_state[2] ),
    .Q_N(_00093_),
    .Q(\top_ihp.wb_uart.uart_rx.state[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.bit_cnt[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1077),
    .D(_02825_),
    .Q_N(_11267_),
    .Q(\top_ihp.wb_uart.uart_tx.bit_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.bit_cnt[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1077),
    .D(_02826_),
    .Q_N(_11266_),
    .Q(\top_ihp.wb_uart.uart_tx.bit_cnt[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.bit_cnt[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1077),
    .D(_02827_),
    .Q_N(_00184_),
    .Q(\top_ihp.wb_uart.uart_tx.bit_cnt[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.bit_cnt[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1081),
    .D(_02828_),
    .Q_N(_13565_),
    .Q(\top_ihp.wb_uart.uart_tx.bit_cnt[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[0]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1073),
    .D(_00037_),
    .Q_N(_13566_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[10]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1076),
    .D(_00038_),
    .Q_N(_13567_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[11]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1076),
    .D(_00039_),
    .Q_N(_13568_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[12]$_DFF_PN0_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1076),
    .D(_00040_),
    .Q_N(_13569_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[13]$_DFF_PN0_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1076),
    .D(_00041_),
    .Q_N(_13570_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[14]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1076),
    .D(_00042_),
    .Q_N(_13571_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[15]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1079),
    .D(_00043_),
    .Q_N(_13572_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[16]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1076),
    .D(_00044_),
    .Q_N(_13573_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[17]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1076),
    .D(_00045_),
    .Q_N(_13574_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[18]$_DFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1077),
    .D(_00046_),
    .Q_N(_13575_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[19]$_DFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1074),
    .D(_00047_),
    .Q_N(_13576_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[1]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1073),
    .D(_00048_),
    .Q_N(_13577_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[20]$_DFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1074),
    .D(_00049_),
    .Q_N(_13578_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[21]$_DFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1074),
    .D(_00050_),
    .Q_N(_13579_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[22]$_DFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1074),
    .D(_00051_),
    .Q_N(_13580_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[23]$_DFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1074),
    .D(_00052_),
    .Q_N(_13581_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[24]$_DFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1074),
    .D(_00053_),
    .Q_N(_13582_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[25]$_DFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1074),
    .D(_00054_),
    .Q_N(_13583_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[26]$_DFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1074),
    .D(_00055_),
    .Q_N(_13584_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[27]$_DFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1080),
    .D(_00056_),
    .Q_N(_13585_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[28]$_DFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1080),
    .D(_00057_),
    .Q_N(_13586_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[29]$_DFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1080),
    .D(_00058_),
    .Q_N(_13587_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[2]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1073),
    .D(_00059_),
    .Q_N(_13588_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[30]$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1075),
    .D(_00060_),
    .Q_N(_13589_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[31]$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1075),
    .D(_00061_),
    .Q_N(_13590_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[3]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1073),
    .D(_00062_),
    .Q_N(_13591_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[4]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1073),
    .D(_00063_),
    .Q_N(_13592_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[5]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1073),
    .D(_00064_),
    .Q_N(_13593_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[6]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1073),
    .D(_00065_),
    .Q_N(_13594_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[7]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1073),
    .D(_00066_),
    .Q_N(_13595_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[8]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1075),
    .D(_00067_),
    .Q_N(_13596_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[9]$_DFF_PN0_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1076),
    .D(_00068_),
    .Q_N(_13597_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.state[0]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1083),
    .D(\top_ihp.wb_uart.uart_tx.next_state[0] ),
    .Q_N(_13598_),
    .Q(\top_ihp.wb_uart.uart_tx.state[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.state[1]$_DFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1083),
    .D(\top_ihp.wb_uart.uart_tx.next_state[1] ),
    .Q_N(_11265_),
    .Q(\top_ihp.wb_uart.uart_tx.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1077),
    .D(_02829_),
    .Q_N(_11264_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1077),
    .D(_02830_),
    .Q_N(_11263_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1078),
    .D(_02831_),
    .Q_N(_11262_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1078),
    .D(_02832_),
    .Q_N(_11261_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1077),
    .D(_02833_),
    .Q_N(_11260_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1083),
    .D(_02834_),
    .Q_N(_11259_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1083),
    .D(_02835_),
    .Q_N(_11258_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1084),
    .D(_02836_),
    .Q_N(_11257_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_ready$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1083),
    .D(_02837_),
    .Q_N(_11256_),
    .Q(\top_ihp.wb_uart.tx_ready ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_reg$_DFF_PN1_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1084),
    .D(_00324_),
    .Q_N(\top_ihp.tx ),
    .Q(_13602_));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[0]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[1]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[2]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[3]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[4]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[5]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[6]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[7]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[0]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[1]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[2]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[3]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[4]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[5]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[6]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout26 (.X(net26),
    .A(_05943_));
 sg13g2_buf_2 fanout27 (.A(_05746_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_03474_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_03096_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_03094_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_03091_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_03089_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_03063_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_03054_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_03049_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_03047_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_03034_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_03014_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_03004_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_11060_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_11058_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_11055_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_11053_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_11027_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_11018_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_11016_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_11011_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_11009_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_10996_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_10973_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_10960_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_10349_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_09698_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_08738_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_08711_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_08688_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_06017_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_06009_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_06008_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_05944_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_05918_),
    .X(net61));
 sg13g2_buf_4 fanout62 (.X(net62),
    .A(_05742_));
 sg13g2_buf_4 fanout63 (.X(net63),
    .A(_05708_));
 sg13g2_buf_2 fanout64 (.A(_04817_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_03539_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_03537_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_03534_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_03532_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_03505_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_03498_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_03496_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_03491_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_03489_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_03472_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_03466_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_03461_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_03458_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_03451_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_03446_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_03444_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_03441_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_03056_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_03052_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_03040_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_03036_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_03030_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_03025_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_03020_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_03018_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_03016_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_03010_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_02980_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_02971_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_02955_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_02926_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_02912_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_02892_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_02879_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_11222_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_11198_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_11174_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_11170_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_11161_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_11158_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_11126_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_11112_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_11014_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_11002_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_10998_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_10993_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_10992_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_10984_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_10980_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_10979_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_10977_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_10975_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_10969_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_10957_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_10845_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_10830_),
    .X(net120));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(_10648_));
 sg13g2_buf_2 fanout122 (.A(_10646_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_10645_),
    .X(net123));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(_10643_));
 sg13g2_buf_2 fanout125 (.A(_10638_),
    .X(net125));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(_10628_));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(_10624_));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(_10623_));
 sg13g2_buf_2 fanout129 (.A(_10609_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_10608_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_10604_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_10597_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_10548_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_10543_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_10536_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_10534_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_10531_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_10514_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_10484_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_10469_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_10440_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_10413_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_10381_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_10327_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_10315_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_10248_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_10237_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_10189_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_10128_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_10015_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_09993_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_09978_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_09906_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_09861_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_09825_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_09697_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_08607_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_08581_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_08555_),
    .X(net159));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(_06238_));
 sg13g2_buf_4 fanout161 (.X(net161),
    .A(_06189_));
 sg13g2_buf_2 fanout162 (.A(_06163_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_06156_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_06149_),
    .X(net164));
 sg13g2_buf_4 fanout165 (.X(net165),
    .A(_06115_));
 sg13g2_buf_2 fanout166 (.A(_06106_),
    .X(net166));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(_06102_));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(_06068_));
 sg13g2_buf_2 fanout169 (.A(_06066_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_06059_),
    .X(net170));
 sg13g2_buf_4 fanout171 (.X(net171),
    .A(_06029_));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(_05999_));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(_05994_));
 sg13g2_buf_2 fanout174 (.A(_05983_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_05965_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_05939_),
    .X(net176));
 sg13g2_buf_4 fanout177 (.X(net177),
    .A(_05924_));
 sg13g2_buf_2 fanout178 (.A(_05923_),
    .X(net178));
 sg13g2_buf_4 fanout179 (.X(net179),
    .A(_05901_));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(_05899_));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(_05896_));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(_05895_));
 sg13g2_buf_4 fanout183 (.X(net183),
    .A(_05893_));
 sg13g2_buf_2 fanout184 (.A(_05889_),
    .X(net184));
 sg13g2_buf_4 fanout185 (.X(net185),
    .A(_05884_));
 sg13g2_buf_2 fanout186 (.A(_05875_),
    .X(net186));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(_05867_));
 sg13g2_buf_2 fanout188 (.A(_05863_),
    .X(net188));
 sg13g2_buf_4 fanout189 (.X(net189),
    .A(_05848_));
 sg13g2_buf_2 fanout190 (.A(_05836_),
    .X(net190));
 sg13g2_buf_4 fanout191 (.X(net191),
    .A(_05833_));
 sg13g2_buf_2 fanout192 (.A(_05812_),
    .X(net192));
 sg13g2_buf_4 fanout193 (.X(net193),
    .A(_05805_));
 sg13g2_buf_4 fanout194 (.X(net194),
    .A(_05799_));
 sg13g2_buf_4 fanout195 (.X(net195),
    .A(_05791_));
 sg13g2_buf_2 fanout196 (.A(_05787_),
    .X(net196));
 sg13g2_buf_4 fanout197 (.X(net197),
    .A(_05715_));
 sg13g2_buf_2 fanout198 (.A(_05684_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_05677_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_05674_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_05652_),
    .X(net201));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(_05629_));
 sg13g2_buf_2 fanout203 (.A(_05531_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_05501_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_05242_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_04946_),
    .X(net206));
 sg13g2_buf_4 fanout207 (.X(net207),
    .A(_04867_));
 sg13g2_buf_4 fanout208 (.X(net208),
    .A(_04844_));
 sg13g2_buf_2 fanout209 (.A(_04823_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_04821_),
    .X(net210));
 sg13g2_buf_4 fanout211 (.X(net211),
    .A(_04394_));
 sg13g2_buf_4 fanout212 (.X(net212),
    .A(_04393_));
 sg13g2_buf_4 fanout213 (.X(net213),
    .A(_04392_));
 sg13g2_buf_4 fanout214 (.X(net214),
    .A(_04389_));
 sg13g2_buf_4 fanout215 (.X(net215),
    .A(_04388_));
 sg13g2_buf_4 fanout216 (.X(net216),
    .A(_04387_));
 sg13g2_buf_4 fanout217 (.X(net217),
    .A(_04327_));
 sg13g2_buf_4 fanout218 (.X(net218),
    .A(_04272_));
 sg13g2_buf_4 fanout219 (.X(net219),
    .A(_04217_));
 sg13g2_buf_2 fanout220 (.A(_03510_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_03494_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_03482_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_03479_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_03477_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_03470_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_03468_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_03464_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_03456_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_03453_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_03448_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_03128_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_03123_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_03108_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_03105_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_03084_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_03080_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_03068_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_03066_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_03060_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_03059_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_03038_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_03031_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_03028_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_03023_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_03008_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_03002_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_02999_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_02963_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_02956_),
    .X(net249));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(_02954_));
 sg13g2_buf_2 fanout251 (.A(_02943_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_02939_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_02929_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_02915_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_02911_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_02894_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_02887_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_02875_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_02869_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_02868_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_02848_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_02843_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_11249_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_11244_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_11241_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_11213_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_11205_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_11199_),
    .X(net268));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(_11197_));
 sg13g2_buf_2 fanout270 (.A(_11139_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_11129_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_11115_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_11111_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_11091_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_11090_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_11077_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_11072_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_11069_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_11046_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_11041_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_11031_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_11024_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_11021_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_11000_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_10987_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_10967_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_10958_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_10956_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_10939_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_10936_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_10927_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_10924_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_10915_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_10914_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_10901_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_10900_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_10889_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_10888_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_10874_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_10873_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_10858_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_10848_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_10834_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_10829_),
    .X(net304));
 sg13g2_buf_4 fanout305 (.X(net305),
    .A(_10647_));
 sg13g2_buf_2 fanout306 (.A(_10644_),
    .X(net306));
 sg13g2_buf_4 fanout307 (.X(net307),
    .A(_10642_));
 sg13g2_buf_2 fanout308 (.A(_10639_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_10636_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_10633_),
    .X(net310));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(_10631_));
 sg13g2_buf_2 fanout312 (.A(_10630_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_10629_),
    .X(net313));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(_10626_));
 sg13g2_buf_2 fanout315 (.A(_10606_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_10499_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_10281_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_10260_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_10236_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_10217_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_10204_),
    .X(net321));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(_10188_));
 sg13g2_buf_2 fanout323 (.A(_10169_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_10153_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_10127_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_10085_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_10060_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_10039_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_09992_),
    .X(net329));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(_09977_));
 sg13g2_buf_2 fanout331 (.A(_09942_),
    .X(net331));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(_09905_));
 sg13g2_buf_2 fanout333 (.A(_06310_),
    .X(net333));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(_06276_));
 sg13g2_buf_2 fanout335 (.A(_06271_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_06172_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_06143_),
    .X(net337));
 sg13g2_buf_4 fanout338 (.X(net338),
    .A(_06141_));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(_06139_));
 sg13g2_buf_4 fanout340 (.X(net340),
    .A(_06086_));
 sg13g2_buf_2 fanout341 (.A(_06080_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_06065_),
    .X(net342));
 sg13g2_buf_4 fanout343 (.X(net343),
    .A(_06063_));
 sg13g2_buf_2 fanout344 (.A(_06052_),
    .X(net344));
 sg13g2_buf_4 fanout345 (.X(net345),
    .A(_06046_));
 sg13g2_buf_4 fanout346 (.X(net346),
    .A(_06042_));
 sg13g2_buf_2 fanout347 (.A(_06040_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_06020_),
    .X(net348));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(_06018_));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(_06002_));
 sg13g2_buf_2 fanout351 (.A(_05986_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_05981_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_05978_),
    .X(net353));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(_05966_));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(_05961_));
 sg13g2_buf_2 fanout356 (.A(_05960_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_05954_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_05951_),
    .X(net358));
 sg13g2_buf_4 fanout359 (.X(net359),
    .A(_05949_));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(_05937_));
 sg13g2_buf_4 fanout361 (.X(net361),
    .A(_05935_));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(_05934_));
 sg13g2_buf_4 fanout363 (.X(net363),
    .A(_05932_));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(_05929_));
 sg13g2_buf_2 fanout365 (.A(_05927_),
    .X(net365));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(_05919_));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(_05911_));
 sg13g2_buf_2 fanout368 (.A(_05903_),
    .X(net368));
 sg13g2_buf_4 fanout369 (.X(net369),
    .A(_05900_));
 sg13g2_buf_2 fanout370 (.A(_05898_),
    .X(net370));
 sg13g2_buf_4 fanout371 (.X(net371),
    .A(_05892_));
 sg13g2_buf_4 fanout372 (.X(net372),
    .A(_05888_));
 sg13g2_buf_2 fanout373 (.A(_05887_),
    .X(net373));
 sg13g2_buf_4 fanout374 (.X(net374),
    .A(_05883_));
 sg13g2_buf_2 fanout375 (.A(_05872_),
    .X(net375));
 sg13g2_buf_4 fanout376 (.X(net376),
    .A(_05870_));
 sg13g2_buf_2 fanout377 (.A(_05869_),
    .X(net377));
 sg13g2_buf_4 fanout378 (.X(net378),
    .A(_05864_));
 sg13g2_buf_4 fanout379 (.X(net379),
    .A(_05861_));
 sg13g2_buf_4 fanout380 (.X(net380),
    .A(_05857_));
 sg13g2_buf_4 fanout381 (.X(net381),
    .A(_05855_));
 sg13g2_buf_4 fanout382 (.X(net382),
    .A(_05854_));
 sg13g2_buf_4 fanout383 (.X(net383),
    .A(_05847_));
 sg13g2_buf_4 fanout384 (.X(net384),
    .A(_05844_));
 sg13g2_buf_2 fanout385 (.A(_05843_),
    .X(net385));
 sg13g2_buf_4 fanout386 (.X(net386),
    .A(_05841_));
 sg13g2_buf_4 fanout387 (.X(net387),
    .A(_05839_));
 sg13g2_buf_2 fanout388 (.A(_05835_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_05830_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_05828_),
    .X(net390));
 sg13g2_buf_4 fanout391 (.X(net391),
    .A(_05814_));
 sg13g2_buf_4 fanout392 (.X(net392),
    .A(_05810_));
 sg13g2_buf_2 fanout393 (.A(_05809_),
    .X(net393));
 sg13g2_buf_4 fanout394 (.X(net394),
    .A(_05802_));
 sg13g2_buf_4 fanout395 (.X(net395),
    .A(_05800_));
 sg13g2_buf_4 fanout396 (.X(net396),
    .A(_05796_));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(_05795_));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(_05793_));
 sg13g2_buf_4 fanout399 (.X(net399),
    .A(_05790_));
 sg13g2_buf_2 fanout400 (.A(_05783_),
    .X(net400));
 sg13g2_buf_4 fanout401 (.X(net401),
    .A(_05778_));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(_05776_));
 sg13g2_buf_2 fanout403 (.A(_05736_),
    .X(net403));
 sg13g2_buf_4 fanout404 (.X(net404),
    .A(_05733_));
 sg13g2_buf_4 fanout405 (.X(net405),
    .A(_05729_));
 sg13g2_buf_4 fanout406 (.X(net406),
    .A(_05726_));
 sg13g2_buf_4 fanout407 (.X(net407),
    .A(_05722_));
 sg13g2_buf_2 fanout408 (.A(_05719_),
    .X(net408));
 sg13g2_buf_4 fanout409 (.X(net409),
    .A(_05714_));
 sg13g2_buf_4 fanout410 (.X(net410),
    .A(_05711_));
 sg13g2_buf_2 fanout411 (.A(_05681_),
    .X(net411));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(_05670_));
 sg13g2_buf_2 fanout413 (.A(_05665_),
    .X(net413));
 sg13g2_buf_4 fanout414 (.X(net414),
    .A(_05660_));
 sg13g2_buf_2 fanout415 (.A(_05648_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_05645_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_05641_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_05636_),
    .X(net418));
 sg13g2_buf_4 fanout419 (.X(net419),
    .A(_05628_));
 sg13g2_buf_2 fanout420 (.A(_05626_),
    .X(net420));
 sg13g2_buf_4 fanout421 (.X(net421),
    .A(_05618_));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(_05615_));
 sg13g2_buf_4 fanout423 (.X(net423),
    .A(_05609_));
 sg13g2_buf_4 fanout424 (.X(net424),
    .A(_05606_));
 sg13g2_buf_4 fanout425 (.X(net425),
    .A(_05602_));
 sg13g2_buf_4 fanout426 (.X(net426),
    .A(_05596_));
 sg13g2_buf_4 fanout427 (.X(net427),
    .A(_05574_));
 sg13g2_buf_2 fanout428 (.A(_05571_),
    .X(net428));
 sg13g2_buf_4 fanout429 (.X(net429),
    .A(_05530_));
 sg13g2_buf_2 fanout430 (.A(_05515_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_05507_),
    .X(net431));
 sg13g2_buf_4 fanout432 (.X(net432),
    .A(_05500_));
 sg13g2_buf_4 fanout433 (.X(net433),
    .A(_05483_));
 sg13g2_buf_2 fanout434 (.A(_05473_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_05461_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_05456_),
    .X(net436));
 sg13g2_buf_4 fanout437 (.X(net437),
    .A(_05440_));
 sg13g2_buf_2 fanout438 (.A(_05430_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_05047_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_05035_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_04992_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_04983_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_04945_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_04937_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_04018_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_04015_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_04006_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_04003_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_03993_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_03938_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_03935_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_03926_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_03923_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_03913_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_03858_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_03855_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_03846_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_03843_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_03833_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_03776_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_03773_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_03764_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_03761_),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_03751_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_03574_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_03571_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_03562_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_03559_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_03549_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_03543_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_03480_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_03475_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(_03459_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(_03454_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_03438_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_03381_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_03378_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_03369_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_03366_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_03356_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_03299_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_03296_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_03287_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_03284_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_03274_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_03258_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_03255_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_03246_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_03243_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_03233_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_03176_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_03173_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_03164_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_03161_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_03151_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_03107_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_03058_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_03001_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_02874_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_02867_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_02862_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_11068_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_11023_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_10809_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_10806_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_10797_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_10794_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_10784_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_10690_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_10687_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_10678_),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_10675_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_10665_),
    .X(net513));
 sg13g2_buf_4 fanout514 (.X(net514),
    .A(_10641_));
 sg13g2_buf_4 fanout515 (.X(net515),
    .A(_10640_));
 sg13g2_buf_4 fanout516 (.X(net516),
    .A(_10627_));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(_10622_));
 sg13g2_buf_2 fanout518 (.A(_10612_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_10557_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_10554_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_10544_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_10540_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_10528_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_10527_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_10269_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_10262_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_10249_),
    .X(net527));
 sg13g2_buf_4 fanout528 (.X(net528),
    .A(_10203_));
 sg13g2_buf_2 fanout529 (.A(_10062_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_10040_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_09757_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_08685_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_06146_),
    .X(net533));
 sg13g2_buf_4 fanout534 (.X(net534),
    .A(_06062_));
 sg13g2_buf_4 fanout535 (.X(net535),
    .A(_06001_));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(_05914_));
 sg13g2_buf_2 fanout537 (.A(_05905_),
    .X(net537));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(_05885_));
 sg13g2_buf_4 fanout539 (.X(net539),
    .A(_05873_));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(_05782_));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(_05770_));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(_05617_));
 sg13g2_buf_2 fanout543 (.A(_05551_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_05548_),
    .X(net544));
 sg13g2_buf_4 fanout545 (.X(net545),
    .A(_05520_));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(_05514_));
 sg13g2_buf_2 fanout547 (.A(_05506_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_05492_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_05489_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_05486_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_05482_),
    .X(net551));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(_05472_));
 sg13g2_buf_2 fanout553 (.A(_05439_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_05429_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_05208_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_04322_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_04320_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_04319_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_04267_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_04265_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_04264_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_04210_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_04205_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_04195_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_03994_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_03992_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_03978_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_03975_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_03966_),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(_03963_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_03953_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_03914_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_03912_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_03898_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_03895_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_03886_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_03883_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_03873_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_03834_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_03832_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_03817_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_03814_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_03805_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_03802_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_03792_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_03752_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_03750_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_03696_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_03693_),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_03684_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_03681_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_03671_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_03656_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_03653_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_03644_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_03641_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_03631_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(_03615_),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_03612_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_03603_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_03600_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_03590_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_03550_),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_03548_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_03529_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_03526_),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_03519_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_03516_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_03513_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_03501_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_03439_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_03437_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_03422_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_03419_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_03410_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_03407_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_03397_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_03357_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_03355_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_03341_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_03338_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_03329_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_03326_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_03316_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_03275_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_03273_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_03234_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_03232_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_03218_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_03215_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_03206_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_03203_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_03193_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_03152_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_03150_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_02842_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_11182_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_11179_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_11168_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_11165_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_11153_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_10785_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_10783_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_10730_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_10727_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_10718_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_10715_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_10705_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_10666_),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_10664_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_10621_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_10600_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_10591_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_10589_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_10586_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_10577_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_10576_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_10575_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_10526_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_09758_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_09756_),
    .X(net661));
 sg13g2_buf_4 fanout662 (.X(net662),
    .A(_06094_));
 sg13g2_buf_2 fanout663 (.A(_06091_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_06057_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_05913_),
    .X(net665));
 sg13g2_buf_4 fanout666 (.X(net666),
    .A(_05821_));
 sg13g2_buf_2 fanout667 (.A(_05784_),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(_05543_),
    .X(net668));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(_05519_));
 sg13g2_buf_4 fanout670 (.X(net670),
    .A(_05491_));
 sg13g2_buf_2 fanout671 (.A(_05488_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_05485_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_05413_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_04058_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_04055_),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(_04046_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_04043_),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_04033_),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(_03954_),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_03952_),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(_03874_),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(_03872_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_03793_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(_03791_),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(_03736_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(_03733_),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_03724_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_03721_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_03711_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(_03672_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_03670_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(_03632_),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_03630_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_03591_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(_03589_),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_03502_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_03500_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(_03398_),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(_03396_),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(_03317_),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_03315_),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(_03194_),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(_03192_),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(_11154_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_11152_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_10881_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(_10831_),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(_10826_),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(_10770_),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(_10767_),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(_10758_),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(_10755_),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(_10746_),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(_10745_),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(_10706_),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(_10704_),
    .X(net716));
 sg13g2_buf_4 fanout717 (.X(net717),
    .A(_10657_));
 sg13g2_buf_2 fanout718 (.A(_10654_),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(_05970_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(_05825_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_05598_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_05586_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_05535_),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(_05523_),
    .X(net724));
 sg13g2_buf_4 fanout725 (.X(net725),
    .A(_05518_));
 sg13g2_buf_2 fanout726 (.A(_05479_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(_05469_),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(_05452_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(_05388_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_04034_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_04032_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_03712_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_03710_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(_10744_),
    .X(net734));
 sg13g2_buf_4 fanout735 (.X(net735),
    .A(_10662_));
 sg13g2_buf_2 fanout736 (.A(_10653_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_05198_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_04323_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_04268_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_04211_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_10870_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_10430_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_07537_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_07518_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_07435_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_06304_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_06175_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_05537_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_05495_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_05487_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_05416_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_05398_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_05394_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_05380_),
    .X(net754));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(_05345_));
 sg13g2_buf_2 fanout756 (.A(_05333_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(_05256_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_05232_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_04967_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_04088_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_03113_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_10988_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_10619_),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_10520_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_10392_),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_09752_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_09726_),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_08808_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_08807_),
    .X(net769));
 sg13g2_buf_4 fanout770 (.X(net770),
    .A(_07565_));
 sg13g2_buf_2 fanout771 (.A(_07531_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_07505_),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(_07475_),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_05512_),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(_05212_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(_05188_),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(_04996_),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(_04993_),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(_04962_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(_04576_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_04569_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_04093_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_04087_),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(_10822_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(_10570_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_09949_),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(_09917_),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(_09875_),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(_08806_),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(_08214_),
    .X(net790));
 sg13g2_buf_4 fanout791 (.X(net791),
    .A(_07634_));
 sg13g2_buf_2 fanout792 (.A(_07559_),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(_07541_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(_07540_),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_07534_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(_07515_),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_07504_));
 sg13g2_buf_2 fanout798 (.A(_07474_),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(_07455_),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(_07444_),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(_06023_),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(_04948_),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(_04086_),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(_04075_),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(_09925_),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(_08827_),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(_08805_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_08224_),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(_08213_),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(_07721_),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(_07677_),
    .X(net811));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(_07599_));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(_07595_));
 sg13g2_buf_2 fanout814 (.A(_07577_),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(_07570_),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(_07556_),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(_07550_),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(_07548_),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(_07547_),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(_07542_),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_07532_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(_07525_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(_07512_),
    .X(net823));
 sg13g2_buf_4 fanout824 (.X(net824),
    .A(_07508_));
 sg13g2_buf_2 fanout825 (.A(_07493_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_07481_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_07478_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_07471_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_07465_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_07462_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_07454_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_04568_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_04495_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_04459_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(_04085_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_08640_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_07978_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_07644_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_07602_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_07563_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_07549_),
    .X(net841));
 sg13g2_buf_4 fanout842 (.X(net842),
    .A(_07520_));
 sg13g2_buf_2 fanout843 (.A(_07492_),
    .X(net843));
 sg13g2_buf_4 fanout844 (.X(net844),
    .A(_07488_));
 sg13g2_buf_2 fanout845 (.A(_07461_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_07449_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_04621_),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_04516_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_04508_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_04504_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_04473_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_04469_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_04443_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_09615_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_09609_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_08825_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_07977_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_07682_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_07628_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_07555_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_07539_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_07485_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_07448_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_07438_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_04542_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_04534_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_04531_),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(_04510_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_04491_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(_04488_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_04468_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_04455_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_04452_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(_04450_),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(_04446_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_04442_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_09632_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_09614_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_09608_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_09493_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_08965_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_08832_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_08207_),
    .X(net883));
 sg13g2_buf_4 fanout884 (.X(net884),
    .A(_07603_));
 sg13g2_buf_2 fanout885 (.A(_07498_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_04868_),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(_04845_),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(_09612_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(_09607_),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_09519_),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_08784_),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(_07708_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(_07497_),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_04862_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_04848_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(_04815_),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_04400_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_09864_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(_09622_),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(_09605_),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_09070_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(_08904_),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(_08900_),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(_08770_),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(_08372_),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(_04146_),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(_04133_),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(_04131_),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(_04122_),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(_04111_),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(_04109_),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_10009_),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(_09870_),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(_09869_),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_09865_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_09863_),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(_09748_),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(_09655_),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(_09621_),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_09604_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_09600_),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(_09487_),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(_09169_),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(_09099_),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(_09040_),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(_09026_),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(_08975_),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(_08947_),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(_08939_),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(_08938_),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(_08913_),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(_08903_),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(_08899_),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(_08888_),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(_08880_),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_08875_),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(_08860_),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(_08846_),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_07987_),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(_05415_),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(_05353_),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(_04583_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_04566_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(_09909_),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_09908_),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(_09856_),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(_09848_),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_09819_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_09693_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(_09620_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(_09618_),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(_09599_),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_09593_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_09082_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(_09025_),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_08969_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_08956_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_08954_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_08946_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_08940_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_08937_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_08923_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_08915_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_08912_),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(_08902_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(_08898_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_08854_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_08845_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_08838_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(_08777_),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_08310_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(_08195_),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_07986_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_07982_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(_05364_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_05030_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_04985_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_04971_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_04966_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_04959_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_04565_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_04402_),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(_04396_),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(_04079_),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(_09849_),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(_09798_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_09788_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(_09707_),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(_09676_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_09657_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(_09653_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_09631_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_09627_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_09617_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_09596_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_09592_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_09180_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_09015_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_08998_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_08968_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_08953_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_08936_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_08935_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_08908_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_08895_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_08891_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(_08889_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_08885_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(_08873_),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(_08865_),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(_08858_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(_08853_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_08849_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_08841_),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_08837_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(_08812_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_08221_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_08194_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_07985_),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_05374_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(_04078_),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(_09820_),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(_09815_),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_09784_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_09689_),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(_09678_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(_09675_),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_09661_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_09616_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_09602_),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_09495_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(_08952_),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(_08881_),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_08877_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_08872_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_08867_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(_08861_),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(_08843_),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(_08840_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_08834_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_08772_),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(_08475_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(_08307_),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(_08290_),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(_08122_),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(_08050_),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_07984_),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(_07980_),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(_07960_),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(_04110_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(_09594_),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(_09590_),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(_08856_),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(_08855_),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_08489_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(_08479_),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_08276_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(_08208_),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_08197_),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_08169_),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(_08163_),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(_08123_),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(_08036_),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(_08033_),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(_08029_),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(_08019_),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(_08014_),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(_08012_),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(_08010_),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(_07995_),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(_07994_),
    .X(net1071));
 sg13g2_buf_2 fanout1072 (.A(_08493_),
    .X(net1072));
 sg13g2_buf_4 fanout1073 (.X(net1073),
    .A(net1075));
 sg13g2_buf_4 fanout1074 (.X(net1074),
    .A(net1075));
 sg13g2_buf_2 fanout1075 (.A(net1098),
    .X(net1075));
 sg13g2_buf_4 fanout1076 (.X(net1076),
    .A(net1079));
 sg13g2_buf_4 fanout1077 (.X(net1077),
    .A(net1079));
 sg13g2_buf_2 fanout1078 (.A(net1079),
    .X(net1078));
 sg13g2_buf_1 fanout1079 (.A(net1098),
    .X(net1079));
 sg13g2_buf_4 fanout1080 (.X(net1080),
    .A(net1081));
 sg13g2_buf_2 fanout1081 (.A(net1085),
    .X(net1081));
 sg13g2_buf_4 fanout1082 (.X(net1082),
    .A(net1085));
 sg13g2_buf_4 fanout1083 (.X(net1083),
    .A(net1084));
 sg13g2_buf_4 fanout1084 (.X(net1084),
    .A(net1085));
 sg13g2_buf_1 fanout1085 (.A(net1098),
    .X(net1085));
 sg13g2_buf_4 fanout1086 (.X(net1086),
    .A(net1089));
 sg13g2_buf_2 fanout1087 (.A(net1089),
    .X(net1087));
 sg13g2_buf_4 fanout1088 (.X(net1088),
    .A(net1089));
 sg13g2_buf_2 fanout1089 (.A(net1097),
    .X(net1089));
 sg13g2_buf_4 fanout1090 (.X(net1090),
    .A(net1097));
 sg13g2_buf_4 fanout1091 (.X(net1091),
    .A(net1097));
 sg13g2_buf_4 fanout1092 (.X(net1092),
    .A(net1096));
 sg13g2_buf_2 fanout1093 (.A(net1096),
    .X(net1093));
 sg13g2_buf_4 fanout1094 (.X(net1094),
    .A(net1096));
 sg13g2_buf_4 fanout1095 (.X(net1095),
    .A(net1096));
 sg13g2_buf_1 fanout1096 (.A(net1097),
    .X(net1096));
 sg13g2_buf_1 fanout1097 (.A(net1098),
    .X(net1097));
 sg13g2_buf_1 fanout1098 (.A(net1207),
    .X(net1098));
 sg13g2_buf_4 fanout1099 (.X(net1099),
    .A(net1100));
 sg13g2_buf_4 fanout1100 (.X(net1100),
    .A(net1101));
 sg13g2_buf_4 fanout1101 (.X(net1101),
    .A(net1110));
 sg13g2_buf_4 fanout1102 (.X(net1102),
    .A(net1103));
 sg13g2_buf_4 fanout1103 (.X(net1103),
    .A(net1107));
 sg13g2_buf_4 fanout1104 (.X(net1104),
    .A(net1106));
 sg13g2_buf_4 fanout1105 (.X(net1105),
    .A(net1106));
 sg13g2_buf_4 fanout1106 (.X(net1106),
    .A(net1107));
 sg13g2_buf_2 fanout1107 (.A(net1110),
    .X(net1107));
 sg13g2_buf_4 fanout1108 (.X(net1108),
    .A(net1109));
 sg13g2_buf_4 fanout1109 (.X(net1109),
    .A(net1110));
 sg13g2_buf_2 fanout1110 (.A(net1207),
    .X(net1110));
 sg13g2_buf_4 fanout1111 (.X(net1111),
    .A(net1112));
 sg13g2_buf_2 fanout1112 (.A(net1113),
    .X(net1112));
 sg13g2_buf_4 fanout1113 (.X(net1113),
    .A(net1117));
 sg13g2_buf_4 fanout1114 (.X(net1114),
    .A(net1116));
 sg13g2_buf_2 fanout1115 (.A(net1116),
    .X(net1115));
 sg13g2_buf_4 fanout1116 (.X(net1116),
    .A(net1117));
 sg13g2_buf_2 fanout1117 (.A(net1149),
    .X(net1117));
 sg13g2_buf_4 fanout1118 (.X(net1118),
    .A(net1122));
 sg13g2_buf_2 fanout1119 (.A(net1122),
    .X(net1119));
 sg13g2_buf_4 fanout1120 (.X(net1120),
    .A(net1121));
 sg13g2_buf_4 fanout1121 (.X(net1121),
    .A(net1122));
 sg13g2_buf_1 fanout1122 (.A(net1149),
    .X(net1122));
 sg13g2_buf_4 fanout1123 (.X(net1123),
    .A(net1125));
 sg13g2_buf_4 fanout1124 (.X(net1124),
    .A(net1125));
 sg13g2_buf_2 fanout1125 (.A(net1129),
    .X(net1125));
 sg13g2_buf_4 fanout1126 (.X(net1126),
    .A(net1128));
 sg13g2_buf_2 fanout1127 (.A(net1128),
    .X(net1127));
 sg13g2_buf_4 fanout1128 (.X(net1128),
    .A(net1129));
 sg13g2_buf_1 fanout1129 (.A(net1133),
    .X(net1129));
 sg13g2_buf_4 fanout1130 (.X(net1130),
    .A(net1131));
 sg13g2_buf_4 fanout1131 (.X(net1131),
    .A(net1132));
 sg13g2_buf_4 fanout1132 (.X(net1132),
    .A(net1133));
 sg13g2_buf_2 fanout1133 (.A(net1149),
    .X(net1133));
 sg13g2_buf_4 fanout1134 (.X(net1134),
    .A(net1138));
 sg13g2_buf_2 fanout1135 (.A(net1138),
    .X(net1135));
 sg13g2_buf_4 fanout1136 (.X(net1136),
    .A(net1138));
 sg13g2_buf_2 fanout1137 (.A(net1138),
    .X(net1137));
 sg13g2_buf_1 fanout1138 (.A(net1149),
    .X(net1138));
 sg13g2_buf_4 fanout1139 (.X(net1139),
    .A(net1140));
 sg13g2_buf_4 fanout1140 (.X(net1140),
    .A(net1142));
 sg13g2_buf_4 fanout1141 (.X(net1141),
    .A(net1142));
 sg13g2_buf_2 fanout1142 (.A(net1149),
    .X(net1142));
 sg13g2_buf_4 fanout1143 (.X(net1143),
    .A(net1148));
 sg13g2_buf_4 fanout1144 (.X(net1144),
    .A(net1145));
 sg13g2_buf_4 fanout1145 (.X(net1145),
    .A(net1148));
 sg13g2_buf_4 fanout1146 (.X(net1146),
    .A(net1147));
 sg13g2_buf_2 fanout1147 (.A(net1148),
    .X(net1147));
 sg13g2_buf_2 fanout1148 (.A(net1149),
    .X(net1148));
 sg13g2_buf_2 fanout1149 (.A(net1207),
    .X(net1149));
 sg13g2_buf_4 fanout1150 (.X(net1150),
    .A(net1151));
 sg13g2_buf_2 fanout1151 (.A(net1156),
    .X(net1151));
 sg13g2_buf_4 fanout1152 (.X(net1152),
    .A(net1156));
 sg13g2_buf_4 fanout1153 (.X(net1153),
    .A(net1156));
 sg13g2_buf_4 fanout1154 (.X(net1154),
    .A(net1155));
 sg13g2_buf_4 fanout1155 (.X(net1155),
    .A(net1156));
 sg13g2_buf_2 fanout1156 (.A(net1207),
    .X(net1156));
 sg13g2_buf_4 fanout1157 (.X(net1157),
    .A(net1158));
 sg13g2_buf_4 fanout1158 (.X(net1158),
    .A(net1164));
 sg13g2_buf_4 fanout1159 (.X(net1159),
    .A(net1164));
 sg13g2_buf_4 fanout1160 (.X(net1160),
    .A(net1161));
 sg13g2_buf_4 fanout1161 (.X(net1161),
    .A(net1162));
 sg13g2_buf_4 fanout1162 (.X(net1162),
    .A(net1163));
 sg13g2_buf_2 fanout1163 (.A(net1164),
    .X(net1163));
 sg13g2_buf_2 fanout1164 (.A(net1207),
    .X(net1164));
 sg13g2_buf_4 fanout1165 (.X(net1165),
    .A(net1169));
 sg13g2_buf_4 fanout1166 (.X(net1166),
    .A(net1169));
 sg13g2_buf_4 fanout1167 (.X(net1167),
    .A(net1168));
 sg13g2_buf_4 fanout1168 (.X(net1168),
    .A(net1169));
 sg13g2_buf_2 fanout1169 (.A(net1185),
    .X(net1169));
 sg13g2_buf_4 fanout1170 (.X(net1170),
    .A(net1174));
 sg13g2_buf_2 fanout1171 (.A(net1174),
    .X(net1171));
 sg13g2_buf_4 fanout1172 (.X(net1172),
    .A(net1174));
 sg13g2_buf_4 fanout1173 (.X(net1173),
    .A(net1174));
 sg13g2_buf_1 fanout1174 (.A(net1185),
    .X(net1174));
 sg13g2_buf_4 fanout1175 (.X(net1175),
    .A(net1178));
 sg13g2_buf_4 fanout1176 (.X(net1176),
    .A(net1178));
 sg13g2_buf_4 fanout1177 (.X(net1177),
    .A(net1178));
 sg13g2_buf_2 fanout1178 (.A(net1185),
    .X(net1178));
 sg13g2_buf_4 fanout1179 (.X(net1179),
    .A(net1180));
 sg13g2_buf_4 fanout1180 (.X(net1180),
    .A(net1184));
 sg13g2_buf_2 fanout1181 (.A(net1184),
    .X(net1181));
 sg13g2_buf_4 fanout1182 (.X(net1182),
    .A(net1184));
 sg13g2_buf_2 fanout1183 (.A(net1184),
    .X(net1183));
 sg13g2_buf_1 fanout1184 (.A(net1185),
    .X(net1184));
 sg13g2_buf_1 fanout1185 (.A(net1206),
    .X(net1185));
 sg13g2_buf_4 fanout1186 (.X(net1186),
    .A(net1190));
 sg13g2_buf_2 fanout1187 (.A(net1190),
    .X(net1187));
 sg13g2_buf_4 fanout1188 (.X(net1188),
    .A(net1190));
 sg13g2_buf_2 fanout1189 (.A(net1190),
    .X(net1189));
 sg13g2_buf_1 fanout1190 (.A(net1206),
    .X(net1190));
 sg13g2_buf_4 fanout1191 (.X(net1191),
    .A(net1192));
 sg13g2_buf_4 fanout1192 (.X(net1192),
    .A(net1195));
 sg13g2_buf_4 fanout1193 (.X(net1193),
    .A(net1195));
 sg13g2_buf_4 fanout1194 (.X(net1194),
    .A(net1195));
 sg13g2_buf_2 fanout1195 (.A(net1206),
    .X(net1195));
 sg13g2_buf_4 fanout1196 (.X(net1196),
    .A(net1197));
 sg13g2_buf_4 fanout1197 (.X(net1197),
    .A(net1205));
 sg13g2_buf_4 fanout1198 (.X(net1198),
    .A(net1199));
 sg13g2_buf_2 fanout1199 (.A(net1205),
    .X(net1199));
 sg13g2_buf_4 fanout1200 (.X(net1200),
    .A(net1202));
 sg13g2_buf_4 fanout1201 (.X(net1201),
    .A(net1202));
 sg13g2_buf_2 fanout1202 (.A(net1205),
    .X(net1202));
 sg13g2_buf_4 fanout1203 (.X(net1203),
    .A(net1205));
 sg13g2_buf_4 fanout1204 (.X(net1204),
    .A(net1205));
 sg13g2_buf_1 fanout1205 (.A(net1206),
    .X(net1205));
 sg13g2_buf_1 fanout1206 (.A(net1207),
    .X(net1206));
 sg13g2_buf_2 fanout1207 (.A(net1),
    .X(net1207));
 sg13g2_buf_4 fanout1208 (.X(net1208),
    .A(net1210));
 sg13g2_buf_4 fanout1209 (.X(net1209),
    .A(net1210));
 sg13g2_buf_2 fanout1210 (.A(net1218),
    .X(net1210));
 sg13g2_buf_4 fanout1211 (.X(net1211),
    .A(net1212));
 sg13g2_buf_4 fanout1212 (.X(net1212),
    .A(net1218));
 sg13g2_buf_4 fanout1213 (.X(net1213),
    .A(net1214));
 sg13g2_buf_4 fanout1214 (.X(net1214),
    .A(net1217));
 sg13g2_buf_4 fanout1215 (.X(net1215),
    .A(net1216));
 sg13g2_buf_2 fanout1216 (.A(net1217),
    .X(net1216));
 sg13g2_buf_2 fanout1217 (.A(net1218),
    .X(net1217));
 sg13g2_buf_1 fanout1218 (.A(net1247),
    .X(net1218));
 sg13g2_buf_4 fanout1219 (.X(net1219),
    .A(net1228));
 sg13g2_buf_2 fanout1220 (.A(net1228),
    .X(net1220));
 sg13g2_buf_4 fanout1221 (.X(net1221),
    .A(net1222));
 sg13g2_buf_4 fanout1222 (.X(net1222),
    .A(net1228));
 sg13g2_buf_4 fanout1223 (.X(net1223),
    .A(net1227));
 sg13g2_buf_2 fanout1224 (.A(net1227),
    .X(net1224));
 sg13g2_buf_4 fanout1225 (.X(net1225),
    .A(net1226));
 sg13g2_buf_4 fanout1226 (.X(net1226),
    .A(net1227));
 sg13g2_buf_2 fanout1227 (.A(net1228),
    .X(net1227));
 sg13g2_buf_1 fanout1228 (.A(net1247),
    .X(net1228));
 sg13g2_buf_4 fanout1229 (.X(net1229),
    .A(net1231));
 sg13g2_buf_4 fanout1230 (.X(net1230),
    .A(net1231));
 sg13g2_buf_2 fanout1231 (.A(net1233),
    .X(net1231));
 sg13g2_buf_4 fanout1232 (.X(net1232),
    .A(net1233));
 sg13g2_buf_2 fanout1233 (.A(net1238),
    .X(net1233));
 sg13g2_buf_4 fanout1234 (.X(net1234),
    .A(net1238));
 sg13g2_buf_4 fanout1235 (.X(net1235),
    .A(net1238));
 sg13g2_buf_4 fanout1236 (.X(net1236),
    .A(net1237));
 sg13g2_buf_4 fanout1237 (.X(net1237),
    .A(net1238));
 sg13g2_buf_1 fanout1238 (.A(net1247),
    .X(net1238));
 sg13g2_buf_4 fanout1239 (.X(net1239),
    .A(net1242));
 sg13g2_buf_4 fanout1240 (.X(net1240),
    .A(net1242));
 sg13g2_buf_2 fanout1241 (.A(net1242),
    .X(net1241));
 sg13g2_buf_1 fanout1242 (.A(net1247),
    .X(net1242));
 sg13g2_buf_4 fanout1243 (.X(net1243),
    .A(net1246));
 sg13g2_buf_4 fanout1244 (.X(net1244),
    .A(net1246));
 sg13g2_buf_2 fanout1245 (.A(net1246),
    .X(net1245));
 sg13g2_buf_2 fanout1246 (.A(net1247),
    .X(net1246));
 sg13g2_buf_1 fanout1247 (.A(net1430),
    .X(net1247));
 sg13g2_buf_4 fanout1248 (.X(net1248),
    .A(net1252));
 sg13g2_buf_4 fanout1249 (.X(net1249),
    .A(net1252));
 sg13g2_buf_4 fanout1250 (.X(net1250),
    .A(net1251));
 sg13g2_buf_4 fanout1251 (.X(net1251),
    .A(net1252));
 sg13g2_buf_2 fanout1252 (.A(net1258),
    .X(net1252));
 sg13g2_buf_4 fanout1253 (.X(net1253),
    .A(net1258));
 sg13g2_buf_2 fanout1254 (.A(net1258),
    .X(net1254));
 sg13g2_buf_4 fanout1255 (.X(net1255),
    .A(net1257));
 sg13g2_buf_4 fanout1256 (.X(net1256),
    .A(net1257));
 sg13g2_buf_2 fanout1257 (.A(net1258),
    .X(net1257));
 sg13g2_buf_1 fanout1258 (.A(net1274),
    .X(net1258));
 sg13g2_buf_4 fanout1259 (.X(net1259),
    .A(net1262));
 sg13g2_buf_4 fanout1260 (.X(net1260),
    .A(net1262));
 sg13g2_buf_2 fanout1261 (.A(net1262),
    .X(net1261));
 sg13g2_buf_2 fanout1262 (.A(net1274),
    .X(net1262));
 sg13g2_buf_4 fanout1263 (.X(net1263),
    .A(net1266));
 sg13g2_buf_2 fanout1264 (.A(net1266),
    .X(net1264));
 sg13g2_buf_4 fanout1265 (.X(net1265),
    .A(net1266));
 sg13g2_buf_1 fanout1266 (.A(net1274),
    .X(net1266));
 sg13g2_buf_4 fanout1267 (.X(net1267),
    .A(net1268));
 sg13g2_buf_4 fanout1268 (.X(net1268),
    .A(net1273));
 sg13g2_buf_4 fanout1269 (.X(net1269),
    .A(net1272));
 sg13g2_buf_4 fanout1270 (.X(net1270),
    .A(net1272));
 sg13g2_buf_2 fanout1271 (.A(net1272),
    .X(net1271));
 sg13g2_buf_2 fanout1272 (.A(net1273),
    .X(net1272));
 sg13g2_buf_2 fanout1273 (.A(net1274),
    .X(net1273));
 sg13g2_buf_1 fanout1274 (.A(net1430),
    .X(net1274));
 sg13g2_buf_4 fanout1275 (.X(net1275),
    .A(net1278));
 sg13g2_buf_4 fanout1276 (.X(net1276),
    .A(net1277));
 sg13g2_buf_4 fanout1277 (.X(net1277),
    .A(net1278));
 sg13g2_buf_2 fanout1278 (.A(net1296),
    .X(net1278));
 sg13g2_buf_4 fanout1279 (.X(net1279),
    .A(net1280));
 sg13g2_buf_4 fanout1280 (.X(net1280),
    .A(net1296));
 sg13g2_buf_4 fanout1281 (.X(net1281),
    .A(net1283));
 sg13g2_buf_4 fanout1282 (.X(net1282),
    .A(net1283));
 sg13g2_buf_2 fanout1283 (.A(net1296),
    .X(net1283));
 sg13g2_buf_4 fanout1284 (.X(net1284),
    .A(net1287));
 sg13g2_buf_4 fanout1285 (.X(net1285),
    .A(net1287));
 sg13g2_buf_2 fanout1286 (.A(net1287),
    .X(net1286));
 sg13g2_buf_2 fanout1287 (.A(net1296),
    .X(net1287));
 sg13g2_buf_4 fanout1288 (.X(net1288),
    .A(net1295));
 sg13g2_buf_2 fanout1289 (.A(net1295),
    .X(net1289));
 sg13g2_buf_4 fanout1290 (.X(net1290),
    .A(net1295));
 sg13g2_buf_4 fanout1291 (.X(net1291),
    .A(net1294));
 sg13g2_buf_4 fanout1292 (.X(net1292),
    .A(net1294));
 sg13g2_buf_2 fanout1293 (.A(net1294),
    .X(net1293));
 sg13g2_buf_1 fanout1294 (.A(net1295),
    .X(net1294));
 sg13g2_buf_1 fanout1295 (.A(net1296),
    .X(net1295));
 sg13g2_buf_1 fanout1296 (.A(net1430),
    .X(net1296));
 sg13g2_buf_4 fanout1297 (.X(net1297),
    .A(net1298));
 sg13g2_buf_4 fanout1298 (.X(net1298),
    .A(net1300));
 sg13g2_buf_4 fanout1299 (.X(net1299),
    .A(net1300));
 sg13g2_buf_2 fanout1300 (.A(net1312),
    .X(net1300));
 sg13g2_buf_4 fanout1301 (.X(net1301),
    .A(net1303));
 sg13g2_buf_4 fanout1302 (.X(net1302),
    .A(net1303));
 sg13g2_buf_2 fanout1303 (.A(net1312),
    .X(net1303));
 sg13g2_buf_4 fanout1304 (.X(net1304),
    .A(net1306));
 sg13g2_buf_4 fanout1305 (.X(net1305),
    .A(net1306));
 sg13g2_buf_2 fanout1306 (.A(net1312),
    .X(net1306));
 sg13g2_buf_4 fanout1307 (.X(net1307),
    .A(net1311));
 sg13g2_buf_2 fanout1308 (.A(net1311),
    .X(net1308));
 sg13g2_buf_4 fanout1309 (.X(net1309),
    .A(net1311));
 sg13g2_buf_2 fanout1310 (.A(net1311),
    .X(net1310));
 sg13g2_buf_1 fanout1311 (.A(net1312),
    .X(net1311));
 sg13g2_buf_1 fanout1312 (.A(net1363),
    .X(net1312));
 sg13g2_buf_4 fanout1313 (.X(net1313),
    .A(net1316));
 sg13g2_buf_2 fanout1314 (.A(net1316),
    .X(net1314));
 sg13g2_buf_4 fanout1315 (.X(net1315),
    .A(net1316));
 sg13g2_buf_2 fanout1316 (.A(net1328),
    .X(net1316));
 sg13g2_buf_4 fanout1317 (.X(net1317),
    .A(net1320));
 sg13g2_buf_2 fanout1318 (.A(net1320),
    .X(net1318));
 sg13g2_buf_4 fanout1319 (.X(net1319),
    .A(net1320));
 sg13g2_buf_2 fanout1320 (.A(net1328),
    .X(net1320));
 sg13g2_buf_4 fanout1321 (.X(net1321),
    .A(net1323));
 sg13g2_buf_4 fanout1322 (.X(net1322),
    .A(net1323));
 sg13g2_buf_2 fanout1323 (.A(net1328),
    .X(net1323));
 sg13g2_buf_4 fanout1324 (.X(net1324),
    .A(net1327));
 sg13g2_buf_4 fanout1325 (.X(net1325),
    .A(net1327));
 sg13g2_buf_2 fanout1326 (.A(net1327),
    .X(net1326));
 sg13g2_buf_2 fanout1327 (.A(net1328),
    .X(net1327));
 sg13g2_buf_1 fanout1328 (.A(net1363),
    .X(net1328));
 sg13g2_buf_4 fanout1329 (.X(net1329),
    .A(net1331));
 sg13g2_buf_4 fanout1330 (.X(net1330),
    .A(net1331));
 sg13g2_buf_2 fanout1331 (.A(net1345),
    .X(net1331));
 sg13g2_buf_4 fanout1332 (.X(net1332),
    .A(net1335));
 sg13g2_buf_4 fanout1333 (.X(net1333),
    .A(net1335));
 sg13g2_buf_2 fanout1334 (.A(net1335),
    .X(net1334));
 sg13g2_buf_1 fanout1335 (.A(net1345),
    .X(net1335));
 sg13g2_buf_4 fanout1336 (.X(net1336),
    .A(net1340));
 sg13g2_buf_2 fanout1337 (.A(net1340),
    .X(net1337));
 sg13g2_buf_4 fanout1338 (.X(net1338),
    .A(net1339));
 sg13g2_buf_4 fanout1339 (.X(net1339),
    .A(net1340));
 sg13g2_buf_1 fanout1340 (.A(net1345),
    .X(net1340));
 sg13g2_buf_4 fanout1341 (.X(net1341),
    .A(net1344));
 sg13g2_buf_4 fanout1342 (.X(net1342),
    .A(net1344));
 sg13g2_buf_4 fanout1343 (.X(net1343),
    .A(net1344));
 sg13g2_buf_2 fanout1344 (.A(net1345),
    .X(net1344));
 sg13g2_buf_1 fanout1345 (.A(net1363),
    .X(net1345));
 sg13g2_buf_4 fanout1346 (.X(net1346),
    .A(net1348));
 sg13g2_buf_4 fanout1347 (.X(net1347),
    .A(net1348));
 sg13g2_buf_2 fanout1348 (.A(net1362),
    .X(net1348));
 sg13g2_buf_4 fanout1349 (.X(net1349),
    .A(net1353));
 sg13g2_buf_2 fanout1350 (.A(net1353),
    .X(net1350));
 sg13g2_buf_4 fanout1351 (.X(net1351),
    .A(net1353));
 sg13g2_buf_2 fanout1352 (.A(net1353),
    .X(net1352));
 sg13g2_buf_1 fanout1353 (.A(net1362),
    .X(net1353));
 sg13g2_buf_4 fanout1354 (.X(net1354),
    .A(net1357));
 sg13g2_buf_4 fanout1355 (.X(net1355),
    .A(net1357));
 sg13g2_buf_2 fanout1356 (.A(net1357),
    .X(net1356));
 sg13g2_buf_1 fanout1357 (.A(net1362),
    .X(net1357));
 sg13g2_buf_4 fanout1358 (.X(net1358),
    .A(net1361));
 sg13g2_buf_4 fanout1359 (.X(net1359),
    .A(net1361));
 sg13g2_buf_4 fanout1360 (.X(net1360),
    .A(net1361));
 sg13g2_buf_2 fanout1361 (.A(net1362),
    .X(net1361));
 sg13g2_buf_1 fanout1362 (.A(net1363),
    .X(net1362));
 sg13g2_buf_1 fanout1363 (.A(net1430),
    .X(net1363));
 sg13g2_buf_4 fanout1364 (.X(net1364),
    .A(net1370));
 sg13g2_buf_4 fanout1365 (.X(net1365),
    .A(net1370));
 sg13g2_buf_4 fanout1366 (.X(net1366),
    .A(net1369));
 sg13g2_buf_2 fanout1367 (.A(net1369),
    .X(net1367));
 sg13g2_buf_4 fanout1368 (.X(net1368),
    .A(net1369));
 sg13g2_buf_2 fanout1369 (.A(net1370),
    .X(net1369));
 sg13g2_buf_2 fanout1370 (.A(net1394),
    .X(net1370));
 sg13g2_buf_4 fanout1371 (.X(net1371),
    .A(net1374));
 sg13g2_buf_4 fanout1372 (.X(net1372),
    .A(net1374));
 sg13g2_buf_2 fanout1373 (.A(net1374),
    .X(net1373));
 sg13g2_buf_1 fanout1374 (.A(net1394),
    .X(net1374));
 sg13g2_buf_4 fanout1375 (.X(net1375),
    .A(net1377));
 sg13g2_buf_4 fanout1376 (.X(net1376),
    .A(net1377));
 sg13g2_buf_2 fanout1377 (.A(net1394),
    .X(net1377));
 sg13g2_buf_4 fanout1378 (.X(net1378),
    .A(net1380));
 sg13g2_buf_4 fanout1379 (.X(net1379),
    .A(net1380));
 sg13g2_buf_4 fanout1380 (.X(net1380),
    .A(net1385));
 sg13g2_buf_4 fanout1381 (.X(net1381),
    .A(net1385));
 sg13g2_buf_2 fanout1382 (.A(net1385),
    .X(net1382));
 sg13g2_buf_4 fanout1383 (.X(net1383),
    .A(net1384));
 sg13g2_buf_4 fanout1384 (.X(net1384),
    .A(net1385));
 sg13g2_buf_1 fanout1385 (.A(net1394),
    .X(net1385));
 sg13g2_buf_4 fanout1386 (.X(net1386),
    .A(net1389));
 sg13g2_buf_2 fanout1387 (.A(net1389),
    .X(net1387));
 sg13g2_buf_4 fanout1388 (.X(net1388),
    .A(net1389));
 sg13g2_buf_2 fanout1389 (.A(net1394),
    .X(net1389));
 sg13g2_buf_4 fanout1390 (.X(net1390),
    .A(net1393));
 sg13g2_buf_2 fanout1391 (.A(net1393),
    .X(net1391));
 sg13g2_buf_4 fanout1392 (.X(net1392),
    .A(net1393));
 sg13g2_buf_2 fanout1393 (.A(net1394),
    .X(net1393));
 sg13g2_buf_1 fanout1394 (.A(net1430),
    .X(net1394));
 sg13g2_buf_4 fanout1395 (.X(net1395),
    .A(net1398));
 sg13g2_buf_4 fanout1396 (.X(net1396),
    .A(net1398));
 sg13g2_buf_2 fanout1397 (.A(net1398),
    .X(net1397));
 sg13g2_buf_2 fanout1398 (.A(net1401),
    .X(net1398));
 sg13g2_buf_4 fanout1399 (.X(net1399),
    .A(net1401));
 sg13g2_buf_4 fanout1400 (.X(net1400),
    .A(net1401));
 sg13g2_buf_2 fanout1401 (.A(net1429),
    .X(net1401));
 sg13g2_buf_4 fanout1402 (.X(net1402),
    .A(net1406));
 sg13g2_buf_2 fanout1403 (.A(net1406),
    .X(net1403));
 sg13g2_buf_4 fanout1404 (.X(net1404),
    .A(net1406));
 sg13g2_buf_2 fanout1405 (.A(net1406),
    .X(net1405));
 sg13g2_buf_1 fanout1406 (.A(net1429),
    .X(net1406));
 sg13g2_buf_4 fanout1407 (.X(net1407),
    .A(net1410));
 sg13g2_buf_4 fanout1408 (.X(net1408),
    .A(net1410));
 sg13g2_buf_2 fanout1409 (.A(net1410),
    .X(net1409));
 sg13g2_buf_2 fanout1410 (.A(net1429),
    .X(net1410));
 sg13g2_buf_4 fanout1411 (.X(net1411),
    .A(net1415));
 sg13g2_buf_2 fanout1412 (.A(net1415),
    .X(net1412));
 sg13g2_buf_4 fanout1413 (.X(net1413),
    .A(net1415));
 sg13g2_buf_2 fanout1414 (.A(net1415),
    .X(net1414));
 sg13g2_buf_1 fanout1415 (.A(net1428),
    .X(net1415));
 sg13g2_buf_4 fanout1416 (.X(net1416),
    .A(net1420));
 sg13g2_buf_2 fanout1417 (.A(net1420),
    .X(net1417));
 sg13g2_buf_4 fanout1418 (.X(net1418),
    .A(net1420));
 sg13g2_buf_2 fanout1419 (.A(net1420),
    .X(net1419));
 sg13g2_buf_1 fanout1420 (.A(net1428),
    .X(net1420));
 sg13g2_buf_4 fanout1421 (.X(net1421),
    .A(net1423));
 sg13g2_buf_4 fanout1422 (.X(net1422),
    .A(net1423));
 sg13g2_buf_4 fanout1423 (.X(net1423),
    .A(net1428));
 sg13g2_buf_4 fanout1424 (.X(net1424),
    .A(net1427));
 sg13g2_buf_2 fanout1425 (.A(net1427),
    .X(net1425));
 sg13g2_buf_4 fanout1426 (.X(net1426),
    .A(net1427));
 sg13g2_buf_1 fanout1427 (.A(net1428),
    .X(net1427));
 sg13g2_buf_1 fanout1428 (.A(net1429),
    .X(net1428));
 sg13g2_buf_1 fanout1429 (.A(net1430),
    .X(net1429));
 sg13g2_buf_2 fanout1430 (.A(net1),
    .X(net1430));
 sg13g2_tiehi _24629__1431 (.L_HI(net1431));
 sg13g2_tiehi _24630__1432 (.L_HI(net1432));
 sg13g2_tiehi _24631__1433 (.L_HI(net1433));
 sg13g2_tiehi _24632__1434 (.L_HI(net1434));
 sg13g2_tiehi _24633__1435 (.L_HI(net1435));
 sg13g2_tiehi _24634__1436 (.L_HI(net1436));
 sg13g2_tiehi _24635__1437 (.L_HI(net1437));
 sg13g2_tiehi _24636__1438 (.L_HI(net1438));
 sg13g2_tiehi \top_ihp.oisc.mem_addr_lowbits[0]$_DFF_P__1439  (.L_HI(net1439));
 sg13g2_tiehi \top_ihp.oisc.mem_addr_lowbits[1]$_DFF_P__1440  (.L_HI(net1440));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[0]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[1]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[2]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[3]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[4]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[5]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[6]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[7]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \top_ihp.oisc.regs[16][0]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \top_ihp.oisc.regs[16][10]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \top_ihp.oisc.regs[16][11]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \top_ihp.oisc.regs[16][12]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \top_ihp.oisc.regs[16][13]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \top_ihp.oisc.regs[16][14]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \top_ihp.oisc.regs[16][15]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \top_ihp.oisc.regs[16][16]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \top_ihp.oisc.regs[16][17]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \top_ihp.oisc.regs[16][18]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \top_ihp.oisc.regs[16][19]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \top_ihp.oisc.regs[16][1]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \top_ihp.oisc.regs[16][20]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \top_ihp.oisc.regs[16][21]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \top_ihp.oisc.regs[16][22]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \top_ihp.oisc.regs[16][23]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \top_ihp.oisc.regs[16][24]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \top_ihp.oisc.regs[16][25]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \top_ihp.oisc.regs[16][26]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \top_ihp.oisc.regs[16][27]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \top_ihp.oisc.regs[16][28]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \top_ihp.oisc.regs[16][29]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \top_ihp.oisc.regs[16][2]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \top_ihp.oisc.regs[16][30]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \top_ihp.oisc.regs[16][31]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \top_ihp.oisc.regs[16][3]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \top_ihp.oisc.regs[16][4]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \top_ihp.oisc.regs[16][5]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \top_ihp.oisc.regs[16][6]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \top_ihp.oisc.regs[16][7]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \top_ihp.oisc.regs[16][8]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \top_ihp.oisc.regs[16][9]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \top_ihp.oisc.regs[17][0]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \top_ihp.oisc.regs[17][10]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \top_ihp.oisc.regs[17][11]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \top_ihp.oisc.regs[17][12]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \top_ihp.oisc.regs[17][13]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \top_ihp.oisc.regs[17][14]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \top_ihp.oisc.regs[17][15]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \top_ihp.oisc.regs[17][16]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \top_ihp.oisc.regs[17][17]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \top_ihp.oisc.regs[17][18]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \top_ihp.oisc.regs[17][19]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \top_ihp.oisc.regs[17][1]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \top_ihp.oisc.regs[17][20]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \top_ihp.oisc.regs[17][21]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \top_ihp.oisc.regs[17][22]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \top_ihp.oisc.regs[17][23]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \top_ihp.oisc.regs[17][24]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \top_ihp.oisc.regs[17][25]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \top_ihp.oisc.regs[17][26]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \top_ihp.oisc.regs[17][27]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \top_ihp.oisc.regs[17][28]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \top_ihp.oisc.regs[17][29]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \top_ihp.oisc.regs[17][2]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \top_ihp.oisc.regs[17][30]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \top_ihp.oisc.regs[17][31]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \top_ihp.oisc.regs[17][3]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \top_ihp.oisc.regs[17][4]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \top_ihp.oisc.regs[17][5]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \top_ihp.oisc.regs[17][6]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \top_ihp.oisc.regs[17][7]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \top_ihp.oisc.regs[17][8]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \top_ihp.oisc.regs[17][9]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \top_ihp.oisc.regs[18][0]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \top_ihp.oisc.regs[18][10]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \top_ihp.oisc.regs[18][11]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \top_ihp.oisc.regs[18][12]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \top_ihp.oisc.regs[18][13]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \top_ihp.oisc.regs[18][14]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \top_ihp.oisc.regs[18][15]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \top_ihp.oisc.regs[18][16]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \top_ihp.oisc.regs[18][17]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \top_ihp.oisc.regs[18][18]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \top_ihp.oisc.regs[18][19]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \top_ihp.oisc.regs[18][1]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \top_ihp.oisc.regs[18][20]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \top_ihp.oisc.regs[18][21]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \top_ihp.oisc.regs[18][22]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \top_ihp.oisc.regs[18][23]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \top_ihp.oisc.regs[18][24]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \top_ihp.oisc.regs[18][25]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \top_ihp.oisc.regs[18][26]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \top_ihp.oisc.regs[18][27]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \top_ihp.oisc.regs[18][28]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \top_ihp.oisc.regs[18][29]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \top_ihp.oisc.regs[18][2]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \top_ihp.oisc.regs[18][30]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \top_ihp.oisc.regs[18][31]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \top_ihp.oisc.regs[18][3]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \top_ihp.oisc.regs[18][4]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \top_ihp.oisc.regs[18][5]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \top_ihp.oisc.regs[18][6]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \top_ihp.oisc.regs[18][7]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \top_ihp.oisc.regs[18][8]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \top_ihp.oisc.regs[18][9]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \top_ihp.oisc.regs[19][0]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \top_ihp.oisc.regs[19][10]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \top_ihp.oisc.regs[19][11]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \top_ihp.oisc.regs[19][12]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \top_ihp.oisc.regs[19][13]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \top_ihp.oisc.regs[19][14]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \top_ihp.oisc.regs[19][15]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \top_ihp.oisc.regs[19][16]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \top_ihp.oisc.regs[19][17]$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \top_ihp.oisc.regs[19][18]$_DFFE_PP__1554  (.L_HI(net1554));
 sg13g2_tiehi \top_ihp.oisc.regs[19][19]$_DFFE_PP__1555  (.L_HI(net1555));
 sg13g2_tiehi \top_ihp.oisc.regs[19][1]$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \top_ihp.oisc.regs[19][20]$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \top_ihp.oisc.regs[19][21]$_DFFE_PP__1558  (.L_HI(net1558));
 sg13g2_tiehi \top_ihp.oisc.regs[19][22]$_DFFE_PP__1559  (.L_HI(net1559));
 sg13g2_tiehi \top_ihp.oisc.regs[19][23]$_DFFE_PP__1560  (.L_HI(net1560));
 sg13g2_tiehi \top_ihp.oisc.regs[19][24]$_DFFE_PP__1561  (.L_HI(net1561));
 sg13g2_tiehi \top_ihp.oisc.regs[19][25]$_DFFE_PP__1562  (.L_HI(net1562));
 sg13g2_tiehi \top_ihp.oisc.regs[19][26]$_DFFE_PP__1563  (.L_HI(net1563));
 sg13g2_tiehi \top_ihp.oisc.regs[19][27]$_DFFE_PP__1564  (.L_HI(net1564));
 sg13g2_tiehi \top_ihp.oisc.regs[19][28]$_DFFE_PP__1565  (.L_HI(net1565));
 sg13g2_tiehi \top_ihp.oisc.regs[19][29]$_DFFE_PP__1566  (.L_HI(net1566));
 sg13g2_tiehi \top_ihp.oisc.regs[19][2]$_DFFE_PP__1567  (.L_HI(net1567));
 sg13g2_tiehi \top_ihp.oisc.regs[19][30]$_DFFE_PP__1568  (.L_HI(net1568));
 sg13g2_tiehi \top_ihp.oisc.regs[19][31]$_DFFE_PP__1569  (.L_HI(net1569));
 sg13g2_tiehi \top_ihp.oisc.regs[19][3]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \top_ihp.oisc.regs[19][4]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \top_ihp.oisc.regs[19][5]$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \top_ihp.oisc.regs[19][6]$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \top_ihp.oisc.regs[19][7]$_DFFE_PP__1574  (.L_HI(net1574));
 sg13g2_tiehi \top_ihp.oisc.regs[19][8]$_DFFE_PP__1575  (.L_HI(net1575));
 sg13g2_tiehi \top_ihp.oisc.regs[19][9]$_DFFE_PP__1576  (.L_HI(net1576));
 sg13g2_tiehi \top_ihp.oisc.regs[20][0]$_DFFE_PP__1577  (.L_HI(net1577));
 sg13g2_tiehi \top_ihp.oisc.regs[20][10]$_DFFE_PP__1578  (.L_HI(net1578));
 sg13g2_tiehi \top_ihp.oisc.regs[20][11]$_DFFE_PP__1579  (.L_HI(net1579));
 sg13g2_tiehi \top_ihp.oisc.regs[20][12]$_DFFE_PP__1580  (.L_HI(net1580));
 sg13g2_tiehi \top_ihp.oisc.regs[20][13]$_DFFE_PP__1581  (.L_HI(net1581));
 sg13g2_tiehi \top_ihp.oisc.regs[20][14]$_DFFE_PP__1582  (.L_HI(net1582));
 sg13g2_tiehi \top_ihp.oisc.regs[20][15]$_DFFE_PP__1583  (.L_HI(net1583));
 sg13g2_tiehi \top_ihp.oisc.regs[20][16]$_DFFE_PP__1584  (.L_HI(net1584));
 sg13g2_tiehi \top_ihp.oisc.regs[20][17]$_DFFE_PP__1585  (.L_HI(net1585));
 sg13g2_tiehi \top_ihp.oisc.regs[20][18]$_DFFE_PP__1586  (.L_HI(net1586));
 sg13g2_tiehi \top_ihp.oisc.regs[20][19]$_DFFE_PP__1587  (.L_HI(net1587));
 sg13g2_tiehi \top_ihp.oisc.regs[20][1]$_DFFE_PP__1588  (.L_HI(net1588));
 sg13g2_tiehi \top_ihp.oisc.regs[20][20]$_DFFE_PP__1589  (.L_HI(net1589));
 sg13g2_tiehi \top_ihp.oisc.regs[20][21]$_DFFE_PP__1590  (.L_HI(net1590));
 sg13g2_tiehi \top_ihp.oisc.regs[20][22]$_DFFE_PP__1591  (.L_HI(net1591));
 sg13g2_tiehi \top_ihp.oisc.regs[20][23]$_DFFE_PP__1592  (.L_HI(net1592));
 sg13g2_tiehi \top_ihp.oisc.regs[20][24]$_DFFE_PP__1593  (.L_HI(net1593));
 sg13g2_tiehi \top_ihp.oisc.regs[20][25]$_DFFE_PP__1594  (.L_HI(net1594));
 sg13g2_tiehi \top_ihp.oisc.regs[20][26]$_DFFE_PP__1595  (.L_HI(net1595));
 sg13g2_tiehi \top_ihp.oisc.regs[20][27]$_DFFE_PP__1596  (.L_HI(net1596));
 sg13g2_tiehi \top_ihp.oisc.regs[20][28]$_DFFE_PP__1597  (.L_HI(net1597));
 sg13g2_tiehi \top_ihp.oisc.regs[20][29]$_DFFE_PP__1598  (.L_HI(net1598));
 sg13g2_tiehi \top_ihp.oisc.regs[20][2]$_DFFE_PP__1599  (.L_HI(net1599));
 sg13g2_tiehi \top_ihp.oisc.regs[20][30]$_DFFE_PP__1600  (.L_HI(net1600));
 sg13g2_tiehi \top_ihp.oisc.regs[20][31]$_DFFE_PP__1601  (.L_HI(net1601));
 sg13g2_tiehi \top_ihp.oisc.regs[20][3]$_DFFE_PP__1602  (.L_HI(net1602));
 sg13g2_tiehi \top_ihp.oisc.regs[20][4]$_DFFE_PP__1603  (.L_HI(net1603));
 sg13g2_tiehi \top_ihp.oisc.regs[20][5]$_DFFE_PP__1604  (.L_HI(net1604));
 sg13g2_tiehi \top_ihp.oisc.regs[20][6]$_DFFE_PP__1605  (.L_HI(net1605));
 sg13g2_tiehi \top_ihp.oisc.regs[20][7]$_DFFE_PP__1606  (.L_HI(net1606));
 sg13g2_tiehi \top_ihp.oisc.regs[20][8]$_DFFE_PP__1607  (.L_HI(net1607));
 sg13g2_tiehi \top_ihp.oisc.regs[20][9]$_DFFE_PP__1608  (.L_HI(net1608));
 sg13g2_tiehi \top_ihp.oisc.regs[21][0]$_DFFE_PP__1609  (.L_HI(net1609));
 sg13g2_tiehi \top_ihp.oisc.regs[21][10]$_DFFE_PP__1610  (.L_HI(net1610));
 sg13g2_tiehi \top_ihp.oisc.regs[21][11]$_DFFE_PP__1611  (.L_HI(net1611));
 sg13g2_tiehi \top_ihp.oisc.regs[21][12]$_DFFE_PP__1612  (.L_HI(net1612));
 sg13g2_tiehi \top_ihp.oisc.regs[21][13]$_DFFE_PP__1613  (.L_HI(net1613));
 sg13g2_tiehi \top_ihp.oisc.regs[21][14]$_DFFE_PP__1614  (.L_HI(net1614));
 sg13g2_tiehi \top_ihp.oisc.regs[21][15]$_DFFE_PP__1615  (.L_HI(net1615));
 sg13g2_tiehi \top_ihp.oisc.regs[21][16]$_DFFE_PP__1616  (.L_HI(net1616));
 sg13g2_tiehi \top_ihp.oisc.regs[21][17]$_DFFE_PP__1617  (.L_HI(net1617));
 sg13g2_tiehi \top_ihp.oisc.regs[21][18]$_DFFE_PP__1618  (.L_HI(net1618));
 sg13g2_tiehi \top_ihp.oisc.regs[21][19]$_DFFE_PP__1619  (.L_HI(net1619));
 sg13g2_tiehi \top_ihp.oisc.regs[21][1]$_DFFE_PP__1620  (.L_HI(net1620));
 sg13g2_tiehi \top_ihp.oisc.regs[21][20]$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \top_ihp.oisc.regs[21][21]$_DFFE_PP__1622  (.L_HI(net1622));
 sg13g2_tiehi \top_ihp.oisc.regs[21][22]$_DFFE_PP__1623  (.L_HI(net1623));
 sg13g2_tiehi \top_ihp.oisc.regs[21][23]$_DFFE_PP__1624  (.L_HI(net1624));
 sg13g2_tiehi \top_ihp.oisc.regs[21][24]$_DFFE_PP__1625  (.L_HI(net1625));
 sg13g2_tiehi \top_ihp.oisc.regs[21][25]$_DFFE_PP__1626  (.L_HI(net1626));
 sg13g2_tiehi \top_ihp.oisc.regs[21][26]$_DFFE_PP__1627  (.L_HI(net1627));
 sg13g2_tiehi \top_ihp.oisc.regs[21][27]$_DFFE_PP__1628  (.L_HI(net1628));
 sg13g2_tiehi \top_ihp.oisc.regs[21][28]$_DFFE_PP__1629  (.L_HI(net1629));
 sg13g2_tiehi \top_ihp.oisc.regs[21][29]$_DFFE_PP__1630  (.L_HI(net1630));
 sg13g2_tiehi \top_ihp.oisc.regs[21][2]$_DFFE_PP__1631  (.L_HI(net1631));
 sg13g2_tiehi \top_ihp.oisc.regs[21][30]$_DFFE_PP__1632  (.L_HI(net1632));
 sg13g2_tiehi \top_ihp.oisc.regs[21][31]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \top_ihp.oisc.regs[21][3]$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \top_ihp.oisc.regs[21][4]$_DFFE_PP__1635  (.L_HI(net1635));
 sg13g2_tiehi \top_ihp.oisc.regs[21][5]$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \top_ihp.oisc.regs[21][6]$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \top_ihp.oisc.regs[21][7]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \top_ihp.oisc.regs[21][8]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \top_ihp.oisc.regs[21][9]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \top_ihp.oisc.regs[22][0]$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \top_ihp.oisc.regs[22][10]$_DFFE_PP__1642  (.L_HI(net1642));
 sg13g2_tiehi \top_ihp.oisc.regs[22][11]$_DFFE_PP__1643  (.L_HI(net1643));
 sg13g2_tiehi \top_ihp.oisc.regs[22][12]$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \top_ihp.oisc.regs[22][13]$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \top_ihp.oisc.regs[22][14]$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \top_ihp.oisc.regs[22][15]$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \top_ihp.oisc.regs[22][16]$_DFFE_PP__1648  (.L_HI(net1648));
 sg13g2_tiehi \top_ihp.oisc.regs[22][17]$_DFFE_PP__1649  (.L_HI(net1649));
 sg13g2_tiehi \top_ihp.oisc.regs[22][18]$_DFFE_PP__1650  (.L_HI(net1650));
 sg13g2_tiehi \top_ihp.oisc.regs[22][19]$_DFFE_PP__1651  (.L_HI(net1651));
 sg13g2_tiehi \top_ihp.oisc.regs[22][1]$_DFFE_PP__1652  (.L_HI(net1652));
 sg13g2_tiehi \top_ihp.oisc.regs[22][20]$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \top_ihp.oisc.regs[22][21]$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \top_ihp.oisc.regs[22][22]$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \top_ihp.oisc.regs[22][23]$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \top_ihp.oisc.regs[22][24]$_DFFE_PP__1657  (.L_HI(net1657));
 sg13g2_tiehi \top_ihp.oisc.regs[22][25]$_DFFE_PP__1658  (.L_HI(net1658));
 sg13g2_tiehi \top_ihp.oisc.regs[22][26]$_DFFE_PP__1659  (.L_HI(net1659));
 sg13g2_tiehi \top_ihp.oisc.regs[22][27]$_DFFE_PP__1660  (.L_HI(net1660));
 sg13g2_tiehi \top_ihp.oisc.regs[22][28]$_DFFE_PP__1661  (.L_HI(net1661));
 sg13g2_tiehi \top_ihp.oisc.regs[22][29]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \top_ihp.oisc.regs[22][2]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \top_ihp.oisc.regs[22][30]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \top_ihp.oisc.regs[22][31]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \top_ihp.oisc.regs[22][3]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \top_ihp.oisc.regs[22][4]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \top_ihp.oisc.regs[22][5]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \top_ihp.oisc.regs[22][6]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \top_ihp.oisc.regs[22][7]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \top_ihp.oisc.regs[22][8]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \top_ihp.oisc.regs[22][9]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \top_ihp.oisc.regs[23][0]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \top_ihp.oisc.regs[23][10]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \top_ihp.oisc.regs[23][11]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \top_ihp.oisc.regs[23][12]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \top_ihp.oisc.regs[23][13]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \top_ihp.oisc.regs[23][14]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \top_ihp.oisc.regs[23][15]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \top_ihp.oisc.regs[23][16]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \top_ihp.oisc.regs[23][17]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \top_ihp.oisc.regs[23][18]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \top_ihp.oisc.regs[23][19]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \top_ihp.oisc.regs[23][1]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \top_ihp.oisc.regs[23][20]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \top_ihp.oisc.regs[23][21]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \top_ihp.oisc.regs[23][22]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \top_ihp.oisc.regs[23][23]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \top_ihp.oisc.regs[23][24]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \top_ihp.oisc.regs[23][25]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \top_ihp.oisc.regs[23][26]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \top_ihp.oisc.regs[23][27]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \top_ihp.oisc.regs[23][28]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \top_ihp.oisc.regs[23][29]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \top_ihp.oisc.regs[23][2]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \top_ihp.oisc.regs[23][30]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \top_ihp.oisc.regs[23][31]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \top_ihp.oisc.regs[23][3]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \top_ihp.oisc.regs[23][4]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \top_ihp.oisc.regs[23][5]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \top_ihp.oisc.regs[23][6]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \top_ihp.oisc.regs[23][7]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \top_ihp.oisc.regs[23][8]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \top_ihp.oisc.regs[23][9]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \top_ihp.oisc.regs[24][0]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \top_ihp.oisc.regs[24][10]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \top_ihp.oisc.regs[24][11]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \top_ihp.oisc.regs[24][12]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \top_ihp.oisc.regs[24][13]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \top_ihp.oisc.regs[24][14]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \top_ihp.oisc.regs[24][15]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \top_ihp.oisc.regs[24][16]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \top_ihp.oisc.regs[24][17]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \top_ihp.oisc.regs[24][18]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \top_ihp.oisc.regs[24][19]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \top_ihp.oisc.regs[24][1]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \top_ihp.oisc.regs[24][20]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \top_ihp.oisc.regs[24][21]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \top_ihp.oisc.regs[24][22]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \top_ihp.oisc.regs[24][23]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \top_ihp.oisc.regs[24][24]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \top_ihp.oisc.regs[24][25]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \top_ihp.oisc.regs[24][26]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \top_ihp.oisc.regs[24][27]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \top_ihp.oisc.regs[24][28]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \top_ihp.oisc.regs[24][29]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \top_ihp.oisc.regs[24][2]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \top_ihp.oisc.regs[24][30]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \top_ihp.oisc.regs[24][31]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \top_ihp.oisc.regs[24][3]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \top_ihp.oisc.regs[24][4]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \top_ihp.oisc.regs[24][5]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \top_ihp.oisc.regs[24][6]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \top_ihp.oisc.regs[24][7]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \top_ihp.oisc.regs[24][8]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \top_ihp.oisc.regs[24][9]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \top_ihp.oisc.regs[25][0]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \top_ihp.oisc.regs[25][10]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \top_ihp.oisc.regs[25][11]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \top_ihp.oisc.regs[25][12]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \top_ihp.oisc.regs[25][13]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \top_ihp.oisc.regs[25][14]$_DFFE_PP__1742  (.L_HI(net1742));
 sg13g2_tiehi \top_ihp.oisc.regs[25][15]$_DFFE_PP__1743  (.L_HI(net1743));
 sg13g2_tiehi \top_ihp.oisc.regs[25][16]$_DFFE_PP__1744  (.L_HI(net1744));
 sg13g2_tiehi \top_ihp.oisc.regs[25][17]$_DFFE_PP__1745  (.L_HI(net1745));
 sg13g2_tiehi \top_ihp.oisc.regs[25][18]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \top_ihp.oisc.regs[25][19]$_DFFE_PP__1747  (.L_HI(net1747));
 sg13g2_tiehi \top_ihp.oisc.regs[25][1]$_DFFE_PP__1748  (.L_HI(net1748));
 sg13g2_tiehi \top_ihp.oisc.regs[25][20]$_DFFE_PP__1749  (.L_HI(net1749));
 sg13g2_tiehi \top_ihp.oisc.regs[25][21]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \top_ihp.oisc.regs[25][22]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \top_ihp.oisc.regs[25][23]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \top_ihp.oisc.regs[25][24]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \top_ihp.oisc.regs[25][25]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \top_ihp.oisc.regs[25][26]$_DFFE_PP__1755  (.L_HI(net1755));
 sg13g2_tiehi \top_ihp.oisc.regs[25][27]$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \top_ihp.oisc.regs[25][28]$_DFFE_PP__1757  (.L_HI(net1757));
 sg13g2_tiehi \top_ihp.oisc.regs[25][29]$_DFFE_PP__1758  (.L_HI(net1758));
 sg13g2_tiehi \top_ihp.oisc.regs[25][2]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \top_ihp.oisc.regs[25][30]$_DFFE_PP__1760  (.L_HI(net1760));
 sg13g2_tiehi \top_ihp.oisc.regs[25][31]$_DFFE_PP__1761  (.L_HI(net1761));
 sg13g2_tiehi \top_ihp.oisc.regs[25][3]$_DFFE_PP__1762  (.L_HI(net1762));
 sg13g2_tiehi \top_ihp.oisc.regs[25][4]$_DFFE_PP__1763  (.L_HI(net1763));
 sg13g2_tiehi \top_ihp.oisc.regs[25][5]$_DFFE_PP__1764  (.L_HI(net1764));
 sg13g2_tiehi \top_ihp.oisc.regs[25][6]$_DFFE_PP__1765  (.L_HI(net1765));
 sg13g2_tiehi \top_ihp.oisc.regs[25][7]$_DFFE_PP__1766  (.L_HI(net1766));
 sg13g2_tiehi \top_ihp.oisc.regs[25][8]$_DFFE_PP__1767  (.L_HI(net1767));
 sg13g2_tiehi \top_ihp.oisc.regs[25][9]$_DFFE_PP__1768  (.L_HI(net1768));
 sg13g2_tiehi \top_ihp.oisc.regs[26][0]$_DFFE_PP__1769  (.L_HI(net1769));
 sg13g2_tiehi \top_ihp.oisc.regs[26][10]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \top_ihp.oisc.regs[26][11]$_DFFE_PP__1771  (.L_HI(net1771));
 sg13g2_tiehi \top_ihp.oisc.regs[26][12]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \top_ihp.oisc.regs[26][13]$_DFFE_PP__1773  (.L_HI(net1773));
 sg13g2_tiehi \top_ihp.oisc.regs[26][14]$_DFFE_PP__1774  (.L_HI(net1774));
 sg13g2_tiehi \top_ihp.oisc.regs[26][15]$_DFFE_PP__1775  (.L_HI(net1775));
 sg13g2_tiehi \top_ihp.oisc.regs[26][16]$_DFFE_PP__1776  (.L_HI(net1776));
 sg13g2_tiehi \top_ihp.oisc.regs[26][17]$_DFFE_PP__1777  (.L_HI(net1777));
 sg13g2_tiehi \top_ihp.oisc.regs[26][18]$_DFFE_PP__1778  (.L_HI(net1778));
 sg13g2_tiehi \top_ihp.oisc.regs[26][19]$_DFFE_PP__1779  (.L_HI(net1779));
 sg13g2_tiehi \top_ihp.oisc.regs[26][1]$_DFFE_PP__1780  (.L_HI(net1780));
 sg13g2_tiehi \top_ihp.oisc.regs[26][20]$_DFFE_PP__1781  (.L_HI(net1781));
 sg13g2_tiehi \top_ihp.oisc.regs[26][21]$_DFFE_PP__1782  (.L_HI(net1782));
 sg13g2_tiehi \top_ihp.oisc.regs[26][22]$_DFFE_PP__1783  (.L_HI(net1783));
 sg13g2_tiehi \top_ihp.oisc.regs[26][23]$_DFFE_PP__1784  (.L_HI(net1784));
 sg13g2_tiehi \top_ihp.oisc.regs[26][24]$_DFFE_PP__1785  (.L_HI(net1785));
 sg13g2_tiehi \top_ihp.oisc.regs[26][25]$_DFFE_PP__1786  (.L_HI(net1786));
 sg13g2_tiehi \top_ihp.oisc.regs[26][26]$_DFFE_PP__1787  (.L_HI(net1787));
 sg13g2_tiehi \top_ihp.oisc.regs[26][27]$_DFFE_PP__1788  (.L_HI(net1788));
 sg13g2_tiehi \top_ihp.oisc.regs[26][28]$_DFFE_PP__1789  (.L_HI(net1789));
 sg13g2_tiehi \top_ihp.oisc.regs[26][29]$_DFFE_PP__1790  (.L_HI(net1790));
 sg13g2_tiehi \top_ihp.oisc.regs[26][2]$_DFFE_PP__1791  (.L_HI(net1791));
 sg13g2_tiehi \top_ihp.oisc.regs[26][30]$_DFFE_PP__1792  (.L_HI(net1792));
 sg13g2_tiehi \top_ihp.oisc.regs[26][31]$_DFFE_PP__1793  (.L_HI(net1793));
 sg13g2_tiehi \top_ihp.oisc.regs[26][3]$_DFFE_PP__1794  (.L_HI(net1794));
 sg13g2_tiehi \top_ihp.oisc.regs[26][4]$_DFFE_PP__1795  (.L_HI(net1795));
 sg13g2_tiehi \top_ihp.oisc.regs[26][5]$_DFFE_PP__1796  (.L_HI(net1796));
 sg13g2_tiehi \top_ihp.oisc.regs[26][6]$_DFFE_PP__1797  (.L_HI(net1797));
 sg13g2_tiehi \top_ihp.oisc.regs[26][7]$_DFFE_PP__1798  (.L_HI(net1798));
 sg13g2_tiehi \top_ihp.oisc.regs[26][8]$_DFFE_PP__1799  (.L_HI(net1799));
 sg13g2_tiehi \top_ihp.oisc.regs[26][9]$_DFFE_PP__1800  (.L_HI(net1800));
 sg13g2_tiehi \top_ihp.oisc.regs[27][0]$_DFFE_PP__1801  (.L_HI(net1801));
 sg13g2_tiehi \top_ihp.oisc.regs[27][10]$_DFFE_PP__1802  (.L_HI(net1802));
 sg13g2_tiehi \top_ihp.oisc.regs[27][11]$_DFFE_PP__1803  (.L_HI(net1803));
 sg13g2_tiehi \top_ihp.oisc.regs[27][12]$_DFFE_PP__1804  (.L_HI(net1804));
 sg13g2_tiehi \top_ihp.oisc.regs[27][13]$_DFFE_PP__1805  (.L_HI(net1805));
 sg13g2_tiehi \top_ihp.oisc.regs[27][14]$_DFFE_PP__1806  (.L_HI(net1806));
 sg13g2_tiehi \top_ihp.oisc.regs[27][15]$_DFFE_PP__1807  (.L_HI(net1807));
 sg13g2_tiehi \top_ihp.oisc.regs[27][16]$_DFFE_PP__1808  (.L_HI(net1808));
 sg13g2_tiehi \top_ihp.oisc.regs[27][17]$_DFFE_PP__1809  (.L_HI(net1809));
 sg13g2_tiehi \top_ihp.oisc.regs[27][18]$_DFFE_PP__1810  (.L_HI(net1810));
 sg13g2_tiehi \top_ihp.oisc.regs[27][19]$_DFFE_PP__1811  (.L_HI(net1811));
 sg13g2_tiehi \top_ihp.oisc.regs[27][1]$_DFFE_PP__1812  (.L_HI(net1812));
 sg13g2_tiehi \top_ihp.oisc.regs[27][20]$_DFFE_PP__1813  (.L_HI(net1813));
 sg13g2_tiehi \top_ihp.oisc.regs[27][21]$_DFFE_PP__1814  (.L_HI(net1814));
 sg13g2_tiehi \top_ihp.oisc.regs[27][22]$_DFFE_PP__1815  (.L_HI(net1815));
 sg13g2_tiehi \top_ihp.oisc.regs[27][23]$_DFFE_PP__1816  (.L_HI(net1816));
 sg13g2_tiehi \top_ihp.oisc.regs[27][24]$_DFFE_PP__1817  (.L_HI(net1817));
 sg13g2_tiehi \top_ihp.oisc.regs[27][25]$_DFFE_PP__1818  (.L_HI(net1818));
 sg13g2_tiehi \top_ihp.oisc.regs[27][26]$_DFFE_PP__1819  (.L_HI(net1819));
 sg13g2_tiehi \top_ihp.oisc.regs[27][27]$_DFFE_PP__1820  (.L_HI(net1820));
 sg13g2_tiehi \top_ihp.oisc.regs[27][28]$_DFFE_PP__1821  (.L_HI(net1821));
 sg13g2_tiehi \top_ihp.oisc.regs[27][29]$_DFFE_PP__1822  (.L_HI(net1822));
 sg13g2_tiehi \top_ihp.oisc.regs[27][2]$_DFFE_PP__1823  (.L_HI(net1823));
 sg13g2_tiehi \top_ihp.oisc.regs[27][30]$_DFFE_PP__1824  (.L_HI(net1824));
 sg13g2_tiehi \top_ihp.oisc.regs[27][31]$_DFFE_PP__1825  (.L_HI(net1825));
 sg13g2_tiehi \top_ihp.oisc.regs[27][3]$_DFFE_PP__1826  (.L_HI(net1826));
 sg13g2_tiehi \top_ihp.oisc.regs[27][4]$_DFFE_PP__1827  (.L_HI(net1827));
 sg13g2_tiehi \top_ihp.oisc.regs[27][5]$_DFFE_PP__1828  (.L_HI(net1828));
 sg13g2_tiehi \top_ihp.oisc.regs[27][6]$_DFFE_PP__1829  (.L_HI(net1829));
 sg13g2_tiehi \top_ihp.oisc.regs[27][7]$_DFFE_PP__1830  (.L_HI(net1830));
 sg13g2_tiehi \top_ihp.oisc.regs[27][8]$_DFFE_PP__1831  (.L_HI(net1831));
 sg13g2_tiehi \top_ihp.oisc.regs[27][9]$_DFFE_PP__1832  (.L_HI(net1832));
 sg13g2_tiehi \top_ihp.oisc.regs[28][0]$_DFFE_PP__1833  (.L_HI(net1833));
 sg13g2_tiehi \top_ihp.oisc.regs[28][10]$_DFFE_PP__1834  (.L_HI(net1834));
 sg13g2_tiehi \top_ihp.oisc.regs[28][11]$_DFFE_PP__1835  (.L_HI(net1835));
 sg13g2_tiehi \top_ihp.oisc.regs[28][12]$_DFFE_PP__1836  (.L_HI(net1836));
 sg13g2_tiehi \top_ihp.oisc.regs[28][13]$_DFFE_PP__1837  (.L_HI(net1837));
 sg13g2_tiehi \top_ihp.oisc.regs[28][14]$_DFFE_PP__1838  (.L_HI(net1838));
 sg13g2_tiehi \top_ihp.oisc.regs[28][15]$_DFFE_PP__1839  (.L_HI(net1839));
 sg13g2_tiehi \top_ihp.oisc.regs[28][16]$_DFFE_PP__1840  (.L_HI(net1840));
 sg13g2_tiehi \top_ihp.oisc.regs[28][17]$_DFFE_PP__1841  (.L_HI(net1841));
 sg13g2_tiehi \top_ihp.oisc.regs[28][18]$_DFFE_PP__1842  (.L_HI(net1842));
 sg13g2_tiehi \top_ihp.oisc.regs[28][19]$_DFFE_PP__1843  (.L_HI(net1843));
 sg13g2_tiehi \top_ihp.oisc.regs[28][1]$_DFFE_PP__1844  (.L_HI(net1844));
 sg13g2_tiehi \top_ihp.oisc.regs[28][20]$_DFFE_PP__1845  (.L_HI(net1845));
 sg13g2_tiehi \top_ihp.oisc.regs[28][21]$_DFFE_PP__1846  (.L_HI(net1846));
 sg13g2_tiehi \top_ihp.oisc.regs[28][22]$_DFFE_PP__1847  (.L_HI(net1847));
 sg13g2_tiehi \top_ihp.oisc.regs[28][23]$_DFFE_PP__1848  (.L_HI(net1848));
 sg13g2_tiehi \top_ihp.oisc.regs[28][24]$_DFFE_PP__1849  (.L_HI(net1849));
 sg13g2_tiehi \top_ihp.oisc.regs[28][25]$_DFFE_PP__1850  (.L_HI(net1850));
 sg13g2_tiehi \top_ihp.oisc.regs[28][26]$_DFFE_PP__1851  (.L_HI(net1851));
 sg13g2_tiehi \top_ihp.oisc.regs[28][27]$_DFFE_PP__1852  (.L_HI(net1852));
 sg13g2_tiehi \top_ihp.oisc.regs[28][28]$_DFFE_PP__1853  (.L_HI(net1853));
 sg13g2_tiehi \top_ihp.oisc.regs[28][29]$_DFFE_PP__1854  (.L_HI(net1854));
 sg13g2_tiehi \top_ihp.oisc.regs[28][2]$_DFFE_PP__1855  (.L_HI(net1855));
 sg13g2_tiehi \top_ihp.oisc.regs[28][30]$_DFFE_PP__1856  (.L_HI(net1856));
 sg13g2_tiehi \top_ihp.oisc.regs[28][31]$_DFFE_PP__1857  (.L_HI(net1857));
 sg13g2_tiehi \top_ihp.oisc.regs[28][3]$_DFFE_PP__1858  (.L_HI(net1858));
 sg13g2_tiehi \top_ihp.oisc.regs[28][4]$_DFFE_PP__1859  (.L_HI(net1859));
 sg13g2_tiehi \top_ihp.oisc.regs[28][5]$_DFFE_PP__1860  (.L_HI(net1860));
 sg13g2_tiehi \top_ihp.oisc.regs[28][6]$_DFFE_PP__1861  (.L_HI(net1861));
 sg13g2_tiehi \top_ihp.oisc.regs[28][7]$_DFFE_PP__1862  (.L_HI(net1862));
 sg13g2_tiehi \top_ihp.oisc.regs[28][8]$_DFFE_PP__1863  (.L_HI(net1863));
 sg13g2_tiehi \top_ihp.oisc.regs[28][9]$_DFFE_PP__1864  (.L_HI(net1864));
 sg13g2_tiehi \top_ihp.oisc.regs[29][0]$_DFFE_PP__1865  (.L_HI(net1865));
 sg13g2_tiehi \top_ihp.oisc.regs[29][10]$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \top_ihp.oisc.regs[29][11]$_DFFE_PP__1867  (.L_HI(net1867));
 sg13g2_tiehi \top_ihp.oisc.regs[29][12]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \top_ihp.oisc.regs[29][13]$_DFFE_PP__1869  (.L_HI(net1869));
 sg13g2_tiehi \top_ihp.oisc.regs[29][14]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \top_ihp.oisc.regs[29][15]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \top_ihp.oisc.regs[29][16]$_DFFE_PP__1872  (.L_HI(net1872));
 sg13g2_tiehi \top_ihp.oisc.regs[29][17]$_DFFE_PP__1873  (.L_HI(net1873));
 sg13g2_tiehi \top_ihp.oisc.regs[29][18]$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \top_ihp.oisc.regs[29][19]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \top_ihp.oisc.regs[29][1]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \top_ihp.oisc.regs[29][20]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \top_ihp.oisc.regs[29][21]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \top_ihp.oisc.regs[29][22]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \top_ihp.oisc.regs[29][23]$_DFFE_PP__1880  (.L_HI(net1880));
 sg13g2_tiehi \top_ihp.oisc.regs[29][24]$_DFFE_PP__1881  (.L_HI(net1881));
 sg13g2_tiehi \top_ihp.oisc.regs[29][25]$_DFFE_PP__1882  (.L_HI(net1882));
 sg13g2_tiehi \top_ihp.oisc.regs[29][26]$_DFFE_PP__1883  (.L_HI(net1883));
 sg13g2_tiehi \top_ihp.oisc.regs[29][27]$_DFFE_PP__1884  (.L_HI(net1884));
 sg13g2_tiehi \top_ihp.oisc.regs[29][28]$_DFFE_PP__1885  (.L_HI(net1885));
 sg13g2_tiehi \top_ihp.oisc.regs[29][29]$_DFFE_PP__1886  (.L_HI(net1886));
 sg13g2_tiehi \top_ihp.oisc.regs[29][2]$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \top_ihp.oisc.regs[29][30]$_DFFE_PP__1888  (.L_HI(net1888));
 sg13g2_tiehi \top_ihp.oisc.regs[29][31]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \top_ihp.oisc.regs[29][3]$_DFFE_PP__1890  (.L_HI(net1890));
 sg13g2_tiehi \top_ihp.oisc.regs[29][4]$_DFFE_PP__1891  (.L_HI(net1891));
 sg13g2_tiehi \top_ihp.oisc.regs[29][5]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \top_ihp.oisc.regs[29][6]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \top_ihp.oisc.regs[29][7]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \top_ihp.oisc.regs[29][8]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \top_ihp.oisc.regs[29][9]$_DFFE_PP__1896  (.L_HI(net1896));
 sg13g2_tiehi \top_ihp.oisc.regs[30][0]$_DFFE_PP__1897  (.L_HI(net1897));
 sg13g2_tiehi \top_ihp.oisc.regs[30][10]$_DFFE_PP__1898  (.L_HI(net1898));
 sg13g2_tiehi \top_ihp.oisc.regs[30][11]$_DFFE_PP__1899  (.L_HI(net1899));
 sg13g2_tiehi \top_ihp.oisc.regs[30][12]$_DFFE_PP__1900  (.L_HI(net1900));
 sg13g2_tiehi \top_ihp.oisc.regs[30][13]$_DFFE_PP__1901  (.L_HI(net1901));
 sg13g2_tiehi \top_ihp.oisc.regs[30][14]$_DFFE_PP__1902  (.L_HI(net1902));
 sg13g2_tiehi \top_ihp.oisc.regs[30][15]$_DFFE_PP__1903  (.L_HI(net1903));
 sg13g2_tiehi \top_ihp.oisc.regs[30][16]$_DFFE_PP__1904  (.L_HI(net1904));
 sg13g2_tiehi \top_ihp.oisc.regs[30][17]$_DFFE_PP__1905  (.L_HI(net1905));
 sg13g2_tiehi \top_ihp.oisc.regs[30][18]$_DFFE_PP__1906  (.L_HI(net1906));
 sg13g2_tiehi \top_ihp.oisc.regs[30][19]$_DFFE_PP__1907  (.L_HI(net1907));
 sg13g2_tiehi \top_ihp.oisc.regs[30][1]$_DFFE_PP__1908  (.L_HI(net1908));
 sg13g2_tiehi \top_ihp.oisc.regs[30][20]$_DFFE_PP__1909  (.L_HI(net1909));
 sg13g2_tiehi \top_ihp.oisc.regs[30][21]$_DFFE_PP__1910  (.L_HI(net1910));
 sg13g2_tiehi \top_ihp.oisc.regs[30][22]$_DFFE_PP__1911  (.L_HI(net1911));
 sg13g2_tiehi \top_ihp.oisc.regs[30][23]$_DFFE_PP__1912  (.L_HI(net1912));
 sg13g2_tiehi \top_ihp.oisc.regs[30][24]$_DFFE_PP__1913  (.L_HI(net1913));
 sg13g2_tiehi \top_ihp.oisc.regs[30][25]$_DFFE_PP__1914  (.L_HI(net1914));
 sg13g2_tiehi \top_ihp.oisc.regs[30][26]$_DFFE_PP__1915  (.L_HI(net1915));
 sg13g2_tiehi \top_ihp.oisc.regs[30][27]$_DFFE_PP__1916  (.L_HI(net1916));
 sg13g2_tiehi \top_ihp.oisc.regs[30][28]$_DFFE_PP__1917  (.L_HI(net1917));
 sg13g2_tiehi \top_ihp.oisc.regs[30][29]$_DFFE_PP__1918  (.L_HI(net1918));
 sg13g2_tiehi \top_ihp.oisc.regs[30][2]$_DFFE_PP__1919  (.L_HI(net1919));
 sg13g2_tiehi \top_ihp.oisc.regs[30][30]$_DFFE_PP__1920  (.L_HI(net1920));
 sg13g2_tiehi \top_ihp.oisc.regs[30][31]$_DFFE_PP__1921  (.L_HI(net1921));
 sg13g2_tiehi \top_ihp.oisc.regs[30][3]$_DFFE_PP__1922  (.L_HI(net1922));
 sg13g2_tiehi \top_ihp.oisc.regs[30][4]$_DFFE_PP__1923  (.L_HI(net1923));
 sg13g2_tiehi \top_ihp.oisc.regs[30][5]$_DFFE_PP__1924  (.L_HI(net1924));
 sg13g2_tiehi \top_ihp.oisc.regs[30][6]$_DFFE_PP__1925  (.L_HI(net1925));
 sg13g2_tiehi \top_ihp.oisc.regs[30][7]$_DFFE_PP__1926  (.L_HI(net1926));
 sg13g2_tiehi \top_ihp.oisc.regs[30][8]$_DFFE_PP__1927  (.L_HI(net1927));
 sg13g2_tiehi \top_ihp.oisc.regs[30][9]$_DFFE_PP__1928  (.L_HI(net1928));
 sg13g2_tiehi \top_ihp.oisc.regs[31][0]$_DFFE_PP__1929  (.L_HI(net1929));
 sg13g2_tiehi \top_ihp.oisc.regs[31][10]$_DFFE_PP__1930  (.L_HI(net1930));
 sg13g2_tiehi \top_ihp.oisc.regs[31][11]$_DFFE_PP__1931  (.L_HI(net1931));
 sg13g2_tiehi \top_ihp.oisc.regs[31][12]$_DFFE_PP__1932  (.L_HI(net1932));
 sg13g2_tiehi \top_ihp.oisc.regs[31][13]$_DFFE_PP__1933  (.L_HI(net1933));
 sg13g2_tiehi \top_ihp.oisc.regs[31][14]$_DFFE_PP__1934  (.L_HI(net1934));
 sg13g2_tiehi \top_ihp.oisc.regs[31][15]$_DFFE_PP__1935  (.L_HI(net1935));
 sg13g2_tiehi \top_ihp.oisc.regs[31][16]$_DFFE_PP__1936  (.L_HI(net1936));
 sg13g2_tiehi \top_ihp.oisc.regs[31][17]$_DFFE_PP__1937  (.L_HI(net1937));
 sg13g2_tiehi \top_ihp.oisc.regs[31][18]$_DFFE_PP__1938  (.L_HI(net1938));
 sg13g2_tiehi \top_ihp.oisc.regs[31][19]$_DFFE_PP__1939  (.L_HI(net1939));
 sg13g2_tiehi \top_ihp.oisc.regs[31][1]$_DFFE_PP__1940  (.L_HI(net1940));
 sg13g2_tiehi \top_ihp.oisc.regs[31][20]$_DFFE_PP__1941  (.L_HI(net1941));
 sg13g2_tiehi \top_ihp.oisc.regs[31][21]$_DFFE_PP__1942  (.L_HI(net1942));
 sg13g2_tiehi \top_ihp.oisc.regs[31][22]$_DFFE_PP__1943  (.L_HI(net1943));
 sg13g2_tiehi \top_ihp.oisc.regs[31][23]$_DFFE_PP__1944  (.L_HI(net1944));
 sg13g2_tiehi \top_ihp.oisc.regs[31][24]$_DFFE_PP__1945  (.L_HI(net1945));
 sg13g2_tiehi \top_ihp.oisc.regs[31][25]$_DFFE_PP__1946  (.L_HI(net1946));
 sg13g2_tiehi \top_ihp.oisc.regs[31][26]$_DFFE_PP__1947  (.L_HI(net1947));
 sg13g2_tiehi \top_ihp.oisc.regs[31][27]$_DFFE_PP__1948  (.L_HI(net1948));
 sg13g2_tiehi \top_ihp.oisc.regs[31][28]$_DFFE_PP__1949  (.L_HI(net1949));
 sg13g2_tiehi \top_ihp.oisc.regs[31][29]$_DFFE_PP__1950  (.L_HI(net1950));
 sg13g2_tiehi \top_ihp.oisc.regs[31][2]$_DFFE_PP__1951  (.L_HI(net1951));
 sg13g2_tiehi \top_ihp.oisc.regs[31][30]$_DFFE_PP__1952  (.L_HI(net1952));
 sg13g2_tiehi \top_ihp.oisc.regs[31][31]$_DFFE_PP__1953  (.L_HI(net1953));
 sg13g2_tiehi \top_ihp.oisc.regs[31][3]$_DFFE_PP__1954  (.L_HI(net1954));
 sg13g2_tiehi \top_ihp.oisc.regs[31][4]$_DFFE_PP__1955  (.L_HI(net1955));
 sg13g2_tiehi \top_ihp.oisc.regs[31][5]$_DFFE_PP__1956  (.L_HI(net1956));
 sg13g2_tiehi \top_ihp.oisc.regs[31][6]$_DFFE_PP__1957  (.L_HI(net1957));
 sg13g2_tiehi \top_ihp.oisc.regs[31][7]$_DFFE_PP__1958  (.L_HI(net1958));
 sg13g2_tiehi \top_ihp.oisc.regs[31][8]$_DFFE_PP__1959  (.L_HI(net1959));
 sg13g2_tiehi \top_ihp.oisc.regs[31][9]$_DFFE_PP__1960  (.L_HI(net1960));
 sg13g2_tiehi \top_ihp.oisc.regs[32][0]$_DFFE_PP__1961  (.L_HI(net1961));
 sg13g2_tiehi \top_ihp.oisc.regs[32][10]$_DFFE_PP__1962  (.L_HI(net1962));
 sg13g2_tiehi \top_ihp.oisc.regs[32][11]$_DFFE_PP__1963  (.L_HI(net1963));
 sg13g2_tiehi \top_ihp.oisc.regs[32][12]$_DFFE_PP__1964  (.L_HI(net1964));
 sg13g2_tiehi \top_ihp.oisc.regs[32][13]$_DFFE_PP__1965  (.L_HI(net1965));
 sg13g2_tiehi \top_ihp.oisc.regs[32][14]$_DFFE_PP__1966  (.L_HI(net1966));
 sg13g2_tiehi \top_ihp.oisc.regs[32][15]$_DFFE_PP__1967  (.L_HI(net1967));
 sg13g2_tiehi \top_ihp.oisc.regs[32][16]$_DFFE_PP__1968  (.L_HI(net1968));
 sg13g2_tiehi \top_ihp.oisc.regs[32][17]$_DFFE_PP__1969  (.L_HI(net1969));
 sg13g2_tiehi \top_ihp.oisc.regs[32][18]$_DFFE_PP__1970  (.L_HI(net1970));
 sg13g2_tiehi \top_ihp.oisc.regs[32][19]$_DFFE_PP__1971  (.L_HI(net1971));
 sg13g2_tiehi \top_ihp.oisc.regs[32][1]$_DFFE_PP__1972  (.L_HI(net1972));
 sg13g2_tiehi \top_ihp.oisc.regs[32][20]$_DFFE_PP__1973  (.L_HI(net1973));
 sg13g2_tiehi \top_ihp.oisc.regs[32][21]$_DFFE_PP__1974  (.L_HI(net1974));
 sg13g2_tiehi \top_ihp.oisc.regs[32][22]$_DFFE_PP__1975  (.L_HI(net1975));
 sg13g2_tiehi \top_ihp.oisc.regs[32][23]$_DFFE_PP__1976  (.L_HI(net1976));
 sg13g2_tiehi \top_ihp.oisc.regs[32][24]$_DFFE_PP__1977  (.L_HI(net1977));
 sg13g2_tiehi \top_ihp.oisc.regs[32][25]$_DFFE_PP__1978  (.L_HI(net1978));
 sg13g2_tiehi \top_ihp.oisc.regs[32][26]$_DFFE_PP__1979  (.L_HI(net1979));
 sg13g2_tiehi \top_ihp.oisc.regs[32][27]$_DFFE_PP__1980  (.L_HI(net1980));
 sg13g2_tiehi \top_ihp.oisc.regs[32][28]$_DFFE_PP__1981  (.L_HI(net1981));
 sg13g2_tiehi \top_ihp.oisc.regs[32][29]$_DFFE_PP__1982  (.L_HI(net1982));
 sg13g2_tiehi \top_ihp.oisc.regs[32][2]$_DFFE_PP__1983  (.L_HI(net1983));
 sg13g2_tiehi \top_ihp.oisc.regs[32][30]$_DFFE_PP__1984  (.L_HI(net1984));
 sg13g2_tiehi \top_ihp.oisc.regs[32][31]$_DFFE_PP__1985  (.L_HI(net1985));
 sg13g2_tiehi \top_ihp.oisc.regs[32][3]$_DFFE_PP__1986  (.L_HI(net1986));
 sg13g2_tiehi \top_ihp.oisc.regs[32][4]$_DFFE_PP__1987  (.L_HI(net1987));
 sg13g2_tiehi \top_ihp.oisc.regs[32][5]$_DFFE_PP__1988  (.L_HI(net1988));
 sg13g2_tiehi \top_ihp.oisc.regs[32][6]$_DFFE_PP__1989  (.L_HI(net1989));
 sg13g2_tiehi \top_ihp.oisc.regs[32][7]$_DFFE_PP__1990  (.L_HI(net1990));
 sg13g2_tiehi \top_ihp.oisc.regs[32][8]$_DFFE_PP__1991  (.L_HI(net1991));
 sg13g2_tiehi \top_ihp.oisc.regs[32][9]$_DFFE_PP__1992  (.L_HI(net1992));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[0]$_SDFFCE_PN0P__1993  (.L_HI(net1993));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[1]$_SDFFCE_PN0P__1994  (.L_HI(net1994));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[2]$_SDFFCE_PN0P__1995  (.L_HI(net1995));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[3]$_SDFFCE_PN0P__1996  (.L_HI(net1996));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[4]$_SDFFCE_PN0P__1997  (.L_HI(net1997));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[5]$_SDFFCE_PN0P__1998  (.L_HI(net1998));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[6]$_SDFFCE_PN0P__1999  (.L_HI(net1999));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[7]$_SDFFCE_PN0P__2000  (.L_HI(net2000));
 sg13g2_tiehi \top_ihp.wb_emem.last_bit$_DFFE_PP__2001  (.L_HI(net2001));
 sg13g2_tiehi \top_ihp.wb_emem.last_wait$_DFFE_PP__2002  (.L_HI(net2002));
 sg13g2_tiehi \top_ihp.wb_emem.nbits[3]$_SDFFCE_NP1P__2003  (.L_HI(net2003));
 sg13g2_tiehi \top_ihp.wb_emem.nbits[4]$_SDFFCE_NP0P__2004  (.L_HI(net2004));
 sg13g2_tiehi \top_ihp.wb_emem.nbits[5]$_SDFFCE_NP0P__2005  (.L_HI(net2005));
 sg13g2_tiehi \top_ihp.wb_emem.nbits[6]$_SDFFCE_NP0P__2006  (.L_HI(net2006));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[0]$_SDFFCE_PN0P__2007  (.L_HI(net2007));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[1]$_SDFFCE_PN0P__2008  (.L_HI(net2008));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[2]$_SDFFCE_PN0P__2009  (.L_HI(net2009));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[3]$_SDFFCE_PN0P__2010  (.L_HI(net2010));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[4]$_SDFFCE_PN0P__2011  (.L_HI(net2011));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[5]$_SDFFCE_PN0P__2012  (.L_HI(net2012));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[6]$_SDFFCE_PN0P__2013  (.L_HI(net2013));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[7]$_SDFFCE_PN0P__2014  (.L_HI(net2014));
 sg13g2_tiehi \top_ihp.wb_uart.ack_o$_SDFFCE_PP0P__2015  (.L_HI(net2015));
 sg13g2_inv_1 net1791_2 (.Y(net2017),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 net1791_3 (.Y(net2018),
    .A(clknet_leaf_64_clk));
 sg13g2_inv_1 net1791_4 (.Y(net2019),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 net1791_5 (.Y(net2020),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 net1791_6 (.Y(net2021),
    .A(clknet_leaf_61_clk));
 sg13g2_inv_1 net1791_7 (.Y(net2022),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 net1791_8 (.Y(net2023),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 net1791_9 (.Y(net2024),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 net1791_10 (.Y(net2025),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 net1791_11 (.Y(net2026),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 net1791_12 (.Y(net2027),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 net1791_13 (.Y(net2028),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 net1791_14 (.Y(net2029),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 net1791_15 (.Y(net2030),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 net1791_16 (.Y(net2031),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _17 (.Y(net2032),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _17_18 (.Y(net2033),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _17_19 (.Y(net2034),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _17_20 (.Y(net2035),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _17_21 (.Y(net2036),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _17_22 (.Y(net2037),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _17_23 (.Y(net2038),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _17_24 (.Y(net2039),
    .A(clknet_leaf_55_clk));
 sg13g2_inv_1 _17_25 (.Y(net2040),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _17_26 (.Y(net2041),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _17_27 (.Y(net2042),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _17_28 (.Y(net2043),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _17_29 (.Y(net2044),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _17_30 (.Y(net2045),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _17_31 (.Y(net2046),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _17_32 (.Y(net2047),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _17_33 (.Y(net2048),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _17_34 (.Y(net2049),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _17_35 (.Y(net2050),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _17_36 (.Y(net2051),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _17_37 (.Y(net2052),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _17_38 (.Y(net2053),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _17_39 (.Y(net2054),
    .A(clknet_leaf_61_clk));
 sg13g2_inv_1 _17_40 (.Y(net2055),
    .A(clknet_leaf_61_clk));
 sg13g2_inv_1 _17_41 (.Y(net2056),
    .A(clknet_leaf_62_clk));
 sg13g2_inv_1 _17_42 (.Y(net2057),
    .A(clknet_leaf_61_clk));
 sg13g2_inv_1 _17_43 (.Y(net2058),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 _17_44 (.Y(net2059),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 _17_45 (.Y(net2060),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _17_46 (.Y(net2061),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _17_47 (.Y(net2062),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _17_48 (.Y(net2063),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _17_49 (.Y(net2064),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 _17_50 (.Y(net2065),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _17_51 (.Y(net2066),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 _17_52 (.Y(net2067),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 _17_53 (.Y(net2068),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 _17_54 (.Y(net2069),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 _17_55 (.Y(net2070),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 _17_56 (.Y(net2071),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 _17_57 (.Y(net2072),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _17_58 (.Y(net2073),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _17_59 (.Y(net2074),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _17_60 (.Y(net2075),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 _17_61 (.Y(net2076),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 _17_62 (.Y(net2077),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _17_63 (.Y(net2078),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _17_64 (.Y(net2079),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _17_65 (.Y(net2080),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _17_66 (.Y(net2081),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _17_67 (.Y(net2082),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _17_68 (.Y(net2083),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _17_69 (.Y(net2084),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _17_70 (.Y(net2085),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _17_71 (.Y(net2086),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _17_72 (.Y(net2087),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 _17_73 (.Y(net2088),
    .A(clknet_leaf_20_clk));
 sg13g2_inv_1 _17_74 (.Y(net2089),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _17_75 (.Y(net2090),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _17_76 (.Y(net2091),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _17_77 (.Y(net2092),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _17_78 (.Y(net2093),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _17_79 (.Y(net2094),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _17_80 (.Y(net2095),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _17_81 (.Y(net2096),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _17_82 (.Y(net2097),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _17_83 (.Y(net2098),
    .A(clknet_leaf_20_clk));
 sg13g2_inv_1 _17_84 (.Y(net2099),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _17_85 (.Y(net2100),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _17_86 (.Y(net2101),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _17_87 (.Y(net2102),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _17_88 (.Y(net2103),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _17_89 (.Y(net2104),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _17_90 (.Y(net2105),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _17_91 (.Y(net2106),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _17_92 (.Y(net2107),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 _17_93 (.Y(net2108),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 _17_94 (.Y(net2109),
    .A(clknet_leaf_20_clk));
 sg13g2_inv_1 _17_95 (.Y(net2110),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 _17_96 (.Y(net2111),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _17_97 (.Y(net2112),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _17_98 (.Y(net2113),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _17_99 (.Y(net2114),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 _17_100 (.Y(net2115),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _17_101 (.Y(net2116),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 _17_102 (.Y(net2117),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _17_103 (.Y(net2118),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _17_104 (.Y(net2119),
    .A(clknet_leaf_20_clk));
 sg13g2_inv_1 _17_105 (.Y(net2120),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _17_106 (.Y(net2121),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _17_107 (.Y(net2122),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _17_108 (.Y(net2123),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _17_109 (.Y(net2124),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _17_110 (.Y(net2125),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _17_111 (.Y(net2126),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _17_112 (.Y(net2127),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _17_113 (.Y(net2128),
    .A(clknet_leaf_20_clk));
 sg13g2_inv_1 _17_114 (.Y(net2129),
    .A(clknet_leaf_20_clk));
 sg13g2_inv_1 _17_115 (.Y(net2130),
    .A(clknet_leaf_20_clk));
 sg13g2_inv_1 _17_116 (.Y(net2131),
    .A(clknet_leaf_20_clk));
 sg13g2_inv_1 _17_117 (.Y(net2132),
    .A(clknet_leaf_59_clk));
 sg13g2_inv_1 _17_118 (.Y(net2133),
    .A(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_8 clkbuf_leaf_311_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_8 clkbuf_leaf_312_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_8 clkbuf_leaf_313_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_313_clk));
 sg13g2_buf_8 clkbuf_leaf_314_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_314_clk));
 sg13g2_buf_8 clkbuf_leaf_315_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_315_clk));
 sg13g2_buf_8 clkbuf_leaf_316_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_316_clk));
 sg13g2_buf_8 clkbuf_leaf_317_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_317_clk));
 sg13g2_buf_8 clkbuf_leaf_318_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_318_clk));
 sg13g2_buf_8 clkbuf_leaf_319_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_319_clk));
 sg13g2_buf_8 clkbuf_leaf_320_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_320_clk));
 sg13g2_buf_8 clkbuf_leaf_321_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_321_clk));
 sg13g2_buf_8 clkbuf_leaf_322_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_322_clk));
 sg13g2_buf_8 clkbuf_leaf_323_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_323_clk));
 sg13g2_buf_8 clkbuf_leaf_324_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_324_clk));
 sg13g2_buf_8 clkbuf_leaf_325_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_325_clk));
 sg13g2_buf_8 clkbuf_leaf_326_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_326_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_0__f_clk (.X(clknet_6_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_1__f_clk (.X(clknet_6_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_2__f_clk (.X(clknet_6_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_3__f_clk (.X(clknet_6_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_4__f_clk (.X(clknet_6_4__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_5__f_clk (.X(clknet_6_5__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_6__f_clk (.X(clknet_6_6__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_7__f_clk (.X(clknet_6_7__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_8__f_clk (.X(clknet_6_8__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_9__f_clk (.X(clknet_6_9__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_10__f_clk (.X(clknet_6_10__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_11__f_clk (.X(clknet_6_11__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_12__f_clk (.X(clknet_6_12__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_13__f_clk (.X(clknet_6_13__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_14__f_clk (.X(clknet_6_14__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_15__f_clk (.X(clknet_6_15__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_16__f_clk (.X(clknet_6_16__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_17__f_clk (.X(clknet_6_17__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_18__f_clk (.X(clknet_6_18__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_19__f_clk (.X(clknet_6_19__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_20__f_clk (.X(clknet_6_20__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_21__f_clk (.X(clknet_6_21__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_22__f_clk (.X(clknet_6_22__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_23__f_clk (.X(clknet_6_23__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_24__f_clk (.X(clknet_6_24__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_25__f_clk (.X(clknet_6_25__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_26__f_clk (.X(clknet_6_26__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_27__f_clk (.X(clknet_6_27__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_28__f_clk (.X(clknet_6_28__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_29__f_clk (.X(clknet_6_29__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_30__f_clk (.X(clknet_6_30__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_31__f_clk (.X(clknet_6_31__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_32__f_clk (.X(clknet_6_32__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_33__f_clk (.X(clknet_6_33__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_34__f_clk (.X(clknet_6_34__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_35__f_clk (.X(clknet_6_35__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_36__f_clk (.X(clknet_6_36__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_37__f_clk (.X(clknet_6_37__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_38__f_clk (.X(clknet_6_38__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_39__f_clk (.X(clknet_6_39__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_40__f_clk (.X(clknet_6_40__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_41__f_clk (.X(clknet_6_41__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_42__f_clk (.X(clknet_6_42__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_43__f_clk (.X(clknet_6_43__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_44__f_clk (.X(clknet_6_44__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_45__f_clk (.X(clknet_6_45__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_46__f_clk (.X(clknet_6_46__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_47__f_clk (.X(clknet_6_47__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_48__f_clk (.X(clknet_6_48__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_49__f_clk (.X(clknet_6_49__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_50__f_clk (.X(clknet_6_50__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_51__f_clk (.X(clknet_6_51__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_52__f_clk (.X(clknet_6_52__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_53__f_clk (.X(clknet_6_53__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_54__f_clk (.X(clknet_6_54__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_55__f_clk (.X(clknet_6_55__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_56__f_clk (.X(clknet_6_56__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_57__f_clk (.X(clknet_6_57__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_58__f_clk (.X(clknet_6_58__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_59__f_clk (.X(clknet_6_59__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_60__f_clk (.X(clknet_6_60__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_61__f_clk (.X(clknet_6_61__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_62__f_clk (.X(clknet_6_62__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_63__f_clk (.X(clknet_6_63__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_1__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_2__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_3__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_4__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_5__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_6__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_6_9__leaf_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_6_10__leaf_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_6_11__leaf_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_6_12__leaf_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_6_13__leaf_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_6_14__leaf_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload14 (.A(clknet_6_17__leaf_clk));
 sg13g2_buf_8 clkload15 (.A(clknet_6_18__leaf_clk));
 sg13g2_buf_8 clkload16 (.A(clknet_6_19__leaf_clk));
 sg13g2_buf_8 clkload17 (.A(clknet_6_20__leaf_clk));
 sg13g2_buf_8 clkload18 (.A(clknet_6_21__leaf_clk));
 sg13g2_buf_8 clkload19 (.A(clknet_6_22__leaf_clk));
 sg13g2_buf_8 clkload20 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload21 (.A(clknet_6_25__leaf_clk));
 sg13g2_buf_8 clkload22 (.A(clknet_6_26__leaf_clk));
 sg13g2_buf_8 clkload23 (.A(clknet_6_27__leaf_clk));
 sg13g2_buf_8 clkload24 (.A(clknet_6_28__leaf_clk));
 sg13g2_buf_8 clkload25 (.A(clknet_6_29__leaf_clk));
 sg13g2_buf_8 clkload26 (.A(clknet_6_30__leaf_clk));
 sg13g2_buf_8 clkload27 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload28 (.A(clknet_6_33__leaf_clk));
 sg13g2_buf_8 clkload29 (.A(clknet_6_34__leaf_clk));
 sg13g2_buf_8 clkload30 (.A(clknet_6_35__leaf_clk));
 sg13g2_buf_8 clkload31 (.A(clknet_6_36__leaf_clk));
 sg13g2_buf_8 clkload32 (.A(clknet_6_37__leaf_clk));
 sg13g2_buf_8 clkload33 (.A(clknet_6_38__leaf_clk));
 sg13g2_buf_8 clkload34 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload35 (.A(clknet_6_41__leaf_clk));
 sg13g2_buf_8 clkload36 (.A(clknet_6_42__leaf_clk));
 sg13g2_buf_8 clkload37 (.A(clknet_6_43__leaf_clk));
 sg13g2_buf_8 clkload38 (.A(clknet_6_44__leaf_clk));
 sg13g2_buf_8 clkload39 (.A(clknet_6_45__leaf_clk));
 sg13g2_buf_8 clkload40 (.A(clknet_6_46__leaf_clk));
 sg13g2_buf_8 clkload41 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload42 (.A(clknet_6_49__leaf_clk));
 sg13g2_buf_8 clkload43 (.A(clknet_6_50__leaf_clk));
 sg13g2_buf_8 clkload44 (.A(clknet_6_51__leaf_clk));
 sg13g2_buf_8 clkload45 (.A(clknet_6_52__leaf_clk));
 sg13g2_buf_8 clkload46 (.A(clknet_6_53__leaf_clk));
 sg13g2_buf_8 clkload47 (.A(clknet_6_54__leaf_clk));
 sg13g2_buf_8 clkload48 (.A(clknet_6_55__leaf_clk));
 sg13g2_inv_1 clkload49 (.A(clknet_leaf_326_clk));
 sg13g2_inv_2 clkload50 (.A(clknet_leaf_39_clk));
 sg13g2_buf_16 clkload51 (.A(clknet_leaf_58_clk));
 sg13g2_inv_2 clkload52 (.A(clknet_leaf_38_clk));
 sg13g2_inv_4 clkload53 (.A(clknet_leaf_40_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00366_));
 sg13g2_antennanp ANTENNA_2 (.A(_00394_));
 sg13g2_antennanp ANTENNA_3 (.A(_00406_));
 sg13g2_antennanp ANTENNA_4 (.A(_00406_));
 sg13g2_antennanp ANTENNA_5 (.A(_00408_));
 sg13g2_antennanp ANTENNA_6 (.A(_00411_));
 sg13g2_antennanp ANTENNA_7 (.A(_00412_));
 sg13g2_antennanp ANTENNA_8 (.A(_00413_));
 sg13g2_antennanp ANTENNA_9 (.A(_00413_));
 sg13g2_antennanp ANTENNA_10 (.A(_00417_));
 sg13g2_antennanp ANTENNA_11 (.A(_03004_));
 sg13g2_antennanp ANTENNA_12 (.A(_03004_));
 sg13g2_antennanp ANTENNA_13 (.A(_03004_));
 sg13g2_antennanp ANTENNA_14 (.A(_03056_));
 sg13g2_antennanp ANTENNA_15 (.A(_03056_));
 sg13g2_antennanp ANTENNA_16 (.A(_03056_));
 sg13g2_antennanp ANTENNA_17 (.A(_03063_));
 sg13g2_antennanp ANTENNA_18 (.A(_03063_));
 sg13g2_antennanp ANTENNA_19 (.A(_03063_));
 sg13g2_antennanp ANTENNA_20 (.A(_03063_));
 sg13g2_antennanp ANTENNA_21 (.A(_03145_));
 sg13g2_antennanp ANTENNA_22 (.A(_03441_));
 sg13g2_antennanp ANTENNA_23 (.A(_03441_));
 sg13g2_antennanp ANTENNA_24 (.A(_03441_));
 sg13g2_antennanp ANTENNA_25 (.A(_03441_));
 sg13g2_antennanp ANTENNA_26 (.A(_03441_));
 sg13g2_antennanp ANTENNA_27 (.A(_03441_));
 sg13g2_antennanp ANTENNA_28 (.A(_03441_));
 sg13g2_antennanp ANTENNA_29 (.A(_03441_));
 sg13g2_antennanp ANTENNA_30 (.A(_03441_));
 sg13g2_antennanp ANTENNA_31 (.A(_03441_));
 sg13g2_antennanp ANTENNA_32 (.A(_03446_));
 sg13g2_antennanp ANTENNA_33 (.A(_03446_));
 sg13g2_antennanp ANTENNA_34 (.A(_03446_));
 sg13g2_antennanp ANTENNA_35 (.A(_03451_));
 sg13g2_antennanp ANTENNA_36 (.A(_03451_));
 sg13g2_antennanp ANTENNA_37 (.A(_03451_));
 sg13g2_antennanp ANTENNA_38 (.A(_03451_));
 sg13g2_antennanp ANTENNA_39 (.A(_03451_));
 sg13g2_antennanp ANTENNA_40 (.A(_03464_));
 sg13g2_antennanp ANTENNA_41 (.A(_03464_));
 sg13g2_antennanp ANTENNA_42 (.A(_03464_));
 sg13g2_antennanp ANTENNA_43 (.A(_03464_));
 sg13g2_antennanp ANTENNA_44 (.A(_03464_));
 sg13g2_antennanp ANTENNA_45 (.A(_03464_));
 sg13g2_antennanp ANTENNA_46 (.A(_03464_));
 sg13g2_antennanp ANTENNA_47 (.A(_03464_));
 sg13g2_antennanp ANTENNA_48 (.A(_03464_));
 sg13g2_antennanp ANTENNA_49 (.A(_03464_));
 sg13g2_antennanp ANTENNA_50 (.A(_03534_));
 sg13g2_antennanp ANTENNA_51 (.A(_03534_));
 sg13g2_antennanp ANTENNA_52 (.A(_03534_));
 sg13g2_antennanp ANTENNA_53 (.A(_03534_));
 sg13g2_antennanp ANTENNA_54 (.A(_03534_));
 sg13g2_antennanp ANTENNA_55 (.A(_03534_));
 sg13g2_antennanp ANTENNA_56 (.A(_03537_));
 sg13g2_antennanp ANTENNA_57 (.A(_03537_));
 sg13g2_antennanp ANTENNA_58 (.A(_03537_));
 sg13g2_antennanp ANTENNA_59 (.A(_03537_));
 sg13g2_antennanp ANTENNA_60 (.A(_03543_));
 sg13g2_antennanp ANTENNA_61 (.A(_03543_));
 sg13g2_antennanp ANTENNA_62 (.A(_03543_));
 sg13g2_antennanp ANTENNA_63 (.A(_03543_));
 sg13g2_antennanp ANTENNA_64 (.A(_04085_));
 sg13g2_antennanp ANTENNA_65 (.A(_04085_));
 sg13g2_antennanp ANTENNA_66 (.A(_04085_));
 sg13g2_antennanp ANTENNA_67 (.A(_04086_));
 sg13g2_antennanp ANTENNA_68 (.A(_04086_));
 sg13g2_antennanp ANTENNA_69 (.A(_04086_));
 sg13g2_antennanp ANTENNA_70 (.A(_04088_));
 sg13g2_antennanp ANTENNA_71 (.A(_04088_));
 sg13g2_antennanp ANTENNA_72 (.A(_04088_));
 sg13g2_antennanp ANTENNA_73 (.A(_04088_));
 sg13g2_antennanp ANTENNA_74 (.A(_04107_));
 sg13g2_antennanp ANTENNA_75 (.A(_04743_));
 sg13g2_antennanp ANTENNA_76 (.A(_04743_));
 sg13g2_antennanp ANTENNA_77 (.A(_05388_));
 sg13g2_antennanp ANTENNA_78 (.A(_05388_));
 sg13g2_antennanp ANTENNA_79 (.A(_05388_));
 sg13g2_antennanp ANTENNA_80 (.A(_05412_));
 sg13g2_antennanp ANTENNA_81 (.A(_05412_));
 sg13g2_antennanp ANTENNA_82 (.A(_05412_));
 sg13g2_antennanp ANTENNA_83 (.A(_05412_));
 sg13g2_antennanp ANTENNA_84 (.A(_05412_));
 sg13g2_antennanp ANTENNA_85 (.A(_05412_));
 sg13g2_antennanp ANTENNA_86 (.A(_05430_));
 sg13g2_antennanp ANTENNA_87 (.A(_05430_));
 sg13g2_antennanp ANTENNA_88 (.A(_05430_));
 sg13g2_antennanp ANTENNA_89 (.A(_05430_));
 sg13g2_antennanp ANTENNA_90 (.A(_05430_));
 sg13g2_antennanp ANTENNA_91 (.A(_05430_));
 sg13g2_antennanp ANTENNA_92 (.A(_05430_));
 sg13g2_antennanp ANTENNA_93 (.A(_05430_));
 sg13g2_antennanp ANTENNA_94 (.A(_05430_));
 sg13g2_antennanp ANTENNA_95 (.A(_05430_));
 sg13g2_antennanp ANTENNA_96 (.A(_05436_));
 sg13g2_antennanp ANTENNA_97 (.A(_05436_));
 sg13g2_antennanp ANTENNA_98 (.A(_05436_));
 sg13g2_antennanp ANTENNA_99 (.A(_05436_));
 sg13g2_antennanp ANTENNA_100 (.A(_05458_));
 sg13g2_antennanp ANTENNA_101 (.A(_05458_));
 sg13g2_antennanp ANTENNA_102 (.A(_05458_));
 sg13g2_antennanp ANTENNA_103 (.A(_05458_));
 sg13g2_antennanp ANTENNA_104 (.A(_05458_));
 sg13g2_antennanp ANTENNA_105 (.A(_05458_));
 sg13g2_antennanp ANTENNA_106 (.A(_05458_));
 sg13g2_antennanp ANTENNA_107 (.A(_05458_));
 sg13g2_antennanp ANTENNA_108 (.A(_05458_));
 sg13g2_antennanp ANTENNA_109 (.A(_05458_));
 sg13g2_antennanp ANTENNA_110 (.A(_05469_));
 sg13g2_antennanp ANTENNA_111 (.A(_05469_));
 sg13g2_antennanp ANTENNA_112 (.A(_05469_));
 sg13g2_antennanp ANTENNA_113 (.A(_05469_));
 sg13g2_antennanp ANTENNA_114 (.A(_05469_));
 sg13g2_antennanp ANTENNA_115 (.A(_05495_));
 sg13g2_antennanp ANTENNA_116 (.A(_05495_));
 sg13g2_antennanp ANTENNA_117 (.A(_05495_));
 sg13g2_antennanp ANTENNA_118 (.A(_05518_));
 sg13g2_antennanp ANTENNA_119 (.A(_05518_));
 sg13g2_antennanp ANTENNA_120 (.A(_05518_));
 sg13g2_antennanp ANTENNA_121 (.A(_05518_));
 sg13g2_antennanp ANTENNA_122 (.A(_05518_));
 sg13g2_antennanp ANTENNA_123 (.A(_05518_));
 sg13g2_antennanp ANTENNA_124 (.A(_05518_));
 sg13g2_antennanp ANTENNA_125 (.A(_05518_));
 sg13g2_antennanp ANTENNA_126 (.A(_05518_));
 sg13g2_antennanp ANTENNA_127 (.A(_05518_));
 sg13g2_antennanp ANTENNA_128 (.A(_05531_));
 sg13g2_antennanp ANTENNA_129 (.A(_05531_));
 sg13g2_antennanp ANTENNA_130 (.A(_05531_));
 sg13g2_antennanp ANTENNA_131 (.A(_05531_));
 sg13g2_antennanp ANTENNA_132 (.A(_05531_));
 sg13g2_antennanp ANTENNA_133 (.A(_05531_));
 sg13g2_antennanp ANTENNA_134 (.A(_05531_));
 sg13g2_antennanp ANTENNA_135 (.A(_05531_));
 sg13g2_antennanp ANTENNA_136 (.A(_05582_));
 sg13g2_antennanp ANTENNA_137 (.A(_05582_));
 sg13g2_antennanp ANTENNA_138 (.A(_05582_));
 sg13g2_antennanp ANTENNA_139 (.A(_05582_));
 sg13g2_antennanp ANTENNA_140 (.A(_05582_));
 sg13g2_antennanp ANTENNA_141 (.A(_05582_));
 sg13g2_antennanp ANTENNA_142 (.A(_05582_));
 sg13g2_antennanp ANTENNA_143 (.A(_05582_));
 sg13g2_antennanp ANTENNA_144 (.A(_05582_));
 sg13g2_antennanp ANTENNA_145 (.A(_05582_));
 sg13g2_antennanp ANTENNA_146 (.A(_05582_));
 sg13g2_antennanp ANTENNA_147 (.A(_05582_));
 sg13g2_antennanp ANTENNA_148 (.A(_05592_));
 sg13g2_antennanp ANTENNA_149 (.A(_05621_));
 sg13g2_antennanp ANTENNA_150 (.A(_05631_));
 sg13g2_antennanp ANTENNA_151 (.A(_05639_));
 sg13g2_antennanp ANTENNA_152 (.A(_05645_));
 sg13g2_antennanp ANTENNA_153 (.A(_05645_));
 sg13g2_antennanp ANTENNA_154 (.A(_05645_));
 sg13g2_antennanp ANTENNA_155 (.A(_05645_));
 sg13g2_antennanp ANTENNA_156 (.A(_05684_));
 sg13g2_antennanp ANTENNA_157 (.A(_05684_));
 sg13g2_antennanp ANTENNA_158 (.A(_05684_));
 sg13g2_antennanp ANTENNA_159 (.A(_05684_));
 sg13g2_antennanp ANTENNA_160 (.A(_05689_));
 sg13g2_antennanp ANTENNA_161 (.A(_05719_));
 sg13g2_antennanp ANTENNA_162 (.A(_05719_));
 sg13g2_antennanp ANTENNA_163 (.A(_05719_));
 sg13g2_antennanp ANTENNA_164 (.A(_05719_));
 sg13g2_antennanp ANTENNA_165 (.A(_05719_));
 sg13g2_antennanp ANTENNA_166 (.A(_05729_));
 sg13g2_antennanp ANTENNA_167 (.A(_05729_));
 sg13g2_antennanp ANTENNA_168 (.A(_05729_));
 sg13g2_antennanp ANTENNA_169 (.A(_05735_));
 sg13g2_antennanp ANTENNA_170 (.A(_05735_));
 sg13g2_antennanp ANTENNA_171 (.A(_05735_));
 sg13g2_antennanp ANTENNA_172 (.A(_05735_));
 sg13g2_antennanp ANTENNA_173 (.A(_05735_));
 sg13g2_antennanp ANTENNA_174 (.A(_05735_));
 sg13g2_antennanp ANTENNA_175 (.A(_05735_));
 sg13g2_antennanp ANTENNA_176 (.A(_05735_));
 sg13g2_antennanp ANTENNA_177 (.A(_05735_));
 sg13g2_antennanp ANTENNA_178 (.A(_05735_));
 sg13g2_antennanp ANTENNA_179 (.A(_05735_));
 sg13g2_antennanp ANTENNA_180 (.A(_05735_));
 sg13g2_antennanp ANTENNA_181 (.A(_05735_));
 sg13g2_antennanp ANTENNA_182 (.A(_05735_));
 sg13g2_antennanp ANTENNA_183 (.A(_05739_));
 sg13g2_antennanp ANTENNA_184 (.A(_05773_));
 sg13g2_antennanp ANTENNA_185 (.A(_05781_));
 sg13g2_antennanp ANTENNA_186 (.A(_05782_));
 sg13g2_antennanp ANTENNA_187 (.A(_05782_));
 sg13g2_antennanp ANTENNA_188 (.A(_05782_));
 sg13g2_antennanp ANTENNA_189 (.A(_05785_));
 sg13g2_antennanp ANTENNA_190 (.A(_05807_));
 sg13g2_antennanp ANTENNA_191 (.A(_05825_));
 sg13g2_antennanp ANTENNA_192 (.A(_05825_));
 sg13g2_antennanp ANTENNA_193 (.A(_05825_));
 sg13g2_antennanp ANTENNA_194 (.A(_05829_));
 sg13g2_antennanp ANTENNA_195 (.A(_05839_));
 sg13g2_antennanp ANTENNA_196 (.A(_05839_));
 sg13g2_antennanp ANTENNA_197 (.A(_05839_));
 sg13g2_antennanp ANTENNA_198 (.A(_05841_));
 sg13g2_antennanp ANTENNA_199 (.A(_05841_));
 sg13g2_antennanp ANTENNA_200 (.A(_05841_));
 sg13g2_antennanp ANTENNA_201 (.A(_05851_));
 sg13g2_antennanp ANTENNA_202 (.A(_05858_));
 sg13g2_antennanp ANTENNA_203 (.A(_05860_));
 sg13g2_antennanp ANTENNA_204 (.A(_05866_));
 sg13g2_antennanp ANTENNA_205 (.A(_05869_));
 sg13g2_antennanp ANTENNA_206 (.A(_05869_));
 sg13g2_antennanp ANTENNA_207 (.A(_05869_));
 sg13g2_antennanp ANTENNA_208 (.A(_05869_));
 sg13g2_antennanp ANTENNA_209 (.A(_05877_));
 sg13g2_antennanp ANTENNA_210 (.A(_05889_));
 sg13g2_antennanp ANTENNA_211 (.A(_05889_));
 sg13g2_antennanp ANTENNA_212 (.A(_05889_));
 sg13g2_antennanp ANTENNA_213 (.A(_05900_));
 sg13g2_antennanp ANTENNA_214 (.A(_05900_));
 sg13g2_antennanp ANTENNA_215 (.A(_05900_));
 sg13g2_antennanp ANTENNA_216 (.A(_05934_));
 sg13g2_antennanp ANTENNA_217 (.A(_05934_));
 sg13g2_antennanp ANTENNA_218 (.A(_05934_));
 sg13g2_antennanp ANTENNA_219 (.A(_05937_));
 sg13g2_antennanp ANTENNA_220 (.A(_05937_));
 sg13g2_antennanp ANTENNA_221 (.A(_05937_));
 sg13g2_antennanp ANTENNA_222 (.A(_05942_));
 sg13g2_antennanp ANTENNA_223 (.A(_05960_));
 sg13g2_antennanp ANTENNA_224 (.A(_05960_));
 sg13g2_antennanp ANTENNA_225 (.A(_05960_));
 sg13g2_antennanp ANTENNA_226 (.A(_05977_));
 sg13g2_antennanp ANTENNA_227 (.A(_05999_));
 sg13g2_antennanp ANTENNA_228 (.A(_05999_));
 sg13g2_antennanp ANTENNA_229 (.A(_05999_));
 sg13g2_antennanp ANTENNA_230 (.A(_05999_));
 sg13g2_antennanp ANTENNA_231 (.A(_05999_));
 sg13g2_antennanp ANTENNA_232 (.A(_05999_));
 sg13g2_antennanp ANTENNA_233 (.A(_05999_));
 sg13g2_antennanp ANTENNA_234 (.A(_05999_));
 sg13g2_antennanp ANTENNA_235 (.A(_06023_));
 sg13g2_antennanp ANTENNA_236 (.A(_06023_));
 sg13g2_antennanp ANTENNA_237 (.A(_06023_));
 sg13g2_antennanp ANTENNA_238 (.A(_06027_));
 sg13g2_antennanp ANTENNA_239 (.A(_06038_));
 sg13g2_antennanp ANTENNA_240 (.A(_06045_));
 sg13g2_antennanp ANTENNA_241 (.A(_06053_));
 sg13g2_antennanp ANTENNA_242 (.A(_06065_));
 sg13g2_antennanp ANTENNA_243 (.A(_06065_));
 sg13g2_antennanp ANTENNA_244 (.A(_06065_));
 sg13g2_antennanp ANTENNA_245 (.A(_06102_));
 sg13g2_antennanp ANTENNA_246 (.A(_06102_));
 sg13g2_antennanp ANTENNA_247 (.A(_06102_));
 sg13g2_antennanp ANTENNA_248 (.A(_06139_));
 sg13g2_antennanp ANTENNA_249 (.A(_06139_));
 sg13g2_antennanp ANTENNA_250 (.A(_06139_));
 sg13g2_antennanp ANTENNA_251 (.A(_06146_));
 sg13g2_antennanp ANTENNA_252 (.A(_06146_));
 sg13g2_antennanp ANTENNA_253 (.A(_06146_));
 sg13g2_antennanp ANTENNA_254 (.A(_06152_));
 sg13g2_antennanp ANTENNA_255 (.A(_06163_));
 sg13g2_antennanp ANTENNA_256 (.A(_06163_));
 sg13g2_antennanp ANTENNA_257 (.A(_06163_));
 sg13g2_antennanp ANTENNA_258 (.A(_06163_));
 sg13g2_antennanp ANTENNA_259 (.A(_06195_));
 sg13g2_antennanp ANTENNA_260 (.A(_06216_));
 sg13g2_antennanp ANTENNA_261 (.A(_06236_));
 sg13g2_antennanp ANTENNA_262 (.A(_06247_));
 sg13g2_antennanp ANTENNA_263 (.A(_06259_));
 sg13g2_antennanp ANTENNA_264 (.A(_06285_));
 sg13g2_antennanp ANTENNA_265 (.A(_06303_));
 sg13g2_antennanp ANTENNA_266 (.A(_06303_));
 sg13g2_antennanp ANTENNA_267 (.A(_06303_));
 sg13g2_antennanp ANTENNA_268 (.A(_06318_));
 sg13g2_antennanp ANTENNA_269 (.A(_06325_));
 sg13g2_antennanp ANTENNA_270 (.A(_06328_));
 sg13g2_antennanp ANTENNA_271 (.A(_06337_));
 sg13g2_antennanp ANTENNA_272 (.A(_06350_));
 sg13g2_antennanp ANTENNA_273 (.A(_06355_));
 sg13g2_antennanp ANTENNA_274 (.A(_06370_));
 sg13g2_antennanp ANTENNA_275 (.A(_06380_));
 sg13g2_antennanp ANTENNA_276 (.A(_06385_));
 sg13g2_antennanp ANTENNA_277 (.A(_06391_));
 sg13g2_antennanp ANTENNA_278 (.A(_06423_));
 sg13g2_antennanp ANTENNA_279 (.A(_06435_));
 sg13g2_antennanp ANTENNA_280 (.A(_06438_));
 sg13g2_antennanp ANTENNA_281 (.A(_06464_));
 sg13g2_antennanp ANTENNA_282 (.A(_06475_));
 sg13g2_antennanp ANTENNA_283 (.A(_06525_));
 sg13g2_antennanp ANTENNA_284 (.A(_06530_));
 sg13g2_antennanp ANTENNA_285 (.A(_06532_));
 sg13g2_antennanp ANTENNA_286 (.A(_06582_));
 sg13g2_antennanp ANTENNA_287 (.A(_06591_));
 sg13g2_antennanp ANTENNA_288 (.A(_06605_));
 sg13g2_antennanp ANTENNA_289 (.A(_06653_));
 sg13g2_antennanp ANTENNA_290 (.A(_06660_));
 sg13g2_antennanp ANTENNA_291 (.A(_06667_));
 sg13g2_antennanp ANTENNA_292 (.A(_06671_));
 sg13g2_antennanp ANTENNA_293 (.A(_06697_));
 sg13g2_antennanp ANTENNA_294 (.A(_06701_));
 sg13g2_antennanp ANTENNA_295 (.A(_06703_));
 sg13g2_antennanp ANTENNA_296 (.A(_06751_));
 sg13g2_antennanp ANTENNA_297 (.A(_06772_));
 sg13g2_antennanp ANTENNA_298 (.A(_06813_));
 sg13g2_antennanp ANTENNA_299 (.A(_06815_));
 sg13g2_antennanp ANTENNA_300 (.A(_06816_));
 sg13g2_antennanp ANTENNA_301 (.A(_06829_));
 sg13g2_antennanp ANTENNA_302 (.A(_06850_));
 sg13g2_antennanp ANTENNA_303 (.A(_06854_));
 sg13g2_antennanp ANTENNA_304 (.A(_06869_));
 sg13g2_antennanp ANTENNA_305 (.A(_06870_));
 sg13g2_antennanp ANTENNA_306 (.A(_06875_));
 sg13g2_antennanp ANTENNA_307 (.A(_06881_));
 sg13g2_antennanp ANTENNA_308 (.A(_06901_));
 sg13g2_antennanp ANTENNA_309 (.A(_06921_));
 sg13g2_antennanp ANTENNA_310 (.A(_06932_));
 sg13g2_antennanp ANTENNA_311 (.A(_06936_));
 sg13g2_antennanp ANTENNA_312 (.A(_06959_));
 sg13g2_antennanp ANTENNA_313 (.A(_06993_));
 sg13g2_antennanp ANTENNA_314 (.A(_06998_));
 sg13g2_antennanp ANTENNA_315 (.A(_07008_));
 sg13g2_antennanp ANTENNA_316 (.A(_07035_));
 sg13g2_antennanp ANTENNA_317 (.A(_07036_));
 sg13g2_antennanp ANTENNA_318 (.A(_07047_));
 sg13g2_antennanp ANTENNA_319 (.A(_07060_));
 sg13g2_antennanp ANTENNA_320 (.A(_07069_));
 sg13g2_antennanp ANTENNA_321 (.A(_07074_));
 sg13g2_antennanp ANTENNA_322 (.A(_07080_));
 sg13g2_antennanp ANTENNA_323 (.A(_07107_));
 sg13g2_antennanp ANTENNA_324 (.A(_07108_));
 sg13g2_antennanp ANTENNA_325 (.A(_07111_));
 sg13g2_antennanp ANTENNA_326 (.A(_07119_));
 sg13g2_antennanp ANTENNA_327 (.A(_07139_));
 sg13g2_antennanp ANTENNA_328 (.A(_07146_));
 sg13g2_antennanp ANTENNA_329 (.A(_07191_));
 sg13g2_antennanp ANTENNA_330 (.A(_07212_));
 sg13g2_antennanp ANTENNA_331 (.A(_07217_));
 sg13g2_antennanp ANTENNA_332 (.A(_07254_));
 sg13g2_antennanp ANTENNA_333 (.A(_07282_));
 sg13g2_antennanp ANTENNA_334 (.A(_07284_));
 sg13g2_antennanp ANTENNA_335 (.A(_07288_));
 sg13g2_antennanp ANTENNA_336 (.A(_07302_));
 sg13g2_antennanp ANTENNA_337 (.A(_07312_));
 sg13g2_antennanp ANTENNA_338 (.A(_07363_));
 sg13g2_antennanp ANTENNA_339 (.A(_07375_));
 sg13g2_antennanp ANTENNA_340 (.A(_07403_));
 sg13g2_antennanp ANTENNA_341 (.A(_07420_));
 sg13g2_antennanp ANTENNA_342 (.A(_07428_));
 sg13g2_antennanp ANTENNA_343 (.A(_07454_));
 sg13g2_antennanp ANTENNA_344 (.A(_07454_));
 sg13g2_antennanp ANTENNA_345 (.A(_07454_));
 sg13g2_antennanp ANTENNA_346 (.A(_07460_));
 sg13g2_antennanp ANTENNA_347 (.A(_07460_));
 sg13g2_antennanp ANTENNA_348 (.A(_07460_));
 sg13g2_antennanp ANTENNA_349 (.A(_07460_));
 sg13g2_antennanp ANTENNA_350 (.A(_07460_));
 sg13g2_antennanp ANTENNA_351 (.A(_07491_));
 sg13g2_antennanp ANTENNA_352 (.A(_07491_));
 sg13g2_antennanp ANTENNA_353 (.A(_07491_));
 sg13g2_antennanp ANTENNA_354 (.A(_07491_));
 sg13g2_antennanp ANTENNA_355 (.A(_07491_));
 sg13g2_antennanp ANTENNA_356 (.A(_07491_));
 sg13g2_antennanp ANTENNA_357 (.A(_07491_));
 sg13g2_antennanp ANTENNA_358 (.A(_07491_));
 sg13g2_antennanp ANTENNA_359 (.A(_07491_));
 sg13g2_antennanp ANTENNA_360 (.A(_07491_));
 sg13g2_antennanp ANTENNA_361 (.A(_07496_));
 sg13g2_antennanp ANTENNA_362 (.A(_07496_));
 sg13g2_antennanp ANTENNA_363 (.A(_07496_));
 sg13g2_antennanp ANTENNA_364 (.A(_07496_));
 sg13g2_antennanp ANTENNA_365 (.A(_07609_));
 sg13g2_antennanp ANTENNA_366 (.A(_07622_));
 sg13g2_antennanp ANTENNA_367 (.A(_07636_));
 sg13g2_antennanp ANTENNA_368 (.A(_07704_));
 sg13g2_antennanp ANTENNA_369 (.A(_07730_));
 sg13g2_antennanp ANTENNA_370 (.A(_07758_));
 sg13g2_antennanp ANTENNA_371 (.A(_07758_));
 sg13g2_antennanp ANTENNA_372 (.A(_07809_));
 sg13g2_antennanp ANTENNA_373 (.A(_07809_));
 sg13g2_antennanp ANTENNA_374 (.A(_07822_));
 sg13g2_antennanp ANTENNA_375 (.A(_07835_));
 sg13g2_antennanp ANTENNA_376 (.A(_07835_));
 sg13g2_antennanp ANTENNA_377 (.A(_07914_));
 sg13g2_antennanp ANTENNA_378 (.A(_07926_));
 sg13g2_antennanp ANTENNA_379 (.A(_07939_));
 sg13g2_antennanp ANTENNA_380 (.A(_07952_));
 sg13g2_antennanp ANTENNA_381 (.A(_08033_));
 sg13g2_antennanp ANTENNA_382 (.A(_08033_));
 sg13g2_antennanp ANTENNA_383 (.A(_08169_));
 sg13g2_antennanp ANTENNA_384 (.A(_08169_));
 sg13g2_antennanp ANTENNA_385 (.A(_08814_));
 sg13g2_antennanp ANTENNA_386 (.A(_08814_));
 sg13g2_antennanp ANTENNA_387 (.A(_08814_));
 sg13g2_antennanp ANTENNA_388 (.A(_08814_));
 sg13g2_antennanp ANTENNA_389 (.A(_08814_));
 sg13g2_antennanp ANTENNA_390 (.A(_09280_));
 sg13g2_antennanp ANTENNA_391 (.A(_09280_));
 sg13g2_antennanp ANTENNA_392 (.A(_09280_));
 sg13g2_antennanp ANTENNA_393 (.A(_09280_));
 sg13g2_antennanp ANTENNA_394 (.A(_09280_));
 sg13g2_antennanp ANTENNA_395 (.A(_09724_));
 sg13g2_antennanp ANTENNA_396 (.A(_09825_));
 sg13g2_antennanp ANTENNA_397 (.A(_09825_));
 sg13g2_antennanp ANTENNA_398 (.A(_09825_));
 sg13g2_antennanp ANTENNA_399 (.A(_09991_));
 sg13g2_antennanp ANTENNA_400 (.A(_09991_));
 sg13g2_antennanp ANTENNA_401 (.A(_09991_));
 sg13g2_antennanp ANTENNA_402 (.A(_10085_));
 sg13g2_antennanp ANTENNA_403 (.A(_10085_));
 sg13g2_antennanp ANTENNA_404 (.A(_10085_));
 sg13g2_antennanp ANTENNA_405 (.A(_10247_));
 sg13g2_antennanp ANTENNA_406 (.A(_10247_));
 sg13g2_antennanp ANTENNA_407 (.A(_10247_));
 sg13g2_antennanp ANTENNA_408 (.A(_10518_));
 sg13g2_antennanp ANTENNA_409 (.A(_10591_));
 sg13g2_antennanp ANTENNA_410 (.A(_10591_));
 sg13g2_antennanp ANTENNA_411 (.A(_10591_));
 sg13g2_antennanp ANTENNA_412 (.A(_10604_));
 sg13g2_antennanp ANTENNA_413 (.A(_10604_));
 sg13g2_antennanp ANTENNA_414 (.A(_10604_));
 sg13g2_antennanp ANTENNA_415 (.A(_10604_));
 sg13g2_antennanp ANTENNA_416 (.A(_10617_));
 sg13g2_antennanp ANTENNA_417 (.A(_10636_));
 sg13g2_antennanp ANTENNA_418 (.A(_10636_));
 sg13g2_antennanp ANTENNA_419 (.A(_10636_));
 sg13g2_antennanp ANTENNA_420 (.A(_10636_));
 sg13g2_antennanp ANTENNA_421 (.A(_10636_));
 sg13g2_antennanp ANTENNA_422 (.A(_10636_));
 sg13g2_antennanp ANTENNA_423 (.A(_10646_));
 sg13g2_antennanp ANTENNA_424 (.A(_10646_));
 sg13g2_antennanp ANTENNA_425 (.A(_10646_));
 sg13g2_antennanp ANTENNA_426 (.A(_10647_));
 sg13g2_antennanp ANTENNA_427 (.A(_10647_));
 sg13g2_antennanp ANTENNA_428 (.A(_10647_));
 sg13g2_antennanp ANTENNA_429 (.A(_10952_));
 sg13g2_antennanp ANTENNA_430 (.A(_10963_));
 sg13g2_antennanp ANTENNA_431 (.A(_11055_));
 sg13g2_antennanp ANTENNA_432 (.A(_11055_));
 sg13g2_antennanp ANTENNA_433 (.A(_11055_));
 sg13g2_antennanp ANTENNA_434 (.A(_11058_));
 sg13g2_antennanp ANTENNA_435 (.A(_11058_));
 sg13g2_antennanp ANTENNA_436 (.A(_11058_));
 sg13g2_antennanp ANTENNA_437 (.A(_11058_));
 sg13g2_antennanp ANTENNA_438 (.A(_11058_));
 sg13g2_antennanp ANTENNA_439 (.A(_11058_));
 sg13g2_antennanp ANTENNA_440 (.A(_11058_));
 sg13g2_antennanp ANTENNA_441 (.A(_11058_));
 sg13g2_antennanp ANTENNA_442 (.A(_11058_));
 sg13g2_antennanp ANTENNA_443 (.A(_11058_));
 sg13g2_antennanp ANTENNA_444 (.A(_11240_));
 sg13g2_antennanp ANTENNA_445 (.A(_11240_));
 sg13g2_antennanp ANTENNA_446 (.A(_11240_));
 sg13g2_antennanp ANTENNA_447 (.A(_11240_));
 sg13g2_antennanp ANTENNA_448 (.A(_11240_));
 sg13g2_antennanp ANTENNA_449 (.A(_11240_));
 sg13g2_antennanp ANTENNA_450 (.A(_11240_));
 sg13g2_antennanp ANTENNA_451 (.A(_11240_));
 sg13g2_antennanp ANTENNA_452 (.A(_11240_));
 sg13g2_antennanp ANTENNA_453 (.A(_11243_));
 sg13g2_antennanp ANTENNA_454 (.A(_11243_));
 sg13g2_antennanp ANTENNA_455 (.A(_11243_));
 sg13g2_antennanp ANTENNA_456 (.A(_11243_));
 sg13g2_antennanp ANTENNA_457 (.A(_11243_));
 sg13g2_antennanp ANTENNA_458 (.A(_11243_));
 sg13g2_antennanp ANTENNA_459 (.A(_11243_));
 sg13g2_antennanp ANTENNA_460 (.A(_11243_));
 sg13g2_antennanp ANTENNA_461 (.A(_11243_));
 sg13g2_antennanp ANTENNA_462 (.A(\top_ihp.oisc.op_a[22] ));
 sg13g2_antennanp ANTENNA_463 (.A(\top_ihp.oisc.op_a[27] ));
 sg13g2_antennanp ANTENNA_464 (.A(\top_ihp.oisc.op_a[6] ));
 sg13g2_antennanp ANTENNA_465 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_466 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_467 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_468 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_469 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_470 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_471 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_472 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_473 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_474 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_475 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_476 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_477 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_478 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_479 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_480 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_481 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_482 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_483 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_484 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_485 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_486 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_487 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_488 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_489 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_490 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_491 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_492 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_493 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_494 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_495 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_496 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_497 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_498 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_499 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_500 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_501 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_502 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_503 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_504 (.A(\top_ihp.oisc.regs[4][19] ));
 sg13g2_antennanp ANTENNA_505 (.A(\top_ihp.oisc.regs[4][19] ));
 sg13g2_antennanp ANTENNA_506 (.A(\top_ihp.oisc.regs[4][19] ));
 sg13g2_antennanp ANTENNA_507 (.A(\top_ihp.oisc.regs[4][19] ));
 sg13g2_antennanp ANTENNA_508 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_509 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_510 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_511 (.A(\top_ihp.tx ));
 sg13g2_antennanp ANTENNA_512 (.A(net1));
 sg13g2_antennanp ANTENNA_513 (.A(net1));
 sg13g2_antennanp ANTENNA_514 (.A(net1));
 sg13g2_antennanp ANTENNA_515 (.A(net5));
 sg13g2_antennanp ANTENNA_516 (.A(net10));
 sg13g2_antennanp ANTENNA_517 (.A(net37));
 sg13g2_antennanp ANTENNA_518 (.A(net37));
 sg13g2_antennanp ANTENNA_519 (.A(net37));
 sg13g2_antennanp ANTENNA_520 (.A(net37));
 sg13g2_antennanp ANTENNA_521 (.A(net37));
 sg13g2_antennanp ANTENNA_522 (.A(net37));
 sg13g2_antennanp ANTENNA_523 (.A(net37));
 sg13g2_antennanp ANTENNA_524 (.A(net37));
 sg13g2_antennanp ANTENNA_525 (.A(net37));
 sg13g2_antennanp ANTENNA_526 (.A(net67));
 sg13g2_antennanp ANTENNA_527 (.A(net67));
 sg13g2_antennanp ANTENNA_528 (.A(net67));
 sg13g2_antennanp ANTENNA_529 (.A(net67));
 sg13g2_antennanp ANTENNA_530 (.A(net67));
 sg13g2_antennanp ANTENNA_531 (.A(net67));
 sg13g2_antennanp ANTENNA_532 (.A(net67));
 sg13g2_antennanp ANTENNA_533 (.A(net67));
 sg13g2_antennanp ANTENNA_534 (.A(net77));
 sg13g2_antennanp ANTENNA_535 (.A(net77));
 sg13g2_antennanp ANTENNA_536 (.A(net77));
 sg13g2_antennanp ANTENNA_537 (.A(net77));
 sg13g2_antennanp ANTENNA_538 (.A(net77));
 sg13g2_antennanp ANTENNA_539 (.A(net77));
 sg13g2_antennanp ANTENNA_540 (.A(net77));
 sg13g2_antennanp ANTENNA_541 (.A(net77));
 sg13g2_antennanp ANTENNA_542 (.A(net77));
 sg13g2_antennanp ANTENNA_543 (.A(net91));
 sg13g2_antennanp ANTENNA_544 (.A(net91));
 sg13g2_antennanp ANTENNA_545 (.A(net91));
 sg13g2_antennanp ANTENNA_546 (.A(net91));
 sg13g2_antennanp ANTENNA_547 (.A(net91));
 sg13g2_antennanp ANTENNA_548 (.A(net91));
 sg13g2_antennanp ANTENNA_549 (.A(net91));
 sg13g2_antennanp ANTENNA_550 (.A(net91));
 sg13g2_antennanp ANTENNA_551 (.A(net91));
 sg13g2_antennanp ANTENNA_552 (.A(net111));
 sg13g2_antennanp ANTENNA_553 (.A(net111));
 sg13g2_antennanp ANTENNA_554 (.A(net111));
 sg13g2_antennanp ANTENNA_555 (.A(net111));
 sg13g2_antennanp ANTENNA_556 (.A(net111));
 sg13g2_antennanp ANTENNA_557 (.A(net111));
 sg13g2_antennanp ANTENNA_558 (.A(net111));
 sg13g2_antennanp ANTENNA_559 (.A(net111));
 sg13g2_antennanp ANTENNA_560 (.A(net111));
 sg13g2_antennanp ANTENNA_561 (.A(net146));
 sg13g2_antennanp ANTENNA_562 (.A(net146));
 sg13g2_antennanp ANTENNA_563 (.A(net146));
 sg13g2_antennanp ANTENNA_564 (.A(net146));
 sg13g2_antennanp ANTENNA_565 (.A(net146));
 sg13g2_antennanp ANTENNA_566 (.A(net146));
 sg13g2_antennanp ANTENNA_567 (.A(net146));
 sg13g2_antennanp ANTENNA_568 (.A(net146));
 sg13g2_antennanp ANTENNA_569 (.A(net146));
 sg13g2_antennanp ANTENNA_570 (.A(net155));
 sg13g2_antennanp ANTENNA_571 (.A(net155));
 sg13g2_antennanp ANTENNA_572 (.A(net155));
 sg13g2_antennanp ANTENNA_573 (.A(net155));
 sg13g2_antennanp ANTENNA_574 (.A(net155));
 sg13g2_antennanp ANTENNA_575 (.A(net155));
 sg13g2_antennanp ANTENNA_576 (.A(net155));
 sg13g2_antennanp ANTENNA_577 (.A(net155));
 sg13g2_antennanp ANTENNA_578 (.A(net155));
 sg13g2_antennanp ANTENNA_579 (.A(net155));
 sg13g2_antennanp ANTENNA_580 (.A(net155));
 sg13g2_antennanp ANTENNA_581 (.A(net191));
 sg13g2_antennanp ANTENNA_582 (.A(net191));
 sg13g2_antennanp ANTENNA_583 (.A(net191));
 sg13g2_antennanp ANTENNA_584 (.A(net191));
 sg13g2_antennanp ANTENNA_585 (.A(net191));
 sg13g2_antennanp ANTENNA_586 (.A(net191));
 sg13g2_antennanp ANTENNA_587 (.A(net191));
 sg13g2_antennanp ANTENNA_588 (.A(net191));
 sg13g2_antennanp ANTENNA_589 (.A(net191));
 sg13g2_antennanp ANTENNA_590 (.A(net191));
 sg13g2_antennanp ANTENNA_591 (.A(net191));
 sg13g2_antennanp ANTENNA_592 (.A(net191));
 sg13g2_antennanp ANTENNA_593 (.A(net191));
 sg13g2_antennanp ANTENNA_594 (.A(net191));
 sg13g2_antennanp ANTENNA_595 (.A(net191));
 sg13g2_antennanp ANTENNA_596 (.A(net191));
 sg13g2_antennanp ANTENNA_597 (.A(net191));
 sg13g2_antennanp ANTENNA_598 (.A(net191));
 sg13g2_antennanp ANTENNA_599 (.A(net191));
 sg13g2_antennanp ANTENNA_600 (.A(net191));
 sg13g2_antennanp ANTENNA_601 (.A(net191));
 sg13g2_antennanp ANTENNA_602 (.A(net191));
 sg13g2_antennanp ANTENNA_603 (.A(net194));
 sg13g2_antennanp ANTENNA_604 (.A(net194));
 sg13g2_antennanp ANTENNA_605 (.A(net194));
 sg13g2_antennanp ANTENNA_606 (.A(net194));
 sg13g2_antennanp ANTENNA_607 (.A(net194));
 sg13g2_antennanp ANTENNA_608 (.A(net194));
 sg13g2_antennanp ANTENNA_609 (.A(net194));
 sg13g2_antennanp ANTENNA_610 (.A(net194));
 sg13g2_antennanp ANTENNA_611 (.A(net194));
 sg13g2_antennanp ANTENNA_612 (.A(net194));
 sg13g2_antennanp ANTENNA_613 (.A(net194));
 sg13g2_antennanp ANTENNA_614 (.A(net194));
 sg13g2_antennanp ANTENNA_615 (.A(net194));
 sg13g2_antennanp ANTENNA_616 (.A(net194));
 sg13g2_antennanp ANTENNA_617 (.A(net194));
 sg13g2_antennanp ANTENNA_618 (.A(net194));
 sg13g2_antennanp ANTENNA_619 (.A(net194));
 sg13g2_antennanp ANTENNA_620 (.A(net194));
 sg13g2_antennanp ANTENNA_621 (.A(net244));
 sg13g2_antennanp ANTENNA_622 (.A(net244));
 sg13g2_antennanp ANTENNA_623 (.A(net244));
 sg13g2_antennanp ANTENNA_624 (.A(net244));
 sg13g2_antennanp ANTENNA_625 (.A(net244));
 sg13g2_antennanp ANTENNA_626 (.A(net244));
 sg13g2_antennanp ANTENNA_627 (.A(net244));
 sg13g2_antennanp ANTENNA_628 (.A(net244));
 sg13g2_antennanp ANTENNA_629 (.A(net244));
 sg13g2_antennanp ANTENNA_630 (.A(net250));
 sg13g2_antennanp ANTENNA_631 (.A(net250));
 sg13g2_antennanp ANTENNA_632 (.A(net250));
 sg13g2_antennanp ANTENNA_633 (.A(net250));
 sg13g2_antennanp ANTENNA_634 (.A(net250));
 sg13g2_antennanp ANTENNA_635 (.A(net250));
 sg13g2_antennanp ANTENNA_636 (.A(net250));
 sg13g2_antennanp ANTENNA_637 (.A(net250));
 sg13g2_antennanp ANTENNA_638 (.A(net292));
 sg13g2_antennanp ANTENNA_639 (.A(net292));
 sg13g2_antennanp ANTENNA_640 (.A(net292));
 sg13g2_antennanp ANTENNA_641 (.A(net292));
 sg13g2_antennanp ANTENNA_642 (.A(net292));
 sg13g2_antennanp ANTENNA_643 (.A(net292));
 sg13g2_antennanp ANTENNA_644 (.A(net292));
 sg13g2_antennanp ANTENNA_645 (.A(net292));
 sg13g2_antennanp ANTENNA_646 (.A(net292));
 sg13g2_antennanp ANTENNA_647 (.A(net307));
 sg13g2_antennanp ANTENNA_648 (.A(net307));
 sg13g2_antennanp ANTENNA_649 (.A(net307));
 sg13g2_antennanp ANTENNA_650 (.A(net307));
 sg13g2_antennanp ANTENNA_651 (.A(net307));
 sg13g2_antennanp ANTENNA_652 (.A(net307));
 sg13g2_antennanp ANTENNA_653 (.A(net307));
 sg13g2_antennanp ANTENNA_654 (.A(net307));
 sg13g2_antennanp ANTENNA_655 (.A(net307));
 sg13g2_antennanp ANTENNA_656 (.A(net307));
 sg13g2_antennanp ANTENNA_657 (.A(net307));
 sg13g2_antennanp ANTENNA_658 (.A(net308));
 sg13g2_antennanp ANTENNA_659 (.A(net308));
 sg13g2_antennanp ANTENNA_660 (.A(net308));
 sg13g2_antennanp ANTENNA_661 (.A(net308));
 sg13g2_antennanp ANTENNA_662 (.A(net308));
 sg13g2_antennanp ANTENNA_663 (.A(net308));
 sg13g2_antennanp ANTENNA_664 (.A(net308));
 sg13g2_antennanp ANTENNA_665 (.A(net308));
 sg13g2_antennanp ANTENNA_666 (.A(net308));
 sg13g2_antennanp ANTENNA_667 (.A(net317));
 sg13g2_antennanp ANTENNA_668 (.A(net317));
 sg13g2_antennanp ANTENNA_669 (.A(net317));
 sg13g2_antennanp ANTENNA_670 (.A(net317));
 sg13g2_antennanp ANTENNA_671 (.A(net317));
 sg13g2_antennanp ANTENNA_672 (.A(net317));
 sg13g2_antennanp ANTENNA_673 (.A(net317));
 sg13g2_antennanp ANTENNA_674 (.A(net317));
 sg13g2_antennanp ANTENNA_675 (.A(net317));
 sg13g2_antennanp ANTENNA_676 (.A(net356));
 sg13g2_antennanp ANTENNA_677 (.A(net356));
 sg13g2_antennanp ANTENNA_678 (.A(net356));
 sg13g2_antennanp ANTENNA_679 (.A(net356));
 sg13g2_antennanp ANTENNA_680 (.A(net356));
 sg13g2_antennanp ANTENNA_681 (.A(net356));
 sg13g2_antennanp ANTENNA_682 (.A(net356));
 sg13g2_antennanp ANTENNA_683 (.A(net356));
 sg13g2_antennanp ANTENNA_684 (.A(net357));
 sg13g2_antennanp ANTENNA_685 (.A(net357));
 sg13g2_antennanp ANTENNA_686 (.A(net357));
 sg13g2_antennanp ANTENNA_687 (.A(net357));
 sg13g2_antennanp ANTENNA_688 (.A(net357));
 sg13g2_antennanp ANTENNA_689 (.A(net357));
 sg13g2_antennanp ANTENNA_690 (.A(net357));
 sg13g2_antennanp ANTENNA_691 (.A(net357));
 sg13g2_antennanp ANTENNA_692 (.A(net357));
 sg13g2_antennanp ANTENNA_693 (.A(net357));
 sg13g2_antennanp ANTENNA_694 (.A(net357));
 sg13g2_antennanp ANTENNA_695 (.A(net357));
 sg13g2_antennanp ANTENNA_696 (.A(net357));
 sg13g2_antennanp ANTENNA_697 (.A(net357));
 sg13g2_antennanp ANTENNA_698 (.A(net361));
 sg13g2_antennanp ANTENNA_699 (.A(net361));
 sg13g2_antennanp ANTENNA_700 (.A(net361));
 sg13g2_antennanp ANTENNA_701 (.A(net361));
 sg13g2_antennanp ANTENNA_702 (.A(net361));
 sg13g2_antennanp ANTENNA_703 (.A(net361));
 sg13g2_antennanp ANTENNA_704 (.A(net361));
 sg13g2_antennanp ANTENNA_705 (.A(net361));
 sg13g2_antennanp ANTENNA_706 (.A(net361));
 sg13g2_antennanp ANTENNA_707 (.A(net361));
 sg13g2_antennanp ANTENNA_708 (.A(net361));
 sg13g2_antennanp ANTENNA_709 (.A(net361));
 sg13g2_antennanp ANTENNA_710 (.A(net361));
 sg13g2_antennanp ANTENNA_711 (.A(net361));
 sg13g2_antennanp ANTENNA_712 (.A(net361));
 sg13g2_antennanp ANTENNA_713 (.A(net361));
 sg13g2_antennanp ANTENNA_714 (.A(net361));
 sg13g2_antennanp ANTENNA_715 (.A(net361));
 sg13g2_antennanp ANTENNA_716 (.A(net361));
 sg13g2_antennanp ANTENNA_717 (.A(net361));
 sg13g2_antennanp ANTENNA_718 (.A(net369));
 sg13g2_antennanp ANTENNA_719 (.A(net369));
 sg13g2_antennanp ANTENNA_720 (.A(net369));
 sg13g2_antennanp ANTENNA_721 (.A(net369));
 sg13g2_antennanp ANTENNA_722 (.A(net369));
 sg13g2_antennanp ANTENNA_723 (.A(net369));
 sg13g2_antennanp ANTENNA_724 (.A(net369));
 sg13g2_antennanp ANTENNA_725 (.A(net369));
 sg13g2_antennanp ANTENNA_726 (.A(net369));
 sg13g2_antennanp ANTENNA_727 (.A(net369));
 sg13g2_antennanp ANTENNA_728 (.A(net369));
 sg13g2_antennanp ANTENNA_729 (.A(net369));
 sg13g2_antennanp ANTENNA_730 (.A(net369));
 sg13g2_antennanp ANTENNA_731 (.A(net369));
 sg13g2_antennanp ANTENNA_732 (.A(net369));
 sg13g2_antennanp ANTENNA_733 (.A(net369));
 sg13g2_antennanp ANTENNA_734 (.A(net369));
 sg13g2_antennanp ANTENNA_735 (.A(net369));
 sg13g2_antennanp ANTENNA_736 (.A(net369));
 sg13g2_antennanp ANTENNA_737 (.A(net369));
 sg13g2_antennanp ANTENNA_738 (.A(net378));
 sg13g2_antennanp ANTENNA_739 (.A(net378));
 sg13g2_antennanp ANTENNA_740 (.A(net378));
 sg13g2_antennanp ANTENNA_741 (.A(net378));
 sg13g2_antennanp ANTENNA_742 (.A(net378));
 sg13g2_antennanp ANTENNA_743 (.A(net378));
 sg13g2_antennanp ANTENNA_744 (.A(net378));
 sg13g2_antennanp ANTENNA_745 (.A(net378));
 sg13g2_antennanp ANTENNA_746 (.A(net381));
 sg13g2_antennanp ANTENNA_747 (.A(net381));
 sg13g2_antennanp ANTENNA_748 (.A(net381));
 sg13g2_antennanp ANTENNA_749 (.A(net381));
 sg13g2_antennanp ANTENNA_750 (.A(net381));
 sg13g2_antennanp ANTENNA_751 (.A(net381));
 sg13g2_antennanp ANTENNA_752 (.A(net381));
 sg13g2_antennanp ANTENNA_753 (.A(net381));
 sg13g2_antennanp ANTENNA_754 (.A(net381));
 sg13g2_antennanp ANTENNA_755 (.A(net381));
 sg13g2_antennanp ANTENNA_756 (.A(net381));
 sg13g2_antennanp ANTENNA_757 (.A(net381));
 sg13g2_antennanp ANTENNA_758 (.A(net381));
 sg13g2_antennanp ANTENNA_759 (.A(net381));
 sg13g2_antennanp ANTENNA_760 (.A(net383));
 sg13g2_antennanp ANTENNA_761 (.A(net383));
 sg13g2_antennanp ANTENNA_762 (.A(net383));
 sg13g2_antennanp ANTENNA_763 (.A(net383));
 sg13g2_antennanp ANTENNA_764 (.A(net383));
 sg13g2_antennanp ANTENNA_765 (.A(net383));
 sg13g2_antennanp ANTENNA_766 (.A(net383));
 sg13g2_antennanp ANTENNA_767 (.A(net383));
 sg13g2_antennanp ANTENNA_768 (.A(net384));
 sg13g2_antennanp ANTENNA_769 (.A(net384));
 sg13g2_antennanp ANTENNA_770 (.A(net384));
 sg13g2_antennanp ANTENNA_771 (.A(net384));
 sg13g2_antennanp ANTENNA_772 (.A(net384));
 sg13g2_antennanp ANTENNA_773 (.A(net384));
 sg13g2_antennanp ANTENNA_774 (.A(net384));
 sg13g2_antennanp ANTENNA_775 (.A(net384));
 sg13g2_antennanp ANTENNA_776 (.A(net397));
 sg13g2_antennanp ANTENNA_777 (.A(net397));
 sg13g2_antennanp ANTENNA_778 (.A(net397));
 sg13g2_antennanp ANTENNA_779 (.A(net397));
 sg13g2_antennanp ANTENNA_780 (.A(net397));
 sg13g2_antennanp ANTENNA_781 (.A(net397));
 sg13g2_antennanp ANTENNA_782 (.A(net397));
 sg13g2_antennanp ANTENNA_783 (.A(net397));
 sg13g2_antennanp ANTENNA_784 (.A(net397));
 sg13g2_antennanp ANTENNA_785 (.A(net397));
 sg13g2_antennanp ANTENNA_786 (.A(net397));
 sg13g2_antennanp ANTENNA_787 (.A(net397));
 sg13g2_antennanp ANTENNA_788 (.A(net397));
 sg13g2_antennanp ANTENNA_789 (.A(net397));
 sg13g2_antennanp ANTENNA_790 (.A(net397));
 sg13g2_antennanp ANTENNA_791 (.A(net412));
 sg13g2_antennanp ANTENNA_792 (.A(net412));
 sg13g2_antennanp ANTENNA_793 (.A(net412));
 sg13g2_antennanp ANTENNA_794 (.A(net412));
 sg13g2_antennanp ANTENNA_795 (.A(net412));
 sg13g2_antennanp ANTENNA_796 (.A(net412));
 sg13g2_antennanp ANTENNA_797 (.A(net412));
 sg13g2_antennanp ANTENNA_798 (.A(net412));
 sg13g2_antennanp ANTENNA_799 (.A(net412));
 sg13g2_antennanp ANTENNA_800 (.A(net412));
 sg13g2_antennanp ANTENNA_801 (.A(net412));
 sg13g2_antennanp ANTENNA_802 (.A(net412));
 sg13g2_antennanp ANTENNA_803 (.A(net412));
 sg13g2_antennanp ANTENNA_804 (.A(net412));
 sg13g2_antennanp ANTENNA_805 (.A(net412));
 sg13g2_antennanp ANTENNA_806 (.A(net427));
 sg13g2_antennanp ANTENNA_807 (.A(net427));
 sg13g2_antennanp ANTENNA_808 (.A(net427));
 sg13g2_antennanp ANTENNA_809 (.A(net427));
 sg13g2_antennanp ANTENNA_810 (.A(net427));
 sg13g2_antennanp ANTENNA_811 (.A(net427));
 sg13g2_antennanp ANTENNA_812 (.A(net427));
 sg13g2_antennanp ANTENNA_813 (.A(net427));
 sg13g2_antennanp ANTENNA_814 (.A(net427));
 sg13g2_antennanp ANTENNA_815 (.A(net427));
 sg13g2_antennanp ANTENNA_816 (.A(net427));
 sg13g2_antennanp ANTENNA_817 (.A(net427));
 sg13g2_antennanp ANTENNA_818 (.A(net427));
 sg13g2_antennanp ANTENNA_819 (.A(net427));
 sg13g2_antennanp ANTENNA_820 (.A(net427));
 sg13g2_antennanp ANTENNA_821 (.A(net427));
 sg13g2_antennanp ANTENNA_822 (.A(net427));
 sg13g2_antennanp ANTENNA_823 (.A(net427));
 sg13g2_antennanp ANTENNA_824 (.A(net427));
 sg13g2_antennanp ANTENNA_825 (.A(net427));
 sg13g2_antennanp ANTENNA_826 (.A(net427));
 sg13g2_antennanp ANTENNA_827 (.A(net427));
 sg13g2_antennanp ANTENNA_828 (.A(net427));
 sg13g2_antennanp ANTENNA_829 (.A(net436));
 sg13g2_antennanp ANTENNA_830 (.A(net436));
 sg13g2_antennanp ANTENNA_831 (.A(net436));
 sg13g2_antennanp ANTENNA_832 (.A(net436));
 sg13g2_antennanp ANTENNA_833 (.A(net436));
 sg13g2_antennanp ANTENNA_834 (.A(net436));
 sg13g2_antennanp ANTENNA_835 (.A(net436));
 sg13g2_antennanp ANTENNA_836 (.A(net436));
 sg13g2_antennanp ANTENNA_837 (.A(net498));
 sg13g2_antennanp ANTENNA_838 (.A(net498));
 sg13g2_antennanp ANTENNA_839 (.A(net498));
 sg13g2_antennanp ANTENNA_840 (.A(net498));
 sg13g2_antennanp ANTENNA_841 (.A(net498));
 sg13g2_antennanp ANTENNA_842 (.A(net498));
 sg13g2_antennanp ANTENNA_843 (.A(net498));
 sg13g2_antennanp ANTENNA_844 (.A(net498));
 sg13g2_antennanp ANTENNA_845 (.A(net498));
 sg13g2_antennanp ANTENNA_846 (.A(net525));
 sg13g2_antennanp ANTENNA_847 (.A(net525));
 sg13g2_antennanp ANTENNA_848 (.A(net525));
 sg13g2_antennanp ANTENNA_849 (.A(net525));
 sg13g2_antennanp ANTENNA_850 (.A(net525));
 sg13g2_antennanp ANTENNA_851 (.A(net525));
 sg13g2_antennanp ANTENNA_852 (.A(net525));
 sg13g2_antennanp ANTENNA_853 (.A(net525));
 sg13g2_antennanp ANTENNA_854 (.A(net725));
 sg13g2_antennanp ANTENNA_855 (.A(net725));
 sg13g2_antennanp ANTENNA_856 (.A(net725));
 sg13g2_antennanp ANTENNA_857 (.A(net725));
 sg13g2_antennanp ANTENNA_858 (.A(net725));
 sg13g2_antennanp ANTENNA_859 (.A(net725));
 sg13g2_antennanp ANTENNA_860 (.A(net725));
 sg13g2_antennanp ANTENNA_861 (.A(net725));
 sg13g2_antennanp ANTENNA_862 (.A(net725));
 sg13g2_antennanp ANTENNA_863 (.A(net749));
 sg13g2_antennanp ANTENNA_864 (.A(net749));
 sg13g2_antennanp ANTENNA_865 (.A(net749));
 sg13g2_antennanp ANTENNA_866 (.A(net749));
 sg13g2_antennanp ANTENNA_867 (.A(net749));
 sg13g2_antennanp ANTENNA_868 (.A(net749));
 sg13g2_antennanp ANTENNA_869 (.A(net749));
 sg13g2_antennanp ANTENNA_870 (.A(net749));
 sg13g2_antennanp ANTENNA_871 (.A(net803));
 sg13g2_antennanp ANTENNA_872 (.A(net803));
 sg13g2_antennanp ANTENNA_873 (.A(net803));
 sg13g2_antennanp ANTENNA_874 (.A(net803));
 sg13g2_antennanp ANTENNA_875 (.A(net803));
 sg13g2_antennanp ANTENNA_876 (.A(net803));
 sg13g2_antennanp ANTENNA_877 (.A(net803));
 sg13g2_antennanp ANTENNA_878 (.A(net803));
 sg13g2_antennanp ANTENNA_879 (.A(net803));
 sg13g2_antennanp ANTENNA_880 (.A(net1061));
 sg13g2_antennanp ANTENNA_881 (.A(net1061));
 sg13g2_antennanp ANTENNA_882 (.A(net1061));
 sg13g2_antennanp ANTENNA_883 (.A(net1061));
 sg13g2_antennanp ANTENNA_884 (.A(net1061));
 sg13g2_antennanp ANTENNA_885 (.A(net1061));
 sg13g2_antennanp ANTENNA_886 (.A(net1061));
 sg13g2_antennanp ANTENNA_887 (.A(net1061));
 sg13g2_antennanp ANTENNA_888 (.A(net1061));
 sg13g2_antennanp ANTENNA_889 (.A(net1207));
 sg13g2_antennanp ANTENNA_890 (.A(net1207));
 sg13g2_antennanp ANTENNA_891 (.A(net1207));
 sg13g2_antennanp ANTENNA_892 (.A(net1207));
 sg13g2_antennanp ANTENNA_893 (.A(net1207));
 sg13g2_antennanp ANTENNA_894 (.A(net1207));
 sg13g2_antennanp ANTENNA_895 (.A(_00366_));
 sg13g2_antennanp ANTENNA_896 (.A(_00366_));
 sg13g2_antennanp ANTENNA_897 (.A(_00394_));
 sg13g2_antennanp ANTENNA_898 (.A(_00394_));
 sg13g2_antennanp ANTENNA_899 (.A(_00394_));
 sg13g2_antennanp ANTENNA_900 (.A(_00406_));
 sg13g2_antennanp ANTENNA_901 (.A(_00406_));
 sg13g2_antennanp ANTENNA_902 (.A(_00408_));
 sg13g2_antennanp ANTENNA_903 (.A(_00411_));
 sg13g2_antennanp ANTENNA_904 (.A(_00412_));
 sg13g2_antennanp ANTENNA_905 (.A(_00413_));
 sg13g2_antennanp ANTENNA_906 (.A(_00413_));
 sg13g2_antennanp ANTENNA_907 (.A(_00417_));
 sg13g2_antennanp ANTENNA_908 (.A(_03004_));
 sg13g2_antennanp ANTENNA_909 (.A(_03004_));
 sg13g2_antennanp ANTENNA_910 (.A(_03004_));
 sg13g2_antennanp ANTENNA_911 (.A(_03038_));
 sg13g2_antennanp ANTENNA_912 (.A(_03038_));
 sg13g2_antennanp ANTENNA_913 (.A(_03038_));
 sg13g2_antennanp ANTENNA_914 (.A(_03038_));
 sg13g2_antennanp ANTENNA_915 (.A(_03063_));
 sg13g2_antennanp ANTENNA_916 (.A(_03063_));
 sg13g2_antennanp ANTENNA_917 (.A(_03063_));
 sg13g2_antennanp ANTENNA_918 (.A(_03063_));
 sg13g2_antennanp ANTENNA_919 (.A(_03145_));
 sg13g2_antennanp ANTENNA_920 (.A(_03451_));
 sg13g2_antennanp ANTENNA_921 (.A(_03451_));
 sg13g2_antennanp ANTENNA_922 (.A(_03451_));
 sg13g2_antennanp ANTENNA_923 (.A(_03451_));
 sg13g2_antennanp ANTENNA_924 (.A(_03451_));
 sg13g2_antennanp ANTENNA_925 (.A(_03451_));
 sg13g2_antennanp ANTENNA_926 (.A(_04085_));
 sg13g2_antennanp ANTENNA_927 (.A(_04085_));
 sg13g2_antennanp ANTENNA_928 (.A(_04085_));
 sg13g2_antennanp ANTENNA_929 (.A(_04085_));
 sg13g2_antennanp ANTENNA_930 (.A(_04086_));
 sg13g2_antennanp ANTENNA_931 (.A(_04086_));
 sg13g2_antennanp ANTENNA_932 (.A(_04086_));
 sg13g2_antennanp ANTENNA_933 (.A(_04107_));
 sg13g2_antennanp ANTENNA_934 (.A(_04743_));
 sg13g2_antennanp ANTENNA_935 (.A(_04743_));
 sg13g2_antennanp ANTENNA_936 (.A(_05436_));
 sg13g2_antennanp ANTENNA_937 (.A(_05436_));
 sg13g2_antennanp ANTENNA_938 (.A(_05436_));
 sg13g2_antennanp ANTENNA_939 (.A(_05436_));
 sg13g2_antennanp ANTENNA_940 (.A(_05495_));
 sg13g2_antennanp ANTENNA_941 (.A(_05495_));
 sg13g2_antennanp ANTENNA_942 (.A(_05531_));
 sg13g2_antennanp ANTENNA_943 (.A(_05531_));
 sg13g2_antennanp ANTENNA_944 (.A(_05531_));
 sg13g2_antennanp ANTENNA_945 (.A(_05531_));
 sg13g2_antennanp ANTENNA_946 (.A(_05531_));
 sg13g2_antennanp ANTENNA_947 (.A(_05531_));
 sg13g2_antennanp ANTENNA_948 (.A(_05531_));
 sg13g2_antennanp ANTENNA_949 (.A(_05531_));
 sg13g2_antennanp ANTENNA_950 (.A(_05582_));
 sg13g2_antennanp ANTENNA_951 (.A(_05582_));
 sg13g2_antennanp ANTENNA_952 (.A(_05582_));
 sg13g2_antennanp ANTENNA_953 (.A(_05582_));
 sg13g2_antennanp ANTENNA_954 (.A(_05582_));
 sg13g2_antennanp ANTENNA_955 (.A(_05582_));
 sg13g2_antennanp ANTENNA_956 (.A(_05582_));
 sg13g2_antennanp ANTENNA_957 (.A(_05592_));
 sg13g2_antennanp ANTENNA_958 (.A(_05621_));
 sg13g2_antennanp ANTENNA_959 (.A(_05631_));
 sg13g2_antennanp ANTENNA_960 (.A(_05639_));
 sg13g2_antennanp ANTENNA_961 (.A(_05648_));
 sg13g2_antennanp ANTENNA_962 (.A(_05648_));
 sg13g2_antennanp ANTENNA_963 (.A(_05648_));
 sg13g2_antennanp ANTENNA_964 (.A(_05689_));
 sg13g2_antennanp ANTENNA_965 (.A(_05719_));
 sg13g2_antennanp ANTENNA_966 (.A(_05719_));
 sg13g2_antennanp ANTENNA_967 (.A(_05719_));
 sg13g2_antennanp ANTENNA_968 (.A(_05719_));
 sg13g2_antennanp ANTENNA_969 (.A(_05719_));
 sg13g2_antennanp ANTENNA_970 (.A(_05729_));
 sg13g2_antennanp ANTENNA_971 (.A(_05729_));
 sg13g2_antennanp ANTENNA_972 (.A(_05729_));
 sg13g2_antennanp ANTENNA_973 (.A(_05735_));
 sg13g2_antennanp ANTENNA_974 (.A(_05735_));
 sg13g2_antennanp ANTENNA_975 (.A(_05735_));
 sg13g2_antennanp ANTENNA_976 (.A(_05735_));
 sg13g2_antennanp ANTENNA_977 (.A(_05735_));
 sg13g2_antennanp ANTENNA_978 (.A(_05735_));
 sg13g2_antennanp ANTENNA_979 (.A(_05735_));
 sg13g2_antennanp ANTENNA_980 (.A(_05735_));
 sg13g2_antennanp ANTENNA_981 (.A(_05739_));
 sg13g2_antennanp ANTENNA_982 (.A(_05773_));
 sg13g2_antennanp ANTENNA_983 (.A(_05781_));
 sg13g2_antennanp ANTENNA_984 (.A(_05782_));
 sg13g2_antennanp ANTENNA_985 (.A(_05782_));
 sg13g2_antennanp ANTENNA_986 (.A(_05782_));
 sg13g2_antennanp ANTENNA_987 (.A(_05785_));
 sg13g2_antennanp ANTENNA_988 (.A(_05807_));
 sg13g2_antennanp ANTENNA_989 (.A(_05825_));
 sg13g2_antennanp ANTENNA_990 (.A(_05825_));
 sg13g2_antennanp ANTENNA_991 (.A(_05825_));
 sg13g2_antennanp ANTENNA_992 (.A(_05829_));
 sg13g2_antennanp ANTENNA_993 (.A(_05841_));
 sg13g2_antennanp ANTENNA_994 (.A(_05841_));
 sg13g2_antennanp ANTENNA_995 (.A(_05841_));
 sg13g2_antennanp ANTENNA_996 (.A(_05851_));
 sg13g2_antennanp ANTENNA_997 (.A(_05858_));
 sg13g2_antennanp ANTENNA_998 (.A(_05866_));
 sg13g2_antennanp ANTENNA_999 (.A(_05869_));
 sg13g2_antennanp ANTENNA_1000 (.A(_05869_));
 sg13g2_antennanp ANTENNA_1001 (.A(_05869_));
 sg13g2_antennanp ANTENNA_1002 (.A(_05877_));
 sg13g2_antennanp ANTENNA_1003 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1004 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1005 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1006 (.A(_05934_));
 sg13g2_antennanp ANTENNA_1007 (.A(_05934_));
 sg13g2_antennanp ANTENNA_1008 (.A(_05934_));
 sg13g2_antennanp ANTENNA_1009 (.A(_05942_));
 sg13g2_antennanp ANTENNA_1010 (.A(_05960_));
 sg13g2_antennanp ANTENNA_1011 (.A(_05960_));
 sg13g2_antennanp ANTENNA_1012 (.A(_05960_));
 sg13g2_antennanp ANTENNA_1013 (.A(_05977_));
 sg13g2_antennanp ANTENNA_1014 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1015 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1016 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1017 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1018 (.A(_06027_));
 sg13g2_antennanp ANTENNA_1019 (.A(_06038_));
 sg13g2_antennanp ANTENNA_1020 (.A(_06045_));
 sg13g2_antennanp ANTENNA_1021 (.A(_06053_));
 sg13g2_antennanp ANTENNA_1022 (.A(_06065_));
 sg13g2_antennanp ANTENNA_1023 (.A(_06065_));
 sg13g2_antennanp ANTENNA_1024 (.A(_06065_));
 sg13g2_antennanp ANTENNA_1025 (.A(_06102_));
 sg13g2_antennanp ANTENNA_1026 (.A(_06102_));
 sg13g2_antennanp ANTENNA_1027 (.A(_06102_));
 sg13g2_antennanp ANTENNA_1028 (.A(_06102_));
 sg13g2_antennanp ANTENNA_1029 (.A(_06102_));
 sg13g2_antennanp ANTENNA_1030 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1031 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1032 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1033 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1034 (.A(_06152_));
 sg13g2_antennanp ANTENNA_1035 (.A(_06163_));
 sg13g2_antennanp ANTENNA_1036 (.A(_06163_));
 sg13g2_antennanp ANTENNA_1037 (.A(_06163_));
 sg13g2_antennanp ANTENNA_1038 (.A(_06183_));
 sg13g2_antennanp ANTENNA_1039 (.A(_06183_));
 sg13g2_antennanp ANTENNA_1040 (.A(_06183_));
 sg13g2_antennanp ANTENNA_1041 (.A(_06183_));
 sg13g2_antennanp ANTENNA_1042 (.A(_06195_));
 sg13g2_antennanp ANTENNA_1043 (.A(_06216_));
 sg13g2_antennanp ANTENNA_1044 (.A(_06236_));
 sg13g2_antennanp ANTENNA_1045 (.A(_06247_));
 sg13g2_antennanp ANTENNA_1046 (.A(_06259_));
 sg13g2_antennanp ANTENNA_1047 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1048 (.A(_06303_));
 sg13g2_antennanp ANTENNA_1049 (.A(_06318_));
 sg13g2_antennanp ANTENNA_1050 (.A(_06337_));
 sg13g2_antennanp ANTENNA_1051 (.A(_06350_));
 sg13g2_antennanp ANTENNA_1052 (.A(_06355_));
 sg13g2_antennanp ANTENNA_1053 (.A(_06370_));
 sg13g2_antennanp ANTENNA_1054 (.A(_06385_));
 sg13g2_antennanp ANTENNA_1055 (.A(_06391_));
 sg13g2_antennanp ANTENNA_1056 (.A(_06423_));
 sg13g2_antennanp ANTENNA_1057 (.A(_06435_));
 sg13g2_antennanp ANTENNA_1058 (.A(_06438_));
 sg13g2_antennanp ANTENNA_1059 (.A(_06464_));
 sg13g2_antennanp ANTENNA_1060 (.A(_06475_));
 sg13g2_antennanp ANTENNA_1061 (.A(_06525_));
 sg13g2_antennanp ANTENNA_1062 (.A(_06530_));
 sg13g2_antennanp ANTENNA_1063 (.A(_06532_));
 sg13g2_antennanp ANTENNA_1064 (.A(_06582_));
 sg13g2_antennanp ANTENNA_1065 (.A(_06605_));
 sg13g2_antennanp ANTENNA_1066 (.A(_06653_));
 sg13g2_antennanp ANTENNA_1067 (.A(_06660_));
 sg13g2_antennanp ANTENNA_1068 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1069 (.A(_06671_));
 sg13g2_antennanp ANTENNA_1070 (.A(_06697_));
 sg13g2_antennanp ANTENNA_1071 (.A(_06701_));
 sg13g2_antennanp ANTENNA_1072 (.A(_06703_));
 sg13g2_antennanp ANTENNA_1073 (.A(_06751_));
 sg13g2_antennanp ANTENNA_1074 (.A(_06772_));
 sg13g2_antennanp ANTENNA_1075 (.A(_06772_));
 sg13g2_antennanp ANTENNA_1076 (.A(_06813_));
 sg13g2_antennanp ANTENNA_1077 (.A(_06815_));
 sg13g2_antennanp ANTENNA_1078 (.A(_06815_));
 sg13g2_antennanp ANTENNA_1079 (.A(_06816_));
 sg13g2_antennanp ANTENNA_1080 (.A(_06829_));
 sg13g2_antennanp ANTENNA_1081 (.A(_06850_));
 sg13g2_antennanp ANTENNA_1082 (.A(_06854_));
 sg13g2_antennanp ANTENNA_1083 (.A(_06869_));
 sg13g2_antennanp ANTENNA_1084 (.A(_06870_));
 sg13g2_antennanp ANTENNA_1085 (.A(_06875_));
 sg13g2_antennanp ANTENNA_1086 (.A(_06881_));
 sg13g2_antennanp ANTENNA_1087 (.A(_06901_));
 sg13g2_antennanp ANTENNA_1088 (.A(_06921_));
 sg13g2_antennanp ANTENNA_1089 (.A(_06932_));
 sg13g2_antennanp ANTENNA_1090 (.A(_06936_));
 sg13g2_antennanp ANTENNA_1091 (.A(_06959_));
 sg13g2_antennanp ANTENNA_1092 (.A(_06993_));
 sg13g2_antennanp ANTENNA_1093 (.A(_06998_));
 sg13g2_antennanp ANTENNA_1094 (.A(_07008_));
 sg13g2_antennanp ANTENNA_1095 (.A(_07035_));
 sg13g2_antennanp ANTENNA_1096 (.A(_07036_));
 sg13g2_antennanp ANTENNA_1097 (.A(_07047_));
 sg13g2_antennanp ANTENNA_1098 (.A(_07060_));
 sg13g2_antennanp ANTENNA_1099 (.A(_07069_));
 sg13g2_antennanp ANTENNA_1100 (.A(_07074_));
 sg13g2_antennanp ANTENNA_1101 (.A(_07080_));
 sg13g2_antennanp ANTENNA_1102 (.A(_07108_));
 sg13g2_antennanp ANTENNA_1103 (.A(_07111_));
 sg13g2_antennanp ANTENNA_1104 (.A(_07139_));
 sg13g2_antennanp ANTENNA_1105 (.A(_07146_));
 sg13g2_antennanp ANTENNA_1106 (.A(_07191_));
 sg13g2_antennanp ANTENNA_1107 (.A(_07212_));
 sg13g2_antennanp ANTENNA_1108 (.A(_07217_));
 sg13g2_antennanp ANTENNA_1109 (.A(_07254_));
 sg13g2_antennanp ANTENNA_1110 (.A(_07282_));
 sg13g2_antennanp ANTENNA_1111 (.A(_07284_));
 sg13g2_antennanp ANTENNA_1112 (.A(_07288_));
 sg13g2_antennanp ANTENNA_1113 (.A(_07302_));
 sg13g2_antennanp ANTENNA_1114 (.A(_07312_));
 sg13g2_antennanp ANTENNA_1115 (.A(_07363_));
 sg13g2_antennanp ANTENNA_1116 (.A(_07375_));
 sg13g2_antennanp ANTENNA_1117 (.A(_07403_));
 sg13g2_antennanp ANTENNA_1118 (.A(_07420_));
 sg13g2_antennanp ANTENNA_1119 (.A(_07420_));
 sg13g2_antennanp ANTENNA_1120 (.A(_07428_));
 sg13g2_antennanp ANTENNA_1121 (.A(_07460_));
 sg13g2_antennanp ANTENNA_1122 (.A(_07460_));
 sg13g2_antennanp ANTENNA_1123 (.A(_07460_));
 sg13g2_antennanp ANTENNA_1124 (.A(_07460_));
 sg13g2_antennanp ANTENNA_1125 (.A(_07460_));
 sg13g2_antennanp ANTENNA_1126 (.A(_07491_));
 sg13g2_antennanp ANTENNA_1127 (.A(_07491_));
 sg13g2_antennanp ANTENNA_1128 (.A(_07491_));
 sg13g2_antennanp ANTENNA_1129 (.A(_07491_));
 sg13g2_antennanp ANTENNA_1130 (.A(_07491_));
 sg13g2_antennanp ANTENNA_1131 (.A(_07491_));
 sg13g2_antennanp ANTENNA_1132 (.A(_07496_));
 sg13g2_antennanp ANTENNA_1133 (.A(_07496_));
 sg13g2_antennanp ANTENNA_1134 (.A(_07496_));
 sg13g2_antennanp ANTENNA_1135 (.A(_07496_));
 sg13g2_antennanp ANTENNA_1136 (.A(_07609_));
 sg13g2_antennanp ANTENNA_1137 (.A(_07622_));
 sg13g2_antennanp ANTENNA_1138 (.A(_07636_));
 sg13g2_antennanp ANTENNA_1139 (.A(_07704_));
 sg13g2_antennanp ANTENNA_1140 (.A(_07704_));
 sg13g2_antennanp ANTENNA_1141 (.A(_07730_));
 sg13g2_antennanp ANTENNA_1142 (.A(_07758_));
 sg13g2_antennanp ANTENNA_1143 (.A(_07822_));
 sg13g2_antennanp ANTENNA_1144 (.A(_07835_));
 sg13g2_antennanp ANTENNA_1145 (.A(_07835_));
 sg13g2_antennanp ANTENNA_1146 (.A(_07914_));
 sg13g2_antennanp ANTENNA_1147 (.A(_07926_));
 sg13g2_antennanp ANTENNA_1148 (.A(_07939_));
 sg13g2_antennanp ANTENNA_1149 (.A(_07952_));
 sg13g2_antennanp ANTENNA_1150 (.A(_08169_));
 sg13g2_antennanp ANTENNA_1151 (.A(_08169_));
 sg13g2_antennanp ANTENNA_1152 (.A(_09280_));
 sg13g2_antennanp ANTENNA_1153 (.A(_09280_));
 sg13g2_antennanp ANTENNA_1154 (.A(_09280_));
 sg13g2_antennanp ANTENNA_1155 (.A(_09280_));
 sg13g2_antennanp ANTENNA_1156 (.A(_09280_));
 sg13g2_antennanp ANTENNA_1157 (.A(_09724_));
 sg13g2_antennanp ANTENNA_1158 (.A(_09825_));
 sg13g2_antennanp ANTENNA_1159 (.A(_09825_));
 sg13g2_antennanp ANTENNA_1160 (.A(_09825_));
 sg13g2_antennanp ANTENNA_1161 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1162 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1163 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1164 (.A(_10247_));
 sg13g2_antennanp ANTENNA_1165 (.A(_10247_));
 sg13g2_antennanp ANTENNA_1166 (.A(_10247_));
 sg13g2_antennanp ANTENNA_1167 (.A(_10518_));
 sg13g2_antennanp ANTENNA_1168 (.A(_10604_));
 sg13g2_antennanp ANTENNA_1169 (.A(_10604_));
 sg13g2_antennanp ANTENNA_1170 (.A(_10604_));
 sg13g2_antennanp ANTENNA_1171 (.A(_10604_));
 sg13g2_antennanp ANTENNA_1172 (.A(_10617_));
 sg13g2_antennanp ANTENNA_1173 (.A(_10636_));
 sg13g2_antennanp ANTENNA_1174 (.A(_10636_));
 sg13g2_antennanp ANTENNA_1175 (.A(_10636_));
 sg13g2_antennanp ANTENNA_1176 (.A(_10636_));
 sg13g2_antennanp ANTENNA_1177 (.A(_10636_));
 sg13g2_antennanp ANTENNA_1178 (.A(_10636_));
 sg13g2_antennanp ANTENNA_1179 (.A(_10636_));
 sg13g2_antennanp ANTENNA_1180 (.A(_10636_));
 sg13g2_antennanp ANTENNA_1181 (.A(_10636_));
 sg13g2_antennanp ANTENNA_1182 (.A(_10647_));
 sg13g2_antennanp ANTENNA_1183 (.A(_10647_));
 sg13g2_antennanp ANTENNA_1184 (.A(_10647_));
 sg13g2_antennanp ANTENNA_1185 (.A(_10952_));
 sg13g2_antennanp ANTENNA_1186 (.A(_10963_));
 sg13g2_antennanp ANTENNA_1187 (.A(_11060_));
 sg13g2_antennanp ANTENNA_1188 (.A(_11060_));
 sg13g2_antennanp ANTENNA_1189 (.A(_11060_));
 sg13g2_antennanp ANTENNA_1190 (.A(_11060_));
 sg13g2_antennanp ANTENNA_1191 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1192 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1193 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1194 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1195 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1196 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1197 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1198 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1199 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1200 (.A(\top_ihp.oisc.op_a[22] ));
 sg13g2_antennanp ANTENNA_1201 (.A(\top_ihp.oisc.op_a[27] ));
 sg13g2_antennanp ANTENNA_1202 (.A(\top_ihp.oisc.op_a[6] ));
 sg13g2_antennanp ANTENNA_1203 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_1204 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_1205 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_1206 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_1207 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_1208 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_1209 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_1210 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_1211 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_1212 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_1213 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_1214 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_1215 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_1216 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_1217 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_1218 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_1219 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_1220 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_1221 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_1222 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_1223 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_1224 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_1225 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_1226 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_1227 (.A(\top_ihp.tx ));
 sg13g2_antennanp ANTENNA_1228 (.A(net1));
 sg13g2_antennanp ANTENNA_1229 (.A(net1));
 sg13g2_antennanp ANTENNA_1230 (.A(net1));
 sg13g2_antennanp ANTENNA_1231 (.A(net5));
 sg13g2_antennanp ANTENNA_1232 (.A(net10));
 sg13g2_antennanp ANTENNA_1233 (.A(net63));
 sg13g2_antennanp ANTENNA_1234 (.A(net63));
 sg13g2_antennanp ANTENNA_1235 (.A(net63));
 sg13g2_antennanp ANTENNA_1236 (.A(net63));
 sg13g2_antennanp ANTENNA_1237 (.A(net63));
 sg13g2_antennanp ANTENNA_1238 (.A(net63));
 sg13g2_antennanp ANTENNA_1239 (.A(net63));
 sg13g2_antennanp ANTENNA_1240 (.A(net63));
 sg13g2_antennanp ANTENNA_1241 (.A(net63));
 sg13g2_antennanp ANTENNA_1242 (.A(net63));
 sg13g2_antennanp ANTENNA_1243 (.A(net63));
 sg13g2_antennanp ANTENNA_1244 (.A(net63));
 sg13g2_antennanp ANTENNA_1245 (.A(net63));
 sg13g2_antennanp ANTENNA_1246 (.A(net63));
 sg13g2_antennanp ANTENNA_1247 (.A(net63));
 sg13g2_antennanp ANTENNA_1248 (.A(net63));
 sg13g2_antennanp ANTENNA_1249 (.A(net63));
 sg13g2_antennanp ANTENNA_1250 (.A(net63));
 sg13g2_antennanp ANTENNA_1251 (.A(net63));
 sg13g2_antennanp ANTENNA_1252 (.A(net67));
 sg13g2_antennanp ANTENNA_1253 (.A(net67));
 sg13g2_antennanp ANTENNA_1254 (.A(net67));
 sg13g2_antennanp ANTENNA_1255 (.A(net67));
 sg13g2_antennanp ANTENNA_1256 (.A(net67));
 sg13g2_antennanp ANTENNA_1257 (.A(net67));
 sg13g2_antennanp ANTENNA_1258 (.A(net67));
 sg13g2_antennanp ANTENNA_1259 (.A(net67));
 sg13g2_antennanp ANTENNA_1260 (.A(net67));
 sg13g2_antennanp ANTENNA_1261 (.A(net67));
 sg13g2_antennanp ANTENNA_1262 (.A(net67));
 sg13g2_antennanp ANTENNA_1263 (.A(net77));
 sg13g2_antennanp ANTENNA_1264 (.A(net77));
 sg13g2_antennanp ANTENNA_1265 (.A(net77));
 sg13g2_antennanp ANTENNA_1266 (.A(net77));
 sg13g2_antennanp ANTENNA_1267 (.A(net77));
 sg13g2_antennanp ANTENNA_1268 (.A(net77));
 sg13g2_antennanp ANTENNA_1269 (.A(net77));
 sg13g2_antennanp ANTENNA_1270 (.A(net77));
 sg13g2_antennanp ANTENNA_1271 (.A(net77));
 sg13g2_antennanp ANTENNA_1272 (.A(net91));
 sg13g2_antennanp ANTENNA_1273 (.A(net91));
 sg13g2_antennanp ANTENNA_1274 (.A(net91));
 sg13g2_antennanp ANTENNA_1275 (.A(net91));
 sg13g2_antennanp ANTENNA_1276 (.A(net91));
 sg13g2_antennanp ANTENNA_1277 (.A(net91));
 sg13g2_antennanp ANTENNA_1278 (.A(net91));
 sg13g2_antennanp ANTENNA_1279 (.A(net91));
 sg13g2_antennanp ANTENNA_1280 (.A(net91));
 sg13g2_antennanp ANTENNA_1281 (.A(net146));
 sg13g2_antennanp ANTENNA_1282 (.A(net146));
 sg13g2_antennanp ANTENNA_1283 (.A(net146));
 sg13g2_antennanp ANTENNA_1284 (.A(net146));
 sg13g2_antennanp ANTENNA_1285 (.A(net146));
 sg13g2_antennanp ANTENNA_1286 (.A(net146));
 sg13g2_antennanp ANTENNA_1287 (.A(net146));
 sg13g2_antennanp ANTENNA_1288 (.A(net146));
 sg13g2_antennanp ANTENNA_1289 (.A(net146));
 sg13g2_antennanp ANTENNA_1290 (.A(net155));
 sg13g2_antennanp ANTENNA_1291 (.A(net155));
 sg13g2_antennanp ANTENNA_1292 (.A(net155));
 sg13g2_antennanp ANTENNA_1293 (.A(net155));
 sg13g2_antennanp ANTENNA_1294 (.A(net155));
 sg13g2_antennanp ANTENNA_1295 (.A(net155));
 sg13g2_antennanp ANTENNA_1296 (.A(net155));
 sg13g2_antennanp ANTENNA_1297 (.A(net155));
 sg13g2_antennanp ANTENNA_1298 (.A(net155));
 sg13g2_antennanp ANTENNA_1299 (.A(net155));
 sg13g2_antennanp ANTENNA_1300 (.A(net155));
 sg13g2_antennanp ANTENNA_1301 (.A(net191));
 sg13g2_antennanp ANTENNA_1302 (.A(net191));
 sg13g2_antennanp ANTENNA_1303 (.A(net191));
 sg13g2_antennanp ANTENNA_1304 (.A(net191));
 sg13g2_antennanp ANTENNA_1305 (.A(net191));
 sg13g2_antennanp ANTENNA_1306 (.A(net191));
 sg13g2_antennanp ANTENNA_1307 (.A(net191));
 sg13g2_antennanp ANTENNA_1308 (.A(net191));
 sg13g2_antennanp ANTENNA_1309 (.A(net194));
 sg13g2_antennanp ANTENNA_1310 (.A(net194));
 sg13g2_antennanp ANTENNA_1311 (.A(net194));
 sg13g2_antennanp ANTENNA_1312 (.A(net194));
 sg13g2_antennanp ANTENNA_1313 (.A(net194));
 sg13g2_antennanp ANTENNA_1314 (.A(net194));
 sg13g2_antennanp ANTENNA_1315 (.A(net194));
 sg13g2_antennanp ANTENNA_1316 (.A(net194));
 sg13g2_antennanp ANTENNA_1317 (.A(net292));
 sg13g2_antennanp ANTENNA_1318 (.A(net292));
 sg13g2_antennanp ANTENNA_1319 (.A(net292));
 sg13g2_antennanp ANTENNA_1320 (.A(net292));
 sg13g2_antennanp ANTENNA_1321 (.A(net292));
 sg13g2_antennanp ANTENNA_1322 (.A(net292));
 sg13g2_antennanp ANTENNA_1323 (.A(net292));
 sg13g2_antennanp ANTENNA_1324 (.A(net292));
 sg13g2_antennanp ANTENNA_1325 (.A(net292));
 sg13g2_antennanp ANTENNA_1326 (.A(net308));
 sg13g2_antennanp ANTENNA_1327 (.A(net308));
 sg13g2_antennanp ANTENNA_1328 (.A(net308));
 sg13g2_antennanp ANTENNA_1329 (.A(net308));
 sg13g2_antennanp ANTENNA_1330 (.A(net308));
 sg13g2_antennanp ANTENNA_1331 (.A(net308));
 sg13g2_antennanp ANTENNA_1332 (.A(net308));
 sg13g2_antennanp ANTENNA_1333 (.A(net308));
 sg13g2_antennanp ANTENNA_1334 (.A(net317));
 sg13g2_antennanp ANTENNA_1335 (.A(net317));
 sg13g2_antennanp ANTENNA_1336 (.A(net317));
 sg13g2_antennanp ANTENNA_1337 (.A(net317));
 sg13g2_antennanp ANTENNA_1338 (.A(net317));
 sg13g2_antennanp ANTENNA_1339 (.A(net317));
 sg13g2_antennanp ANTENNA_1340 (.A(net317));
 sg13g2_antennanp ANTENNA_1341 (.A(net317));
 sg13g2_antennanp ANTENNA_1342 (.A(net317));
 sg13g2_antennanp ANTENNA_1343 (.A(net340));
 sg13g2_antennanp ANTENNA_1344 (.A(net340));
 sg13g2_antennanp ANTENNA_1345 (.A(net340));
 sg13g2_antennanp ANTENNA_1346 (.A(net340));
 sg13g2_antennanp ANTENNA_1347 (.A(net340));
 sg13g2_antennanp ANTENNA_1348 (.A(net340));
 sg13g2_antennanp ANTENNA_1349 (.A(net340));
 sg13g2_antennanp ANTENNA_1350 (.A(net340));
 sg13g2_antennanp ANTENNA_1351 (.A(net340));
 sg13g2_antennanp ANTENNA_1352 (.A(net369));
 sg13g2_antennanp ANTENNA_1353 (.A(net369));
 sg13g2_antennanp ANTENNA_1354 (.A(net369));
 sg13g2_antennanp ANTENNA_1355 (.A(net369));
 sg13g2_antennanp ANTENNA_1356 (.A(net369));
 sg13g2_antennanp ANTENNA_1357 (.A(net369));
 sg13g2_antennanp ANTENNA_1358 (.A(net369));
 sg13g2_antennanp ANTENNA_1359 (.A(net369));
 sg13g2_antennanp ANTENNA_1360 (.A(net378));
 sg13g2_antennanp ANTENNA_1361 (.A(net378));
 sg13g2_antennanp ANTENNA_1362 (.A(net378));
 sg13g2_antennanp ANTENNA_1363 (.A(net378));
 sg13g2_antennanp ANTENNA_1364 (.A(net378));
 sg13g2_antennanp ANTENNA_1365 (.A(net378));
 sg13g2_antennanp ANTENNA_1366 (.A(net378));
 sg13g2_antennanp ANTENNA_1367 (.A(net378));
 sg13g2_antennanp ANTENNA_1368 (.A(net378));
 sg13g2_antennanp ANTENNA_1369 (.A(net378));
 sg13g2_antennanp ANTENNA_1370 (.A(net378));
 sg13g2_antennanp ANTENNA_1371 (.A(net378));
 sg13g2_antennanp ANTENNA_1372 (.A(net384));
 sg13g2_antennanp ANTENNA_1373 (.A(net384));
 sg13g2_antennanp ANTENNA_1374 (.A(net384));
 sg13g2_antennanp ANTENNA_1375 (.A(net384));
 sg13g2_antennanp ANTENNA_1376 (.A(net384));
 sg13g2_antennanp ANTENNA_1377 (.A(net384));
 sg13g2_antennanp ANTENNA_1378 (.A(net384));
 sg13g2_antennanp ANTENNA_1379 (.A(net384));
 sg13g2_antennanp ANTENNA_1380 (.A(net384));
 sg13g2_antennanp ANTENNA_1381 (.A(net384));
 sg13g2_antennanp ANTENNA_1382 (.A(net384));
 sg13g2_antennanp ANTENNA_1383 (.A(net384));
 sg13g2_antennanp ANTENNA_1384 (.A(net412));
 sg13g2_antennanp ANTENNA_1385 (.A(net412));
 sg13g2_antennanp ANTENNA_1386 (.A(net412));
 sg13g2_antennanp ANTENNA_1387 (.A(net412));
 sg13g2_antennanp ANTENNA_1388 (.A(net412));
 sg13g2_antennanp ANTENNA_1389 (.A(net412));
 sg13g2_antennanp ANTENNA_1390 (.A(net412));
 sg13g2_antennanp ANTENNA_1391 (.A(net412));
 sg13g2_antennanp ANTENNA_1392 (.A(net435));
 sg13g2_antennanp ANTENNA_1393 (.A(net435));
 sg13g2_antennanp ANTENNA_1394 (.A(net435));
 sg13g2_antennanp ANTENNA_1395 (.A(net435));
 sg13g2_antennanp ANTENNA_1396 (.A(net435));
 sg13g2_antennanp ANTENNA_1397 (.A(net435));
 sg13g2_antennanp ANTENNA_1398 (.A(net435));
 sg13g2_antennanp ANTENNA_1399 (.A(net435));
 sg13g2_antennanp ANTENNA_1400 (.A(net436));
 sg13g2_antennanp ANTENNA_1401 (.A(net436));
 sg13g2_antennanp ANTENNA_1402 (.A(net436));
 sg13g2_antennanp ANTENNA_1403 (.A(net436));
 sg13g2_antennanp ANTENNA_1404 (.A(net436));
 sg13g2_antennanp ANTENNA_1405 (.A(net436));
 sg13g2_antennanp ANTENNA_1406 (.A(net436));
 sg13g2_antennanp ANTENNA_1407 (.A(net436));
 sg13g2_antennanp ANTENNA_1408 (.A(net498));
 sg13g2_antennanp ANTENNA_1409 (.A(net498));
 sg13g2_antennanp ANTENNA_1410 (.A(net498));
 sg13g2_antennanp ANTENNA_1411 (.A(net498));
 sg13g2_antennanp ANTENNA_1412 (.A(net498));
 sg13g2_antennanp ANTENNA_1413 (.A(net498));
 sg13g2_antennanp ANTENNA_1414 (.A(net498));
 sg13g2_antennanp ANTENNA_1415 (.A(net498));
 sg13g2_antennanp ANTENNA_1416 (.A(net498));
 sg13g2_antennanp ANTENNA_1417 (.A(net525));
 sg13g2_antennanp ANTENNA_1418 (.A(net525));
 sg13g2_antennanp ANTENNA_1419 (.A(net525));
 sg13g2_antennanp ANTENNA_1420 (.A(net525));
 sg13g2_antennanp ANTENNA_1421 (.A(net525));
 sg13g2_antennanp ANTENNA_1422 (.A(net525));
 sg13g2_antennanp ANTENNA_1423 (.A(net525));
 sg13g2_antennanp ANTENNA_1424 (.A(net525));
 sg13g2_antennanp ANTENNA_1425 (.A(net525));
 sg13g2_antennanp ANTENNA_1426 (.A(net525));
 sg13g2_antennanp ANTENNA_1427 (.A(net1207));
 sg13g2_antennanp ANTENNA_1428 (.A(net1207));
 sg13g2_antennanp ANTENNA_1429 (.A(net1207));
 sg13g2_antennanp ANTENNA_1430 (.A(net1207));
 sg13g2_antennanp ANTENNA_1431 (.A(net1207));
 sg13g2_antennanp ANTENNA_1432 (.A(net1207));
 sg13g2_antennanp ANTENNA_1433 (.A(net1207));
 sg13g2_antennanp ANTENNA_1434 (.A(net1430));
 sg13g2_antennanp ANTENNA_1435 (.A(net1430));
 sg13g2_antennanp ANTENNA_1436 (.A(net1430));
 sg13g2_antennanp ANTENNA_1437 (.A(net1430));
 sg13g2_antennanp ANTENNA_1438 (.A(net1430));
 sg13g2_antennanp ANTENNA_1439 (.A(net1430));
 sg13g2_antennanp ANTENNA_1440 (.A(net1430));
 sg13g2_antennanp ANTENNA_1441 (.A(_00366_));
 sg13g2_antennanp ANTENNA_1442 (.A(_00366_));
 sg13g2_antennanp ANTENNA_1443 (.A(_00394_));
 sg13g2_antennanp ANTENNA_1444 (.A(_00394_));
 sg13g2_antennanp ANTENNA_1445 (.A(_00406_));
 sg13g2_antennanp ANTENNA_1446 (.A(_00406_));
 sg13g2_antennanp ANTENNA_1447 (.A(_00408_));
 sg13g2_antennanp ANTENNA_1448 (.A(_00411_));
 sg13g2_antennanp ANTENNA_1449 (.A(_00412_));
 sg13g2_antennanp ANTENNA_1450 (.A(_00413_));
 sg13g2_antennanp ANTENNA_1451 (.A(_00413_));
 sg13g2_antennanp ANTENNA_1452 (.A(_00417_));
 sg13g2_antennanp ANTENNA_1453 (.A(_03004_));
 sg13g2_antennanp ANTENNA_1454 (.A(_03004_));
 sg13g2_antennanp ANTENNA_1455 (.A(_03004_));
 sg13g2_antennanp ANTENNA_1456 (.A(_03063_));
 sg13g2_antennanp ANTENNA_1457 (.A(_03063_));
 sg13g2_antennanp ANTENNA_1458 (.A(_03063_));
 sg13g2_antennanp ANTENNA_1459 (.A(_03063_));
 sg13g2_antennanp ANTENNA_1460 (.A(_03145_));
 sg13g2_antennanp ANTENNA_1461 (.A(_03451_));
 sg13g2_antennanp ANTENNA_1462 (.A(_03451_));
 sg13g2_antennanp ANTENNA_1463 (.A(_03451_));
 sg13g2_antennanp ANTENNA_1464 (.A(_03451_));
 sg13g2_antennanp ANTENNA_1465 (.A(_03451_));
 sg13g2_antennanp ANTENNA_1466 (.A(_03451_));
 sg13g2_antennanp ANTENNA_1467 (.A(_04085_));
 sg13g2_antennanp ANTENNA_1468 (.A(_04085_));
 sg13g2_antennanp ANTENNA_1469 (.A(_04085_));
 sg13g2_antennanp ANTENNA_1470 (.A(_04086_));
 sg13g2_antennanp ANTENNA_1471 (.A(_04086_));
 sg13g2_antennanp ANTENNA_1472 (.A(_04086_));
 sg13g2_antennanp ANTENNA_1473 (.A(_04107_));
 sg13g2_antennanp ANTENNA_1474 (.A(_04743_));
 sg13g2_antennanp ANTENNA_1475 (.A(_04743_));
 sg13g2_antennanp ANTENNA_1476 (.A(_05412_));
 sg13g2_antennanp ANTENNA_1477 (.A(_05412_));
 sg13g2_antennanp ANTENNA_1478 (.A(_05412_));
 sg13g2_antennanp ANTENNA_1479 (.A(_05412_));
 sg13g2_antennanp ANTENNA_1480 (.A(_05412_));
 sg13g2_antennanp ANTENNA_1481 (.A(_05412_));
 sg13g2_antennanp ANTENNA_1482 (.A(_05436_));
 sg13g2_antennanp ANTENNA_1483 (.A(_05436_));
 sg13g2_antennanp ANTENNA_1484 (.A(_05436_));
 sg13g2_antennanp ANTENNA_1485 (.A(_05436_));
 sg13g2_antennanp ANTENNA_1486 (.A(_05495_));
 sg13g2_antennanp ANTENNA_1487 (.A(_05495_));
 sg13g2_antennanp ANTENNA_1488 (.A(_05495_));
 sg13g2_antennanp ANTENNA_1489 (.A(_05592_));
 sg13g2_antennanp ANTENNA_1490 (.A(_05621_));
 sg13g2_antennanp ANTENNA_1491 (.A(_05631_));
 sg13g2_antennanp ANTENNA_1492 (.A(_05639_));
 sg13g2_antennanp ANTENNA_1493 (.A(_05648_));
 sg13g2_antennanp ANTENNA_1494 (.A(_05648_));
 sg13g2_antennanp ANTENNA_1495 (.A(_05648_));
 sg13g2_antennanp ANTENNA_1496 (.A(_05689_));
 sg13g2_antennanp ANTENNA_1497 (.A(_05719_));
 sg13g2_antennanp ANTENNA_1498 (.A(_05719_));
 sg13g2_antennanp ANTENNA_1499 (.A(_05719_));
 sg13g2_antennanp ANTENNA_1500 (.A(_05719_));
 sg13g2_antennanp ANTENNA_1501 (.A(_05719_));
 sg13g2_antennanp ANTENNA_1502 (.A(_05729_));
 sg13g2_antennanp ANTENNA_1503 (.A(_05729_));
 sg13g2_antennanp ANTENNA_1504 (.A(_05729_));
 sg13g2_antennanp ANTENNA_1505 (.A(_05739_));
 sg13g2_antennanp ANTENNA_1506 (.A(_05773_));
 sg13g2_antennanp ANTENNA_1507 (.A(_05781_));
 sg13g2_antennanp ANTENNA_1508 (.A(_05785_));
 sg13g2_antennanp ANTENNA_1509 (.A(_05807_));
 sg13g2_antennanp ANTENNA_1510 (.A(_05825_));
 sg13g2_antennanp ANTENNA_1511 (.A(_05825_));
 sg13g2_antennanp ANTENNA_1512 (.A(_05825_));
 sg13g2_antennanp ANTENNA_1513 (.A(_05829_));
 sg13g2_antennanp ANTENNA_1514 (.A(_05858_));
 sg13g2_antennanp ANTENNA_1515 (.A(_05866_));
 sg13g2_antennanp ANTENNA_1516 (.A(_05877_));
 sg13g2_antennanp ANTENNA_1517 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1518 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1519 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1520 (.A(_05942_));
 sg13g2_antennanp ANTENNA_1521 (.A(_05960_));
 sg13g2_antennanp ANTENNA_1522 (.A(_05960_));
 sg13g2_antennanp ANTENNA_1523 (.A(_05960_));
 sg13g2_antennanp ANTENNA_1524 (.A(_05977_));
 sg13g2_antennanp ANTENNA_1525 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1526 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1527 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1528 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1529 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1530 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1531 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1532 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1533 (.A(_06027_));
 sg13g2_antennanp ANTENNA_1534 (.A(_06038_));
 sg13g2_antennanp ANTENNA_1535 (.A(_06045_));
 sg13g2_antennanp ANTENNA_1536 (.A(_06053_));
 sg13g2_antennanp ANTENNA_1537 (.A(_06065_));
 sg13g2_antennanp ANTENNA_1538 (.A(_06065_));
 sg13g2_antennanp ANTENNA_1539 (.A(_06065_));
 sg13g2_antennanp ANTENNA_1540 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1541 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1542 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1543 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1544 (.A(_06152_));
 sg13g2_antennanp ANTENNA_1545 (.A(_06163_));
 sg13g2_antennanp ANTENNA_1546 (.A(_06163_));
 sg13g2_antennanp ANTENNA_1547 (.A(_06163_));
 sg13g2_antennanp ANTENNA_1548 (.A(_06183_));
 sg13g2_antennanp ANTENNA_1549 (.A(_06183_));
 sg13g2_antennanp ANTENNA_1550 (.A(_06183_));
 sg13g2_antennanp ANTENNA_1551 (.A(_06183_));
 sg13g2_antennanp ANTENNA_1552 (.A(_06195_));
 sg13g2_antennanp ANTENNA_1553 (.A(_06216_));
 sg13g2_antennanp ANTENNA_1554 (.A(_06236_));
 sg13g2_antennanp ANTENNA_1555 (.A(_06247_));
 sg13g2_antennanp ANTENNA_1556 (.A(_06259_));
 sg13g2_antennanp ANTENNA_1557 (.A(_06285_));
 sg13g2_antennanp ANTENNA_1558 (.A(_06303_));
 sg13g2_antennanp ANTENNA_1559 (.A(_06318_));
 sg13g2_antennanp ANTENNA_1560 (.A(_06337_));
 sg13g2_antennanp ANTENNA_1561 (.A(_06350_));
 sg13g2_antennanp ANTENNA_1562 (.A(_06355_));
 sg13g2_antennanp ANTENNA_1563 (.A(_06370_));
 sg13g2_antennanp ANTENNA_1564 (.A(_06380_));
 sg13g2_antennanp ANTENNA_1565 (.A(_06385_));
 sg13g2_antennanp ANTENNA_1566 (.A(_06391_));
 sg13g2_antennanp ANTENNA_1567 (.A(_06423_));
 sg13g2_antennanp ANTENNA_1568 (.A(_06435_));
 sg13g2_antennanp ANTENNA_1569 (.A(_06438_));
 sg13g2_antennanp ANTENNA_1570 (.A(_06464_));
 sg13g2_antennanp ANTENNA_1571 (.A(_06475_));
 sg13g2_antennanp ANTENNA_1572 (.A(_06525_));
 sg13g2_antennanp ANTENNA_1573 (.A(_06530_));
 sg13g2_antennanp ANTENNA_1574 (.A(_06532_));
 sg13g2_antennanp ANTENNA_1575 (.A(_06582_));
 sg13g2_antennanp ANTENNA_1576 (.A(_06605_));
 sg13g2_antennanp ANTENNA_1577 (.A(_06653_));
 sg13g2_antennanp ANTENNA_1578 (.A(_06660_));
 sg13g2_antennanp ANTENNA_1579 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1580 (.A(_06671_));
 sg13g2_antennanp ANTENNA_1581 (.A(_06697_));
 sg13g2_antennanp ANTENNA_1582 (.A(_06701_));
 sg13g2_antennanp ANTENNA_1583 (.A(_06703_));
 sg13g2_antennanp ANTENNA_1584 (.A(_06751_));
 sg13g2_antennanp ANTENNA_1585 (.A(_06772_));
 sg13g2_antennanp ANTENNA_1586 (.A(_06813_));
 sg13g2_antennanp ANTENNA_1587 (.A(_06815_));
 sg13g2_antennanp ANTENNA_1588 (.A(_06816_));
 sg13g2_antennanp ANTENNA_1589 (.A(_06829_));
 sg13g2_antennanp ANTENNA_1590 (.A(_06850_));
 sg13g2_antennanp ANTENNA_1591 (.A(_06854_));
 sg13g2_antennanp ANTENNA_1592 (.A(_06869_));
 sg13g2_antennanp ANTENNA_1593 (.A(_06870_));
 sg13g2_antennanp ANTENNA_1594 (.A(_06875_));
 sg13g2_antennanp ANTENNA_1595 (.A(_06881_));
 sg13g2_antennanp ANTENNA_1596 (.A(_06901_));
 sg13g2_antennanp ANTENNA_1597 (.A(_06921_));
 sg13g2_antennanp ANTENNA_1598 (.A(_06932_));
 sg13g2_antennanp ANTENNA_1599 (.A(_06936_));
 sg13g2_antennanp ANTENNA_1600 (.A(_06936_));
 sg13g2_antennanp ANTENNA_1601 (.A(_06959_));
 sg13g2_antennanp ANTENNA_1602 (.A(_06993_));
 sg13g2_antennanp ANTENNA_1603 (.A(_06998_));
 sg13g2_antennanp ANTENNA_1604 (.A(_07008_));
 sg13g2_antennanp ANTENNA_1605 (.A(_07035_));
 sg13g2_antennanp ANTENNA_1606 (.A(_07036_));
 sg13g2_antennanp ANTENNA_1607 (.A(_07047_));
 sg13g2_antennanp ANTENNA_1608 (.A(_07060_));
 sg13g2_antennanp ANTENNA_1609 (.A(_07069_));
 sg13g2_antennanp ANTENNA_1610 (.A(_07074_));
 sg13g2_antennanp ANTENNA_1611 (.A(_07080_));
 sg13g2_antennanp ANTENNA_1612 (.A(_07108_));
 sg13g2_antennanp ANTENNA_1613 (.A(_07139_));
 sg13g2_antennanp ANTENNA_1614 (.A(_07146_));
 sg13g2_antennanp ANTENNA_1615 (.A(_07191_));
 sg13g2_antennanp ANTENNA_1616 (.A(_07212_));
 sg13g2_antennanp ANTENNA_1617 (.A(_07217_));
 sg13g2_antennanp ANTENNA_1618 (.A(_07254_));
 sg13g2_antennanp ANTENNA_1619 (.A(_07282_));
 sg13g2_antennanp ANTENNA_1620 (.A(_07284_));
 sg13g2_antennanp ANTENNA_1621 (.A(_07288_));
 sg13g2_antennanp ANTENNA_1622 (.A(_07288_));
 sg13g2_antennanp ANTENNA_1623 (.A(_07302_));
 sg13g2_antennanp ANTENNA_1624 (.A(_07312_));
 sg13g2_antennanp ANTENNA_1625 (.A(_07363_));
 sg13g2_antennanp ANTENNA_1626 (.A(_07375_));
 sg13g2_antennanp ANTENNA_1627 (.A(_07403_));
 sg13g2_antennanp ANTENNA_1628 (.A(_07420_));
 sg13g2_antennanp ANTENNA_1629 (.A(_07420_));
 sg13g2_antennanp ANTENNA_1630 (.A(_07428_));
 sg13g2_antennanp ANTENNA_1631 (.A(_07460_));
 sg13g2_antennanp ANTENNA_1632 (.A(_07460_));
 sg13g2_antennanp ANTENNA_1633 (.A(_07460_));
 sg13g2_antennanp ANTENNA_1634 (.A(_07460_));
 sg13g2_antennanp ANTENNA_1635 (.A(_07460_));
 sg13g2_antennanp ANTENNA_1636 (.A(_07460_));
 sg13g2_antennanp ANTENNA_1637 (.A(_07491_));
 sg13g2_antennanp ANTENNA_1638 (.A(_07491_));
 sg13g2_antennanp ANTENNA_1639 (.A(_07491_));
 sg13g2_antennanp ANTENNA_1640 (.A(_07491_));
 sg13g2_antennanp ANTENNA_1641 (.A(_07491_));
 sg13g2_antennanp ANTENNA_1642 (.A(_07491_));
 sg13g2_antennanp ANTENNA_1643 (.A(_07496_));
 sg13g2_antennanp ANTENNA_1644 (.A(_07496_));
 sg13g2_antennanp ANTENNA_1645 (.A(_07496_));
 sg13g2_antennanp ANTENNA_1646 (.A(_07496_));
 sg13g2_antennanp ANTENNA_1647 (.A(_07609_));
 sg13g2_antennanp ANTENNA_1648 (.A(_07622_));
 sg13g2_antennanp ANTENNA_1649 (.A(_07636_));
 sg13g2_antennanp ANTENNA_1650 (.A(_07704_));
 sg13g2_antennanp ANTENNA_1651 (.A(_07704_));
 sg13g2_antennanp ANTENNA_1652 (.A(_07730_));
 sg13g2_antennanp ANTENNA_1653 (.A(_07758_));
 sg13g2_antennanp ANTENNA_1654 (.A(_07822_));
 sg13g2_antennanp ANTENNA_1655 (.A(_07835_));
 sg13g2_antennanp ANTENNA_1656 (.A(_07835_));
 sg13g2_antennanp ANTENNA_1657 (.A(_07914_));
 sg13g2_antennanp ANTENNA_1658 (.A(_07926_));
 sg13g2_antennanp ANTENNA_1659 (.A(_07939_));
 sg13g2_antennanp ANTENNA_1660 (.A(_07939_));
 sg13g2_antennanp ANTENNA_1661 (.A(_07952_));
 sg13g2_antennanp ANTENNA_1662 (.A(_08169_));
 sg13g2_antennanp ANTENNA_1663 (.A(_08169_));
 sg13g2_antennanp ANTENNA_1664 (.A(_09280_));
 sg13g2_antennanp ANTENNA_1665 (.A(_09280_));
 sg13g2_antennanp ANTENNA_1666 (.A(_09280_));
 sg13g2_antennanp ANTENNA_1667 (.A(_09280_));
 sg13g2_antennanp ANTENNA_1668 (.A(_09280_));
 sg13g2_antennanp ANTENNA_1669 (.A(_09724_));
 sg13g2_antennanp ANTENNA_1670 (.A(_09825_));
 sg13g2_antennanp ANTENNA_1671 (.A(_09825_));
 sg13g2_antennanp ANTENNA_1672 (.A(_09825_));
 sg13g2_antennanp ANTENNA_1673 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1674 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1675 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1676 (.A(_10247_));
 sg13g2_antennanp ANTENNA_1677 (.A(_10247_));
 sg13g2_antennanp ANTENNA_1678 (.A(_10247_));
 sg13g2_antennanp ANTENNA_1679 (.A(_10518_));
 sg13g2_antennanp ANTENNA_1680 (.A(_10604_));
 sg13g2_antennanp ANTENNA_1681 (.A(_10604_));
 sg13g2_antennanp ANTENNA_1682 (.A(_10604_));
 sg13g2_antennanp ANTENNA_1683 (.A(_10604_));
 sg13g2_antennanp ANTENNA_1684 (.A(_10617_));
 sg13g2_antennanp ANTENNA_1685 (.A(_10952_));
 sg13g2_antennanp ANTENNA_1686 (.A(_10963_));
 sg13g2_antennanp ANTENNA_1687 (.A(_11000_));
 sg13g2_antennanp ANTENNA_1688 (.A(_11000_));
 sg13g2_antennanp ANTENNA_1689 (.A(_11000_));
 sg13g2_antennanp ANTENNA_1690 (.A(_11060_));
 sg13g2_antennanp ANTENNA_1691 (.A(_11060_));
 sg13g2_antennanp ANTENNA_1692 (.A(_11060_));
 sg13g2_antennanp ANTENNA_1693 (.A(_11060_));
 sg13g2_antennanp ANTENNA_1694 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1695 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1696 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1697 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1698 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1699 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1700 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1701 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1702 (.A(_11243_));
 sg13g2_antennanp ANTENNA_1703 (.A(\top_ihp.oisc.op_a[22] ));
 sg13g2_antennanp ANTENNA_1704 (.A(\top_ihp.oisc.op_a[27] ));
 sg13g2_antennanp ANTENNA_1705 (.A(\top_ihp.oisc.op_a[6] ));
 sg13g2_antennanp ANTENNA_1706 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_1707 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_1708 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_1709 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_1710 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_1711 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_1712 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_1713 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_1714 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_1715 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_1716 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_1717 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_1718 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_1719 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_1720 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_1721 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_1722 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_1723 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_1724 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_1725 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_1726 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_1727 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_1728 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_1729 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_1730 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_1731 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_1732 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_1733 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_1734 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_1735 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_1736 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_1737 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_1738 (.A(\top_ihp.tx ));
 sg13g2_antennanp ANTENNA_1739 (.A(net1));
 sg13g2_antennanp ANTENNA_1740 (.A(net1));
 sg13g2_antennanp ANTENNA_1741 (.A(net1));
 sg13g2_antennanp ANTENNA_1742 (.A(net5));
 sg13g2_antennanp ANTENNA_1743 (.A(net10));
 sg13g2_antennanp ANTENNA_1744 (.A(net67));
 sg13g2_antennanp ANTENNA_1745 (.A(net67));
 sg13g2_antennanp ANTENNA_1746 (.A(net67));
 sg13g2_antennanp ANTENNA_1747 (.A(net67));
 sg13g2_antennanp ANTENNA_1748 (.A(net67));
 sg13g2_antennanp ANTENNA_1749 (.A(net67));
 sg13g2_antennanp ANTENNA_1750 (.A(net67));
 sg13g2_antennanp ANTENNA_1751 (.A(net67));
 sg13g2_antennanp ANTENNA_1752 (.A(net67));
 sg13g2_antennanp ANTENNA_1753 (.A(net67));
 sg13g2_antennanp ANTENNA_1754 (.A(net67));
 sg13g2_antennanp ANTENNA_1755 (.A(net67));
 sg13g2_antennanp ANTENNA_1756 (.A(net67));
 sg13g2_antennanp ANTENNA_1757 (.A(net67));
 sg13g2_antennanp ANTENNA_1758 (.A(net67));
 sg13g2_antennanp ANTENNA_1759 (.A(net67));
 sg13g2_antennanp ANTENNA_1760 (.A(net67));
 sg13g2_antennanp ANTENNA_1761 (.A(net67));
 sg13g2_antennanp ANTENNA_1762 (.A(net77));
 sg13g2_antennanp ANTENNA_1763 (.A(net77));
 sg13g2_antennanp ANTENNA_1764 (.A(net77));
 sg13g2_antennanp ANTENNA_1765 (.A(net77));
 sg13g2_antennanp ANTENNA_1766 (.A(net77));
 sg13g2_antennanp ANTENNA_1767 (.A(net77));
 sg13g2_antennanp ANTENNA_1768 (.A(net77));
 sg13g2_antennanp ANTENNA_1769 (.A(net77));
 sg13g2_antennanp ANTENNA_1770 (.A(net77));
 sg13g2_antennanp ANTENNA_1771 (.A(net91));
 sg13g2_antennanp ANTENNA_1772 (.A(net91));
 sg13g2_antennanp ANTENNA_1773 (.A(net91));
 sg13g2_antennanp ANTENNA_1774 (.A(net91));
 sg13g2_antennanp ANTENNA_1775 (.A(net91));
 sg13g2_antennanp ANTENNA_1776 (.A(net91));
 sg13g2_antennanp ANTENNA_1777 (.A(net91));
 sg13g2_antennanp ANTENNA_1778 (.A(net91));
 sg13g2_antennanp ANTENNA_1779 (.A(net91));
 sg13g2_antennanp ANTENNA_1780 (.A(net146));
 sg13g2_antennanp ANTENNA_1781 (.A(net146));
 sg13g2_antennanp ANTENNA_1782 (.A(net146));
 sg13g2_antennanp ANTENNA_1783 (.A(net146));
 sg13g2_antennanp ANTENNA_1784 (.A(net146));
 sg13g2_antennanp ANTENNA_1785 (.A(net146));
 sg13g2_antennanp ANTENNA_1786 (.A(net146));
 sg13g2_antennanp ANTENNA_1787 (.A(net146));
 sg13g2_antennanp ANTENNA_1788 (.A(net146));
 sg13g2_antennanp ANTENNA_1789 (.A(net146));
 sg13g2_antennanp ANTENNA_1790 (.A(net146));
 sg13g2_antennanp ANTENNA_1791 (.A(net146));
 sg13g2_antennanp ANTENNA_1792 (.A(net155));
 sg13g2_antennanp ANTENNA_1793 (.A(net155));
 sg13g2_antennanp ANTENNA_1794 (.A(net155));
 sg13g2_antennanp ANTENNA_1795 (.A(net155));
 sg13g2_antennanp ANTENNA_1796 (.A(net155));
 sg13g2_antennanp ANTENNA_1797 (.A(net155));
 sg13g2_antennanp ANTENNA_1798 (.A(net155));
 sg13g2_antennanp ANTENNA_1799 (.A(net155));
 sg13g2_antennanp ANTENNA_1800 (.A(net155));
 sg13g2_antennanp ANTENNA_1801 (.A(net155));
 sg13g2_antennanp ANTENNA_1802 (.A(net155));
 sg13g2_antennanp ANTENNA_1803 (.A(net292));
 sg13g2_antennanp ANTENNA_1804 (.A(net292));
 sg13g2_antennanp ANTENNA_1805 (.A(net292));
 sg13g2_antennanp ANTENNA_1806 (.A(net292));
 sg13g2_antennanp ANTENNA_1807 (.A(net292));
 sg13g2_antennanp ANTENNA_1808 (.A(net292));
 sg13g2_antennanp ANTENNA_1809 (.A(net292));
 sg13g2_antennanp ANTENNA_1810 (.A(net292));
 sg13g2_antennanp ANTENNA_1811 (.A(net292));
 sg13g2_antennanp ANTENNA_1812 (.A(net308));
 sg13g2_antennanp ANTENNA_1813 (.A(net308));
 sg13g2_antennanp ANTENNA_1814 (.A(net308));
 sg13g2_antennanp ANTENNA_1815 (.A(net308));
 sg13g2_antennanp ANTENNA_1816 (.A(net308));
 sg13g2_antennanp ANTENNA_1817 (.A(net308));
 sg13g2_antennanp ANTENNA_1818 (.A(net308));
 sg13g2_antennanp ANTENNA_1819 (.A(net308));
 sg13g2_antennanp ANTENNA_1820 (.A(net317));
 sg13g2_antennanp ANTENNA_1821 (.A(net317));
 sg13g2_antennanp ANTENNA_1822 (.A(net317));
 sg13g2_antennanp ANTENNA_1823 (.A(net317));
 sg13g2_antennanp ANTENNA_1824 (.A(net317));
 sg13g2_antennanp ANTENNA_1825 (.A(net317));
 sg13g2_antennanp ANTENNA_1826 (.A(net317));
 sg13g2_antennanp ANTENNA_1827 (.A(net317));
 sg13g2_antennanp ANTENNA_1828 (.A(net317));
 sg13g2_antennanp ANTENNA_1829 (.A(net397));
 sg13g2_antennanp ANTENNA_1830 (.A(net397));
 sg13g2_antennanp ANTENNA_1831 (.A(net397));
 sg13g2_antennanp ANTENNA_1832 (.A(net397));
 sg13g2_antennanp ANTENNA_1833 (.A(net397));
 sg13g2_antennanp ANTENNA_1834 (.A(net397));
 sg13g2_antennanp ANTENNA_1835 (.A(net397));
 sg13g2_antennanp ANTENNA_1836 (.A(net397));
 sg13g2_antennanp ANTENNA_1837 (.A(net397));
 sg13g2_antennanp ANTENNA_1838 (.A(net412));
 sg13g2_antennanp ANTENNA_1839 (.A(net412));
 sg13g2_antennanp ANTENNA_1840 (.A(net412));
 sg13g2_antennanp ANTENNA_1841 (.A(net412));
 sg13g2_antennanp ANTENNA_1842 (.A(net412));
 sg13g2_antennanp ANTENNA_1843 (.A(net412));
 sg13g2_antennanp ANTENNA_1844 (.A(net412));
 sg13g2_antennanp ANTENNA_1845 (.A(net412));
 sg13g2_antennanp ANTENNA_1846 (.A(net436));
 sg13g2_antennanp ANTENNA_1847 (.A(net436));
 sg13g2_antennanp ANTENNA_1848 (.A(net436));
 sg13g2_antennanp ANTENNA_1849 (.A(net436));
 sg13g2_antennanp ANTENNA_1850 (.A(net436));
 sg13g2_antennanp ANTENNA_1851 (.A(net436));
 sg13g2_antennanp ANTENNA_1852 (.A(net436));
 sg13g2_antennanp ANTENNA_1853 (.A(net436));
 sg13g2_antennanp ANTENNA_1854 (.A(net436));
 sg13g2_antennanp ANTENNA_1855 (.A(net498));
 sg13g2_antennanp ANTENNA_1856 (.A(net498));
 sg13g2_antennanp ANTENNA_1857 (.A(net498));
 sg13g2_antennanp ANTENNA_1858 (.A(net498));
 sg13g2_antennanp ANTENNA_1859 (.A(net498));
 sg13g2_antennanp ANTENNA_1860 (.A(net498));
 sg13g2_antennanp ANTENNA_1861 (.A(net498));
 sg13g2_antennanp ANTENNA_1862 (.A(net498));
 sg13g2_antennanp ANTENNA_1863 (.A(net498));
 sg13g2_antennanp ANTENNA_1864 (.A(net525));
 sg13g2_antennanp ANTENNA_1865 (.A(net525));
 sg13g2_antennanp ANTENNA_1866 (.A(net525));
 sg13g2_antennanp ANTENNA_1867 (.A(net525));
 sg13g2_antennanp ANTENNA_1868 (.A(net525));
 sg13g2_antennanp ANTENNA_1869 (.A(net525));
 sg13g2_antennanp ANTENNA_1870 (.A(net525));
 sg13g2_antennanp ANTENNA_1871 (.A(net525));
 sg13g2_antennanp ANTENNA_1872 (.A(net525));
 sg13g2_antennanp ANTENNA_1873 (.A(net525));
 sg13g2_antennanp ANTENNA_1874 (.A(net1207));
 sg13g2_antennanp ANTENNA_1875 (.A(net1207));
 sg13g2_antennanp ANTENNA_1876 (.A(net1207));
 sg13g2_antennanp ANTENNA_1877 (.A(net1207));
 sg13g2_antennanp ANTENNA_1878 (.A(net1207));
 sg13g2_antennanp ANTENNA_1879 (.A(net1207));
 sg13g2_antennanp ANTENNA_1880 (.A(net1207));
 sg13g2_antennanp ANTENNA_1881 (.A(net1430));
 sg13g2_antennanp ANTENNA_1882 (.A(net1430));
 sg13g2_antennanp ANTENNA_1883 (.A(net1430));
 sg13g2_antennanp ANTENNA_1884 (.A(net1430));
 sg13g2_antennanp ANTENNA_1885 (.A(net1430));
 sg13g2_antennanp ANTENNA_1886 (.A(net1430));
 sg13g2_antennanp ANTENNA_1887 (.A(net1430));
 sg13g2_antennanp ANTENNA_1888 (.A(net1430));
 sg13g2_antennanp ANTENNA_1889 (.A(net1430));
 sg13g2_antennanp ANTENNA_1890 (.A(net1430));
 sg13g2_antennanp ANTENNA_1891 (.A(net1430));
 sg13g2_antennanp ANTENNA_1892 (.A(net1430));
 sg13g2_antennanp ANTENNA_1893 (.A(net1430));
 sg13g2_antennanp ANTENNA_1894 (.A(net1430));
 sg13g2_antennanp ANTENNA_1895 (.A(net1430));
 sg13g2_antennanp ANTENNA_1896 (.A(net1430));
 sg13g2_antennanp ANTENNA_1897 (.A(net1430));
 sg13g2_antennanp ANTENNA_1898 (.A(_00366_));
 sg13g2_antennanp ANTENNA_1899 (.A(_00366_));
 sg13g2_antennanp ANTENNA_1900 (.A(_00394_));
 sg13g2_antennanp ANTENNA_1901 (.A(_00394_));
 sg13g2_antennanp ANTENNA_1902 (.A(_00406_));
 sg13g2_antennanp ANTENNA_1903 (.A(_00406_));
 sg13g2_antennanp ANTENNA_1904 (.A(_00408_));
 sg13g2_antennanp ANTENNA_1905 (.A(_00411_));
 sg13g2_antennanp ANTENNA_1906 (.A(_00412_));
 sg13g2_antennanp ANTENNA_1907 (.A(_00413_));
 sg13g2_antennanp ANTENNA_1908 (.A(_00413_));
 sg13g2_antennanp ANTENNA_1909 (.A(_00417_));
 sg13g2_antennanp ANTENNA_1910 (.A(_03004_));
 sg13g2_antennanp ANTENNA_1911 (.A(_03004_));
 sg13g2_antennanp ANTENNA_1912 (.A(_03004_));
 sg13g2_antennanp ANTENNA_1913 (.A(_03145_));
 sg13g2_antennanp ANTENNA_1914 (.A(_03451_));
 sg13g2_antennanp ANTENNA_1915 (.A(_03451_));
 sg13g2_antennanp ANTENNA_1916 (.A(_03451_));
 sg13g2_antennanp ANTENNA_1917 (.A(_03451_));
 sg13g2_antennanp ANTENNA_1918 (.A(_03451_));
 sg13g2_antennanp ANTENNA_1919 (.A(_03451_));
 sg13g2_antennanp ANTENNA_1920 (.A(_04085_));
 sg13g2_antennanp ANTENNA_1921 (.A(_04085_));
 sg13g2_antennanp ANTENNA_1922 (.A(_04085_));
 sg13g2_antennanp ANTENNA_1923 (.A(_04086_));
 sg13g2_antennanp ANTENNA_1924 (.A(_04086_));
 sg13g2_antennanp ANTENNA_1925 (.A(_04086_));
 sg13g2_antennanp ANTENNA_1926 (.A(_04107_));
 sg13g2_antennanp ANTENNA_1927 (.A(_04743_));
 sg13g2_antennanp ANTENNA_1928 (.A(_04743_));
 sg13g2_antennanp ANTENNA_1929 (.A(_05412_));
 sg13g2_antennanp ANTENNA_1930 (.A(_05412_));
 sg13g2_antennanp ANTENNA_1931 (.A(_05412_));
 sg13g2_antennanp ANTENNA_1932 (.A(_05412_));
 sg13g2_antennanp ANTENNA_1933 (.A(_05412_));
 sg13g2_antennanp ANTENNA_1934 (.A(_05412_));
 sg13g2_antennanp ANTENNA_1935 (.A(_05436_));
 sg13g2_antennanp ANTENNA_1936 (.A(_05436_));
 sg13g2_antennanp ANTENNA_1937 (.A(_05436_));
 sg13g2_antennanp ANTENNA_1938 (.A(_05436_));
 sg13g2_antennanp ANTENNA_1939 (.A(_05495_));
 sg13g2_antennanp ANTENNA_1940 (.A(_05495_));
 sg13g2_antennanp ANTENNA_1941 (.A(_05495_));
 sg13g2_antennanp ANTENNA_1942 (.A(_05592_));
 sg13g2_antennanp ANTENNA_1943 (.A(_05621_));
 sg13g2_antennanp ANTENNA_1944 (.A(_05631_));
 sg13g2_antennanp ANTENNA_1945 (.A(_05639_));
 sg13g2_antennanp ANTENNA_1946 (.A(_05689_));
 sg13g2_antennanp ANTENNA_1947 (.A(_05719_));
 sg13g2_antennanp ANTENNA_1948 (.A(_05719_));
 sg13g2_antennanp ANTENNA_1949 (.A(_05719_));
 sg13g2_antennanp ANTENNA_1950 (.A(_05719_));
 sg13g2_antennanp ANTENNA_1951 (.A(_05719_));
 sg13g2_antennanp ANTENNA_1952 (.A(_05739_));
 sg13g2_antennanp ANTENNA_1953 (.A(_05773_));
 sg13g2_antennanp ANTENNA_1954 (.A(_05781_));
 sg13g2_antennanp ANTENNA_1955 (.A(_05785_));
 sg13g2_antennanp ANTENNA_1956 (.A(_05807_));
 sg13g2_antennanp ANTENNA_1957 (.A(_05825_));
 sg13g2_antennanp ANTENNA_1958 (.A(_05825_));
 sg13g2_antennanp ANTENNA_1959 (.A(_05825_));
 sg13g2_antennanp ANTENNA_1960 (.A(_05825_));
 sg13g2_antennanp ANTENNA_1961 (.A(_05825_));
 sg13g2_antennanp ANTENNA_1962 (.A(_05825_));
 sg13g2_antennanp ANTENNA_1963 (.A(_05829_));
 sg13g2_antennanp ANTENNA_1964 (.A(_05858_));
 sg13g2_antennanp ANTENNA_1965 (.A(_05866_));
 sg13g2_antennanp ANTENNA_1966 (.A(_05877_));
 sg13g2_antennanp ANTENNA_1967 (.A(_05889_));
 sg13g2_antennanp ANTENNA_1968 (.A(_05889_));
 sg13g2_antennanp ANTENNA_1969 (.A(_05889_));
 sg13g2_antennanp ANTENNA_1970 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1971 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1972 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1973 (.A(_05942_));
 sg13g2_antennanp ANTENNA_1974 (.A(_05977_));
 sg13g2_antennanp ANTENNA_1975 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1976 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1977 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1978 (.A(_05999_));
 sg13g2_antennanp ANTENNA_1979 (.A(_06027_));
 sg13g2_antennanp ANTENNA_1980 (.A(_06038_));
 sg13g2_antennanp ANTENNA_1981 (.A(_06045_));
 sg13g2_antennanp ANTENNA_1982 (.A(_06053_));
 sg13g2_antennanp ANTENNA_1983 (.A(_06065_));
 sg13g2_antennanp ANTENNA_1984 (.A(_06065_));
 sg13g2_antennanp ANTENNA_1985 (.A(_06065_));
 sg13g2_antennanp ANTENNA_1986 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1987 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1988 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1989 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1990 (.A(_06152_));
 sg13g2_antennanp ANTENNA_1991 (.A(_06163_));
 sg13g2_antennanp ANTENNA_1992 (.A(_06163_));
 sg13g2_antennanp ANTENNA_1993 (.A(_06163_));
 sg13g2_antennanp ANTENNA_1994 (.A(_06183_));
 sg13g2_antennanp ANTENNA_1995 (.A(_06183_));
 sg13g2_antennanp ANTENNA_1996 (.A(_06183_));
 sg13g2_antennanp ANTENNA_1997 (.A(_06183_));
 sg13g2_antennanp ANTENNA_1998 (.A(_06195_));
 sg13g2_antennanp ANTENNA_1999 (.A(_06216_));
 sg13g2_antennanp ANTENNA_2000 (.A(_06216_));
 sg13g2_antennanp ANTENNA_2001 (.A(_06236_));
 sg13g2_antennanp ANTENNA_2002 (.A(_06247_));
 sg13g2_antennanp ANTENNA_2003 (.A(_06259_));
 sg13g2_antennanp ANTENNA_2004 (.A(_06285_));
 sg13g2_antennanp ANTENNA_2005 (.A(_06303_));
 sg13g2_antennanp ANTENNA_2006 (.A(_06318_));
 sg13g2_antennanp ANTENNA_2007 (.A(_06337_));
 sg13g2_antennanp ANTENNA_2008 (.A(_06350_));
 sg13g2_antennanp ANTENNA_2009 (.A(_06355_));
 sg13g2_antennanp ANTENNA_2010 (.A(_06370_));
 sg13g2_antennanp ANTENNA_2011 (.A(_06380_));
 sg13g2_antennanp ANTENNA_2012 (.A(_06385_));
 sg13g2_antennanp ANTENNA_2013 (.A(_06391_));
 sg13g2_antennanp ANTENNA_2014 (.A(_06423_));
 sg13g2_antennanp ANTENNA_2015 (.A(_06435_));
 sg13g2_antennanp ANTENNA_2016 (.A(_06438_));
 sg13g2_antennanp ANTENNA_2017 (.A(_06464_));
 sg13g2_antennanp ANTENNA_2018 (.A(_06475_));
 sg13g2_antennanp ANTENNA_2019 (.A(_06525_));
 sg13g2_antennanp ANTENNA_2020 (.A(_06530_));
 sg13g2_antennanp ANTENNA_2021 (.A(_06532_));
 sg13g2_antennanp ANTENNA_2022 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2023 (.A(_06605_));
 sg13g2_antennanp ANTENNA_2024 (.A(_06653_));
 sg13g2_antennanp ANTENNA_2025 (.A(_06660_));
 sg13g2_antennanp ANTENNA_2026 (.A(_06667_));
 sg13g2_antennanp ANTENNA_2027 (.A(_06671_));
 sg13g2_antennanp ANTENNA_2028 (.A(_06697_));
 sg13g2_antennanp ANTENNA_2029 (.A(_06701_));
 sg13g2_antennanp ANTENNA_2030 (.A(_06703_));
 sg13g2_antennanp ANTENNA_2031 (.A(_06751_));
 sg13g2_antennanp ANTENNA_2032 (.A(_06772_));
 sg13g2_antennanp ANTENNA_2033 (.A(_06813_));
 sg13g2_antennanp ANTENNA_2034 (.A(_06815_));
 sg13g2_antennanp ANTENNA_2035 (.A(_06816_));
 sg13g2_antennanp ANTENNA_2036 (.A(_06829_));
 sg13g2_antennanp ANTENNA_2037 (.A(_06850_));
 sg13g2_antennanp ANTENNA_2038 (.A(_06854_));
 sg13g2_antennanp ANTENNA_2039 (.A(_06854_));
 sg13g2_antennanp ANTENNA_2040 (.A(_06869_));
 sg13g2_antennanp ANTENNA_2041 (.A(_06870_));
 sg13g2_antennanp ANTENNA_2042 (.A(_06875_));
 sg13g2_antennanp ANTENNA_2043 (.A(_06881_));
 sg13g2_antennanp ANTENNA_2044 (.A(_06901_));
 sg13g2_antennanp ANTENNA_2045 (.A(_06921_));
 sg13g2_antennanp ANTENNA_2046 (.A(_06932_));
 sg13g2_antennanp ANTENNA_2047 (.A(_06936_));
 sg13g2_antennanp ANTENNA_2048 (.A(_06936_));
 sg13g2_antennanp ANTENNA_2049 (.A(_06959_));
 sg13g2_antennanp ANTENNA_2050 (.A(_06993_));
 sg13g2_antennanp ANTENNA_2051 (.A(_06998_));
 sg13g2_antennanp ANTENNA_2052 (.A(_07008_));
 sg13g2_antennanp ANTENNA_2053 (.A(_07035_));
 sg13g2_antennanp ANTENNA_2054 (.A(_07036_));
 sg13g2_antennanp ANTENNA_2055 (.A(_07047_));
 sg13g2_antennanp ANTENNA_2056 (.A(_07060_));
 sg13g2_antennanp ANTENNA_2057 (.A(_07069_));
 sg13g2_antennanp ANTENNA_2058 (.A(_07074_));
 sg13g2_antennanp ANTENNA_2059 (.A(_07080_));
 sg13g2_antennanp ANTENNA_2060 (.A(_07108_));
 sg13g2_antennanp ANTENNA_2061 (.A(_07139_));
 sg13g2_antennanp ANTENNA_2062 (.A(_07146_));
 sg13g2_antennanp ANTENNA_2063 (.A(_07191_));
 sg13g2_antennanp ANTENNA_2064 (.A(_07212_));
 sg13g2_antennanp ANTENNA_2065 (.A(_07217_));
 sg13g2_antennanp ANTENNA_2066 (.A(_07282_));
 sg13g2_antennanp ANTENNA_2067 (.A(_07284_));
 sg13g2_antennanp ANTENNA_2068 (.A(_07288_));
 sg13g2_antennanp ANTENNA_2069 (.A(_07288_));
 sg13g2_antennanp ANTENNA_2070 (.A(_07302_));
 sg13g2_antennanp ANTENNA_2071 (.A(_07312_));
 sg13g2_antennanp ANTENNA_2072 (.A(_07363_));
 sg13g2_antennanp ANTENNA_2073 (.A(_07375_));
 sg13g2_antennanp ANTENNA_2074 (.A(_07403_));
 sg13g2_antennanp ANTENNA_2075 (.A(_07428_));
 sg13g2_antennanp ANTENNA_2076 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2077 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2078 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2079 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2080 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2081 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2082 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2083 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2084 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2085 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2086 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2087 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2088 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2089 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2090 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2091 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2092 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2093 (.A(_07496_));
 sg13g2_antennanp ANTENNA_2094 (.A(_07496_));
 sg13g2_antennanp ANTENNA_2095 (.A(_07496_));
 sg13g2_antennanp ANTENNA_2096 (.A(_07496_));
 sg13g2_antennanp ANTENNA_2097 (.A(_07609_));
 sg13g2_antennanp ANTENNA_2098 (.A(_07622_));
 sg13g2_antennanp ANTENNA_2099 (.A(_07636_));
 sg13g2_antennanp ANTENNA_2100 (.A(_07704_));
 sg13g2_antennanp ANTENNA_2101 (.A(_07704_));
 sg13g2_antennanp ANTENNA_2102 (.A(_07730_));
 sg13g2_antennanp ANTENNA_2103 (.A(_07758_));
 sg13g2_antennanp ANTENNA_2104 (.A(_07822_));
 sg13g2_antennanp ANTENNA_2105 (.A(_07835_));
 sg13g2_antennanp ANTENNA_2106 (.A(_07835_));
 sg13g2_antennanp ANTENNA_2107 (.A(_07914_));
 sg13g2_antennanp ANTENNA_2108 (.A(_07926_));
 sg13g2_antennanp ANTENNA_2109 (.A(_07939_));
 sg13g2_antennanp ANTENNA_2110 (.A(_07952_));
 sg13g2_antennanp ANTENNA_2111 (.A(_08169_));
 sg13g2_antennanp ANTENNA_2112 (.A(_08169_));
 sg13g2_antennanp ANTENNA_2113 (.A(_09280_));
 sg13g2_antennanp ANTENNA_2114 (.A(_09280_));
 sg13g2_antennanp ANTENNA_2115 (.A(_09280_));
 sg13g2_antennanp ANTENNA_2116 (.A(_09280_));
 sg13g2_antennanp ANTENNA_2117 (.A(_09280_));
 sg13g2_antennanp ANTENNA_2118 (.A(_09724_));
 sg13g2_antennanp ANTENNA_2119 (.A(_09825_));
 sg13g2_antennanp ANTENNA_2120 (.A(_09825_));
 sg13g2_antennanp ANTENNA_2121 (.A(_09825_));
 sg13g2_antennanp ANTENNA_2122 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2123 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2124 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2125 (.A(_10247_));
 sg13g2_antennanp ANTENNA_2126 (.A(_10247_));
 sg13g2_antennanp ANTENNA_2127 (.A(_10247_));
 sg13g2_antennanp ANTENNA_2128 (.A(_10518_));
 sg13g2_antennanp ANTENNA_2129 (.A(_10518_));
 sg13g2_antennanp ANTENNA_2130 (.A(_10604_));
 sg13g2_antennanp ANTENNA_2131 (.A(_10604_));
 sg13g2_antennanp ANTENNA_2132 (.A(_10604_));
 sg13g2_antennanp ANTENNA_2133 (.A(_10604_));
 sg13g2_antennanp ANTENNA_2134 (.A(_10617_));
 sg13g2_antennanp ANTENNA_2135 (.A(_10952_));
 sg13g2_antennanp ANTENNA_2136 (.A(_10963_));
 sg13g2_antennanp ANTENNA_2137 (.A(_11000_));
 sg13g2_antennanp ANTENNA_2138 (.A(_11000_));
 sg13g2_antennanp ANTENNA_2139 (.A(_11000_));
 sg13g2_antennanp ANTENNA_2140 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2141 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2142 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2143 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2144 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2145 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2146 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2147 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2148 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2149 (.A(\top_ihp.oisc.op_a[22] ));
 sg13g2_antennanp ANTENNA_2150 (.A(\top_ihp.oisc.op_a[27] ));
 sg13g2_antennanp ANTENNA_2151 (.A(\top_ihp.oisc.op_a[6] ));
 sg13g2_antennanp ANTENNA_2152 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_2153 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_2154 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_2155 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_2156 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_2157 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_2158 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_2159 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_2160 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_2161 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_2162 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_2163 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_2164 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_2165 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_2166 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_2167 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_2168 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_2169 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_2170 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_2171 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_2172 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_2173 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_2174 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_2175 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_2176 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_2177 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_2178 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_2179 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_2180 (.A(\top_ihp.tx ));
 sg13g2_antennanp ANTENNA_2181 (.A(net1));
 sg13g2_antennanp ANTENNA_2182 (.A(net1));
 sg13g2_antennanp ANTENNA_2183 (.A(net1));
 sg13g2_antennanp ANTENNA_2184 (.A(net5));
 sg13g2_antennanp ANTENNA_2185 (.A(net10));
 sg13g2_antennanp ANTENNA_2186 (.A(net77));
 sg13g2_antennanp ANTENNA_2187 (.A(net77));
 sg13g2_antennanp ANTENNA_2188 (.A(net77));
 sg13g2_antennanp ANTENNA_2189 (.A(net77));
 sg13g2_antennanp ANTENNA_2190 (.A(net77));
 sg13g2_antennanp ANTENNA_2191 (.A(net77));
 sg13g2_antennanp ANTENNA_2192 (.A(net77));
 sg13g2_antennanp ANTENNA_2193 (.A(net77));
 sg13g2_antennanp ANTENNA_2194 (.A(net77));
 sg13g2_antennanp ANTENNA_2195 (.A(net91));
 sg13g2_antennanp ANTENNA_2196 (.A(net91));
 sg13g2_antennanp ANTENNA_2197 (.A(net91));
 sg13g2_antennanp ANTENNA_2198 (.A(net91));
 sg13g2_antennanp ANTENNA_2199 (.A(net91));
 sg13g2_antennanp ANTENNA_2200 (.A(net91));
 sg13g2_antennanp ANTENNA_2201 (.A(net91));
 sg13g2_antennanp ANTENNA_2202 (.A(net91));
 sg13g2_antennanp ANTENNA_2203 (.A(net91));
 sg13g2_antennanp ANTENNA_2204 (.A(net146));
 sg13g2_antennanp ANTENNA_2205 (.A(net146));
 sg13g2_antennanp ANTENNA_2206 (.A(net146));
 sg13g2_antennanp ANTENNA_2207 (.A(net146));
 sg13g2_antennanp ANTENNA_2208 (.A(net146));
 sg13g2_antennanp ANTENNA_2209 (.A(net146));
 sg13g2_antennanp ANTENNA_2210 (.A(net146));
 sg13g2_antennanp ANTENNA_2211 (.A(net146));
 sg13g2_antennanp ANTENNA_2212 (.A(net146));
 sg13g2_antennanp ANTENNA_2213 (.A(net146));
 sg13g2_antennanp ANTENNA_2214 (.A(net146));
 sg13g2_antennanp ANTENNA_2215 (.A(net146));
 sg13g2_antennanp ANTENNA_2216 (.A(net155));
 sg13g2_antennanp ANTENNA_2217 (.A(net155));
 sg13g2_antennanp ANTENNA_2218 (.A(net155));
 sg13g2_antennanp ANTENNA_2219 (.A(net155));
 sg13g2_antennanp ANTENNA_2220 (.A(net155));
 sg13g2_antennanp ANTENNA_2221 (.A(net155));
 sg13g2_antennanp ANTENNA_2222 (.A(net155));
 sg13g2_antennanp ANTENNA_2223 (.A(net155));
 sg13g2_antennanp ANTENNA_2224 (.A(net155));
 sg13g2_antennanp ANTENNA_2225 (.A(net155));
 sg13g2_antennanp ANTENNA_2226 (.A(net155));
 sg13g2_antennanp ANTENNA_2227 (.A(net292));
 sg13g2_antennanp ANTENNA_2228 (.A(net292));
 sg13g2_antennanp ANTENNA_2229 (.A(net292));
 sg13g2_antennanp ANTENNA_2230 (.A(net292));
 sg13g2_antennanp ANTENNA_2231 (.A(net292));
 sg13g2_antennanp ANTENNA_2232 (.A(net292));
 sg13g2_antennanp ANTENNA_2233 (.A(net292));
 sg13g2_antennanp ANTENNA_2234 (.A(net292));
 sg13g2_antennanp ANTENNA_2235 (.A(net308));
 sg13g2_antennanp ANTENNA_2236 (.A(net308));
 sg13g2_antennanp ANTENNA_2237 (.A(net308));
 sg13g2_antennanp ANTENNA_2238 (.A(net308));
 sg13g2_antennanp ANTENNA_2239 (.A(net308));
 sg13g2_antennanp ANTENNA_2240 (.A(net308));
 sg13g2_antennanp ANTENNA_2241 (.A(net308));
 sg13g2_antennanp ANTENNA_2242 (.A(net308));
 sg13g2_antennanp ANTENNA_2243 (.A(net308));
 sg13g2_antennanp ANTENNA_2244 (.A(net317));
 sg13g2_antennanp ANTENNA_2245 (.A(net317));
 sg13g2_antennanp ANTENNA_2246 (.A(net317));
 sg13g2_antennanp ANTENNA_2247 (.A(net317));
 sg13g2_antennanp ANTENNA_2248 (.A(net317));
 sg13g2_antennanp ANTENNA_2249 (.A(net317));
 sg13g2_antennanp ANTENNA_2250 (.A(net317));
 sg13g2_antennanp ANTENNA_2251 (.A(net317));
 sg13g2_antennanp ANTENNA_2252 (.A(net317));
 sg13g2_antennanp ANTENNA_2253 (.A(net397));
 sg13g2_antennanp ANTENNA_2254 (.A(net397));
 sg13g2_antennanp ANTENNA_2255 (.A(net397));
 sg13g2_antennanp ANTENNA_2256 (.A(net397));
 sg13g2_antennanp ANTENNA_2257 (.A(net397));
 sg13g2_antennanp ANTENNA_2258 (.A(net397));
 sg13g2_antennanp ANTENNA_2259 (.A(net397));
 sg13g2_antennanp ANTENNA_2260 (.A(net397));
 sg13g2_antennanp ANTENNA_2261 (.A(net397));
 sg13g2_antennanp ANTENNA_2262 (.A(net498));
 sg13g2_antennanp ANTENNA_2263 (.A(net498));
 sg13g2_antennanp ANTENNA_2264 (.A(net498));
 sg13g2_antennanp ANTENNA_2265 (.A(net498));
 sg13g2_antennanp ANTENNA_2266 (.A(net498));
 sg13g2_antennanp ANTENNA_2267 (.A(net498));
 sg13g2_antennanp ANTENNA_2268 (.A(net498));
 sg13g2_antennanp ANTENNA_2269 (.A(net498));
 sg13g2_antennanp ANTENNA_2270 (.A(net498));
 sg13g2_antennanp ANTENNA_2271 (.A(net525));
 sg13g2_antennanp ANTENNA_2272 (.A(net525));
 sg13g2_antennanp ANTENNA_2273 (.A(net525));
 sg13g2_antennanp ANTENNA_2274 (.A(net525));
 sg13g2_antennanp ANTENNA_2275 (.A(net525));
 sg13g2_antennanp ANTENNA_2276 (.A(net525));
 sg13g2_antennanp ANTENNA_2277 (.A(net525));
 sg13g2_antennanp ANTENNA_2278 (.A(net525));
 sg13g2_antennanp ANTENNA_2279 (.A(net525));
 sg13g2_antennanp ANTENNA_2280 (.A(net525));
 sg13g2_antennanp ANTENNA_2281 (.A(net525));
 sg13g2_antennanp ANTENNA_2282 (.A(net525));
 sg13g2_antennanp ANTENNA_2283 (.A(net525));
 sg13g2_antennanp ANTENNA_2284 (.A(net525));
 sg13g2_antennanp ANTENNA_2285 (.A(net525));
 sg13g2_antennanp ANTENNA_2286 (.A(net803));
 sg13g2_antennanp ANTENNA_2287 (.A(net803));
 sg13g2_antennanp ANTENNA_2288 (.A(net803));
 sg13g2_antennanp ANTENNA_2289 (.A(net803));
 sg13g2_antennanp ANTENNA_2290 (.A(net803));
 sg13g2_antennanp ANTENNA_2291 (.A(net803));
 sg13g2_antennanp ANTENNA_2292 (.A(net803));
 sg13g2_antennanp ANTENNA_2293 (.A(net803));
 sg13g2_antennanp ANTENNA_2294 (.A(net803));
 sg13g2_antennanp ANTENNA_2295 (.A(net1207));
 sg13g2_antennanp ANTENNA_2296 (.A(net1207));
 sg13g2_antennanp ANTENNA_2297 (.A(net1207));
 sg13g2_antennanp ANTENNA_2298 (.A(net1207));
 sg13g2_antennanp ANTENNA_2299 (.A(net1207));
 sg13g2_antennanp ANTENNA_2300 (.A(net1207));
 sg13g2_antennanp ANTENNA_2301 (.A(net1207));
 sg13g2_antennanp ANTENNA_2302 (.A(net1430));
 sg13g2_antennanp ANTENNA_2303 (.A(net1430));
 sg13g2_antennanp ANTENNA_2304 (.A(net1430));
 sg13g2_antennanp ANTENNA_2305 (.A(net1430));
 sg13g2_antennanp ANTENNA_2306 (.A(net1430));
 sg13g2_antennanp ANTENNA_2307 (.A(net1430));
 sg13g2_antennanp ANTENNA_2308 (.A(net1430));
 sg13g2_antennanp ANTENNA_2309 (.A(_00366_));
 sg13g2_antennanp ANTENNA_2310 (.A(_00366_));
 sg13g2_antennanp ANTENNA_2311 (.A(_00394_));
 sg13g2_antennanp ANTENNA_2312 (.A(_00394_));
 sg13g2_antennanp ANTENNA_2313 (.A(_00408_));
 sg13g2_antennanp ANTENNA_2314 (.A(_00411_));
 sg13g2_antennanp ANTENNA_2315 (.A(_00412_));
 sg13g2_antennanp ANTENNA_2316 (.A(_00413_));
 sg13g2_antennanp ANTENNA_2317 (.A(_00413_));
 sg13g2_antennanp ANTENNA_2318 (.A(_00417_));
 sg13g2_antennanp ANTENNA_2319 (.A(_03004_));
 sg13g2_antennanp ANTENNA_2320 (.A(_03004_));
 sg13g2_antennanp ANTENNA_2321 (.A(_03004_));
 sg13g2_antennanp ANTENNA_2322 (.A(_03145_));
 sg13g2_antennanp ANTENNA_2323 (.A(_03451_));
 sg13g2_antennanp ANTENNA_2324 (.A(_03451_));
 sg13g2_antennanp ANTENNA_2325 (.A(_03451_));
 sg13g2_antennanp ANTENNA_2326 (.A(_03451_));
 sg13g2_antennanp ANTENNA_2327 (.A(_03451_));
 sg13g2_antennanp ANTENNA_2328 (.A(_03451_));
 sg13g2_antennanp ANTENNA_2329 (.A(_04085_));
 sg13g2_antennanp ANTENNA_2330 (.A(_04085_));
 sg13g2_antennanp ANTENNA_2331 (.A(_04085_));
 sg13g2_antennanp ANTENNA_2332 (.A(_04086_));
 sg13g2_antennanp ANTENNA_2333 (.A(_04086_));
 sg13g2_antennanp ANTENNA_2334 (.A(_04086_));
 sg13g2_antennanp ANTENNA_2335 (.A(_04107_));
 sg13g2_antennanp ANTENNA_2336 (.A(_04743_));
 sg13g2_antennanp ANTENNA_2337 (.A(_04743_));
 sg13g2_antennanp ANTENNA_2338 (.A(_05412_));
 sg13g2_antennanp ANTENNA_2339 (.A(_05412_));
 sg13g2_antennanp ANTENNA_2340 (.A(_05412_));
 sg13g2_antennanp ANTENNA_2341 (.A(_05412_));
 sg13g2_antennanp ANTENNA_2342 (.A(_05412_));
 sg13g2_antennanp ANTENNA_2343 (.A(_05412_));
 sg13g2_antennanp ANTENNA_2344 (.A(_05412_));
 sg13g2_antennanp ANTENNA_2345 (.A(_05412_));
 sg13g2_antennanp ANTENNA_2346 (.A(_05430_));
 sg13g2_antennanp ANTENNA_2347 (.A(_05430_));
 sg13g2_antennanp ANTENNA_2348 (.A(_05430_));
 sg13g2_antennanp ANTENNA_2349 (.A(_05430_));
 sg13g2_antennanp ANTENNA_2350 (.A(_05430_));
 sg13g2_antennanp ANTENNA_2351 (.A(_05430_));
 sg13g2_antennanp ANTENNA_2352 (.A(_05430_));
 sg13g2_antennanp ANTENNA_2353 (.A(_05430_));
 sg13g2_antennanp ANTENNA_2354 (.A(_05430_));
 sg13g2_antennanp ANTENNA_2355 (.A(_05430_));
 sg13g2_antennanp ANTENNA_2356 (.A(_05436_));
 sg13g2_antennanp ANTENNA_2357 (.A(_05436_));
 sg13g2_antennanp ANTENNA_2358 (.A(_05436_));
 sg13g2_antennanp ANTENNA_2359 (.A(_05436_));
 sg13g2_antennanp ANTENNA_2360 (.A(_05495_));
 sg13g2_antennanp ANTENNA_2361 (.A(_05495_));
 sg13g2_antennanp ANTENNA_2362 (.A(_05495_));
 sg13g2_antennanp ANTENNA_2363 (.A(_05592_));
 sg13g2_antennanp ANTENNA_2364 (.A(_05621_));
 sg13g2_antennanp ANTENNA_2365 (.A(_05631_));
 sg13g2_antennanp ANTENNA_2366 (.A(_05639_));
 sg13g2_antennanp ANTENNA_2367 (.A(_05648_));
 sg13g2_antennanp ANTENNA_2368 (.A(_05648_));
 sg13g2_antennanp ANTENNA_2369 (.A(_05648_));
 sg13g2_antennanp ANTENNA_2370 (.A(_05689_));
 sg13g2_antennanp ANTENNA_2371 (.A(_05719_));
 sg13g2_antennanp ANTENNA_2372 (.A(_05719_));
 sg13g2_antennanp ANTENNA_2373 (.A(_05719_));
 sg13g2_antennanp ANTENNA_2374 (.A(_05719_));
 sg13g2_antennanp ANTENNA_2375 (.A(_05719_));
 sg13g2_antennanp ANTENNA_2376 (.A(_05739_));
 sg13g2_antennanp ANTENNA_2377 (.A(_05773_));
 sg13g2_antennanp ANTENNA_2378 (.A(_05781_));
 sg13g2_antennanp ANTENNA_2379 (.A(_05782_));
 sg13g2_antennanp ANTENNA_2380 (.A(_05782_));
 sg13g2_antennanp ANTENNA_2381 (.A(_05782_));
 sg13g2_antennanp ANTENNA_2382 (.A(_05785_));
 sg13g2_antennanp ANTENNA_2383 (.A(_05807_));
 sg13g2_antennanp ANTENNA_2384 (.A(_05825_));
 sg13g2_antennanp ANTENNA_2385 (.A(_05825_));
 sg13g2_antennanp ANTENNA_2386 (.A(_05825_));
 sg13g2_antennanp ANTENNA_2387 (.A(_05825_));
 sg13g2_antennanp ANTENNA_2388 (.A(_05825_));
 sg13g2_antennanp ANTENNA_2389 (.A(_05825_));
 sg13g2_antennanp ANTENNA_2390 (.A(_05829_));
 sg13g2_antennanp ANTENNA_2391 (.A(_05858_));
 sg13g2_antennanp ANTENNA_2392 (.A(_05866_));
 sg13g2_antennanp ANTENNA_2393 (.A(_05877_));
 sg13g2_antennanp ANTENNA_2394 (.A(_05900_));
 sg13g2_antennanp ANTENNA_2395 (.A(_05900_));
 sg13g2_antennanp ANTENNA_2396 (.A(_05900_));
 sg13g2_antennanp ANTENNA_2397 (.A(_05942_));
 sg13g2_antennanp ANTENNA_2398 (.A(_05977_));
 sg13g2_antennanp ANTENNA_2399 (.A(_05999_));
 sg13g2_antennanp ANTENNA_2400 (.A(_05999_));
 sg13g2_antennanp ANTENNA_2401 (.A(_05999_));
 sg13g2_antennanp ANTENNA_2402 (.A(_05999_));
 sg13g2_antennanp ANTENNA_2403 (.A(_06027_));
 sg13g2_antennanp ANTENNA_2404 (.A(_06038_));
 sg13g2_antennanp ANTENNA_2405 (.A(_06045_));
 sg13g2_antennanp ANTENNA_2406 (.A(_06053_));
 sg13g2_antennanp ANTENNA_2407 (.A(_06065_));
 sg13g2_antennanp ANTENNA_2408 (.A(_06065_));
 sg13g2_antennanp ANTENNA_2409 (.A(_06065_));
 sg13g2_antennanp ANTENNA_2410 (.A(_06146_));
 sg13g2_antennanp ANTENNA_2411 (.A(_06146_));
 sg13g2_antennanp ANTENNA_2412 (.A(_06146_));
 sg13g2_antennanp ANTENNA_2413 (.A(_06146_));
 sg13g2_antennanp ANTENNA_2414 (.A(_06152_));
 sg13g2_antennanp ANTENNA_2415 (.A(_06163_));
 sg13g2_antennanp ANTENNA_2416 (.A(_06163_));
 sg13g2_antennanp ANTENNA_2417 (.A(_06163_));
 sg13g2_antennanp ANTENNA_2418 (.A(_06183_));
 sg13g2_antennanp ANTENNA_2419 (.A(_06183_));
 sg13g2_antennanp ANTENNA_2420 (.A(_06183_));
 sg13g2_antennanp ANTENNA_2421 (.A(_06183_));
 sg13g2_antennanp ANTENNA_2422 (.A(_06195_));
 sg13g2_antennanp ANTENNA_2423 (.A(_06216_));
 sg13g2_antennanp ANTENNA_2424 (.A(_06236_));
 sg13g2_antennanp ANTENNA_2425 (.A(_06247_));
 sg13g2_antennanp ANTENNA_2426 (.A(_06259_));
 sg13g2_antennanp ANTENNA_2427 (.A(_06285_));
 sg13g2_antennanp ANTENNA_2428 (.A(_06303_));
 sg13g2_antennanp ANTENNA_2429 (.A(_06318_));
 sg13g2_antennanp ANTENNA_2430 (.A(_06337_));
 sg13g2_antennanp ANTENNA_2431 (.A(_06350_));
 sg13g2_antennanp ANTENNA_2432 (.A(_06355_));
 sg13g2_antennanp ANTENNA_2433 (.A(_06370_));
 sg13g2_antennanp ANTENNA_2434 (.A(_06380_));
 sg13g2_antennanp ANTENNA_2435 (.A(_06380_));
 sg13g2_antennanp ANTENNA_2436 (.A(_06385_));
 sg13g2_antennanp ANTENNA_2437 (.A(_06391_));
 sg13g2_antennanp ANTENNA_2438 (.A(_06423_));
 sg13g2_antennanp ANTENNA_2439 (.A(_06435_));
 sg13g2_antennanp ANTENNA_2440 (.A(_06438_));
 sg13g2_antennanp ANTENNA_2441 (.A(_06464_));
 sg13g2_antennanp ANTENNA_2442 (.A(_06475_));
 sg13g2_antennanp ANTENNA_2443 (.A(_06525_));
 sg13g2_antennanp ANTENNA_2444 (.A(_06530_));
 sg13g2_antennanp ANTENNA_2445 (.A(_06532_));
 sg13g2_antennanp ANTENNA_2446 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2447 (.A(_06605_));
 sg13g2_antennanp ANTENNA_2448 (.A(_06653_));
 sg13g2_antennanp ANTENNA_2449 (.A(_06660_));
 sg13g2_antennanp ANTENNA_2450 (.A(_06667_));
 sg13g2_antennanp ANTENNA_2451 (.A(_06671_));
 sg13g2_antennanp ANTENNA_2452 (.A(_06671_));
 sg13g2_antennanp ANTENNA_2453 (.A(_06697_));
 sg13g2_antennanp ANTENNA_2454 (.A(_06701_));
 sg13g2_antennanp ANTENNA_2455 (.A(_06703_));
 sg13g2_antennanp ANTENNA_2456 (.A(_06751_));
 sg13g2_antennanp ANTENNA_2457 (.A(_06772_));
 sg13g2_antennanp ANTENNA_2458 (.A(_06813_));
 sg13g2_antennanp ANTENNA_2459 (.A(_06815_));
 sg13g2_antennanp ANTENNA_2460 (.A(_06816_));
 sg13g2_antennanp ANTENNA_2461 (.A(_06829_));
 sg13g2_antennanp ANTENNA_2462 (.A(_06850_));
 sg13g2_antennanp ANTENNA_2463 (.A(_06854_));
 sg13g2_antennanp ANTENNA_2464 (.A(_06854_));
 sg13g2_antennanp ANTENNA_2465 (.A(_06869_));
 sg13g2_antennanp ANTENNA_2466 (.A(_06870_));
 sg13g2_antennanp ANTENNA_2467 (.A(_06875_));
 sg13g2_antennanp ANTENNA_2468 (.A(_06881_));
 sg13g2_antennanp ANTENNA_2469 (.A(_06901_));
 sg13g2_antennanp ANTENNA_2470 (.A(_06932_));
 sg13g2_antennanp ANTENNA_2471 (.A(_06936_));
 sg13g2_antennanp ANTENNA_2472 (.A(_06959_));
 sg13g2_antennanp ANTENNA_2473 (.A(_06993_));
 sg13g2_antennanp ANTENNA_2474 (.A(_06998_));
 sg13g2_antennanp ANTENNA_2475 (.A(_07008_));
 sg13g2_antennanp ANTENNA_2476 (.A(_07035_));
 sg13g2_antennanp ANTENNA_2477 (.A(_07036_));
 sg13g2_antennanp ANTENNA_2478 (.A(_07047_));
 sg13g2_antennanp ANTENNA_2479 (.A(_07060_));
 sg13g2_antennanp ANTENNA_2480 (.A(_07069_));
 sg13g2_antennanp ANTENNA_2481 (.A(_07074_));
 sg13g2_antennanp ANTENNA_2482 (.A(_07080_));
 sg13g2_antennanp ANTENNA_2483 (.A(_07108_));
 sg13g2_antennanp ANTENNA_2484 (.A(_07146_));
 sg13g2_antennanp ANTENNA_2485 (.A(_07191_));
 sg13g2_antennanp ANTENNA_2486 (.A(_07212_));
 sg13g2_antennanp ANTENNA_2487 (.A(_07217_));
 sg13g2_antennanp ANTENNA_2488 (.A(_07282_));
 sg13g2_antennanp ANTENNA_2489 (.A(_07284_));
 sg13g2_antennanp ANTENNA_2490 (.A(_07288_));
 sg13g2_antennanp ANTENNA_2491 (.A(_07302_));
 sg13g2_antennanp ANTENNA_2492 (.A(_07312_));
 sg13g2_antennanp ANTENNA_2493 (.A(_07363_));
 sg13g2_antennanp ANTENNA_2494 (.A(_07375_));
 sg13g2_antennanp ANTENNA_2495 (.A(_07403_));
 sg13g2_antennanp ANTENNA_2496 (.A(_07428_));
 sg13g2_antennanp ANTENNA_2497 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2498 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2499 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2500 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2501 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2502 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2503 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2504 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2505 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2506 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2507 (.A(_07460_));
 sg13g2_antennanp ANTENNA_2508 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2509 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2510 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2511 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2512 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2513 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2514 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2515 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2516 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2517 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2518 (.A(_07491_));
 sg13g2_antennanp ANTENNA_2519 (.A(_07496_));
 sg13g2_antennanp ANTENNA_2520 (.A(_07496_));
 sg13g2_antennanp ANTENNA_2521 (.A(_07496_));
 sg13g2_antennanp ANTENNA_2522 (.A(_07496_));
 sg13g2_antennanp ANTENNA_2523 (.A(_07609_));
 sg13g2_antennanp ANTENNA_2524 (.A(_07622_));
 sg13g2_antennanp ANTENNA_2525 (.A(_07636_));
 sg13g2_antennanp ANTENNA_2526 (.A(_07704_));
 sg13g2_antennanp ANTENNA_2527 (.A(_07704_));
 sg13g2_antennanp ANTENNA_2528 (.A(_07730_));
 sg13g2_antennanp ANTENNA_2529 (.A(_07730_));
 sg13g2_antennanp ANTENNA_2530 (.A(_07758_));
 sg13g2_antennanp ANTENNA_2531 (.A(_07822_));
 sg13g2_antennanp ANTENNA_2532 (.A(_07835_));
 sg13g2_antennanp ANTENNA_2533 (.A(_07835_));
 sg13g2_antennanp ANTENNA_2534 (.A(_07914_));
 sg13g2_antennanp ANTENNA_2535 (.A(_07926_));
 sg13g2_antennanp ANTENNA_2536 (.A(_07939_));
 sg13g2_antennanp ANTENNA_2537 (.A(_07939_));
 sg13g2_antennanp ANTENNA_2538 (.A(_07952_));
 sg13g2_antennanp ANTENNA_2539 (.A(_08169_));
 sg13g2_antennanp ANTENNA_2540 (.A(_08169_));
 sg13g2_antennanp ANTENNA_2541 (.A(_09280_));
 sg13g2_antennanp ANTENNA_2542 (.A(_09280_));
 sg13g2_antennanp ANTENNA_2543 (.A(_09280_));
 sg13g2_antennanp ANTENNA_2544 (.A(_09280_));
 sg13g2_antennanp ANTENNA_2545 (.A(_09280_));
 sg13g2_antennanp ANTENNA_2546 (.A(_09724_));
 sg13g2_antennanp ANTENNA_2547 (.A(_09825_));
 sg13g2_antennanp ANTENNA_2548 (.A(_09825_));
 sg13g2_antennanp ANTENNA_2549 (.A(_09825_));
 sg13g2_antennanp ANTENNA_2550 (.A(_10247_));
 sg13g2_antennanp ANTENNA_2551 (.A(_10247_));
 sg13g2_antennanp ANTENNA_2552 (.A(_10247_));
 sg13g2_antennanp ANTENNA_2553 (.A(_10518_));
 sg13g2_antennanp ANTENNA_2554 (.A(_10604_));
 sg13g2_antennanp ANTENNA_2555 (.A(_10604_));
 sg13g2_antennanp ANTENNA_2556 (.A(_10604_));
 sg13g2_antennanp ANTENNA_2557 (.A(_10604_));
 sg13g2_antennanp ANTENNA_2558 (.A(_10617_));
 sg13g2_antennanp ANTENNA_2559 (.A(_10952_));
 sg13g2_antennanp ANTENNA_2560 (.A(_10963_));
 sg13g2_antennanp ANTENNA_2561 (.A(_11000_));
 sg13g2_antennanp ANTENNA_2562 (.A(_11000_));
 sg13g2_antennanp ANTENNA_2563 (.A(_11000_));
 sg13g2_antennanp ANTENNA_2564 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2565 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2566 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2567 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2568 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2569 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2570 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2571 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2572 (.A(_11243_));
 sg13g2_antennanp ANTENNA_2573 (.A(\top_ihp.oisc.op_a[22] ));
 sg13g2_antennanp ANTENNA_2574 (.A(\top_ihp.oisc.op_a[27] ));
 sg13g2_antennanp ANTENNA_2575 (.A(\top_ihp.oisc.op_a[6] ));
 sg13g2_antennanp ANTENNA_2576 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_2577 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_2578 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_2579 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_2580 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_2581 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_2582 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_2583 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_2584 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_2585 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_2586 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_2587 (.A(\top_ihp.oisc.regs[32][16] ));
 sg13g2_antennanp ANTENNA_2588 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_2589 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_2590 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_2591 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_2592 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_2593 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_2594 (.A(\top_ihp.oisc.regs[32][29] ));
 sg13g2_antennanp ANTENNA_2595 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_2596 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_2597 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_2598 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_2599 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_2600 (.A(\top_ihp.oisc.regs[63][5] ));
 sg13g2_antennanp ANTENNA_2601 (.A(\top_ihp.tx ));
 sg13g2_antennanp ANTENNA_2602 (.A(net1));
 sg13g2_antennanp ANTENNA_2603 (.A(net1));
 sg13g2_antennanp ANTENNA_2604 (.A(net1));
 sg13g2_antennanp ANTENNA_2605 (.A(net1));
 sg13g2_antennanp ANTENNA_2606 (.A(net5));
 sg13g2_antennanp ANTENNA_2607 (.A(net10));
 sg13g2_antennanp ANTENNA_2608 (.A(net77));
 sg13g2_antennanp ANTENNA_2609 (.A(net77));
 sg13g2_antennanp ANTENNA_2610 (.A(net77));
 sg13g2_antennanp ANTENNA_2611 (.A(net77));
 sg13g2_antennanp ANTENNA_2612 (.A(net77));
 sg13g2_antennanp ANTENNA_2613 (.A(net77));
 sg13g2_antennanp ANTENNA_2614 (.A(net77));
 sg13g2_antennanp ANTENNA_2615 (.A(net77));
 sg13g2_antennanp ANTENNA_2616 (.A(net91));
 sg13g2_antennanp ANTENNA_2617 (.A(net91));
 sg13g2_antennanp ANTENNA_2618 (.A(net91));
 sg13g2_antennanp ANTENNA_2619 (.A(net91));
 sg13g2_antennanp ANTENNA_2620 (.A(net91));
 sg13g2_antennanp ANTENNA_2621 (.A(net91));
 sg13g2_antennanp ANTENNA_2622 (.A(net91));
 sg13g2_antennanp ANTENNA_2623 (.A(net91));
 sg13g2_antennanp ANTENNA_2624 (.A(net91));
 sg13g2_antennanp ANTENNA_2625 (.A(net91));
 sg13g2_antennanp ANTENNA_2626 (.A(net91));
 sg13g2_antennanp ANTENNA_2627 (.A(net91));
 sg13g2_antennanp ANTENNA_2628 (.A(net91));
 sg13g2_antennanp ANTENNA_2629 (.A(net91));
 sg13g2_antennanp ANTENNA_2630 (.A(net146));
 sg13g2_antennanp ANTENNA_2631 (.A(net146));
 sg13g2_antennanp ANTENNA_2632 (.A(net146));
 sg13g2_antennanp ANTENNA_2633 (.A(net146));
 sg13g2_antennanp ANTENNA_2634 (.A(net146));
 sg13g2_antennanp ANTENNA_2635 (.A(net146));
 sg13g2_antennanp ANTENNA_2636 (.A(net146));
 sg13g2_antennanp ANTENNA_2637 (.A(net146));
 sg13g2_antennanp ANTENNA_2638 (.A(net146));
 sg13g2_antennanp ANTENNA_2639 (.A(net146));
 sg13g2_antennanp ANTENNA_2640 (.A(net146));
 sg13g2_antennanp ANTENNA_2641 (.A(net146));
 sg13g2_antennanp ANTENNA_2642 (.A(net155));
 sg13g2_antennanp ANTENNA_2643 (.A(net155));
 sg13g2_antennanp ANTENNA_2644 (.A(net155));
 sg13g2_antennanp ANTENNA_2645 (.A(net155));
 sg13g2_antennanp ANTENNA_2646 (.A(net155));
 sg13g2_antennanp ANTENNA_2647 (.A(net155));
 sg13g2_antennanp ANTENNA_2648 (.A(net155));
 sg13g2_antennanp ANTENNA_2649 (.A(net155));
 sg13g2_antennanp ANTENNA_2650 (.A(net155));
 sg13g2_antennanp ANTENNA_2651 (.A(net155));
 sg13g2_antennanp ANTENNA_2652 (.A(net155));
 sg13g2_antennanp ANTENNA_2653 (.A(net292));
 sg13g2_antennanp ANTENNA_2654 (.A(net292));
 sg13g2_antennanp ANTENNA_2655 (.A(net292));
 sg13g2_antennanp ANTENNA_2656 (.A(net292));
 sg13g2_antennanp ANTENNA_2657 (.A(net292));
 sg13g2_antennanp ANTENNA_2658 (.A(net292));
 sg13g2_antennanp ANTENNA_2659 (.A(net292));
 sg13g2_antennanp ANTENNA_2660 (.A(net292));
 sg13g2_antennanp ANTENNA_2661 (.A(net292));
 sg13g2_antennanp ANTENNA_2662 (.A(net317));
 sg13g2_antennanp ANTENNA_2663 (.A(net317));
 sg13g2_antennanp ANTENNA_2664 (.A(net317));
 sg13g2_antennanp ANTENNA_2665 (.A(net317));
 sg13g2_antennanp ANTENNA_2666 (.A(net317));
 sg13g2_antennanp ANTENNA_2667 (.A(net317));
 sg13g2_antennanp ANTENNA_2668 (.A(net317));
 sg13g2_antennanp ANTENNA_2669 (.A(net317));
 sg13g2_antennanp ANTENNA_2670 (.A(net317));
 sg13g2_antennanp ANTENNA_2671 (.A(net317));
 sg13g2_antennanp ANTENNA_2672 (.A(net317));
 sg13g2_antennanp ANTENNA_2673 (.A(net317));
 sg13g2_antennanp ANTENNA_2674 (.A(net397));
 sg13g2_antennanp ANTENNA_2675 (.A(net397));
 sg13g2_antennanp ANTENNA_2676 (.A(net397));
 sg13g2_antennanp ANTENNA_2677 (.A(net397));
 sg13g2_antennanp ANTENNA_2678 (.A(net397));
 sg13g2_antennanp ANTENNA_2679 (.A(net397));
 sg13g2_antennanp ANTENNA_2680 (.A(net397));
 sg13g2_antennanp ANTENNA_2681 (.A(net397));
 sg13g2_antennanp ANTENNA_2682 (.A(net397));
 sg13g2_antennanp ANTENNA_2683 (.A(net397));
 sg13g2_antennanp ANTENNA_2684 (.A(net397));
 sg13g2_antennanp ANTENNA_2685 (.A(net397));
 sg13g2_antennanp ANTENNA_2686 (.A(net397));
 sg13g2_antennanp ANTENNA_2687 (.A(net498));
 sg13g2_antennanp ANTENNA_2688 (.A(net498));
 sg13g2_antennanp ANTENNA_2689 (.A(net498));
 sg13g2_antennanp ANTENNA_2690 (.A(net498));
 sg13g2_antennanp ANTENNA_2691 (.A(net498));
 sg13g2_antennanp ANTENNA_2692 (.A(net498));
 sg13g2_antennanp ANTENNA_2693 (.A(net498));
 sg13g2_antennanp ANTENNA_2694 (.A(net498));
 sg13g2_antennanp ANTENNA_2695 (.A(net498));
 sg13g2_antennanp ANTENNA_2696 (.A(net525));
 sg13g2_antennanp ANTENNA_2697 (.A(net525));
 sg13g2_antennanp ANTENNA_2698 (.A(net525));
 sg13g2_antennanp ANTENNA_2699 (.A(net525));
 sg13g2_antennanp ANTENNA_2700 (.A(net525));
 sg13g2_antennanp ANTENNA_2701 (.A(net525));
 sg13g2_antennanp ANTENNA_2702 (.A(net525));
 sg13g2_antennanp ANTENNA_2703 (.A(net525));
 sg13g2_antennanp ANTENNA_2704 (.A(net525));
 sg13g2_antennanp ANTENNA_2705 (.A(net525));
 sg13g2_antennanp ANTENNA_2706 (.A(net525));
 sg13g2_antennanp ANTENNA_2707 (.A(net803));
 sg13g2_antennanp ANTENNA_2708 (.A(net803));
 sg13g2_antennanp ANTENNA_2709 (.A(net803));
 sg13g2_antennanp ANTENNA_2710 (.A(net803));
 sg13g2_antennanp ANTENNA_2711 (.A(net803));
 sg13g2_antennanp ANTENNA_2712 (.A(net803));
 sg13g2_antennanp ANTENNA_2713 (.A(net803));
 sg13g2_antennanp ANTENNA_2714 (.A(net803));
 sg13g2_antennanp ANTENNA_2715 (.A(net803));
 sg13g2_antennanp ANTENNA_2716 (.A(net1207));
 sg13g2_antennanp ANTENNA_2717 (.A(net1207));
 sg13g2_antennanp ANTENNA_2718 (.A(net1207));
 sg13g2_antennanp ANTENNA_2719 (.A(net1207));
 sg13g2_antennanp ANTENNA_2720 (.A(net1207));
 sg13g2_antennanp ANTENNA_2721 (.A(net1207));
 sg13g2_antennanp ANTENNA_2722 (.A(net1207));
 sg13g2_antennanp ANTENNA_2723 (.A(net1430));
 sg13g2_antennanp ANTENNA_2724 (.A(net1430));
 sg13g2_antennanp ANTENNA_2725 (.A(net1430));
 sg13g2_antennanp ANTENNA_2726 (.A(net1430));
 sg13g2_antennanp ANTENNA_2727 (.A(net1430));
 sg13g2_antennanp ANTENNA_2728 (.A(net1430));
 sg13g2_antennanp ANTENNA_2729 (.A(net1430));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_4 FILLER_0_175 ();
 sg13g2_fill_1 FILLER_0_179 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_decap_8 FILLER_0_213 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_fill_2 FILLER_0_227 ();
 sg13g2_fill_1 FILLER_0_229 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_decap_8 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_270 ();
 sg13g2_fill_2 FILLER_0_277 ();
 sg13g2_fill_1 FILLER_0_279 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_313 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_decap_4 FILLER_0_327 ();
 sg13g2_fill_1 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_decap_4 FILLER_0_407 ();
 sg13g2_fill_2 FILLER_0_411 ();
 sg13g2_decap_8 FILLER_0_423 ();
 sg13g2_decap_8 FILLER_0_430 ();
 sg13g2_fill_2 FILLER_0_437 ();
 sg13g2_fill_1 FILLER_0_439 ();
 sg13g2_fill_1 FILLER_0_445 ();
 sg13g2_decap_8 FILLER_0_456 ();
 sg13g2_decap_8 FILLER_0_463 ();
 sg13g2_decap_8 FILLER_0_470 ();
 sg13g2_decap_8 FILLER_0_477 ();
 sg13g2_fill_2 FILLER_0_484 ();
 sg13g2_decap_8 FILLER_0_512 ();
 sg13g2_decap_8 FILLER_0_519 ();
 sg13g2_decap_8 FILLER_0_526 ();
 sg13g2_decap_8 FILLER_0_533 ();
 sg13g2_decap_8 FILLER_0_540 ();
 sg13g2_decap_8 FILLER_0_547 ();
 sg13g2_decap_8 FILLER_0_554 ();
 sg13g2_decap_8 FILLER_0_561 ();
 sg13g2_decap_8 FILLER_0_568 ();
 sg13g2_decap_8 FILLER_0_575 ();
 sg13g2_decap_8 FILLER_0_582 ();
 sg13g2_fill_1 FILLER_0_589 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_fill_2 FILLER_0_609 ();
 sg13g2_fill_1 FILLER_0_611 ();
 sg13g2_decap_8 FILLER_0_638 ();
 sg13g2_decap_8 FILLER_0_645 ();
 sg13g2_decap_8 FILLER_0_652 ();
 sg13g2_decap_8 FILLER_0_659 ();
 sg13g2_decap_8 FILLER_0_666 ();
 sg13g2_decap_4 FILLER_0_673 ();
 sg13g2_fill_1 FILLER_0_677 ();
 sg13g2_decap_8 FILLER_0_704 ();
 sg13g2_decap_4 FILLER_0_711 ();
 sg13g2_decap_4 FILLER_0_745 ();
 sg13g2_fill_2 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_785 ();
 sg13g2_decap_8 FILLER_0_792 ();
 sg13g2_decap_8 FILLER_0_799 ();
 sg13g2_decap_8 FILLER_0_806 ();
 sg13g2_decap_4 FILLER_0_813 ();
 sg13g2_fill_1 FILLER_0_817 ();
 sg13g2_decap_4 FILLER_0_822 ();
 sg13g2_fill_1 FILLER_0_856 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_fill_2 FILLER_0_896 ();
 sg13g2_fill_1 FILLER_0_898 ();
 sg13g2_decap_8 FILLER_0_929 ();
 sg13g2_decap_8 FILLER_0_936 ();
 sg13g2_decap_8 FILLER_0_943 ();
 sg13g2_fill_2 FILLER_0_950 ();
 sg13g2_fill_1 FILLER_0_952 ();
 sg13g2_fill_1 FILLER_0_957 ();
 sg13g2_decap_8 FILLER_0_962 ();
 sg13g2_decap_8 FILLER_0_969 ();
 sg13g2_decap_8 FILLER_0_976 ();
 sg13g2_decap_8 FILLER_0_983 ();
 sg13g2_decap_8 FILLER_0_990 ();
 sg13g2_decap_8 FILLER_0_997 ();
 sg13g2_decap_8 FILLER_0_1004 ();
 sg13g2_decap_8 FILLER_0_1011 ();
 sg13g2_decap_8 FILLER_0_1018 ();
 sg13g2_decap_4 FILLER_0_1025 ();
 sg13g2_decap_8 FILLER_0_1033 ();
 sg13g2_decap_8 FILLER_0_1040 ();
 sg13g2_decap_8 FILLER_0_1047 ();
 sg13g2_decap_8 FILLER_0_1054 ();
 sg13g2_decap_8 FILLER_0_1061 ();
 sg13g2_fill_2 FILLER_0_1068 ();
 sg13g2_fill_1 FILLER_0_1070 ();
 sg13g2_decap_4 FILLER_0_1075 ();
 sg13g2_fill_2 FILLER_0_1079 ();
 sg13g2_decap_8 FILLER_0_1107 ();
 sg13g2_decap_8 FILLER_0_1114 ();
 sg13g2_decap_8 FILLER_0_1121 ();
 sg13g2_decap_8 FILLER_0_1128 ();
 sg13g2_decap_8 FILLER_0_1135 ();
 sg13g2_decap_8 FILLER_0_1142 ();
 sg13g2_decap_4 FILLER_0_1149 ();
 sg13g2_decap_8 FILLER_0_1179 ();
 sg13g2_decap_8 FILLER_0_1186 ();
 sg13g2_decap_8 FILLER_0_1193 ();
 sg13g2_decap_8 FILLER_0_1200 ();
 sg13g2_decap_8 FILLER_0_1207 ();
 sg13g2_decap_4 FILLER_0_1214 ();
 sg13g2_fill_1 FILLER_0_1218 ();
 sg13g2_decap_8 FILLER_0_1223 ();
 sg13g2_decap_8 FILLER_0_1260 ();
 sg13g2_decap_8 FILLER_0_1267 ();
 sg13g2_decap_8 FILLER_0_1274 ();
 sg13g2_decap_8 FILLER_0_1281 ();
 sg13g2_decap_4 FILLER_0_1288 ();
 sg13g2_fill_1 FILLER_0_1292 ();
 sg13g2_decap_8 FILLER_0_1323 ();
 sg13g2_decap_8 FILLER_0_1330 ();
 sg13g2_decap_8 FILLER_0_1337 ();
 sg13g2_decap_8 FILLER_0_1344 ();
 sg13g2_decap_8 FILLER_0_1351 ();
 sg13g2_decap_8 FILLER_0_1358 ();
 sg13g2_decap_8 FILLER_0_1365 ();
 sg13g2_decap_8 FILLER_0_1372 ();
 sg13g2_decap_8 FILLER_0_1379 ();
 sg13g2_decap_8 FILLER_0_1386 ();
 sg13g2_decap_8 FILLER_0_1393 ();
 sg13g2_fill_2 FILLER_0_1400 ();
 sg13g2_fill_1 FILLER_0_1402 ();
 sg13g2_decap_8 FILLER_0_1438 ();
 sg13g2_fill_2 FILLER_0_1445 ();
 sg13g2_fill_1 FILLER_0_1447 ();
 sg13g2_decap_8 FILLER_0_1474 ();
 sg13g2_decap_4 FILLER_0_1481 ();
 sg13g2_decap_8 FILLER_0_1511 ();
 sg13g2_decap_8 FILLER_0_1518 ();
 sg13g2_decap_8 FILLER_0_1525 ();
 sg13g2_decap_8 FILLER_0_1532 ();
 sg13g2_decap_8 FILLER_0_1539 ();
 sg13g2_decap_8 FILLER_0_1546 ();
 sg13g2_decap_8 FILLER_0_1553 ();
 sg13g2_decap_8 FILLER_0_1560 ();
 sg13g2_decap_8 FILLER_0_1567 ();
 sg13g2_decap_8 FILLER_0_1574 ();
 sg13g2_decap_8 FILLER_0_1581 ();
 sg13g2_fill_2 FILLER_0_1588 ();
 sg13g2_decap_8 FILLER_0_1620 ();
 sg13g2_decap_4 FILLER_0_1657 ();
 sg13g2_fill_2 FILLER_0_1661 ();
 sg13g2_decap_8 FILLER_0_1684 ();
 sg13g2_decap_8 FILLER_0_1691 ();
 sg13g2_fill_2 FILLER_0_1698 ();
 sg13g2_fill_1 FILLER_0_1700 ();
 sg13g2_fill_1 FILLER_0_1716 ();
 sg13g2_fill_1 FILLER_0_1727 ();
 sg13g2_decap_8 FILLER_0_1747 ();
 sg13g2_decap_8 FILLER_0_1754 ();
 sg13g2_decap_8 FILLER_0_1761 ();
 sg13g2_decap_4 FILLER_0_1768 ();
 sg13g2_fill_1 FILLER_0_1772 ();
 sg13g2_decap_8 FILLER_0_1777 ();
 sg13g2_decap_8 FILLER_0_1784 ();
 sg13g2_decap_8 FILLER_0_1791 ();
 sg13g2_decap_8 FILLER_0_1798 ();
 sg13g2_decap_8 FILLER_0_1805 ();
 sg13g2_decap_8 FILLER_0_1812 ();
 sg13g2_decap_8 FILLER_0_1819 ();
 sg13g2_decap_8 FILLER_0_1826 ();
 sg13g2_decap_8 FILLER_0_1833 ();
 sg13g2_decap_8 FILLER_0_1840 ();
 sg13g2_decap_8 FILLER_0_1847 ();
 sg13g2_decap_8 FILLER_0_1854 ();
 sg13g2_decap_8 FILLER_0_1861 ();
 sg13g2_decap_8 FILLER_0_1868 ();
 sg13g2_decap_8 FILLER_0_1875 ();
 sg13g2_decap_8 FILLER_0_1882 ();
 sg13g2_decap_8 FILLER_0_1889 ();
 sg13g2_decap_8 FILLER_0_1896 ();
 sg13g2_decap_8 FILLER_0_1903 ();
 sg13g2_decap_8 FILLER_0_1910 ();
 sg13g2_decap_8 FILLER_0_1917 ();
 sg13g2_decap_8 FILLER_0_1924 ();
 sg13g2_decap_8 FILLER_0_1931 ();
 sg13g2_decap_8 FILLER_0_1938 ();
 sg13g2_decap_8 FILLER_0_1945 ();
 sg13g2_decap_8 FILLER_0_1952 ();
 sg13g2_decap_8 FILLER_0_1959 ();
 sg13g2_decap_8 FILLER_0_1966 ();
 sg13g2_decap_8 FILLER_0_1973 ();
 sg13g2_decap_8 FILLER_0_1980 ();
 sg13g2_decap_8 FILLER_0_1987 ();
 sg13g2_decap_8 FILLER_0_1994 ();
 sg13g2_decap_8 FILLER_0_2001 ();
 sg13g2_decap_8 FILLER_0_2008 ();
 sg13g2_decap_8 FILLER_0_2015 ();
 sg13g2_decap_8 FILLER_0_2022 ();
 sg13g2_decap_8 FILLER_0_2029 ();
 sg13g2_decap_8 FILLER_0_2036 ();
 sg13g2_decap_8 FILLER_0_2043 ();
 sg13g2_decap_8 FILLER_0_2050 ();
 sg13g2_decap_8 FILLER_0_2057 ();
 sg13g2_fill_2 FILLER_0_2064 ();
 sg13g2_fill_1 FILLER_0_2066 ();
 sg13g2_decap_8 FILLER_0_2071 ();
 sg13g2_decap_8 FILLER_0_2078 ();
 sg13g2_fill_2 FILLER_0_2085 ();
 sg13g2_fill_1 FILLER_0_2087 ();
 sg13g2_decap_8 FILLER_0_2092 ();
 sg13g2_decap_8 FILLER_0_2099 ();
 sg13g2_decap_4 FILLER_0_2106 ();
 sg13g2_decap_8 FILLER_0_2166 ();
 sg13g2_decap_8 FILLER_0_2173 ();
 sg13g2_decap_8 FILLER_0_2180 ();
 sg13g2_decap_8 FILLER_0_2187 ();
 sg13g2_decap_8 FILLER_0_2194 ();
 sg13g2_decap_8 FILLER_0_2201 ();
 sg13g2_decap_8 FILLER_0_2208 ();
 sg13g2_decap_8 FILLER_0_2215 ();
 sg13g2_decap_8 FILLER_0_2222 ();
 sg13g2_decap_8 FILLER_0_2229 ();
 sg13g2_decap_8 FILLER_0_2236 ();
 sg13g2_decap_8 FILLER_0_2243 ();
 sg13g2_decap_8 FILLER_0_2250 ();
 sg13g2_decap_8 FILLER_0_2257 ();
 sg13g2_decap_8 FILLER_0_2264 ();
 sg13g2_decap_8 FILLER_0_2271 ();
 sg13g2_decap_8 FILLER_0_2278 ();
 sg13g2_decap_8 FILLER_0_2285 ();
 sg13g2_decap_4 FILLER_0_2292 ();
 sg13g2_decap_8 FILLER_0_2303 ();
 sg13g2_decap_8 FILLER_0_2310 ();
 sg13g2_decap_8 FILLER_0_2317 ();
 sg13g2_decap_8 FILLER_0_2324 ();
 sg13g2_decap_8 FILLER_0_2331 ();
 sg13g2_decap_8 FILLER_0_2338 ();
 sg13g2_decap_8 FILLER_0_2345 ();
 sg13g2_decap_8 FILLER_0_2352 ();
 sg13g2_decap_8 FILLER_0_2359 ();
 sg13g2_decap_4 FILLER_0_2366 ();
 sg13g2_decap_8 FILLER_0_2374 ();
 sg13g2_decap_8 FILLER_0_2381 ();
 sg13g2_decap_8 FILLER_0_2388 ();
 sg13g2_decap_8 FILLER_0_2395 ();
 sg13g2_decap_8 FILLER_0_2402 ();
 sg13g2_decap_8 FILLER_0_2435 ();
 sg13g2_decap_8 FILLER_0_2442 ();
 sg13g2_decap_8 FILLER_0_2449 ();
 sg13g2_decap_8 FILLER_0_2456 ();
 sg13g2_decap_8 FILLER_0_2463 ();
 sg13g2_decap_8 FILLER_0_2470 ();
 sg13g2_decap_8 FILLER_0_2477 ();
 sg13g2_decap_8 FILLER_0_2484 ();
 sg13g2_decap_8 FILLER_0_2491 ();
 sg13g2_decap_8 FILLER_0_2498 ();
 sg13g2_decap_8 FILLER_0_2505 ();
 sg13g2_decap_4 FILLER_0_2516 ();
 sg13g2_fill_2 FILLER_0_2520 ();
 sg13g2_decap_8 FILLER_0_2526 ();
 sg13g2_decap_8 FILLER_0_2533 ();
 sg13g2_decap_8 FILLER_0_2540 ();
 sg13g2_decap_8 FILLER_0_2547 ();
 sg13g2_decap_8 FILLER_0_2554 ();
 sg13g2_decap_8 FILLER_0_2561 ();
 sg13g2_decap_8 FILLER_0_2568 ();
 sg13g2_decap_8 FILLER_0_2575 ();
 sg13g2_decap_8 FILLER_0_2582 ();
 sg13g2_decap_8 FILLER_0_2589 ();
 sg13g2_decap_8 FILLER_0_2596 ();
 sg13g2_decap_8 FILLER_0_2603 ();
 sg13g2_decap_8 FILLER_0_2610 ();
 sg13g2_decap_8 FILLER_0_2617 ();
 sg13g2_decap_8 FILLER_0_2624 ();
 sg13g2_decap_8 FILLER_0_2631 ();
 sg13g2_decap_8 FILLER_0_2638 ();
 sg13g2_decap_8 FILLER_0_2645 ();
 sg13g2_decap_8 FILLER_0_2652 ();
 sg13g2_decap_8 FILLER_0_2659 ();
 sg13g2_decap_4 FILLER_0_2666 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_4 FILLER_1_56 ();
 sg13g2_decap_4 FILLER_1_86 ();
 sg13g2_decap_8 FILLER_1_142 ();
 sg13g2_decap_8 FILLER_1_149 ();
 sg13g2_decap_8 FILLER_1_156 ();
 sg13g2_decap_8 FILLER_1_163 ();
 sg13g2_decap_4 FILLER_1_170 ();
 sg13g2_fill_1 FILLER_1_174 ();
 sg13g2_fill_2 FILLER_1_211 ();
 sg13g2_fill_1 FILLER_1_213 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_fill_2 FILLER_1_231 ();
 sg13g2_fill_1 FILLER_1_233 ();
 sg13g2_decap_8 FILLER_1_260 ();
 sg13g2_decap_4 FILLER_1_267 ();
 sg13g2_fill_2 FILLER_1_271 ();
 sg13g2_decap_4 FILLER_1_283 ();
 sg13g2_fill_1 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_317 ();
 sg13g2_decap_8 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_fill_2 FILLER_1_391 ();
 sg13g2_fill_2 FILLER_1_419 ();
 sg13g2_fill_1 FILLER_1_421 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_decap_4 FILLER_1_439 ();
 sg13g2_fill_2 FILLER_1_448 ();
 sg13g2_decap_4 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_fill_2 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_fill_2 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_551 ();
 sg13g2_decap_8 FILLER_1_558 ();
 sg13g2_decap_4 FILLER_1_565 ();
 sg13g2_fill_2 FILLER_1_569 ();
 sg13g2_fill_2 FILLER_1_581 ();
 sg13g2_fill_2 FILLER_1_588 ();
 sg13g2_fill_1 FILLER_1_590 ();
 sg13g2_fill_1 FILLER_1_617 ();
 sg13g2_fill_1 FILLER_1_644 ();
 sg13g2_fill_2 FILLER_1_671 ();
 sg13g2_fill_1 FILLER_1_673 ();
 sg13g2_decap_4 FILLER_1_708 ();
 sg13g2_fill_1 FILLER_1_712 ();
 sg13g2_fill_1 FILLER_1_790 ();
 sg13g2_decap_4 FILLER_1_821 ();
 sg13g2_fill_2 FILLER_1_825 ();
 sg13g2_decap_4 FILLER_1_831 ();
 sg13g2_fill_2 FILLER_1_835 ();
 sg13g2_fill_2 FILLER_1_858 ();
 sg13g2_fill_1 FILLER_1_860 ();
 sg13g2_decap_8 FILLER_1_867 ();
 sg13g2_decap_4 FILLER_1_874 ();
 sg13g2_fill_2 FILLER_1_878 ();
 sg13g2_decap_8 FILLER_1_884 ();
 sg13g2_decap_8 FILLER_1_891 ();
 sg13g2_fill_2 FILLER_1_898 ();
 sg13g2_decap_8 FILLER_1_904 ();
 sg13g2_decap_8 FILLER_1_911 ();
 sg13g2_fill_2 FILLER_1_961 ();
 sg13g2_fill_1 FILLER_1_997 ();
 sg13g2_fill_2 FILLER_1_1050 ();
 sg13g2_fill_1 FILLER_1_1052 ();
 sg13g2_fill_2 FILLER_1_1079 ();
 sg13g2_fill_1 FILLER_1_1081 ();
 sg13g2_decap_8 FILLER_1_1116 ();
 sg13g2_fill_2 FILLER_1_1123 ();
 sg13g2_fill_1 FILLER_1_1125 ();
 sg13g2_fill_2 FILLER_1_1152 ();
 sg13g2_fill_1 FILLER_1_1206 ();
 sg13g2_decap_8 FILLER_1_1241 ();
 sg13g2_decap_8 FILLER_1_1248 ();
 sg13g2_decap_8 FILLER_1_1255 ();
 sg13g2_fill_1 FILLER_1_1262 ();
 sg13g2_fill_1 FILLER_1_1315 ();
 sg13g2_fill_1 FILLER_1_1342 ();
 sg13g2_fill_1 FILLER_1_1369 ();
 sg13g2_fill_1 FILLER_1_1396 ();
 sg13g2_decap_4 FILLER_1_1431 ();
 sg13g2_fill_1 FILLER_1_1435 ();
 sg13g2_fill_1 FILLER_1_1440 ();
 sg13g2_fill_1 FILLER_1_1445 ();
 sg13g2_fill_2 FILLER_1_1450 ();
 sg13g2_fill_2 FILLER_1_1478 ();
 sg13g2_decap_8 FILLER_1_1510 ();
 sg13g2_decap_4 FILLER_1_1517 ();
 sg13g2_fill_2 FILLER_1_1521 ();
 sg13g2_fill_2 FILLER_1_1553 ();
 sg13g2_fill_2 FILLER_1_1628 ();
 sg13g2_fill_1 FILLER_1_1630 ();
 sg13g2_decap_8 FILLER_1_1696 ();
 sg13g2_decap_4 FILLER_1_1703 ();
 sg13g2_fill_2 FILLER_1_1720 ();
 sg13g2_decap_8 FILLER_1_1748 ();
 sg13g2_decap_4 FILLER_1_1755 ();
 sg13g2_fill_2 FILLER_1_1841 ();
 sg13g2_decap_4 FILLER_1_1934 ();
 sg13g2_fill_1 FILLER_1_1938 ();
 sg13g2_fill_2 FILLER_1_1944 ();
 sg13g2_fill_1 FILLER_1_1946 ();
 sg13g2_fill_2 FILLER_1_1952 ();
 sg13g2_fill_1 FILLER_1_1954 ();
 sg13g2_decap_8 FILLER_1_1959 ();
 sg13g2_decap_4 FILLER_1_1966 ();
 sg13g2_fill_2 FILLER_1_1975 ();
 sg13g2_decap_8 FILLER_1_1981 ();
 sg13g2_decap_8 FILLER_1_1988 ();
 sg13g2_decap_4 FILLER_1_1999 ();
 sg13g2_fill_1 FILLER_1_2003 ();
 sg13g2_decap_8 FILLER_1_2030 ();
 sg13g2_decap_8 FILLER_1_2037 ();
 sg13g2_decap_8 FILLER_1_2044 ();
 sg13g2_decap_8 FILLER_1_2051 ();
 sg13g2_fill_2 FILLER_1_2114 ();
 sg13g2_fill_1 FILLER_1_2116 ();
 sg13g2_fill_1 FILLER_1_2138 ();
 sg13g2_decap_8 FILLER_1_2174 ();
 sg13g2_decap_8 FILLER_1_2181 ();
 sg13g2_fill_2 FILLER_1_2188 ();
 sg13g2_fill_2 FILLER_1_2195 ();
 sg13g2_fill_1 FILLER_1_2197 ();
 sg13g2_decap_8 FILLER_1_2224 ();
 sg13g2_fill_2 FILLER_1_2231 ();
 sg13g2_decap_4 FILLER_1_2267 ();
 sg13g2_decap_8 FILLER_1_2275 ();
 sg13g2_fill_2 FILLER_1_2282 ();
 sg13g2_fill_1 FILLER_1_2284 ();
 sg13g2_decap_4 FILLER_1_2353 ();
 sg13g2_fill_2 FILLER_1_2357 ();
 sg13g2_decap_4 FILLER_1_2389 ();
 sg13g2_decap_8 FILLER_1_2431 ();
 sg13g2_decap_4 FILLER_1_2438 ();
 sg13g2_fill_1 FILLER_1_2442 ();
 sg13g2_decap_8 FILLER_1_2447 ();
 sg13g2_decap_8 FILLER_1_2454 ();
 sg13g2_fill_1 FILLER_1_2461 ();
 sg13g2_decap_8 FILLER_1_2540 ();
 sg13g2_decap_8 FILLER_1_2547 ();
 sg13g2_decap_8 FILLER_1_2584 ();
 sg13g2_decap_8 FILLER_1_2591 ();
 sg13g2_decap_8 FILLER_1_2598 ();
 sg13g2_decap_8 FILLER_1_2605 ();
 sg13g2_decap_8 FILLER_1_2612 ();
 sg13g2_decap_8 FILLER_1_2619 ();
 sg13g2_decap_8 FILLER_1_2626 ();
 sg13g2_decap_8 FILLER_1_2633 ();
 sg13g2_decap_8 FILLER_1_2640 ();
 sg13g2_decap_8 FILLER_1_2647 ();
 sg13g2_decap_8 FILLER_1_2654 ();
 sg13g2_decap_8 FILLER_1_2661 ();
 sg13g2_fill_2 FILLER_1_2668 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_4 FILLER_2_56 ();
 sg13g2_fill_1 FILLER_2_90 ();
 sg13g2_fill_2 FILLER_2_95 ();
 sg13g2_fill_1 FILLER_2_97 ();
 sg13g2_fill_2 FILLER_2_106 ();
 sg13g2_fill_2 FILLER_2_112 ();
 sg13g2_fill_1 FILLER_2_114 ();
 sg13g2_fill_1 FILLER_2_119 ();
 sg13g2_fill_2 FILLER_2_124 ();
 sg13g2_fill_1 FILLER_2_131 ();
 sg13g2_fill_2 FILLER_2_136 ();
 sg13g2_decap_8 FILLER_2_142 ();
 sg13g2_decap_8 FILLER_2_149 ();
 sg13g2_decap_8 FILLER_2_156 ();
 sg13g2_decap_8 FILLER_2_163 ();
 sg13g2_fill_2 FILLER_2_170 ();
 sg13g2_decap_8 FILLER_2_185 ();
 sg13g2_fill_2 FILLER_2_202 ();
 sg13g2_fill_2 FILLER_2_208 ();
 sg13g2_decap_8 FILLER_2_215 ();
 sg13g2_fill_1 FILLER_2_237 ();
 sg13g2_fill_1 FILLER_2_248 ();
 sg13g2_fill_1 FILLER_2_253 ();
 sg13g2_fill_1 FILLER_2_262 ();
 sg13g2_decap_4 FILLER_2_268 ();
 sg13g2_decap_4 FILLER_2_295 ();
 sg13g2_fill_2 FILLER_2_299 ();
 sg13g2_fill_1 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_316 ();
 sg13g2_fill_1 FILLER_2_323 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_fill_1 FILLER_2_446 ();
 sg13g2_fill_2 FILLER_2_478 ();
 sg13g2_fill_1 FILLER_2_480 ();
 sg13g2_decap_8 FILLER_2_521 ();
 sg13g2_fill_2 FILLER_2_528 ();
 sg13g2_fill_1 FILLER_2_530 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_fill_1 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_fill_2 FILLER_2_637 ();
 sg13g2_fill_1 FILLER_2_639 ();
 sg13g2_decap_8 FILLER_2_671 ();
 sg13g2_decap_8 FILLER_2_678 ();
 sg13g2_fill_1 FILLER_2_685 ();
 sg13g2_decap_8 FILLER_2_694 ();
 sg13g2_decap_8 FILLER_2_701 ();
 sg13g2_decap_8 FILLER_2_708 ();
 sg13g2_fill_1 FILLER_2_715 ();
 sg13g2_decap_4 FILLER_2_720 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_4 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_817 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_fill_2 FILLER_2_837 ();
 sg13g2_fill_1 FILLER_2_839 ();
 sg13g2_fill_1 FILLER_2_866 ();
 sg13g2_fill_1 FILLER_2_919 ();
 sg13g2_decap_4 FILLER_2_980 ();
 sg13g2_fill_1 FILLER_2_984 ();
 sg13g2_fill_2 FILLER_2_989 ();
 sg13g2_fill_1 FILLER_2_995 ();
 sg13g2_fill_2 FILLER_2_1078 ();
 sg13g2_fill_1 FILLER_2_1080 ();
 sg13g2_fill_2 FILLER_2_1102 ();
 sg13g2_fill_1 FILLER_2_1104 ();
 sg13g2_decap_8 FILLER_2_1131 ();
 sg13g2_decap_8 FILLER_2_1138 ();
 sg13g2_fill_1 FILLER_2_1145 ();
 sg13g2_fill_2 FILLER_2_1156 ();
 sg13g2_fill_1 FILLER_2_1158 ();
 sg13g2_fill_2 FILLER_2_1171 ();
 sg13g2_fill_1 FILLER_2_1173 ();
 sg13g2_fill_2 FILLER_2_1178 ();
 sg13g2_fill_1 FILLER_2_1210 ();
 sg13g2_fill_1 FILLER_2_1215 ();
 sg13g2_fill_1 FILLER_2_1246 ();
 sg13g2_fill_2 FILLER_2_1320 ();
 sg13g2_fill_1 FILLER_2_1326 ();
 sg13g2_fill_2 FILLER_2_1331 ();
 sg13g2_decap_8 FILLER_2_1343 ();
 sg13g2_decap_8 FILLER_2_1350 ();
 sg13g2_decap_8 FILLER_2_1357 ();
 sg13g2_decap_4 FILLER_2_1364 ();
 sg13g2_fill_1 FILLER_2_1372 ();
 sg13g2_fill_2 FILLER_2_1425 ();
 sg13g2_fill_2 FILLER_2_1453 ();
 sg13g2_decap_8 FILLER_2_1463 ();
 sg13g2_decap_8 FILLER_2_1470 ();
 sg13g2_fill_2 FILLER_2_1477 ();
 sg13g2_fill_1 FILLER_2_1479 ();
 sg13g2_fill_1 FILLER_2_1511 ();
 sg13g2_decap_8 FILLER_2_1576 ();
 sg13g2_fill_2 FILLER_2_1583 ();
 sg13g2_fill_2 FILLER_2_1593 ();
 sg13g2_fill_1 FILLER_2_1595 ();
 sg13g2_decap_4 FILLER_2_1626 ();
 sg13g2_fill_1 FILLER_2_1630 ();
 sg13g2_decap_8 FILLER_2_1643 ();
 sg13g2_decap_8 FILLER_2_1650 ();
 sg13g2_decap_8 FILLER_2_1657 ();
 sg13g2_decap_8 FILLER_2_1664 ();
 sg13g2_decap_4 FILLER_2_1671 ();
 sg13g2_fill_1 FILLER_2_1679 ();
 sg13g2_fill_1 FILLER_2_1723 ();
 sg13g2_decap_8 FILLER_2_1750 ();
 sg13g2_decap_8 FILLER_2_1757 ();
 sg13g2_decap_8 FILLER_2_1768 ();
 sg13g2_fill_2 FILLER_2_1775 ();
 sg13g2_fill_1 FILLER_2_1777 ();
 sg13g2_decap_8 FILLER_2_1804 ();
 sg13g2_decap_8 FILLER_2_1811 ();
 sg13g2_decap_4 FILLER_2_1818 ();
 sg13g2_decap_8 FILLER_2_1862 ();
 sg13g2_decap_8 FILLER_2_1869 ();
 sg13g2_fill_2 FILLER_2_1876 ();
 sg13g2_fill_1 FILLER_2_1878 ();
 sg13g2_decap_8 FILLER_2_1888 ();
 sg13g2_decap_8 FILLER_2_1895 ();
 sg13g2_decap_4 FILLER_2_1902 ();
 sg13g2_fill_1 FILLER_2_1967 ();
 sg13g2_fill_2 FILLER_2_2020 ();
 sg13g2_fill_1 FILLER_2_2022 ();
 sg13g2_decap_8 FILLER_2_2075 ();
 sg13g2_decap_8 FILLER_2_2082 ();
 sg13g2_decap_8 FILLER_2_2089 ();
 sg13g2_fill_2 FILLER_2_2113 ();
 sg13g2_fill_1 FILLER_2_2115 ();
 sg13g2_fill_2 FILLER_2_2289 ();
 sg13g2_fill_2 FILLER_2_2299 ();
 sg13g2_fill_1 FILLER_2_2305 ();
 sg13g2_fill_2 FILLER_2_2332 ();
 sg13g2_fill_2 FILLER_2_2338 ();
 sg13g2_fill_1 FILLER_2_2345 ();
 sg13g2_decap_8 FILLER_2_2372 ();
 sg13g2_fill_2 FILLER_2_2379 ();
 sg13g2_fill_1 FILLER_2_2381 ();
 sg13g2_decap_8 FILLER_2_2416 ();
 sg13g2_decap_8 FILLER_2_2423 ();
 sg13g2_fill_2 FILLER_2_2494 ();
 sg13g2_decap_4 FILLER_2_2500 ();
 sg13g2_fill_1 FILLER_2_2504 ();
 sg13g2_decap_4 FILLER_2_2531 ();
 sg13g2_fill_1 FILLER_2_2535 ();
 sg13g2_fill_2 FILLER_2_2562 ();
 sg13g2_fill_1 FILLER_2_2564 ();
 sg13g2_decap_8 FILLER_2_2569 ();
 sg13g2_decap_8 FILLER_2_2576 ();
 sg13g2_decap_8 FILLER_2_2583 ();
 sg13g2_decap_8 FILLER_2_2590 ();
 sg13g2_decap_8 FILLER_2_2597 ();
 sg13g2_decap_8 FILLER_2_2604 ();
 sg13g2_decap_8 FILLER_2_2611 ();
 sg13g2_decap_8 FILLER_2_2618 ();
 sg13g2_decap_8 FILLER_2_2625 ();
 sg13g2_decap_8 FILLER_2_2632 ();
 sg13g2_decap_8 FILLER_2_2639 ();
 sg13g2_decap_8 FILLER_2_2646 ();
 sg13g2_decap_8 FILLER_2_2653 ();
 sg13g2_decap_8 FILLER_2_2660 ();
 sg13g2_fill_2 FILLER_2_2667 ();
 sg13g2_fill_1 FILLER_2_2669 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_4 FILLER_3_35 ();
 sg13g2_decap_4 FILLER_3_43 ();
 sg13g2_decap_4 FILLER_3_91 ();
 sg13g2_fill_1 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_159 ();
 sg13g2_decap_8 FILLER_3_166 ();
 sg13g2_fill_2 FILLER_3_173 ();
 sg13g2_fill_1 FILLER_3_175 ();
 sg13g2_fill_2 FILLER_3_215 ();
 sg13g2_fill_1 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_4 FILLER_3_242 ();
 sg13g2_decap_4 FILLER_3_250 ();
 sg13g2_fill_1 FILLER_3_254 ();
 sg13g2_fill_2 FILLER_3_265 ();
 sg13g2_fill_1 FILLER_3_267 ();
 sg13g2_decap_8 FILLER_3_304 ();
 sg13g2_decap_8 FILLER_3_311 ();
 sg13g2_decap_8 FILLER_3_318 ();
 sg13g2_decap_8 FILLER_3_325 ();
 sg13g2_decap_8 FILLER_3_332 ();
 sg13g2_decap_8 FILLER_3_339 ();
 sg13g2_decap_8 FILLER_3_346 ();
 sg13g2_decap_8 FILLER_3_353 ();
 sg13g2_decap_8 FILLER_3_360 ();
 sg13g2_decap_4 FILLER_3_367 ();
 sg13g2_decap_4 FILLER_3_407 ();
 sg13g2_fill_1 FILLER_3_411 ();
 sg13g2_decap_4 FILLER_3_433 ();
 sg13g2_fill_2 FILLER_3_437 ();
 sg13g2_fill_2 FILLER_3_449 ();
 sg13g2_fill_2 FILLER_3_469 ();
 sg13g2_fill_1 FILLER_3_471 ();
 sg13g2_decap_4 FILLER_3_485 ();
 sg13g2_fill_1 FILLER_3_489 ();
 sg13g2_fill_2 FILLER_3_500 ();
 sg13g2_fill_1 FILLER_3_502 ();
 sg13g2_fill_2 FILLER_3_506 ();
 sg13g2_fill_1 FILLER_3_508 ();
 sg13g2_fill_1 FILLER_3_514 ();
 sg13g2_fill_1 FILLER_3_543 ();
 sg13g2_decap_8 FILLER_3_548 ();
 sg13g2_fill_2 FILLER_3_584 ();
 sg13g2_fill_2 FILLER_3_590 ();
 sg13g2_decap_8 FILLER_3_610 ();
 sg13g2_decap_8 FILLER_3_617 ();
 sg13g2_decap_8 FILLER_3_624 ();
 sg13g2_decap_8 FILLER_3_631 ();
 sg13g2_fill_2 FILLER_3_638 ();
 sg13g2_decap_8 FILLER_3_650 ();
 sg13g2_decap_8 FILLER_3_657 ();
 sg13g2_fill_1 FILLER_3_664 ();
 sg13g2_decap_8 FILLER_3_670 ();
 sg13g2_fill_2 FILLER_3_677 ();
 sg13g2_fill_1 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_688 ();
 sg13g2_decap_8 FILLER_3_695 ();
 sg13g2_fill_2 FILLER_3_702 ();
 sg13g2_fill_1 FILLER_3_736 ();
 sg13g2_fill_1 FILLER_3_741 ();
 sg13g2_decap_8 FILLER_3_748 ();
 sg13g2_decap_8 FILLER_3_755 ();
 sg13g2_decap_8 FILLER_3_762 ();
 sg13g2_decap_8 FILLER_3_769 ();
 sg13g2_decap_8 FILLER_3_776 ();
 sg13g2_fill_1 FILLER_3_783 ();
 sg13g2_fill_1 FILLER_3_820 ();
 sg13g2_decap_4 FILLER_3_907 ();
 sg13g2_decap_4 FILLER_3_915 ();
 sg13g2_fill_2 FILLER_3_925 ();
 sg13g2_fill_1 FILLER_3_927 ();
 sg13g2_decap_4 FILLER_3_936 ();
 sg13g2_fill_1 FILLER_3_940 ();
 sg13g2_fill_2 FILLER_3_947 ();
 sg13g2_fill_1 FILLER_3_975 ();
 sg13g2_fill_1 FILLER_3_1002 ();
 sg13g2_decap_8 FILLER_3_1015 ();
 sg13g2_decap_8 FILLER_3_1022 ();
 sg13g2_fill_1 FILLER_3_1029 ();
 sg13g2_decap_4 FILLER_3_1034 ();
 sg13g2_fill_1 FILLER_3_1047 ();
 sg13g2_fill_1 FILLER_3_1053 ();
 sg13g2_fill_1 FILLER_3_1080 ();
 sg13g2_fill_2 FILLER_3_1107 ();
 sg13g2_decap_8 FILLER_3_1114 ();
 sg13g2_decap_8 FILLER_3_1147 ();
 sg13g2_decap_8 FILLER_3_1154 ();
 sg13g2_fill_2 FILLER_3_1161 ();
 sg13g2_decap_8 FILLER_3_1176 ();
 sg13g2_fill_1 FILLER_3_1183 ();
 sg13g2_fill_2 FILLER_3_1236 ();
 sg13g2_decap_8 FILLER_3_1244 ();
 sg13g2_decap_4 FILLER_3_1251 ();
 sg13g2_fill_1 FILLER_3_1259 ();
 sg13g2_decap_8 FILLER_3_1264 ();
 sg13g2_fill_2 FILLER_3_1271 ();
 sg13g2_fill_1 FILLER_3_1277 ();
 sg13g2_fill_2 FILLER_3_1286 ();
 sg13g2_fill_1 FILLER_3_1288 ();
 sg13g2_decap_8 FILLER_3_1315 ();
 sg13g2_decap_8 FILLER_3_1322 ();
 sg13g2_decap_8 FILLER_3_1329 ();
 sg13g2_decap_8 FILLER_3_1367 ();
 sg13g2_fill_2 FILLER_3_1374 ();
 sg13g2_decap_4 FILLER_3_1380 ();
 sg13g2_decap_8 FILLER_3_1388 ();
 sg13g2_decap_4 FILLER_3_1395 ();
 sg13g2_decap_8 FILLER_3_1429 ();
 sg13g2_decap_8 FILLER_3_1436 ();
 sg13g2_decap_8 FILLER_3_1449 ();
 sg13g2_decap_8 FILLER_3_1456 ();
 sg13g2_decap_8 FILLER_3_1463 ();
 sg13g2_decap_4 FILLER_3_1470 ();
 sg13g2_fill_2 FILLER_3_1474 ();
 sg13g2_decap_8 FILLER_3_1506 ();
 sg13g2_decap_4 FILLER_3_1513 ();
 sg13g2_decap_4 FILLER_3_1547 ();
 sg13g2_decap_4 FILLER_3_1559 ();
 sg13g2_decap_8 FILLER_3_1567 ();
 sg13g2_decap_8 FILLER_3_1574 ();
 sg13g2_decap_8 FILLER_3_1581 ();
 sg13g2_decap_8 FILLER_3_1588 ();
 sg13g2_decap_8 FILLER_3_1595 ();
 sg13g2_decap_8 FILLER_3_1602 ();
 sg13g2_fill_1 FILLER_3_1609 ();
 sg13g2_decap_8 FILLER_3_1627 ();
 sg13g2_decap_4 FILLER_3_1634 ();
 sg13g2_fill_1 FILLER_3_1638 ();
 sg13g2_fill_1 FILLER_3_1652 ();
 sg13g2_decap_8 FILLER_3_1666 ();
 sg13g2_decap_8 FILLER_3_1673 ();
 sg13g2_fill_2 FILLER_3_1680 ();
 sg13g2_fill_2 FILLER_3_1708 ();
 sg13g2_fill_1 FILLER_3_1710 ();
 sg13g2_fill_2 FILLER_3_1715 ();
 sg13g2_fill_1 FILLER_3_1717 ();
 sg13g2_fill_2 FILLER_3_1724 ();
 sg13g2_fill_1 FILLER_3_1756 ();
 sg13g2_decap_8 FILLER_3_1761 ();
 sg13g2_decap_8 FILLER_3_1768 ();
 sg13g2_decap_8 FILLER_3_1810 ();
 sg13g2_fill_2 FILLER_3_1817 ();
 sg13g2_decap_4 FILLER_3_1845 ();
 sg13g2_fill_1 FILLER_3_1881 ();
 sg13g2_decap_8 FILLER_3_1908 ();
 sg13g2_fill_2 FILLER_3_1915 ();
 sg13g2_fill_1 FILLER_3_1917 ();
 sg13g2_decap_8 FILLER_3_2096 ();
 sg13g2_decap_8 FILLER_3_2103 ();
 sg13g2_decap_8 FILLER_3_2110 ();
 sg13g2_fill_2 FILLER_3_2117 ();
 sg13g2_fill_1 FILLER_3_2119 ();
 sg13g2_decap_8 FILLER_3_2125 ();
 sg13g2_decap_4 FILLER_3_2132 ();
 sg13g2_fill_2 FILLER_3_2136 ();
 sg13g2_decap_8 FILLER_3_2143 ();
 sg13g2_decap_8 FILLER_3_2150 ();
 sg13g2_decap_4 FILLER_3_2157 ();
 sg13g2_fill_1 FILLER_3_2161 ();
 sg13g2_fill_1 FILLER_3_2171 ();
 sg13g2_decap_4 FILLER_3_2176 ();
 sg13g2_fill_2 FILLER_3_2180 ();
 sg13g2_fill_1 FILLER_3_2212 ();
 sg13g2_decap_8 FILLER_3_2217 ();
 sg13g2_fill_1 FILLER_3_2238 ();
 sg13g2_fill_2 FILLER_3_2279 ();
 sg13g2_fill_1 FILLER_3_2281 ();
 sg13g2_fill_2 FILLER_3_2308 ();
 sg13g2_fill_2 FILLER_3_2314 ();
 sg13g2_decap_4 FILLER_3_2320 ();
 sg13g2_fill_1 FILLER_3_2324 ();
 sg13g2_fill_2 FILLER_3_2364 ();
 sg13g2_fill_1 FILLER_3_2366 ();
 sg13g2_fill_1 FILLER_3_2406 ();
 sg13g2_decap_8 FILLER_3_2433 ();
 sg13g2_decap_8 FILLER_3_2440 ();
 sg13g2_decap_8 FILLER_3_2447 ();
 sg13g2_fill_2 FILLER_3_2454 ();
 sg13g2_fill_1 FILLER_3_2456 ();
 sg13g2_decap_8 FILLER_3_2510 ();
 sg13g2_decap_8 FILLER_3_2517 ();
 sg13g2_decap_4 FILLER_3_2524 ();
 sg13g2_fill_1 FILLER_3_2528 ();
 sg13g2_decap_8 FILLER_3_2568 ();
 sg13g2_decap_8 FILLER_3_2575 ();
 sg13g2_decap_8 FILLER_3_2582 ();
 sg13g2_decap_8 FILLER_3_2589 ();
 sg13g2_decap_8 FILLER_3_2596 ();
 sg13g2_decap_8 FILLER_3_2603 ();
 sg13g2_decap_8 FILLER_3_2610 ();
 sg13g2_decap_8 FILLER_3_2617 ();
 sg13g2_decap_8 FILLER_3_2624 ();
 sg13g2_decap_8 FILLER_3_2631 ();
 sg13g2_decap_8 FILLER_3_2638 ();
 sg13g2_decap_8 FILLER_3_2645 ();
 sg13g2_decap_8 FILLER_3_2652 ();
 sg13g2_decap_8 FILLER_3_2659 ();
 sg13g2_decap_4 FILLER_3_2666 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_36 ();
 sg13g2_fill_1 FILLER_4_38 ();
 sg13g2_fill_1 FILLER_4_65 ();
 sg13g2_fill_2 FILLER_4_126 ();
 sg13g2_fill_1 FILLER_4_128 ();
 sg13g2_decap_4 FILLER_4_139 ();
 sg13g2_decap_8 FILLER_4_169 ();
 sg13g2_decap_4 FILLER_4_176 ();
 sg13g2_fill_1 FILLER_4_180 ();
 sg13g2_fill_1 FILLER_4_211 ();
 sg13g2_decap_4 FILLER_4_222 ();
 sg13g2_decap_8 FILLER_4_262 ();
 sg13g2_fill_2 FILLER_4_269 ();
 sg13g2_fill_1 FILLER_4_271 ();
 sg13g2_fill_2 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_365 ();
 sg13g2_fill_2 FILLER_4_372 ();
 sg13g2_fill_1 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_4 FILLER_4_409 ();
 sg13g2_fill_2 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_fill_2 FILLER_4_448 ();
 sg13g2_fill_1 FILLER_4_450 ();
 sg13g2_fill_2 FILLER_4_456 ();
 sg13g2_decap_4 FILLER_4_463 ();
 sg13g2_fill_2 FILLER_4_467 ();
 sg13g2_fill_1 FILLER_4_488 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_4 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_583 ();
 sg13g2_decap_8 FILLER_4_590 ();
 sg13g2_fill_2 FILLER_4_597 ();
 sg13g2_fill_1 FILLER_4_599 ();
 sg13g2_fill_1 FILLER_4_610 ();
 sg13g2_decap_4 FILLER_4_637 ();
 sg13g2_fill_1 FILLER_4_645 ();
 sg13g2_decap_8 FILLER_4_650 ();
 sg13g2_decap_8 FILLER_4_657 ();
 sg13g2_decap_8 FILLER_4_664 ();
 sg13g2_fill_2 FILLER_4_671 ();
 sg13g2_decap_4 FILLER_4_707 ();
 sg13g2_fill_1 FILLER_4_711 ();
 sg13g2_decap_4 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_772 ();
 sg13g2_fill_2 FILLER_4_784 ();
 sg13g2_decap_4 FILLER_4_791 ();
 sg13g2_fill_2 FILLER_4_799 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_fill_2 FILLER_4_812 ();
 sg13g2_fill_1 FILLER_4_814 ();
 sg13g2_fill_1 FILLER_4_849 ();
 sg13g2_decap_4 FILLER_4_880 ();
 sg13g2_fill_2 FILLER_4_884 ();
 sg13g2_fill_2 FILLER_4_890 ();
 sg13g2_decap_8 FILLER_4_896 ();
 sg13g2_decap_8 FILLER_4_903 ();
 sg13g2_decap_8 FILLER_4_910 ();
 sg13g2_decap_4 FILLER_4_923 ();
 sg13g2_fill_1 FILLER_4_927 ();
 sg13g2_decap_8 FILLER_4_993 ();
 sg13g2_decap_8 FILLER_4_1000 ();
 sg13g2_decap_8 FILLER_4_1007 ();
 sg13g2_decap_4 FILLER_4_1014 ();
 sg13g2_decap_4 FILLER_4_1044 ();
 sg13g2_fill_1 FILLER_4_1048 ();
 sg13g2_fill_1 FILLER_4_1053 ();
 sg13g2_fill_1 FILLER_4_1059 ();
 sg13g2_decap_8 FILLER_4_1077 ();
 sg13g2_decap_8 FILLER_4_1084 ();
 sg13g2_fill_1 FILLER_4_1096 ();
 sg13g2_decap_4 FILLER_4_1118 ();
 sg13g2_fill_1 FILLER_4_1122 ();
 sg13g2_fill_2 FILLER_4_1128 ();
 sg13g2_decap_8 FILLER_4_1134 ();
 sg13g2_decap_8 FILLER_4_1141 ();
 sg13g2_decap_8 FILLER_4_1148 ();
 sg13g2_fill_2 FILLER_4_1155 ();
 sg13g2_fill_1 FILLER_4_1157 ();
 sg13g2_decap_8 FILLER_4_1194 ();
 sg13g2_decap_8 FILLER_4_1201 ();
 sg13g2_decap_8 FILLER_4_1212 ();
 sg13g2_fill_2 FILLER_4_1219 ();
 sg13g2_decap_8 FILLER_4_1251 ();
 sg13g2_decap_8 FILLER_4_1258 ();
 sg13g2_decap_8 FILLER_4_1265 ();
 sg13g2_decap_8 FILLER_4_1272 ();
 sg13g2_decap_8 FILLER_4_1279 ();
 sg13g2_fill_1 FILLER_4_1286 ();
 sg13g2_decap_8 FILLER_4_1292 ();
 sg13g2_decap_4 FILLER_4_1299 ();
 sg13g2_decap_4 FILLER_4_1307 ();
 sg13g2_fill_1 FILLER_4_1311 ();
 sg13g2_decap_4 FILLER_4_1315 ();
 sg13g2_fill_2 FILLER_4_1319 ();
 sg13g2_decap_8 FILLER_4_1356 ();
 sg13g2_decap_8 FILLER_4_1363 ();
 sg13g2_decap_4 FILLER_4_1370 ();
 sg13g2_fill_1 FILLER_4_1374 ();
 sg13g2_fill_1 FILLER_4_1385 ();
 sg13g2_fill_1 FILLER_4_1391 ();
 sg13g2_decap_8 FILLER_4_1396 ();
 sg13g2_decap_4 FILLER_4_1403 ();
 sg13g2_fill_2 FILLER_4_1407 ();
 sg13g2_fill_2 FILLER_4_1418 ();
 sg13g2_fill_2 FILLER_4_1430 ();
 sg13g2_fill_2 FILLER_4_1458 ();
 sg13g2_fill_2 FILLER_4_1486 ();
 sg13g2_decap_4 FILLER_4_1514 ();
 sg13g2_decap_4 FILLER_4_1528 ();
 sg13g2_fill_1 FILLER_4_1532 ();
 sg13g2_fill_2 FILLER_4_1537 ();
 sg13g2_fill_1 FILLER_4_1539 ();
 sg13g2_decap_8 FILLER_4_1574 ();
 sg13g2_decap_8 FILLER_4_1581 ();
 sg13g2_fill_1 FILLER_4_1588 ();
 sg13g2_decap_8 FILLER_4_1629 ();
 sg13g2_decap_8 FILLER_4_1636 ();
 sg13g2_decap_8 FILLER_4_1643 ();
 sg13g2_fill_2 FILLER_4_1702 ();
 sg13g2_fill_1 FILLER_4_1708 ();
 sg13g2_fill_2 FILLER_4_1721 ();
 sg13g2_decap_4 FILLER_4_1764 ();
 sg13g2_fill_1 FILLER_4_1768 ();
 sg13g2_fill_2 FILLER_4_1774 ();
 sg13g2_fill_2 FILLER_4_1780 ();
 sg13g2_decap_8 FILLER_4_1800 ();
 sg13g2_decap_8 FILLER_4_1807 ();
 sg13g2_decap_4 FILLER_4_1814 ();
 sg13g2_fill_2 FILLER_4_1818 ();
 sg13g2_fill_1 FILLER_4_1829 ();
 sg13g2_decap_8 FILLER_4_1847 ();
 sg13g2_fill_2 FILLER_4_1854 ();
 sg13g2_decap_8 FILLER_4_1887 ();
 sg13g2_decap_4 FILLER_4_1894 ();
 sg13g2_fill_1 FILLER_4_1898 ();
 sg13g2_fill_1 FILLER_4_1907 ();
 sg13g2_fill_1 FILLER_4_1952 ();
 sg13g2_fill_1 FILLER_4_1966 ();
 sg13g2_decap_4 FILLER_4_1998 ();
 sg13g2_fill_1 FILLER_4_2002 ();
 sg13g2_fill_1 FILLER_4_2027 ();
 sg13g2_fill_1 FILLER_4_2055 ();
 sg13g2_decap_4 FILLER_4_2068 ();
 sg13g2_fill_1 FILLER_4_2072 ();
 sg13g2_fill_2 FILLER_4_2086 ();
 sg13g2_decap_8 FILLER_4_2128 ();
 sg13g2_decap_8 FILLER_4_2135 ();
 sg13g2_decap_8 FILLER_4_2151 ();
 sg13g2_decap_4 FILLER_4_2158 ();
 sg13g2_fill_1 FILLER_4_2194 ();
 sg13g2_decap_4 FILLER_4_2200 ();
 sg13g2_fill_1 FILLER_4_2208 ();
 sg13g2_fill_1 FILLER_4_2215 ();
 sg13g2_fill_1 FILLER_4_2220 ();
 sg13g2_fill_1 FILLER_4_2226 ();
 sg13g2_fill_2 FILLER_4_2230 ();
 sg13g2_fill_1 FILLER_4_2249 ();
 sg13g2_fill_1 FILLER_4_2257 ();
 sg13g2_fill_2 FILLER_4_2262 ();
 sg13g2_fill_2 FILLER_4_2270 ();
 sg13g2_fill_1 FILLER_4_2272 ();
 sg13g2_fill_2 FILLER_4_2276 ();
 sg13g2_fill_1 FILLER_4_2294 ();
 sg13g2_fill_2 FILLER_4_2305 ();
 sg13g2_decap_8 FILLER_4_2316 ();
 sg13g2_decap_8 FILLER_4_2323 ();
 sg13g2_fill_1 FILLER_4_2330 ();
 sg13g2_fill_1 FILLER_4_2375 ();
 sg13g2_fill_2 FILLER_4_2395 ();
 sg13g2_fill_1 FILLER_4_2397 ();
 sg13g2_fill_2 FILLER_4_2424 ();
 sg13g2_fill_1 FILLER_4_2426 ();
 sg13g2_decap_4 FILLER_4_2431 ();
 sg13g2_fill_1 FILLER_4_2461 ();
 sg13g2_fill_1 FILLER_4_2512 ();
 sg13g2_decap_4 FILLER_4_2517 ();
 sg13g2_fill_1 FILLER_4_2535 ();
 sg13g2_decap_8 FILLER_4_2571 ();
 sg13g2_decap_8 FILLER_4_2578 ();
 sg13g2_decap_4 FILLER_4_2585 ();
 sg13g2_decap_8 FILLER_4_2615 ();
 sg13g2_decap_8 FILLER_4_2622 ();
 sg13g2_decap_8 FILLER_4_2629 ();
 sg13g2_decap_8 FILLER_4_2636 ();
 sg13g2_decap_8 FILLER_4_2643 ();
 sg13g2_decap_8 FILLER_4_2650 ();
 sg13g2_decap_8 FILLER_4_2657 ();
 sg13g2_decap_4 FILLER_4_2664 ();
 sg13g2_fill_2 FILLER_4_2668 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_7 ();
 sg13g2_fill_2 FILLER_5_58 ();
 sg13g2_fill_2 FILLER_5_64 ();
 sg13g2_fill_1 FILLER_5_88 ();
 sg13g2_fill_2 FILLER_5_92 ();
 sg13g2_fill_1 FILLER_5_94 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_126 ();
 sg13g2_decap_4 FILLER_5_148 ();
 sg13g2_fill_2 FILLER_5_152 ();
 sg13g2_decap_8 FILLER_5_157 ();
 sg13g2_decap_8 FILLER_5_164 ();
 sg13g2_decap_8 FILLER_5_171 ();
 sg13g2_decap_8 FILLER_5_178 ();
 sg13g2_decap_8 FILLER_5_185 ();
 sg13g2_decap_8 FILLER_5_202 ();
 sg13g2_fill_1 FILLER_5_209 ();
 sg13g2_decap_8 FILLER_5_220 ();
 sg13g2_fill_1 FILLER_5_227 ();
 sg13g2_fill_1 FILLER_5_257 ();
 sg13g2_fill_2 FILLER_5_263 ();
 sg13g2_fill_1 FILLER_5_265 ();
 sg13g2_fill_1 FILLER_5_286 ();
 sg13g2_decap_8 FILLER_5_338 ();
 sg13g2_decap_8 FILLER_5_345 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_359 ();
 sg13g2_decap_8 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_4 FILLER_5_380 ();
 sg13g2_fill_2 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_fill_2 FILLER_5_401 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_4 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_431 ();
 sg13g2_decap_8 FILLER_5_437 ();
 sg13g2_decap_8 FILLER_5_444 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_4 FILLER_5_497 ();
 sg13g2_fill_1 FILLER_5_540 ();
 sg13g2_decap_8 FILLER_5_545 ();
 sg13g2_decap_8 FILLER_5_552 ();
 sg13g2_decap_8 FILLER_5_559 ();
 sg13g2_decap_8 FILLER_5_566 ();
 sg13g2_decap_8 FILLER_5_573 ();
 sg13g2_fill_2 FILLER_5_580 ();
 sg13g2_fill_1 FILLER_5_582 ();
 sg13g2_fill_2 FILLER_5_601 ();
 sg13g2_fill_1 FILLER_5_603 ();
 sg13g2_decap_8 FILLER_5_617 ();
 sg13g2_decap_8 FILLER_5_624 ();
 sg13g2_decap_8 FILLER_5_631 ();
 sg13g2_fill_2 FILLER_5_638 ();
 sg13g2_fill_1 FILLER_5_640 ();
 sg13g2_fill_2 FILLER_5_672 ();
 sg13g2_fill_1 FILLER_5_716 ();
 sg13g2_fill_2 FILLER_5_740 ();
 sg13g2_fill_1 FILLER_5_742 ();
 sg13g2_fill_2 FILLER_5_747 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_4 FILLER_5_819 ();
 sg13g2_fill_1 FILLER_5_823 ();
 sg13g2_fill_2 FILLER_5_851 ();
 sg13g2_fill_2 FILLER_5_863 ();
 sg13g2_fill_1 FILLER_5_869 ();
 sg13g2_decap_8 FILLER_5_876 ();
 sg13g2_decap_8 FILLER_5_883 ();
 sg13g2_decap_8 FILLER_5_890 ();
 sg13g2_decap_4 FILLER_5_909 ();
 sg13g2_fill_1 FILLER_5_913 ();
 sg13g2_fill_2 FILLER_5_940 ();
 sg13g2_fill_1 FILLER_5_942 ();
 sg13g2_decap_8 FILLER_5_987 ();
 sg13g2_decap_8 FILLER_5_994 ();
 sg13g2_fill_2 FILLER_5_1001 ();
 sg13g2_decap_8 FILLER_5_1008 ();
 sg13g2_decap_8 FILLER_5_1015 ();
 sg13g2_fill_2 FILLER_5_1061 ();
 sg13g2_fill_1 FILLER_5_1063 ();
 sg13g2_fill_1 FILLER_5_1079 ();
 sg13g2_decap_4 FILLER_5_1084 ();
 sg13g2_decap_8 FILLER_5_1092 ();
 sg13g2_decap_8 FILLER_5_1099 ();
 sg13g2_decap_4 FILLER_5_1106 ();
 sg13g2_fill_1 FILLER_5_1110 ();
 sg13g2_decap_8 FILLER_5_1117 ();
 sg13g2_decap_8 FILLER_5_1124 ();
 sg13g2_decap_4 FILLER_5_1131 ();
 sg13g2_fill_2 FILLER_5_1135 ();
 sg13g2_decap_4 FILLER_5_1147 ();
 sg13g2_fill_1 FILLER_5_1151 ();
 sg13g2_decap_8 FILLER_5_1178 ();
 sg13g2_decap_4 FILLER_5_1185 ();
 sg13g2_fill_1 FILLER_5_1189 ();
 sg13g2_decap_4 FILLER_5_1204 ();
 sg13g2_fill_2 FILLER_5_1208 ();
 sg13g2_decap_8 FILLER_5_1214 ();
 sg13g2_decap_4 FILLER_5_1221 ();
 sg13g2_fill_2 FILLER_5_1225 ();
 sg13g2_decap_8 FILLER_5_1239 ();
 sg13g2_decap_8 FILLER_5_1246 ();
 sg13g2_decap_4 FILLER_5_1263 ();
 sg13g2_fill_2 FILLER_5_1267 ();
 sg13g2_decap_8 FILLER_5_1274 ();
 sg13g2_decap_8 FILLER_5_1281 ();
 sg13g2_decap_4 FILLER_5_1288 ();
 sg13g2_fill_2 FILLER_5_1292 ();
 sg13g2_decap_4 FILLER_5_1297 ();
 sg13g2_fill_1 FILLER_5_1306 ();
 sg13g2_fill_1 FILLER_5_1311 ();
 sg13g2_fill_2 FILLER_5_1344 ();
 sg13g2_fill_1 FILLER_5_1346 ();
 sg13g2_decap_8 FILLER_5_1356 ();
 sg13g2_fill_2 FILLER_5_1363 ();
 sg13g2_decap_8 FILLER_5_1456 ();
 sg13g2_fill_1 FILLER_5_1463 ();
 sg13g2_decap_8 FILLER_5_1472 ();
 sg13g2_decap_8 FILLER_5_1479 ();
 sg13g2_fill_2 FILLER_5_1486 ();
 sg13g2_decap_4 FILLER_5_1496 ();
 sg13g2_decap_8 FILLER_5_1508 ();
 sg13g2_decap_4 FILLER_5_1515 ();
 sg13g2_fill_1 FILLER_5_1529 ();
 sg13g2_fill_2 FILLER_5_1546 ();
 sg13g2_fill_1 FILLER_5_1548 ();
 sg13g2_fill_1 FILLER_5_1561 ();
 sg13g2_decap_4 FILLER_5_1592 ();
 sg13g2_decap_8 FILLER_5_1604 ();
 sg13g2_decap_4 FILLER_5_1611 ();
 sg13g2_fill_2 FILLER_5_1615 ();
 sg13g2_fill_1 FILLER_5_1630 ();
 sg13g2_decap_8 FILLER_5_1637 ();
 sg13g2_decap_8 FILLER_5_1644 ();
 sg13g2_fill_2 FILLER_5_1651 ();
 sg13g2_fill_1 FILLER_5_1653 ();
 sg13g2_decap_4 FILLER_5_1688 ();
 sg13g2_fill_1 FILLER_5_1731 ();
 sg13g2_fill_2 FILLER_5_1745 ();
 sg13g2_fill_2 FILLER_5_1752 ();
 sg13g2_fill_1 FILLER_5_1754 ();
 sg13g2_fill_1 FILLER_5_1797 ();
 sg13g2_decap_8 FILLER_5_1801 ();
 sg13g2_fill_2 FILLER_5_1808 ();
 sg13g2_decap_8 FILLER_5_1818 ();
 sg13g2_decap_4 FILLER_5_1825 ();
 sg13g2_fill_2 FILLER_5_1829 ();
 sg13g2_decap_8 FILLER_5_1862 ();
 sg13g2_fill_2 FILLER_5_1869 ();
 sg13g2_fill_1 FILLER_5_1871 ();
 sg13g2_fill_2 FILLER_5_1912 ();
 sg13g2_fill_1 FILLER_5_1947 ();
 sg13g2_decap_8 FILLER_5_1953 ();
 sg13g2_decap_8 FILLER_5_1960 ();
 sg13g2_decap_4 FILLER_5_1972 ();
 sg13g2_decap_8 FILLER_5_1980 ();
 sg13g2_decap_4 FILLER_5_1993 ();
 sg13g2_fill_1 FILLER_5_1997 ();
 sg13g2_fill_2 FILLER_5_2010 ();
 sg13g2_fill_1 FILLER_5_2032 ();
 sg13g2_decap_8 FILLER_5_2076 ();
 sg13g2_decap_4 FILLER_5_2083 ();
 sg13g2_fill_2 FILLER_5_2087 ();
 sg13g2_decap_8 FILLER_5_2120 ();
 sg13g2_decap_8 FILLER_5_2127 ();
 sg13g2_decap_8 FILLER_5_2134 ();
 sg13g2_decap_8 FILLER_5_2141 ();
 sg13g2_decap_8 FILLER_5_2148 ();
 sg13g2_decap_8 FILLER_5_2155 ();
 sg13g2_decap_4 FILLER_5_2162 ();
 sg13g2_fill_2 FILLER_5_2166 ();
 sg13g2_fill_2 FILLER_5_2194 ();
 sg13g2_fill_1 FILLER_5_2196 ();
 sg13g2_fill_2 FILLER_5_2203 ();
 sg13g2_fill_1 FILLER_5_2205 ();
 sg13g2_fill_2 FILLER_5_2263 ();
 sg13g2_decap_4 FILLER_5_2269 ();
 sg13g2_fill_1 FILLER_5_2273 ();
 sg13g2_fill_1 FILLER_5_2312 ();
 sg13g2_decap_8 FILLER_5_2343 ();
 sg13g2_fill_2 FILLER_5_2350 ();
 sg13g2_fill_2 FILLER_5_2357 ();
 sg13g2_fill_2 FILLER_5_2368 ();
 sg13g2_decap_8 FILLER_5_2411 ();
 sg13g2_fill_2 FILLER_5_2418 ();
 sg13g2_fill_2 FILLER_5_2430 ();
 sg13g2_decap_8 FILLER_5_2437 ();
 sg13g2_decap_8 FILLER_5_2444 ();
 sg13g2_fill_2 FILLER_5_2451 ();
 sg13g2_fill_1 FILLER_5_2453 ();
 sg13g2_decap_8 FILLER_5_2459 ();
 sg13g2_decap_8 FILLER_5_2466 ();
 sg13g2_decap_4 FILLER_5_2473 ();
 sg13g2_fill_2 FILLER_5_2477 ();
 sg13g2_decap_4 FILLER_5_2490 ();
 sg13g2_fill_1 FILLER_5_2494 ();
 sg13g2_decap_8 FILLER_5_2499 ();
 sg13g2_fill_2 FILLER_5_2506 ();
 sg13g2_fill_1 FILLER_5_2508 ();
 sg13g2_decap_8 FILLER_5_2514 ();
 sg13g2_decap_8 FILLER_5_2521 ();
 sg13g2_decap_8 FILLER_5_2528 ();
 sg13g2_decap_8 FILLER_5_2535 ();
 sg13g2_decap_8 FILLER_5_2542 ();
 sg13g2_decap_8 FILLER_5_2549 ();
 sg13g2_decap_4 FILLER_5_2556 ();
 sg13g2_fill_1 FILLER_5_2560 ();
 sg13g2_decap_8 FILLER_5_2565 ();
 sg13g2_decap_8 FILLER_5_2607 ();
 sg13g2_decap_8 FILLER_5_2614 ();
 sg13g2_decap_8 FILLER_5_2621 ();
 sg13g2_decap_8 FILLER_5_2628 ();
 sg13g2_decap_8 FILLER_5_2635 ();
 sg13g2_decap_8 FILLER_5_2642 ();
 sg13g2_decap_8 FILLER_5_2649 ();
 sg13g2_decap_8 FILLER_5_2656 ();
 sg13g2_decap_8 FILLER_5_2663 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_18 ();
 sg13g2_decap_8 FILLER_6_53 ();
 sg13g2_fill_1 FILLER_6_60 ();
 sg13g2_decap_8 FILLER_6_94 ();
 sg13g2_decap_8 FILLER_6_101 ();
 sg13g2_decap_8 FILLER_6_108 ();
 sg13g2_decap_8 FILLER_6_115 ();
 sg13g2_fill_2 FILLER_6_122 ();
 sg13g2_decap_8 FILLER_6_148 ();
 sg13g2_decap_8 FILLER_6_155 ();
 sg13g2_decap_8 FILLER_6_162 ();
 sg13g2_decap_8 FILLER_6_169 ();
 sg13g2_decap_8 FILLER_6_176 ();
 sg13g2_decap_8 FILLER_6_183 ();
 sg13g2_decap_8 FILLER_6_190 ();
 sg13g2_decap_8 FILLER_6_197 ();
 sg13g2_decap_8 FILLER_6_204 ();
 sg13g2_decap_8 FILLER_6_211 ();
 sg13g2_decap_8 FILLER_6_218 ();
 sg13g2_decap_8 FILLER_6_225 ();
 sg13g2_fill_2 FILLER_6_232 ();
 sg13g2_decap_4 FILLER_6_244 ();
 sg13g2_decap_8 FILLER_6_263 ();
 sg13g2_decap_8 FILLER_6_270 ();
 sg13g2_decap_8 FILLER_6_281 ();
 sg13g2_decap_4 FILLER_6_288 ();
 sg13g2_fill_2 FILLER_6_292 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_fill_2 FILLER_6_333 ();
 sg13g2_fill_1 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_fill_1 FILLER_6_379 ();
 sg13g2_fill_2 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_6_423 ();
 sg13g2_fill_1 FILLER_6_430 ();
 sg13g2_decap_4 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_498 ();
 sg13g2_fill_2 FILLER_6_505 ();
 sg13g2_fill_1 FILLER_6_507 ();
 sg13g2_decap_8 FILLER_6_552 ();
 sg13g2_decap_4 FILLER_6_559 ();
 sg13g2_fill_2 FILLER_6_563 ();
 sg13g2_fill_1 FILLER_6_575 ();
 sg13g2_fill_2 FILLER_6_606 ();
 sg13g2_decap_4 FILLER_6_634 ();
 sg13g2_fill_1 FILLER_6_678 ();
 sg13g2_fill_1 FILLER_6_683 ();
 sg13g2_fill_2 FILLER_6_705 ();
 sg13g2_decap_8 FILLER_6_713 ();
 sg13g2_decap_8 FILLER_6_720 ();
 sg13g2_decap_8 FILLER_6_727 ();
 sg13g2_decap_8 FILLER_6_734 ();
 sg13g2_decap_8 FILLER_6_741 ();
 sg13g2_decap_4 FILLER_6_748 ();
 sg13g2_fill_1 FILLER_6_752 ();
 sg13g2_decap_4 FILLER_6_765 ();
 sg13g2_fill_1 FILLER_6_769 ();
 sg13g2_fill_2 FILLER_6_806 ();
 sg13g2_fill_1 FILLER_6_808 ();
 sg13g2_decap_8 FILLER_6_815 ();
 sg13g2_decap_8 FILLER_6_822 ();
 sg13g2_fill_2 FILLER_6_849 ();
 sg13g2_fill_2 FILLER_6_856 ();
 sg13g2_fill_1 FILLER_6_858 ();
 sg13g2_fill_2 FILLER_6_880 ();
 sg13g2_fill_1 FILLER_6_882 ();
 sg13g2_fill_1 FILLER_6_945 ();
 sg13g2_fill_2 FILLER_6_965 ();
 sg13g2_decap_8 FILLER_6_1001 ();
 sg13g2_decap_4 FILLER_6_1008 ();
 sg13g2_fill_2 FILLER_6_1012 ();
 sg13g2_decap_8 FILLER_6_1019 ();
 sg13g2_decap_8 FILLER_6_1026 ();
 sg13g2_fill_2 FILLER_6_1033 ();
 sg13g2_fill_1 FILLER_6_1035 ();
 sg13g2_decap_4 FILLER_6_1042 ();
 sg13g2_fill_2 FILLER_6_1061 ();
 sg13g2_fill_1 FILLER_6_1063 ();
 sg13g2_decap_8 FILLER_6_1090 ();
 sg13g2_fill_2 FILLER_6_1097 ();
 sg13g2_fill_1 FILLER_6_1099 ();
 sg13g2_decap_8 FILLER_6_1157 ();
 sg13g2_decap_4 FILLER_6_1164 ();
 sg13g2_fill_1 FILLER_6_1168 ();
 sg13g2_decap_4 FILLER_6_1179 ();
 sg13g2_fill_2 FILLER_6_1183 ();
 sg13g2_fill_2 FILLER_6_1191 ();
 sg13g2_decap_8 FILLER_6_1225 ();
 sg13g2_fill_2 FILLER_6_1232 ();
 sg13g2_fill_1 FILLER_6_1234 ();
 sg13g2_fill_1 FILLER_6_1240 ();
 sg13g2_fill_2 FILLER_6_1272 ();
 sg13g2_decap_8 FILLER_6_1279 ();
 sg13g2_fill_2 FILLER_6_1286 ();
 sg13g2_fill_1 FILLER_6_1324 ();
 sg13g2_fill_1 FILLER_6_1337 ();
 sg13g2_decap_8 FILLER_6_1342 ();
 sg13g2_decap_8 FILLER_6_1375 ();
 sg13g2_decap_8 FILLER_6_1382 ();
 sg13g2_fill_2 FILLER_6_1389 ();
 sg13g2_fill_1 FILLER_6_1391 ();
 sg13g2_decap_4 FILLER_6_1400 ();
 sg13g2_decap_4 FILLER_6_1417 ();
 sg13g2_fill_1 FILLER_6_1425 ();
 sg13g2_decap_8 FILLER_6_1430 ();
 sg13g2_fill_2 FILLER_6_1437 ();
 sg13g2_fill_1 FILLER_6_1439 ();
 sg13g2_decap_8 FILLER_6_1466 ();
 sg13g2_decap_8 FILLER_6_1473 ();
 sg13g2_fill_2 FILLER_6_1480 ();
 sg13g2_fill_1 FILLER_6_1482 ();
 sg13g2_fill_1 FILLER_6_1489 ();
 sg13g2_fill_2 FILLER_6_1552 ();
 sg13g2_decap_4 FILLER_6_1571 ();
 sg13g2_fill_2 FILLER_6_1575 ();
 sg13g2_decap_4 FILLER_6_1590 ();
 sg13g2_fill_2 FILLER_6_1594 ();
 sg13g2_decap_8 FILLER_6_1618 ();
 sg13g2_decap_4 FILLER_6_1629 ();
 sg13g2_fill_1 FILLER_6_1633 ();
 sg13g2_decap_4 FILLER_6_1660 ();
 sg13g2_fill_2 FILLER_6_1664 ();
 sg13g2_decap_8 FILLER_6_1679 ();
 sg13g2_fill_2 FILLER_6_1686 ();
 sg13g2_fill_1 FILLER_6_1688 ();
 sg13g2_fill_2 FILLER_6_1721 ();
 sg13g2_fill_2 FILLER_6_1787 ();
 sg13g2_fill_1 FILLER_6_1789 ();
 sg13g2_fill_2 FILLER_6_1796 ();
 sg13g2_decap_8 FILLER_6_1804 ();
 sg13g2_decap_4 FILLER_6_1811 ();
 sg13g2_fill_2 FILLER_6_1841 ();
 sg13g2_fill_2 FILLER_6_1861 ();
 sg13g2_fill_2 FILLER_6_1869 ();
 sg13g2_fill_1 FILLER_6_1871 ();
 sg13g2_decap_4 FILLER_6_1884 ();
 sg13g2_fill_2 FILLER_6_1888 ();
 sg13g2_fill_2 FILLER_6_1958 ();
 sg13g2_fill_1 FILLER_6_1960 ();
 sg13g2_decap_8 FILLER_6_1966 ();
 sg13g2_decap_8 FILLER_6_1973 ();
 sg13g2_fill_1 FILLER_6_1980 ();
 sg13g2_fill_2 FILLER_6_1985 ();
 sg13g2_fill_1 FILLER_6_1987 ();
 sg13g2_fill_1 FILLER_6_2000 ();
 sg13g2_fill_1 FILLER_6_2010 ();
 sg13g2_decap_8 FILLER_6_2017 ();
 sg13g2_fill_2 FILLER_6_2024 ();
 sg13g2_fill_1 FILLER_6_2026 ();
 sg13g2_fill_2 FILLER_6_2066 ();
 sg13g2_decap_8 FILLER_6_2077 ();
 sg13g2_fill_1 FILLER_6_2084 ();
 sg13g2_fill_2 FILLER_6_2116 ();
 sg13g2_fill_1 FILLER_6_2118 ();
 sg13g2_fill_2 FILLER_6_2155 ();
 sg13g2_decap_8 FILLER_6_2162 ();
 sg13g2_fill_2 FILLER_6_2169 ();
 sg13g2_fill_2 FILLER_6_2176 ();
 sg13g2_decap_8 FILLER_6_2188 ();
 sg13g2_fill_1 FILLER_6_2195 ();
 sg13g2_fill_2 FILLER_6_2222 ();
 sg13g2_fill_1 FILLER_6_2250 ();
 sg13g2_decap_8 FILLER_6_2270 ();
 sg13g2_decap_4 FILLER_6_2277 ();
 sg13g2_decap_8 FILLER_6_2284 ();
 sg13g2_fill_2 FILLER_6_2291 ();
 sg13g2_decap_8 FILLER_6_2328 ();
 sg13g2_decap_8 FILLER_6_2335 ();
 sg13g2_decap_8 FILLER_6_2342 ();
 sg13g2_fill_1 FILLER_6_2349 ();
 sg13g2_fill_2 FILLER_6_2379 ();
 sg13g2_fill_1 FILLER_6_2381 ();
 sg13g2_fill_2 FILLER_6_2387 ();
 sg13g2_fill_2 FILLER_6_2395 ();
 sg13g2_decap_4 FILLER_6_2405 ();
 sg13g2_decap_8 FILLER_6_2439 ();
 sg13g2_decap_4 FILLER_6_2446 ();
 sg13g2_fill_1 FILLER_6_2450 ();
 sg13g2_decap_8 FILLER_6_2457 ();
 sg13g2_decap_8 FILLER_6_2464 ();
 sg13g2_fill_1 FILLER_6_2471 ();
 sg13g2_fill_1 FILLER_6_2504 ();
 sg13g2_decap_8 FILLER_6_2531 ();
 sg13g2_decap_4 FILLER_6_2538 ();
 sg13g2_fill_1 FILLER_6_2542 ();
 sg13g2_decap_4 FILLER_6_2569 ();
 sg13g2_fill_1 FILLER_6_2573 ();
 sg13g2_fill_2 FILLER_6_2579 ();
 sg13g2_fill_1 FILLER_6_2581 ();
 sg13g2_decap_8 FILLER_6_2591 ();
 sg13g2_decap_8 FILLER_6_2598 ();
 sg13g2_decap_8 FILLER_6_2605 ();
 sg13g2_decap_8 FILLER_6_2612 ();
 sg13g2_decap_8 FILLER_6_2619 ();
 sg13g2_decap_8 FILLER_6_2626 ();
 sg13g2_decap_8 FILLER_6_2633 ();
 sg13g2_decap_8 FILLER_6_2640 ();
 sg13g2_decap_8 FILLER_6_2647 ();
 sg13g2_decap_8 FILLER_6_2654 ();
 sg13g2_decap_8 FILLER_6_2661 ();
 sg13g2_fill_2 FILLER_6_2668 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_4 FILLER_7_28 ();
 sg13g2_fill_1 FILLER_7_32 ();
 sg13g2_fill_1 FILLER_7_43 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_4 FILLER_7_63 ();
 sg13g2_fill_1 FILLER_7_67 ();
 sg13g2_decap_8 FILLER_7_81 ();
 sg13g2_fill_2 FILLER_7_88 ();
 sg13g2_decap_8 FILLER_7_120 ();
 sg13g2_fill_1 FILLER_7_127 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_fill_2 FILLER_7_168 ();
 sg13g2_fill_1 FILLER_7_199 ();
 sg13g2_fill_1 FILLER_7_205 ();
 sg13g2_fill_1 FILLER_7_216 ();
 sg13g2_decap_8 FILLER_7_221 ();
 sg13g2_decap_4 FILLER_7_228 ();
 sg13g2_fill_1 FILLER_7_232 ();
 sg13g2_decap_4 FILLER_7_269 ();
 sg13g2_decap_8 FILLER_7_305 ();
 sg13g2_decap_8 FILLER_7_312 ();
 sg13g2_fill_1 FILLER_7_355 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_fill_2 FILLER_7_402 ();
 sg13g2_fill_1 FILLER_7_407 ();
 sg13g2_fill_1 FILLER_7_474 ();
 sg13g2_decap_8 FILLER_7_479 ();
 sg13g2_decap_4 FILLER_7_486 ();
 sg13g2_fill_2 FILLER_7_490 ();
 sg13g2_fill_2 FILLER_7_498 ();
 sg13g2_decap_8 FILLER_7_505 ();
 sg13g2_decap_8 FILLER_7_512 ();
 sg13g2_fill_1 FILLER_7_539 ();
 sg13g2_fill_1 FILLER_7_545 ();
 sg13g2_fill_2 FILLER_7_572 ();
 sg13g2_decap_4 FILLER_7_600 ();
 sg13g2_decap_4 FILLER_7_640 ();
 sg13g2_fill_2 FILLER_7_644 ();
 sg13g2_fill_1 FILLER_7_655 ();
 sg13g2_decap_8 FILLER_7_661 ();
 sg13g2_decap_8 FILLER_7_668 ();
 sg13g2_decap_8 FILLER_7_675 ();
 sg13g2_fill_1 FILLER_7_682 ();
 sg13g2_fill_1 FILLER_7_733 ();
 sg13g2_fill_2 FILLER_7_747 ();
 sg13g2_decap_8 FILLER_7_762 ();
 sg13g2_decap_8 FILLER_7_769 ();
 sg13g2_decap_4 FILLER_7_776 ();
 sg13g2_fill_2 FILLER_7_822 ();
 sg13g2_decap_8 FILLER_7_828 ();
 sg13g2_fill_2 FILLER_7_877 ();
 sg13g2_decap_4 FILLER_7_919 ();
 sg13g2_fill_2 FILLER_7_923 ();
 sg13g2_decap_8 FILLER_7_929 ();
 sg13g2_decap_8 FILLER_7_940 ();
 sg13g2_decap_8 FILLER_7_947 ();
 sg13g2_fill_2 FILLER_7_954 ();
 sg13g2_fill_1 FILLER_7_956 ();
 sg13g2_fill_2 FILLER_7_991 ();
 sg13g2_fill_1 FILLER_7_993 ();
 sg13g2_fill_1 FILLER_7_1052 ();
 sg13g2_fill_1 FILLER_7_1067 ();
 sg13g2_decap_8 FILLER_7_1094 ();
 sg13g2_fill_2 FILLER_7_1101 ();
 sg13g2_fill_1 FILLER_7_1114 ();
 sg13g2_fill_1 FILLER_7_1120 ();
 sg13g2_fill_2 FILLER_7_1126 ();
 sg13g2_fill_2 FILLER_7_1133 ();
 sg13g2_fill_1 FILLER_7_1156 ();
 sg13g2_decap_8 FILLER_7_1199 ();
 sg13g2_fill_1 FILLER_7_1206 ();
 sg13g2_fill_1 FILLER_7_1233 ();
 sg13g2_fill_2 FILLER_7_1323 ();
 sg13g2_fill_1 FILLER_7_1331 ();
 sg13g2_fill_1 FILLER_7_1342 ();
 sg13g2_fill_1 FILLER_7_1369 ();
 sg13g2_fill_1 FILLER_7_1374 ();
 sg13g2_fill_1 FILLER_7_1432 ();
 sg13g2_decap_8 FILLER_7_1438 ();
 sg13g2_decap_4 FILLER_7_1445 ();
 sg13g2_decap_8 FILLER_7_1481 ();
 sg13g2_fill_2 FILLER_7_1514 ();
 sg13g2_fill_2 FILLER_7_1522 ();
 sg13g2_fill_2 FILLER_7_1530 ();
 sg13g2_fill_2 FILLER_7_1570 ();
 sg13g2_fill_1 FILLER_7_1572 ();
 sg13g2_fill_2 FILLER_7_1664 ();
 sg13g2_fill_1 FILLER_7_1666 ();
 sg13g2_fill_1 FILLER_7_1703 ();
 sg13g2_fill_1 FILLER_7_1847 ();
 sg13g2_decap_8 FILLER_7_1856 ();
 sg13g2_decap_4 FILLER_7_1863 ();
 sg13g2_fill_2 FILLER_7_1867 ();
 sg13g2_decap_4 FILLER_7_1891 ();
 sg13g2_decap_8 FILLER_7_1921 ();
 sg13g2_fill_2 FILLER_7_1928 ();
 sg13g2_fill_1 FILLER_7_1930 ();
 sg13g2_fill_1 FILLER_7_1936 ();
 sg13g2_fill_1 FILLER_7_1942 ();
 sg13g2_fill_1 FILLER_7_1953 ();
 sg13g2_decap_4 FILLER_7_1959 ();
 sg13g2_fill_1 FILLER_7_1963 ();
 sg13g2_fill_2 FILLER_7_1990 ();
 sg13g2_fill_2 FILLER_7_2029 ();
 sg13g2_fill_1 FILLER_7_2070 ();
 sg13g2_fill_2 FILLER_7_2097 ();
 sg13g2_fill_1 FILLER_7_2099 ();
 sg13g2_decap_8 FILLER_7_2104 ();
 sg13g2_decap_8 FILLER_7_2111 ();
 sg13g2_decap_4 FILLER_7_2122 ();
 sg13g2_decap_4 FILLER_7_2132 ();
 sg13g2_fill_2 FILLER_7_2136 ();
 sg13g2_fill_1 FILLER_7_2164 ();
 sg13g2_decap_4 FILLER_7_2174 ();
 sg13g2_fill_2 FILLER_7_2184 ();
 sg13g2_decap_4 FILLER_7_2192 ();
 sg13g2_decap_8 FILLER_7_2200 ();
 sg13g2_decap_8 FILLER_7_2207 ();
 sg13g2_decap_4 FILLER_7_2214 ();
 sg13g2_fill_1 FILLER_7_2218 ();
 sg13g2_fill_1 FILLER_7_2269 ();
 sg13g2_decap_8 FILLER_7_2276 ();
 sg13g2_decap_8 FILLER_7_2283 ();
 sg13g2_decap_4 FILLER_7_2290 ();
 sg13g2_fill_1 FILLER_7_2303 ();
 sg13g2_fill_1 FILLER_7_2339 ();
 sg13g2_fill_1 FILLER_7_2346 ();
 sg13g2_fill_1 FILLER_7_2359 ();
 sg13g2_decap_8 FILLER_7_2379 ();
 sg13g2_fill_2 FILLER_7_2386 ();
 sg13g2_decap_4 FILLER_7_2394 ();
 sg13g2_fill_1 FILLER_7_2398 ();
 sg13g2_decap_8 FILLER_7_2408 ();
 sg13g2_decap_4 FILLER_7_2415 ();
 sg13g2_fill_1 FILLER_7_2419 ();
 sg13g2_fill_1 FILLER_7_2454 ();
 sg13g2_fill_2 FILLER_7_2486 ();
 sg13g2_decap_4 FILLER_7_2498 ();
 sg13g2_fill_1 FILLER_7_2507 ();
 sg13g2_fill_1 FILLER_7_2512 ();
 sg13g2_fill_1 FILLER_7_2518 ();
 sg13g2_fill_1 FILLER_7_2545 ();
 sg13g2_decap_8 FILLER_7_2620 ();
 sg13g2_decap_8 FILLER_7_2627 ();
 sg13g2_decap_8 FILLER_7_2634 ();
 sg13g2_decap_8 FILLER_7_2641 ();
 sg13g2_decap_8 FILLER_7_2648 ();
 sg13g2_decap_8 FILLER_7_2655 ();
 sg13g2_decap_8 FILLER_7_2662 ();
 sg13g2_fill_1 FILLER_7_2669 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_2 ();
 sg13g2_fill_1 FILLER_8_29 ();
 sg13g2_decap_8 FILLER_8_81 ();
 sg13g2_fill_1 FILLER_8_88 ();
 sg13g2_fill_1 FILLER_8_101 ();
 sg13g2_decap_8 FILLER_8_115 ();
 sg13g2_decap_4 FILLER_8_122 ();
 sg13g2_fill_1 FILLER_8_126 ();
 sg13g2_decap_4 FILLER_8_131 ();
 sg13g2_decap_8 FILLER_8_165 ();
 sg13g2_decap_8 FILLER_8_172 ();
 sg13g2_fill_2 FILLER_8_179 ();
 sg13g2_fill_1 FILLER_8_181 ();
 sg13g2_decap_4 FILLER_8_192 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_fill_1 FILLER_8_303 ();
 sg13g2_fill_1 FILLER_8_309 ();
 sg13g2_fill_2 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_369 ();
 sg13g2_decap_4 FILLER_8_411 ();
 sg13g2_decap_4 FILLER_8_419 ();
 sg13g2_decap_4 FILLER_8_453 ();
 sg13g2_fill_2 FILLER_8_462 ();
 sg13g2_fill_1 FILLER_8_464 ();
 sg13g2_fill_1 FILLER_8_470 ();
 sg13g2_fill_1 FILLER_8_475 ();
 sg13g2_fill_1 FILLER_8_490 ();
 sg13g2_fill_2 FILLER_8_497 ();
 sg13g2_fill_1 FILLER_8_499 ();
 sg13g2_decap_8 FILLER_8_505 ();
 sg13g2_fill_1 FILLER_8_512 ();
 sg13g2_fill_2 FILLER_8_526 ();
 sg13g2_fill_1 FILLER_8_528 ();
 sg13g2_decap_8 FILLER_8_618 ();
 sg13g2_decap_8 FILLER_8_625 ();
 sg13g2_decap_8 FILLER_8_632 ();
 sg13g2_decap_8 FILLER_8_639 ();
 sg13g2_fill_1 FILLER_8_646 ();
 sg13g2_decap_8 FILLER_8_652 ();
 sg13g2_decap_4 FILLER_8_659 ();
 sg13g2_fill_2 FILLER_8_663 ();
 sg13g2_decap_4 FILLER_8_669 ();
 sg13g2_decap_4 FILLER_8_686 ();
 sg13g2_fill_2 FILLER_8_690 ();
 sg13g2_decap_4 FILLER_8_698 ();
 sg13g2_decap_8 FILLER_8_754 ();
 sg13g2_decap_4 FILLER_8_761 ();
 sg13g2_fill_1 FILLER_8_765 ();
 sg13g2_fill_2 FILLER_8_826 ();
 sg13g2_fill_2 FILLER_8_832 ();
 sg13g2_fill_1 FILLER_8_866 ();
 sg13g2_fill_2 FILLER_8_878 ();
 sg13g2_fill_1 FILLER_8_880 ();
 sg13g2_fill_2 FILLER_8_885 ();
 sg13g2_decap_8 FILLER_8_923 ();
 sg13g2_decap_4 FILLER_8_930 ();
 sg13g2_fill_1 FILLER_8_934 ();
 sg13g2_decap_8 FILLER_8_943 ();
 sg13g2_fill_2 FILLER_8_954 ();
 sg13g2_fill_1 FILLER_8_956 ();
 sg13g2_decap_4 FILLER_8_963 ();
 sg13g2_decap_8 FILLER_8_985 ();
 sg13g2_fill_1 FILLER_8_992 ();
 sg13g2_fill_1 FILLER_8_1001 ();
 sg13g2_fill_2 FILLER_8_1007 ();
 sg13g2_fill_1 FILLER_8_1025 ();
 sg13g2_fill_1 FILLER_8_1034 ();
 sg13g2_fill_1 FILLER_8_1051 ();
 sg13g2_fill_1 FILLER_8_1080 ();
 sg13g2_fill_2 FILLER_8_1096 ();
 sg13g2_fill_1 FILLER_8_1106 ();
 sg13g2_decap_8 FILLER_8_1130 ();
 sg13g2_decap_8 FILLER_8_1137 ();
 sg13g2_fill_2 FILLER_8_1144 ();
 sg13g2_fill_2 FILLER_8_1158 ();
 sg13g2_fill_1 FILLER_8_1160 ();
 sg13g2_fill_2 FILLER_8_1179 ();
 sg13g2_fill_1 FILLER_8_1181 ();
 sg13g2_decap_8 FILLER_8_1188 ();
 sg13g2_decap_8 FILLER_8_1195 ();
 sg13g2_fill_2 FILLER_8_1202 ();
 sg13g2_fill_1 FILLER_8_1204 ();
 sg13g2_fill_2 FILLER_8_1209 ();
 sg13g2_decap_8 FILLER_8_1221 ();
 sg13g2_fill_2 FILLER_8_1228 ();
 sg13g2_fill_1 FILLER_8_1230 ();
 sg13g2_fill_2 FILLER_8_1273 ();
 sg13g2_fill_1 FILLER_8_1275 ();
 sg13g2_fill_1 FILLER_8_1309 ();
 sg13g2_decap_4 FILLER_8_1337 ();
 sg13g2_fill_1 FILLER_8_1341 ();
 sg13g2_decap_4 FILLER_8_1347 ();
 sg13g2_fill_1 FILLER_8_1351 ();
 sg13g2_decap_4 FILLER_8_1356 ();
 sg13g2_fill_2 FILLER_8_1366 ();
 sg13g2_fill_1 FILLER_8_1368 ();
 sg13g2_decap_4 FILLER_8_1392 ();
 sg13g2_fill_2 FILLER_8_1396 ();
 sg13g2_decap_8 FILLER_8_1413 ();
 sg13g2_decap_8 FILLER_8_1420 ();
 sg13g2_decap_8 FILLER_8_1437 ();
 sg13g2_fill_1 FILLER_8_1444 ();
 sg13g2_fill_2 FILLER_8_1454 ();
 sg13g2_fill_1 FILLER_8_1456 ();
 sg13g2_fill_2 FILLER_8_1460 ();
 sg13g2_fill_1 FILLER_8_1462 ();
 sg13g2_decap_8 FILLER_8_1469 ();
 sg13g2_decap_8 FILLER_8_1476 ();
 sg13g2_fill_2 FILLER_8_1483 ();
 sg13g2_decap_4 FILLER_8_1489 ();
 sg13g2_fill_1 FILLER_8_1493 ();
 sg13g2_decap_8 FILLER_8_1498 ();
 sg13g2_decap_4 FILLER_8_1505 ();
 sg13g2_fill_1 FILLER_8_1543 ();
 sg13g2_decap_8 FILLER_8_1560 ();
 sg13g2_decap_8 FILLER_8_1567 ();
 sg13g2_fill_1 FILLER_8_1594 ();
 sg13g2_fill_2 FILLER_8_1608 ();
 sg13g2_decap_8 FILLER_8_1619 ();
 sg13g2_fill_2 FILLER_8_1631 ();
 sg13g2_fill_2 FILLER_8_1638 ();
 sg13g2_fill_1 FILLER_8_1675 ();
 sg13g2_decap_4 FILLER_8_1691 ();
 sg13g2_fill_1 FILLER_8_1695 ();
 sg13g2_fill_1 FILLER_8_1714 ();
 sg13g2_fill_2 FILLER_8_1721 ();
 sg13g2_fill_2 FILLER_8_1732 ();
 sg13g2_fill_2 FILLER_8_1748 ();
 sg13g2_fill_2 FILLER_8_1767 ();
 sg13g2_fill_1 FILLER_8_1769 ();
 sg13g2_decap_4 FILLER_8_1785 ();
 sg13g2_fill_2 FILLER_8_1794 ();
 sg13g2_fill_1 FILLER_8_1802 ();
 sg13g2_decap_8 FILLER_8_1816 ();
 sg13g2_fill_2 FILLER_8_1823 ();
 sg13g2_fill_1 FILLER_8_1825 ();
 sg13g2_decap_8 FILLER_8_1836 ();
 sg13g2_decap_8 FILLER_8_1843 ();
 sg13g2_decap_8 FILLER_8_1850 ();
 sg13g2_decap_4 FILLER_8_1857 ();
 sg13g2_fill_2 FILLER_8_1861 ();
 sg13g2_decap_4 FILLER_8_1889 ();
 sg13g2_fill_1 FILLER_8_1893 ();
 sg13g2_decap_8 FILLER_8_1899 ();
 sg13g2_decap_8 FILLER_8_1906 ();
 sg13g2_fill_2 FILLER_8_1913 ();
 sg13g2_fill_1 FILLER_8_1915 ();
 sg13g2_fill_1 FILLER_8_2024 ();
 sg13g2_decap_4 FILLER_8_2030 ();
 sg13g2_fill_2 FILLER_8_2034 ();
 sg13g2_fill_2 FILLER_8_2045 ();
 sg13g2_fill_2 FILLER_8_2056 ();
 sg13g2_fill_1 FILLER_8_2084 ();
 sg13g2_decap_8 FILLER_8_2097 ();
 sg13g2_decap_8 FILLER_8_2104 ();
 sg13g2_decap_8 FILLER_8_2148 ();
 sg13g2_decap_4 FILLER_8_2155 ();
 sg13g2_decap_8 FILLER_8_2168 ();
 sg13g2_fill_2 FILLER_8_2175 ();
 sg13g2_fill_1 FILLER_8_2177 ();
 sg13g2_fill_2 FILLER_8_2238 ();
 sg13g2_decap_8 FILLER_8_2281 ();
 sg13g2_fill_2 FILLER_8_2288 ();
 sg13g2_fill_1 FILLER_8_2290 ();
 sg13g2_decap_4 FILLER_8_2340 ();
 sg13g2_fill_1 FILLER_8_2344 ();
 sg13g2_decap_4 FILLER_8_2351 ();
 sg13g2_fill_2 FILLER_8_2355 ();
 sg13g2_fill_2 FILLER_8_2387 ();
 sg13g2_fill_1 FILLER_8_2389 ();
 sg13g2_fill_2 FILLER_8_2398 ();
 sg13g2_fill_1 FILLER_8_2400 ();
 sg13g2_decap_4 FILLER_8_2416 ();
 sg13g2_fill_2 FILLER_8_2438 ();
 sg13g2_fill_1 FILLER_8_2440 ();
 sg13g2_fill_2 FILLER_8_2457 ();
 sg13g2_fill_2 FILLER_8_2497 ();
 sg13g2_decap_8 FILLER_8_2505 ();
 sg13g2_fill_2 FILLER_8_2512 ();
 sg13g2_decap_8 FILLER_8_2518 ();
 sg13g2_decap_8 FILLER_8_2525 ();
 sg13g2_decap_8 FILLER_8_2532 ();
 sg13g2_fill_2 FILLER_8_2539 ();
 sg13g2_fill_1 FILLER_8_2555 ();
 sg13g2_fill_2 FILLER_8_2560 ();
 sg13g2_fill_1 FILLER_8_2562 ();
 sg13g2_fill_2 FILLER_8_2593 ();
 sg13g2_decap_8 FILLER_8_2621 ();
 sg13g2_decap_8 FILLER_8_2628 ();
 sg13g2_decap_8 FILLER_8_2635 ();
 sg13g2_decap_8 FILLER_8_2642 ();
 sg13g2_decap_8 FILLER_8_2649 ();
 sg13g2_decap_8 FILLER_8_2656 ();
 sg13g2_decap_8 FILLER_8_2663 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_2 ();
 sg13g2_decap_4 FILLER_9_46 ();
 sg13g2_fill_2 FILLER_9_50 ();
 sg13g2_decap_4 FILLER_9_57 ();
 sg13g2_decap_8 FILLER_9_69 ();
 sg13g2_decap_8 FILLER_9_76 ();
 sg13g2_decap_8 FILLER_9_83 ();
 sg13g2_decap_8 FILLER_9_132 ();
 sg13g2_fill_2 FILLER_9_139 ();
 sg13g2_fill_1 FILLER_9_141 ();
 sg13g2_decap_8 FILLER_9_150 ();
 sg13g2_decap_8 FILLER_9_157 ();
 sg13g2_decap_8 FILLER_9_164 ();
 sg13g2_fill_2 FILLER_9_171 ();
 sg13g2_fill_2 FILLER_9_199 ();
 sg13g2_decap_4 FILLER_9_276 ();
 sg13g2_fill_1 FILLER_9_285 ();
 sg13g2_fill_1 FILLER_9_312 ();
 sg13g2_fill_1 FILLER_9_331 ();
 sg13g2_fill_1 FILLER_9_358 ();
 sg13g2_fill_2 FILLER_9_390 ();
 sg13g2_fill_2 FILLER_9_402 ();
 sg13g2_fill_1 FILLER_9_404 ();
 sg13g2_decap_4 FILLER_9_416 ();
 sg13g2_fill_2 FILLER_9_432 ();
 sg13g2_fill_1 FILLER_9_434 ();
 sg13g2_fill_1 FILLER_9_454 ();
 sg13g2_fill_1 FILLER_9_459 ();
 sg13g2_decap_8 FILLER_9_496 ();
 sg13g2_decap_8 FILLER_9_503 ();
 sg13g2_decap_8 FILLER_9_510 ();
 sg13g2_decap_8 FILLER_9_517 ();
 sg13g2_decap_8 FILLER_9_524 ();
 sg13g2_fill_2 FILLER_9_531 ();
 sg13g2_fill_1 FILLER_9_533 ();
 sg13g2_fill_1 FILLER_9_544 ();
 sg13g2_decap_8 FILLER_9_549 ();
 sg13g2_decap_8 FILLER_9_556 ();
 sg13g2_decap_8 FILLER_9_563 ();
 sg13g2_decap_4 FILLER_9_570 ();
 sg13g2_fill_2 FILLER_9_574 ();
 sg13g2_fill_1 FILLER_9_596 ();
 sg13g2_fill_2 FILLER_9_607 ();
 sg13g2_fill_1 FILLER_9_609 ();
 sg13g2_fill_2 FILLER_9_618 ();
 sg13g2_decap_8 FILLER_9_625 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_fill_1 FILLER_9_668 ();
 sg13g2_decap_8 FILLER_9_674 ();
 sg13g2_decap_8 FILLER_9_681 ();
 sg13g2_fill_1 FILLER_9_688 ();
 sg13g2_fill_1 FILLER_9_715 ();
 sg13g2_decap_8 FILLER_9_755 ();
 sg13g2_fill_2 FILLER_9_762 ();
 sg13g2_fill_1 FILLER_9_764 ();
 sg13g2_decap_8 FILLER_9_813 ();
 sg13g2_fill_1 FILLER_9_847 ();
 sg13g2_decap_4 FILLER_9_861 ();
 sg13g2_fill_1 FILLER_9_865 ();
 sg13g2_decap_8 FILLER_9_878 ();
 sg13g2_decap_4 FILLER_9_885 ();
 sg13g2_fill_1 FILLER_9_889 ();
 sg13g2_decap_8 FILLER_9_907 ();
 sg13g2_decap_4 FILLER_9_927 ();
 sg13g2_fill_1 FILLER_9_931 ();
 sg13g2_decap_4 FILLER_9_936 ();
 sg13g2_fill_1 FILLER_9_940 ();
 sg13g2_decap_4 FILLER_9_946 ();
 sg13g2_fill_2 FILLER_9_950 ();
 sg13g2_fill_2 FILLER_9_957 ();
 sg13g2_fill_1 FILLER_9_959 ();
 sg13g2_decap_8 FILLER_9_1017 ();
 sg13g2_decap_4 FILLER_9_1024 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_fill_2 FILLER_9_1042 ();
 sg13g2_fill_2 FILLER_9_1097 ();
 sg13g2_fill_1 FILLER_9_1115 ();
 sg13g2_fill_2 FILLER_9_1119 ();
 sg13g2_decap_8 FILLER_9_1129 ();
 sg13g2_fill_1 FILLER_9_1136 ();
 sg13g2_fill_2 FILLER_9_1163 ();
 sg13g2_decap_4 FILLER_9_1170 ();
 sg13g2_fill_2 FILLER_9_1174 ();
 sg13g2_decap_8 FILLER_9_1184 ();
 sg13g2_decap_8 FILLER_9_1191 ();
 sg13g2_decap_8 FILLER_9_1198 ();
 sg13g2_decap_4 FILLER_9_1205 ();
 sg13g2_fill_2 FILLER_9_1217 ();
 sg13g2_fill_2 FILLER_9_1236 ();
 sg13g2_fill_2 FILLER_9_1256 ();
 sg13g2_fill_1 FILLER_9_1275 ();
 sg13g2_fill_2 FILLER_9_1292 ();
 sg13g2_fill_1 FILLER_9_1299 ();
 sg13g2_fill_1 FILLER_9_1311 ();
 sg13g2_decap_4 FILLER_9_1368 ();
 sg13g2_fill_1 FILLER_9_1377 ();
 sg13g2_decap_4 FILLER_9_1394 ();
 sg13g2_fill_2 FILLER_9_1398 ();
 sg13g2_decap_4 FILLER_9_1412 ();
 sg13g2_fill_1 FILLER_9_1416 ();
 sg13g2_fill_2 FILLER_9_1426 ();
 sg13g2_fill_2 FILLER_9_1454 ();
 sg13g2_fill_1 FILLER_9_1456 ();
 sg13g2_fill_2 FILLER_9_1463 ();
 sg13g2_decap_4 FILLER_9_1492 ();
 sg13g2_decap_4 FILLER_9_1501 ();
 sg13g2_decap_8 FILLER_9_1517 ();
 sg13g2_fill_2 FILLER_9_1524 ();
 sg13g2_decap_8 FILLER_9_1561 ();
 sg13g2_fill_2 FILLER_9_1583 ();
 sg13g2_fill_1 FILLER_9_1585 ();
 sg13g2_decap_8 FILLER_9_1601 ();
 sg13g2_fill_2 FILLER_9_1608 ();
 sg13g2_fill_1 FILLER_9_1610 ();
 sg13g2_fill_1 FILLER_9_1637 ();
 sg13g2_decap_8 FILLER_9_1642 ();
 sg13g2_decap_4 FILLER_9_1649 ();
 sg13g2_decap_8 FILLER_9_1681 ();
 sg13g2_fill_2 FILLER_9_1688 ();
 sg13g2_fill_1 FILLER_9_1690 ();
 sg13g2_decap_8 FILLER_9_1696 ();
 sg13g2_decap_8 FILLER_9_1703 ();
 sg13g2_decap_8 FILLER_9_1710 ();
 sg13g2_decap_4 FILLER_9_1717 ();
 sg13g2_fill_2 FILLER_9_1721 ();
 sg13g2_decap_8 FILLER_9_1726 ();
 sg13g2_fill_2 FILLER_9_1733 ();
 sg13g2_decap_8 FILLER_9_1748 ();
 sg13g2_decap_8 FILLER_9_1755 ();
 sg13g2_fill_2 FILLER_9_1762 ();
 sg13g2_fill_1 FILLER_9_1764 ();
 sg13g2_decap_8 FILLER_9_1782 ();
 sg13g2_decap_8 FILLER_9_1789 ();
 sg13g2_decap_8 FILLER_9_1796 ();
 sg13g2_decap_4 FILLER_9_1803 ();
 sg13g2_fill_1 FILLER_9_1807 ();
 sg13g2_fill_2 FILLER_9_1813 ();
 sg13g2_fill_1 FILLER_9_1827 ();
 sg13g2_decap_4 FILLER_9_1881 ();
 sg13g2_decap_8 FILLER_9_1889 ();
 sg13g2_decap_4 FILLER_9_1928 ();
 sg13g2_fill_1 FILLER_9_1932 ();
 sg13g2_fill_1 FILLER_9_1939 ();
 sg13g2_decap_8 FILLER_9_1950 ();
 sg13g2_fill_2 FILLER_9_1957 ();
 sg13g2_fill_1 FILLER_9_1959 ();
 sg13g2_fill_2 FILLER_9_1990 ();
 sg13g2_fill_2 FILLER_9_2003 ();
 sg13g2_fill_2 FILLER_9_2037 ();
 sg13g2_fill_1 FILLER_9_2054 ();
 sg13g2_fill_2 FILLER_9_2061 ();
 sg13g2_decap_4 FILLER_9_2135 ();
 sg13g2_decap_8 FILLER_9_2143 ();
 sg13g2_fill_1 FILLER_9_2150 ();
 sg13g2_fill_2 FILLER_9_2165 ();
 sg13g2_fill_1 FILLER_9_2167 ();
 sg13g2_fill_2 FILLER_9_2173 ();
 sg13g2_fill_2 FILLER_9_2187 ();
 sg13g2_fill_1 FILLER_9_2204 ();
 sg13g2_decap_8 FILLER_9_2214 ();
 sg13g2_decap_8 FILLER_9_2239 ();
 sg13g2_fill_1 FILLER_9_2249 ();
 sg13g2_fill_2 FILLER_9_2255 ();
 sg13g2_fill_1 FILLER_9_2312 ();
 sg13g2_decap_8 FILLER_9_2317 ();
 sg13g2_decap_8 FILLER_9_2324 ();
 sg13g2_fill_1 FILLER_9_2331 ();
 sg13g2_decap_8 FILLER_9_2337 ();
 sg13g2_decap_8 FILLER_9_2344 ();
 sg13g2_decap_8 FILLER_9_2351 ();
 sg13g2_fill_2 FILLER_9_2420 ();
 sg13g2_fill_1 FILLER_9_2422 ();
 sg13g2_fill_2 FILLER_9_2489 ();
 sg13g2_decap_4 FILLER_9_2517 ();
 sg13g2_decap_4 FILLER_9_2555 ();
 sg13g2_fill_2 FILLER_9_2559 ();
 sg13g2_decap_8 FILLER_9_2605 ();
 sg13g2_decap_8 FILLER_9_2612 ();
 sg13g2_decap_8 FILLER_9_2619 ();
 sg13g2_decap_8 FILLER_9_2626 ();
 sg13g2_decap_8 FILLER_9_2633 ();
 sg13g2_decap_8 FILLER_9_2640 ();
 sg13g2_decap_8 FILLER_9_2647 ();
 sg13g2_decap_8 FILLER_9_2654 ();
 sg13g2_decap_8 FILLER_9_2661 ();
 sg13g2_fill_2 FILLER_9_2668 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_11 ();
 sg13g2_decap_4 FILLER_10_24 ();
 sg13g2_fill_2 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_43 ();
 sg13g2_decap_4 FILLER_10_50 ();
 sg13g2_decap_8 FILLER_10_67 ();
 sg13g2_decap_8 FILLER_10_74 ();
 sg13g2_decap_8 FILLER_10_81 ();
 sg13g2_fill_2 FILLER_10_88 ();
 sg13g2_fill_2 FILLER_10_100 ();
 sg13g2_fill_1 FILLER_10_102 ();
 sg13g2_decap_8 FILLER_10_108 ();
 sg13g2_decap_8 FILLER_10_115 ();
 sg13g2_decap_8 FILLER_10_122 ();
 sg13g2_decap_8 FILLER_10_129 ();
 sg13g2_decap_8 FILLER_10_136 ();
 sg13g2_decap_8 FILLER_10_143 ();
 sg13g2_decap_8 FILLER_10_150 ();
 sg13g2_decap_8 FILLER_10_157 ();
 sg13g2_decap_8 FILLER_10_164 ();
 sg13g2_decap_8 FILLER_10_171 ();
 sg13g2_decap_8 FILLER_10_178 ();
 sg13g2_fill_1 FILLER_10_185 ();
 sg13g2_fill_1 FILLER_10_196 ();
 sg13g2_fill_2 FILLER_10_201 ();
 sg13g2_fill_1 FILLER_10_203 ();
 sg13g2_fill_1 FILLER_10_214 ();
 sg13g2_fill_2 FILLER_10_241 ();
 sg13g2_fill_1 FILLER_10_243 ();
 sg13g2_decap_4 FILLER_10_264 ();
 sg13g2_fill_2 FILLER_10_303 ();
 sg13g2_decap_8 FILLER_10_309 ();
 sg13g2_fill_2 FILLER_10_316 ();
 sg13g2_decap_8 FILLER_10_328 ();
 sg13g2_decap_8 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_fill_1 FILLER_10_370 ();
 sg13g2_fill_2 FILLER_10_385 ();
 sg13g2_fill_1 FILLER_10_397 ();
 sg13g2_decap_4 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_10_411 ();
 sg13g2_decap_8 FILLER_10_418 ();
 sg13g2_decap_8 FILLER_10_425 ();
 sg13g2_decap_8 FILLER_10_432 ();
 sg13g2_decap_4 FILLER_10_439 ();
 sg13g2_fill_1 FILLER_10_443 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_fill_2 FILLER_10_455 ();
 sg13g2_fill_1 FILLER_10_461 ();
 sg13g2_decap_8 FILLER_10_466 ();
 sg13g2_fill_2 FILLER_10_473 ();
 sg13g2_fill_1 FILLER_10_479 ();
 sg13g2_fill_1 FILLER_10_485 ();
 sg13g2_fill_2 FILLER_10_491 ();
 sg13g2_fill_2 FILLER_10_499 ();
 sg13g2_fill_1 FILLER_10_501 ();
 sg13g2_fill_1 FILLER_10_510 ();
 sg13g2_decap_8 FILLER_10_520 ();
 sg13g2_decap_4 FILLER_10_537 ();
 sg13g2_decap_8 FILLER_10_549 ();
 sg13g2_decap_8 FILLER_10_556 ();
 sg13g2_decap_8 FILLER_10_563 ();
 sg13g2_decap_8 FILLER_10_570 ();
 sg13g2_decap_8 FILLER_10_577 ();
 sg13g2_decap_8 FILLER_10_584 ();
 sg13g2_decap_8 FILLER_10_612 ();
 sg13g2_decap_8 FILLER_10_619 ();
 sg13g2_decap_8 FILLER_10_626 ();
 sg13g2_fill_1 FILLER_10_633 ();
 sg13g2_decap_8 FILLER_10_648 ();
 sg13g2_decap_8 FILLER_10_655 ();
 sg13g2_fill_2 FILLER_10_667 ();
 sg13g2_decap_8 FILLER_10_673 ();
 sg13g2_decap_8 FILLER_10_680 ();
 sg13g2_decap_8 FILLER_10_687 ();
 sg13g2_decap_8 FILLER_10_694 ();
 sg13g2_fill_2 FILLER_10_701 ();
 sg13g2_fill_1 FILLER_10_703 ();
 sg13g2_decap_8 FILLER_10_757 ();
 sg13g2_decap_8 FILLER_10_764 ();
 sg13g2_fill_1 FILLER_10_771 ();
 sg13g2_decap_8 FILLER_10_780 ();
 sg13g2_decap_8 FILLER_10_787 ();
 sg13g2_decap_8 FILLER_10_794 ();
 sg13g2_decap_8 FILLER_10_801 ();
 sg13g2_decap_8 FILLER_10_808 ();
 sg13g2_decap_8 FILLER_10_815 ();
 sg13g2_decap_8 FILLER_10_822 ();
 sg13g2_decap_8 FILLER_10_829 ();
 sg13g2_fill_2 FILLER_10_836 ();
 sg13g2_fill_1 FILLER_10_838 ();
 sg13g2_fill_1 FILLER_10_874 ();
 sg13g2_decap_4 FILLER_10_918 ();
 sg13g2_fill_2 FILLER_10_922 ();
 sg13g2_decap_8 FILLER_10_932 ();
 sg13g2_decap_8 FILLER_10_939 ();
 sg13g2_decap_4 FILLER_10_946 ();
 sg13g2_decap_8 FILLER_10_953 ();
 sg13g2_decap_4 FILLER_10_973 ();
 sg13g2_fill_2 FILLER_10_977 ();
 sg13g2_fill_2 FILLER_10_988 ();
 sg13g2_decap_4 FILLER_10_1031 ();
 sg13g2_fill_1 FILLER_10_1035 ();
 sg13g2_fill_2 FILLER_10_1048 ();
 sg13g2_fill_1 FILLER_10_1062 ();
 sg13g2_fill_1 FILLER_10_1098 ();
 sg13g2_decap_8 FILLER_10_1123 ();
 sg13g2_decap_8 FILLER_10_1130 ();
 sg13g2_fill_2 FILLER_10_1140 ();
 sg13g2_fill_1 FILLER_10_1142 ();
 sg13g2_decap_8 FILLER_10_1190 ();
 sg13g2_fill_2 FILLER_10_1197 ();
 sg13g2_decap_8 FILLER_10_1208 ();
 sg13g2_decap_4 FILLER_10_1215 ();
 sg13g2_fill_1 FILLER_10_1219 ();
 sg13g2_fill_2 FILLER_10_1230 ();
 sg13g2_fill_2 FILLER_10_1236 ();
 sg13g2_fill_1 FILLER_10_1238 ();
 sg13g2_fill_1 FILLER_10_1265 ();
 sg13g2_fill_2 FILLER_10_1292 ();
 sg13g2_fill_2 FILLER_10_1298 ();
 sg13g2_decap_4 FILLER_10_1322 ();
 sg13g2_decap_4 FILLER_10_1332 ();
 sg13g2_fill_1 FILLER_10_1336 ();
 sg13g2_decap_8 FILLER_10_1342 ();
 sg13g2_decap_8 FILLER_10_1349 ();
 sg13g2_decap_8 FILLER_10_1356 ();
 sg13g2_fill_1 FILLER_10_1363 ();
 sg13g2_decap_8 FILLER_10_1396 ();
 sg13g2_decap_8 FILLER_10_1403 ();
 sg13g2_fill_1 FILLER_10_1410 ();
 sg13g2_decap_8 FILLER_10_1419 ();
 sg13g2_decap_8 FILLER_10_1426 ();
 sg13g2_decap_8 FILLER_10_1437 ();
 sg13g2_decap_8 FILLER_10_1444 ();
 sg13g2_decap_8 FILLER_10_1451 ();
 sg13g2_decap_8 FILLER_10_1458 ();
 sg13g2_fill_2 FILLER_10_1471 ();
 sg13g2_decap_8 FILLER_10_1491 ();
 sg13g2_decap_8 FILLER_10_1498 ();
 sg13g2_decap_4 FILLER_10_1505 ();
 sg13g2_fill_1 FILLER_10_1509 ();
 sg13g2_decap_8 FILLER_10_1515 ();
 sg13g2_decap_4 FILLER_10_1522 ();
 sg13g2_fill_1 FILLER_10_1526 ();
 sg13g2_decap_8 FILLER_10_1559 ();
 sg13g2_decap_8 FILLER_10_1566 ();
 sg13g2_decap_4 FILLER_10_1573 ();
 sg13g2_decap_8 FILLER_10_1603 ();
 sg13g2_decap_4 FILLER_10_1610 ();
 sg13g2_decap_4 FILLER_10_1648 ();
 sg13g2_fill_1 FILLER_10_1652 ();
 sg13g2_decap_8 FILLER_10_1674 ();
 sg13g2_decap_8 FILLER_10_1681 ();
 sg13g2_decap_4 FILLER_10_1688 ();
 sg13g2_fill_2 FILLER_10_1692 ();
 sg13g2_decap_8 FILLER_10_1704 ();
 sg13g2_decap_8 FILLER_10_1711 ();
 sg13g2_decap_8 FILLER_10_1718 ();
 sg13g2_decap_8 FILLER_10_1725 ();
 sg13g2_fill_2 FILLER_10_1762 ();
 sg13g2_decap_4 FILLER_10_1781 ();
 sg13g2_decap_8 FILLER_10_1795 ();
 sg13g2_decap_8 FILLER_10_1802 ();
 sg13g2_decap_8 FILLER_10_1809 ();
 sg13g2_decap_8 FILLER_10_1816 ();
 sg13g2_fill_2 FILLER_10_1832 ();
 sg13g2_fill_1 FILLER_10_1834 ();
 sg13g2_fill_1 FILLER_10_1840 ();
 sg13g2_decap_8 FILLER_10_1846 ();
 sg13g2_decap_8 FILLER_10_1853 ();
 sg13g2_decap_8 FILLER_10_1860 ();
 sg13g2_decap_8 FILLER_10_1867 ();
 sg13g2_fill_2 FILLER_10_1874 ();
 sg13g2_fill_1 FILLER_10_1876 ();
 sg13g2_fill_2 FILLER_10_1886 ();
 sg13g2_decap_4 FILLER_10_1894 ();
 sg13g2_decap_8 FILLER_10_1912 ();
 sg13g2_decap_8 FILLER_10_1919 ();
 sg13g2_decap_4 FILLER_10_1926 ();
 sg13g2_decap_8 FILLER_10_1939 ();
 sg13g2_decap_4 FILLER_10_1946 ();
 sg13g2_fill_2 FILLER_10_1950 ();
 sg13g2_fill_2 FILLER_10_1958 ();
 sg13g2_decap_8 FILLER_10_2012 ();
 sg13g2_decap_8 FILLER_10_2019 ();
 sg13g2_decap_8 FILLER_10_2026 ();
 sg13g2_fill_1 FILLER_10_2033 ();
 sg13g2_fill_1 FILLER_10_2057 ();
 sg13g2_fill_1 FILLER_10_2066 ();
 sg13g2_decap_4 FILLER_10_2072 ();
 sg13g2_fill_2 FILLER_10_2080 ();
 sg13g2_fill_2 FILLER_10_2095 ();
 sg13g2_fill_1 FILLER_10_2097 ();
 sg13g2_fill_2 FILLER_10_2106 ();
 sg13g2_fill_1 FILLER_10_2108 ();
 sg13g2_fill_2 FILLER_10_2118 ();
 sg13g2_fill_1 FILLER_10_2120 ();
 sg13g2_decap_8 FILLER_10_2134 ();
 sg13g2_decap_4 FILLER_10_2141 ();
 sg13g2_fill_1 FILLER_10_2145 ();
 sg13g2_fill_2 FILLER_10_2182 ();
 sg13g2_fill_1 FILLER_10_2213 ();
 sg13g2_fill_2 FILLER_10_2252 ();
 sg13g2_fill_2 FILLER_10_2262 ();
 sg13g2_fill_1 FILLER_10_2273 ();
 sg13g2_decap_8 FILLER_10_2297 ();
 sg13g2_decap_8 FILLER_10_2304 ();
 sg13g2_decap_8 FILLER_10_2311 ();
 sg13g2_decap_4 FILLER_10_2318 ();
 sg13g2_decap_4 FILLER_10_2326 ();
 sg13g2_decap_8 FILLER_10_2334 ();
 sg13g2_fill_1 FILLER_10_2341 ();
 sg13g2_fill_1 FILLER_10_2360 ();
 sg13g2_fill_2 FILLER_10_2392 ();
 sg13g2_fill_2 FILLER_10_2399 ();
 sg13g2_fill_1 FILLER_10_2401 ();
 sg13g2_decap_8 FILLER_10_2406 ();
 sg13g2_fill_1 FILLER_10_2413 ();
 sg13g2_decap_8 FILLER_10_2422 ();
 sg13g2_fill_2 FILLER_10_2429 ();
 sg13g2_fill_1 FILLER_10_2431 ();
 sg13g2_decap_4 FILLER_10_2438 ();
 sg13g2_fill_2 FILLER_10_2446 ();
 sg13g2_fill_1 FILLER_10_2474 ();
 sg13g2_fill_1 FILLER_10_2489 ();
 sg13g2_decap_8 FILLER_10_2503 ();
 sg13g2_decap_8 FILLER_10_2510 ();
 sg13g2_decap_4 FILLER_10_2522 ();
 sg13g2_decap_8 FILLER_10_2531 ();
 sg13g2_decap_8 FILLER_10_2538 ();
 sg13g2_fill_2 FILLER_10_2545 ();
 sg13g2_fill_1 FILLER_10_2547 ();
 sg13g2_decap_8 FILLER_10_2557 ();
 sg13g2_decap_8 FILLER_10_2564 ();
 sg13g2_fill_2 FILLER_10_2571 ();
 sg13g2_fill_1 FILLER_10_2573 ();
 sg13g2_decap_8 FILLER_10_2583 ();
 sg13g2_decap_8 FILLER_10_2590 ();
 sg13g2_decap_8 FILLER_10_2597 ();
 sg13g2_decap_8 FILLER_10_2604 ();
 sg13g2_decap_8 FILLER_10_2611 ();
 sg13g2_decap_8 FILLER_10_2618 ();
 sg13g2_decap_8 FILLER_10_2625 ();
 sg13g2_decap_8 FILLER_10_2632 ();
 sg13g2_decap_8 FILLER_10_2639 ();
 sg13g2_decap_8 FILLER_10_2646 ();
 sg13g2_decap_8 FILLER_10_2653 ();
 sg13g2_decap_8 FILLER_10_2660 ();
 sg13g2_fill_2 FILLER_10_2667 ();
 sg13g2_fill_1 FILLER_10_2669 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_4 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_72 ();
 sg13g2_decap_4 FILLER_11_100 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_fill_2 FILLER_11_119 ();
 sg13g2_fill_1 FILLER_11_121 ();
 sg13g2_decap_8 FILLER_11_127 ();
 sg13g2_decap_8 FILLER_11_134 ();
 sg13g2_fill_1 FILLER_11_141 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_4 FILLER_11_203 ();
 sg13g2_fill_1 FILLER_11_207 ();
 sg13g2_decap_4 FILLER_11_218 ();
 sg13g2_fill_2 FILLER_11_222 ();
 sg13g2_decap_8 FILLER_11_229 ();
 sg13g2_decap_8 FILLER_11_236 ();
 sg13g2_decap_8 FILLER_11_243 ();
 sg13g2_decap_8 FILLER_11_250 ();
 sg13g2_decap_8 FILLER_11_281 ();
 sg13g2_fill_1 FILLER_11_288 ();
 sg13g2_decap_4 FILLER_11_293 ();
 sg13g2_fill_1 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_365 ();
 sg13g2_decap_4 FILLER_11_372 ();
 sg13g2_fill_1 FILLER_11_376 ();
 sg13g2_decap_4 FILLER_11_384 ();
 sg13g2_fill_2 FILLER_11_388 ();
 sg13g2_decap_4 FILLER_11_396 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_decap_4 FILLER_11_410 ();
 sg13g2_fill_2 FILLER_11_414 ();
 sg13g2_decap_8 FILLER_11_442 ();
 sg13g2_decap_4 FILLER_11_449 ();
 sg13g2_fill_2 FILLER_11_459 ();
 sg13g2_decap_8 FILLER_11_470 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_fill_2 FILLER_11_574 ();
 sg13g2_fill_2 FILLER_11_612 ();
 sg13g2_decap_8 FILLER_11_640 ();
 sg13g2_decap_8 FILLER_11_647 ();
 sg13g2_fill_1 FILLER_11_654 ();
 sg13g2_decap_8 FILLER_11_685 ();
 sg13g2_decap_4 FILLER_11_692 ();
 sg13g2_decap_4 FILLER_11_713 ();
 sg13g2_decap_8 FILLER_11_724 ();
 sg13g2_decap_8 FILLER_11_731 ();
 sg13g2_decap_8 FILLER_11_738 ();
 sg13g2_decap_8 FILLER_11_745 ();
 sg13g2_decap_4 FILLER_11_752 ();
 sg13g2_decap_8 FILLER_11_760 ();
 sg13g2_decap_4 FILLER_11_767 ();
 sg13g2_decap_8 FILLER_11_801 ();
 sg13g2_decap_4 FILLER_11_808 ();
 sg13g2_fill_2 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_818 ();
 sg13g2_decap_4 FILLER_11_838 ();
 sg13g2_decap_8 FILLER_11_846 ();
 sg13g2_fill_2 FILLER_11_853 ();
 sg13g2_fill_2 FILLER_11_863 ();
 sg13g2_fill_1 FILLER_11_865 ();
 sg13g2_decap_8 FILLER_11_872 ();
 sg13g2_fill_1 FILLER_11_879 ();
 sg13g2_decap_8 FILLER_11_884 ();
 sg13g2_decap_4 FILLER_11_891 ();
 sg13g2_fill_1 FILLER_11_895 ();
 sg13g2_decap_4 FILLER_11_900 ();
 sg13g2_decap_8 FILLER_11_908 ();
 sg13g2_decap_8 FILLER_11_915 ();
 sg13g2_decap_4 FILLER_11_922 ();
 sg13g2_fill_1 FILLER_11_926 ();
 sg13g2_fill_1 FILLER_11_931 ();
 sg13g2_decap_8 FILLER_11_966 ();
 sg13g2_decap_8 FILLER_11_973 ();
 sg13g2_decap_8 FILLER_11_980 ();
 sg13g2_decap_8 FILLER_11_987 ();
 sg13g2_fill_1 FILLER_11_994 ();
 sg13g2_fill_1 FILLER_11_1011 ();
 sg13g2_fill_1 FILLER_11_1017 ();
 sg13g2_decap_8 FILLER_11_1053 ();
 sg13g2_fill_1 FILLER_11_1060 ();
 sg13g2_fill_2 FILLER_11_1070 ();
 sg13g2_decap_4 FILLER_11_1091 ();
 sg13g2_fill_1 FILLER_11_1095 ();
 sg13g2_decap_8 FILLER_11_1122 ();
 sg13g2_decap_8 FILLER_11_1129 ();
 sg13g2_fill_1 FILLER_11_1136 ();
 sg13g2_decap_4 FILLER_11_1142 ();
 sg13g2_fill_1 FILLER_11_1146 ();
 sg13g2_fill_2 FILLER_11_1184 ();
 sg13g2_fill_1 FILLER_11_1186 ();
 sg13g2_fill_1 FILLER_11_1247 ();
 sg13g2_fill_2 FILLER_11_1266 ();
 sg13g2_fill_1 FILLER_11_1268 ();
 sg13g2_decap_8 FILLER_11_1278 ();
 sg13g2_fill_1 FILLER_11_1285 ();
 sg13g2_decap_8 FILLER_11_1292 ();
 sg13g2_fill_1 FILLER_11_1299 ();
 sg13g2_fill_2 FILLER_11_1306 ();
 sg13g2_fill_2 FILLER_11_1338 ();
 sg13g2_decap_4 FILLER_11_1372 ();
 sg13g2_fill_2 FILLER_11_1376 ();
 sg13g2_decap_4 FILLER_11_1402 ();
 sg13g2_fill_2 FILLER_11_1406 ();
 sg13g2_fill_2 FILLER_11_1439 ();
 sg13g2_decap_8 FILLER_11_1485 ();
 sg13g2_decap_4 FILLER_11_1492 ();
 sg13g2_fill_1 FILLER_11_1496 ();
 sg13g2_fill_2 FILLER_11_1505 ();
 sg13g2_decap_8 FILLER_11_1520 ();
 sg13g2_decap_8 FILLER_11_1527 ();
 sg13g2_fill_1 FILLER_11_1534 ();
 sg13g2_decap_4 FILLER_11_1556 ();
 sg13g2_fill_2 FILLER_11_1560 ();
 sg13g2_decap_8 FILLER_11_1575 ();
 sg13g2_decap_8 FILLER_11_1582 ();
 sg13g2_fill_2 FILLER_11_1589 ();
 sg13g2_fill_1 FILLER_11_1591 ();
 sg13g2_decap_8 FILLER_11_1601 ();
 sg13g2_decap_8 FILLER_11_1608 ();
 sg13g2_decap_8 FILLER_11_1615 ();
 sg13g2_fill_1 FILLER_11_1622 ();
 sg13g2_decap_8 FILLER_11_1650 ();
 sg13g2_decap_4 FILLER_11_1657 ();
 sg13g2_fill_1 FILLER_11_1692 ();
 sg13g2_fill_2 FILLER_11_1785 ();
 sg13g2_fill_2 FILLER_11_1790 ();
 sg13g2_decap_4 FILLER_11_1797 ();
 sg13g2_fill_1 FILLER_11_1801 ();
 sg13g2_fill_2 FILLER_11_1807 ();
 sg13g2_fill_1 FILLER_11_1809 ();
 sg13g2_decap_4 FILLER_11_1815 ();
 sg13g2_fill_2 FILLER_11_1819 ();
 sg13g2_fill_1 FILLER_11_1854 ();
 sg13g2_decap_4 FILLER_11_1859 ();
 sg13g2_fill_2 FILLER_11_1863 ();
 sg13g2_fill_1 FILLER_11_1886 ();
 sg13g2_fill_2 FILLER_11_1893 ();
 sg13g2_fill_1 FILLER_11_1895 ();
 sg13g2_decap_4 FILLER_11_1944 ();
 sg13g2_fill_1 FILLER_11_1948 ();
 sg13g2_fill_1 FILLER_11_1957 ();
 sg13g2_fill_2 FILLER_11_1964 ();
 sg13g2_decap_8 FILLER_11_1972 ();
 sg13g2_fill_1 FILLER_11_1979 ();
 sg13g2_decap_8 FILLER_11_1985 ();
 sg13g2_fill_1 FILLER_11_1997 ();
 sg13g2_fill_2 FILLER_11_2029 ();
 sg13g2_decap_4 FILLER_11_2074 ();
 sg13g2_fill_2 FILLER_11_2078 ();
 sg13g2_decap_4 FILLER_11_2084 ();
 sg13g2_decap_8 FILLER_11_2098 ();
 sg13g2_decap_8 FILLER_11_2105 ();
 sg13g2_decap_4 FILLER_11_2112 ();
 sg13g2_fill_1 FILLER_11_2116 ();
 sg13g2_decap_8 FILLER_11_2129 ();
 sg13g2_decap_8 FILLER_11_2136 ();
 sg13g2_decap_8 FILLER_11_2143 ();
 sg13g2_decap_4 FILLER_11_2154 ();
 sg13g2_decap_4 FILLER_11_2204 ();
 sg13g2_fill_1 FILLER_11_2208 ();
 sg13g2_decap_4 FILLER_11_2213 ();
 sg13g2_fill_1 FILLER_11_2217 ();
 sg13g2_decap_4 FILLER_11_2227 ();
 sg13g2_decap_8 FILLER_11_2257 ();
 sg13g2_fill_1 FILLER_11_2270 ();
 sg13g2_decap_4 FILLER_11_2303 ();
 sg13g2_fill_1 FILLER_11_2307 ();
 sg13g2_decap_4 FILLER_11_2312 ();
 sg13g2_fill_2 FILLER_11_2316 ();
 sg13g2_fill_2 FILLER_11_2323 ();
 sg13g2_fill_2 FILLER_11_2387 ();
 sg13g2_fill_1 FILLER_11_2389 ();
 sg13g2_decap_4 FILLER_11_2400 ();
 sg13g2_fill_1 FILLER_11_2404 ();
 sg13g2_fill_2 FILLER_11_2409 ();
 sg13g2_fill_1 FILLER_11_2419 ();
 sg13g2_decap_8 FILLER_11_2425 ();
 sg13g2_fill_2 FILLER_11_2438 ();
 sg13g2_fill_1 FILLER_11_2440 ();
 sg13g2_fill_1 FILLER_11_2493 ();
 sg13g2_decap_4 FILLER_11_2510 ();
 sg13g2_decap_8 FILLER_11_2544 ();
 sg13g2_fill_2 FILLER_11_2577 ();
 sg13g2_decap_4 FILLER_11_2610 ();
 sg13g2_decap_8 FILLER_11_2644 ();
 sg13g2_decap_8 FILLER_11_2651 ();
 sg13g2_decap_8 FILLER_11_2658 ();
 sg13g2_decap_4 FILLER_11_2665 ();
 sg13g2_fill_1 FILLER_11_2669 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_9 ();
 sg13g2_decap_4 FILLER_12_39 ();
 sg13g2_fill_1 FILLER_12_43 ();
 sg13g2_fill_1 FILLER_12_86 ();
 sg13g2_decap_8 FILLER_12_136 ();
 sg13g2_decap_8 FILLER_12_143 ();
 sg13g2_decap_8 FILLER_12_186 ();
 sg13g2_decap_8 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_214 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_fill_2 FILLER_12_228 ();
 sg13g2_fill_1 FILLER_12_230 ();
 sg13g2_decap_8 FILLER_12_244 ();
 sg13g2_decap_8 FILLER_12_251 ();
 sg13g2_fill_1 FILLER_12_258 ();
 sg13g2_decap_8 FILLER_12_272 ();
 sg13g2_decap_8 FILLER_12_279 ();
 sg13g2_decap_8 FILLER_12_286 ();
 sg13g2_decap_8 FILLER_12_293 ();
 sg13g2_decap_4 FILLER_12_300 ();
 sg13g2_fill_2 FILLER_12_304 ();
 sg13g2_decap_8 FILLER_12_332 ();
 sg13g2_decap_8 FILLER_12_339 ();
 sg13g2_decap_8 FILLER_12_346 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_fill_2 FILLER_12_360 ();
 sg13g2_fill_1 FILLER_12_362 ();
 sg13g2_fill_1 FILLER_12_393 ();
 sg13g2_fill_1 FILLER_12_399 ();
 sg13g2_fill_1 FILLER_12_461 ();
 sg13g2_decap_8 FILLER_12_468 ();
 sg13g2_fill_2 FILLER_12_499 ();
 sg13g2_decap_4 FILLER_12_543 ();
 sg13g2_fill_2 FILLER_12_547 ();
 sg13g2_decap_8 FILLER_12_585 ();
 sg13g2_fill_1 FILLER_12_592 ();
 sg13g2_decap_8 FILLER_12_638 ();
 sg13g2_fill_2 FILLER_12_645 ();
 sg13g2_fill_1 FILLER_12_647 ();
 sg13g2_fill_1 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_688 ();
 sg13g2_fill_1 FILLER_12_695 ();
 sg13g2_decap_4 FILLER_12_731 ();
 sg13g2_fill_1 FILLER_12_735 ();
 sg13g2_fill_2 FILLER_12_749 ();
 sg13g2_decap_4 FILLER_12_801 ();
 sg13g2_fill_1 FILLER_12_805 ();
 sg13g2_fill_2 FILLER_12_862 ();
 sg13g2_fill_1 FILLER_12_864 ();
 sg13g2_fill_1 FILLER_12_936 ();
 sg13g2_fill_1 FILLER_12_961 ();
 sg13g2_decap_4 FILLER_12_970 ();
 sg13g2_fill_1 FILLER_12_974 ();
 sg13g2_fill_2 FILLER_12_1027 ();
 sg13g2_decap_8 FILLER_12_1109 ();
 sg13g2_fill_1 FILLER_12_1116 ();
 sg13g2_decap_4 FILLER_12_1126 ();
 sg13g2_fill_1 FILLER_12_1136 ();
 sg13g2_decap_8 FILLER_12_1140 ();
 sg13g2_decap_8 FILLER_12_1147 ();
 sg13g2_decap_8 FILLER_12_1167 ();
 sg13g2_decap_8 FILLER_12_1174 ();
 sg13g2_decap_4 FILLER_12_1181 ();
 sg13g2_fill_1 FILLER_12_1185 ();
 sg13g2_fill_2 FILLER_12_1212 ();
 sg13g2_fill_1 FILLER_12_1214 ();
 sg13g2_decap_8 FILLER_12_1261 ();
 sg13g2_decap_8 FILLER_12_1268 ();
 sg13g2_decap_8 FILLER_12_1275 ();
 sg13g2_fill_2 FILLER_12_1282 ();
 sg13g2_decap_8 FILLER_12_1295 ();
 sg13g2_decap_8 FILLER_12_1302 ();
 sg13g2_decap_4 FILLER_12_1309 ();
 sg13g2_decap_8 FILLER_12_1327 ();
 sg13g2_fill_1 FILLER_12_1334 ();
 sg13g2_decap_4 FILLER_12_1344 ();
 sg13g2_decap_8 FILLER_12_1356 ();
 sg13g2_fill_1 FILLER_12_1363 ();
 sg13g2_fill_2 FILLER_12_1372 ();
 sg13g2_fill_2 FILLER_12_1401 ();
 sg13g2_decap_8 FILLER_12_1407 ();
 sg13g2_decap_8 FILLER_12_1414 ();
 sg13g2_decap_8 FILLER_12_1421 ();
 sg13g2_fill_1 FILLER_12_1428 ();
 sg13g2_decap_8 FILLER_12_1433 ();
 sg13g2_decap_8 FILLER_12_1440 ();
 sg13g2_decap_8 FILLER_12_1447 ();
 sg13g2_fill_2 FILLER_12_1454 ();
 sg13g2_fill_1 FILLER_12_1501 ();
 sg13g2_fill_1 FILLER_12_1574 ();
 sg13g2_decap_8 FILLER_12_1601 ();
 sg13g2_decap_4 FILLER_12_1608 ();
 sg13g2_fill_2 FILLER_12_1612 ();
 sg13g2_decap_8 FILLER_12_1644 ();
 sg13g2_decap_8 FILLER_12_1651 ();
 sg13g2_decap_4 FILLER_12_1666 ();
 sg13g2_decap_8 FILLER_12_1674 ();
 sg13g2_decap_4 FILLER_12_1681 ();
 sg13g2_decap_8 FILLER_12_1729 ();
 sg13g2_decap_4 FILLER_12_1736 ();
 sg13g2_fill_1 FILLER_12_1749 ();
 sg13g2_fill_2 FILLER_12_1793 ();
 sg13g2_fill_2 FILLER_12_1826 ();
 sg13g2_fill_2 FILLER_12_1833 ();
 sg13g2_fill_1 FILLER_12_1835 ();
 sg13g2_fill_1 FILLER_12_1862 ();
 sg13g2_fill_1 FILLER_12_1889 ();
 sg13g2_fill_2 FILLER_12_1896 ();
 sg13g2_decap_4 FILLER_12_1924 ();
 sg13g2_fill_2 FILLER_12_1963 ();
 sg13g2_fill_1 FILLER_12_1965 ();
 sg13g2_fill_1 FILLER_12_2015 ();
 sg13g2_fill_2 FILLER_12_2021 ();
 sg13g2_fill_1 FILLER_12_2023 ();
 sg13g2_fill_2 FILLER_12_2028 ();
 sg13g2_decap_8 FILLER_12_2035 ();
 sg13g2_decap_8 FILLER_12_2042 ();
 sg13g2_decap_8 FILLER_12_2107 ();
 sg13g2_decap_8 FILLER_12_2123 ();
 sg13g2_decap_4 FILLER_12_2130 ();
 sg13g2_fill_1 FILLER_12_2139 ();
 sg13g2_fill_2 FILLER_12_2149 ();
 sg13g2_decap_8 FILLER_12_2219 ();
 sg13g2_decap_4 FILLER_12_2226 ();
 sg13g2_decap_4 FILLER_12_2234 ();
 sg13g2_fill_2 FILLER_12_2238 ();
 sg13g2_decap_8 FILLER_12_2244 ();
 sg13g2_decap_8 FILLER_12_2251 ();
 sg13g2_decap_8 FILLER_12_2258 ();
 sg13g2_decap_4 FILLER_12_2265 ();
 sg13g2_fill_2 FILLER_12_2269 ();
 sg13g2_fill_2 FILLER_12_2289 ();
 sg13g2_fill_1 FILLER_12_2296 ();
 sg13g2_decap_8 FILLER_12_2354 ();
 sg13g2_fill_1 FILLER_12_2361 ();
 sg13g2_decap_8 FILLER_12_2368 ();
 sg13g2_fill_2 FILLER_12_2378 ();
 sg13g2_fill_2 FILLER_12_2392 ();
 sg13g2_fill_1 FILLER_12_2394 ();
 sg13g2_decap_4 FILLER_12_2431 ();
 sg13g2_fill_2 FILLER_12_2441 ();
 sg13g2_decap_8 FILLER_12_2456 ();
 sg13g2_decap_8 FILLER_12_2463 ();
 sg13g2_decap_8 FILLER_12_2470 ();
 sg13g2_fill_2 FILLER_12_2477 ();
 sg13g2_fill_1 FILLER_12_2479 ();
 sg13g2_decap_8 FILLER_12_2517 ();
 sg13g2_decap_8 FILLER_12_2524 ();
 sg13g2_fill_2 FILLER_12_2531 ();
 sg13g2_fill_2 FILLER_12_2537 ();
 sg13g2_fill_1 FILLER_12_2539 ();
 sg13g2_decap_4 FILLER_12_2552 ();
 sg13g2_fill_1 FILLER_12_2556 ();
 sg13g2_decap_4 FILLER_12_2565 ();
 sg13g2_fill_2 FILLER_12_2569 ();
 sg13g2_decap_4 FILLER_12_2606 ();
 sg13g2_decap_8 FILLER_12_2614 ();
 sg13g2_decap_8 FILLER_12_2621 ();
 sg13g2_decap_8 FILLER_12_2628 ();
 sg13g2_decap_8 FILLER_12_2635 ();
 sg13g2_decap_8 FILLER_12_2642 ();
 sg13g2_decap_8 FILLER_12_2649 ();
 sg13g2_decap_8 FILLER_12_2656 ();
 sg13g2_decap_8 FILLER_12_2663 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_41 ();
 sg13g2_fill_1 FILLER_13_51 ();
 sg13g2_fill_1 FILLER_13_58 ();
 sg13g2_fill_1 FILLER_13_62 ();
 sg13g2_fill_1 FILLER_13_72 ();
 sg13g2_fill_2 FILLER_13_76 ();
 sg13g2_decap_8 FILLER_13_104 ();
 sg13g2_decap_8 FILLER_13_137 ();
 sg13g2_fill_2 FILLER_13_170 ();
 sg13g2_fill_1 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_204 ();
 sg13g2_decap_4 FILLER_13_211 ();
 sg13g2_decap_8 FILLER_13_251 ();
 sg13g2_decap_8 FILLER_13_258 ();
 sg13g2_fill_2 FILLER_13_265 ();
 sg13g2_decap_8 FILLER_13_293 ();
 sg13g2_decap_8 FILLER_13_300 ();
 sg13g2_decap_4 FILLER_13_307 ();
 sg13g2_fill_1 FILLER_13_311 ();
 sg13g2_decap_8 FILLER_13_338 ();
 sg13g2_fill_1 FILLER_13_345 ();
 sg13g2_fill_2 FILLER_13_372 ();
 sg13g2_fill_1 FILLER_13_374 ();
 sg13g2_fill_1 FILLER_13_395 ();
 sg13g2_fill_2 FILLER_13_402 ();
 sg13g2_fill_1 FILLER_13_419 ();
 sg13g2_fill_1 FILLER_13_424 ();
 sg13g2_fill_2 FILLER_13_462 ();
 sg13g2_decap_4 FILLER_13_468 ();
 sg13g2_fill_2 FILLER_13_472 ();
 sg13g2_decap_4 FILLER_13_478 ();
 sg13g2_fill_1 FILLER_13_482 ();
 sg13g2_fill_2 FILLER_13_487 ();
 sg13g2_fill_2 FILLER_13_530 ();
 sg13g2_decap_8 FILLER_13_535 ();
 sg13g2_fill_2 FILLER_13_542 ();
 sg13g2_decap_8 FILLER_13_575 ();
 sg13g2_decap_8 FILLER_13_582 ();
 sg13g2_decap_8 FILLER_13_589 ();
 sg13g2_decap_8 FILLER_13_596 ();
 sg13g2_decap_8 FILLER_13_603 ();
 sg13g2_decap_8 FILLER_13_610 ();
 sg13g2_decap_8 FILLER_13_617 ();
 sg13g2_decap_4 FILLER_13_624 ();
 sg13g2_fill_2 FILLER_13_628 ();
 sg13g2_decap_4 FILLER_13_634 ();
 sg13g2_decap_4 FILLER_13_642 ();
 sg13g2_fill_2 FILLER_13_646 ();
 sg13g2_fill_2 FILLER_13_661 ();
 sg13g2_decap_4 FILLER_13_690 ();
 sg13g2_fill_2 FILLER_13_697 ();
 sg13g2_decap_8 FILLER_13_717 ();
 sg13g2_decap_8 FILLER_13_724 ();
 sg13g2_decap_8 FILLER_13_731 ();
 sg13g2_decap_8 FILLER_13_738 ();
 sg13g2_decap_8 FILLER_13_745 ();
 sg13g2_fill_2 FILLER_13_752 ();
 sg13g2_fill_1 FILLER_13_754 ();
 sg13g2_fill_2 FILLER_13_763 ();
 sg13g2_fill_2 FILLER_13_787 ();
 sg13g2_fill_1 FILLER_13_789 ();
 sg13g2_decap_8 FILLER_13_800 ();
 sg13g2_fill_2 FILLER_13_807 ();
 sg13g2_decap_8 FILLER_13_862 ();
 sg13g2_decap_4 FILLER_13_869 ();
 sg13g2_fill_2 FILLER_13_873 ();
 sg13g2_fill_1 FILLER_13_879 ();
 sg13g2_decap_4 FILLER_13_888 ();
 sg13g2_fill_1 FILLER_13_892 ();
 sg13g2_fill_1 FILLER_13_906 ();
 sg13g2_fill_2 FILLER_13_933 ();
 sg13g2_fill_1 FILLER_13_935 ();
 sg13g2_fill_2 FILLER_13_942 ();
 sg13g2_fill_1 FILLER_13_944 ();
 sg13g2_decap_4 FILLER_13_961 ();
 sg13g2_fill_2 FILLER_13_965 ();
 sg13g2_decap_4 FILLER_13_971 ();
 sg13g2_fill_2 FILLER_13_975 ();
 sg13g2_fill_2 FILLER_13_990 ();
 sg13g2_fill_2 FILLER_13_1030 ();
 sg13g2_decap_4 FILLER_13_1040 ();
 sg13g2_fill_1 FILLER_13_1044 ();
 sg13g2_fill_2 FILLER_13_1099 ();
 sg13g2_decap_8 FILLER_13_1118 ();
 sg13g2_fill_1 FILLER_13_1125 ();
 sg13g2_decap_8 FILLER_13_1157 ();
 sg13g2_decap_8 FILLER_13_1164 ();
 sg13g2_decap_8 FILLER_13_1171 ();
 sg13g2_decap_8 FILLER_13_1178 ();
 sg13g2_decap_8 FILLER_13_1185 ();
 sg13g2_decap_8 FILLER_13_1192 ();
 sg13g2_decap_4 FILLER_13_1208 ();
 sg13g2_fill_1 FILLER_13_1212 ();
 sg13g2_fill_1 FILLER_13_1225 ();
 sg13g2_fill_2 FILLER_13_1234 ();
 sg13g2_fill_1 FILLER_13_1236 ();
 sg13g2_fill_2 FILLER_13_1255 ();
 sg13g2_fill_1 FILLER_13_1257 ();
 sg13g2_fill_1 FILLER_13_1264 ();
 sg13g2_fill_2 FILLER_13_1322 ();
 sg13g2_decap_8 FILLER_13_1350 ();
 sg13g2_decap_8 FILLER_13_1357 ();
 sg13g2_decap_8 FILLER_13_1364 ();
 sg13g2_decap_8 FILLER_13_1371 ();
 sg13g2_fill_2 FILLER_13_1378 ();
 sg13g2_fill_1 FILLER_13_1380 ();
 sg13g2_fill_2 FILLER_13_1412 ();
 sg13g2_fill_1 FILLER_13_1414 ();
 sg13g2_decap_8 FILLER_13_1455 ();
 sg13g2_fill_1 FILLER_13_1534 ();
 sg13g2_fill_1 FILLER_13_1550 ();
 sg13g2_fill_2 FILLER_13_1573 ();
 sg13g2_decap_8 FILLER_13_1601 ();
 sg13g2_decap_8 FILLER_13_1608 ();
 sg13g2_fill_2 FILLER_13_1615 ();
 sg13g2_fill_1 FILLER_13_1617 ();
 sg13g2_decap_8 FILLER_13_1623 ();
 sg13g2_decap_8 FILLER_13_1678 ();
 sg13g2_decap_8 FILLER_13_1685 ();
 sg13g2_fill_1 FILLER_13_1705 ();
 sg13g2_fill_1 FILLER_13_1733 ();
 sg13g2_decap_8 FILLER_13_1755 ();
 sg13g2_decap_4 FILLER_13_1762 ();
 sg13g2_fill_1 FILLER_13_1766 ();
 sg13g2_fill_2 FILLER_13_1798 ();
 sg13g2_fill_1 FILLER_13_1804 ();
 sg13g2_fill_2 FILLER_13_1809 ();
 sg13g2_fill_1 FILLER_13_1811 ();
 sg13g2_fill_2 FILLER_13_1817 ();
 sg13g2_fill_1 FILLER_13_1819 ();
 sg13g2_decap_4 FILLER_13_1850 ();
 sg13g2_fill_2 FILLER_13_1854 ();
 sg13g2_fill_1 FILLER_13_1861 ();
 sg13g2_decap_4 FILLER_13_1875 ();
 sg13g2_fill_1 FILLER_13_1910 ();
 sg13g2_fill_2 FILLER_13_1915 ();
 sg13g2_decap_4 FILLER_13_1922 ();
 sg13g2_fill_2 FILLER_13_1926 ();
 sg13g2_decap_4 FILLER_13_1940 ();
 sg13g2_fill_1 FILLER_13_1944 ();
 sg13g2_fill_1 FILLER_13_1979 ();
 sg13g2_decap_4 FILLER_13_1986 ();
 sg13g2_fill_1 FILLER_13_1990 ();
 sg13g2_fill_2 FILLER_13_2047 ();
 sg13g2_fill_1 FILLER_13_2049 ();
 sg13g2_fill_1 FILLER_13_2055 ();
 sg13g2_fill_2 FILLER_13_2060 ();
 sg13g2_fill_2 FILLER_13_2074 ();
 sg13g2_fill_1 FILLER_13_2076 ();
 sg13g2_fill_1 FILLER_13_2134 ();
 sg13g2_fill_2 FILLER_13_2148 ();
 sg13g2_fill_2 FILLER_13_2164 ();
 sg13g2_fill_1 FILLER_13_2171 ();
 sg13g2_decap_8 FILLER_13_2176 ();
 sg13g2_fill_2 FILLER_13_2183 ();
 sg13g2_decap_8 FILLER_13_2189 ();
 sg13g2_fill_2 FILLER_13_2208 ();
 sg13g2_fill_1 FILLER_13_2210 ();
 sg13g2_fill_2 FILLER_13_2237 ();
 sg13g2_fill_2 FILLER_13_2244 ();
 sg13g2_decap_8 FILLER_13_2275 ();
 sg13g2_decap_4 FILLER_13_2282 ();
 sg13g2_decap_4 FILLER_13_2289 ();
 sg13g2_decap_4 FILLER_13_2315 ();
 sg13g2_fill_2 FILLER_13_2369 ();
 sg13g2_fill_1 FILLER_13_2371 ();
 sg13g2_decap_8 FILLER_13_2407 ();
 sg13g2_decap_4 FILLER_13_2414 ();
 sg13g2_fill_1 FILLER_13_2418 ();
 sg13g2_decap_4 FILLER_13_2450 ();
 sg13g2_fill_2 FILLER_13_2454 ();
 sg13g2_decap_8 FILLER_13_2460 ();
 sg13g2_fill_2 FILLER_13_2467 ();
 sg13g2_fill_1 FILLER_13_2469 ();
 sg13g2_decap_8 FILLER_13_2483 ();
 sg13g2_fill_2 FILLER_13_2490 ();
 sg13g2_fill_1 FILLER_13_2492 ();
 sg13g2_decap_8 FILLER_13_2535 ();
 sg13g2_decap_8 FILLER_13_2542 ();
 sg13g2_decap_8 FILLER_13_2549 ();
 sg13g2_decap_8 FILLER_13_2556 ();
 sg13g2_decap_8 FILLER_13_2563 ();
 sg13g2_decap_8 FILLER_13_2570 ();
 sg13g2_decap_4 FILLER_13_2577 ();
 sg13g2_fill_1 FILLER_13_2581 ();
 sg13g2_decap_4 FILLER_13_2604 ();
 sg13g2_fill_2 FILLER_13_2608 ();
 sg13g2_decap_8 FILLER_13_2636 ();
 sg13g2_decap_8 FILLER_13_2643 ();
 sg13g2_decap_8 FILLER_13_2650 ();
 sg13g2_decap_8 FILLER_13_2657 ();
 sg13g2_decap_4 FILLER_13_2664 ();
 sg13g2_fill_2 FILLER_13_2668 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_7 ();
 sg13g2_fill_1 FILLER_14_36 ();
 sg13g2_fill_1 FILLER_14_43 ();
 sg13g2_decap_8 FILLER_14_78 ();
 sg13g2_decap_8 FILLER_14_85 ();
 sg13g2_decap_8 FILLER_14_92 ();
 sg13g2_decap_8 FILLER_14_99 ();
 sg13g2_decap_8 FILLER_14_106 ();
 sg13g2_fill_2 FILLER_14_113 ();
 sg13g2_fill_1 FILLER_14_115 ();
 sg13g2_decap_8 FILLER_14_142 ();
 sg13g2_fill_2 FILLER_14_149 ();
 sg13g2_decap_4 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_207 ();
 sg13g2_fill_1 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_251 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_decap_8 FILLER_14_290 ();
 sg13g2_decap_8 FILLER_14_297 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_fill_1 FILLER_14_311 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_fill_2 FILLER_14_361 ();
 sg13g2_fill_1 FILLER_14_363 ();
 sg13g2_decap_4 FILLER_14_373 ();
 sg13g2_fill_2 FILLER_14_377 ();
 sg13g2_fill_2 FILLER_14_384 ();
 sg13g2_fill_2 FILLER_14_392 ();
 sg13g2_fill_2 FILLER_14_399 ();
 sg13g2_fill_1 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_415 ();
 sg13g2_fill_2 FILLER_14_422 ();
 sg13g2_fill_1 FILLER_14_450 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_fill_2 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_467 ();
 sg13g2_decap_4 FILLER_14_484 ();
 sg13g2_fill_1 FILLER_14_488 ();
 sg13g2_fill_2 FILLER_14_493 ();
 sg13g2_decap_4 FILLER_14_499 ();
 sg13g2_decap_8 FILLER_14_538 ();
 sg13g2_decap_8 FILLER_14_545 ();
 sg13g2_decap_8 FILLER_14_552 ();
 sg13g2_decap_8 FILLER_14_559 ();
 sg13g2_decap_8 FILLER_14_566 ();
 sg13g2_decap_8 FILLER_14_573 ();
 sg13g2_decap_8 FILLER_14_580 ();
 sg13g2_fill_1 FILLER_14_587 ();
 sg13g2_decap_8 FILLER_14_610 ();
 sg13g2_decap_8 FILLER_14_617 ();
 sg13g2_decap_8 FILLER_14_624 ();
 sg13g2_fill_2 FILLER_14_631 ();
 sg13g2_decap_4 FILLER_14_650 ();
 sg13g2_fill_1 FILLER_14_654 ();
 sg13g2_fill_1 FILLER_14_660 ();
 sg13g2_fill_2 FILLER_14_666 ();
 sg13g2_fill_2 FILLER_14_691 ();
 sg13g2_fill_2 FILLER_14_701 ();
 sg13g2_decap_4 FILLER_14_726 ();
 sg13g2_fill_2 FILLER_14_756 ();
 sg13g2_fill_1 FILLER_14_758 ();
 sg13g2_decap_8 FILLER_14_794 ();
 sg13g2_decap_8 FILLER_14_801 ();
 sg13g2_fill_1 FILLER_14_808 ();
 sg13g2_decap_4 FILLER_14_813 ();
 sg13g2_decap_8 FILLER_14_830 ();
 sg13g2_decap_8 FILLER_14_837 ();
 sg13g2_decap_8 FILLER_14_844 ();
 sg13g2_decap_4 FILLER_14_851 ();
 sg13g2_fill_2 FILLER_14_855 ();
 sg13g2_decap_8 FILLER_14_870 ();
 sg13g2_fill_1 FILLER_14_877 ();
 sg13g2_decap_4 FILLER_14_883 ();
 sg13g2_fill_2 FILLER_14_887 ();
 sg13g2_fill_1 FILLER_14_902 ();
 sg13g2_fill_1 FILLER_14_916 ();
 sg13g2_decap_4 FILLER_14_921 ();
 sg13g2_fill_2 FILLER_14_929 ();
 sg13g2_fill_1 FILLER_14_931 ();
 sg13g2_decap_8 FILLER_14_938 ();
 sg13g2_fill_1 FILLER_14_945 ();
 sg13g2_fill_1 FILLER_14_972 ();
 sg13g2_decap_4 FILLER_14_981 ();
 sg13g2_fill_1 FILLER_14_1019 ();
 sg13g2_fill_2 FILLER_14_1028 ();
 sg13g2_fill_1 FILLER_14_1039 ();
 sg13g2_fill_1 FILLER_14_1066 ();
 sg13g2_fill_2 FILLER_14_1125 ();
 sg13g2_fill_1 FILLER_14_1127 ();
 sg13g2_fill_2 FILLER_14_1140 ();
 sg13g2_fill_1 FILLER_14_1142 ();
 sg13g2_fill_2 FILLER_14_1173 ();
 sg13g2_decap_4 FILLER_14_1180 ();
 sg13g2_fill_1 FILLER_14_1184 ();
 sg13g2_decap_8 FILLER_14_1189 ();
 sg13g2_fill_1 FILLER_14_1196 ();
 sg13g2_fill_2 FILLER_14_1201 ();
 sg13g2_decap_4 FILLER_14_1207 ();
 sg13g2_fill_2 FILLER_14_1215 ();
 sg13g2_decap_8 FILLER_14_1229 ();
 sg13g2_decap_4 FILLER_14_1270 ();
 sg13g2_fill_1 FILLER_14_1274 ();
 sg13g2_decap_8 FILLER_14_1297 ();
 sg13g2_decap_8 FILLER_14_1304 ();
 sg13g2_decap_8 FILLER_14_1311 ();
 sg13g2_decap_4 FILLER_14_1318 ();
 sg13g2_decap_8 FILLER_14_1327 ();
 sg13g2_decap_4 FILLER_14_1334 ();
 sg13g2_fill_1 FILLER_14_1338 ();
 sg13g2_decap_8 FILLER_14_1343 ();
 sg13g2_decap_8 FILLER_14_1350 ();
 sg13g2_decap_8 FILLER_14_1357 ();
 sg13g2_fill_2 FILLER_14_1364 ();
 sg13g2_fill_1 FILLER_14_1366 ();
 sg13g2_decap_8 FILLER_14_1378 ();
 sg13g2_fill_2 FILLER_14_1385 ();
 sg13g2_fill_1 FILLER_14_1394 ();
 sg13g2_decap_4 FILLER_14_1433 ();
 sg13g2_fill_2 FILLER_14_1437 ();
 sg13g2_fill_2 FILLER_14_1471 ();
 sg13g2_decap_8 FILLER_14_1506 ();
 sg13g2_fill_1 FILLER_14_1557 ();
 sg13g2_fill_1 FILLER_14_1561 ();
 sg13g2_decap_8 FILLER_14_1578 ();
 sg13g2_fill_1 FILLER_14_1591 ();
 sg13g2_decap_8 FILLER_14_1601 ();
 sg13g2_fill_1 FILLER_14_1608 ();
 sg13g2_fill_1 FILLER_14_1661 ();
 sg13g2_fill_2 FILLER_14_1665 ();
 sg13g2_fill_2 FILLER_14_1693 ();
 sg13g2_fill_1 FILLER_14_1706 ();
 sg13g2_fill_2 FILLER_14_1734 ();
 sg13g2_decap_8 FILLER_14_1740 ();
 sg13g2_decap_8 FILLER_14_1747 ();
 sg13g2_decap_8 FILLER_14_1754 ();
 sg13g2_decap_8 FILLER_14_1761 ();
 sg13g2_fill_2 FILLER_14_1768 ();
 sg13g2_fill_1 FILLER_14_1778 ();
 sg13g2_fill_2 FILLER_14_1783 ();
 sg13g2_decap_8 FILLER_14_1814 ();
 sg13g2_decap_8 FILLER_14_1821 ();
 sg13g2_decap_8 FILLER_14_1828 ();
 sg13g2_fill_2 FILLER_14_1835 ();
 sg13g2_fill_1 FILLER_14_1837 ();
 sg13g2_decap_8 FILLER_14_1843 ();
 sg13g2_fill_1 FILLER_14_1850 ();
 sg13g2_fill_2 FILLER_14_1886 ();
 sg13g2_fill_1 FILLER_14_1888 ();
 sg13g2_fill_2 FILLER_14_1899 ();
 sg13g2_fill_1 FILLER_14_1901 ();
 sg13g2_decap_8 FILLER_14_1906 ();
 sg13g2_decap_4 FILLER_14_1913 ();
 sg13g2_fill_1 FILLER_14_1947 ();
 sg13g2_fill_1 FILLER_14_1974 ();
 sg13g2_decap_8 FILLER_14_1984 ();
 sg13g2_decap_4 FILLER_14_1991 ();
 sg13g2_decap_8 FILLER_14_2000 ();
 sg13g2_decap_8 FILLER_14_2007 ();
 sg13g2_decap_8 FILLER_14_2014 ();
 sg13g2_decap_8 FILLER_14_2021 ();
 sg13g2_decap_4 FILLER_14_2028 ();
 sg13g2_fill_1 FILLER_14_2032 ();
 sg13g2_decap_4 FILLER_14_2037 ();
 sg13g2_fill_1 FILLER_14_2041 ();
 sg13g2_decap_4 FILLER_14_2051 ();
 sg13g2_fill_1 FILLER_14_2071 ();
 sg13g2_fill_2 FILLER_14_2092 ();
 sg13g2_fill_1 FILLER_14_2094 ();
 sg13g2_fill_2 FILLER_14_2105 ();
 sg13g2_fill_1 FILLER_14_2107 ();
 sg13g2_fill_2 FILLER_14_2134 ();
 sg13g2_fill_2 FILLER_14_2162 ();
 sg13g2_decap_8 FILLER_14_2179 ();
 sg13g2_decap_8 FILLER_14_2186 ();
 sg13g2_decap_8 FILLER_14_2193 ();
 sg13g2_decap_4 FILLER_14_2213 ();
 sg13g2_decap_4 FILLER_14_2262 ();
 sg13g2_fill_1 FILLER_14_2266 ();
 sg13g2_fill_1 FILLER_14_2293 ();
 sg13g2_decap_8 FILLER_14_2331 ();
 sg13g2_decap_8 FILLER_14_2338 ();
 sg13g2_decap_8 FILLER_14_2345 ();
 sg13g2_decap_8 FILLER_14_2352 ();
 sg13g2_decap_4 FILLER_14_2359 ();
 sg13g2_fill_1 FILLER_14_2363 ();
 sg13g2_fill_1 FILLER_14_2420 ();
 sg13g2_fill_2 FILLER_14_2447 ();
 sg13g2_fill_1 FILLER_14_2490 ();
 sg13g2_decap_8 FILLER_14_2495 ();
 sg13g2_decap_8 FILLER_14_2502 ();
 sg13g2_decap_8 FILLER_14_2509 ();
 sg13g2_decap_8 FILLER_14_2516 ();
 sg13g2_decap_8 FILLER_14_2523 ();
 sg13g2_fill_1 FILLER_14_2530 ();
 sg13g2_decap_8 FILLER_14_2557 ();
 sg13g2_decap_8 FILLER_14_2564 ();
 sg13g2_decap_8 FILLER_14_2571 ();
 sg13g2_decap_8 FILLER_14_2578 ();
 sg13g2_fill_1 FILLER_14_2594 ();
 sg13g2_decap_8 FILLER_14_2621 ();
 sg13g2_decap_8 FILLER_14_2628 ();
 sg13g2_decap_8 FILLER_14_2635 ();
 sg13g2_decap_8 FILLER_14_2642 ();
 sg13g2_decap_8 FILLER_14_2649 ();
 sg13g2_decap_8 FILLER_14_2656 ();
 sg13g2_decap_8 FILLER_14_2663 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_fill_2 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_41 ();
 sg13g2_decap_8 FILLER_15_80 ();
 sg13g2_decap_8 FILLER_15_87 ();
 sg13g2_decap_8 FILLER_15_102 ();
 sg13g2_decap_8 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_fill_2 FILLER_15_123 ();
 sg13g2_fill_1 FILLER_15_125 ();
 sg13g2_fill_2 FILLER_15_172 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_fill_1 FILLER_15_179 ();
 sg13g2_fill_2 FILLER_15_183 ();
 sg13g2_fill_2 FILLER_15_195 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_fill_1 FILLER_15_204 ();
 sg13g2_fill_2 FILLER_15_231 ();
 sg13g2_fill_1 FILLER_15_233 ();
 sg13g2_decap_8 FILLER_15_243 ();
 sg13g2_fill_2 FILLER_15_270 ();
 sg13g2_fill_1 FILLER_15_294 ();
 sg13g2_fill_2 FILLER_15_302 ();
 sg13g2_fill_1 FILLER_15_304 ();
 sg13g2_fill_2 FILLER_15_309 ();
 sg13g2_fill_1 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_331 ();
 sg13g2_decap_8 FILLER_15_338 ();
 sg13g2_decap_8 FILLER_15_345 ();
 sg13g2_fill_2 FILLER_15_352 ();
 sg13g2_fill_2 FILLER_15_400 ();
 sg13g2_decap_4 FILLER_15_408 ();
 sg13g2_fill_2 FILLER_15_412 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_8 FILLER_15_424 ();
 sg13g2_fill_1 FILLER_15_440 ();
 sg13g2_decap_8 FILLER_15_447 ();
 sg13g2_fill_2 FILLER_15_454 ();
 sg13g2_fill_1 FILLER_15_456 ();
 sg13g2_fill_1 FILLER_15_464 ();
 sg13g2_decap_8 FILLER_15_500 ();
 sg13g2_decap_8 FILLER_15_507 ();
 sg13g2_decap_8 FILLER_15_519 ();
 sg13g2_decap_4 FILLER_15_526 ();
 sg13g2_fill_2 FILLER_15_530 ();
 sg13g2_fill_1 FILLER_15_558 ();
 sg13g2_fill_1 FILLER_15_589 ();
 sg13g2_fill_2 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_fill_2 FILLER_15_630 ();
 sg13g2_fill_1 FILLER_15_632 ();
 sg13g2_fill_2 FILLER_15_641 ();
 sg13g2_decap_8 FILLER_15_648 ();
 sg13g2_decap_4 FILLER_15_655 ();
 sg13g2_fill_1 FILLER_15_663 ();
 sg13g2_fill_1 FILLER_15_668 ();
 sg13g2_fill_1 FILLER_15_690 ();
 sg13g2_fill_1 FILLER_15_699 ();
 sg13g2_fill_1 FILLER_15_705 ();
 sg13g2_decap_8 FILLER_15_711 ();
 sg13g2_fill_1 FILLER_15_718 ();
 sg13g2_decap_8 FILLER_15_741 ();
 sg13g2_fill_1 FILLER_15_748 ();
 sg13g2_decap_4 FILLER_15_754 ();
 sg13g2_fill_1 FILLER_15_793 ();
 sg13g2_fill_1 FILLER_15_824 ();
 sg13g2_decap_8 FILLER_15_830 ();
 sg13g2_decap_8 FILLER_15_837 ();
 sg13g2_decap_4 FILLER_15_844 ();
 sg13g2_fill_2 FILLER_15_848 ();
 sg13g2_decap_8 FILLER_15_860 ();
 sg13g2_fill_1 FILLER_15_867 ();
 sg13g2_fill_1 FILLER_15_882 ();
 sg13g2_fill_2 FILLER_15_892 ();
 sg13g2_decap_4 FILLER_15_899 ();
 sg13g2_decap_4 FILLER_15_908 ();
 sg13g2_fill_1 FILLER_15_912 ();
 sg13g2_decap_8 FILLER_15_917 ();
 sg13g2_decap_8 FILLER_15_924 ();
 sg13g2_fill_1 FILLER_15_931 ();
 sg13g2_fill_1 FILLER_15_968 ();
 sg13g2_decap_8 FILLER_15_990 ();
 sg13g2_fill_2 FILLER_15_997 ();
 sg13g2_fill_1 FILLER_15_999 ();
 sg13g2_fill_2 FILLER_15_1040 ();
 sg13g2_fill_1 FILLER_15_1042 ();
 sg13g2_fill_1 FILLER_15_1049 ();
 sg13g2_decap_4 FILLER_15_1056 ();
 sg13g2_fill_2 FILLER_15_1066 ();
 sg13g2_decap_4 FILLER_15_1093 ();
 sg13g2_fill_2 FILLER_15_1101 ();
 sg13g2_fill_1 FILLER_15_1134 ();
 sg13g2_decap_4 FILLER_15_1144 ();
 sg13g2_fill_2 FILLER_15_1148 ();
 sg13g2_decap_4 FILLER_15_1154 ();
 sg13g2_fill_2 FILLER_15_1158 ();
 sg13g2_decap_4 FILLER_15_1166 ();
 sg13g2_decap_8 FILLER_15_1232 ();
 sg13g2_fill_2 FILLER_15_1239 ();
 sg13g2_fill_1 FILLER_15_1241 ();
 sg13g2_decap_4 FILLER_15_1252 ();
 sg13g2_fill_2 FILLER_15_1264 ();
 sg13g2_fill_1 FILLER_15_1266 ();
 sg13g2_decap_8 FILLER_15_1308 ();
 sg13g2_fill_2 FILLER_15_1324 ();
 sg13g2_fill_1 FILLER_15_1326 ();
 sg13g2_fill_1 FILLER_15_1358 ();
 sg13g2_fill_2 FILLER_15_1425 ();
 sg13g2_fill_2 FILLER_15_1448 ();
 sg13g2_decap_4 FILLER_15_1456 ();
 sg13g2_fill_2 FILLER_15_1460 ();
 sg13g2_decap_4 FILLER_15_1488 ();
 sg13g2_decap_8 FILLER_15_1498 ();
 sg13g2_decap_8 FILLER_15_1505 ();
 sg13g2_decap_4 FILLER_15_1512 ();
 sg13g2_fill_1 FILLER_15_1525 ();
 sg13g2_fill_1 FILLER_15_1541 ();
 sg13g2_fill_2 FILLER_15_1592 ();
 sg13g2_fill_1 FILLER_15_1594 ();
 sg13g2_decap_8 FILLER_15_1607 ();
 sg13g2_decap_4 FILLER_15_1614 ();
 sg13g2_fill_1 FILLER_15_1618 ();
 sg13g2_decap_8 FILLER_15_1623 ();
 sg13g2_fill_1 FILLER_15_1630 ();
 sg13g2_decap_8 FILLER_15_1645 ();
 sg13g2_decap_4 FILLER_15_1652 ();
 sg13g2_fill_2 FILLER_15_1679 ();
 sg13g2_fill_2 FILLER_15_1688 ();
 sg13g2_decap_8 FILLER_15_1697 ();
 sg13g2_decap_8 FILLER_15_1704 ();
 sg13g2_decap_8 FILLER_15_1711 ();
 sg13g2_fill_2 FILLER_15_1718 ();
 sg13g2_fill_1 FILLER_15_1720 ();
 sg13g2_fill_2 FILLER_15_1727 ();
 sg13g2_decap_8 FILLER_15_1755 ();
 sg13g2_decap_8 FILLER_15_1762 ();
 sg13g2_decap_4 FILLER_15_1769 ();
 sg13g2_fill_2 FILLER_15_1773 ();
 sg13g2_decap_4 FILLER_15_1809 ();
 sg13g2_decap_8 FILLER_15_1822 ();
 sg13g2_decap_8 FILLER_15_1829 ();
 sg13g2_fill_1 FILLER_15_1836 ();
 sg13g2_decap_8 FILLER_15_1863 ();
 sg13g2_decap_4 FILLER_15_1870 ();
 sg13g2_fill_1 FILLER_15_1879 ();
 sg13g2_decap_8 FILLER_15_1884 ();
 sg13g2_fill_2 FILLER_15_1891 ();
 sg13g2_decap_8 FILLER_15_1914 ();
 sg13g2_decap_4 FILLER_15_1921 ();
 sg13g2_fill_1 FILLER_15_1925 ();
 sg13g2_decap_8 FILLER_15_1936 ();
 sg13g2_decap_8 FILLER_15_1943 ();
 sg13g2_fill_2 FILLER_15_1950 ();
 sg13g2_fill_1 FILLER_15_1952 ();
 sg13g2_fill_2 FILLER_15_1984 ();
 sg13g2_fill_1 FILLER_15_1986 ();
 sg13g2_fill_2 FILLER_15_1996 ();
 sg13g2_decap_8 FILLER_15_2003 ();
 sg13g2_decap_8 FILLER_15_2010 ();
 sg13g2_decap_8 FILLER_15_2017 ();
 sg13g2_decap_8 FILLER_15_2024 ();
 sg13g2_fill_2 FILLER_15_2031 ();
 sg13g2_decap_8 FILLER_15_2048 ();
 sg13g2_decap_8 FILLER_15_2055 ();
 sg13g2_decap_8 FILLER_15_2062 ();
 sg13g2_fill_2 FILLER_15_2069 ();
 sg13g2_fill_1 FILLER_15_2074 ();
 sg13g2_decap_8 FILLER_15_2097 ();
 sg13g2_decap_4 FILLER_15_2104 ();
 sg13g2_fill_2 FILLER_15_2117 ();
 sg13g2_fill_1 FILLER_15_2145 ();
 sg13g2_fill_1 FILLER_15_2192 ();
 sg13g2_decap_8 FILLER_15_2197 ();
 sg13g2_fill_2 FILLER_15_2204 ();
 sg13g2_fill_1 FILLER_15_2206 ();
 sg13g2_fill_2 FILLER_15_2210 ();
 sg13g2_fill_1 FILLER_15_2212 ();
 sg13g2_decap_4 FILLER_15_2242 ();
 sg13g2_fill_2 FILLER_15_2284 ();
 sg13g2_fill_2 FILLER_15_2295 ();
 sg13g2_fill_1 FILLER_15_2337 ();
 sg13g2_fill_2 FILLER_15_2343 ();
 sg13g2_fill_2 FILLER_15_2349 ();
 sg13g2_fill_1 FILLER_15_2357 ();
 sg13g2_fill_2 FILLER_15_2364 ();
 sg13g2_fill_2 FILLER_15_2371 ();
 sg13g2_fill_2 FILLER_15_2377 ();
 sg13g2_fill_1 FILLER_15_2420 ();
 sg13g2_fill_1 FILLER_15_2427 ();
 sg13g2_decap_4 FILLER_15_2433 ();
 sg13g2_fill_1 FILLER_15_2437 ();
 sg13g2_decap_8 FILLER_15_2442 ();
 sg13g2_fill_2 FILLER_15_2449 ();
 sg13g2_fill_1 FILLER_15_2451 ();
 sg13g2_fill_2 FILLER_15_2462 ();
 sg13g2_fill_1 FILLER_15_2464 ();
 sg13g2_fill_1 FILLER_15_2469 ();
 sg13g2_fill_2 FILLER_15_2478 ();
 sg13g2_fill_1 FILLER_15_2480 ();
 sg13g2_fill_1 FILLER_15_2490 ();
 sg13g2_decap_8 FILLER_15_2539 ();
 sg13g2_fill_1 FILLER_15_2546 ();
 sg13g2_decap_4 FILLER_15_2582 ();
 sg13g2_decap_8 FILLER_15_2604 ();
 sg13g2_decap_8 FILLER_15_2611 ();
 sg13g2_decap_8 FILLER_15_2618 ();
 sg13g2_decap_8 FILLER_15_2625 ();
 sg13g2_decap_8 FILLER_15_2632 ();
 sg13g2_decap_8 FILLER_15_2639 ();
 sg13g2_decap_8 FILLER_15_2646 ();
 sg13g2_decap_8 FILLER_15_2653 ();
 sg13g2_decap_8 FILLER_15_2660 ();
 sg13g2_fill_2 FILLER_15_2667 ();
 sg13g2_fill_1 FILLER_15_2669 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_16 ();
 sg13g2_fill_2 FILLER_16_25 ();
 sg13g2_fill_2 FILLER_16_33 ();
 sg13g2_fill_2 FILLER_16_43 ();
 sg13g2_fill_1 FILLER_16_45 ();
 sg13g2_decap_8 FILLER_16_78 ();
 sg13g2_decap_4 FILLER_16_85 ();
 sg13g2_fill_2 FILLER_16_89 ();
 sg13g2_decap_8 FILLER_16_117 ();
 sg13g2_decap_8 FILLER_16_124 ();
 sg13g2_decap_8 FILLER_16_131 ();
 sg13g2_decap_8 FILLER_16_138 ();
 sg13g2_decap_8 FILLER_16_145 ();
 sg13g2_decap_8 FILLER_16_152 ();
 sg13g2_decap_8 FILLER_16_159 ();
 sg13g2_decap_8 FILLER_16_166 ();
 sg13g2_decap_8 FILLER_16_173 ();
 sg13g2_decap_8 FILLER_16_180 ();
 sg13g2_fill_2 FILLER_16_187 ();
 sg13g2_fill_2 FILLER_16_194 ();
 sg13g2_fill_1 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_fill_2 FILLER_16_221 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_decap_4 FILLER_16_258 ();
 sg13g2_fill_1 FILLER_16_262 ();
 sg13g2_fill_2 FILLER_16_268 ();
 sg13g2_decap_8 FILLER_16_316 ();
 sg13g2_decap_8 FILLER_16_323 ();
 sg13g2_fill_1 FILLER_16_330 ();
 sg13g2_decap_8 FILLER_16_340 ();
 sg13g2_decap_8 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_fill_2 FILLER_16_361 ();
 sg13g2_fill_1 FILLER_16_363 ();
 sg13g2_fill_2 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_fill_1 FILLER_16_388 ();
 sg13g2_decap_4 FILLER_16_406 ();
 sg13g2_fill_2 FILLER_16_410 ();
 sg13g2_decap_8 FILLER_16_443 ();
 sg13g2_decap_8 FILLER_16_450 ();
 sg13g2_decap_8 FILLER_16_457 ();
 sg13g2_decap_8 FILLER_16_464 ();
 sg13g2_fill_2 FILLER_16_471 ();
 sg13g2_fill_1 FILLER_16_473 ();
 sg13g2_decap_4 FILLER_16_480 ();
 sg13g2_fill_1 FILLER_16_484 ();
 sg13g2_fill_1 FILLER_16_495 ();
 sg13g2_fill_2 FILLER_16_501 ();
 sg13g2_fill_1 FILLER_16_507 ();
 sg13g2_fill_1 FILLER_16_512 ();
 sg13g2_fill_1 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_524 ();
 sg13g2_decap_8 FILLER_16_531 ();
 sg13g2_decap_8 FILLER_16_538 ();
 sg13g2_decap_4 FILLER_16_550 ();
 sg13g2_fill_2 FILLER_16_554 ();
 sg13g2_decap_8 FILLER_16_561 ();
 sg13g2_decap_8 FILLER_16_568 ();
 sg13g2_decap_8 FILLER_16_575 ();
 sg13g2_decap_4 FILLER_16_582 ();
 sg13g2_fill_1 FILLER_16_586 ();
 sg13g2_decap_8 FILLER_16_592 ();
 sg13g2_decap_4 FILLER_16_608 ();
 sg13g2_fill_2 FILLER_16_612 ();
 sg13g2_decap_4 FILLER_16_619 ();
 sg13g2_fill_2 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_633 ();
 sg13g2_decap_8 FILLER_16_640 ();
 sg13g2_decap_8 FILLER_16_647 ();
 sg13g2_decap_4 FILLER_16_654 ();
 sg13g2_fill_1 FILLER_16_658 ();
 sg13g2_fill_2 FILLER_16_674 ();
 sg13g2_fill_1 FILLER_16_676 ();
 sg13g2_decap_8 FILLER_16_691 ();
 sg13g2_decap_4 FILLER_16_698 ();
 sg13g2_fill_2 FILLER_16_702 ();
 sg13g2_decap_4 FILLER_16_708 ();
 sg13g2_fill_1 FILLER_16_743 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_fill_2 FILLER_16_763 ();
 sg13g2_fill_1 FILLER_16_765 ();
 sg13g2_decap_4 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_778 ();
 sg13g2_fill_1 FILLER_16_785 ();
 sg13g2_decap_8 FILLER_16_792 ();
 sg13g2_decap_8 FILLER_16_799 ();
 sg13g2_fill_1 FILLER_16_806 ();
 sg13g2_fill_1 FILLER_16_841 ();
 sg13g2_fill_2 FILLER_16_848 ();
 sg13g2_fill_2 FILLER_16_871 ();
 sg13g2_fill_2 FILLER_16_899 ();
 sg13g2_fill_1 FILLER_16_901 ();
 sg13g2_decap_8 FILLER_16_907 ();
 sg13g2_decap_8 FILLER_16_914 ();
 sg13g2_decap_8 FILLER_16_921 ();
 sg13g2_decap_8 FILLER_16_928 ();
 sg13g2_fill_2 FILLER_16_935 ();
 sg13g2_decap_4 FILLER_16_946 ();
 sg13g2_fill_1 FILLER_16_950 ();
 sg13g2_fill_2 FILLER_16_959 ();
 sg13g2_fill_1 FILLER_16_961 ();
 sg13g2_decap_8 FILLER_16_991 ();
 sg13g2_decap_4 FILLER_16_998 ();
 sg13g2_fill_2 FILLER_16_1021 ();
 sg13g2_fill_1 FILLER_16_1023 ();
 sg13g2_fill_2 FILLER_16_1062 ();
 sg13g2_fill_1 FILLER_16_1064 ();
 sg13g2_fill_1 FILLER_16_1070 ();
 sg13g2_decap_8 FILLER_16_1076 ();
 sg13g2_decap_8 FILLER_16_1083 ();
 sg13g2_decap_4 FILLER_16_1090 ();
 sg13g2_fill_1 FILLER_16_1094 ();
 sg13g2_decap_8 FILLER_16_1108 ();
 sg13g2_fill_1 FILLER_16_1115 ();
 sg13g2_fill_1 FILLER_16_1122 ();
 sg13g2_decap_4 FILLER_16_1149 ();
 sg13g2_fill_2 FILLER_16_1174 ();
 sg13g2_fill_1 FILLER_16_1176 ();
 sg13g2_fill_2 FILLER_16_1267 ();
 sg13g2_decap_4 FILLER_16_1272 ();
 sg13g2_fill_1 FILLER_16_1276 ();
 sg13g2_fill_1 FILLER_16_1303 ();
 sg13g2_fill_2 FILLER_16_1310 ();
 sg13g2_fill_1 FILLER_16_1312 ();
 sg13g2_fill_2 FILLER_16_1339 ();
 sg13g2_fill_1 FILLER_16_1345 ();
 sg13g2_fill_1 FILLER_16_1351 ();
 sg13g2_fill_1 FILLER_16_1366 ();
 sg13g2_fill_2 FILLER_16_1384 ();
 sg13g2_fill_2 FILLER_16_1392 ();
 sg13g2_decap_8 FILLER_16_1434 ();
 sg13g2_fill_1 FILLER_16_1441 ();
 sg13g2_fill_1 FILLER_16_1445 ();
 sg13g2_decap_8 FILLER_16_1452 ();
 sg13g2_fill_1 FILLER_16_1463 ();
 sg13g2_fill_2 FILLER_16_1490 ();
 sg13g2_decap_8 FILLER_16_1499 ();
 sg13g2_decap_4 FILLER_16_1506 ();
 sg13g2_fill_1 FILLER_16_1519 ();
 sg13g2_fill_2 FILLER_16_1561 ();
 sg13g2_fill_1 FILLER_16_1572 ();
 sg13g2_fill_1 FILLER_16_1578 ();
 sg13g2_fill_2 FILLER_16_1635 ();
 sg13g2_fill_1 FILLER_16_1637 ();
 sg13g2_fill_2 FILLER_16_1680 ();
 sg13g2_fill_1 FILLER_16_1682 ();
 sg13g2_decap_4 FILLER_16_1709 ();
 sg13g2_fill_2 FILLER_16_1713 ();
 sg13g2_fill_1 FILLER_16_1745 ();
 sg13g2_decap_8 FILLER_16_1755 ();
 sg13g2_decap_8 FILLER_16_1762 ();
 sg13g2_decap_8 FILLER_16_1769 ();
 sg13g2_decap_4 FILLER_16_1776 ();
 sg13g2_fill_2 FILLER_16_1780 ();
 sg13g2_fill_1 FILLER_16_1791 ();
 sg13g2_decap_4 FILLER_16_1844 ();
 sg13g2_fill_1 FILLER_16_1848 ();
 sg13g2_decap_8 FILLER_16_1854 ();
 sg13g2_fill_2 FILLER_16_1861 ();
 sg13g2_fill_1 FILLER_16_1863 ();
 sg13g2_decap_8 FILLER_16_1890 ();
 sg13g2_decap_8 FILLER_16_1897 ();
 sg13g2_fill_2 FILLER_16_1904 ();
 sg13g2_fill_1 FILLER_16_1906 ();
 sg13g2_decap_8 FILLER_16_1922 ();
 sg13g2_decap_4 FILLER_16_1929 ();
 sg13g2_fill_1 FILLER_16_1933 ();
 sg13g2_decap_8 FILLER_16_1939 ();
 sg13g2_decap_8 FILLER_16_1946 ();
 sg13g2_decap_8 FILLER_16_1953 ();
 sg13g2_decap_4 FILLER_16_1964 ();
 sg13g2_fill_2 FILLER_16_1968 ();
 sg13g2_fill_2 FILLER_16_1979 ();
 sg13g2_fill_1 FILLER_16_1981 ();
 sg13g2_decap_8 FILLER_16_2013 ();
 sg13g2_decap_4 FILLER_16_2020 ();
 sg13g2_fill_2 FILLER_16_2024 ();
 sg13g2_decap_8 FILLER_16_2052 ();
 sg13g2_fill_2 FILLER_16_2059 ();
 sg13g2_fill_1 FILLER_16_2061 ();
 sg13g2_fill_1 FILLER_16_2071 ();
 sg13g2_decap_8 FILLER_16_2104 ();
 sg13g2_decap_8 FILLER_16_2111 ();
 sg13g2_fill_1 FILLER_16_2118 ();
 sg13g2_decap_8 FILLER_16_2128 ();
 sg13g2_decap_8 FILLER_16_2135 ();
 sg13g2_decap_8 FILLER_16_2142 ();
 sg13g2_fill_1 FILLER_16_2149 ();
 sg13g2_fill_2 FILLER_16_2179 ();
 sg13g2_fill_2 FILLER_16_2213 ();
 sg13g2_fill_1 FILLER_16_2220 ();
 sg13g2_fill_1 FILLER_16_2227 ();
 sg13g2_fill_1 FILLER_16_2232 ();
 sg13g2_decap_4 FILLER_16_2277 ();
 sg13g2_fill_2 FILLER_16_2281 ();
 sg13g2_fill_1 FILLER_16_2385 ();
 sg13g2_fill_2 FILLER_16_2395 ();
 sg13g2_fill_1 FILLER_16_2406 ();
 sg13g2_decap_8 FILLER_16_2437 ();
 sg13g2_decap_4 FILLER_16_2444 ();
 sg13g2_fill_1 FILLER_16_2448 ();
 sg13g2_fill_2 FILLER_16_2475 ();
 sg13g2_fill_1 FILLER_16_2477 ();
 sg13g2_decap_4 FILLER_16_2496 ();
 sg13g2_fill_1 FILLER_16_2500 ();
 sg13g2_decap_4 FILLER_16_2510 ();
 sg13g2_fill_1 FILLER_16_2514 ();
 sg13g2_decap_8 FILLER_16_2528 ();
 sg13g2_decap_8 FILLER_16_2535 ();
 sg13g2_fill_2 FILLER_16_2542 ();
 sg13g2_decap_8 FILLER_16_2549 ();
 sg13g2_decap_8 FILLER_16_2556 ();
 sg13g2_decap_4 FILLER_16_2563 ();
 sg13g2_fill_1 FILLER_16_2567 ();
 sg13g2_decap_8 FILLER_16_2635 ();
 sg13g2_decap_8 FILLER_16_2642 ();
 sg13g2_decap_8 FILLER_16_2649 ();
 sg13g2_decap_8 FILLER_16_2656 ();
 sg13g2_decap_8 FILLER_16_2663 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_45 ();
 sg13g2_fill_2 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_55 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_fill_2 FILLER_17_84 ();
 sg13g2_fill_1 FILLER_17_95 ();
 sg13g2_fill_1 FILLER_17_101 ();
 sg13g2_fill_1 FILLER_17_106 ();
 sg13g2_fill_1 FILLER_17_115 ();
 sg13g2_fill_2 FILLER_17_121 ();
 sg13g2_fill_1 FILLER_17_123 ();
 sg13g2_fill_1 FILLER_17_171 ();
 sg13g2_fill_2 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_281 ();
 sg13g2_decap_8 FILLER_17_288 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_4 FILLER_17_353 ();
 sg13g2_fill_1 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_4 FILLER_17_370 ();
 sg13g2_decap_4 FILLER_17_380 ();
 sg13g2_fill_2 FILLER_17_384 ();
 sg13g2_fill_1 FILLER_17_391 ();
 sg13g2_fill_2 FILLER_17_398 ();
 sg13g2_fill_1 FILLER_17_400 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_2 FILLER_17_408 ();
 sg13g2_decap_4 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_460 ();
 sg13g2_decap_4 FILLER_17_467 ();
 sg13g2_fill_1 FILLER_17_504 ();
 sg13g2_fill_2 FILLER_17_521 ();
 sg13g2_decap_8 FILLER_17_531 ();
 sg13g2_fill_1 FILLER_17_538 ();
 sg13g2_decap_8 FILLER_17_570 ();
 sg13g2_decap_8 FILLER_17_577 ();
 sg13g2_decap_8 FILLER_17_584 ();
 sg13g2_fill_2 FILLER_17_591 ();
 sg13g2_fill_1 FILLER_17_593 ();
 sg13g2_fill_2 FILLER_17_599 ();
 sg13g2_decap_8 FILLER_17_627 ();
 sg13g2_decap_8 FILLER_17_634 ();
 sg13g2_decap_8 FILLER_17_641 ();
 sg13g2_fill_2 FILLER_17_648 ();
 sg13g2_fill_1 FILLER_17_650 ();
 sg13g2_fill_2 FILLER_17_659 ();
 sg13g2_decap_8 FILLER_17_674 ();
 sg13g2_decap_4 FILLER_17_685 ();
 sg13g2_fill_2 FILLER_17_689 ();
 sg13g2_decap_4 FILLER_17_696 ();
 sg13g2_decap_8 FILLER_17_711 ();
 sg13g2_fill_1 FILLER_17_718 ();
 sg13g2_fill_1 FILLER_17_731 ();
 sg13g2_decap_8 FILLER_17_741 ();
 sg13g2_decap_8 FILLER_17_768 ();
 sg13g2_fill_1 FILLER_17_775 ();
 sg13g2_decap_8 FILLER_17_786 ();
 sg13g2_decap_8 FILLER_17_793 ();
 sg13g2_decap_8 FILLER_17_800 ();
 sg13g2_decap_8 FILLER_17_807 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_fill_2 FILLER_17_847 ();
 sg13g2_fill_1 FILLER_17_849 ();
 sg13g2_fill_2 FILLER_17_889 ();
 sg13g2_fill_1 FILLER_17_891 ();
 sg13g2_decap_8 FILLER_17_904 ();
 sg13g2_decap_4 FILLER_17_925 ();
 sg13g2_fill_1 FILLER_17_929 ();
 sg13g2_fill_2 FILLER_17_935 ();
 sg13g2_fill_1 FILLER_17_937 ();
 sg13g2_decap_8 FILLER_17_977 ();
 sg13g2_decap_4 FILLER_17_984 ();
 sg13g2_fill_2 FILLER_17_1022 ();
 sg13g2_fill_1 FILLER_17_1024 ();
 sg13g2_decap_8 FILLER_17_1068 ();
 sg13g2_decap_4 FILLER_17_1075 ();
 sg13g2_fill_1 FILLER_17_1079 ();
 sg13g2_fill_1 FILLER_17_1105 ();
 sg13g2_decap_4 FILLER_17_1130 ();
 sg13g2_decap_8 FILLER_17_1140 ();
 sg13g2_decap_4 FILLER_17_1147 ();
 sg13g2_fill_2 FILLER_17_1151 ();
 sg13g2_decap_8 FILLER_17_1198 ();
 sg13g2_decap_4 FILLER_17_1205 ();
 sg13g2_decap_8 FILLER_17_1214 ();
 sg13g2_decap_8 FILLER_17_1227 ();
 sg13g2_fill_2 FILLER_17_1234 ();
 sg13g2_decap_8 FILLER_17_1274 ();
 sg13g2_decap_8 FILLER_17_1281 ();
 sg13g2_decap_8 FILLER_17_1291 ();
 sg13g2_decap_8 FILLER_17_1298 ();
 sg13g2_fill_1 FILLER_17_1310 ();
 sg13g2_decap_4 FILLER_17_1319 ();
 sg13g2_fill_2 FILLER_17_1331 ();
 sg13g2_fill_1 FILLER_17_1333 ();
 sg13g2_decap_4 FILLER_17_1338 ();
 sg13g2_fill_1 FILLER_17_1342 ();
 sg13g2_fill_2 FILLER_17_1374 ();
 sg13g2_fill_1 FILLER_17_1382 ();
 sg13g2_fill_1 FILLER_17_1401 ();
 sg13g2_fill_2 FILLER_17_1414 ();
 sg13g2_fill_2 FILLER_17_1446 ();
 sg13g2_fill_1 FILLER_17_1448 ();
 sg13g2_fill_1 FILLER_17_1537 ();
 sg13g2_decap_8 FILLER_17_1554 ();
 sg13g2_fill_2 FILLER_17_1561 ();
 sg13g2_fill_1 FILLER_17_1566 ();
 sg13g2_fill_1 FILLER_17_1623 ();
 sg13g2_decap_8 FILLER_17_1633 ();
 sg13g2_fill_2 FILLER_17_1640 ();
 sg13g2_fill_1 FILLER_17_1666 ();
 sg13g2_decap_8 FILLER_17_1672 ();
 sg13g2_fill_2 FILLER_17_1679 ();
 sg13g2_fill_1 FILLER_17_1681 ();
 sg13g2_fill_2 FILLER_17_1734 ();
 sg13g2_fill_1 FILLER_17_1792 ();
 sg13g2_fill_1 FILLER_17_1812 ();
 sg13g2_fill_2 FILLER_17_1824 ();
 sg13g2_fill_2 FILLER_17_1835 ();
 sg13g2_fill_1 FILLER_17_1837 ();
 sg13g2_decap_8 FILLER_17_1841 ();
 sg13g2_decap_8 FILLER_17_1848 ();
 sg13g2_decap_4 FILLER_17_1855 ();
 sg13g2_fill_2 FILLER_17_1894 ();
 sg13g2_fill_1 FILLER_17_1927 ();
 sg13g2_decap_4 FILLER_17_1934 ();
 sg13g2_fill_2 FILLER_17_1938 ();
 sg13g2_fill_1 FILLER_17_1945 ();
 sg13g2_fill_1 FILLER_17_1950 ();
 sg13g2_fill_1 FILLER_17_1982 ();
 sg13g2_fill_1 FILLER_17_1988 ();
 sg13g2_fill_2 FILLER_17_2015 ();
 sg13g2_fill_1 FILLER_17_2047 ();
 sg13g2_fill_1 FILLER_17_2053 ();
 sg13g2_fill_1 FILLER_17_2062 ();
 sg13g2_fill_1 FILLER_17_2080 ();
 sg13g2_decap_8 FILLER_17_2124 ();
 sg13g2_fill_1 FILLER_17_2131 ();
 sg13g2_decap_8 FILLER_17_2136 ();
 sg13g2_decap_4 FILLER_17_2143 ();
 sg13g2_fill_2 FILLER_17_2229 ();
 sg13g2_fill_1 FILLER_17_2231 ();
 sg13g2_decap_8 FILLER_17_2254 ();
 sg13g2_decap_8 FILLER_17_2261 ();
 sg13g2_decap_8 FILLER_17_2268 ();
 sg13g2_decap_8 FILLER_17_2275 ();
 sg13g2_decap_8 FILLER_17_2282 ();
 sg13g2_fill_2 FILLER_17_2292 ();
 sg13g2_fill_2 FILLER_17_2302 ();
 sg13g2_fill_1 FILLER_17_2304 ();
 sg13g2_decap_8 FILLER_17_2362 ();
 sg13g2_decap_4 FILLER_17_2369 ();
 sg13g2_fill_2 FILLER_17_2373 ();
 sg13g2_decap_8 FILLER_17_2414 ();
 sg13g2_fill_2 FILLER_17_2421 ();
 sg13g2_decap_4 FILLER_17_2457 ();
 sg13g2_fill_1 FILLER_17_2504 ();
 sg13g2_decap_8 FILLER_17_2510 ();
 sg13g2_decap_8 FILLER_17_2517 ();
 sg13g2_decap_8 FILLER_17_2524 ();
 sg13g2_decap_4 FILLER_17_2531 ();
 sg13g2_fill_2 FILLER_17_2535 ();
 sg13g2_fill_2 FILLER_17_2563 ();
 sg13g2_decap_8 FILLER_17_2574 ();
 sg13g2_decap_8 FILLER_17_2620 ();
 sg13g2_decap_8 FILLER_17_2627 ();
 sg13g2_decap_8 FILLER_17_2634 ();
 sg13g2_decap_8 FILLER_17_2641 ();
 sg13g2_decap_8 FILLER_17_2648 ();
 sg13g2_decap_8 FILLER_17_2655 ();
 sg13g2_decap_8 FILLER_17_2662 ();
 sg13g2_fill_1 FILLER_17_2669 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_48 ();
 sg13g2_decap_8 FILLER_18_53 ();
 sg13g2_decap_8 FILLER_18_60 ();
 sg13g2_decap_8 FILLER_18_67 ();
 sg13g2_decap_8 FILLER_18_74 ();
 sg13g2_decap_4 FILLER_18_81 ();
 sg13g2_fill_2 FILLER_18_123 ();
 sg13g2_fill_1 FILLER_18_125 ();
 sg13g2_decap_4 FILLER_18_139 ();
 sg13g2_fill_1 FILLER_18_143 ();
 sg13g2_decap_8 FILLER_18_159 ();
 sg13g2_decap_4 FILLER_18_166 ();
 sg13g2_decap_8 FILLER_18_180 ();
 sg13g2_decap_8 FILLER_18_187 ();
 sg13g2_fill_2 FILLER_18_194 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_4 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_243 ();
 sg13g2_decap_8 FILLER_18_250 ();
 sg13g2_decap_8 FILLER_18_257 ();
 sg13g2_decap_8 FILLER_18_264 ();
 sg13g2_fill_2 FILLER_18_271 ();
 sg13g2_decap_4 FILLER_18_277 ();
 sg13g2_fill_2 FILLER_18_281 ();
 sg13g2_decap_8 FILLER_18_293 ();
 sg13g2_fill_1 FILLER_18_300 ();
 sg13g2_fill_1 FILLER_18_340 ();
 sg13g2_fill_2 FILLER_18_346 ();
 sg13g2_fill_1 FILLER_18_353 ();
 sg13g2_fill_2 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_decap_4 FILLER_18_382 ();
 sg13g2_decap_4 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_fill_1 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_443 ();
 sg13g2_decap_4 FILLER_18_450 ();
 sg13g2_fill_1 FILLER_18_454 ();
 sg13g2_fill_2 FILLER_18_463 ();
 sg13g2_fill_1 FILLER_18_465 ();
 sg13g2_fill_2 FILLER_18_482 ();
 sg13g2_fill_2 FILLER_18_489 ();
 sg13g2_fill_2 FILLER_18_495 ();
 sg13g2_fill_1 FILLER_18_497 ();
 sg13g2_decap_4 FILLER_18_504 ();
 sg13g2_fill_1 FILLER_18_522 ();
 sg13g2_decap_4 FILLER_18_535 ();
 sg13g2_decap_8 FILLER_18_622 ();
 sg13g2_decap_8 FILLER_18_629 ();
 sg13g2_decap_8 FILLER_18_636 ();
 sg13g2_fill_2 FILLER_18_643 ();
 sg13g2_decap_4 FILLER_18_662 ();
 sg13g2_decap_4 FILLER_18_681 ();
 sg13g2_fill_1 FILLER_18_690 ();
 sg13g2_fill_1 FILLER_18_709 ();
 sg13g2_decap_4 FILLER_18_715 ();
 sg13g2_fill_1 FILLER_18_719 ();
 sg13g2_decap_4 FILLER_18_733 ();
 sg13g2_fill_1 FILLER_18_737 ();
 sg13g2_decap_8 FILLER_18_746 ();
 sg13g2_decap_8 FILLER_18_753 ();
 sg13g2_decap_4 FILLER_18_760 ();
 sg13g2_decap_8 FILLER_18_794 ();
 sg13g2_decap_8 FILLER_18_801 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_fill_2 FILLER_18_815 ();
 sg13g2_fill_2 FILLER_18_851 ();
 sg13g2_fill_1 FILLER_18_853 ();
 sg13g2_fill_2 FILLER_18_931 ();
 sg13g2_fill_1 FILLER_18_933 ();
 sg13g2_decap_8 FILLER_18_964 ();
 sg13g2_fill_2 FILLER_18_971 ();
 sg13g2_decap_8 FILLER_18_1003 ();
 sg13g2_decap_8 FILLER_18_1010 ();
 sg13g2_decap_4 FILLER_18_1017 ();
 sg13g2_fill_2 FILLER_18_1021 ();
 sg13g2_fill_2 FILLER_18_1049 ();
 sg13g2_fill_1 FILLER_18_1051 ();
 sg13g2_decap_8 FILLER_18_1065 ();
 sg13g2_fill_2 FILLER_18_1072 ();
 sg13g2_fill_1 FILLER_18_1105 ();
 sg13g2_decap_4 FILLER_18_1109 ();
 sg13g2_decap_8 FILLER_18_1121 ();
 sg13g2_decap_8 FILLER_18_1128 ();
 sg13g2_decap_8 FILLER_18_1135 ();
 sg13g2_decap_8 FILLER_18_1142 ();
 sg13g2_decap_4 FILLER_18_1149 ();
 sg13g2_fill_2 FILLER_18_1153 ();
 sg13g2_decap_8 FILLER_18_1159 ();
 sg13g2_decap_8 FILLER_18_1166 ();
 sg13g2_decap_4 FILLER_18_1173 ();
 sg13g2_fill_2 FILLER_18_1177 ();
 sg13g2_decap_8 FILLER_18_1183 ();
 sg13g2_decap_8 FILLER_18_1190 ();
 sg13g2_decap_8 FILLER_18_1197 ();
 sg13g2_decap_8 FILLER_18_1204 ();
 sg13g2_decap_8 FILLER_18_1211 ();
 sg13g2_decap_8 FILLER_18_1218 ();
 sg13g2_decap_8 FILLER_18_1225 ();
 sg13g2_decap_8 FILLER_18_1232 ();
 sg13g2_decap_8 FILLER_18_1239 ();
 sg13g2_decap_8 FILLER_18_1246 ();
 sg13g2_decap_8 FILLER_18_1253 ();
 sg13g2_decap_8 FILLER_18_1260 ();
 sg13g2_decap_4 FILLER_18_1267 ();
 sg13g2_fill_1 FILLER_18_1271 ();
 sg13g2_decap_8 FILLER_18_1276 ();
 sg13g2_fill_2 FILLER_18_1283 ();
 sg13g2_decap_8 FILLER_18_1297 ();
 sg13g2_decap_8 FILLER_18_1304 ();
 sg13g2_fill_2 FILLER_18_1311 ();
 sg13g2_fill_1 FILLER_18_1313 ();
 sg13g2_fill_2 FILLER_18_1319 ();
 sg13g2_fill_2 FILLER_18_1326 ();
 sg13g2_fill_1 FILLER_18_1359 ();
 sg13g2_decap_8 FILLER_18_1382 ();
 sg13g2_decap_8 FILLER_18_1389 ();
 sg13g2_decap_8 FILLER_18_1396 ();
 sg13g2_decap_8 FILLER_18_1403 ();
 sg13g2_decap_4 FILLER_18_1410 ();
 sg13g2_fill_2 FILLER_18_1418 ();
 sg13g2_decap_8 FILLER_18_1429 ();
 sg13g2_decap_8 FILLER_18_1436 ();
 sg13g2_fill_2 FILLER_18_1470 ();
 sg13g2_fill_1 FILLER_18_1477 ();
 sg13g2_fill_2 FILLER_18_1521 ();
 sg13g2_decap_4 FILLER_18_1528 ();
 sg13g2_fill_2 FILLER_18_1532 ();
 sg13g2_fill_1 FILLER_18_1549 ();
 sg13g2_decap_4 FILLER_18_1557 ();
 sg13g2_fill_1 FILLER_18_1561 ();
 sg13g2_decap_4 FILLER_18_1571 ();
 sg13g2_fill_2 FILLER_18_1595 ();
 sg13g2_decap_8 FILLER_18_1615 ();
 sg13g2_decap_8 FILLER_18_1622 ();
 sg13g2_fill_1 FILLER_18_1629 ();
 sg13g2_decap_8 FILLER_18_1642 ();
 sg13g2_decap_4 FILLER_18_1649 ();
 sg13g2_fill_1 FILLER_18_1653 ();
 sg13g2_decap_4 FILLER_18_1660 ();
 sg13g2_fill_1 FILLER_18_1664 ();
 sg13g2_decap_8 FILLER_18_1691 ();
 sg13g2_fill_2 FILLER_18_1698 ();
 sg13g2_fill_1 FILLER_18_1700 ();
 sg13g2_decap_8 FILLER_18_1731 ();
 sg13g2_decap_8 FILLER_18_1742 ();
 sg13g2_fill_2 FILLER_18_1749 ();
 sg13g2_fill_1 FILLER_18_1751 ();
 sg13g2_fill_1 FILLER_18_1793 ();
 sg13g2_fill_2 FILLER_18_1853 ();
 sg13g2_decap_8 FILLER_18_1860 ();
 sg13g2_fill_2 FILLER_18_1867 ();
 sg13g2_fill_2 FILLER_18_1878 ();
 sg13g2_decap_8 FILLER_18_1893 ();
 sg13g2_decap_8 FILLER_18_1900 ();
 sg13g2_decap_4 FILLER_18_1907 ();
 sg13g2_decap_4 FILLER_18_1937 ();
 sg13g2_fill_1 FILLER_18_1941 ();
 sg13g2_fill_1 FILLER_18_1994 ();
 sg13g2_decap_4 FILLER_18_2018 ();
 sg13g2_fill_2 FILLER_18_2022 ();
 sg13g2_fill_1 FILLER_18_2033 ();
 sg13g2_fill_1 FILLER_18_2040 ();
 sg13g2_fill_2 FILLER_18_2045 ();
 sg13g2_fill_1 FILLER_18_2047 ();
 sg13g2_fill_2 FILLER_18_2056 ();
 sg13g2_fill_1 FILLER_18_2058 ();
 sg13g2_fill_2 FILLER_18_2068 ();
 sg13g2_fill_1 FILLER_18_2070 ();
 sg13g2_fill_2 FILLER_18_2097 ();
 sg13g2_fill_1 FILLER_18_2099 ();
 sg13g2_decap_4 FILLER_18_2104 ();
 sg13g2_decap_4 FILLER_18_2113 ();
 sg13g2_fill_1 FILLER_18_2117 ();
 sg13g2_fill_1 FILLER_18_2122 ();
 sg13g2_decap_8 FILLER_18_2146 ();
 sg13g2_decap_8 FILLER_18_2153 ();
 sg13g2_fill_1 FILLER_18_2160 ();
 sg13g2_fill_1 FILLER_18_2168 ();
 sg13g2_fill_2 FILLER_18_2183 ();
 sg13g2_fill_2 FILLER_18_2194 ();
 sg13g2_fill_1 FILLER_18_2196 ();
 sg13g2_decap_8 FILLER_18_2201 ();
 sg13g2_decap_8 FILLER_18_2208 ();
 sg13g2_decap_8 FILLER_18_2215 ();
 sg13g2_decap_4 FILLER_18_2222 ();
 sg13g2_decap_8 FILLER_18_2257 ();
 sg13g2_decap_8 FILLER_18_2264 ();
 sg13g2_decap_4 FILLER_18_2271 ();
 sg13g2_fill_2 FILLER_18_2275 ();
 sg13g2_fill_1 FILLER_18_2282 ();
 sg13g2_decap_4 FILLER_18_2317 ();
 sg13g2_decap_8 FILLER_18_2324 ();
 sg13g2_decap_8 FILLER_18_2331 ();
 sg13g2_decap_4 FILLER_18_2338 ();
 sg13g2_fill_1 FILLER_18_2342 ();
 sg13g2_decap_8 FILLER_18_2349 ();
 sg13g2_decap_8 FILLER_18_2356 ();
 sg13g2_fill_1 FILLER_18_2363 ();
 sg13g2_decap_8 FILLER_18_2382 ();
 sg13g2_decap_8 FILLER_18_2389 ();
 sg13g2_decap_8 FILLER_18_2396 ();
 sg13g2_decap_8 FILLER_18_2403 ();
 sg13g2_decap_8 FILLER_18_2410 ();
 sg13g2_decap_8 FILLER_18_2417 ();
 sg13g2_decap_4 FILLER_18_2424 ();
 sg13g2_decap_8 FILLER_18_2433 ();
 sg13g2_fill_2 FILLER_18_2440 ();
 sg13g2_fill_1 FILLER_18_2442 ();
 sg13g2_decap_8 FILLER_18_2461 ();
 sg13g2_decap_8 FILLER_18_2468 ();
 sg13g2_decap_4 FILLER_18_2475 ();
 sg13g2_fill_1 FILLER_18_2479 ();
 sg13g2_decap_8 FILLER_18_2532 ();
 sg13g2_fill_2 FILLER_18_2539 ();
 sg13g2_fill_1 FILLER_18_2541 ();
 sg13g2_decap_8 FILLER_18_2552 ();
 sg13g2_decap_8 FILLER_18_2559 ();
 sg13g2_decap_8 FILLER_18_2566 ();
 sg13g2_decap_4 FILLER_18_2573 ();
 sg13g2_fill_2 FILLER_18_2594 ();
 sg13g2_fill_1 FILLER_18_2596 ();
 sg13g2_decap_8 FILLER_18_2623 ();
 sg13g2_decap_8 FILLER_18_2630 ();
 sg13g2_decap_8 FILLER_18_2637 ();
 sg13g2_decap_8 FILLER_18_2644 ();
 sg13g2_decap_8 FILLER_18_2651 ();
 sg13g2_decap_8 FILLER_18_2658 ();
 sg13g2_decap_4 FILLER_18_2665 ();
 sg13g2_fill_1 FILLER_18_2669 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_4 FILLER_19_21 ();
 sg13g2_fill_2 FILLER_19_25 ();
 sg13g2_decap_4 FILLER_19_37 ();
 sg13g2_fill_1 FILLER_19_41 ();
 sg13g2_fill_2 FILLER_19_48 ();
 sg13g2_fill_1 FILLER_19_50 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_4 FILLER_19_91 ();
 sg13g2_fill_1 FILLER_19_95 ();
 sg13g2_fill_1 FILLER_19_104 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_fill_1 FILLER_19_116 ();
 sg13g2_fill_2 FILLER_19_127 ();
 sg13g2_decap_8 FILLER_19_150 ();
 sg13g2_decap_4 FILLER_19_157 ();
 sg13g2_fill_2 FILLER_19_161 ();
 sg13g2_fill_2 FILLER_19_209 ();
 sg13g2_decap_4 FILLER_19_237 ();
 sg13g2_fill_1 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_297 ();
 sg13g2_decap_8 FILLER_19_304 ();
 sg13g2_fill_2 FILLER_19_311 ();
 sg13g2_fill_2 FILLER_19_333 ();
 sg13g2_fill_1 FILLER_19_335 ();
 sg13g2_decap_4 FILLER_19_362 ();
 sg13g2_fill_1 FILLER_19_366 ();
 sg13g2_decap_4 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_403 ();
 sg13g2_fill_1 FILLER_19_410 ();
 sg13g2_fill_2 FILLER_19_420 ();
 sg13g2_fill_2 FILLER_19_431 ();
 sg13g2_fill_1 FILLER_19_433 ();
 sg13g2_decap_8 FILLER_19_442 ();
 sg13g2_decap_4 FILLER_19_449 ();
 sg13g2_fill_1 FILLER_19_483 ();
 sg13g2_fill_2 FILLER_19_489 ();
 sg13g2_fill_1 FILLER_19_491 ();
 sg13g2_decap_4 FILLER_19_521 ();
 sg13g2_fill_1 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_529 ();
 sg13g2_decap_8 FILLER_19_536 ();
 sg13g2_fill_2 FILLER_19_543 ();
 sg13g2_fill_1 FILLER_19_545 ();
 sg13g2_fill_1 FILLER_19_567 ();
 sg13g2_fill_2 FILLER_19_572 ();
 sg13g2_fill_1 FILLER_19_599 ();
 sg13g2_fill_1 FILLER_19_608 ();
 sg13g2_decap_4 FILLER_19_617 ();
 sg13g2_fill_2 FILLER_19_621 ();
 sg13g2_decap_8 FILLER_19_627 ();
 sg13g2_decap_8 FILLER_19_634 ();
 sg13g2_fill_2 FILLER_19_641 ();
 sg13g2_fill_1 FILLER_19_643 ();
 sg13g2_decap_8 FILLER_19_674 ();
 sg13g2_fill_1 FILLER_19_700 ();
 sg13g2_fill_2 FILLER_19_714 ();
 sg13g2_fill_1 FILLER_19_716 ();
 sg13g2_decap_4 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_751 ();
 sg13g2_fill_2 FILLER_19_758 ();
 sg13g2_decap_8 FILLER_19_808 ();
 sg13g2_decap_4 FILLER_19_815 ();
 sg13g2_fill_2 FILLER_19_819 ();
 sg13g2_fill_2 FILLER_19_851 ();
 sg13g2_fill_1 FILLER_19_853 ();
 sg13g2_decap_8 FILLER_19_901 ();
 sg13g2_fill_2 FILLER_19_908 ();
 sg13g2_fill_1 FILLER_19_910 ();
 sg13g2_decap_4 FILLER_19_919 ();
 sg13g2_fill_1 FILLER_19_923 ();
 sg13g2_decap_8 FILLER_19_936 ();
 sg13g2_decap_4 FILLER_19_943 ();
 sg13g2_fill_2 FILLER_19_947 ();
 sg13g2_fill_1 FILLER_19_953 ();
 sg13g2_decap_8 FILLER_19_984 ();
 sg13g2_fill_1 FILLER_19_991 ();
 sg13g2_decap_4 FILLER_19_997 ();
 sg13g2_fill_2 FILLER_19_1015 ();
 sg13g2_fill_1 FILLER_19_1017 ();
 sg13g2_fill_1 FILLER_19_1035 ();
 sg13g2_decap_4 FILLER_19_1067 ();
 sg13g2_fill_1 FILLER_19_1071 ();
 sg13g2_decap_8 FILLER_19_1078 ();
 sg13g2_fill_2 FILLER_19_1085 ();
 sg13g2_fill_1 FILLER_19_1087 ();
 sg13g2_fill_1 FILLER_19_1096 ();
 sg13g2_decap_4 FILLER_19_1149 ();
 sg13g2_fill_1 FILLER_19_1153 ();
 sg13g2_decap_8 FILLER_19_1159 ();
 sg13g2_decap_8 FILLER_19_1166 ();
 sg13g2_decap_8 FILLER_19_1173 ();
 sg13g2_decap_4 FILLER_19_1180 ();
 sg13g2_fill_2 FILLER_19_1184 ();
 sg13g2_decap_8 FILLER_19_1199 ();
 sg13g2_decap_4 FILLER_19_1206 ();
 sg13g2_fill_2 FILLER_19_1210 ();
 sg13g2_decap_4 FILLER_19_1243 ();
 sg13g2_fill_1 FILLER_19_1247 ();
 sg13g2_decap_8 FILLER_19_1253 ();
 sg13g2_decap_8 FILLER_19_1264 ();
 sg13g2_decap_8 FILLER_19_1271 ();
 sg13g2_decap_8 FILLER_19_1278 ();
 sg13g2_decap_8 FILLER_19_1285 ();
 sg13g2_decap_8 FILLER_19_1292 ();
 sg13g2_decap_8 FILLER_19_1308 ();
 sg13g2_decap_4 FILLER_19_1315 ();
 sg13g2_decap_8 FILLER_19_1323 ();
 sg13g2_decap_4 FILLER_19_1330 ();
 sg13g2_fill_2 FILLER_19_1364 ();
 sg13g2_decap_4 FILLER_19_1371 ();
 sg13g2_fill_2 FILLER_19_1375 ();
 sg13g2_decap_8 FILLER_19_1381 ();
 sg13g2_fill_2 FILLER_19_1388 ();
 sg13g2_decap_8 FILLER_19_1399 ();
 sg13g2_fill_1 FILLER_19_1406 ();
 sg13g2_decap_8 FILLER_19_1433 ();
 sg13g2_decap_4 FILLER_19_1440 ();
 sg13g2_fill_2 FILLER_19_1444 ();
 sg13g2_fill_2 FILLER_19_1462 ();
 sg13g2_fill_1 FILLER_19_1472 ();
 sg13g2_fill_1 FILLER_19_1479 ();
 sg13g2_fill_2 FILLER_19_1512 ();
 sg13g2_fill_1 FILLER_19_1569 ();
 sg13g2_fill_2 FILLER_19_1597 ();
 sg13g2_decap_8 FILLER_19_1656 ();
 sg13g2_decap_8 FILLER_19_1663 ();
 sg13g2_decap_8 FILLER_19_1670 ();
 sg13g2_decap_8 FILLER_19_1677 ();
 sg13g2_decap_8 FILLER_19_1684 ();
 sg13g2_decap_8 FILLER_19_1691 ();
 sg13g2_fill_2 FILLER_19_1698 ();
 sg13g2_decap_8 FILLER_19_1713 ();
 sg13g2_fill_1 FILLER_19_1720 ();
 sg13g2_decap_8 FILLER_19_1725 ();
 sg13g2_decap_8 FILLER_19_1732 ();
 sg13g2_fill_2 FILLER_19_1773 ();
 sg13g2_decap_8 FILLER_19_1788 ();
 sg13g2_decap_8 FILLER_19_1795 ();
 sg13g2_fill_2 FILLER_19_1802 ();
 sg13g2_decap_8 FILLER_19_1847 ();
 sg13g2_decap_8 FILLER_19_1854 ();
 sg13g2_decap_8 FILLER_19_1861 ();
 sg13g2_decap_8 FILLER_19_1868 ();
 sg13g2_fill_1 FILLER_19_1875 ();
 sg13g2_decap_8 FILLER_19_1907 ();
 sg13g2_decap_8 FILLER_19_1914 ();
 sg13g2_fill_2 FILLER_19_1926 ();
 sg13g2_fill_1 FILLER_19_1928 ();
 sg13g2_decap_8 FILLER_19_1933 ();
 sg13g2_fill_1 FILLER_19_1945 ();
 sg13g2_decap_8 FILLER_19_1950 ();
 sg13g2_decap_8 FILLER_19_1957 ();
 sg13g2_decap_8 FILLER_19_1964 ();
 sg13g2_decap_8 FILLER_19_1971 ();
 sg13g2_fill_2 FILLER_19_1978 ();
 sg13g2_fill_1 FILLER_19_1988 ();
 sg13g2_fill_2 FILLER_19_2003 ();
 sg13g2_fill_1 FILLER_19_2005 ();
 sg13g2_decap_8 FILLER_19_2011 ();
 sg13g2_decap_8 FILLER_19_2018 ();
 sg13g2_decap_8 FILLER_19_2025 ();
 sg13g2_decap_4 FILLER_19_2032 ();
 sg13g2_fill_2 FILLER_19_2036 ();
 sg13g2_decap_8 FILLER_19_2042 ();
 sg13g2_decap_8 FILLER_19_2049 ();
 sg13g2_decap_4 FILLER_19_2056 ();
 sg13g2_fill_1 FILLER_19_2060 ();
 sg13g2_decap_8 FILLER_19_2117 ();
 sg13g2_decap_8 FILLER_19_2124 ();
 sg13g2_decap_8 FILLER_19_2131 ();
 sg13g2_decap_4 FILLER_19_2138 ();
 sg13g2_fill_2 FILLER_19_2142 ();
 sg13g2_decap_8 FILLER_19_2179 ();
 sg13g2_decap_4 FILLER_19_2197 ();
 sg13g2_fill_2 FILLER_19_2201 ();
 sg13g2_decap_8 FILLER_19_2209 ();
 sg13g2_decap_8 FILLER_19_2216 ();
 sg13g2_fill_2 FILLER_19_2223 ();
 sg13g2_fill_1 FILLER_19_2225 ();
 sg13g2_fill_1 FILLER_19_2252 ();
 sg13g2_decap_4 FILLER_19_2266 ();
 sg13g2_fill_1 FILLER_19_2270 ();
 sg13g2_decap_8 FILLER_19_2307 ();
 sg13g2_decap_8 FILLER_19_2374 ();
 sg13g2_decap_4 FILLER_19_2381 ();
 sg13g2_fill_1 FILLER_19_2385 ();
 sg13g2_decap_8 FILLER_19_2396 ();
 sg13g2_decap_8 FILLER_19_2403 ();
 sg13g2_decap_8 FILLER_19_2410 ();
 sg13g2_decap_4 FILLER_19_2417 ();
 sg13g2_fill_1 FILLER_19_2460 ();
 sg13g2_decap_8 FILLER_19_2465 ();
 sg13g2_decap_8 FILLER_19_2472 ();
 sg13g2_decap_8 FILLER_19_2479 ();
 sg13g2_decap_8 FILLER_19_2486 ();
 sg13g2_decap_8 FILLER_19_2493 ();
 sg13g2_fill_2 FILLER_19_2500 ();
 sg13g2_decap_8 FILLER_19_2528 ();
 sg13g2_decap_4 FILLER_19_2535 ();
 sg13g2_decap_8 FILLER_19_2609 ();
 sg13g2_decap_8 FILLER_19_2616 ();
 sg13g2_decap_8 FILLER_19_2623 ();
 sg13g2_decap_8 FILLER_19_2630 ();
 sg13g2_decap_8 FILLER_19_2637 ();
 sg13g2_decap_8 FILLER_19_2644 ();
 sg13g2_decap_8 FILLER_19_2651 ();
 sg13g2_decap_8 FILLER_19_2658 ();
 sg13g2_decap_4 FILLER_19_2665 ();
 sg13g2_fill_1 FILLER_19_2669 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_14 ();
 sg13g2_fill_1 FILLER_20_79 ();
 sg13g2_fill_1 FILLER_20_84 ();
 sg13g2_fill_2 FILLER_20_150 ();
 sg13g2_decap_8 FILLER_20_156 ();
 sg13g2_decap_8 FILLER_20_163 ();
 sg13g2_decap_8 FILLER_20_170 ();
 sg13g2_decap_8 FILLER_20_177 ();
 sg13g2_decap_4 FILLER_20_184 ();
 sg13g2_fill_1 FILLER_20_188 ();
 sg13g2_decap_4 FILLER_20_199 ();
 sg13g2_fill_1 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_4 FILLER_20_235 ();
 sg13g2_fill_1 FILLER_20_239 ();
 sg13g2_fill_2 FILLER_20_284 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_decap_8 FILLER_20_292 ();
 sg13g2_decap_8 FILLER_20_299 ();
 sg13g2_decap_8 FILLER_20_306 ();
 sg13g2_decap_8 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_320 ();
 sg13g2_fill_1 FILLER_20_327 ();
 sg13g2_fill_1 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_fill_1 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_425 ();
 sg13g2_decap_8 FILLER_20_432 ();
 sg13g2_fill_2 FILLER_20_439 ();
 sg13g2_fill_1 FILLER_20_441 ();
 sg13g2_fill_2 FILLER_20_468 ();
 sg13g2_fill_1 FILLER_20_484 ();
 sg13g2_decap_4 FILLER_20_489 ();
 sg13g2_fill_2 FILLER_20_493 ();
 sg13g2_fill_1 FILLER_20_522 ();
 sg13g2_fill_2 FILLER_20_555 ();
 sg13g2_fill_1 FILLER_20_580 ();
 sg13g2_fill_2 FILLER_20_587 ();
 sg13g2_decap_4 FILLER_20_605 ();
 sg13g2_decap_8 FILLER_20_614 ();
 sg13g2_decap_8 FILLER_20_621 ();
 sg13g2_decap_8 FILLER_20_628 ();
 sg13g2_fill_2 FILLER_20_635 ();
 sg13g2_fill_1 FILLER_20_645 ();
 sg13g2_fill_2 FILLER_20_673 ();
 sg13g2_fill_1 FILLER_20_675 ();
 sg13g2_fill_1 FILLER_20_686 ();
 sg13g2_fill_2 FILLER_20_707 ();
 sg13g2_fill_1 FILLER_20_709 ();
 sg13g2_decap_8 FILLER_20_715 ();
 sg13g2_decap_8 FILLER_20_722 ();
 sg13g2_decap_8 FILLER_20_729 ();
 sg13g2_decap_4 FILLER_20_736 ();
 sg13g2_decap_8 FILLER_20_753 ();
 sg13g2_decap_8 FILLER_20_760 ();
 sg13g2_fill_2 FILLER_20_767 ();
 sg13g2_fill_1 FILLER_20_769 ();
 sg13g2_fill_1 FILLER_20_778 ();
 sg13g2_fill_1 FILLER_20_784 ();
 sg13g2_fill_1 FILLER_20_793 ();
 sg13g2_fill_2 FILLER_20_840 ();
 sg13g2_fill_2 FILLER_20_848 ();
 sg13g2_fill_1 FILLER_20_850 ();
 sg13g2_decap_8 FILLER_20_861 ();
 sg13g2_decap_4 FILLER_20_868 ();
 sg13g2_fill_1 FILLER_20_872 ();
 sg13g2_decap_4 FILLER_20_877 ();
 sg13g2_fill_2 FILLER_20_897 ();
 sg13g2_decap_4 FILLER_20_909 ();
 sg13g2_decap_8 FILLER_20_939 ();
 sg13g2_decap_8 FILLER_20_946 ();
 sg13g2_decap_8 FILLER_20_962 ();
 sg13g2_decap_4 FILLER_20_969 ();
 sg13g2_fill_1 FILLER_20_973 ();
 sg13g2_decap_8 FILLER_20_980 ();
 sg13g2_decap_8 FILLER_20_987 ();
 sg13g2_decap_8 FILLER_20_994 ();
 sg13g2_fill_1 FILLER_20_1001 ();
 sg13g2_decap_8 FILLER_20_1008 ();
 sg13g2_fill_2 FILLER_20_1015 ();
 sg13g2_fill_1 FILLER_20_1017 ();
 sg13g2_decap_8 FILLER_20_1035 ();
 sg13g2_decap_8 FILLER_20_1042 ();
 sg13g2_decap_4 FILLER_20_1049 ();
 sg13g2_fill_1 FILLER_20_1053 ();
 sg13g2_fill_1 FILLER_20_1064 ();
 sg13g2_fill_1 FILLER_20_1071 ();
 sg13g2_decap_8 FILLER_20_1078 ();
 sg13g2_decap_8 FILLER_20_1085 ();
 sg13g2_fill_2 FILLER_20_1092 ();
 sg13g2_decap_4 FILLER_20_1108 ();
 sg13g2_fill_1 FILLER_20_1120 ();
 sg13g2_fill_1 FILLER_20_1182 ();
 sg13g2_fill_1 FILLER_20_1192 ();
 sg13g2_fill_1 FILLER_20_1199 ();
 sg13g2_fill_2 FILLER_20_1206 ();
 sg13g2_decap_8 FILLER_20_1275 ();
 sg13g2_decap_8 FILLER_20_1282 ();
 sg13g2_decap_4 FILLER_20_1326 ();
 sg13g2_fill_2 FILLER_20_1330 ();
 sg13g2_fill_1 FILLER_20_1337 ();
 sg13g2_fill_2 FILLER_20_1342 ();
 sg13g2_decap_4 FILLER_20_1354 ();
 sg13g2_fill_2 FILLER_20_1384 ();
 sg13g2_fill_2 FILLER_20_1391 ();
 sg13g2_fill_1 FILLER_20_1393 ();
 sg13g2_fill_1 FILLER_20_1402 ();
 sg13g2_fill_2 FILLER_20_1408 ();
 sg13g2_fill_1 FILLER_20_1410 ();
 sg13g2_fill_1 FILLER_20_1419 ();
 sg13g2_fill_1 FILLER_20_1446 ();
 sg13g2_fill_1 FILLER_20_1452 ();
 sg13g2_fill_1 FILLER_20_1479 ();
 sg13g2_fill_2 FILLER_20_1484 ();
 sg13g2_fill_2 FILLER_20_1524 ();
 sg13g2_fill_2 FILLER_20_1539 ();
 sg13g2_fill_2 FILLER_20_1583 ();
 sg13g2_fill_2 FILLER_20_1604 ();
 sg13g2_fill_2 FILLER_20_1620 ();
 sg13g2_fill_1 FILLER_20_1627 ();
 sg13g2_decap_8 FILLER_20_1638 ();
 sg13g2_fill_1 FILLER_20_1645 ();
 sg13g2_fill_1 FILLER_20_1677 ();
 sg13g2_decap_8 FILLER_20_1742 ();
 sg13g2_decap_8 FILLER_20_1749 ();
 sg13g2_decap_8 FILLER_20_1756 ();
 sg13g2_fill_2 FILLER_20_1763 ();
 sg13g2_fill_2 FILLER_20_1771 ();
 sg13g2_decap_8 FILLER_20_1783 ();
 sg13g2_decap_8 FILLER_20_1790 ();
 sg13g2_decap_4 FILLER_20_1797 ();
 sg13g2_fill_1 FILLER_20_1846 ();
 sg13g2_fill_2 FILLER_20_1852 ();
 sg13g2_decap_4 FILLER_20_1859 ();
 sg13g2_fill_1 FILLER_20_1863 ();
 sg13g2_decap_4 FILLER_20_1894 ();
 sg13g2_decap_4 FILLER_20_1902 ();
 sg13g2_decap_8 FILLER_20_1914 ();
 sg13g2_decap_8 FILLER_20_1921 ();
 sg13g2_decap_8 FILLER_20_1928 ();
 sg13g2_decap_8 FILLER_20_1935 ();
 sg13g2_decap_8 FILLER_20_1942 ();
 sg13g2_decap_8 FILLER_20_1949 ();
 sg13g2_decap_8 FILLER_20_1956 ();
 sg13g2_fill_2 FILLER_20_1963 ();
 sg13g2_decap_8 FILLER_20_1978 ();
 sg13g2_decap_4 FILLER_20_1985 ();
 sg13g2_fill_2 FILLER_20_1993 ();
 sg13g2_decap_4 FILLER_20_1999 ();
 sg13g2_fill_1 FILLER_20_2033 ();
 sg13g2_decap_8 FILLER_20_2066 ();
 sg13g2_decap_8 FILLER_20_2077 ();
 sg13g2_fill_2 FILLER_20_2084 ();
 sg13g2_fill_1 FILLER_20_2086 ();
 sg13g2_decap_8 FILLER_20_2099 ();
 sg13g2_fill_1 FILLER_20_2106 ();
 sg13g2_fill_2 FILLER_20_2112 ();
 sg13g2_fill_1 FILLER_20_2114 ();
 sg13g2_decap_4 FILLER_20_2119 ();
 sg13g2_fill_1 FILLER_20_2123 ();
 sg13g2_decap_4 FILLER_20_2137 ();
 sg13g2_fill_2 FILLER_20_2141 ();
 sg13g2_fill_1 FILLER_20_2147 ();
 sg13g2_fill_1 FILLER_20_2152 ();
 sg13g2_fill_2 FILLER_20_2191 ();
 sg13g2_fill_1 FILLER_20_2229 ();
 sg13g2_decap_4 FILLER_20_2235 ();
 sg13g2_fill_2 FILLER_20_2243 ();
 sg13g2_fill_1 FILLER_20_2251 ();
 sg13g2_decap_8 FILLER_20_2265 ();
 sg13g2_decap_8 FILLER_20_2272 ();
 sg13g2_decap_8 FILLER_20_2279 ();
 sg13g2_fill_2 FILLER_20_2286 ();
 sg13g2_fill_1 FILLER_20_2288 ();
 sg13g2_decap_8 FILLER_20_2299 ();
 sg13g2_fill_2 FILLER_20_2306 ();
 sg13g2_decap_8 FILLER_20_2329 ();
 sg13g2_decap_8 FILLER_20_2336 ();
 sg13g2_fill_1 FILLER_20_2343 ();
 sg13g2_decap_4 FILLER_20_2348 ();
 sg13g2_fill_2 FILLER_20_2352 ();
 sg13g2_decap_4 FILLER_20_2358 ();
 sg13g2_fill_2 FILLER_20_2388 ();
 sg13g2_fill_1 FILLER_20_2390 ();
 sg13g2_decap_8 FILLER_20_2417 ();
 sg13g2_decap_8 FILLER_20_2424 ();
 sg13g2_decap_8 FILLER_20_2431 ();
 sg13g2_decap_8 FILLER_20_2438 ();
 sg13g2_decap_8 FILLER_20_2445 ();
 sg13g2_fill_1 FILLER_20_2452 ();
 sg13g2_decap_8 FILLER_20_2484 ();
 sg13g2_fill_1 FILLER_20_2491 ();
 sg13g2_decap_8 FILLER_20_2513 ();
 sg13g2_fill_2 FILLER_20_2520 ();
 sg13g2_fill_1 FILLER_20_2522 ();
 sg13g2_fill_1 FILLER_20_2538 ();
 sg13g2_decap_4 FILLER_20_2565 ();
 sg13g2_fill_1 FILLER_20_2569 ();
 sg13g2_fill_1 FILLER_20_2578 ();
 sg13g2_decap_8 FILLER_20_2588 ();
 sg13g2_decap_8 FILLER_20_2595 ();
 sg13g2_decap_8 FILLER_20_2602 ();
 sg13g2_decap_8 FILLER_20_2609 ();
 sg13g2_decap_8 FILLER_20_2616 ();
 sg13g2_decap_8 FILLER_20_2623 ();
 sg13g2_decap_8 FILLER_20_2630 ();
 sg13g2_decap_8 FILLER_20_2637 ();
 sg13g2_decap_8 FILLER_20_2644 ();
 sg13g2_decap_8 FILLER_20_2651 ();
 sg13g2_decap_8 FILLER_20_2658 ();
 sg13g2_decap_4 FILLER_20_2665 ();
 sg13g2_fill_1 FILLER_20_2669 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_55 ();
 sg13g2_fill_1 FILLER_21_57 ();
 sg13g2_decap_8 FILLER_21_62 ();
 sg13g2_decap_8 FILLER_21_69 ();
 sg13g2_decap_8 FILLER_21_76 ();
 sg13g2_decap_8 FILLER_21_83 ();
 sg13g2_decap_8 FILLER_21_95 ();
 sg13g2_decap_8 FILLER_21_102 ();
 sg13g2_decap_4 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_159 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_decap_8 FILLER_21_177 ();
 sg13g2_fill_1 FILLER_21_184 ();
 sg13g2_decap_8 FILLER_21_195 ();
 sg13g2_decap_8 FILLER_21_202 ();
 sg13g2_decap_8 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_216 ();
 sg13g2_decap_8 FILLER_21_223 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_decap_4 FILLER_21_237 ();
 sg13g2_fill_2 FILLER_21_241 ();
 sg13g2_fill_2 FILLER_21_253 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_decap_8 FILLER_21_261 ();
 sg13g2_decap_4 FILLER_21_268 ();
 sg13g2_fill_1 FILLER_21_272 ();
 sg13g2_decap_4 FILLER_21_283 ();
 sg13g2_fill_2 FILLER_21_297 ();
 sg13g2_fill_1 FILLER_21_299 ();
 sg13g2_decap_8 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_4 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_359 ();
 sg13g2_decap_8 FILLER_21_366 ();
 sg13g2_decap_4 FILLER_21_373 ();
 sg13g2_fill_1 FILLER_21_377 ();
 sg13g2_decap_4 FILLER_21_394 ();
 sg13g2_fill_1 FILLER_21_398 ();
 sg13g2_fill_1 FILLER_21_411 ();
 sg13g2_decap_4 FILLER_21_415 ();
 sg13g2_fill_1 FILLER_21_419 ();
 sg13g2_fill_1 FILLER_21_423 ();
 sg13g2_decap_4 FILLER_21_435 ();
 sg13g2_fill_2 FILLER_21_439 ();
 sg13g2_fill_2 FILLER_21_449 ();
 sg13g2_fill_1 FILLER_21_451 ();
 sg13g2_fill_1 FILLER_21_483 ();
 sg13g2_fill_2 FILLER_21_529 ();
 sg13g2_fill_2 FILLER_21_558 ();
 sg13g2_fill_1 FILLER_21_569 ();
 sg13g2_fill_2 FILLER_21_579 ();
 sg13g2_fill_1 FILLER_21_585 ();
 sg13g2_fill_1 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_622 ();
 sg13g2_decap_8 FILLER_21_629 ();
 sg13g2_fill_2 FILLER_21_636 ();
 sg13g2_fill_1 FILLER_21_649 ();
 sg13g2_fill_2 FILLER_21_665 ();
 sg13g2_fill_2 FILLER_21_674 ();
 sg13g2_fill_1 FILLER_21_676 ();
 sg13g2_decap_4 FILLER_21_682 ();
 sg13g2_fill_1 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_696 ();
 sg13g2_decap_8 FILLER_21_703 ();
 sg13g2_decap_8 FILLER_21_710 ();
 sg13g2_decap_4 FILLER_21_717 ();
 sg13g2_decap_8 FILLER_21_726 ();
 sg13g2_decap_8 FILLER_21_733 ();
 sg13g2_fill_2 FILLER_21_740 ();
 sg13g2_fill_2 FILLER_21_778 ();
 sg13g2_decap_8 FILLER_21_823 ();
 sg13g2_decap_8 FILLER_21_830 ();
 sg13g2_fill_2 FILLER_21_837 ();
 sg13g2_decap_8 FILLER_21_845 ();
 sg13g2_decap_8 FILLER_21_852 ();
 sg13g2_fill_2 FILLER_21_859 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_fill_1 FILLER_21_909 ();
 sg13g2_decap_8 FILLER_21_936 ();
 sg13g2_decap_8 FILLER_21_943 ();
 sg13g2_decap_8 FILLER_21_960 ();
 sg13g2_fill_1 FILLER_21_967 ();
 sg13g2_decap_4 FILLER_21_973 ();
 sg13g2_fill_1 FILLER_21_981 ();
 sg13g2_fill_2 FILLER_21_1008 ();
 sg13g2_decap_4 FILLER_21_1036 ();
 sg13g2_fill_2 FILLER_21_1071 ();
 sg13g2_fill_2 FILLER_21_1077 ();
 sg13g2_fill_1 FILLER_21_1091 ();
 sg13g2_fill_2 FILLER_21_1134 ();
 sg13g2_fill_1 FILLER_21_1144 ();
 sg13g2_decap_4 FILLER_21_1154 ();
 sg13g2_fill_1 FILLER_21_1158 ();
 sg13g2_decap_8 FILLER_21_1246 ();
 sg13g2_fill_2 FILLER_21_1253 ();
 sg13g2_fill_1 FILLER_21_1255 ();
 sg13g2_fill_2 FILLER_21_1260 ();
 sg13g2_fill_1 FILLER_21_1262 ();
 sg13g2_fill_2 FILLER_21_1323 ();
 sg13g2_fill_1 FILLER_21_1325 ();
 sg13g2_fill_2 FILLER_21_1339 ();
 sg13g2_fill_1 FILLER_21_1341 ();
 sg13g2_fill_2 FILLER_21_1372 ();
 sg13g2_fill_1 FILLER_21_1374 ();
 sg13g2_fill_2 FILLER_21_1381 ();
 sg13g2_fill_1 FILLER_21_1383 ();
 sg13g2_fill_2 FILLER_21_1390 ();
 sg13g2_fill_1 FILLER_21_1409 ();
 sg13g2_fill_1 FILLER_21_1415 ();
 sg13g2_fill_1 FILLER_21_1422 ();
 sg13g2_fill_1 FILLER_21_1428 ();
 sg13g2_fill_2 FILLER_21_1434 ();
 sg13g2_fill_1 FILLER_21_1436 ();
 sg13g2_decap_8 FILLER_21_1443 ();
 sg13g2_decap_4 FILLER_21_1450 ();
 sg13g2_fill_1 FILLER_21_1454 ();
 sg13g2_fill_2 FILLER_21_1460 ();
 sg13g2_fill_2 FILLER_21_1468 ();
 sg13g2_fill_2 FILLER_21_1475 ();
 sg13g2_fill_2 FILLER_21_1550 ();
 sg13g2_fill_2 FILLER_21_1575 ();
 sg13g2_fill_2 FILLER_21_1581 ();
 sg13g2_fill_2 FILLER_21_1609 ();
 sg13g2_fill_1 FILLER_21_1611 ();
 sg13g2_fill_2 FILLER_21_1638 ();
 sg13g2_fill_1 FILLER_21_1640 ();
 sg13g2_fill_1 FILLER_21_1645 ();
 sg13g2_fill_1 FILLER_21_1651 ();
 sg13g2_fill_1 FILLER_21_1661 ();
 sg13g2_decap_8 FILLER_21_1666 ();
 sg13g2_decap_8 FILLER_21_1673 ();
 sg13g2_fill_2 FILLER_21_1680 ();
 sg13g2_fill_1 FILLER_21_1682 ();
 sg13g2_decap_4 FILLER_21_1688 ();
 sg13g2_decap_8 FILLER_21_1697 ();
 sg13g2_decap_4 FILLER_21_1712 ();
 sg13g2_fill_1 FILLER_21_1716 ();
 sg13g2_decap_8 FILLER_21_1752 ();
 sg13g2_fill_2 FILLER_21_1759 ();
 sg13g2_fill_1 FILLER_21_1761 ();
 sg13g2_fill_2 FILLER_21_1774 ();
 sg13g2_decap_8 FILLER_21_1784 ();
 sg13g2_fill_2 FILLER_21_1791 ();
 sg13g2_fill_1 FILLER_21_1793 ();
 sg13g2_decap_8 FILLER_21_1798 ();
 sg13g2_decap_4 FILLER_21_1805 ();
 sg13g2_fill_2 FILLER_21_1827 ();
 sg13g2_fill_1 FILLER_21_1829 ();
 sg13g2_decap_4 FILLER_21_1835 ();
 sg13g2_decap_4 FILLER_21_1845 ();
 sg13g2_fill_2 FILLER_21_1849 ();
 sg13g2_fill_1 FILLER_21_1880 ();
 sg13g2_fill_1 FILLER_21_1886 ();
 sg13g2_decap_8 FILLER_21_1894 ();
 sg13g2_fill_2 FILLER_21_1901 ();
 sg13g2_fill_2 FILLER_21_1908 ();
 sg13g2_decap_8 FILLER_21_1914 ();
 sg13g2_decap_4 FILLER_21_1921 ();
 sg13g2_fill_2 FILLER_21_1925 ();
 sg13g2_fill_1 FILLER_21_1957 ();
 sg13g2_fill_1 FILLER_21_1989 ();
 sg13g2_fill_2 FILLER_21_1994 ();
 sg13g2_fill_1 FILLER_21_1996 ();
 sg13g2_fill_2 FILLER_21_2029 ();
 sg13g2_decap_8 FILLER_21_2072 ();
 sg13g2_decap_4 FILLER_21_2079 ();
 sg13g2_fill_1 FILLER_21_2083 ();
 sg13g2_decap_8 FILLER_21_2097 ();
 sg13g2_decap_4 FILLER_21_2104 ();
 sg13g2_fill_1 FILLER_21_2108 ();
 sg13g2_decap_8 FILLER_21_2135 ();
 sg13g2_decap_8 FILLER_21_2142 ();
 sg13g2_decap_8 FILLER_21_2149 ();
 sg13g2_decap_8 FILLER_21_2156 ();
 sg13g2_decap_8 FILLER_21_2163 ();
 sg13g2_decap_8 FILLER_21_2175 ();
 sg13g2_fill_1 FILLER_21_2182 ();
 sg13g2_decap_4 FILLER_21_2188 ();
 sg13g2_fill_1 FILLER_21_2192 ();
 sg13g2_decap_8 FILLER_21_2204 ();
 sg13g2_decap_8 FILLER_21_2211 ();
 sg13g2_fill_2 FILLER_21_2218 ();
 sg13g2_fill_1 FILLER_21_2246 ();
 sg13g2_fill_2 FILLER_21_2294 ();
 sg13g2_fill_2 FILLER_21_2327 ();
 sg13g2_decap_8 FILLER_21_2334 ();
 sg13g2_decap_8 FILLER_21_2341 ();
 sg13g2_fill_2 FILLER_21_2348 ();
 sg13g2_decap_8 FILLER_21_2381 ();
 sg13g2_fill_1 FILLER_21_2388 ();
 sg13g2_fill_1 FILLER_21_2401 ();
 sg13g2_fill_1 FILLER_21_2408 ();
 sg13g2_fill_1 FILLER_21_2413 ();
 sg13g2_fill_1 FILLER_21_2454 ();
 sg13g2_fill_2 FILLER_21_2460 ();
 sg13g2_fill_1 FILLER_21_2462 ();
 sg13g2_decap_8 FILLER_21_2526 ();
 sg13g2_decap_8 FILLER_21_2533 ();
 sg13g2_fill_2 FILLER_21_2540 ();
 sg13g2_fill_1 FILLER_21_2542 ();
 sg13g2_decap_8 FILLER_21_2549 ();
 sg13g2_decap_8 FILLER_21_2556 ();
 sg13g2_decap_4 FILLER_21_2563 ();
 sg13g2_fill_1 FILLER_21_2567 ();
 sg13g2_decap_4 FILLER_21_2572 ();
 sg13g2_fill_2 FILLER_21_2576 ();
 sg13g2_fill_1 FILLER_21_2617 ();
 sg13g2_decap_8 FILLER_21_2622 ();
 sg13g2_decap_8 FILLER_21_2629 ();
 sg13g2_decap_8 FILLER_21_2636 ();
 sg13g2_decap_8 FILLER_21_2643 ();
 sg13g2_decap_8 FILLER_21_2650 ();
 sg13g2_decap_8 FILLER_21_2657 ();
 sg13g2_decap_4 FILLER_21_2664 ();
 sg13g2_fill_2 FILLER_21_2668 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_decap_4 FILLER_22_38 ();
 sg13g2_fill_2 FILLER_22_42 ();
 sg13g2_decap_4 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_66 ();
 sg13g2_decap_8 FILLER_22_73 ();
 sg13g2_decap_8 FILLER_22_80 ();
 sg13g2_fill_1 FILLER_22_87 ();
 sg13g2_decap_8 FILLER_22_101 ();
 sg13g2_decap_8 FILLER_22_108 ();
 sg13g2_decap_4 FILLER_22_115 ();
 sg13g2_decap_8 FILLER_22_155 ();
 sg13g2_fill_1 FILLER_22_162 ();
 sg13g2_decap_8 FILLER_22_194 ();
 sg13g2_fill_2 FILLER_22_201 ();
 sg13g2_decap_8 FILLER_22_239 ();
 sg13g2_fill_2 FILLER_22_246 ();
 sg13g2_fill_1 FILLER_22_258 ();
 sg13g2_fill_1 FILLER_22_273 ();
 sg13g2_fill_1 FILLER_22_279 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_decap_8 FILLER_22_323 ();
 sg13g2_decap_8 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_fill_1 FILLER_22_379 ();
 sg13g2_fill_1 FILLER_22_384 ();
 sg13g2_decap_4 FILLER_22_393 ();
 sg13g2_fill_2 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_438 ();
 sg13g2_decap_4 FILLER_22_444 ();
 sg13g2_fill_2 FILLER_22_448 ();
 sg13g2_fill_1 FILLER_22_458 ();
 sg13g2_fill_2 FILLER_22_464 ();
 sg13g2_fill_2 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_475 ();
 sg13g2_fill_2 FILLER_22_482 ();
 sg13g2_fill_2 FILLER_22_491 ();
 sg13g2_fill_1 FILLER_22_493 ();
 sg13g2_decap_4 FILLER_22_563 ();
 sg13g2_decap_4 FILLER_22_572 ();
 sg13g2_fill_2 FILLER_22_576 ();
 sg13g2_decap_8 FILLER_22_624 ();
 sg13g2_decap_4 FILLER_22_631 ();
 sg13g2_fill_1 FILLER_22_638 ();
 sg13g2_fill_2 FILLER_22_661 ();
 sg13g2_fill_1 FILLER_22_663 ();
 sg13g2_fill_2 FILLER_22_672 ();
 sg13g2_fill_1 FILLER_22_674 ();
 sg13g2_fill_2 FILLER_22_715 ();
 sg13g2_decap_8 FILLER_22_748 ();
 sg13g2_decap_4 FILLER_22_755 ();
 sg13g2_fill_1 FILLER_22_759 ();
 sg13g2_decap_8 FILLER_22_765 ();
 sg13g2_decap_8 FILLER_22_772 ();
 sg13g2_fill_1 FILLER_22_779 ();
 sg13g2_fill_2 FILLER_22_784 ();
 sg13g2_fill_1 FILLER_22_786 ();
 sg13g2_decap_8 FILLER_22_817 ();
 sg13g2_decap_8 FILLER_22_824 ();
 sg13g2_fill_2 FILLER_22_831 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_decap_8 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_22_868 ();
 sg13g2_fill_2 FILLER_22_875 ();
 sg13g2_fill_1 FILLER_22_877 ();
 sg13g2_decap_4 FILLER_22_882 ();
 sg13g2_fill_2 FILLER_22_886 ();
 sg13g2_decap_4 FILLER_22_891 ();
 sg13g2_fill_1 FILLER_22_895 ();
 sg13g2_decap_4 FILLER_22_904 ();
 sg13g2_fill_2 FILLER_22_948 ();
 sg13g2_fill_2 FILLER_22_984 ();
 sg13g2_fill_2 FILLER_22_998 ();
 sg13g2_fill_2 FILLER_22_1003 ();
 sg13g2_fill_2 FILLER_22_1011 ();
 sg13g2_decap_4 FILLER_22_1044 ();
 sg13g2_decap_4 FILLER_22_1057 ();
 sg13g2_fill_1 FILLER_22_1072 ();
 sg13g2_fill_2 FILLER_22_1078 ();
 sg13g2_decap_8 FILLER_22_1084 ();
 sg13g2_fill_2 FILLER_22_1091 ();
 sg13g2_fill_1 FILLER_22_1093 ();
 sg13g2_decap_8 FILLER_22_1103 ();
 sg13g2_fill_1 FILLER_22_1110 ();
 sg13g2_decap_8 FILLER_22_1117 ();
 sg13g2_decap_8 FILLER_22_1124 ();
 sg13g2_fill_1 FILLER_22_1142 ();
 sg13g2_decap_4 FILLER_22_1149 ();
 sg13g2_fill_2 FILLER_22_1158 ();
 sg13g2_decap_4 FILLER_22_1166 ();
 sg13g2_fill_2 FILLER_22_1175 ();
 sg13g2_decap_4 FILLER_22_1182 ();
 sg13g2_fill_2 FILLER_22_1192 ();
 sg13g2_decap_8 FILLER_22_1211 ();
 sg13g2_decap_8 FILLER_22_1218 ();
 sg13g2_decap_4 FILLER_22_1225 ();
 sg13g2_fill_1 FILLER_22_1229 ();
 sg13g2_decap_8 FILLER_22_1286 ();
 sg13g2_fill_2 FILLER_22_1293 ();
 sg13g2_fill_2 FILLER_22_1336 ();
 sg13g2_decap_4 FILLER_22_1364 ();
 sg13g2_fill_1 FILLER_22_1368 ();
 sg13g2_fill_1 FILLER_22_1373 ();
 sg13g2_fill_1 FILLER_22_1380 ();
 sg13g2_fill_1 FILLER_22_1387 ();
 sg13g2_fill_1 FILLER_22_1394 ();
 sg13g2_fill_1 FILLER_22_1400 ();
 sg13g2_fill_2 FILLER_22_1407 ();
 sg13g2_fill_2 FILLER_22_1419 ();
 sg13g2_decap_8 FILLER_22_1468 ();
 sg13g2_decap_4 FILLER_22_1475 ();
 sg13g2_fill_2 FILLER_22_1479 ();
 sg13g2_fill_1 FILLER_22_1539 ();
 sg13g2_fill_1 FILLER_22_1545 ();
 sg13g2_decap_4 FILLER_22_1607 ();
 sg13g2_fill_2 FILLER_22_1642 ();
 sg13g2_fill_1 FILLER_22_1644 ();
 sg13g2_decap_8 FILLER_22_1675 ();
 sg13g2_decap_8 FILLER_22_1713 ();
 sg13g2_fill_2 FILLER_22_1758 ();
 sg13g2_fill_2 FILLER_22_1768 ();
 sg13g2_fill_1 FILLER_22_1770 ();
 sg13g2_decap_4 FILLER_22_1774 ();
 sg13g2_fill_2 FILLER_22_1778 ();
 sg13g2_decap_4 FILLER_22_1790 ();
 sg13g2_fill_2 FILLER_22_1794 ();
 sg13g2_decap_4 FILLER_22_1801 ();
 sg13g2_fill_2 FILLER_22_1836 ();
 sg13g2_fill_2 FILLER_22_1869 ();
 sg13g2_decap_4 FILLER_22_1944 ();
 sg13g2_fill_2 FILLER_22_1948 ();
 sg13g2_fill_1 FILLER_22_1956 ();
 sg13g2_fill_2 FILLER_22_1983 ();
 sg13g2_decap_4 FILLER_22_1990 ();
 sg13g2_fill_1 FILLER_22_1994 ();
 sg13g2_decap_8 FILLER_22_2000 ();
 sg13g2_decap_4 FILLER_22_2007 ();
 sg13g2_decap_8 FILLER_22_2024 ();
 sg13g2_fill_2 FILLER_22_2031 ();
 sg13g2_decap_8 FILLER_22_2037 ();
 sg13g2_decap_4 FILLER_22_2044 ();
 sg13g2_decap_8 FILLER_22_2052 ();
 sg13g2_fill_2 FILLER_22_2071 ();
 sg13g2_fill_2 FILLER_22_2103 ();
 sg13g2_fill_1 FILLER_22_2105 ();
 sg13g2_fill_2 FILLER_22_2112 ();
 sg13g2_fill_1 FILLER_22_2114 ();
 sg13g2_decap_8 FILLER_22_2120 ();
 sg13g2_fill_2 FILLER_22_2144 ();
 sg13g2_fill_1 FILLER_22_2146 ();
 sg13g2_decap_4 FILLER_22_2151 ();
 sg13g2_decap_4 FILLER_22_2161 ();
 sg13g2_fill_2 FILLER_22_2165 ();
 sg13g2_decap_8 FILLER_22_2207 ();
 sg13g2_decap_4 FILLER_22_2214 ();
 sg13g2_fill_1 FILLER_22_2218 ();
 sg13g2_fill_2 FILLER_22_2233 ();
 sg13g2_fill_1 FILLER_22_2235 ();
 sg13g2_fill_1 FILLER_22_2240 ();
 sg13g2_fill_1 FILLER_22_2247 ();
 sg13g2_fill_2 FILLER_22_2258 ();
 sg13g2_fill_1 FILLER_22_2260 ();
 sg13g2_fill_1 FILLER_22_2322 ();
 sg13g2_fill_1 FILLER_22_2349 ();
 sg13g2_decap_8 FILLER_22_2355 ();
 sg13g2_decap_8 FILLER_22_2362 ();
 sg13g2_fill_1 FILLER_22_2369 ();
 sg13g2_decap_8 FILLER_22_2373 ();
 sg13g2_fill_2 FILLER_22_2380 ();
 sg13g2_decap_4 FILLER_22_2388 ();
 sg13g2_fill_1 FILLER_22_2392 ();
 sg13g2_fill_2 FILLER_22_2461 ();
 sg13g2_fill_1 FILLER_22_2469 ();
 sg13g2_fill_1 FILLER_22_2486 ();
 sg13g2_fill_2 FILLER_22_2499 ();
 sg13g2_fill_2 FILLER_22_2536 ();
 sg13g2_decap_8 FILLER_22_2544 ();
 sg13g2_fill_2 FILLER_22_2551 ();
 sg13g2_fill_1 FILLER_22_2553 ();
 sg13g2_fill_1 FILLER_22_2620 ();
 sg13g2_decap_8 FILLER_22_2647 ();
 sg13g2_decap_8 FILLER_22_2654 ();
 sg13g2_decap_8 FILLER_22_2661 ();
 sg13g2_fill_2 FILLER_22_2668 ();
 sg13g2_fill_2 FILLER_23_30 ();
 sg13g2_fill_1 FILLER_23_36 ();
 sg13g2_decap_8 FILLER_23_41 ();
 sg13g2_decap_8 FILLER_23_48 ();
 sg13g2_decap_8 FILLER_23_55 ();
 sg13g2_decap_8 FILLER_23_62 ();
 sg13g2_decap_8 FILLER_23_69 ();
 sg13g2_decap_8 FILLER_23_76 ();
 sg13g2_decap_8 FILLER_23_83 ();
 sg13g2_decap_8 FILLER_23_90 ();
 sg13g2_decap_8 FILLER_23_97 ();
 sg13g2_fill_2 FILLER_23_104 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_decap_8 FILLER_23_137 ();
 sg13g2_fill_1 FILLER_23_180 ();
 sg13g2_fill_2 FILLER_23_188 ();
 sg13g2_fill_2 FILLER_23_195 ();
 sg13g2_decap_8 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_240 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_fill_2 FILLER_23_284 ();
 sg13g2_fill_1 FILLER_23_286 ();
 sg13g2_decap_4 FILLER_23_302 ();
 sg13g2_fill_2 FILLER_23_306 ();
 sg13g2_decap_8 FILLER_23_313 ();
 sg13g2_decap_8 FILLER_23_320 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_fill_1 FILLER_23_368 ();
 sg13g2_decap_4 FILLER_23_375 ();
 sg13g2_fill_1 FILLER_23_389 ();
 sg13g2_fill_1 FILLER_23_414 ();
 sg13g2_decap_8 FILLER_23_419 ();
 sg13g2_fill_1 FILLER_23_440 ();
 sg13g2_decap_8 FILLER_23_451 ();
 sg13g2_fill_2 FILLER_23_458 ();
 sg13g2_fill_1 FILLER_23_460 ();
 sg13g2_decap_8 FILLER_23_465 ();
 sg13g2_fill_2 FILLER_23_472 ();
 sg13g2_fill_1 FILLER_23_474 ();
 sg13g2_decap_8 FILLER_23_480 ();
 sg13g2_decap_8 FILLER_23_487 ();
 sg13g2_decap_8 FILLER_23_494 ();
 sg13g2_decap_8 FILLER_23_501 ();
 sg13g2_fill_2 FILLER_23_508 ();
 sg13g2_fill_1 FILLER_23_510 ();
 sg13g2_decap_8 FILLER_23_515 ();
 sg13g2_fill_2 FILLER_23_522 ();
 sg13g2_fill_1 FILLER_23_524 ();
 sg13g2_fill_2 FILLER_23_556 ();
 sg13g2_fill_1 FILLER_23_558 ();
 sg13g2_decap_4 FILLER_23_593 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_4 FILLER_23_616 ();
 sg13g2_fill_1 FILLER_23_620 ();
 sg13g2_fill_1 FILLER_23_626 ();
 sg13g2_fill_1 FILLER_23_632 ();
 sg13g2_fill_2 FILLER_23_638 ();
 sg13g2_fill_1 FILLER_23_670 ();
 sg13g2_fill_2 FILLER_23_676 ();
 sg13g2_fill_2 FILLER_23_689 ();
 sg13g2_fill_1 FILLER_23_691 ();
 sg13g2_decap_4 FILLER_23_717 ();
 sg13g2_decap_8 FILLER_23_726 ();
 sg13g2_decap_8 FILLER_23_733 ();
 sg13g2_decap_8 FILLER_23_740 ();
 sg13g2_decap_8 FILLER_23_747 ();
 sg13g2_decap_8 FILLER_23_754 ();
 sg13g2_decap_8 FILLER_23_761 ();
 sg13g2_decap_8 FILLER_23_768 ();
 sg13g2_fill_1 FILLER_23_775 ();
 sg13g2_decap_8 FILLER_23_806 ();
 sg13g2_decap_8 FILLER_23_813 ();
 sg13g2_decap_8 FILLER_23_820 ();
 sg13g2_decap_4 FILLER_23_827 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_23_868 ();
 sg13g2_fill_2 FILLER_23_875 ();
 sg13g2_decap_4 FILLER_23_881 ();
 sg13g2_fill_2 FILLER_23_927 ();
 sg13g2_fill_1 FILLER_23_929 ();
 sg13g2_decap_4 FILLER_23_956 ();
 sg13g2_fill_1 FILLER_23_960 ();
 sg13g2_fill_2 FILLER_23_975 ();
 sg13g2_fill_2 FILLER_23_982 ();
 sg13g2_fill_1 FILLER_23_984 ();
 sg13g2_fill_1 FILLER_23_1044 ();
 sg13g2_fill_1 FILLER_23_1085 ();
 sg13g2_fill_1 FILLER_23_1111 ();
 sg13g2_decap_8 FILLER_23_1121 ();
 sg13g2_decap_8 FILLER_23_1128 ();
 sg13g2_fill_1 FILLER_23_1135 ();
 sg13g2_fill_2 FILLER_23_1167 ();
 sg13g2_decap_8 FILLER_23_1182 ();
 sg13g2_decap_4 FILLER_23_1189 ();
 sg13g2_fill_1 FILLER_23_1193 ();
 sg13g2_decap_8 FILLER_23_1199 ();
 sg13g2_decap_8 FILLER_23_1206 ();
 sg13g2_decap_8 FILLER_23_1213 ();
 sg13g2_fill_2 FILLER_23_1220 ();
 sg13g2_decap_8 FILLER_23_1226 ();
 sg13g2_fill_1 FILLER_23_1233 ();
 sg13g2_fill_2 FILLER_23_1239 ();
 sg13g2_fill_1 FILLER_23_1241 ();
 sg13g2_decap_8 FILLER_23_1290 ();
 sg13g2_decap_4 FILLER_23_1297 ();
 sg13g2_decap_4 FILLER_23_1305 ();
 sg13g2_fill_2 FILLER_23_1309 ();
 sg13g2_fill_2 FILLER_23_1317 ();
 sg13g2_fill_1 FILLER_23_1319 ();
 sg13g2_fill_2 FILLER_23_1326 ();
 sg13g2_fill_1 FILLER_23_1328 ();
 sg13g2_fill_1 FILLER_23_1370 ();
 sg13g2_fill_1 FILLER_23_1420 ();
 sg13g2_fill_2 FILLER_23_1431 ();
 sg13g2_fill_1 FILLER_23_1433 ();
 sg13g2_fill_1 FILLER_23_1446 ();
 sg13g2_fill_2 FILLER_23_1505 ();
 sg13g2_fill_1 FILLER_23_1507 ();
 sg13g2_decap_4 FILLER_23_1517 ();
 sg13g2_fill_2 FILLER_23_1521 ();
 sg13g2_fill_1 FILLER_23_1533 ();
 sg13g2_fill_1 FILLER_23_1599 ();
 sg13g2_decap_8 FILLER_23_1604 ();
 sg13g2_fill_1 FILLER_23_1615 ();
 sg13g2_fill_2 FILLER_23_1620 ();
 sg13g2_fill_2 FILLER_23_1627 ();
 sg13g2_fill_1 FILLER_23_1629 ();
 sg13g2_decap_8 FILLER_23_1635 ();
 sg13g2_fill_1 FILLER_23_1642 ();
 sg13g2_decap_8 FILLER_23_1682 ();
 sg13g2_decap_8 FILLER_23_1689 ();
 sg13g2_decap_8 FILLER_23_1700 ();
 sg13g2_decap_8 FILLER_23_1707 ();
 sg13g2_decap_8 FILLER_23_1714 ();
 sg13g2_fill_2 FILLER_23_1721 ();
 sg13g2_fill_1 FILLER_23_1723 ();
 sg13g2_decap_4 FILLER_23_1768 ();
 sg13g2_fill_1 FILLER_23_1807 ();
 sg13g2_decap_4 FILLER_23_1813 ();
 sg13g2_fill_2 FILLER_23_1817 ();
 sg13g2_fill_2 FILLER_23_1823 ();
 sg13g2_fill_2 FILLER_23_1851 ();
 sg13g2_decap_8 FILLER_23_1857 ();
 sg13g2_fill_2 FILLER_23_1864 ();
 sg13g2_decap_8 FILLER_23_1877 ();
 sg13g2_decap_4 FILLER_23_1884 ();
 sg13g2_fill_1 FILLER_23_1888 ();
 sg13g2_decap_8 FILLER_23_1898 ();
 sg13g2_decap_4 FILLER_23_1905 ();
 sg13g2_fill_2 FILLER_23_1909 ();
 sg13g2_fill_2 FILLER_23_1925 ();
 sg13g2_decap_8 FILLER_23_1962 ();
 sg13g2_decap_4 FILLER_23_1969 ();
 sg13g2_fill_1 FILLER_23_1973 ();
 sg13g2_decap_4 FILLER_23_1990 ();
 sg13g2_fill_1 FILLER_23_1994 ();
 sg13g2_fill_2 FILLER_23_2027 ();
 sg13g2_fill_1 FILLER_23_2029 ();
 sg13g2_decap_8 FILLER_23_2034 ();
 sg13g2_decap_8 FILLER_23_2041 ();
 sg13g2_fill_2 FILLER_23_2048 ();
 sg13g2_fill_1 FILLER_23_2055 ();
 sg13g2_fill_1 FILLER_23_2164 ();
 sg13g2_fill_2 FILLER_23_2191 ();
 sg13g2_fill_2 FILLER_23_2199 ();
 sg13g2_fill_1 FILLER_23_2201 ();
 sg13g2_fill_2 FILLER_23_2207 ();
 sg13g2_fill_2 FILLER_23_2214 ();
 sg13g2_fill_1 FILLER_23_2216 ();
 sg13g2_decap_8 FILLER_23_2230 ();
 sg13g2_decap_4 FILLER_23_2237 ();
 sg13g2_fill_1 FILLER_23_2241 ();
 sg13g2_fill_2 FILLER_23_2248 ();
 sg13g2_fill_2 FILLER_23_2275 ();
 sg13g2_fill_1 FILLER_23_2417 ();
 sg13g2_fill_1 FILLER_23_2424 ();
 sg13g2_fill_1 FILLER_23_2440 ();
 sg13g2_fill_1 FILLER_23_2448 ();
 sg13g2_decap_8 FILLER_23_2514 ();
 sg13g2_fill_1 FILLER_23_2521 ();
 sg13g2_decap_8 FILLER_23_2597 ();
 sg13g2_decap_8 FILLER_23_2604 ();
 sg13g2_decap_8 FILLER_23_2611 ();
 sg13g2_decap_8 FILLER_23_2618 ();
 sg13g2_fill_2 FILLER_23_2625 ();
 sg13g2_fill_1 FILLER_23_2627 ();
 sg13g2_decap_8 FILLER_23_2632 ();
 sg13g2_decap_8 FILLER_23_2639 ();
 sg13g2_decap_8 FILLER_23_2646 ();
 sg13g2_decap_8 FILLER_23_2653 ();
 sg13g2_decap_8 FILLER_23_2660 ();
 sg13g2_fill_2 FILLER_23_2667 ();
 sg13g2_fill_1 FILLER_23_2669 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_4 FILLER_24_35 ();
 sg13g2_fill_1 FILLER_24_39 ();
 sg13g2_fill_2 FILLER_24_66 ();
 sg13g2_decap_4 FILLER_24_106 ();
 sg13g2_decap_8 FILLER_24_115 ();
 sg13g2_fill_2 FILLER_24_122 ();
 sg13g2_fill_1 FILLER_24_124 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_4 FILLER_24_161 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_177 ();
 sg13g2_fill_1 FILLER_24_209 ();
 sg13g2_decap_8 FILLER_24_230 ();
 sg13g2_fill_2 FILLER_24_237 ();
 sg13g2_fill_1 FILLER_24_239 ();
 sg13g2_decap_8 FILLER_24_279 ();
 sg13g2_fill_2 FILLER_24_286 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_fill_1 FILLER_24_299 ();
 sg13g2_fill_1 FILLER_24_307 ();
 sg13g2_decap_8 FILLER_24_313 ();
 sg13g2_fill_2 FILLER_24_320 ();
 sg13g2_decap_8 FILLER_24_358 ();
 sg13g2_decap_8 FILLER_24_365 ();
 sg13g2_fill_1 FILLER_24_411 ();
 sg13g2_fill_2 FILLER_24_415 ();
 sg13g2_fill_2 FILLER_24_443 ();
 sg13g2_fill_2 FILLER_24_451 ();
 sg13g2_fill_1 FILLER_24_453 ();
 sg13g2_decap_8 FILLER_24_467 ();
 sg13g2_fill_1 FILLER_24_474 ();
 sg13g2_decap_8 FILLER_24_488 ();
 sg13g2_fill_2 FILLER_24_495 ();
 sg13g2_fill_2 FILLER_24_501 ();
 sg13g2_fill_1 FILLER_24_503 ();
 sg13g2_decap_4 FILLER_24_515 ();
 sg13g2_fill_1 FILLER_24_550 ();
 sg13g2_fill_1 FILLER_24_563 ();
 sg13g2_fill_2 FILLER_24_569 ();
 sg13g2_fill_1 FILLER_24_579 ();
 sg13g2_decap_4 FILLER_24_592 ();
 sg13g2_decap_8 FILLER_24_606 ();
 sg13g2_fill_2 FILLER_24_613 ();
 sg13g2_decap_4 FILLER_24_627 ();
 sg13g2_fill_2 FILLER_24_667 ();
 sg13g2_fill_2 FILLER_24_673 ();
 sg13g2_fill_1 FILLER_24_675 ();
 sg13g2_fill_1 FILLER_24_690 ();
 sg13g2_fill_2 FILLER_24_716 ();
 sg13g2_decap_8 FILLER_24_722 ();
 sg13g2_decap_8 FILLER_24_755 ();
 sg13g2_decap_8 FILLER_24_762 ();
 sg13g2_decap_8 FILLER_24_769 ();
 sg13g2_fill_1 FILLER_24_776 ();
 sg13g2_decap_8 FILLER_24_811 ();
 sg13g2_fill_1 FILLER_24_818 ();
 sg13g2_decap_4 FILLER_24_897 ();
 sg13g2_fill_1 FILLER_24_909 ();
 sg13g2_fill_1 FILLER_24_923 ();
 sg13g2_decap_8 FILLER_24_929 ();
 sg13g2_fill_1 FILLER_24_936 ();
 sg13g2_decap_8 FILLER_24_941 ();
 sg13g2_decap_8 FILLER_24_948 ();
 sg13g2_decap_4 FILLER_24_955 ();
 sg13g2_fill_2 FILLER_24_959 ();
 sg13g2_decap_8 FILLER_24_966 ();
 sg13g2_decap_8 FILLER_24_973 ();
 sg13g2_decap_4 FILLER_24_980 ();
 sg13g2_fill_1 FILLER_24_1031 ();
 sg13g2_decap_8 FILLER_24_1042 ();
 sg13g2_fill_2 FILLER_24_1049 ();
 sg13g2_fill_2 FILLER_24_1059 ();
 sg13g2_decap_8 FILLER_24_1091 ();
 sg13g2_decap_8 FILLER_24_1103 ();
 sg13g2_fill_1 FILLER_24_1110 ();
 sg13g2_decap_8 FILLER_24_1137 ();
 sg13g2_decap_8 FILLER_24_1148 ();
 sg13g2_decap_8 FILLER_24_1186 ();
 sg13g2_fill_1 FILLER_24_1193 ();
 sg13g2_decap_8 FILLER_24_1200 ();
 sg13g2_decap_8 FILLER_24_1207 ();
 sg13g2_decap_8 FILLER_24_1214 ();
 sg13g2_decap_8 FILLER_24_1221 ();
 sg13g2_fill_2 FILLER_24_1228 ();
 sg13g2_fill_1 FILLER_24_1230 ();
 sg13g2_fill_1 FILLER_24_1235 ();
 sg13g2_fill_1 FILLER_24_1254 ();
 sg13g2_decap_8 FILLER_24_1290 ();
 sg13g2_decap_8 FILLER_24_1297 ();
 sg13g2_decap_8 FILLER_24_1304 ();
 sg13g2_decap_8 FILLER_24_1311 ();
 sg13g2_decap_8 FILLER_24_1318 ();
 sg13g2_decap_8 FILLER_24_1325 ();
 sg13g2_decap_8 FILLER_24_1332 ();
 sg13g2_decap_8 FILLER_24_1339 ();
 sg13g2_decap_8 FILLER_24_1346 ();
 sg13g2_decap_8 FILLER_24_1353 ();
 sg13g2_decap_4 FILLER_24_1360 ();
 sg13g2_fill_1 FILLER_24_1364 ();
 sg13g2_decap_4 FILLER_24_1370 ();
 sg13g2_fill_1 FILLER_24_1379 ();
 sg13g2_decap_4 FILLER_24_1390 ();
 sg13g2_fill_2 FILLER_24_1394 ();
 sg13g2_decap_4 FILLER_24_1409 ();
 sg13g2_decap_4 FILLER_24_1483 ();
 sg13g2_fill_2 FILLER_24_1487 ();
 sg13g2_decap_8 FILLER_24_1520 ();
 sg13g2_decap_8 FILLER_24_1527 ();
 sg13g2_fill_2 FILLER_24_1534 ();
 sg13g2_fill_2 FILLER_24_1544 ();
 sg13g2_fill_1 FILLER_24_1546 ();
 sg13g2_fill_2 FILLER_24_1562 ();
 sg13g2_fill_1 FILLER_24_1564 ();
 sg13g2_decap_8 FILLER_24_1617 ();
 sg13g2_decap_8 FILLER_24_1624 ();
 sg13g2_decap_8 FILLER_24_1631 ();
 sg13g2_decap_8 FILLER_24_1638 ();
 sg13g2_fill_2 FILLER_24_1645 ();
 sg13g2_fill_1 FILLER_24_1647 ();
 sg13g2_decap_4 FILLER_24_1652 ();
 sg13g2_fill_1 FILLER_24_1656 ();
 sg13g2_decap_4 FILLER_24_1683 ();
 sg13g2_fill_2 FILLER_24_1687 ();
 sg13g2_fill_2 FILLER_24_1693 ();
 sg13g2_fill_2 FILLER_24_1708 ();
 sg13g2_fill_1 FILLER_24_1710 ();
 sg13g2_decap_4 FILLER_24_1720 ();
 sg13g2_decap_4 FILLER_24_1730 ();
 sg13g2_fill_2 FILLER_24_1734 ();
 sg13g2_decap_8 FILLER_24_1745 ();
 sg13g2_decap_8 FILLER_24_1752 ();
 sg13g2_decap_8 FILLER_24_1759 ();
 sg13g2_decap_4 FILLER_24_1792 ();
 sg13g2_fill_2 FILLER_24_1796 ();
 sg13g2_decap_4 FILLER_24_1813 ();
 sg13g2_fill_2 FILLER_24_1829 ();
 sg13g2_decap_4 FILLER_24_1836 ();
 sg13g2_fill_1 FILLER_24_1840 ();
 sg13g2_decap_8 FILLER_24_1845 ();
 sg13g2_decap_4 FILLER_24_1852 ();
 sg13g2_fill_1 FILLER_24_1856 ();
 sg13g2_decap_8 FILLER_24_1862 ();
 sg13g2_fill_1 FILLER_24_1869 ();
 sg13g2_decap_8 FILLER_24_1906 ();
 sg13g2_decap_4 FILLER_24_1922 ();
 sg13g2_fill_1 FILLER_24_1926 ();
 sg13g2_fill_2 FILLER_24_1957 ();
 sg13g2_fill_1 FILLER_24_1959 ();
 sg13g2_decap_8 FILLER_24_1966 ();
 sg13g2_decap_8 FILLER_24_1973 ();
 sg13g2_fill_2 FILLER_24_1980 ();
 sg13g2_fill_1 FILLER_24_1982 ();
 sg13g2_decap_8 FILLER_24_2018 ();
 sg13g2_fill_2 FILLER_24_2025 ();
 sg13g2_decap_8 FILLER_24_2031 ();
 sg13g2_decap_8 FILLER_24_2038 ();
 sg13g2_decap_8 FILLER_24_2045 ();
 sg13g2_decap_4 FILLER_24_2110 ();
 sg13g2_fill_2 FILLER_24_2114 ();
 sg13g2_decap_4 FILLER_24_2120 ();
 sg13g2_fill_2 FILLER_24_2132 ();
 sg13g2_decap_8 FILLER_24_2234 ();
 sg13g2_fill_1 FILLER_24_2241 ();
 sg13g2_fill_2 FILLER_24_2246 ();
 sg13g2_decap_8 FILLER_24_2279 ();
 sg13g2_fill_1 FILLER_24_2286 ();
 sg13g2_fill_1 FILLER_24_2292 ();
 sg13g2_fill_1 FILLER_24_2311 ();
 sg13g2_fill_1 FILLER_24_2354 ();
 sg13g2_decap_8 FILLER_24_2361 ();
 sg13g2_fill_2 FILLER_24_2384 ();
 sg13g2_fill_2 FILLER_24_2390 ();
 sg13g2_fill_1 FILLER_24_2392 ();
 sg13g2_decap_8 FILLER_24_2406 ();
 sg13g2_fill_2 FILLER_24_2423 ();
 sg13g2_fill_2 FILLER_24_2435 ();
 sg13g2_fill_1 FILLER_24_2437 ();
 sg13g2_fill_2 FILLER_24_2447 ();
 sg13g2_fill_1 FILLER_24_2463 ();
 sg13g2_decap_8 FILLER_24_2490 ();
 sg13g2_decap_4 FILLER_24_2497 ();
 sg13g2_decap_8 FILLER_24_2531 ();
 sg13g2_decap_8 FILLER_24_2538 ();
 sg13g2_fill_2 FILLER_24_2545 ();
 sg13g2_decap_8 FILLER_24_2556 ();
 sg13g2_decap_8 FILLER_24_2563 ();
 sg13g2_decap_8 FILLER_24_2570 ();
 sg13g2_fill_2 FILLER_24_2577 ();
 sg13g2_decap_8 FILLER_24_2605 ();
 sg13g2_decap_8 FILLER_24_2612 ();
 sg13g2_decap_8 FILLER_24_2619 ();
 sg13g2_decap_8 FILLER_24_2626 ();
 sg13g2_decap_8 FILLER_24_2633 ();
 sg13g2_decap_8 FILLER_24_2640 ();
 sg13g2_decap_8 FILLER_24_2647 ();
 sg13g2_decap_8 FILLER_24_2654 ();
 sg13g2_decap_8 FILLER_24_2661 ();
 sg13g2_fill_2 FILLER_24_2668 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_4 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_100 ();
 sg13g2_decap_8 FILLER_25_111 ();
 sg13g2_decap_8 FILLER_25_118 ();
 sg13g2_decap_4 FILLER_25_125 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_decap_8 FILLER_25_156 ();
 sg13g2_fill_1 FILLER_25_163 ();
 sg13g2_fill_1 FILLER_25_195 ();
 sg13g2_fill_1 FILLER_25_206 ();
 sg13g2_fill_2 FILLER_25_211 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_decap_4 FILLER_25_251 ();
 sg13g2_fill_2 FILLER_25_255 ();
 sg13g2_decap_4 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_fill_1 FILLER_25_285 ();
 sg13g2_fill_1 FILLER_25_293 ();
 sg13g2_decap_4 FILLER_25_320 ();
 sg13g2_fill_2 FILLER_25_324 ();
 sg13g2_fill_2 FILLER_25_333 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_decap_4 FILLER_25_368 ();
 sg13g2_fill_2 FILLER_25_372 ();
 sg13g2_fill_2 FILLER_25_397 ();
 sg13g2_decap_8 FILLER_25_409 ();
 sg13g2_fill_1 FILLER_25_416 ();
 sg13g2_decap_8 FILLER_25_422 ();
 sg13g2_decap_4 FILLER_25_492 ();
 sg13g2_fill_2 FILLER_25_496 ();
 sg13g2_decap_4 FILLER_25_502 ();
 sg13g2_fill_1 FILLER_25_506 ();
 sg13g2_decap_8 FILLER_25_533 ();
 sg13g2_decap_4 FILLER_25_540 ();
 sg13g2_decap_4 FILLER_25_614 ();
 sg13g2_fill_2 FILLER_25_634 ();
 sg13g2_fill_1 FILLER_25_636 ();
 sg13g2_fill_1 FILLER_25_650 ();
 sg13g2_fill_2 FILLER_25_661 ();
 sg13g2_decap_4 FILLER_25_668 ();
 sg13g2_fill_1 FILLER_25_681 ();
 sg13g2_fill_2 FILLER_25_687 ();
 sg13g2_fill_1 FILLER_25_689 ();
 sg13g2_fill_2 FILLER_25_699 ();
 sg13g2_fill_2 FILLER_25_706 ();
 sg13g2_fill_2 FILLER_25_718 ();
 sg13g2_fill_1 FILLER_25_720 ();
 sg13g2_fill_2 FILLER_25_731 ();
 sg13g2_fill_1 FILLER_25_733 ();
 sg13g2_fill_2 FILLER_25_738 ();
 sg13g2_fill_1 FILLER_25_740 ();
 sg13g2_fill_2 FILLER_25_746 ();
 sg13g2_decap_8 FILLER_25_774 ();
 sg13g2_decap_4 FILLER_25_781 ();
 sg13g2_fill_2 FILLER_25_785 ();
 sg13g2_decap_4 FILLER_25_795 ();
 sg13g2_fill_2 FILLER_25_799 ();
 sg13g2_decap_8 FILLER_25_811 ();
 sg13g2_fill_2 FILLER_25_818 ();
 sg13g2_fill_1 FILLER_25_820 ();
 sg13g2_fill_1 FILLER_25_825 ();
 sg13g2_fill_2 FILLER_25_830 ();
 sg13g2_decap_8 FILLER_25_858 ();
 sg13g2_decap_4 FILLER_25_865 ();
 sg13g2_decap_4 FILLER_25_873 ();
 sg13g2_fill_2 FILLER_25_877 ();
 sg13g2_decap_8 FILLER_25_883 ();
 sg13g2_fill_2 FILLER_25_890 ();
 sg13g2_fill_1 FILLER_25_892 ();
 sg13g2_fill_2 FILLER_25_898 ();
 sg13g2_decap_4 FILLER_25_934 ();
 sg13g2_decap_8 FILLER_25_947 ();
 sg13g2_decap_4 FILLER_25_954 ();
 sg13g2_fill_1 FILLER_25_958 ();
 sg13g2_fill_1 FILLER_25_963 ();
 sg13g2_decap_4 FILLER_25_970 ();
 sg13g2_fill_1 FILLER_25_1026 ();
 sg13g2_decap_8 FILLER_25_1053 ();
 sg13g2_fill_2 FILLER_25_1060 ();
 sg13g2_fill_1 FILLER_25_1062 ();
 sg13g2_decap_8 FILLER_25_1089 ();
 sg13g2_decap_8 FILLER_25_1096 ();
 sg13g2_fill_2 FILLER_25_1108 ();
 sg13g2_decap_8 FILLER_25_1114 ();
 sg13g2_decap_8 FILLER_25_1121 ();
 sg13g2_decap_8 FILLER_25_1128 ();
 sg13g2_decap_8 FILLER_25_1135 ();
 sg13g2_decap_8 FILLER_25_1142 ();
 sg13g2_decap_4 FILLER_25_1149 ();
 sg13g2_fill_2 FILLER_25_1153 ();
 sg13g2_decap_4 FILLER_25_1211 ();
 sg13g2_fill_1 FILLER_25_1241 ();
 sg13g2_fill_2 FILLER_25_1251 ();
 sg13g2_fill_2 FILLER_25_1274 ();
 sg13g2_fill_2 FILLER_25_1296 ();
 sg13g2_fill_1 FILLER_25_1298 ();
 sg13g2_decap_8 FILLER_25_1308 ();
 sg13g2_decap_8 FILLER_25_1315 ();
 sg13g2_decap_8 FILLER_25_1322 ();
 sg13g2_fill_1 FILLER_25_1329 ();
 sg13g2_decap_4 FILLER_25_1334 ();
 sg13g2_fill_1 FILLER_25_1338 ();
 sg13g2_fill_1 FILLER_25_1343 ();
 sg13g2_decap_8 FILLER_25_1352 ();
 sg13g2_decap_4 FILLER_25_1359 ();
 sg13g2_decap_8 FILLER_25_1368 ();
 sg13g2_fill_2 FILLER_25_1375 ();
 sg13g2_fill_1 FILLER_25_1377 ();
 sg13g2_fill_2 FILLER_25_1382 ();
 sg13g2_fill_2 FILLER_25_1414 ();
 sg13g2_decap_8 FILLER_25_1421 ();
 sg13g2_fill_1 FILLER_25_1432 ();
 sg13g2_decap_4 FILLER_25_1475 ();
 sg13g2_decap_8 FILLER_25_1523 ();
 sg13g2_fill_1 FILLER_25_1530 ();
 sg13g2_decap_4 FILLER_25_1561 ();
 sg13g2_fill_2 FILLER_25_1565 ();
 sg13g2_decap_8 FILLER_25_1573 ();
 sg13g2_fill_2 FILLER_25_1580 ();
 sg13g2_decap_4 FILLER_25_1595 ();
 sg13g2_decap_8 FILLER_25_1603 ();
 sg13g2_decap_8 FILLER_25_1610 ();
 sg13g2_fill_2 FILLER_25_1617 ();
 sg13g2_decap_8 FILLER_25_1628 ();
 sg13g2_decap_8 FILLER_25_1635 ();
 sg13g2_decap_8 FILLER_25_1642 ();
 sg13g2_decap_8 FILLER_25_1649 ();
 sg13g2_fill_2 FILLER_25_1656 ();
 sg13g2_fill_1 FILLER_25_1658 ();
 sg13g2_decap_8 FILLER_25_1664 ();
 sg13g2_decap_8 FILLER_25_1671 ();
 sg13g2_decap_8 FILLER_25_1678 ();
 sg13g2_decap_4 FILLER_25_1685 ();
 sg13g2_decap_8 FILLER_25_1738 ();
 sg13g2_decap_8 FILLER_25_1745 ();
 sg13g2_fill_2 FILLER_25_1752 ();
 sg13g2_fill_1 FILLER_25_1754 ();
 sg13g2_decap_8 FILLER_25_1759 ();
 sg13g2_decap_8 FILLER_25_1766 ();
 sg13g2_decap_4 FILLER_25_1773 ();
 sg13g2_fill_1 FILLER_25_1782 ();
 sg13g2_fill_2 FILLER_25_1796 ();
 sg13g2_decap_8 FILLER_25_1808 ();
 sg13g2_fill_1 FILLER_25_1820 ();
 sg13g2_fill_1 FILLER_25_1829 ();
 sg13g2_decap_8 FILLER_25_1836 ();
 sg13g2_decap_4 FILLER_25_1843 ();
 sg13g2_fill_2 FILLER_25_1847 ();
 sg13g2_fill_2 FILLER_25_1870 ();
 sg13g2_fill_1 FILLER_25_1898 ();
 sg13g2_decap_8 FILLER_25_1942 ();
 sg13g2_fill_1 FILLER_25_1949 ();
 sg13g2_decap_4 FILLER_25_1955 ();
 sg13g2_fill_2 FILLER_25_1959 ();
 sg13g2_decap_4 FILLER_25_2035 ();
 sg13g2_fill_2 FILLER_25_2039 ();
 sg13g2_decap_4 FILLER_25_2077 ();
 sg13g2_fill_1 FILLER_25_2081 ();
 sg13g2_decap_4 FILLER_25_2086 ();
 sg13g2_fill_1 FILLER_25_2090 ();
 sg13g2_fill_1 FILLER_25_2095 ();
 sg13g2_decap_4 FILLER_25_2122 ();
 sg13g2_fill_1 FILLER_25_2126 ();
 sg13g2_decap_8 FILLER_25_2132 ();
 sg13g2_decap_8 FILLER_25_2139 ();
 sg13g2_fill_1 FILLER_25_2146 ();
 sg13g2_decap_8 FILLER_25_2151 ();
 sg13g2_decap_8 FILLER_25_2158 ();
 sg13g2_decap_8 FILLER_25_2165 ();
 sg13g2_decap_8 FILLER_25_2172 ();
 sg13g2_decap_4 FILLER_25_2188 ();
 sg13g2_fill_2 FILLER_25_2192 ();
 sg13g2_fill_1 FILLER_25_2199 ();
 sg13g2_fill_1 FILLER_25_2226 ();
 sg13g2_fill_1 FILLER_25_2233 ();
 sg13g2_fill_1 FILLER_25_2295 ();
 sg13g2_decap_8 FILLER_25_2305 ();
 sg13g2_fill_2 FILLER_25_2312 ();
 sg13g2_fill_1 FILLER_25_2314 ();
 sg13g2_fill_1 FILLER_25_2357 ();
 sg13g2_fill_2 FILLER_25_2366 ();
 sg13g2_decap_8 FILLER_25_2374 ();
 sg13g2_fill_2 FILLER_25_2385 ();
 sg13g2_fill_1 FILLER_25_2422 ();
 sg13g2_decap_4 FILLER_25_2455 ();
 sg13g2_decap_4 FILLER_25_2464 ();
 sg13g2_fill_2 FILLER_25_2468 ();
 sg13g2_fill_1 FILLER_25_2475 ();
 sg13g2_decap_4 FILLER_25_2507 ();
 sg13g2_decap_8 FILLER_25_2572 ();
 sg13g2_fill_1 FILLER_25_2579 ();
 sg13g2_fill_2 FILLER_25_2584 ();
 sg13g2_fill_2 FILLER_25_2591 ();
 sg13g2_fill_2 FILLER_25_2619 ();
 sg13g2_fill_1 FILLER_25_2621 ();
 sg13g2_decap_8 FILLER_25_2626 ();
 sg13g2_decap_8 FILLER_25_2633 ();
 sg13g2_decap_8 FILLER_25_2640 ();
 sg13g2_decap_8 FILLER_25_2647 ();
 sg13g2_decap_8 FILLER_25_2654 ();
 sg13g2_decap_8 FILLER_25_2661 ();
 sg13g2_fill_2 FILLER_25_2668 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_32 ();
 sg13g2_decap_4 FILLER_26_80 ();
 sg13g2_fill_2 FILLER_26_124 ();
 sg13g2_decap_8 FILLER_26_131 ();
 sg13g2_decap_8 FILLER_26_138 ();
 sg13g2_decap_8 FILLER_26_145 ();
 sg13g2_decap_8 FILLER_26_152 ();
 sg13g2_decap_8 FILLER_26_159 ();
 sg13g2_fill_2 FILLER_26_166 ();
 sg13g2_decap_8 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_183 ();
 sg13g2_fill_1 FILLER_26_185 ();
 sg13g2_fill_2 FILLER_26_190 ();
 sg13g2_fill_1 FILLER_26_192 ();
 sg13g2_decap_4 FILLER_26_222 ();
 sg13g2_fill_1 FILLER_26_226 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_4 FILLER_26_245 ();
 sg13g2_fill_2 FILLER_26_249 ();
 sg13g2_decap_4 FILLER_26_269 ();
 sg13g2_fill_2 FILLER_26_309 ();
 sg13g2_decap_4 FILLER_26_315 ();
 sg13g2_fill_2 FILLER_26_328 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_decap_4 FILLER_26_336 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_fill_2 FILLER_26_351 ();
 sg13g2_fill_2 FILLER_26_358 ();
 sg13g2_fill_1 FILLER_26_360 ();
 sg13g2_fill_1 FILLER_26_366 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_4 FILLER_26_378 ();
 sg13g2_fill_2 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_8 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_26_410 ();
 sg13g2_decap_8 FILLER_26_417 ();
 sg13g2_decap_8 FILLER_26_424 ();
 sg13g2_decap_8 FILLER_26_431 ();
 sg13g2_fill_1 FILLER_26_438 ();
 sg13g2_fill_2 FILLER_26_444 ();
 sg13g2_decap_4 FILLER_26_450 ();
 sg13g2_decap_8 FILLER_26_459 ();
 sg13g2_fill_1 FILLER_26_466 ();
 sg13g2_fill_1 FILLER_26_472 ();
 sg13g2_fill_2 FILLER_26_504 ();
 sg13g2_fill_1 FILLER_26_515 ();
 sg13g2_decap_4 FILLER_26_537 ();
 sg13g2_fill_2 FILLER_26_567 ();
 sg13g2_fill_1 FILLER_26_569 ();
 sg13g2_decap_8 FILLER_26_573 ();
 sg13g2_decap_8 FILLER_26_580 ();
 sg13g2_fill_2 FILLER_26_587 ();
 sg13g2_fill_1 FILLER_26_589 ();
 sg13g2_decap_8 FILLER_26_598 ();
 sg13g2_decap_8 FILLER_26_605 ();
 sg13g2_decap_8 FILLER_26_612 ();
 sg13g2_decap_8 FILLER_26_619 ();
 sg13g2_fill_2 FILLER_26_631 ();
 sg13g2_decap_8 FILLER_26_637 ();
 sg13g2_fill_2 FILLER_26_644 ();
 sg13g2_fill_1 FILLER_26_646 ();
 sg13g2_decap_4 FILLER_26_659 ();
 sg13g2_fill_1 FILLER_26_663 ();
 sg13g2_decap_8 FILLER_26_672 ();
 sg13g2_decap_4 FILLER_26_679 ();
 sg13g2_fill_2 FILLER_26_683 ();
 sg13g2_fill_2 FILLER_26_689 ();
 sg13g2_fill_1 FILLER_26_691 ();
 sg13g2_decap_8 FILLER_26_707 ();
 sg13g2_decap_8 FILLER_26_714 ();
 sg13g2_decap_8 FILLER_26_721 ();
 sg13g2_decap_8 FILLER_26_728 ();
 sg13g2_decap_8 FILLER_26_735 ();
 sg13g2_fill_2 FILLER_26_742 ();
 sg13g2_fill_1 FILLER_26_744 ();
 sg13g2_fill_2 FILLER_26_748 ();
 sg13g2_fill_1 FILLER_26_750 ();
 sg13g2_decap_8 FILLER_26_756 ();
 sg13g2_fill_2 FILLER_26_763 ();
 sg13g2_fill_1 FILLER_26_765 ();
 sg13g2_decap_8 FILLER_26_772 ();
 sg13g2_decap_8 FILLER_26_779 ();
 sg13g2_decap_8 FILLER_26_786 ();
 sg13g2_fill_2 FILLER_26_793 ();
 sg13g2_fill_2 FILLER_26_825 ();
 sg13g2_decap_4 FILLER_26_863 ();
 sg13g2_fill_2 FILLER_26_867 ();
 sg13g2_fill_2 FILLER_26_941 ();
 sg13g2_fill_1 FILLER_26_969 ();
 sg13g2_fill_1 FILLER_26_1000 ();
 sg13g2_fill_1 FILLER_26_1016 ();
 sg13g2_fill_2 FILLER_26_1052 ();
 sg13g2_fill_1 FILLER_26_1054 ();
 sg13g2_decap_8 FILLER_26_1063 ();
 sg13g2_fill_1 FILLER_26_1070 ();
 sg13g2_decap_8 FILLER_26_1074 ();
 sg13g2_decap_8 FILLER_26_1081 ();
 sg13g2_decap_8 FILLER_26_1088 ();
 sg13g2_fill_1 FILLER_26_1095 ();
 sg13g2_fill_2 FILLER_26_1122 ();
 sg13g2_fill_1 FILLER_26_1132 ();
 sg13g2_fill_2 FILLER_26_1142 ();
 sg13g2_decap_8 FILLER_26_1148 ();
 sg13g2_decap_8 FILLER_26_1155 ();
 sg13g2_decap_4 FILLER_26_1162 ();
 sg13g2_fill_2 FILLER_26_1166 ();
 sg13g2_fill_2 FILLER_26_1173 ();
 sg13g2_fill_2 FILLER_26_1179 ();
 sg13g2_fill_1 FILLER_26_1181 ();
 sg13g2_decap_8 FILLER_26_1187 ();
 sg13g2_decap_4 FILLER_26_1194 ();
 sg13g2_fill_2 FILLER_26_1228 ();
 sg13g2_fill_1 FILLER_26_1236 ();
 sg13g2_fill_2 FILLER_26_1252 ();
 sg13g2_fill_1 FILLER_26_1275 ();
 sg13g2_decap_8 FILLER_26_1327 ();
 sg13g2_decap_8 FILLER_26_1334 ();
 sg13g2_decap_8 FILLER_26_1341 ();
 sg13g2_decap_8 FILLER_26_1348 ();
 sg13g2_decap_8 FILLER_26_1355 ();
 sg13g2_decap_8 FILLER_26_1362 ();
 sg13g2_decap_8 FILLER_26_1369 ();
 sg13g2_decap_8 FILLER_26_1376 ();
 sg13g2_decap_8 FILLER_26_1383 ();
 sg13g2_decap_4 FILLER_26_1394 ();
 sg13g2_fill_1 FILLER_26_1398 ();
 sg13g2_decap_8 FILLER_26_1403 ();
 sg13g2_decap_8 FILLER_26_1410 ();
 sg13g2_decap_8 FILLER_26_1417 ();
 sg13g2_decap_8 FILLER_26_1424 ();
 sg13g2_decap_8 FILLER_26_1431 ();
 sg13g2_fill_2 FILLER_26_1441 ();
 sg13g2_decap_4 FILLER_26_1455 ();
 sg13g2_fill_2 FILLER_26_1459 ();
 sg13g2_fill_2 FILLER_26_1465 ();
 sg13g2_decap_8 FILLER_26_1471 ();
 sg13g2_decap_8 FILLER_26_1478 ();
 sg13g2_decap_8 FILLER_26_1485 ();
 sg13g2_decap_8 FILLER_26_1492 ();
 sg13g2_fill_2 FILLER_26_1499 ();
 sg13g2_fill_2 FILLER_26_1505 ();
 sg13g2_fill_1 FILLER_26_1507 ();
 sg13g2_decap_4 FILLER_26_1512 ();
 sg13g2_decap_8 FILLER_26_1519 ();
 sg13g2_fill_1 FILLER_26_1526 ();
 sg13g2_decap_8 FILLER_26_1562 ();
 sg13g2_decap_8 FILLER_26_1569 ();
 sg13g2_decap_8 FILLER_26_1576 ();
 sg13g2_fill_2 FILLER_26_1583 ();
 sg13g2_fill_1 FILLER_26_1585 ();
 sg13g2_decap_8 FILLER_26_1642 ();
 sg13g2_decap_4 FILLER_26_1649 ();
 sg13g2_decap_8 FILLER_26_1691 ();
 sg13g2_fill_1 FILLER_26_1698 ();
 sg13g2_fill_2 FILLER_26_1725 ();
 sg13g2_fill_1 FILLER_26_1761 ();
 sg13g2_fill_2 FILLER_26_1824 ();
 sg13g2_fill_2 FILLER_26_1860 ();
 sg13g2_decap_8 FILLER_26_1872 ();
 sg13g2_decap_8 FILLER_26_1879 ();
 sg13g2_fill_2 FILLER_26_1886 ();
 sg13g2_fill_1 FILLER_26_1888 ();
 sg13g2_decap_8 FILLER_26_1892 ();
 sg13g2_fill_1 FILLER_26_1948 ();
 sg13g2_fill_2 FILLER_26_1967 ();
 sg13g2_decap_4 FILLER_26_1977 ();
 sg13g2_fill_2 FILLER_26_1981 ();
 sg13g2_fill_2 FILLER_26_1988 ();
 sg13g2_decap_8 FILLER_26_2003 ();
 sg13g2_decap_4 FILLER_26_2010 ();
 sg13g2_fill_2 FILLER_26_2014 ();
 sg13g2_fill_2 FILLER_26_2021 ();
 sg13g2_fill_1 FILLER_26_2023 ();
 sg13g2_fill_2 FILLER_26_2034 ();
 sg13g2_decap_8 FILLER_26_2049 ();
 sg13g2_decap_4 FILLER_26_2056 ();
 sg13g2_fill_1 FILLER_26_2060 ();
 sg13g2_decap_8 FILLER_26_2067 ();
 sg13g2_decap_8 FILLER_26_2074 ();
 sg13g2_decap_8 FILLER_26_2081 ();
 sg13g2_decap_4 FILLER_26_2088 ();
 sg13g2_fill_2 FILLER_26_2092 ();
 sg13g2_decap_8 FILLER_26_2138 ();
 sg13g2_decap_8 FILLER_26_2145 ();
 sg13g2_decap_8 FILLER_26_2152 ();
 sg13g2_fill_1 FILLER_26_2159 ();
 sg13g2_decap_4 FILLER_26_2186 ();
 sg13g2_fill_2 FILLER_26_2190 ();
 sg13g2_decap_8 FILLER_26_2196 ();
 sg13g2_decap_4 FILLER_26_2203 ();
 sg13g2_fill_2 FILLER_26_2207 ();
 sg13g2_fill_2 FILLER_26_2214 ();
 sg13g2_fill_1 FILLER_26_2216 ();
 sg13g2_fill_2 FILLER_26_2221 ();
 sg13g2_fill_1 FILLER_26_2223 ();
 sg13g2_decap_8 FILLER_26_2228 ();
 sg13g2_decap_8 FILLER_26_2270 ();
 sg13g2_decap_8 FILLER_26_2285 ();
 sg13g2_decap_8 FILLER_26_2292 ();
 sg13g2_fill_1 FILLER_26_2310 ();
 sg13g2_fill_1 FILLER_26_2328 ();
 sg13g2_fill_2 FILLER_26_2335 ();
 sg13g2_fill_1 FILLER_26_2350 ();
 sg13g2_fill_1 FILLER_26_2371 ();
 sg13g2_decap_8 FILLER_26_2403 ();
 sg13g2_decap_8 FILLER_26_2410 ();
 sg13g2_decap_8 FILLER_26_2417 ();
 sg13g2_fill_1 FILLER_26_2424 ();
 sg13g2_decap_4 FILLER_26_2451 ();
 sg13g2_fill_1 FILLER_26_2455 ();
 sg13g2_decap_8 FILLER_26_2460 ();
 sg13g2_fill_2 FILLER_26_2467 ();
 sg13g2_fill_1 FILLER_26_2469 ();
 sg13g2_decap_8 FILLER_26_2474 ();
 sg13g2_decap_8 FILLER_26_2481 ();
 sg13g2_fill_1 FILLER_26_2488 ();
 sg13g2_fill_1 FILLER_26_2506 ();
 sg13g2_decap_8 FILLER_26_2525 ();
 sg13g2_decap_8 FILLER_26_2532 ();
 sg13g2_decap_4 FILLER_26_2539 ();
 sg13g2_fill_2 FILLER_26_2543 ();
 sg13g2_decap_8 FILLER_26_2554 ();
 sg13g2_decap_8 FILLER_26_2561 ();
 sg13g2_fill_2 FILLER_26_2568 ();
 sg13g2_fill_1 FILLER_26_2579 ();
 sg13g2_fill_1 FILLER_26_2606 ();
 sg13g2_decap_8 FILLER_26_2637 ();
 sg13g2_decap_8 FILLER_26_2644 ();
 sg13g2_decap_8 FILLER_26_2651 ();
 sg13g2_decap_8 FILLER_26_2658 ();
 sg13g2_decap_4 FILLER_26_2665 ();
 sg13g2_fill_1 FILLER_26_2669 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_fill_1 FILLER_27_60 ();
 sg13g2_decap_8 FILLER_27_74 ();
 sg13g2_decap_8 FILLER_27_81 ();
 sg13g2_decap_4 FILLER_27_88 ();
 sg13g2_fill_2 FILLER_27_92 ();
 sg13g2_fill_1 FILLER_27_102 ();
 sg13g2_decap_4 FILLER_27_124 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_4 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_187 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_fill_1 FILLER_27_290 ();
 sg13g2_decap_4 FILLER_27_300 ();
 sg13g2_fill_1 FILLER_27_304 ();
 sg13g2_decap_4 FILLER_27_309 ();
 sg13g2_fill_2 FILLER_27_313 ();
 sg13g2_fill_1 FILLER_27_320 ();
 sg13g2_fill_2 FILLER_27_326 ();
 sg13g2_fill_2 FILLER_27_333 ();
 sg13g2_decap_4 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_fill_2 FILLER_27_401 ();
 sg13g2_fill_2 FILLER_27_417 ();
 sg13g2_fill_1 FILLER_27_419 ();
 sg13g2_decap_8 FILLER_27_425 ();
 sg13g2_decap_8 FILLER_27_432 ();
 sg13g2_decap_8 FILLER_27_449 ();
 sg13g2_decap_8 FILLER_27_456 ();
 sg13g2_decap_8 FILLER_27_463 ();
 sg13g2_fill_1 FILLER_27_476 ();
 sg13g2_fill_1 FILLER_27_480 ();
 sg13g2_fill_1 FILLER_27_486 ();
 sg13g2_fill_1 FILLER_27_494 ();
 sg13g2_fill_1 FILLER_27_499 ();
 sg13g2_fill_2 FILLER_27_504 ();
 sg13g2_decap_4 FILLER_27_532 ();
 sg13g2_fill_2 FILLER_27_536 ();
 sg13g2_decap_8 FILLER_27_551 ();
 sg13g2_fill_1 FILLER_27_558 ();
 sg13g2_decap_8 FILLER_27_579 ();
 sg13g2_decap_4 FILLER_27_586 ();
 sg13g2_decap_8 FILLER_27_603 ();
 sg13g2_decap_8 FILLER_27_610 ();
 sg13g2_fill_2 FILLER_27_617 ();
 sg13g2_fill_1 FILLER_27_619 ();
 sg13g2_decap_4 FILLER_27_632 ();
 sg13g2_fill_1 FILLER_27_636 ();
 sg13g2_decap_8 FILLER_27_660 ();
 sg13g2_fill_2 FILLER_27_667 ();
 sg13g2_fill_1 FILLER_27_669 ();
 sg13g2_decap_8 FILLER_27_673 ();
 sg13g2_fill_2 FILLER_27_680 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_fill_1 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_711 ();
 sg13g2_decap_4 FILLER_27_718 ();
 sg13g2_fill_1 FILLER_27_722 ();
 sg13g2_decap_8 FILLER_27_726 ();
 sg13g2_decap_4 FILLER_27_733 ();
 sg13g2_fill_2 FILLER_27_737 ();
 sg13g2_fill_1 FILLER_27_765 ();
 sg13g2_fill_1 FILLER_27_777 ();
 sg13g2_fill_2 FILLER_27_783 ();
 sg13g2_decap_8 FILLER_27_832 ();
 sg13g2_fill_1 FILLER_27_839 ();
 sg13g2_decap_8 FILLER_27_844 ();
 sg13g2_decap_4 FILLER_27_851 ();
 sg13g2_fill_1 FILLER_27_855 ();
 sg13g2_decap_8 FILLER_27_860 ();
 sg13g2_decap_4 FILLER_27_867 ();
 sg13g2_decap_8 FILLER_27_875 ();
 sg13g2_decap_8 FILLER_27_882 ();
 sg13g2_fill_2 FILLER_27_889 ();
 sg13g2_fill_1 FILLER_27_891 ();
 sg13g2_decap_8 FILLER_27_922 ();
 sg13g2_decap_8 FILLER_27_933 ();
 sg13g2_decap_4 FILLER_27_940 ();
 sg13g2_fill_1 FILLER_27_944 ();
 sg13g2_fill_1 FILLER_27_985 ();
 sg13g2_fill_1 FILLER_27_1005 ();
 sg13g2_fill_2 FILLER_27_1017 ();
 sg13g2_fill_1 FILLER_27_1032 ();
 sg13g2_decap_4 FILLER_27_1052 ();
 sg13g2_fill_2 FILLER_27_1056 ();
 sg13g2_fill_2 FILLER_27_1079 ();
 sg13g2_decap_8 FILLER_27_1089 ();
 sg13g2_fill_1 FILLER_27_1096 ();
 sg13g2_fill_1 FILLER_27_1123 ();
 sg13g2_decap_4 FILLER_27_1127 ();
 sg13g2_fill_1 FILLER_27_1131 ();
 sg13g2_decap_8 FILLER_27_1169 ();
 sg13g2_decap_8 FILLER_27_1176 ();
 sg13g2_decap_8 FILLER_27_1183 ();
 sg13g2_decap_8 FILLER_27_1190 ();
 sg13g2_decap_8 FILLER_27_1197 ();
 sg13g2_decap_8 FILLER_27_1204 ();
 sg13g2_decap_8 FILLER_27_1216 ();
 sg13g2_fill_2 FILLER_27_1229 ();
 sg13g2_fill_2 FILLER_27_1236 ();
 sg13g2_decap_4 FILLER_27_1244 ();
 sg13g2_decap_8 FILLER_27_1321 ();
 sg13g2_decap_4 FILLER_27_1328 ();
 sg13g2_fill_1 FILLER_27_1332 ();
 sg13g2_fill_1 FILLER_27_1341 ();
 sg13g2_fill_2 FILLER_27_1377 ();
 sg13g2_fill_1 FILLER_27_1387 ();
 sg13g2_fill_1 FILLER_27_1392 ();
 sg13g2_fill_2 FILLER_27_1397 ();
 sg13g2_fill_1 FILLER_27_1399 ();
 sg13g2_decap_8 FILLER_27_1404 ();
 sg13g2_decap_8 FILLER_27_1411 ();
 sg13g2_decap_8 FILLER_27_1418 ();
 sg13g2_decap_8 FILLER_27_1425 ();
 sg13g2_decap_8 FILLER_27_1432 ();
 sg13g2_fill_1 FILLER_27_1439 ();
 sg13g2_decap_8 FILLER_27_1445 ();
 sg13g2_decap_8 FILLER_27_1452 ();
 sg13g2_fill_2 FILLER_27_1459 ();
 sg13g2_fill_1 FILLER_27_1461 ();
 sg13g2_decap_8 FILLER_27_1466 ();
 sg13g2_decap_4 FILLER_27_1473 ();
 sg13g2_fill_1 FILLER_27_1477 ();
 sg13g2_decap_8 FILLER_27_1517 ();
 sg13g2_decap_8 FILLER_27_1524 ();
 sg13g2_decap_8 FILLER_27_1531 ();
 sg13g2_fill_1 FILLER_27_1538 ();
 sg13g2_decap_8 FILLER_27_1556 ();
 sg13g2_decap_8 FILLER_27_1563 ();
 sg13g2_decap_4 FILLER_27_1570 ();
 sg13g2_decap_4 FILLER_27_1582 ();
 sg13g2_fill_1 FILLER_27_1590 ();
 sg13g2_decap_8 FILLER_27_1621 ();
 sg13g2_decap_8 FILLER_27_1628 ();
 sg13g2_decap_8 FILLER_27_1635 ();
 sg13g2_decap_4 FILLER_27_1642 ();
 sg13g2_fill_1 FILLER_27_1659 ();
 sg13g2_decap_4 FILLER_27_1665 ();
 sg13g2_decap_8 FILLER_27_1684 ();
 sg13g2_decap_4 FILLER_27_1691 ();
 sg13g2_fill_1 FILLER_27_1695 ();
 sg13g2_fill_2 FILLER_27_1714 ();
 sg13g2_fill_2 FILLER_27_1720 ();
 sg13g2_fill_1 FILLER_27_1722 ();
 sg13g2_decap_8 FILLER_27_1768 ();
 sg13g2_fill_2 FILLER_27_1775 ();
 sg13g2_fill_1 FILLER_27_1777 ();
 sg13g2_fill_2 FILLER_27_1793 ();
 sg13g2_decap_8 FILLER_27_1799 ();
 sg13g2_fill_2 FILLER_27_1842 ();
 sg13g2_fill_1 FILLER_27_1844 ();
 sg13g2_decap_4 FILLER_27_1881 ();
 sg13g2_fill_1 FILLER_27_1885 ();
 sg13g2_fill_2 FILLER_27_1899 ();
 sg13g2_fill_2 FILLER_27_1905 ();
 sg13g2_fill_2 FILLER_27_1915 ();
 sg13g2_fill_1 FILLER_27_1917 ();
 sg13g2_decap_8 FILLER_27_1939 ();
 sg13g2_decap_4 FILLER_27_1952 ();
 sg13g2_fill_2 FILLER_27_1956 ();
 sg13g2_decap_8 FILLER_27_1984 ();
 sg13g2_fill_1 FILLER_27_2000 ();
 sg13g2_fill_1 FILLER_27_2015 ();
 sg13g2_fill_2 FILLER_27_2020 ();
 sg13g2_fill_1 FILLER_27_2022 ();
 sg13g2_decap_4 FILLER_27_2054 ();
 sg13g2_fill_2 FILLER_27_2071 ();
 sg13g2_decap_8 FILLER_27_2079 ();
 sg13g2_decap_8 FILLER_27_2086 ();
 sg13g2_decap_4 FILLER_27_2093 ();
 sg13g2_fill_2 FILLER_27_2097 ();
 sg13g2_decap_8 FILLER_27_2125 ();
 sg13g2_decap_8 FILLER_27_2132 ();
 sg13g2_fill_1 FILLER_27_2139 ();
 sg13g2_decap_8 FILLER_27_2179 ();
 sg13g2_decap_8 FILLER_27_2186 ();
 sg13g2_decap_4 FILLER_27_2193 ();
 sg13g2_fill_1 FILLER_27_2197 ();
 sg13g2_fill_1 FILLER_27_2201 ();
 sg13g2_fill_1 FILLER_27_2208 ();
 sg13g2_decap_8 FILLER_27_2214 ();
 sg13g2_decap_8 FILLER_27_2221 ();
 sg13g2_decap_8 FILLER_27_2228 ();
 sg13g2_decap_4 FILLER_27_2235 ();
 sg13g2_decap_8 FILLER_27_2243 ();
 sg13g2_decap_8 FILLER_27_2250 ();
 sg13g2_fill_1 FILLER_27_2257 ();
 sg13g2_fill_2 FILLER_27_2279 ();
 sg13g2_decap_8 FILLER_27_2291 ();
 sg13g2_fill_2 FILLER_27_2302 ();
 sg13g2_fill_1 FILLER_27_2310 ();
 sg13g2_fill_2 FILLER_27_2324 ();
 sg13g2_fill_2 FILLER_27_2332 ();
 sg13g2_decap_4 FILLER_27_2377 ();
 sg13g2_fill_1 FILLER_27_2381 ();
 sg13g2_decap_8 FILLER_27_2408 ();
 sg13g2_decap_8 FILLER_27_2415 ();
 sg13g2_decap_8 FILLER_27_2422 ();
 sg13g2_fill_1 FILLER_27_2429 ();
 sg13g2_fill_2 FILLER_27_2434 ();
 sg13g2_decap_8 FILLER_27_2440 ();
 sg13g2_decap_8 FILLER_27_2447 ();
 sg13g2_decap_4 FILLER_27_2454 ();
 sg13g2_fill_1 FILLER_27_2458 ();
 sg13g2_decap_8 FILLER_27_2463 ();
 sg13g2_decap_4 FILLER_27_2470 ();
 sg13g2_fill_1 FILLER_27_2474 ();
 sg13g2_fill_1 FILLER_27_2481 ();
 sg13g2_decap_8 FILLER_27_2520 ();
 sg13g2_decap_8 FILLER_27_2527 ();
 sg13g2_decap_8 FILLER_27_2534 ();
 sg13g2_decap_8 FILLER_27_2541 ();
 sg13g2_decap_8 FILLER_27_2548 ();
 sg13g2_decap_8 FILLER_27_2555 ();
 sg13g2_fill_2 FILLER_27_2592 ();
 sg13g2_fill_2 FILLER_27_2611 ();
 sg13g2_fill_1 FILLER_27_2613 ();
 sg13g2_decap_8 FILLER_27_2644 ();
 sg13g2_decap_8 FILLER_27_2651 ();
 sg13g2_decap_8 FILLER_27_2658 ();
 sg13g2_decap_4 FILLER_27_2665 ();
 sg13g2_fill_1 FILLER_27_2669 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_38 ();
 sg13g2_decap_8 FILLER_28_45 ();
 sg13g2_fill_1 FILLER_28_52 ();
 sg13g2_decap_8 FILLER_28_57 ();
 sg13g2_decap_8 FILLER_28_64 ();
 sg13g2_decap_8 FILLER_28_71 ();
 sg13g2_decap_8 FILLER_28_78 ();
 sg13g2_decap_4 FILLER_28_85 ();
 sg13g2_fill_1 FILLER_28_89 ();
 sg13g2_decap_8 FILLER_28_127 ();
 sg13g2_decap_8 FILLER_28_134 ();
 sg13g2_decap_8 FILLER_28_141 ();
 sg13g2_decap_4 FILLER_28_148 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_decap_8 FILLER_28_179 ();
 sg13g2_decap_8 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_fill_2 FILLER_28_287 ();
 sg13g2_fill_1 FILLER_28_289 ();
 sg13g2_decap_8 FILLER_28_295 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_decap_4 FILLER_28_308 ();
 sg13g2_fill_1 FILLER_28_312 ();
 sg13g2_fill_2 FILLER_28_333 ();
 sg13g2_fill_1 FILLER_28_335 ();
 sg13g2_decap_4 FILLER_28_348 ();
 sg13g2_fill_2 FILLER_28_352 ();
 sg13g2_fill_2 FILLER_28_424 ();
 sg13g2_decap_4 FILLER_28_434 ();
 sg13g2_fill_2 FILLER_28_448 ();
 sg13g2_fill_1 FILLER_28_450 ();
 sg13g2_decap_8 FILLER_28_455 ();
 sg13g2_decap_4 FILLER_28_462 ();
 sg13g2_fill_1 FILLER_28_466 ();
 sg13g2_fill_1 FILLER_28_471 ();
 sg13g2_fill_2 FILLER_28_477 ();
 sg13g2_fill_1 FILLER_28_479 ();
 sg13g2_decap_8 FILLER_28_515 ();
 sg13g2_decap_4 FILLER_28_522 ();
 sg13g2_fill_2 FILLER_28_526 ();
 sg13g2_decap_4 FILLER_28_536 ();
 sg13g2_fill_2 FILLER_28_614 ();
 sg13g2_fill_1 FILLER_28_621 ();
 sg13g2_decap_8 FILLER_28_627 ();
 sg13g2_fill_1 FILLER_28_634 ();
 sg13g2_decap_8 FILLER_28_648 ();
 sg13g2_decap_8 FILLER_28_655 ();
 sg13g2_decap_8 FILLER_28_662 ();
 sg13g2_decap_8 FILLER_28_669 ();
 sg13g2_decap_8 FILLER_28_676 ();
 sg13g2_fill_2 FILLER_28_683 ();
 sg13g2_fill_1 FILLER_28_694 ();
 sg13g2_fill_1 FILLER_28_702 ();
 sg13g2_decap_4 FILLER_28_708 ();
 sg13g2_decap_8 FILLER_28_729 ();
 sg13g2_decap_8 FILLER_28_736 ();
 sg13g2_decap_4 FILLER_28_743 ();
 sg13g2_fill_1 FILLER_28_747 ();
 sg13g2_fill_1 FILLER_28_753 ();
 sg13g2_decap_8 FILLER_28_774 ();
 sg13g2_fill_2 FILLER_28_781 ();
 sg13g2_decap_8 FILLER_28_830 ();
 sg13g2_decap_4 FILLER_28_837 ();
 sg13g2_fill_2 FILLER_28_841 ();
 sg13g2_decap_8 FILLER_28_848 ();
 sg13g2_decap_8 FILLER_28_855 ();
 sg13g2_decap_4 FILLER_28_862 ();
 sg13g2_fill_2 FILLER_28_866 ();
 sg13g2_decap_8 FILLER_28_872 ();
 sg13g2_decap_8 FILLER_28_879 ();
 sg13g2_fill_2 FILLER_28_947 ();
 sg13g2_fill_2 FILLER_28_953 ();
 sg13g2_decap_8 FILLER_28_963 ();
 sg13g2_decap_8 FILLER_28_970 ();
 sg13g2_fill_2 FILLER_28_992 ();
 sg13g2_fill_2 FILLER_28_1005 ();
 sg13g2_fill_1 FILLER_28_1030 ();
 sg13g2_fill_1 FILLER_28_1057 ();
 sg13g2_fill_1 FILLER_28_1063 ();
 sg13g2_fill_1 FILLER_28_1069 ();
 sg13g2_decap_8 FILLER_28_1096 ();
 sg13g2_decap_8 FILLER_28_1103 ();
 sg13g2_fill_2 FILLER_28_1110 ();
 sg13g2_decap_4 FILLER_28_1115 ();
 sg13g2_fill_2 FILLER_28_1119 ();
 sg13g2_fill_1 FILLER_28_1139 ();
 sg13g2_decap_8 FILLER_28_1171 ();
 sg13g2_fill_2 FILLER_28_1178 ();
 sg13g2_fill_2 FILLER_28_1185 ();
 sg13g2_decap_8 FILLER_28_1191 ();
 sg13g2_decap_8 FILLER_28_1198 ();
 sg13g2_fill_1 FILLER_28_1205 ();
 sg13g2_decap_8 FILLER_28_1215 ();
 sg13g2_decap_4 FILLER_28_1222 ();
 sg13g2_fill_1 FILLER_28_1226 ();
 sg13g2_decap_8 FILLER_28_1232 ();
 sg13g2_fill_2 FILLER_28_1239 ();
 sg13g2_fill_1 FILLER_28_1247 ();
 sg13g2_fill_2 FILLER_28_1262 ();
 sg13g2_decap_8 FILLER_28_1293 ();
 sg13g2_decap_8 FILLER_28_1340 ();
 sg13g2_fill_2 FILLER_28_1347 ();
 sg13g2_fill_1 FILLER_28_1349 ();
 sg13g2_decap_8 FILLER_28_1354 ();
 sg13g2_decap_8 FILLER_28_1361 ();
 sg13g2_decap_4 FILLER_28_1368 ();
 sg13g2_fill_2 FILLER_28_1372 ();
 sg13g2_decap_4 FILLER_28_1398 ();
 sg13g2_decap_8 FILLER_28_1408 ();
 sg13g2_fill_1 FILLER_28_1415 ();
 sg13g2_decap_4 FILLER_28_1424 ();
 sg13g2_fill_2 FILLER_28_1432 ();
 sg13g2_fill_1 FILLER_28_1434 ();
 sg13g2_decap_8 FILLER_28_1441 ();
 sg13g2_decap_4 FILLER_28_1448 ();
 sg13g2_fill_1 FILLER_28_1452 ();
 sg13g2_decap_4 FILLER_28_1461 ();
 sg13g2_decap_8 FILLER_28_1559 ();
 sg13g2_decap_8 FILLER_28_1566 ();
 sg13g2_decap_8 FILLER_28_1573 ();
 sg13g2_decap_4 FILLER_28_1580 ();
 sg13g2_fill_1 FILLER_28_1584 ();
 sg13g2_fill_1 FILLER_28_1615 ();
 sg13g2_decap_8 FILLER_28_1621 ();
 sg13g2_decap_4 FILLER_28_1628 ();
 sg13g2_fill_2 FILLER_28_1632 ();
 sg13g2_decap_4 FILLER_28_1663 ();
 sg13g2_decap_8 FILLER_28_1686 ();
 sg13g2_decap_4 FILLER_28_1693 ();
 sg13g2_fill_2 FILLER_28_1697 ();
 sg13g2_decap_8 FILLER_28_1760 ();
 sg13g2_decap_4 FILLER_28_1767 ();
 sg13g2_fill_2 FILLER_28_1771 ();
 sg13g2_decap_8 FILLER_28_1779 ();
 sg13g2_decap_8 FILLER_28_1786 ();
 sg13g2_decap_8 FILLER_28_1793 ();
 sg13g2_decap_8 FILLER_28_1800 ();
 sg13g2_fill_1 FILLER_28_1807 ();
 sg13g2_decap_4 FILLER_28_1813 ();
 sg13g2_fill_2 FILLER_28_1817 ();
 sg13g2_fill_2 FILLER_28_1828 ();
 sg13g2_decap_8 FILLER_28_1886 ();
 sg13g2_decap_8 FILLER_28_1893 ();
 sg13g2_fill_2 FILLER_28_1900 ();
 sg13g2_decap_4 FILLER_28_1915 ();
 sg13g2_decap_4 FILLER_28_1958 ();
 sg13g2_decap_8 FILLER_28_1971 ();
 sg13g2_decap_4 FILLER_28_1978 ();
 sg13g2_fill_1 FILLER_28_1982 ();
 sg13g2_fill_2 FILLER_28_1995 ();
 sg13g2_fill_2 FILLER_28_2055 ();
 sg13g2_fill_1 FILLER_28_2057 ();
 sg13g2_fill_1 FILLER_28_2090 ();
 sg13g2_decap_8 FILLER_28_2095 ();
 sg13g2_fill_2 FILLER_28_2102 ();
 sg13g2_decap_8 FILLER_28_2139 ();
 sg13g2_decap_8 FILLER_28_2146 ();
 sg13g2_decap_4 FILLER_28_2153 ();
 sg13g2_fill_1 FILLER_28_2157 ();
 sg13g2_decap_4 FILLER_28_2167 ();
 sg13g2_fill_2 FILLER_28_2171 ();
 sg13g2_decap_8 FILLER_28_2183 ();
 sg13g2_fill_2 FILLER_28_2190 ();
 sg13g2_fill_2 FILLER_28_2213 ();
 sg13g2_decap_4 FILLER_28_2245 ();
 sg13g2_decap_4 FILLER_28_2253 ();
 sg13g2_fill_2 FILLER_28_2257 ();
 sg13g2_decap_4 FILLER_28_2268 ();
 sg13g2_fill_1 FILLER_28_2272 ();
 sg13g2_fill_1 FILLER_28_2277 ();
 sg13g2_fill_2 FILLER_28_2304 ();
 sg13g2_fill_1 FILLER_28_2310 ();
 sg13g2_fill_1 FILLER_28_2325 ();
 sg13g2_fill_1 FILLER_28_2364 ();
 sg13g2_fill_1 FILLER_28_2378 ();
 sg13g2_decap_4 FILLER_28_2397 ();
 sg13g2_fill_1 FILLER_28_2401 ();
 sg13g2_decap_4 FILLER_28_2408 ();
 sg13g2_fill_2 FILLER_28_2412 ();
 sg13g2_decap_8 FILLER_28_2422 ();
 sg13g2_decap_8 FILLER_28_2429 ();
 sg13g2_decap_4 FILLER_28_2436 ();
 sg13g2_fill_2 FILLER_28_2440 ();
 sg13g2_fill_1 FILLER_28_2447 ();
 sg13g2_fill_1 FILLER_28_2478 ();
 sg13g2_decap_8 FILLER_28_2497 ();
 sg13g2_decap_8 FILLER_28_2504 ();
 sg13g2_decap_8 FILLER_28_2511 ();
 sg13g2_decap_8 FILLER_28_2518 ();
 sg13g2_fill_2 FILLER_28_2525 ();
 sg13g2_fill_1 FILLER_28_2527 ();
 sg13g2_decap_4 FILLER_28_2537 ();
 sg13g2_fill_1 FILLER_28_2541 ();
 sg13g2_decap_4 FILLER_28_2568 ();
 sg13g2_fill_1 FILLER_28_2572 ();
 sg13g2_decap_8 FILLER_28_2577 ();
 sg13g2_decap_8 FILLER_28_2584 ();
 sg13g2_fill_1 FILLER_28_2591 ();
 sg13g2_decap_8 FILLER_28_2596 ();
 sg13g2_decap_4 FILLER_28_2603 ();
 sg13g2_fill_1 FILLER_28_2607 ();
 sg13g2_decap_8 FILLER_28_2638 ();
 sg13g2_decap_8 FILLER_28_2645 ();
 sg13g2_decap_8 FILLER_28_2652 ();
 sg13g2_decap_8 FILLER_28_2659 ();
 sg13g2_decap_4 FILLER_28_2666 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_11 ();
 sg13g2_decap_4 FILLER_29_25 ();
 sg13g2_fill_1 FILLER_29_29 ();
 sg13g2_decap_8 FILLER_29_38 ();
 sg13g2_decap_4 FILLER_29_45 ();
 sg13g2_fill_2 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_81 ();
 sg13g2_fill_2 FILLER_29_88 ();
 sg13g2_fill_1 FILLER_29_90 ();
 sg13g2_decap_8 FILLER_29_135 ();
 sg13g2_fill_2 FILLER_29_142 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_162 ();
 sg13g2_decap_8 FILLER_29_169 ();
 sg13g2_decap_8 FILLER_29_176 ();
 sg13g2_decap_8 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_220 ();
 sg13g2_fill_1 FILLER_29_234 ();
 sg13g2_fill_2 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_240 ();
 sg13g2_fill_1 FILLER_29_260 ();
 sg13g2_fill_2 FILLER_29_299 ();
 sg13g2_decap_4 FILLER_29_306 ();
 sg13g2_fill_1 FILLER_29_315 ();
 sg13g2_fill_1 FILLER_29_342 ();
 sg13g2_fill_1 FILLER_29_348 ();
 sg13g2_fill_2 FILLER_29_440 ();
 sg13g2_fill_2 FILLER_29_452 ();
 sg13g2_fill_2 FILLER_29_462 ();
 sg13g2_fill_1 FILLER_29_464 ();
 sg13g2_decap_8 FILLER_29_491 ();
 sg13g2_fill_2 FILLER_29_498 ();
 sg13g2_decap_8 FILLER_29_505 ();
 sg13g2_decap_8 FILLER_29_512 ();
 sg13g2_decap_8 FILLER_29_519 ();
 sg13g2_decap_4 FILLER_29_526 ();
 sg13g2_fill_1 FILLER_29_530 ();
 sg13g2_decap_8 FILLER_29_561 ();
 sg13g2_decap_8 FILLER_29_568 ();
 sg13g2_fill_2 FILLER_29_575 ();
 sg13g2_fill_1 FILLER_29_607 ();
 sg13g2_decap_8 FILLER_29_612 ();
 sg13g2_decap_4 FILLER_29_619 ();
 sg13g2_fill_2 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_640 ();
 sg13g2_decap_8 FILLER_29_647 ();
 sg13g2_decap_4 FILLER_29_654 ();
 sg13g2_fill_1 FILLER_29_658 ();
 sg13g2_decap_8 FILLER_29_669 ();
 sg13g2_decap_4 FILLER_29_676 ();
 sg13g2_fill_1 FILLER_29_680 ();
 sg13g2_fill_1 FILLER_29_694 ();
 sg13g2_fill_1 FILLER_29_701 ();
 sg13g2_fill_1 FILLER_29_711 ();
 sg13g2_fill_1 FILLER_29_727 ();
 sg13g2_fill_2 FILLER_29_744 ();
 sg13g2_fill_2 FILLER_29_751 ();
 sg13g2_decap_8 FILLER_29_779 ();
 sg13g2_fill_2 FILLER_29_786 ();
 sg13g2_fill_1 FILLER_29_788 ();
 sg13g2_fill_2 FILLER_29_793 ();
 sg13g2_decap_8 FILLER_29_799 ();
 sg13g2_decap_4 FILLER_29_806 ();
 sg13g2_decap_4 FILLER_29_819 ();
 sg13g2_fill_2 FILLER_29_875 ();
 sg13g2_decap_8 FILLER_29_881 ();
 sg13g2_fill_1 FILLER_29_888 ();
 sg13g2_decap_4 FILLER_29_901 ();
 sg13g2_decap_8 FILLER_29_958 ();
 sg13g2_fill_1 FILLER_29_965 ();
 sg13g2_fill_2 FILLER_29_972 ();
 sg13g2_fill_1 FILLER_29_977 ();
 sg13g2_fill_1 FILLER_29_1028 ();
 sg13g2_fill_2 FILLER_29_1035 ();
 sg13g2_fill_2 FILLER_29_1042 ();
 sg13g2_fill_2 FILLER_29_1050 ();
 sg13g2_fill_1 FILLER_29_1052 ();
 sg13g2_fill_2 FILLER_29_1063 ();
 sg13g2_fill_1 FILLER_29_1065 ();
 sg13g2_fill_2 FILLER_29_1072 ();
 sg13g2_fill_1 FILLER_29_1074 ();
 sg13g2_fill_2 FILLER_29_1087 ();
 sg13g2_fill_1 FILLER_29_1089 ();
 sg13g2_fill_1 FILLER_29_1132 ();
 sg13g2_fill_1 FILLER_29_1139 ();
 sg13g2_decap_4 FILLER_29_1155 ();
 sg13g2_fill_2 FILLER_29_1256 ();
 sg13g2_decap_4 FILLER_29_1264 ();
 sg13g2_fill_2 FILLER_29_1268 ();
 sg13g2_decap_8 FILLER_29_1289 ();
 sg13g2_decap_8 FILLER_29_1296 ();
 sg13g2_fill_2 FILLER_29_1303 ();
 sg13g2_fill_1 FILLER_29_1305 ();
 sg13g2_decap_4 FILLER_29_1311 ();
 sg13g2_decap_8 FILLER_29_1319 ();
 sg13g2_fill_2 FILLER_29_1326 ();
 sg13g2_fill_1 FILLER_29_1328 ();
 sg13g2_decap_4 FILLER_29_1335 ();
 sg13g2_fill_2 FILLER_29_1343 ();
 sg13g2_fill_2 FILLER_29_1393 ();
 sg13g2_fill_1 FILLER_29_1421 ();
 sg13g2_fill_2 FILLER_29_1448 ();
 sg13g2_decap_8 FILLER_29_1484 ();
 sg13g2_fill_2 FILLER_29_1491 ();
 sg13g2_fill_2 FILLER_29_1501 ();
 sg13g2_fill_1 FILLER_29_1503 ();
 sg13g2_decap_8 FILLER_29_1548 ();
 sg13g2_decap_4 FILLER_29_1555 ();
 sg13g2_fill_1 FILLER_29_1559 ();
 sg13g2_decap_8 FILLER_29_1609 ();
 sg13g2_fill_1 FILLER_29_1664 ();
 sg13g2_fill_2 FILLER_29_1716 ();
 sg13g2_fill_1 FILLER_29_1718 ();
 sg13g2_decap_8 FILLER_29_1728 ();
 sg13g2_decap_8 FILLER_29_1735 ();
 sg13g2_decap_8 FILLER_29_1742 ();
 sg13g2_decap_8 FILLER_29_1749 ();
 sg13g2_fill_2 FILLER_29_1756 ();
 sg13g2_fill_1 FILLER_29_1758 ();
 sg13g2_decap_4 FILLER_29_1799 ();
 sg13g2_fill_1 FILLER_29_1803 ();
 sg13g2_decap_8 FILLER_29_1864 ();
 sg13g2_decap_8 FILLER_29_1871 ();
 sg13g2_fill_2 FILLER_29_1878 ();
 sg13g2_fill_2 FILLER_29_1885 ();
 sg13g2_fill_1 FILLER_29_1887 ();
 sg13g2_decap_8 FILLER_29_1937 ();
 sg13g2_decap_8 FILLER_29_1970 ();
 sg13g2_decap_4 FILLER_29_1977 ();
 sg13g2_fill_1 FILLER_29_1981 ();
 sg13g2_decap_8 FILLER_29_2013 ();
 sg13g2_fill_2 FILLER_29_2020 ();
 sg13g2_fill_1 FILLER_29_2022 ();
 sg13g2_fill_1 FILLER_29_2028 ();
 sg13g2_fill_1 FILLER_29_2050 ();
 sg13g2_decap_4 FILLER_29_2056 ();
 sg13g2_fill_2 FILLER_29_2060 ();
 sg13g2_fill_2 FILLER_29_2099 ();
 sg13g2_fill_1 FILLER_29_2101 ();
 sg13g2_fill_2 FILLER_29_2115 ();
 sg13g2_fill_1 FILLER_29_2117 ();
 sg13g2_decap_8 FILLER_29_2201 ();
 sg13g2_fill_1 FILLER_29_2212 ();
 sg13g2_fill_2 FILLER_29_2217 ();
 sg13g2_decap_8 FILLER_29_2227 ();
 sg13g2_fill_2 FILLER_29_2255 ();
 sg13g2_fill_2 FILLER_29_2266 ();
 sg13g2_fill_2 FILLER_29_2276 ();
 sg13g2_fill_2 FILLER_29_2283 ();
 sg13g2_fill_2 FILLER_29_2311 ();
 sg13g2_decap_8 FILLER_29_2317 ();
 sg13g2_decap_4 FILLER_29_2324 ();
 sg13g2_fill_1 FILLER_29_2328 ();
 sg13g2_fill_1 FILLER_29_2337 ();
 sg13g2_decap_4 FILLER_29_2345 ();
 sg13g2_fill_1 FILLER_29_2349 ();
 sg13g2_fill_1 FILLER_29_2354 ();
 sg13g2_fill_1 FILLER_29_2378 ();
 sg13g2_fill_2 FILLER_29_2405 ();
 sg13g2_fill_2 FILLER_29_2453 ();
 sg13g2_fill_1 FILLER_29_2455 ();
 sg13g2_fill_1 FILLER_29_2491 ();
 sg13g2_fill_1 FILLER_29_2497 ();
 sg13g2_fill_1 FILLER_29_2503 ();
 sg13g2_decap_8 FILLER_29_2530 ();
 sg13g2_fill_1 FILLER_29_2537 ();
 sg13g2_fill_1 FILLER_29_2595 ();
 sg13g2_decap_8 FILLER_29_2626 ();
 sg13g2_decap_8 FILLER_29_2633 ();
 sg13g2_decap_8 FILLER_29_2640 ();
 sg13g2_decap_8 FILLER_29_2647 ();
 sg13g2_decap_8 FILLER_29_2654 ();
 sg13g2_decap_8 FILLER_29_2661 ();
 sg13g2_fill_2 FILLER_29_2668 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_45 ();
 sg13g2_fill_1 FILLER_30_61 ();
 sg13g2_fill_2 FILLER_30_67 ();
 sg13g2_fill_2 FILLER_30_82 ();
 sg13g2_decap_8 FILLER_30_89 ();
 sg13g2_decap_8 FILLER_30_96 ();
 sg13g2_decap_8 FILLER_30_103 ();
 sg13g2_fill_2 FILLER_30_110 ();
 sg13g2_fill_1 FILLER_30_112 ();
 sg13g2_fill_2 FILLER_30_122 ();
 sg13g2_fill_1 FILLER_30_124 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_fill_1 FILLER_30_162 ();
 sg13g2_fill_2 FILLER_30_167 ();
 sg13g2_decap_4 FILLER_30_173 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_decap_4 FILLER_30_183 ();
 sg13g2_fill_1 FILLER_30_187 ();
 sg13g2_decap_8 FILLER_30_218 ();
 sg13g2_decap_4 FILLER_30_225 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_decap_8 FILLER_30_261 ();
 sg13g2_decap_4 FILLER_30_268 ();
 sg13g2_fill_1 FILLER_30_272 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_316 ();
 sg13g2_fill_2 FILLER_30_344 ();
 sg13g2_fill_1 FILLER_30_346 ();
 sg13g2_fill_1 FILLER_30_351 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_1 FILLER_30_368 ();
 sg13g2_fill_2 FILLER_30_373 ();
 sg13g2_fill_2 FILLER_30_379 ();
 sg13g2_fill_1 FILLER_30_381 ();
 sg13g2_fill_1 FILLER_30_393 ();
 sg13g2_fill_2 FILLER_30_398 ();
 sg13g2_fill_1 FILLER_30_400 ();
 sg13g2_fill_1 FILLER_30_426 ();
 sg13g2_decap_8 FILLER_30_471 ();
 sg13g2_decap_4 FILLER_30_478 ();
 sg13g2_fill_2 FILLER_30_482 ();
 sg13g2_decap_8 FILLER_30_489 ();
 sg13g2_fill_1 FILLER_30_496 ();
 sg13g2_fill_2 FILLER_30_507 ();
 sg13g2_decap_8 FILLER_30_518 ();
 sg13g2_decap_8 FILLER_30_525 ();
 sg13g2_decap_4 FILLER_30_532 ();
 sg13g2_fill_1 FILLER_30_541 ();
 sg13g2_decap_8 FILLER_30_546 ();
 sg13g2_decap_8 FILLER_30_553 ();
 sg13g2_decap_8 FILLER_30_560 ();
 sg13g2_decap_4 FILLER_30_567 ();
 sg13g2_fill_2 FILLER_30_571 ();
 sg13g2_fill_2 FILLER_30_582 ();
 sg13g2_decap_4 FILLER_30_624 ();
 sg13g2_decap_8 FILLER_30_638 ();
 sg13g2_decap_8 FILLER_30_645 ();
 sg13g2_decap_4 FILLER_30_652 ();
 sg13g2_fill_1 FILLER_30_661 ();
 sg13g2_decap_8 FILLER_30_666 ();
 sg13g2_fill_1 FILLER_30_673 ();
 sg13g2_fill_2 FILLER_30_682 ();
 sg13g2_fill_1 FILLER_30_684 ();
 sg13g2_fill_2 FILLER_30_689 ();
 sg13g2_fill_1 FILLER_30_727 ();
 sg13g2_decap_4 FILLER_30_736 ();
 sg13g2_fill_1 FILLER_30_740 ();
 sg13g2_decap_4 FILLER_30_746 ();
 sg13g2_fill_2 FILLER_30_750 ();
 sg13g2_fill_1 FILLER_30_757 ();
 sg13g2_decap_8 FILLER_30_772 ();
 sg13g2_fill_2 FILLER_30_779 ();
 sg13g2_fill_1 FILLER_30_781 ();
 sg13g2_fill_2 FILLER_30_795 ();
 sg13g2_fill_1 FILLER_30_797 ();
 sg13g2_decap_8 FILLER_30_835 ();
 sg13g2_decap_8 FILLER_30_842 ();
 sg13g2_decap_8 FILLER_30_849 ();
 sg13g2_fill_1 FILLER_30_860 ();
 sg13g2_decap_8 FILLER_30_865 ();
 sg13g2_fill_2 FILLER_30_881 ();
 sg13g2_fill_1 FILLER_30_883 ();
 sg13g2_decap_4 FILLER_30_932 ();
 sg13g2_fill_1 FILLER_30_962 ();
 sg13g2_fill_2 FILLER_30_1017 ();
 sg13g2_fill_2 FILLER_30_1045 ();
 sg13g2_decap_4 FILLER_30_1055 ();
 sg13g2_decap_8 FILLER_30_1069 ();
 sg13g2_decap_8 FILLER_30_1090 ();
 sg13g2_decap_4 FILLER_30_1102 ();
 sg13g2_fill_2 FILLER_30_1135 ();
 sg13g2_fill_1 FILLER_30_1137 ();
 sg13g2_decap_4 FILLER_30_1182 ();
 sg13g2_fill_2 FILLER_30_1224 ();
 sg13g2_fill_1 FILLER_30_1226 ();
 sg13g2_fill_1 FILLER_30_1278 ();
 sg13g2_fill_2 FILLER_30_1290 ();
 sg13g2_fill_1 FILLER_30_1296 ();
 sg13g2_fill_2 FILLER_30_1305 ();
 sg13g2_fill_1 FILLER_30_1376 ();
 sg13g2_decap_8 FILLER_30_1403 ();
 sg13g2_decap_8 FILLER_30_1410 ();
 sg13g2_decap_4 FILLER_30_1417 ();
 sg13g2_fill_1 FILLER_30_1473 ();
 sg13g2_fill_2 FILLER_30_1478 ();
 sg13g2_fill_1 FILLER_30_1485 ();
 sg13g2_decap_8 FILLER_30_1512 ();
 sg13g2_decap_8 FILLER_30_1519 ();
 sg13g2_fill_2 FILLER_30_1526 ();
 sg13g2_fill_2 FILLER_30_1537 ();
 sg13g2_fill_2 FILLER_30_1544 ();
 sg13g2_fill_1 FILLER_30_1546 ();
 sg13g2_decap_8 FILLER_30_1560 ();
 sg13g2_decap_8 FILLER_30_1567 ();
 sg13g2_decap_8 FILLER_30_1574 ();
 sg13g2_decap_8 FILLER_30_1581 ();
 sg13g2_decap_8 FILLER_30_1593 ();
 sg13g2_decap_8 FILLER_30_1604 ();
 sg13g2_decap_4 FILLER_30_1611 ();
 sg13g2_fill_1 FILLER_30_1615 ();
 sg13g2_fill_1 FILLER_30_1620 ();
 sg13g2_decap_4 FILLER_30_1625 ();
 sg13g2_fill_2 FILLER_30_1629 ();
 sg13g2_fill_1 FILLER_30_1636 ();
 sg13g2_decap_8 FILLER_30_1646 ();
 sg13g2_fill_2 FILLER_30_1653 ();
 sg13g2_decap_4 FILLER_30_1660 ();
 sg13g2_fill_2 FILLER_30_1678 ();
 sg13g2_fill_1 FILLER_30_1760 ();
 sg13g2_fill_1 FILLER_30_1799 ();
 sg13g2_decap_4 FILLER_30_1804 ();
 sg13g2_decap_8 FILLER_30_1811 ();
 sg13g2_fill_2 FILLER_30_1818 ();
 sg13g2_fill_1 FILLER_30_1820 ();
 sg13g2_decap_8 FILLER_30_1846 ();
 sg13g2_decap_4 FILLER_30_1853 ();
 sg13g2_fill_2 FILLER_30_1857 ();
 sg13g2_decap_8 FILLER_30_1865 ();
 sg13g2_fill_1 FILLER_30_1872 ();
 sg13g2_decap_8 FILLER_30_1879 ();
 sg13g2_decap_8 FILLER_30_1886 ();
 sg13g2_fill_1 FILLER_30_1893 ();
 sg13g2_decap_8 FILLER_30_1903 ();
 sg13g2_decap_4 FILLER_30_1910 ();
 sg13g2_decap_8 FILLER_30_1922 ();
 sg13g2_fill_1 FILLER_30_1939 ();
 sg13g2_decap_4 FILLER_30_1948 ();
 sg13g2_fill_1 FILLER_30_1952 ();
 sg13g2_fill_2 FILLER_30_1958 ();
 sg13g2_fill_1 FILLER_30_1960 ();
 sg13g2_decap_8 FILLER_30_1971 ();
 sg13g2_decap_8 FILLER_30_1978 ();
 sg13g2_fill_2 FILLER_30_1985 ();
 sg13g2_fill_1 FILLER_30_1987 ();
 sg13g2_fill_1 FILLER_30_2020 ();
 sg13g2_decap_8 FILLER_30_2031 ();
 sg13g2_decap_4 FILLER_30_2038 ();
 sg13g2_fill_2 FILLER_30_2046 ();
 sg13g2_fill_1 FILLER_30_2048 ();
 sg13g2_decap_4 FILLER_30_2054 ();
 sg13g2_fill_2 FILLER_30_2058 ();
 sg13g2_fill_2 FILLER_30_2065 ();
 sg13g2_fill_1 FILLER_30_2067 ();
 sg13g2_fill_1 FILLER_30_2077 ();
 sg13g2_fill_2 FILLER_30_2082 ();
 sg13g2_fill_1 FILLER_30_2084 ();
 sg13g2_decap_8 FILLER_30_2093 ();
 sg13g2_decap_8 FILLER_30_2139 ();
 sg13g2_decap_4 FILLER_30_2146 ();
 sg13g2_decap_8 FILLER_30_2158 ();
 sg13g2_fill_1 FILLER_30_2165 ();
 sg13g2_fill_2 FILLER_30_2192 ();
 sg13g2_fill_1 FILLER_30_2194 ();
 sg13g2_decap_4 FILLER_30_2208 ();
 sg13g2_fill_1 FILLER_30_2212 ();
 sg13g2_decap_8 FILLER_30_2218 ();
 sg13g2_decap_8 FILLER_30_2225 ();
 sg13g2_fill_1 FILLER_30_2232 ();
 sg13g2_fill_1 FILLER_30_2267 ();
 sg13g2_decap_8 FILLER_30_2299 ();
 sg13g2_fill_2 FILLER_30_2306 ();
 sg13g2_fill_1 FILLER_30_2308 ();
 sg13g2_decap_8 FILLER_30_2335 ();
 sg13g2_decap_8 FILLER_30_2342 ();
 sg13g2_decap_8 FILLER_30_2349 ();
 sg13g2_fill_2 FILLER_30_2356 ();
 sg13g2_fill_2 FILLER_30_2363 ();
 sg13g2_fill_1 FILLER_30_2365 ();
 sg13g2_fill_2 FILLER_30_2370 ();
 sg13g2_decap_8 FILLER_30_2378 ();
 sg13g2_decap_8 FILLER_30_2385 ();
 sg13g2_fill_1 FILLER_30_2392 ();
 sg13g2_decap_8 FILLER_30_2398 ();
 sg13g2_fill_2 FILLER_30_2405 ();
 sg13g2_fill_1 FILLER_30_2407 ();
 sg13g2_fill_2 FILLER_30_2413 ();
 sg13g2_fill_1 FILLER_30_2415 ();
 sg13g2_fill_1 FILLER_30_2420 ();
 sg13g2_decap_8 FILLER_30_2426 ();
 sg13g2_decap_8 FILLER_30_2433 ();
 sg13g2_fill_2 FILLER_30_2440 ();
 sg13g2_fill_1 FILLER_30_2442 ();
 sg13g2_decap_4 FILLER_30_2474 ();
 sg13g2_fill_2 FILLER_30_2483 ();
 sg13g2_fill_1 FILLER_30_2485 ();
 sg13g2_fill_1 FILLER_30_2500 ();
 sg13g2_fill_2 FILLER_30_2506 ();
 sg13g2_fill_2 FILLER_30_2534 ();
 sg13g2_decap_8 FILLER_30_2541 ();
 sg13g2_decap_8 FILLER_30_2548 ();
 sg13g2_decap_8 FILLER_30_2555 ();
 sg13g2_decap_8 FILLER_30_2623 ();
 sg13g2_decap_8 FILLER_30_2630 ();
 sg13g2_decap_8 FILLER_30_2637 ();
 sg13g2_decap_8 FILLER_30_2644 ();
 sg13g2_decap_8 FILLER_30_2651 ();
 sg13g2_decap_8 FILLER_30_2658 ();
 sg13g2_decap_4 FILLER_30_2665 ();
 sg13g2_fill_1 FILLER_30_2669 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_14 ();
 sg13g2_fill_1 FILLER_31_16 ();
 sg13g2_decap_8 FILLER_31_46 ();
 sg13g2_fill_2 FILLER_31_53 ();
 sg13g2_decap_8 FILLER_31_66 ();
 sg13g2_decap_8 FILLER_31_73 ();
 sg13g2_decap_8 FILLER_31_80 ();
 sg13g2_decap_8 FILLER_31_87 ();
 sg13g2_decap_8 FILLER_31_94 ();
 sg13g2_fill_1 FILLER_31_101 ();
 sg13g2_fill_1 FILLER_31_107 ();
 sg13g2_decap_8 FILLER_31_117 ();
 sg13g2_decap_8 FILLER_31_124 ();
 sg13g2_fill_2 FILLER_31_131 ();
 sg13g2_fill_1 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_138 ();
 sg13g2_fill_1 FILLER_31_149 ();
 sg13g2_fill_1 FILLER_31_157 ();
 sg13g2_decap_8 FILLER_31_197 ();
 sg13g2_fill_1 FILLER_31_204 ();
 sg13g2_decap_4 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_fill_1 FILLER_31_220 ();
 sg13g2_decap_8 FILLER_31_254 ();
 sg13g2_decap_8 FILLER_31_275 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_fill_1 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_31_335 ();
 sg13g2_decap_8 FILLER_31_341 ();
 sg13g2_decap_4 FILLER_31_348 ();
 sg13g2_fill_2 FILLER_31_352 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_fill_1 FILLER_31_369 ();
 sg13g2_decap_4 FILLER_31_375 ();
 sg13g2_fill_2 FILLER_31_413 ();
 sg13g2_fill_1 FILLER_31_415 ();
 sg13g2_decap_4 FILLER_31_420 ();
 sg13g2_fill_1 FILLER_31_436 ();
 sg13g2_fill_1 FILLER_31_444 ();
 sg13g2_decap_4 FILLER_31_471 ();
 sg13g2_fill_1 FILLER_31_475 ();
 sg13g2_fill_2 FILLER_31_485 ();
 sg13g2_decap_4 FILLER_31_528 ();
 sg13g2_fill_2 FILLER_31_532 ();
 sg13g2_fill_1 FILLER_31_560 ();
 sg13g2_decap_4 FILLER_31_571 ();
 sg13g2_fill_1 FILLER_31_575 ();
 sg13g2_fill_1 FILLER_31_580 ();
 sg13g2_decap_8 FILLER_31_596 ();
 sg13g2_decap_8 FILLER_31_603 ();
 sg13g2_decap_8 FILLER_31_610 ();
 sg13g2_decap_4 FILLER_31_617 ();
 sg13g2_fill_2 FILLER_31_621 ();
 sg13g2_decap_8 FILLER_31_628 ();
 sg13g2_decap_8 FILLER_31_635 ();
 sg13g2_decap_8 FILLER_31_642 ();
 sg13g2_decap_4 FILLER_31_649 ();
 sg13g2_fill_2 FILLER_31_653 ();
 sg13g2_fill_2 FILLER_31_691 ();
 sg13g2_fill_2 FILLER_31_698 ();
 sg13g2_decap_4 FILLER_31_717 ();
 sg13g2_fill_1 FILLER_31_721 ();
 sg13g2_decap_4 FILLER_31_728 ();
 sg13g2_fill_2 FILLER_31_737 ();
 sg13g2_decap_8 FILLER_31_748 ();
 sg13g2_decap_8 FILLER_31_755 ();
 sg13g2_fill_1 FILLER_31_762 ();
 sg13g2_fill_2 FILLER_31_768 ();
 sg13g2_decap_4 FILLER_31_775 ();
 sg13g2_fill_1 FILLER_31_779 ();
 sg13g2_decap_8 FILLER_31_800 ();
 sg13g2_decap_4 FILLER_31_807 ();
 sg13g2_decap_8 FILLER_31_815 ();
 sg13g2_decap_8 FILLER_31_822 ();
 sg13g2_decap_4 FILLER_31_829 ();
 sg13g2_fill_2 FILLER_31_833 ();
 sg13g2_fill_1 FILLER_31_839 ();
 sg13g2_decap_4 FILLER_31_898 ();
 sg13g2_fill_1 FILLER_31_902 ();
 sg13g2_fill_2 FILLER_31_907 ();
 sg13g2_fill_1 FILLER_31_909 ();
 sg13g2_fill_1 FILLER_31_914 ();
 sg13g2_decap_8 FILLER_31_957 ();
 sg13g2_fill_2 FILLER_31_964 ();
 sg13g2_fill_1 FILLER_31_1002 ();
 sg13g2_fill_1 FILLER_31_1012 ();
 sg13g2_fill_1 FILLER_31_1019 ();
 sg13g2_fill_2 FILLER_31_1056 ();
 sg13g2_fill_2 FILLER_31_1067 ();
 sg13g2_decap_4 FILLER_31_1095 ();
 sg13g2_fill_2 FILLER_31_1099 ();
 sg13g2_fill_2 FILLER_31_1105 ();
 sg13g2_fill_1 FILLER_31_1107 ();
 sg13g2_fill_1 FILLER_31_1139 ();
 sg13g2_fill_1 FILLER_31_1170 ();
 sg13g2_fill_2 FILLER_31_1201 ();
 sg13g2_fill_1 FILLER_31_1208 ();
 sg13g2_decap_8 FILLER_31_1213 ();
 sg13g2_fill_2 FILLER_31_1220 ();
 sg13g2_fill_2 FILLER_31_1244 ();
 sg13g2_fill_2 FILLER_31_1272 ();
 sg13g2_fill_1 FILLER_31_1285 ();
 sg13g2_decap_8 FILLER_31_1322 ();
 sg13g2_fill_2 FILLER_31_1329 ();
 sg13g2_fill_2 FILLER_31_1340 ();
 sg13g2_fill_1 FILLER_31_1347 ();
 sg13g2_fill_2 FILLER_31_1353 ();
 sg13g2_fill_1 FILLER_31_1355 ();
 sg13g2_decap_8 FILLER_31_1362 ();
 sg13g2_decap_4 FILLER_31_1375 ();
 sg13g2_decap_8 FILLER_31_1384 ();
 sg13g2_fill_2 FILLER_31_1391 ();
 sg13g2_fill_2 FILLER_31_1398 ();
 sg13g2_fill_2 FILLER_31_1405 ();
 sg13g2_fill_1 FILLER_31_1407 ();
 sg13g2_decap_8 FILLER_31_1413 ();
 sg13g2_decap_4 FILLER_31_1420 ();
 sg13g2_fill_2 FILLER_31_1424 ();
 sg13g2_decap_4 FILLER_31_1443 ();
 sg13g2_decap_8 FILLER_31_1472 ();
 sg13g2_decap_8 FILLER_31_1479 ();
 sg13g2_decap_8 FILLER_31_1486 ();
 sg13g2_decap_8 FILLER_31_1493 ();
 sg13g2_decap_4 FILLER_31_1530 ();
 sg13g2_fill_1 FILLER_31_1534 ();
 sg13g2_decap_4 FILLER_31_1561 ();
 sg13g2_decap_8 FILLER_31_1569 ();
 sg13g2_decap_8 FILLER_31_1576 ();
 sg13g2_fill_1 FILLER_31_1583 ();
 sg13g2_decap_4 FILLER_31_1589 ();
 sg13g2_decap_4 FILLER_31_1599 ();
 sg13g2_fill_2 FILLER_31_1629 ();
 sg13g2_fill_1 FILLER_31_1631 ();
 sg13g2_decap_4 FILLER_31_1637 ();
 sg13g2_fill_1 FILLER_31_1641 ();
 sg13g2_decap_8 FILLER_31_1681 ();
 sg13g2_decap_8 FILLER_31_1696 ();
 sg13g2_fill_2 FILLER_31_1703 ();
 sg13g2_fill_1 FILLER_31_1705 ();
 sg13g2_decap_4 FILLER_31_1712 ();
 sg13g2_fill_2 FILLER_31_1716 ();
 sg13g2_fill_2 FILLER_31_1722 ();
 sg13g2_fill_1 FILLER_31_1724 ();
 sg13g2_fill_1 FILLER_31_1760 ();
 sg13g2_fill_1 FILLER_31_1768 ();
 sg13g2_fill_2 FILLER_31_1779 ();
 sg13g2_decap_8 FILLER_31_1785 ();
 sg13g2_decap_4 FILLER_31_1792 ();
 sg13g2_fill_1 FILLER_31_1796 ();
 sg13g2_fill_2 FILLER_31_1802 ();
 sg13g2_fill_1 FILLER_31_1804 ();
 sg13g2_decap_8 FILLER_31_1818 ();
 sg13g2_decap_4 FILLER_31_1825 ();
 sg13g2_fill_2 FILLER_31_1834 ();
 sg13g2_fill_1 FILLER_31_1849 ();
 sg13g2_fill_1 FILLER_31_1854 ();
 sg13g2_fill_1 FILLER_31_1881 ();
 sg13g2_decap_8 FILLER_31_1886 ();
 sg13g2_decap_8 FILLER_31_1893 ();
 sg13g2_decap_8 FILLER_31_1900 ();
 sg13g2_fill_1 FILLER_31_1907 ();
 sg13g2_fill_1 FILLER_31_1913 ();
 sg13g2_decap_8 FILLER_31_1940 ();
 sg13g2_decap_8 FILLER_31_1947 ();
 sg13g2_decap_8 FILLER_31_1954 ();
 sg13g2_fill_2 FILLER_31_1961 ();
 sg13g2_decap_4 FILLER_31_1968 ();
 sg13g2_fill_1 FILLER_31_1972 ();
 sg13g2_decap_4 FILLER_31_1978 ();
 sg13g2_fill_1 FILLER_31_1982 ();
 sg13g2_decap_8 FILLER_31_1988 ();
 sg13g2_decap_4 FILLER_31_1995 ();
 sg13g2_decap_4 FILLER_31_2022 ();
 sg13g2_fill_2 FILLER_31_2026 ();
 sg13g2_fill_1 FILLER_31_2040 ();
 sg13g2_fill_1 FILLER_31_2045 ();
 sg13g2_fill_1 FILLER_31_2051 ();
 sg13g2_fill_2 FILLER_31_2078 ();
 sg13g2_fill_1 FILLER_31_2080 ();
 sg13g2_fill_1 FILLER_31_2090 ();
 sg13g2_decap_8 FILLER_31_2101 ();
 sg13g2_decap_8 FILLER_31_2108 ();
 sg13g2_fill_2 FILLER_31_2115 ();
 sg13g2_fill_1 FILLER_31_2117 ();
 sg13g2_fill_1 FILLER_31_2124 ();
 sg13g2_fill_1 FILLER_31_2130 ();
 sg13g2_decap_8 FILLER_31_2135 ();
 sg13g2_decap_4 FILLER_31_2142 ();
 sg13g2_fill_2 FILLER_31_2146 ();
 sg13g2_fill_2 FILLER_31_2153 ();
 sg13g2_fill_1 FILLER_31_2155 ();
 sg13g2_fill_2 FILLER_31_2160 ();
 sg13g2_fill_1 FILLER_31_2162 ();
 sg13g2_decap_8 FILLER_31_2169 ();
 sg13g2_fill_2 FILLER_31_2176 ();
 sg13g2_fill_1 FILLER_31_2184 ();
 sg13g2_fill_2 FILLER_31_2191 ();
 sg13g2_fill_1 FILLER_31_2193 ();
 sg13g2_fill_1 FILLER_31_2198 ();
 sg13g2_decap_8 FILLER_31_2204 ();
 sg13g2_decap_8 FILLER_31_2211 ();
 sg13g2_decap_8 FILLER_31_2218 ();
 sg13g2_fill_2 FILLER_31_2225 ();
 sg13g2_fill_2 FILLER_31_2258 ();
 sg13g2_fill_1 FILLER_31_2290 ();
 sg13g2_fill_2 FILLER_31_2297 ();
 sg13g2_fill_1 FILLER_31_2299 ();
 sg13g2_decap_8 FILLER_31_2309 ();
 sg13g2_fill_2 FILLER_31_2316 ();
 sg13g2_decap_4 FILLER_31_2342 ();
 sg13g2_fill_2 FILLER_31_2452 ();
 sg13g2_decap_8 FILLER_31_2458 ();
 sg13g2_decap_8 FILLER_31_2465 ();
 sg13g2_decap_8 FILLER_31_2472 ();
 sg13g2_decap_8 FILLER_31_2479 ();
 sg13g2_decap_4 FILLER_31_2486 ();
 sg13g2_fill_1 FILLER_31_2523 ();
 sg13g2_decap_8 FILLER_31_2537 ();
 sg13g2_fill_2 FILLER_31_2544 ();
 sg13g2_fill_1 FILLER_31_2546 ();
 sg13g2_fill_1 FILLER_31_2557 ();
 sg13g2_decap_4 FILLER_31_2584 ();
 sg13g2_fill_1 FILLER_31_2592 ();
 sg13g2_decap_8 FILLER_31_2603 ();
 sg13g2_decap_8 FILLER_31_2610 ();
 sg13g2_decap_8 FILLER_31_2617 ();
 sg13g2_decap_8 FILLER_31_2624 ();
 sg13g2_decap_8 FILLER_31_2631 ();
 sg13g2_decap_8 FILLER_31_2638 ();
 sg13g2_decap_8 FILLER_31_2645 ();
 sg13g2_decap_8 FILLER_31_2652 ();
 sg13g2_decap_8 FILLER_31_2659 ();
 sg13g2_decap_4 FILLER_31_2666 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_46 ();
 sg13g2_decap_4 FILLER_32_55 ();
 sg13g2_fill_1 FILLER_32_66 ();
 sg13g2_decap_8 FILLER_32_72 ();
 sg13g2_decap_8 FILLER_32_79 ();
 sg13g2_decap_8 FILLER_32_86 ();
 sg13g2_decap_4 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_97 ();
 sg13g2_fill_1 FILLER_32_127 ();
 sg13g2_fill_2 FILLER_32_162 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_fill_2 FILLER_32_191 ();
 sg13g2_decap_8 FILLER_32_198 ();
 sg13g2_decap_8 FILLER_32_205 ();
 sg13g2_decap_8 FILLER_32_212 ();
 sg13g2_decap_8 FILLER_32_219 ();
 sg13g2_decap_4 FILLER_32_229 ();
 sg13g2_fill_2 FILLER_32_233 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_4 FILLER_32_273 ();
 sg13g2_fill_1 FILLER_32_277 ();
 sg13g2_decap_4 FILLER_32_319 ();
 sg13g2_decap_4 FILLER_32_329 ();
 sg13g2_fill_1 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_346 ();
 sg13g2_decap_8 FILLER_32_353 ();
 sg13g2_decap_4 FILLER_32_360 ();
 sg13g2_fill_2 FILLER_32_364 ();
 sg13g2_decap_4 FILLER_32_371 ();
 sg13g2_fill_2 FILLER_32_375 ();
 sg13g2_fill_2 FILLER_32_387 ();
 sg13g2_decap_4 FILLER_32_397 ();
 sg13g2_fill_1 FILLER_32_401 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_fill_1 FILLER_32_409 ();
 sg13g2_decap_8 FILLER_32_414 ();
 sg13g2_decap_8 FILLER_32_421 ();
 sg13g2_decap_8 FILLER_32_428 ();
 sg13g2_decap_4 FILLER_32_435 ();
 sg13g2_fill_1 FILLER_32_439 ();
 sg13g2_decap_8 FILLER_32_459 ();
 sg13g2_decap_4 FILLER_32_466 ();
 sg13g2_decap_8 FILLER_32_478 ();
 sg13g2_decap_4 FILLER_32_485 ();
 sg13g2_decap_8 FILLER_32_534 ();
 sg13g2_decap_8 FILLER_32_541 ();
 sg13g2_fill_2 FILLER_32_548 ();
 sg13g2_fill_1 FILLER_32_550 ();
 sg13g2_fill_2 FILLER_32_570 ();
 sg13g2_fill_2 FILLER_32_582 ();
 sg13g2_fill_1 FILLER_32_584 ();
 sg13g2_decap_4 FILLER_32_625 ();
 sg13g2_decap_8 FILLER_32_634 ();
 sg13g2_decap_4 FILLER_32_641 ();
 sg13g2_fill_2 FILLER_32_645 ();
 sg13g2_fill_1 FILLER_32_659 ();
 sg13g2_fill_1 FILLER_32_668 ();
 sg13g2_fill_1 FILLER_32_706 ();
 sg13g2_fill_1 FILLER_32_712 ();
 sg13g2_decap_4 FILLER_32_722 ();
 sg13g2_fill_2 FILLER_32_726 ();
 sg13g2_fill_1 FILLER_32_736 ();
 sg13g2_decap_4 FILLER_32_742 ();
 sg13g2_fill_2 FILLER_32_758 ();
 sg13g2_fill_2 FILLER_32_786 ();
 sg13g2_decap_8 FILLER_32_793 ();
 sg13g2_fill_1 FILLER_32_800 ();
 sg13g2_decap_8 FILLER_32_821 ();
 sg13g2_decap_8 FILLER_32_828 ();
 sg13g2_fill_2 FILLER_32_835 ();
 sg13g2_fill_1 FILLER_32_837 ();
 sg13g2_decap_4 FILLER_32_842 ();
 sg13g2_fill_2 FILLER_32_846 ();
 sg13g2_fill_2 FILLER_32_852 ();
 sg13g2_fill_2 FILLER_32_880 ();
 sg13g2_fill_1 FILLER_32_882 ();
 sg13g2_decap_8 FILLER_32_900 ();
 sg13g2_decap_8 FILLER_32_907 ();
 sg13g2_decap_8 FILLER_32_914 ();
 sg13g2_fill_1 FILLER_32_921 ();
 sg13g2_fill_2 FILLER_32_926 ();
 sg13g2_fill_1 FILLER_32_928 ();
 sg13g2_decap_8 FILLER_32_942 ();
 sg13g2_fill_2 FILLER_32_949 ();
 sg13g2_fill_1 FILLER_32_951 ();
 sg13g2_fill_2 FILLER_32_982 ();
 sg13g2_fill_1 FILLER_32_984 ();
 sg13g2_decap_8 FILLER_32_990 ();
 sg13g2_fill_2 FILLER_32_997 ();
 sg13g2_fill_1 FILLER_32_999 ();
 sg13g2_fill_2 FILLER_32_1036 ();
 sg13g2_fill_1 FILLER_32_1043 ();
 sg13g2_fill_2 FILLER_32_1048 ();
 sg13g2_fill_1 FILLER_32_1050 ();
 sg13g2_fill_2 FILLER_32_1055 ();
 sg13g2_decap_4 FILLER_32_1089 ();
 sg13g2_fill_2 FILLER_32_1093 ();
 sg13g2_fill_2 FILLER_32_1101 ();
 sg13g2_fill_1 FILLER_32_1103 ();
 sg13g2_decap_8 FILLER_32_1109 ();
 sg13g2_decap_4 FILLER_32_1116 ();
 sg13g2_decap_8 FILLER_32_1124 ();
 sg13g2_fill_2 FILLER_32_1131 ();
 sg13g2_fill_2 FILLER_32_1179 ();
 sg13g2_fill_1 FILLER_32_1181 ();
 sg13g2_fill_2 FILLER_32_1213 ();
 sg13g2_fill_1 FILLER_32_1215 ();
 sg13g2_fill_1 FILLER_32_1242 ();
 sg13g2_fill_2 FILLER_32_1251 ();
 sg13g2_fill_1 FILLER_32_1253 ();
 sg13g2_decap_8 FILLER_32_1293 ();
 sg13g2_decap_8 FILLER_32_1300 ();
 sg13g2_decap_4 FILLER_32_1307 ();
 sg13g2_fill_1 FILLER_32_1337 ();
 sg13g2_decap_4 FILLER_32_1342 ();
 sg13g2_decap_8 FILLER_32_1359 ();
 sg13g2_decap_4 FILLER_32_1366 ();
 sg13g2_fill_2 FILLER_32_1370 ();
 sg13g2_decap_8 FILLER_32_1378 ();
 sg13g2_fill_2 FILLER_32_1385 ();
 sg13g2_fill_1 FILLER_32_1387 ();
 sg13g2_decap_4 FILLER_32_1392 ();
 sg13g2_fill_1 FILLER_32_1396 ();
 sg13g2_decap_8 FILLER_32_1428 ();
 sg13g2_decap_8 FILLER_32_1435 ();
 sg13g2_decap_8 FILLER_32_1442 ();
 sg13g2_decap_8 FILLER_32_1449 ();
 sg13g2_decap_4 FILLER_32_1456 ();
 sg13g2_fill_2 FILLER_32_1460 ();
 sg13g2_fill_1 FILLER_32_1466 ();
 sg13g2_decap_8 FILLER_32_1478 ();
 sg13g2_decap_8 FILLER_32_1485 ();
 sg13g2_fill_1 FILLER_32_1492 ();
 sg13g2_fill_1 FILLER_32_1509 ();
 sg13g2_fill_1 FILLER_32_1523 ();
 sg13g2_decap_8 FILLER_32_1532 ();
 sg13g2_fill_2 FILLER_32_1539 ();
 sg13g2_fill_1 FILLER_32_1541 ();
 sg13g2_decap_4 FILLER_32_1568 ();
 sg13g2_fill_2 FILLER_32_1572 ();
 sg13g2_decap_8 FILLER_32_1604 ();
 sg13g2_decap_4 FILLER_32_1625 ();
 sg13g2_fill_2 FILLER_32_1629 ();
 sg13g2_decap_8 FILLER_32_1661 ();
 sg13g2_decap_8 FILLER_32_1668 ();
 sg13g2_fill_2 FILLER_32_1675 ();
 sg13g2_fill_1 FILLER_32_1677 ();
 sg13g2_decap_4 FILLER_32_1758 ();
 sg13g2_fill_2 FILLER_32_1762 ();
 sg13g2_fill_1 FILLER_32_1781 ();
 sg13g2_decap_4 FILLER_32_1792 ();
 sg13g2_fill_1 FILLER_32_1800 ();
 sg13g2_decap_8 FILLER_32_1805 ();
 sg13g2_fill_1 FILLER_32_1812 ();
 sg13g2_decap_4 FILLER_32_1839 ();
 sg13g2_fill_2 FILLER_32_1843 ();
 sg13g2_fill_2 FILLER_32_1869 ();
 sg13g2_fill_2 FILLER_32_1875 ();
 sg13g2_fill_1 FILLER_32_1881 ();
 sg13g2_decap_8 FILLER_32_1910 ();
 sg13g2_fill_2 FILLER_32_1922 ();
 sg13g2_fill_1 FILLER_32_1924 ();
 sg13g2_decap_4 FILLER_32_1929 ();
 sg13g2_fill_2 FILLER_32_1946 ();
 sg13g2_decap_4 FILLER_32_1978 ();
 sg13g2_fill_2 FILLER_32_1982 ();
 sg13g2_decap_8 FILLER_32_2020 ();
 sg13g2_decap_8 FILLER_32_2027 ();
 sg13g2_fill_2 FILLER_32_2034 ();
 sg13g2_fill_1 FILLER_32_2073 ();
 sg13g2_fill_1 FILLER_32_2078 ();
 sg13g2_fill_2 FILLER_32_2105 ();
 sg13g2_fill_2 FILLER_32_2112 ();
 sg13g2_fill_1 FILLER_32_2114 ();
 sg13g2_fill_1 FILLER_32_2120 ();
 sg13g2_fill_2 FILLER_32_2147 ();
 sg13g2_fill_1 FILLER_32_2149 ();
 sg13g2_decap_4 FILLER_32_2211 ();
 sg13g2_fill_1 FILLER_32_2215 ();
 sg13g2_fill_1 FILLER_32_2242 ();
 sg13g2_fill_2 FILLER_32_2249 ();
 sg13g2_fill_1 FILLER_32_2275 ();
 sg13g2_fill_1 FILLER_32_2280 ();
 sg13g2_decap_8 FILLER_32_2290 ();
 sg13g2_decap_8 FILLER_32_2297 ();
 sg13g2_decap_4 FILLER_32_2304 ();
 sg13g2_fill_1 FILLER_32_2317 ();
 sg13g2_fill_1 FILLER_32_2356 ();
 sg13g2_decap_8 FILLER_32_2386 ();
 sg13g2_decap_8 FILLER_32_2393 ();
 sg13g2_decap_8 FILLER_32_2400 ();
 sg13g2_fill_1 FILLER_32_2407 ();
 sg13g2_fill_2 FILLER_32_2413 ();
 sg13g2_fill_1 FILLER_32_2415 ();
 sg13g2_fill_1 FILLER_32_2431 ();
 sg13g2_fill_1 FILLER_32_2449 ();
 sg13g2_fill_1 FILLER_32_2455 ();
 sg13g2_fill_1 FILLER_32_2462 ();
 sg13g2_fill_1 FILLER_32_2467 ();
 sg13g2_fill_1 FILLER_32_2473 ();
 sg13g2_fill_2 FILLER_32_2548 ();
 sg13g2_fill_1 FILLER_32_2550 ();
 sg13g2_fill_1 FILLER_32_2577 ();
 sg13g2_decap_4 FILLER_32_2583 ();
 sg13g2_fill_1 FILLER_32_2587 ();
 sg13g2_decap_8 FILLER_32_2593 ();
 sg13g2_decap_8 FILLER_32_2600 ();
 sg13g2_decap_8 FILLER_32_2607 ();
 sg13g2_decap_8 FILLER_32_2614 ();
 sg13g2_decap_8 FILLER_32_2621 ();
 sg13g2_decap_8 FILLER_32_2628 ();
 sg13g2_decap_8 FILLER_32_2635 ();
 sg13g2_decap_8 FILLER_32_2642 ();
 sg13g2_decap_8 FILLER_32_2649 ();
 sg13g2_decap_8 FILLER_32_2656 ();
 sg13g2_decap_8 FILLER_32_2663 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_35 ();
 sg13g2_decap_4 FILLER_33_49 ();
 sg13g2_decap_4 FILLER_33_76 ();
 sg13g2_fill_2 FILLER_33_80 ();
 sg13g2_decap_4 FILLER_33_87 ();
 sg13g2_decap_8 FILLER_33_125 ();
 sg13g2_fill_2 FILLER_33_132 ();
 sg13g2_fill_1 FILLER_33_134 ();
 sg13g2_fill_2 FILLER_33_161 ();
 sg13g2_fill_1 FILLER_33_163 ();
 sg13g2_decap_4 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_181 ();
 sg13g2_fill_1 FILLER_33_195 ();
 sg13g2_decap_8 FILLER_33_205 ();
 sg13g2_decap_4 FILLER_33_212 ();
 sg13g2_fill_1 FILLER_33_216 ();
 sg13g2_decap_8 FILLER_33_222 ();
 sg13g2_decap_8 FILLER_33_229 ();
 sg13g2_decap_4 FILLER_33_236 ();
 sg13g2_fill_2 FILLER_33_243 ();
 sg13g2_decap_4 FILLER_33_252 ();
 sg13g2_fill_1 FILLER_33_256 ();
 sg13g2_fill_2 FILLER_33_266 ();
 sg13g2_decap_4 FILLER_33_273 ();
 sg13g2_fill_2 FILLER_33_277 ();
 sg13g2_decap_8 FILLER_33_317 ();
 sg13g2_decap_8 FILLER_33_324 ();
 sg13g2_decap_4 FILLER_33_331 ();
 sg13g2_decap_4 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_4 FILLER_33_409 ();
 sg13g2_decap_8 FILLER_33_418 ();
 sg13g2_decap_4 FILLER_33_425 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_4 FILLER_33_482 ();
 sg13g2_fill_2 FILLER_33_508 ();
 sg13g2_fill_1 FILLER_33_510 ();
 sg13g2_decap_8 FILLER_33_516 ();
 sg13g2_decap_8 FILLER_33_523 ();
 sg13g2_decap_8 FILLER_33_530 ();
 sg13g2_decap_8 FILLER_33_537 ();
 sg13g2_decap_8 FILLER_33_544 ();
 sg13g2_decap_8 FILLER_33_551 ();
 sg13g2_fill_2 FILLER_33_558 ();
 sg13g2_fill_1 FILLER_33_560 ();
 sg13g2_fill_2 FILLER_33_564 ();
 sg13g2_fill_1 FILLER_33_566 ();
 sg13g2_decap_8 FILLER_33_577 ();
 sg13g2_decap_8 FILLER_33_584 ();
 sg13g2_decap_8 FILLER_33_591 ();
 sg13g2_decap_8 FILLER_33_598 ();
 sg13g2_decap_8 FILLER_33_605 ();
 sg13g2_decap_4 FILLER_33_612 ();
 sg13g2_fill_1 FILLER_33_616 ();
 sg13g2_fill_2 FILLER_33_654 ();
 sg13g2_fill_1 FILLER_33_661 ();
 sg13g2_fill_1 FILLER_33_683 ();
 sg13g2_fill_2 FILLER_33_738 ();
 sg13g2_fill_1 FILLER_33_740 ();
 sg13g2_fill_2 FILLER_33_752 ();
 sg13g2_decap_8 FILLER_33_769 ();
 sg13g2_decap_4 FILLER_33_776 ();
 sg13g2_decap_4 FILLER_33_806 ();
 sg13g2_fill_2 FILLER_33_810 ();
 sg13g2_decap_4 FILLER_33_851 ();
 sg13g2_fill_1 FILLER_33_855 ();
 sg13g2_fill_1 FILLER_33_860 ();
 sg13g2_decap_8 FILLER_33_898 ();
 sg13g2_decap_8 FILLER_33_905 ();
 sg13g2_decap_8 FILLER_33_912 ();
 sg13g2_decap_4 FILLER_33_919 ();
 sg13g2_fill_2 FILLER_33_923 ();
 sg13g2_fill_2 FILLER_33_930 ();
 sg13g2_decap_8 FILLER_33_972 ();
 sg13g2_decap_8 FILLER_33_979 ();
 sg13g2_decap_8 FILLER_33_986 ();
 sg13g2_decap_8 FILLER_33_993 ();
 sg13g2_decap_8 FILLER_33_1000 ();
 sg13g2_fill_1 FILLER_33_1007 ();
 sg13g2_decap_4 FILLER_33_1016 ();
 sg13g2_fill_2 FILLER_33_1020 ();
 sg13g2_decap_4 FILLER_33_1048 ();
 sg13g2_decap_8 FILLER_33_1057 ();
 sg13g2_fill_1 FILLER_33_1064 ();
 sg13g2_decap_8 FILLER_33_1096 ();
 sg13g2_fill_2 FILLER_33_1103 ();
 sg13g2_fill_1 FILLER_33_1105 ();
 sg13g2_decap_8 FILLER_33_1111 ();
 sg13g2_fill_2 FILLER_33_1118 ();
 sg13g2_fill_1 FILLER_33_1120 ();
 sg13g2_decap_8 FILLER_33_1126 ();
 sg13g2_decap_8 FILLER_33_1137 ();
 sg13g2_decap_8 FILLER_33_1144 ();
 sg13g2_fill_1 FILLER_33_1151 ();
 sg13g2_fill_1 FILLER_33_1157 ();
 sg13g2_decap_8 FILLER_33_1168 ();
 sg13g2_fill_2 FILLER_33_1175 ();
 sg13g2_decap_8 FILLER_33_1182 ();
 sg13g2_decap_8 FILLER_33_1189 ();
 sg13g2_decap_8 FILLER_33_1196 ();
 sg13g2_decap_8 FILLER_33_1203 ();
 sg13g2_decap_8 FILLER_33_1210 ();
 sg13g2_decap_8 FILLER_33_1217 ();
 sg13g2_decap_4 FILLER_33_1228 ();
 sg13g2_fill_2 FILLER_33_1232 ();
 sg13g2_fill_2 FILLER_33_1259 ();
 sg13g2_fill_2 FILLER_33_1267 ();
 sg13g2_decap_8 FILLER_33_1295 ();
 sg13g2_decap_8 FILLER_33_1302 ();
 sg13g2_decap_4 FILLER_33_1309 ();
 sg13g2_fill_2 FILLER_33_1313 ();
 sg13g2_decap_8 FILLER_33_1319 ();
 sg13g2_decap_4 FILLER_33_1326 ();
 sg13g2_fill_1 FILLER_33_1330 ();
 sg13g2_decap_4 FILLER_33_1340 ();
 sg13g2_decap_8 FILLER_33_1385 ();
 sg13g2_fill_1 FILLER_33_1392 ();
 sg13g2_fill_2 FILLER_33_1423 ();
 sg13g2_fill_1 FILLER_33_1425 ();
 sg13g2_decap_8 FILLER_33_1447 ();
 sg13g2_decap_8 FILLER_33_1454 ();
 sg13g2_fill_2 FILLER_33_1491 ();
 sg13g2_decap_8 FILLER_33_1531 ();
 sg13g2_decap_4 FILLER_33_1538 ();
 sg13g2_fill_1 FILLER_33_1542 ();
 sg13g2_fill_1 FILLER_33_1552 ();
 sg13g2_fill_1 FILLER_33_1558 ();
 sg13g2_fill_2 FILLER_33_1563 ();
 sg13g2_fill_2 FILLER_33_1570 ();
 sg13g2_fill_2 FILLER_33_1576 ();
 sg13g2_decap_8 FILLER_33_1586 ();
 sg13g2_decap_8 FILLER_33_1593 ();
 sg13g2_decap_8 FILLER_33_1600 ();
 sg13g2_decap_4 FILLER_33_1607 ();
 sg13g2_decap_8 FILLER_33_1637 ();
 sg13g2_decap_8 FILLER_33_1644 ();
 sg13g2_decap_4 FILLER_33_1651 ();
 sg13g2_decap_8 FILLER_33_1668 ();
 sg13g2_decap_4 FILLER_33_1675 ();
 sg13g2_fill_2 FILLER_33_1679 ();
 sg13g2_decap_4 FILLER_33_1685 ();
 sg13g2_decap_8 FILLER_33_1693 ();
 sg13g2_decap_8 FILLER_33_1700 ();
 sg13g2_decap_8 FILLER_33_1707 ();
 sg13g2_decap_8 FILLER_33_1714 ();
 sg13g2_decap_4 FILLER_33_1721 ();
 sg13g2_fill_2 FILLER_33_1725 ();
 sg13g2_decap_8 FILLER_33_1731 ();
 sg13g2_decap_4 FILLER_33_1738 ();
 sg13g2_decap_4 FILLER_33_1747 ();
 sg13g2_fill_1 FILLER_33_1787 ();
 sg13g2_decap_8 FILLER_33_1814 ();
 sg13g2_decap_8 FILLER_33_1821 ();
 sg13g2_decap_8 FILLER_33_1828 ();
 sg13g2_fill_2 FILLER_33_1835 ();
 sg13g2_fill_2 FILLER_33_1849 ();
 sg13g2_decap_4 FILLER_33_1856 ();
 sg13g2_fill_1 FILLER_33_1869 ();
 sg13g2_fill_1 FILLER_33_1916 ();
 sg13g2_decap_8 FILLER_33_1954 ();
 sg13g2_decap_8 FILLER_33_1961 ();
 sg13g2_fill_1 FILLER_33_1968 ();
 sg13g2_decap_4 FILLER_33_1974 ();
 sg13g2_fill_1 FILLER_33_1978 ();
 sg13g2_decap_4 FILLER_33_1983 ();
 sg13g2_fill_1 FILLER_33_1987 ();
 sg13g2_fill_1 FILLER_33_2028 ();
 sg13g2_fill_1 FILLER_33_2064 ();
 sg13g2_decap_4 FILLER_33_2071 ();
 sg13g2_fill_1 FILLER_33_2075 ();
 sg13g2_fill_1 FILLER_33_2102 ();
 sg13g2_fill_1 FILLER_33_2108 ();
 sg13g2_fill_1 FILLER_33_2135 ();
 sg13g2_decap_8 FILLER_33_2154 ();
 sg13g2_decap_4 FILLER_33_2161 ();
 sg13g2_decap_8 FILLER_33_2191 ();
 sg13g2_fill_1 FILLER_33_2198 ();
 sg13g2_decap_4 FILLER_33_2205 ();
 sg13g2_decap_8 FILLER_33_2218 ();
 sg13g2_decap_4 FILLER_33_2225 ();
 sg13g2_fill_1 FILLER_33_2229 ();
 sg13g2_decap_4 FILLER_33_2239 ();
 sg13g2_fill_2 FILLER_33_2274 ();
 sg13g2_fill_2 FILLER_33_2279 ();
 sg13g2_fill_1 FILLER_33_2281 ();
 sg13g2_fill_2 FILLER_33_2300 ();
 sg13g2_fill_1 FILLER_33_2302 ();
 sg13g2_decap_8 FILLER_33_2329 ();
 sg13g2_decap_8 FILLER_33_2336 ();
 sg13g2_decap_8 FILLER_33_2343 ();
 sg13g2_decap_8 FILLER_33_2350 ();
 sg13g2_fill_2 FILLER_33_2378 ();
 sg13g2_fill_1 FILLER_33_2380 ();
 sg13g2_fill_2 FILLER_33_2422 ();
 sg13g2_fill_1 FILLER_33_2424 ();
 sg13g2_decap_8 FILLER_33_2465 ();
 sg13g2_decap_8 FILLER_33_2472 ();
 sg13g2_decap_8 FILLER_33_2479 ();
 sg13g2_decap_4 FILLER_33_2508 ();
 sg13g2_decap_8 FILLER_33_2516 ();
 sg13g2_decap_8 FILLER_33_2523 ();
 sg13g2_decap_8 FILLER_33_2530 ();
 sg13g2_decap_8 FILLER_33_2537 ();
 sg13g2_decap_4 FILLER_33_2544 ();
 sg13g2_decap_8 FILLER_33_2565 ();
 sg13g2_decap_8 FILLER_33_2572 ();
 sg13g2_fill_1 FILLER_33_2579 ();
 sg13g2_decap_8 FILLER_33_2584 ();
 sg13g2_decap_8 FILLER_33_2600 ();
 sg13g2_decap_8 FILLER_33_2607 ();
 sg13g2_fill_2 FILLER_33_2614 ();
 sg13g2_decap_8 FILLER_33_2642 ();
 sg13g2_decap_8 FILLER_33_2649 ();
 sg13g2_decap_8 FILLER_33_2656 ();
 sg13g2_decap_8 FILLER_33_2663 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_45 ();
 sg13g2_fill_1 FILLER_34_47 ();
 sg13g2_decap_4 FILLER_34_80 ();
 sg13g2_fill_1 FILLER_34_122 ();
 sg13g2_decap_8 FILLER_34_128 ();
 sg13g2_decap_4 FILLER_34_135 ();
 sg13g2_decap_4 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_166 ();
 sg13g2_fill_2 FILLER_34_173 ();
 sg13g2_fill_1 FILLER_34_175 ();
 sg13g2_fill_1 FILLER_34_181 ();
 sg13g2_fill_2 FILLER_34_213 ();
 sg13g2_fill_2 FILLER_34_241 ();
 sg13g2_fill_1 FILLER_34_243 ();
 sg13g2_decap_4 FILLER_34_249 ();
 sg13g2_fill_2 FILLER_34_265 ();
 sg13g2_fill_1 FILLER_34_267 ();
 sg13g2_decap_4 FILLER_34_273 ();
 sg13g2_fill_2 FILLER_34_277 ();
 sg13g2_decap_8 FILLER_34_284 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_fill_2 FILLER_34_315 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_fill_1 FILLER_34_431 ();
 sg13g2_decap_4 FILLER_34_436 ();
 sg13g2_decap_4 FILLER_34_445 ();
 sg13g2_fill_2 FILLER_34_449 ();
 sg13g2_decap_8 FILLER_34_454 ();
 sg13g2_fill_2 FILLER_34_461 ();
 sg13g2_decap_8 FILLER_34_467 ();
 sg13g2_decap_8 FILLER_34_474 ();
 sg13g2_decap_8 FILLER_34_481 ();
 sg13g2_decap_8 FILLER_34_488 ();
 sg13g2_decap_8 FILLER_34_495 ();
 sg13g2_fill_2 FILLER_34_502 ();
 sg13g2_decap_8 FILLER_34_508 ();
 sg13g2_fill_2 FILLER_34_550 ();
 sg13g2_fill_1 FILLER_34_552 ();
 sg13g2_decap_8 FILLER_34_588 ();
 sg13g2_decap_8 FILLER_34_595 ();
 sg13g2_decap_8 FILLER_34_602 ();
 sg13g2_decap_4 FILLER_34_609 ();
 sg13g2_fill_1 FILLER_34_613 ();
 sg13g2_fill_1 FILLER_34_617 ();
 sg13g2_fill_2 FILLER_34_622 ();
 sg13g2_fill_1 FILLER_34_630 ();
 sg13g2_fill_2 FILLER_34_635 ();
 sg13g2_fill_1 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_661 ();
 sg13g2_decap_8 FILLER_34_668 ();
 sg13g2_fill_2 FILLER_34_675 ();
 sg13g2_fill_1 FILLER_34_677 ();
 sg13g2_decap_8 FILLER_34_681 ();
 sg13g2_decap_8 FILLER_34_688 ();
 sg13g2_decap_8 FILLER_34_695 ();
 sg13g2_fill_1 FILLER_34_702 ();
 sg13g2_fill_1 FILLER_34_720 ();
 sg13g2_fill_2 FILLER_34_729 ();
 sg13g2_fill_2 FILLER_34_735 ();
 sg13g2_fill_1 FILLER_34_737 ();
 sg13g2_fill_2 FILLER_34_743 ();
 sg13g2_fill_1 FILLER_34_745 ();
 sg13g2_decap_8 FILLER_34_756 ();
 sg13g2_fill_1 FILLER_34_763 ();
 sg13g2_fill_2 FILLER_34_775 ();
 sg13g2_decap_4 FILLER_34_782 ();
 sg13g2_fill_2 FILLER_34_812 ();
 sg13g2_decap_8 FILLER_34_848 ();
 sg13g2_decap_4 FILLER_34_855 ();
 sg13g2_fill_1 FILLER_34_859 ();
 sg13g2_decap_8 FILLER_34_898 ();
 sg13g2_decap_8 FILLER_34_905 ();
 sg13g2_decap_8 FILLER_34_912 ();
 sg13g2_decap_8 FILLER_34_919 ();
 sg13g2_decap_4 FILLER_34_926 ();
 sg13g2_fill_1 FILLER_34_930 ();
 sg13g2_fill_2 FILLER_34_948 ();
 sg13g2_decap_4 FILLER_34_980 ();
 sg13g2_fill_1 FILLER_34_984 ();
 sg13g2_decap_8 FILLER_34_999 ();
 sg13g2_decap_8 FILLER_34_1006 ();
 sg13g2_decap_8 FILLER_34_1013 ();
 sg13g2_fill_2 FILLER_34_1020 ();
 sg13g2_fill_1 FILLER_34_1022 ();
 sg13g2_fill_1 FILLER_34_1040 ();
 sg13g2_decap_8 FILLER_34_1046 ();
 sg13g2_fill_2 FILLER_34_1053 ();
 sg13g2_fill_1 FILLER_34_1055 ();
 sg13g2_decap_8 FILLER_34_1060 ();
 sg13g2_decap_8 FILLER_34_1067 ();
 sg13g2_decap_4 FILLER_34_1074 ();
 sg13g2_fill_2 FILLER_34_1078 ();
 sg13g2_decap_8 FILLER_34_1085 ();
 sg13g2_decap_8 FILLER_34_1092 ();
 sg13g2_decap_8 FILLER_34_1111 ();
 sg13g2_fill_2 FILLER_34_1118 ();
 sg13g2_fill_1 FILLER_34_1120 ();
 sg13g2_decap_8 FILLER_34_1147 ();
 sg13g2_decap_8 FILLER_34_1154 ();
 sg13g2_decap_8 FILLER_34_1161 ();
 sg13g2_decap_8 FILLER_34_1172 ();
 sg13g2_decap_8 FILLER_34_1179 ();
 sg13g2_decap_8 FILLER_34_1186 ();
 sg13g2_decap_8 FILLER_34_1193 ();
 sg13g2_fill_2 FILLER_34_1200 ();
 sg13g2_decap_8 FILLER_34_1206 ();
 sg13g2_decap_8 FILLER_34_1213 ();
 sg13g2_decap_8 FILLER_34_1220 ();
 sg13g2_fill_1 FILLER_34_1227 ();
 sg13g2_decap_4 FILLER_34_1259 ();
 sg13g2_fill_2 FILLER_34_1263 ();
 sg13g2_decap_8 FILLER_34_1269 ();
 sg13g2_fill_2 FILLER_34_1280 ();
 sg13g2_fill_1 FILLER_34_1282 ();
 sg13g2_fill_2 FILLER_34_1288 ();
 sg13g2_fill_1 FILLER_34_1290 ();
 sg13g2_decap_8 FILLER_34_1297 ();
 sg13g2_fill_1 FILLER_34_1334 ();
 sg13g2_decap_4 FILLER_34_1340 ();
 sg13g2_decap_8 FILLER_34_1359 ();
 sg13g2_decap_8 FILLER_34_1366 ();
 sg13g2_fill_1 FILLER_34_1373 ();
 sg13g2_fill_2 FILLER_34_1406 ();
 sg13g2_decap_8 FILLER_34_1412 ();
 sg13g2_fill_2 FILLER_34_1453 ();
 sg13g2_decap_4 FILLER_34_1464 ();
 sg13g2_fill_2 FILLER_34_1468 ();
 sg13g2_fill_2 FILLER_34_1474 ();
 sg13g2_fill_1 FILLER_34_1476 ();
 sg13g2_decap_4 FILLER_34_1507 ();
 sg13g2_decap_8 FILLER_34_1515 ();
 sg13g2_decap_4 FILLER_34_1522 ();
 sg13g2_fill_1 FILLER_34_1526 ();
 sg13g2_decap_8 FILLER_34_1553 ();
 sg13g2_fill_2 FILLER_34_1560 ();
 sg13g2_decap_8 FILLER_34_1588 ();
 sg13g2_decap_8 FILLER_34_1595 ();
 sg13g2_decap_8 FILLER_34_1602 ();
 sg13g2_fill_2 FILLER_34_1609 ();
 sg13g2_fill_1 FILLER_34_1611 ();
 sg13g2_decap_8 FILLER_34_1642 ();
 sg13g2_decap_4 FILLER_34_1649 ();
 sg13g2_fill_1 FILLER_34_1653 ();
 sg13g2_fill_1 FILLER_34_1711 ();
 sg13g2_decap_4 FILLER_34_1716 ();
 sg13g2_fill_2 FILLER_34_1725 ();
 sg13g2_fill_1 FILLER_34_1727 ();
 sg13g2_decap_8 FILLER_34_1759 ();
 sg13g2_decap_8 FILLER_34_1766 ();
 sg13g2_fill_2 FILLER_34_1773 ();
 sg13g2_decap_8 FILLER_34_1801 ();
 sg13g2_decap_8 FILLER_34_1808 ();
 sg13g2_decap_8 FILLER_34_1815 ();
 sg13g2_decap_8 FILLER_34_1822 ();
 sg13g2_decap_8 FILLER_34_1829 ();
 sg13g2_decap_8 FILLER_34_1836 ();
 sg13g2_fill_1 FILLER_34_1843 ();
 sg13g2_fill_2 FILLER_34_1866 ();
 sg13g2_fill_1 FILLER_34_1868 ();
 sg13g2_fill_1 FILLER_34_1875 ();
 sg13g2_fill_2 FILLER_34_1941 ();
 sg13g2_fill_1 FILLER_34_1969 ();
 sg13g2_decap_8 FILLER_34_2001 ();
 sg13g2_decap_8 FILLER_34_2008 ();
 sg13g2_decap_8 FILLER_34_2015 ();
 sg13g2_decap_8 FILLER_34_2022 ();
 sg13g2_decap_8 FILLER_34_2029 ();
 sg13g2_decap_4 FILLER_34_2036 ();
 sg13g2_fill_1 FILLER_34_2053 ();
 sg13g2_decap_8 FILLER_34_2059 ();
 sg13g2_decap_8 FILLER_34_2066 ();
 sg13g2_decap_8 FILLER_34_2073 ();
 sg13g2_fill_1 FILLER_34_2080 ();
 sg13g2_decap_8 FILLER_34_2085 ();
 sg13g2_decap_4 FILLER_34_2092 ();
 sg13g2_decap_8 FILLER_34_2100 ();
 sg13g2_decap_8 FILLER_34_2107 ();
 sg13g2_decap_4 FILLER_34_2114 ();
 sg13g2_fill_1 FILLER_34_2118 ();
 sg13g2_decap_8 FILLER_34_2149 ();
 sg13g2_decap_4 FILLER_34_2156 ();
 sg13g2_fill_2 FILLER_34_2160 ();
 sg13g2_decap_8 FILLER_34_2167 ();
 sg13g2_decap_8 FILLER_34_2174 ();
 sg13g2_fill_1 FILLER_34_2181 ();
 sg13g2_decap_8 FILLER_34_2191 ();
 sg13g2_fill_2 FILLER_34_2198 ();
 sg13g2_decap_4 FILLER_34_2204 ();
 sg13g2_fill_1 FILLER_34_2208 ();
 sg13g2_decap_8 FILLER_34_2235 ();
 sg13g2_fill_1 FILLER_34_2250 ();
 sg13g2_decap_8 FILLER_34_2306 ();
 sg13g2_decap_8 FILLER_34_2344 ();
 sg13g2_decap_8 FILLER_34_2351 ();
 sg13g2_decap_8 FILLER_34_2358 ();
 sg13g2_decap_8 FILLER_34_2365 ();
 sg13g2_decap_4 FILLER_34_2372 ();
 sg13g2_fill_2 FILLER_34_2376 ();
 sg13g2_decap_8 FILLER_34_2384 ();
 sg13g2_fill_1 FILLER_34_2391 ();
 sg13g2_decap_8 FILLER_34_2397 ();
 sg13g2_decap_8 FILLER_34_2404 ();
 sg13g2_fill_1 FILLER_34_2411 ();
 sg13g2_fill_2 FILLER_34_2438 ();
 sg13g2_fill_2 FILLER_34_2445 ();
 sg13g2_decap_8 FILLER_34_2479 ();
 sg13g2_decap_8 FILLER_34_2486 ();
 sg13g2_decap_8 FILLER_34_2493 ();
 sg13g2_decap_4 FILLER_34_2500 ();
 sg13g2_fill_2 FILLER_34_2518 ();
 sg13g2_fill_1 FILLER_34_2520 ();
 sg13g2_decap_8 FILLER_34_2547 ();
 sg13g2_decap_4 FILLER_34_2554 ();
 sg13g2_fill_1 FILLER_34_2558 ();
 sg13g2_fill_2 FILLER_34_2590 ();
 sg13g2_fill_1 FILLER_34_2592 ();
 sg13g2_decap_8 FILLER_34_2645 ();
 sg13g2_decap_8 FILLER_34_2652 ();
 sg13g2_decap_8 FILLER_34_2659 ();
 sg13g2_decap_4 FILLER_34_2666 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_46 ();
 sg13g2_fill_1 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_67 ();
 sg13g2_decap_8 FILLER_35_74 ();
 sg13g2_decap_4 FILLER_35_81 ();
 sg13g2_fill_2 FILLER_35_85 ();
 sg13g2_fill_2 FILLER_35_118 ();
 sg13g2_fill_2 FILLER_35_146 ();
 sg13g2_fill_1 FILLER_35_148 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_fill_1 FILLER_35_176 ();
 sg13g2_fill_2 FILLER_35_182 ();
 sg13g2_fill_2 FILLER_35_189 ();
 sg13g2_fill_2 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_230 ();
 sg13g2_decap_4 FILLER_35_237 ();
 sg13g2_fill_1 FILLER_35_241 ();
 sg13g2_decap_8 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_279 ();
 sg13g2_fill_2 FILLER_35_286 ();
 sg13g2_decap_4 FILLER_35_299 ();
 sg13g2_fill_1 FILLER_35_303 ();
 sg13g2_decap_8 FILLER_35_312 ();
 sg13g2_fill_2 FILLER_35_319 ();
 sg13g2_decap_8 FILLER_35_340 ();
 sg13g2_decap_4 FILLER_35_347 ();
 sg13g2_fill_2 FILLER_35_366 ();
 sg13g2_fill_1 FILLER_35_376 ();
 sg13g2_decap_4 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_decap_8 FILLER_35_433 ();
 sg13g2_fill_2 FILLER_35_440 ();
 sg13g2_fill_1 FILLER_35_442 ();
 sg13g2_decap_8 FILLER_35_446 ();
 sg13g2_decap_8 FILLER_35_453 ();
 sg13g2_decap_8 FILLER_35_460 ();
 sg13g2_decap_4 FILLER_35_467 ();
 sg13g2_fill_1 FILLER_35_471 ();
 sg13g2_fill_2 FILLER_35_480 ();
 sg13g2_fill_1 FILLER_35_482 ();
 sg13g2_decap_8 FILLER_35_491 ();
 sg13g2_fill_2 FILLER_35_498 ();
 sg13g2_fill_1 FILLER_35_500 ();
 sg13g2_decap_4 FILLER_35_505 ();
 sg13g2_fill_2 FILLER_35_509 ();
 sg13g2_decap_8 FILLER_35_518 ();
 sg13g2_decap_8 FILLER_35_525 ();
 sg13g2_decap_8 FILLER_35_532 ();
 sg13g2_fill_1 FILLER_35_544 ();
 sg13g2_fill_2 FILLER_35_578 ();
 sg13g2_decap_8 FILLER_35_598 ();
 sg13g2_fill_2 FILLER_35_605 ();
 sg13g2_fill_1 FILLER_35_607 ();
 sg13g2_fill_2 FILLER_35_620 ();
 sg13g2_fill_1 FILLER_35_622 ();
 sg13g2_fill_2 FILLER_35_648 ();
 sg13g2_fill_1 FILLER_35_650 ();
 sg13g2_decap_8 FILLER_35_672 ();
 sg13g2_decap_4 FILLER_35_679 ();
 sg13g2_fill_2 FILLER_35_687 ();
 sg13g2_fill_1 FILLER_35_699 ();
 sg13g2_fill_2 FILLER_35_709 ();
 sg13g2_fill_2 FILLER_35_715 ();
 sg13g2_fill_1 FILLER_35_717 ();
 sg13g2_fill_2 FILLER_35_725 ();
 sg13g2_fill_1 FILLER_35_727 ();
 sg13g2_fill_2 FILLER_35_736 ();
 sg13g2_fill_1 FILLER_35_738 ();
 sg13g2_fill_1 FILLER_35_746 ();
 sg13g2_fill_2 FILLER_35_755 ();
 sg13g2_decap_8 FILLER_35_792 ();
 sg13g2_decap_8 FILLER_35_799 ();
 sg13g2_decap_8 FILLER_35_811 ();
 sg13g2_fill_2 FILLER_35_818 ();
 sg13g2_decap_4 FILLER_35_828 ();
 sg13g2_fill_1 FILLER_35_836 ();
 sg13g2_decap_4 FILLER_35_863 ();
 sg13g2_fill_2 FILLER_35_867 ();
 sg13g2_fill_2 FILLER_35_878 ();
 sg13g2_decap_8 FILLER_35_883 ();
 sg13g2_decap_4 FILLER_35_890 ();
 sg13g2_fill_2 FILLER_35_924 ();
 sg13g2_fill_1 FILLER_35_956 ();
 sg13g2_decap_8 FILLER_35_1006 ();
 sg13g2_fill_1 FILLER_35_1013 ();
 sg13g2_fill_2 FILLER_35_1018 ();
 sg13g2_fill_1 FILLER_35_1020 ();
 sg13g2_fill_2 FILLER_35_1051 ();
 sg13g2_decap_8 FILLER_35_1067 ();
 sg13g2_fill_2 FILLER_35_1074 ();
 sg13g2_fill_2 FILLER_35_1088 ();
 sg13g2_fill_1 FILLER_35_1098 ();
 sg13g2_fill_1 FILLER_35_1108 ();
 sg13g2_decap_8 FILLER_35_1116 ();
 sg13g2_fill_2 FILLER_35_1123 ();
 sg13g2_fill_1 FILLER_35_1125 ();
 sg13g2_decap_8 FILLER_35_1130 ();
 sg13g2_decap_8 FILLER_35_1137 ();
 sg13g2_decap_8 FILLER_35_1149 ();
 sg13g2_fill_1 FILLER_35_1156 ();
 sg13g2_fill_1 FILLER_35_1167 ();
 sg13g2_decap_8 FILLER_35_1178 ();
 sg13g2_decap_8 FILLER_35_1185 ();
 sg13g2_fill_2 FILLER_35_1192 ();
 sg13g2_fill_1 FILLER_35_1194 ();
 sg13g2_decap_4 FILLER_35_1221 ();
 sg13g2_fill_1 FILLER_35_1225 ();
 sg13g2_fill_1 FILLER_35_1231 ();
 sg13g2_decap_8 FILLER_35_1236 ();
 sg13g2_decap_8 FILLER_35_1243 ();
 sg13g2_decap_8 FILLER_35_1250 ();
 sg13g2_decap_8 FILLER_35_1257 ();
 sg13g2_decap_8 FILLER_35_1264 ();
 sg13g2_decap_8 FILLER_35_1271 ();
 sg13g2_decap_4 FILLER_35_1278 ();
 sg13g2_fill_1 FILLER_35_1282 ();
 sg13g2_decap_4 FILLER_35_1313 ();
 sg13g2_fill_2 FILLER_35_1317 ();
 sg13g2_fill_2 FILLER_35_1327 ();
 sg13g2_fill_1 FILLER_35_1333 ();
 sg13g2_fill_2 FILLER_35_1360 ();
 sg13g2_fill_1 FILLER_35_1367 ();
 sg13g2_fill_1 FILLER_35_1374 ();
 sg13g2_fill_1 FILLER_35_1380 ();
 sg13g2_fill_1 FILLER_35_1395 ();
 sg13g2_decap_4 FILLER_35_1420 ();
 sg13g2_fill_1 FILLER_35_1424 ();
 sg13g2_decap_8 FILLER_35_1431 ();
 sg13g2_fill_1 FILLER_35_1438 ();
 sg13g2_fill_1 FILLER_35_1449 ();
 sg13g2_fill_2 FILLER_35_1484 ();
 sg13g2_fill_1 FILLER_35_1496 ();
 sg13g2_decap_8 FILLER_35_1503 ();
 sg13g2_decap_4 FILLER_35_1510 ();
 sg13g2_fill_2 FILLER_35_1514 ();
 sg13g2_fill_2 FILLER_35_1519 ();
 sg13g2_fill_1 FILLER_35_1521 ();
 sg13g2_fill_1 FILLER_35_1533 ();
 sg13g2_fill_1 FILLER_35_1544 ();
 sg13g2_decap_8 FILLER_35_1549 ();
 sg13g2_decap_8 FILLER_35_1556 ();
 sg13g2_decap_4 FILLER_35_1563 ();
 sg13g2_decap_4 FILLER_35_1576 ();
 sg13g2_fill_2 FILLER_35_1580 ();
 sg13g2_fill_1 FILLER_35_1586 ();
 sg13g2_decap_8 FILLER_35_1600 ();
 sg13g2_fill_2 FILLER_35_1607 ();
 sg13g2_fill_2 FILLER_35_1622 ();
 sg13g2_decap_8 FILLER_35_1628 ();
 sg13g2_fill_2 FILLER_35_1635 ();
 sg13g2_decap_8 FILLER_35_1645 ();
 sg13g2_decap_8 FILLER_35_1652 ();
 sg13g2_decap_8 FILLER_35_1659 ();
 sg13g2_decap_8 FILLER_35_1666 ();
 sg13g2_fill_1 FILLER_35_1673 ();
 sg13g2_decap_4 FILLER_35_1687 ();
 sg13g2_fill_2 FILLER_35_1694 ();
 sg13g2_decap_4 FILLER_35_1730 ();
 sg13g2_fill_2 FILLER_35_1788 ();
 sg13g2_fill_1 FILLER_35_1790 ();
 sg13g2_decap_4 FILLER_35_1795 ();
 sg13g2_fill_2 FILLER_35_1799 ();
 sg13g2_fill_1 FILLER_35_1876 ();
 sg13g2_fill_1 FILLER_35_1886 ();
 sg13g2_fill_2 FILLER_35_1892 ();
 sg13g2_decap_8 FILLER_35_1938 ();
 sg13g2_fill_1 FILLER_35_1950 ();
 sg13g2_fill_2 FILLER_35_1955 ();
 sg13g2_fill_1 FILLER_35_1957 ();
 sg13g2_decap_4 FILLER_35_1963 ();
 sg13g2_fill_2 FILLER_35_1967 ();
 sg13g2_decap_8 FILLER_35_2004 ();
 sg13g2_fill_2 FILLER_35_2011 ();
 sg13g2_fill_1 FILLER_35_2013 ();
 sg13g2_decap_8 FILLER_35_2019 ();
 sg13g2_decap_8 FILLER_35_2026 ();
 sg13g2_decap_8 FILLER_35_2033 ();
 sg13g2_fill_2 FILLER_35_2040 ();
 sg13g2_fill_1 FILLER_35_2042 ();
 sg13g2_decap_8 FILLER_35_2054 ();
 sg13g2_decap_8 FILLER_35_2061 ();
 sg13g2_decap_8 FILLER_35_2068 ();
 sg13g2_decap_4 FILLER_35_2075 ();
 sg13g2_decap_4 FILLER_35_2084 ();
 sg13g2_fill_2 FILLER_35_2088 ();
 sg13g2_decap_4 FILLER_35_2094 ();
 sg13g2_decap_8 FILLER_35_2102 ();
 sg13g2_decap_4 FILLER_35_2109 ();
 sg13g2_fill_2 FILLER_35_2113 ();
 sg13g2_decap_4 FILLER_35_2128 ();
 sg13g2_fill_1 FILLER_35_2132 ();
 sg13g2_decap_4 FILLER_35_2142 ();
 sg13g2_fill_2 FILLER_35_2146 ();
 sg13g2_decap_8 FILLER_35_2158 ();
 sg13g2_decap_8 FILLER_35_2165 ();
 sg13g2_decap_8 FILLER_35_2172 ();
 sg13g2_decap_4 FILLER_35_2179 ();
 sg13g2_fill_2 FILLER_35_2183 ();
 sg13g2_decap_8 FILLER_35_2216 ();
 sg13g2_fill_2 FILLER_35_2223 ();
 sg13g2_fill_1 FILLER_35_2225 ();
 sg13g2_decap_8 FILLER_35_2230 ();
 sg13g2_decap_8 FILLER_35_2279 ();
 sg13g2_decap_4 FILLER_35_2286 ();
 sg13g2_fill_2 FILLER_35_2290 ();
 sg13g2_decap_8 FILLER_35_2319 ();
 sg13g2_decap_8 FILLER_35_2326 ();
 sg13g2_decap_8 FILLER_35_2333 ();
 sg13g2_fill_2 FILLER_35_2340 ();
 sg13g2_fill_1 FILLER_35_2342 ();
 sg13g2_decap_4 FILLER_35_2352 ();
 sg13g2_decap_8 FILLER_35_2404 ();
 sg13g2_decap_4 FILLER_35_2411 ();
 sg13g2_fill_1 FILLER_35_2415 ();
 sg13g2_decap_8 FILLER_35_2425 ();
 sg13g2_decap_4 FILLER_35_2432 ();
 sg13g2_fill_2 FILLER_35_2442 ();
 sg13g2_decap_4 FILLER_35_2479 ();
 sg13g2_fill_1 FILLER_35_2483 ();
 sg13g2_decap_8 FILLER_35_2489 ();
 sg13g2_decap_4 FILLER_35_2496 ();
 sg13g2_fill_1 FILLER_35_2500 ();
 sg13g2_decap_8 FILLER_35_2517 ();
 sg13g2_fill_2 FILLER_35_2534 ();
 sg13g2_fill_1 FILLER_35_2541 ();
 sg13g2_fill_1 FILLER_35_2568 ();
 sg13g2_fill_1 FILLER_35_2575 ();
 sg13g2_fill_1 FILLER_35_2581 ();
 sg13g2_fill_2 FILLER_35_2586 ();
 sg13g2_fill_1 FILLER_35_2614 ();
 sg13g2_fill_1 FILLER_35_2619 ();
 sg13g2_fill_1 FILLER_35_2624 ();
 sg13g2_fill_1 FILLER_35_2629 ();
 sg13g2_decap_8 FILLER_35_2634 ();
 sg13g2_decap_8 FILLER_35_2641 ();
 sg13g2_decap_8 FILLER_35_2648 ();
 sg13g2_decap_8 FILLER_35_2655 ();
 sg13g2_decap_8 FILLER_35_2662 ();
 sg13g2_fill_1 FILLER_35_2669 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_9 ();
 sg13g2_decap_4 FILLER_36_39 ();
 sg13g2_fill_1 FILLER_36_43 ();
 sg13g2_fill_1 FILLER_36_52 ();
 sg13g2_fill_2 FILLER_36_58 ();
 sg13g2_decap_8 FILLER_36_64 ();
 sg13g2_decap_8 FILLER_36_71 ();
 sg13g2_decap_8 FILLER_36_78 ();
 sg13g2_decap_8 FILLER_36_85 ();
 sg13g2_decap_8 FILLER_36_92 ();
 sg13g2_decap_8 FILLER_36_99 ();
 sg13g2_decap_8 FILLER_36_106 ();
 sg13g2_fill_1 FILLER_36_113 ();
 sg13g2_decap_8 FILLER_36_118 ();
 sg13g2_fill_2 FILLER_36_125 ();
 sg13g2_decap_4 FILLER_36_131 ();
 sg13g2_fill_2 FILLER_36_135 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_decap_8 FILLER_36_171 ();
 sg13g2_decap_8 FILLER_36_178 ();
 sg13g2_fill_2 FILLER_36_185 ();
 sg13g2_fill_1 FILLER_36_195 ();
 sg13g2_decap_4 FILLER_36_206 ();
 sg13g2_decap_8 FILLER_36_214 ();
 sg13g2_decap_8 FILLER_36_221 ();
 sg13g2_decap_4 FILLER_36_233 ();
 sg13g2_decap_4 FILLER_36_240 ();
 sg13g2_decap_8 FILLER_36_248 ();
 sg13g2_fill_2 FILLER_36_255 ();
 sg13g2_fill_1 FILLER_36_257 ();
 sg13g2_fill_2 FILLER_36_261 ();
 sg13g2_fill_1 FILLER_36_263 ();
 sg13g2_decap_4 FILLER_36_272 ();
 sg13g2_fill_1 FILLER_36_276 ();
 sg13g2_fill_1 FILLER_36_314 ();
 sg13g2_decap_4 FILLER_36_323 ();
 sg13g2_fill_2 FILLER_36_334 ();
 sg13g2_decap_8 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_351 ();
 sg13g2_fill_2 FILLER_36_358 ();
 sg13g2_decap_4 FILLER_36_369 ();
 sg13g2_fill_1 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_8 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_411 ();
 sg13g2_fill_1 FILLER_36_415 ();
 sg13g2_decap_4 FILLER_36_424 ();
 sg13g2_fill_1 FILLER_36_432 ();
 sg13g2_decap_8 FILLER_36_464 ();
 sg13g2_fill_1 FILLER_36_471 ();
 sg13g2_decap_8 FILLER_36_485 ();
 sg13g2_decap_4 FILLER_36_492 ();
 sg13g2_fill_2 FILLER_36_496 ();
 sg13g2_fill_2 FILLER_36_534 ();
 sg13g2_fill_1 FILLER_36_536 ();
 sg13g2_decap_4 FILLER_36_541 ();
 sg13g2_fill_2 FILLER_36_545 ();
 sg13g2_fill_1 FILLER_36_551 ();
 sg13g2_fill_2 FILLER_36_557 ();
 sg13g2_fill_1 FILLER_36_573 ();
 sg13g2_fill_1 FILLER_36_578 ();
 sg13g2_fill_2 FILLER_36_585 ();
 sg13g2_fill_1 FILLER_36_587 ();
 sg13g2_decap_8 FILLER_36_591 ();
 sg13g2_decap_8 FILLER_36_598 ();
 sg13g2_fill_1 FILLER_36_613 ();
 sg13g2_decap_8 FILLER_36_619 ();
 sg13g2_fill_2 FILLER_36_626 ();
 sg13g2_fill_2 FILLER_36_632 ();
 sg13g2_fill_1 FILLER_36_634 ();
 sg13g2_decap_8 FILLER_36_655 ();
 sg13g2_decap_8 FILLER_36_667 ();
 sg13g2_fill_2 FILLER_36_674 ();
 sg13g2_fill_1 FILLER_36_676 ();
 sg13g2_fill_1 FILLER_36_694 ();
 sg13g2_fill_2 FILLER_36_699 ();
 sg13g2_fill_2 FILLER_36_706 ();
 sg13g2_fill_1 FILLER_36_715 ();
 sg13g2_fill_1 FILLER_36_724 ();
 sg13g2_decap_8 FILLER_36_737 ();
 sg13g2_fill_1 FILLER_36_752 ();
 sg13g2_fill_2 FILLER_36_757 ();
 sg13g2_decap_8 FILLER_36_769 ();
 sg13g2_decap_4 FILLER_36_776 ();
 sg13g2_fill_2 FILLER_36_780 ();
 sg13g2_fill_1 FILLER_36_797 ();
 sg13g2_decap_8 FILLER_36_802 ();
 sg13g2_decap_8 FILLER_36_809 ();
 sg13g2_fill_1 FILLER_36_816 ();
 sg13g2_decap_4 FILLER_36_830 ();
 sg13g2_fill_1 FILLER_36_834 ();
 sg13g2_decap_4 FILLER_36_840 ();
 sg13g2_fill_1 FILLER_36_844 ();
 sg13g2_fill_1 FILLER_36_879 ();
 sg13g2_decap_8 FILLER_36_890 ();
 sg13g2_fill_2 FILLER_36_897 ();
 sg13g2_fill_1 FILLER_36_899 ();
 sg13g2_decap_4 FILLER_36_904 ();
 sg13g2_fill_2 FILLER_36_908 ();
 sg13g2_decap_8 FILLER_36_948 ();
 sg13g2_decap_4 FILLER_36_955 ();
 sg13g2_fill_1 FILLER_36_959 ();
 sg13g2_decap_8 FILLER_36_996 ();
 sg13g2_fill_1 FILLER_36_1003 ();
 sg13g2_fill_1 FILLER_36_1012 ();
 sg13g2_fill_1 FILLER_36_1018 ();
 sg13g2_fill_2 FILLER_36_1050 ();
 sg13g2_fill_1 FILLER_36_1058 ();
 sg13g2_fill_2 FILLER_36_1068 ();
 sg13g2_fill_1 FILLER_36_1070 ();
 sg13g2_fill_1 FILLER_36_1135 ();
 sg13g2_decap_4 FILLER_36_1140 ();
 sg13g2_fill_2 FILLER_36_1144 ();
 sg13g2_fill_1 FILLER_36_1172 ();
 sg13g2_fill_1 FILLER_36_1247 ();
 sg13g2_decap_4 FILLER_36_1278 ();
 sg13g2_fill_1 FILLER_36_1282 ();
 sg13g2_decap_8 FILLER_36_1287 ();
 sg13g2_decap_4 FILLER_36_1294 ();
 sg13g2_fill_2 FILLER_36_1298 ();
 sg13g2_decap_4 FILLER_36_1326 ();
 sg13g2_fill_1 FILLER_36_1330 ();
 sg13g2_fill_2 FILLER_36_1391 ();
 sg13g2_fill_1 FILLER_36_1393 ();
 sg13g2_fill_1 FILLER_36_1400 ();
 sg13g2_decap_4 FILLER_36_1430 ();
 sg13g2_fill_1 FILLER_36_1434 ();
 sg13g2_decap_8 FILLER_36_1445 ();
 sg13g2_decap_8 FILLER_36_1478 ();
 sg13g2_decap_8 FILLER_36_1485 ();
 sg13g2_decap_4 FILLER_36_1492 ();
 sg13g2_fill_1 FILLER_36_1496 ();
 sg13g2_decap_8 FILLER_36_1503 ();
 sg13g2_decap_8 FILLER_36_1510 ();
 sg13g2_decap_8 FILLER_36_1517 ();
 sg13g2_decap_8 FILLER_36_1593 ();
 sg13g2_decap_8 FILLER_36_1626 ();
 sg13g2_fill_2 FILLER_36_1633 ();
 sg13g2_fill_1 FILLER_36_1635 ();
 sg13g2_fill_1 FILLER_36_1645 ();
 sg13g2_decap_8 FILLER_36_1672 ();
 sg13g2_decap_4 FILLER_36_1679 ();
 sg13g2_fill_2 FILLER_36_1683 ();
 sg13g2_decap_4 FILLER_36_1702 ();
 sg13g2_fill_1 FILLER_36_1725 ();
 sg13g2_fill_1 FILLER_36_1735 ();
 sg13g2_decap_8 FILLER_36_1762 ();
 sg13g2_decap_8 FILLER_36_1769 ();
 sg13g2_decap_8 FILLER_36_1776 ();
 sg13g2_fill_2 FILLER_36_1783 ();
 sg13g2_fill_1 FILLER_36_1785 ();
 sg13g2_decap_4 FILLER_36_1789 ();
 sg13g2_decap_4 FILLER_36_1801 ();
 sg13g2_fill_2 FILLER_36_1805 ();
 sg13g2_fill_1 FILLER_36_1812 ();
 sg13g2_fill_1 FILLER_36_1839 ();
 sg13g2_fill_2 FILLER_36_1846 ();
 sg13g2_decap_4 FILLER_36_1922 ();
 sg13g2_fill_1 FILLER_36_1934 ();
 sg13g2_fill_1 FILLER_36_1939 ();
 sg13g2_decap_8 FILLER_36_1945 ();
 sg13g2_fill_2 FILLER_36_1952 ();
 sg13g2_fill_2 FILLER_36_2000 ();
 sg13g2_decap_8 FILLER_36_2006 ();
 sg13g2_fill_2 FILLER_36_2013 ();
 sg13g2_fill_1 FILLER_36_2015 ();
 sg13g2_fill_2 FILLER_36_2021 ();
 sg13g2_decap_4 FILLER_36_2032 ();
 sg13g2_fill_2 FILLER_36_2036 ();
 sg13g2_decap_8 FILLER_36_2043 ();
 sg13g2_decap_8 FILLER_36_2050 ();
 sg13g2_fill_2 FILLER_36_2062 ();
 sg13g2_fill_2 FILLER_36_2074 ();
 sg13g2_fill_2 FILLER_36_2106 ();
 sg13g2_decap_4 FILLER_36_2113 ();
 sg13g2_fill_2 FILLER_36_2121 ();
 sg13g2_decap_4 FILLER_36_2136 ();
 sg13g2_decap_8 FILLER_36_2171 ();
 sg13g2_decap_8 FILLER_36_2178 ();
 sg13g2_fill_2 FILLER_36_2185 ();
 sg13g2_fill_1 FILLER_36_2187 ();
 sg13g2_decap_8 FILLER_36_2197 ();
 sg13g2_decap_8 FILLER_36_2204 ();
 sg13g2_fill_1 FILLER_36_2211 ();
 sg13g2_decap_8 FILLER_36_2217 ();
 sg13g2_decap_8 FILLER_36_2224 ();
 sg13g2_fill_2 FILLER_36_2231 ();
 sg13g2_decap_8 FILLER_36_2266 ();
 sg13g2_fill_1 FILLER_36_2273 ();
 sg13g2_decap_8 FILLER_36_2345 ();
 sg13g2_fill_1 FILLER_36_2352 ();
 sg13g2_fill_2 FILLER_36_2364 ();
 sg13g2_decap_8 FILLER_36_2392 ();
 sg13g2_fill_1 FILLER_36_2399 ();
 sg13g2_decap_4 FILLER_36_2431 ();
 sg13g2_fill_2 FILLER_36_2435 ();
 sg13g2_decap_4 FILLER_36_2468 ();
 sg13g2_fill_1 FILLER_36_2472 ();
 sg13g2_decap_8 FILLER_36_2476 ();
 sg13g2_decap_4 FILLER_36_2483 ();
 sg13g2_decap_8 FILLER_36_2492 ();
 sg13g2_decap_4 FILLER_36_2499 ();
 sg13g2_fill_1 FILLER_36_2503 ();
 sg13g2_fill_2 FILLER_36_2559 ();
 sg13g2_fill_1 FILLER_36_2561 ();
 sg13g2_fill_2 FILLER_36_2589 ();
 sg13g2_fill_2 FILLER_36_2596 ();
 sg13g2_fill_1 FILLER_36_2598 ();
 sg13g2_decap_8 FILLER_36_2625 ();
 sg13g2_decap_8 FILLER_36_2632 ();
 sg13g2_decap_8 FILLER_36_2639 ();
 sg13g2_decap_8 FILLER_36_2646 ();
 sg13g2_decap_8 FILLER_36_2653 ();
 sg13g2_decap_8 FILLER_36_2660 ();
 sg13g2_fill_2 FILLER_36_2667 ();
 sg13g2_fill_1 FILLER_36_2669 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_9 ();
 sg13g2_fill_1 FILLER_37_23 ();
 sg13g2_fill_1 FILLER_37_29 ();
 sg13g2_decap_8 FILLER_37_44 ();
 sg13g2_decap_8 FILLER_37_51 ();
 sg13g2_decap_8 FILLER_37_58 ();
 sg13g2_decap_8 FILLER_37_65 ();
 sg13g2_fill_1 FILLER_37_76 ();
 sg13g2_decap_8 FILLER_37_85 ();
 sg13g2_decap_8 FILLER_37_92 ();
 sg13g2_decap_8 FILLER_37_99 ();
 sg13g2_decap_8 FILLER_37_106 ();
 sg13g2_decap_8 FILLER_37_113 ();
 sg13g2_decap_8 FILLER_37_120 ();
 sg13g2_decap_8 FILLER_37_127 ();
 sg13g2_decap_8 FILLER_37_134 ();
 sg13g2_fill_1 FILLER_37_145 ();
 sg13g2_fill_2 FILLER_37_153 ();
 sg13g2_decap_8 FILLER_37_181 ();
 sg13g2_decap_8 FILLER_37_188 ();
 sg13g2_decap_8 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_202 ();
 sg13g2_fill_1 FILLER_37_204 ();
 sg13g2_decap_8 FILLER_37_211 ();
 sg13g2_decap_8 FILLER_37_218 ();
 sg13g2_fill_2 FILLER_37_225 ();
 sg13g2_fill_2 FILLER_37_234 ();
 sg13g2_fill_2 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_244 ();
 sg13g2_decap_8 FILLER_37_253 ();
 sg13g2_decap_8 FILLER_37_260 ();
 sg13g2_fill_2 FILLER_37_267 ();
 sg13g2_decap_4 FILLER_37_276 ();
 sg13g2_fill_1 FILLER_37_301 ();
 sg13g2_fill_1 FILLER_37_307 ();
 sg13g2_decap_4 FILLER_37_315 ();
 sg13g2_fill_1 FILLER_37_319 ();
 sg13g2_fill_1 FILLER_37_352 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_4 FILLER_37_372 ();
 sg13g2_fill_2 FILLER_37_376 ();
 sg13g2_fill_2 FILLER_37_386 ();
 sg13g2_fill_1 FILLER_37_388 ();
 sg13g2_fill_2 FILLER_37_397 ();
 sg13g2_decap_4 FILLER_37_440 ();
 sg13g2_fill_1 FILLER_37_444 ();
 sg13g2_fill_2 FILLER_37_471 ();
 sg13g2_fill_1 FILLER_37_478 ();
 sg13g2_decap_4 FILLER_37_510 ();
 sg13g2_fill_1 FILLER_37_514 ();
 sg13g2_decap_8 FILLER_37_536 ();
 sg13g2_fill_1 FILLER_37_543 ();
 sg13g2_fill_2 FILLER_37_549 ();
 sg13g2_fill_1 FILLER_37_551 ();
 sg13g2_fill_2 FILLER_37_564 ();
 sg13g2_fill_2 FILLER_37_570 ();
 sg13g2_decap_4 FILLER_37_580 ();
 sg13g2_fill_1 FILLER_37_584 ();
 sg13g2_decap_8 FILLER_37_590 ();
 sg13g2_decap_8 FILLER_37_597 ();
 sg13g2_decap_4 FILLER_37_604 ();
 sg13g2_fill_1 FILLER_37_608 ();
 sg13g2_decap_8 FILLER_37_636 ();
 sg13g2_decap_8 FILLER_37_643 ();
 sg13g2_fill_1 FILLER_37_650 ();
 sg13g2_fill_2 FILLER_37_656 ();
 sg13g2_decap_8 FILLER_37_671 ();
 sg13g2_fill_2 FILLER_37_678 ();
 sg13g2_fill_1 FILLER_37_715 ();
 sg13g2_decap_4 FILLER_37_721 ();
 sg13g2_fill_2 FILLER_37_725 ();
 sg13g2_decap_4 FILLER_37_758 ();
 sg13g2_fill_2 FILLER_37_766 ();
 sg13g2_fill_2 FILLER_37_773 ();
 sg13g2_fill_1 FILLER_37_775 ();
 sg13g2_fill_1 FILLER_37_781 ();
 sg13g2_decap_8 FILLER_37_821 ();
 sg13g2_decap_8 FILLER_37_828 ();
 sg13g2_decap_8 FILLER_37_835 ();
 sg13g2_fill_2 FILLER_37_842 ();
 sg13g2_fill_1 FILLER_37_844 ();
 sg13g2_decap_4 FILLER_37_853 ();
 sg13g2_decap_8 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_37_868 ();
 sg13g2_decap_8 FILLER_37_875 ();
 sg13g2_decap_4 FILLER_37_882 ();
 sg13g2_decap_8 FILLER_37_891 ();
 sg13g2_decap_8 FILLER_37_898 ();
 sg13g2_decap_4 FILLER_37_905 ();
 sg13g2_decap_8 FILLER_37_961 ();
 sg13g2_decap_4 FILLER_37_968 ();
 sg13g2_fill_2 FILLER_37_972 ();
 sg13g2_decap_8 FILLER_37_988 ();
 sg13g2_decap_8 FILLER_37_995 ();
 sg13g2_fill_2 FILLER_37_1002 ();
 sg13g2_fill_1 FILLER_37_1004 ();
 sg13g2_decap_8 FILLER_37_1036 ();
 sg13g2_fill_1 FILLER_37_1043 ();
 sg13g2_fill_2 FILLER_37_1053 ();
 sg13g2_fill_1 FILLER_37_1060 ();
 sg13g2_fill_2 FILLER_37_1113 ();
 sg13g2_fill_2 FILLER_37_1144 ();
 sg13g2_fill_2 FILLER_37_1150 ();
 sg13g2_decap_4 FILLER_37_1178 ();
 sg13g2_fill_1 FILLER_37_1182 ();
 sg13g2_fill_1 FILLER_37_1187 ();
 sg13g2_fill_2 FILLER_37_1193 ();
 sg13g2_fill_2 FILLER_37_1209 ();
 sg13g2_fill_1 FILLER_37_1211 ();
 sg13g2_fill_1 FILLER_37_1229 ();
 sg13g2_fill_1 FILLER_37_1235 ();
 sg13g2_decap_8 FILLER_37_1300 ();
 sg13g2_fill_2 FILLER_37_1307 ();
 sg13g2_fill_2 FILLER_37_1335 ();
 sg13g2_decap_8 FILLER_37_1346 ();
 sg13g2_decap_4 FILLER_37_1353 ();
 sg13g2_fill_2 FILLER_37_1357 ();
 sg13g2_fill_1 FILLER_37_1365 ();
 sg13g2_decap_8 FILLER_37_1370 ();
 sg13g2_decap_4 FILLER_37_1377 ();
 sg13g2_fill_2 FILLER_37_1386 ();
 sg13g2_fill_2 FILLER_37_1432 ();
 sg13g2_fill_1 FILLER_37_1434 ();
 sg13g2_fill_2 FILLER_37_1449 ();
 sg13g2_fill_1 FILLER_37_1451 ();
 sg13g2_decap_8 FILLER_37_1456 ();
 sg13g2_decap_8 FILLER_37_1463 ();
 sg13g2_fill_1 FILLER_37_1470 ();
 sg13g2_fill_1 FILLER_37_1501 ();
 sg13g2_decap_8 FILLER_37_1507 ();
 sg13g2_decap_4 FILLER_37_1514 ();
 sg13g2_fill_1 FILLER_37_1518 ();
 sg13g2_decap_4 FILLER_37_1549 ();
 sg13g2_decap_8 FILLER_37_1591 ();
 sg13g2_decap_8 FILLER_37_1598 ();
 sg13g2_fill_2 FILLER_37_1627 ();
 sg13g2_decap_8 FILLER_37_1659 ();
 sg13g2_decap_4 FILLER_37_1666 ();
 sg13g2_fill_1 FILLER_37_1670 ();
 sg13g2_decap_8 FILLER_37_1698 ();
 sg13g2_fill_2 FILLER_37_1710 ();
 sg13g2_fill_1 FILLER_37_1712 ();
 sg13g2_fill_1 FILLER_37_1717 ();
 sg13g2_fill_2 FILLER_37_1748 ();
 sg13g2_fill_1 FILLER_37_1750 ();
 sg13g2_decap_8 FILLER_37_1760 ();
 sg13g2_fill_2 FILLER_37_1767 ();
 sg13g2_decap_4 FILLER_37_1782 ();
 sg13g2_fill_1 FILLER_37_1791 ();
 sg13g2_decap_4 FILLER_37_1810 ();
 sg13g2_fill_1 FILLER_37_1818 ();
 sg13g2_decap_4 FILLER_37_1831 ();
 sg13g2_fill_1 FILLER_37_1835 ();
 sg13g2_fill_2 FILLER_37_1841 ();
 sg13g2_fill_2 FILLER_37_1848 ();
 sg13g2_fill_1 FILLER_37_1850 ();
 sg13g2_fill_1 FILLER_37_1886 ();
 sg13g2_decap_8 FILLER_37_1897 ();
 sg13g2_fill_2 FILLER_37_1904 ();
 sg13g2_fill_2 FILLER_37_1914 ();
 sg13g2_decap_4 FILLER_37_1937 ();
 sg13g2_fill_2 FILLER_37_1941 ();
 sg13g2_decap_8 FILLER_37_1969 ();
 sg13g2_decap_4 FILLER_37_1976 ();
 sg13g2_decap_8 FILLER_37_1988 ();
 sg13g2_fill_1 FILLER_37_1995 ();
 sg13g2_decap_8 FILLER_37_2136 ();
 sg13g2_decap_8 FILLER_37_2143 ();
 sg13g2_decap_8 FILLER_37_2150 ();
 sg13g2_decap_8 FILLER_37_2157 ();
 sg13g2_decap_4 FILLER_37_2164 ();
 sg13g2_fill_2 FILLER_37_2181 ();
 sg13g2_decap_4 FILLER_37_2222 ();
 sg13g2_fill_2 FILLER_37_2226 ();
 sg13g2_fill_1 FILLER_37_2233 ();
 sg13g2_decap_4 FILLER_37_2269 ();
 sg13g2_fill_1 FILLER_37_2273 ();
 sg13g2_decap_4 FILLER_37_2296 ();
 sg13g2_fill_1 FILLER_37_2300 ();
 sg13g2_fill_2 FILLER_37_2310 ();
 sg13g2_decap_4 FILLER_37_2318 ();
 sg13g2_decap_8 FILLER_37_2348 ();
 sg13g2_fill_1 FILLER_37_2355 ();
 sg13g2_fill_2 FILLER_37_2412 ();
 sg13g2_decap_8 FILLER_37_2424 ();
 sg13g2_decap_8 FILLER_37_2431 ();
 sg13g2_fill_2 FILLER_37_2438 ();
 sg13g2_fill_1 FILLER_37_2440 ();
 sg13g2_fill_1 FILLER_37_2476 ();
 sg13g2_fill_2 FILLER_37_2485 ();
 sg13g2_decap_4 FILLER_37_2495 ();
 sg13g2_decap_8 FILLER_37_2507 ();
 sg13g2_decap_4 FILLER_37_2514 ();
 sg13g2_fill_2 FILLER_37_2518 ();
 sg13g2_fill_2 FILLER_37_2549 ();
 sg13g2_decap_8 FILLER_37_2594 ();
 sg13g2_decap_8 FILLER_37_2601 ();
 sg13g2_decap_8 FILLER_37_2608 ();
 sg13g2_decap_8 FILLER_37_2615 ();
 sg13g2_decap_8 FILLER_37_2622 ();
 sg13g2_decap_8 FILLER_37_2629 ();
 sg13g2_decap_8 FILLER_37_2636 ();
 sg13g2_decap_8 FILLER_37_2643 ();
 sg13g2_decap_8 FILLER_37_2650 ();
 sg13g2_decap_8 FILLER_37_2657 ();
 sg13g2_decap_4 FILLER_37_2664 ();
 sg13g2_fill_2 FILLER_37_2668 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_4 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_33 ();
 sg13g2_fill_1 FILLER_38_39 ();
 sg13g2_fill_2 FILLER_38_54 ();
 sg13g2_fill_1 FILLER_38_56 ();
 sg13g2_decap_4 FILLER_38_61 ();
 sg13g2_decap_4 FILLER_38_97 ();
 sg13g2_fill_2 FILLER_38_101 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_fill_2 FILLER_38_154 ();
 sg13g2_fill_2 FILLER_38_170 ();
 sg13g2_fill_1 FILLER_38_172 ();
 sg13g2_fill_1 FILLER_38_207 ();
 sg13g2_decap_4 FILLER_38_258 ();
 sg13g2_fill_1 FILLER_38_262 ();
 sg13g2_fill_2 FILLER_38_366 ();
 sg13g2_decap_4 FILLER_38_397 ();
 sg13g2_fill_1 FILLER_38_401 ();
 sg13g2_decap_4 FILLER_38_407 ();
 sg13g2_fill_2 FILLER_38_411 ();
 sg13g2_decap_4 FILLER_38_422 ();
 sg13g2_fill_1 FILLER_38_426 ();
 sg13g2_decap_4 FILLER_38_435 ();
 sg13g2_fill_1 FILLER_38_439 ();
 sg13g2_fill_1 FILLER_38_444 ();
 sg13g2_decap_8 FILLER_38_509 ();
 sg13g2_decap_8 FILLER_38_516 ();
 sg13g2_decap_8 FILLER_38_523 ();
 sg13g2_decap_4 FILLER_38_530 ();
 sg13g2_decap_8 FILLER_38_569 ();
 sg13g2_decap_8 FILLER_38_576 ();
 sg13g2_decap_8 FILLER_38_583 ();
 sg13g2_decap_4 FILLER_38_590 ();
 sg13g2_fill_2 FILLER_38_594 ();
 sg13g2_decap_8 FILLER_38_601 ();
 sg13g2_decap_4 FILLER_38_608 ();
 sg13g2_fill_1 FILLER_38_612 ();
 sg13g2_decap_4 FILLER_38_638 ();
 sg13g2_fill_1 FILLER_38_647 ();
 sg13g2_decap_8 FILLER_38_669 ();
 sg13g2_fill_2 FILLER_38_676 ();
 sg13g2_fill_1 FILLER_38_678 ();
 sg13g2_fill_1 FILLER_38_703 ();
 sg13g2_decap_8 FILLER_38_714 ();
 sg13g2_decap_8 FILLER_38_721 ();
 sg13g2_fill_1 FILLER_38_728 ();
 sg13g2_fill_2 FILLER_38_740 ();
 sg13g2_fill_1 FILLER_38_764 ();
 sg13g2_fill_1 FILLER_38_774 ();
 sg13g2_fill_2 FILLER_38_801 ();
 sg13g2_decap_8 FILLER_38_816 ();
 sg13g2_decap_8 FILLER_38_823 ();
 sg13g2_decap_8 FILLER_38_830 ();
 sg13g2_decap_4 FILLER_38_837 ();
 sg13g2_fill_2 FILLER_38_841 ();
 sg13g2_decap_8 FILLER_38_869 ();
 sg13g2_decap_8 FILLER_38_876 ();
 sg13g2_decap_4 FILLER_38_883 ();
 sg13g2_decap_8 FILLER_38_913 ();
 sg13g2_decap_8 FILLER_38_920 ();
 sg13g2_decap_4 FILLER_38_927 ();
 sg13g2_decap_8 FILLER_38_983 ();
 sg13g2_decap_4 FILLER_38_990 ();
 sg13g2_fill_1 FILLER_38_994 ();
 sg13g2_decap_4 FILLER_38_1001 ();
 sg13g2_fill_2 FILLER_38_1005 ();
 sg13g2_decap_8 FILLER_38_1015 ();
 sg13g2_decap_8 FILLER_38_1026 ();
 sg13g2_decap_4 FILLER_38_1033 ();
 sg13g2_fill_1 FILLER_38_1037 ();
 sg13g2_fill_2 FILLER_38_1083 ();
 sg13g2_fill_1 FILLER_38_1091 ();
 sg13g2_fill_2 FILLER_38_1104 ();
 sg13g2_fill_1 FILLER_38_1122 ();
 sg13g2_fill_2 FILLER_38_1169 ();
 sg13g2_fill_2 FILLER_38_1177 ();
 sg13g2_fill_1 FILLER_38_1179 ();
 sg13g2_decap_8 FILLER_38_1220 ();
 sg13g2_decap_8 FILLER_38_1227 ();
 sg13g2_decap_8 FILLER_38_1234 ();
 sg13g2_decap_4 FILLER_38_1241 ();
 sg13g2_fill_2 FILLER_38_1245 ();
 sg13g2_decap_4 FILLER_38_1252 ();
 sg13g2_fill_2 FILLER_38_1256 ();
 sg13g2_fill_1 FILLER_38_1262 ();
 sg13g2_fill_2 FILLER_38_1275 ();
 sg13g2_fill_1 FILLER_38_1277 ();
 sg13g2_decap_8 FILLER_38_1283 ();
 sg13g2_fill_2 FILLER_38_1290 ();
 sg13g2_fill_1 FILLER_38_1292 ();
 sg13g2_fill_1 FILLER_38_1297 ();
 sg13g2_fill_1 FILLER_38_1303 ();
 sg13g2_decap_8 FILLER_38_1309 ();
 sg13g2_decap_8 FILLER_38_1329 ();
 sg13g2_decap_4 FILLER_38_1336 ();
 sg13g2_fill_1 FILLER_38_1340 ();
 sg13g2_decap_8 FILLER_38_1350 ();
 sg13g2_decap_8 FILLER_38_1357 ();
 sg13g2_decap_8 FILLER_38_1364 ();
 sg13g2_decap_8 FILLER_38_1371 ();
 sg13g2_fill_2 FILLER_38_1378 ();
 sg13g2_fill_1 FILLER_38_1395 ();
 sg13g2_fill_2 FILLER_38_1401 ();
 sg13g2_fill_1 FILLER_38_1403 ();
 sg13g2_decap_4 FILLER_38_1412 ();
 sg13g2_fill_1 FILLER_38_1416 ();
 sg13g2_decap_4 FILLER_38_1421 ();
 sg13g2_fill_1 FILLER_38_1425 ();
 sg13g2_decap_4 FILLER_38_1430 ();
 sg13g2_decap_8 FILLER_38_1479 ();
 sg13g2_decap_8 FILLER_38_1499 ();
 sg13g2_decap_8 FILLER_38_1506 ();
 sg13g2_fill_2 FILLER_38_1513 ();
 sg13g2_fill_1 FILLER_38_1515 ();
 sg13g2_fill_1 FILLER_38_1555 ();
 sg13g2_fill_1 FILLER_38_1561 ();
 sg13g2_fill_2 FILLER_38_1568 ();
 sg13g2_fill_2 FILLER_38_1591 ();
 sg13g2_fill_1 FILLER_38_1593 ();
 sg13g2_decap_4 FILLER_38_1600 ();
 sg13g2_decap_4 FILLER_38_1635 ();
 sg13g2_fill_2 FILLER_38_1639 ();
 sg13g2_decap_8 FILLER_38_1645 ();
 sg13g2_fill_2 FILLER_38_1652 ();
 sg13g2_fill_1 FILLER_38_1654 ();
 sg13g2_decap_4 FILLER_38_1660 ();
 sg13g2_fill_2 FILLER_38_1664 ();
 sg13g2_fill_2 FILLER_38_1679 ();
 sg13g2_fill_1 FILLER_38_1681 ();
 sg13g2_decap_8 FILLER_38_1712 ();
 sg13g2_decap_8 FILLER_38_1719 ();
 sg13g2_fill_1 FILLER_38_1730 ();
 sg13g2_fill_2 FILLER_38_1742 ();
 sg13g2_fill_1 FILLER_38_1781 ();
 sg13g2_decap_8 FILLER_38_1840 ();
 sg13g2_fill_1 FILLER_38_1847 ();
 sg13g2_fill_1 FILLER_38_1859 ();
 sg13g2_decap_8 FILLER_38_1886 ();
 sg13g2_fill_1 FILLER_38_1893 ();
 sg13g2_fill_2 FILLER_38_1902 ();
 sg13g2_fill_1 FILLER_38_1904 ();
 sg13g2_fill_1 FILLER_38_1918 ();
 sg13g2_decap_8 FILLER_38_1963 ();
 sg13g2_decap_8 FILLER_38_1970 ();
 sg13g2_decap_8 FILLER_38_1977 ();
 sg13g2_decap_8 FILLER_38_1984 ();
 sg13g2_fill_1 FILLER_38_1991 ();
 sg13g2_fill_1 FILLER_38_2032 ();
 sg13g2_decap_8 FILLER_38_2038 ();
 sg13g2_decap_8 FILLER_38_2045 ();
 sg13g2_fill_1 FILLER_38_2052 ();
 sg13g2_decap_4 FILLER_38_2058 ();
 sg13g2_fill_1 FILLER_38_2062 ();
 sg13g2_fill_2 FILLER_38_2067 ();
 sg13g2_fill_1 FILLER_38_2069 ();
 sg13g2_decap_4 FILLER_38_2086 ();
 sg13g2_fill_2 FILLER_38_2090 ();
 sg13g2_fill_2 FILLER_38_2097 ();
 sg13g2_fill_1 FILLER_38_2099 ();
 sg13g2_fill_2 FILLER_38_2106 ();
 sg13g2_fill_1 FILLER_38_2108 ();
 sg13g2_fill_2 FILLER_38_2146 ();
 sg13g2_fill_1 FILLER_38_2148 ();
 sg13g2_decap_4 FILLER_38_2157 ();
 sg13g2_fill_1 FILLER_38_2161 ();
 sg13g2_fill_2 FILLER_38_2188 ();
 sg13g2_fill_1 FILLER_38_2196 ();
 sg13g2_fill_2 FILLER_38_2234 ();
 sg13g2_fill_2 FILLER_38_2252 ();
 sg13g2_decap_4 FILLER_38_2258 ();
 sg13g2_fill_1 FILLER_38_2262 ();
 sg13g2_fill_2 FILLER_38_2301 ();
 sg13g2_decap_8 FILLER_38_2324 ();
 sg13g2_decap_4 FILLER_38_2331 ();
 sg13g2_fill_1 FILLER_38_2335 ();
 sg13g2_decap_8 FILLER_38_2371 ();
 sg13g2_fill_2 FILLER_38_2378 ();
 sg13g2_fill_2 FILLER_38_2392 ();
 sg13g2_fill_1 FILLER_38_2394 ();
 sg13g2_decap_4 FILLER_38_2399 ();
 sg13g2_decap_4 FILLER_38_2407 ();
 sg13g2_decap_8 FILLER_38_2430 ();
 sg13g2_decap_8 FILLER_38_2437 ();
 sg13g2_fill_1 FILLER_38_2444 ();
 sg13g2_decap_4 FILLER_38_2449 ();
 sg13g2_decap_8 FILLER_38_2488 ();
 sg13g2_decap_4 FILLER_38_2495 ();
 sg13g2_decap_8 FILLER_38_2503 ();
 sg13g2_decap_4 FILLER_38_2510 ();
 sg13g2_fill_1 FILLER_38_2514 ();
 sg13g2_decap_8 FILLER_38_2524 ();
 sg13g2_decap_4 FILLER_38_2531 ();
 sg13g2_decap_8 FILLER_38_2544 ();
 sg13g2_decap_8 FILLER_38_2551 ();
 sg13g2_fill_1 FILLER_38_2558 ();
 sg13g2_fill_2 FILLER_38_2564 ();
 sg13g2_fill_1 FILLER_38_2566 ();
 sg13g2_decap_8 FILLER_38_2571 ();
 sg13g2_decap_8 FILLER_38_2578 ();
 sg13g2_decap_8 FILLER_38_2585 ();
 sg13g2_decap_8 FILLER_38_2592 ();
 sg13g2_decap_8 FILLER_38_2599 ();
 sg13g2_decap_8 FILLER_38_2606 ();
 sg13g2_decap_8 FILLER_38_2613 ();
 sg13g2_decap_8 FILLER_38_2620 ();
 sg13g2_decap_8 FILLER_38_2631 ();
 sg13g2_decap_8 FILLER_38_2638 ();
 sg13g2_decap_8 FILLER_38_2645 ();
 sg13g2_decap_8 FILLER_38_2652 ();
 sg13g2_decap_8 FILLER_38_2659 ();
 sg13g2_decap_4 FILLER_38_2666 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_fill_2 FILLER_39_175 ();
 sg13g2_fill_1 FILLER_39_177 ();
 sg13g2_decap_4 FILLER_39_207 ();
 sg13g2_fill_1 FILLER_39_211 ();
 sg13g2_decap_4 FILLER_39_264 ();
 sg13g2_decap_8 FILLER_39_272 ();
 sg13g2_decap_8 FILLER_39_279 ();
 sg13g2_decap_8 FILLER_39_286 ();
 sg13g2_decap_8 FILLER_39_293 ();
 sg13g2_fill_1 FILLER_39_300 ();
 sg13g2_fill_1 FILLER_39_309 ();
 sg13g2_decap_4 FILLER_39_315 ();
 sg13g2_fill_1 FILLER_39_319 ();
 sg13g2_fill_2 FILLER_39_331 ();
 sg13g2_decap_8 FILLER_39_354 ();
 sg13g2_decap_8 FILLER_39_361 ();
 sg13g2_decap_8 FILLER_39_368 ();
 sg13g2_decap_8 FILLER_39_375 ();
 sg13g2_fill_1 FILLER_39_382 ();
 sg13g2_fill_2 FILLER_39_393 ();
 sg13g2_fill_2 FILLER_39_400 ();
 sg13g2_fill_1 FILLER_39_402 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_4 FILLER_39_424 ();
 sg13g2_fill_2 FILLER_39_428 ();
 sg13g2_decap_8 FILLER_39_435 ();
 sg13g2_decap_4 FILLER_39_442 ();
 sg13g2_fill_2 FILLER_39_460 ();
 sg13g2_fill_1 FILLER_39_462 ();
 sg13g2_decap_4 FILLER_39_518 ();
 sg13g2_decap_8 FILLER_39_526 ();
 sg13g2_decap_8 FILLER_39_533 ();
 sg13g2_decap_8 FILLER_39_540 ();
 sg13g2_decap_8 FILLER_39_547 ();
 sg13g2_decap_8 FILLER_39_554 ();
 sg13g2_decap_8 FILLER_39_561 ();
 sg13g2_decap_8 FILLER_39_568 ();
 sg13g2_fill_2 FILLER_39_575 ();
 sg13g2_decap_4 FILLER_39_612 ();
 sg13g2_fill_1 FILLER_39_616 ();
 sg13g2_decap_8 FILLER_39_633 ();
 sg13g2_fill_2 FILLER_39_640 ();
 sg13g2_fill_1 FILLER_39_653 ();
 sg13g2_fill_2 FILLER_39_674 ();
 sg13g2_decap_8 FILLER_39_715 ();
 sg13g2_decap_8 FILLER_39_722 ();
 sg13g2_decap_8 FILLER_39_729 ();
 sg13g2_fill_1 FILLER_39_736 ();
 sg13g2_fill_2 FILLER_39_774 ();
 sg13g2_decap_4 FILLER_39_786 ();
 sg13g2_fill_1 FILLER_39_790 ();
 sg13g2_fill_2 FILLER_39_804 ();
 sg13g2_decap_4 FILLER_39_835 ();
 sg13g2_decap_8 FILLER_39_865 ();
 sg13g2_decap_4 FILLER_39_872 ();
 sg13g2_fill_1 FILLER_39_876 ();
 sg13g2_fill_1 FILLER_39_903 ();
 sg13g2_fill_2 FILLER_39_917 ();
 sg13g2_fill_1 FILLER_39_919 ();
 sg13g2_decap_8 FILLER_39_926 ();
 sg13g2_decap_8 FILLER_39_933 ();
 sg13g2_decap_8 FILLER_39_940 ();
 sg13g2_fill_1 FILLER_39_947 ();
 sg13g2_decap_8 FILLER_39_953 ();
 sg13g2_decap_8 FILLER_39_960 ();
 sg13g2_fill_1 FILLER_39_967 ();
 sg13g2_fill_2 FILLER_39_998 ();
 sg13g2_fill_1 FILLER_39_1000 ();
 sg13g2_fill_1 FILLER_39_1051 ();
 sg13g2_fill_2 FILLER_39_1061 ();
 sg13g2_decap_4 FILLER_39_1076 ();
 sg13g2_fill_2 FILLER_39_1080 ();
 sg13g2_fill_2 FILLER_39_1100 ();
 sg13g2_fill_1 FILLER_39_1118 ();
 sg13g2_fill_2 FILLER_39_1158 ();
 sg13g2_fill_1 FILLER_39_1160 ();
 sg13g2_decap_8 FILLER_39_1192 ();
 sg13g2_decap_8 FILLER_39_1199 ();
 sg13g2_decap_8 FILLER_39_1206 ();
 sg13g2_decap_4 FILLER_39_1213 ();
 sg13g2_fill_1 FILLER_39_1217 ();
 sg13g2_decap_8 FILLER_39_1226 ();
 sg13g2_decap_8 FILLER_39_1233 ();
 sg13g2_decap_8 FILLER_39_1245 ();
 sg13g2_decap_4 FILLER_39_1252 ();
 sg13g2_decap_8 FILLER_39_1260 ();
 sg13g2_decap_8 FILLER_39_1267 ();
 sg13g2_fill_1 FILLER_39_1274 ();
 sg13g2_fill_2 FILLER_39_1280 ();
 sg13g2_fill_1 FILLER_39_1329 ();
 sg13g2_decap_8 FILLER_39_1364 ();
 sg13g2_decap_8 FILLER_39_1371 ();
 sg13g2_decap_4 FILLER_39_1378 ();
 sg13g2_fill_1 FILLER_39_1405 ();
 sg13g2_fill_2 FILLER_39_1412 ();
 sg13g2_fill_2 FILLER_39_1440 ();
 sg13g2_decap_8 FILLER_39_1448 ();
 sg13g2_fill_2 FILLER_39_1485 ();
 sg13g2_fill_2 FILLER_39_1513 ();
 sg13g2_fill_2 FILLER_39_1519 ();
 sg13g2_fill_1 FILLER_39_1521 ();
 sg13g2_decap_8 FILLER_39_1527 ();
 sg13g2_fill_1 FILLER_39_1538 ();
 sg13g2_fill_2 FILLER_39_1597 ();
 sg13g2_decap_8 FILLER_39_1629 ();
 sg13g2_decap_4 FILLER_39_1636 ();
 sg13g2_fill_1 FILLER_39_1640 ();
 sg13g2_decap_4 FILLER_39_1676 ();
 sg13g2_fill_1 FILLER_39_1680 ();
 sg13g2_decap_4 FILLER_39_1686 ();
 sg13g2_fill_1 FILLER_39_1690 ();
 sg13g2_decap_8 FILLER_39_1701 ();
 sg13g2_decap_4 FILLER_39_1708 ();
 sg13g2_fill_1 FILLER_39_1712 ();
 sg13g2_fill_2 FILLER_39_1752 ();
 sg13g2_fill_1 FILLER_39_1754 ();
 sg13g2_decap_8 FILLER_39_1761 ();
 sg13g2_decap_4 FILLER_39_1772 ();
 sg13g2_fill_1 FILLER_39_1781 ();
 sg13g2_decap_4 FILLER_39_1787 ();
 sg13g2_fill_1 FILLER_39_1791 ();
 sg13g2_decap_8 FILLER_39_1804 ();
 sg13g2_decap_4 FILLER_39_1811 ();
 sg13g2_decap_4 FILLER_39_1819 ();
 sg13g2_fill_1 FILLER_39_1823 ();
 sg13g2_decap_8 FILLER_39_1873 ();
 sg13g2_fill_1 FILLER_39_1885 ();
 sg13g2_fill_2 FILLER_39_1926 ();
 sg13g2_fill_1 FILLER_39_1928 ();
 sg13g2_fill_1 FILLER_39_1935 ();
 sg13g2_fill_2 FILLER_39_1976 ();
 sg13g2_decap_4 FILLER_39_1986 ();
 sg13g2_decap_4 FILLER_39_1994 ();
 sg13g2_decap_8 FILLER_39_2007 ();
 sg13g2_decap_8 FILLER_39_2014 ();
 sg13g2_decap_8 FILLER_39_2021 ();
 sg13g2_decap_4 FILLER_39_2028 ();
 sg13g2_fill_1 FILLER_39_2032 ();
 sg13g2_decap_4 FILLER_39_2038 ();
 sg13g2_fill_1 FILLER_39_2042 ();
 sg13g2_fill_1 FILLER_39_2095 ();
 sg13g2_decap_8 FILLER_39_2101 ();
 sg13g2_decap_8 FILLER_39_2108 ();
 sg13g2_decap_8 FILLER_39_2115 ();
 sg13g2_decap_8 FILLER_39_2122 ();
 sg13g2_decap_8 FILLER_39_2129 ();
 sg13g2_decap_8 FILLER_39_2136 ();
 sg13g2_fill_1 FILLER_39_2149 ();
 sg13g2_decap_8 FILLER_39_2154 ();
 sg13g2_fill_1 FILLER_39_2187 ();
 sg13g2_decap_4 FILLER_39_2224 ();
 sg13g2_decap_8 FILLER_39_2243 ();
 sg13g2_decap_8 FILLER_39_2250 ();
 sg13g2_decap_4 FILLER_39_2257 ();
 sg13g2_decap_8 FILLER_39_2292 ();
 sg13g2_decap_8 FILLER_39_2299 ();
 sg13g2_decap_8 FILLER_39_2346 ();
 sg13g2_decap_4 FILLER_39_2353 ();
 sg13g2_decap_8 FILLER_39_2361 ();
 sg13g2_decap_8 FILLER_39_2368 ();
 sg13g2_fill_1 FILLER_39_2375 ();
 sg13g2_fill_1 FILLER_39_2428 ();
 sg13g2_fill_1 FILLER_39_2455 ();
 sg13g2_fill_2 FILLER_39_2461 ();
 sg13g2_decap_8 FILLER_39_2478 ();
 sg13g2_decap_4 FILLER_39_2533 ();
 sg13g2_decap_8 FILLER_39_2585 ();
 sg13g2_decap_8 FILLER_39_2596 ();
 sg13g2_decap_8 FILLER_39_2603 ();
 sg13g2_decap_8 FILLER_39_2610 ();
 sg13g2_decap_8 FILLER_39_2647 ();
 sg13g2_decap_8 FILLER_39_2654 ();
 sg13g2_decap_8 FILLER_39_2661 ();
 sg13g2_fill_2 FILLER_39_2668 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_decap_4 FILLER_40_46 ();
 sg13g2_fill_2 FILLER_40_50 ();
 sg13g2_decap_8 FILLER_40_94 ();
 sg13g2_decap_4 FILLER_40_101 ();
 sg13g2_fill_1 FILLER_40_105 ();
 sg13g2_fill_1 FILLER_40_124 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_fill_1 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_199 ();
 sg13g2_decap_8 FILLER_40_206 ();
 sg13g2_decap_8 FILLER_40_213 ();
 sg13g2_fill_1 FILLER_40_224 ();
 sg13g2_fill_1 FILLER_40_232 ();
 sg13g2_fill_1 FILLER_40_244 ();
 sg13g2_decap_4 FILLER_40_276 ();
 sg13g2_fill_2 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_296 ();
 sg13g2_fill_2 FILLER_40_303 ();
 sg13g2_fill_2 FILLER_40_314 ();
 sg13g2_fill_1 FILLER_40_316 ();
 sg13g2_fill_1 FILLER_40_321 ();
 sg13g2_fill_2 FILLER_40_326 ();
 sg13g2_decap_4 FILLER_40_344 ();
 sg13g2_decap_8 FILLER_40_352 ();
 sg13g2_decap_8 FILLER_40_359 ();
 sg13g2_fill_2 FILLER_40_366 ();
 sg13g2_fill_1 FILLER_40_368 ();
 sg13g2_fill_2 FILLER_40_387 ();
 sg13g2_fill_1 FILLER_40_389 ();
 sg13g2_fill_1 FILLER_40_411 ();
 sg13g2_decap_4 FILLER_40_417 ();
 sg13g2_fill_2 FILLER_40_434 ();
 sg13g2_fill_2 FILLER_40_441 ();
 sg13g2_fill_2 FILLER_40_474 ();
 sg13g2_fill_1 FILLER_40_476 ();
 sg13g2_fill_2 FILLER_40_483 ();
 sg13g2_decap_8 FILLER_40_511 ();
 sg13g2_decap_8 FILLER_40_530 ();
 sg13g2_decap_8 FILLER_40_537 ();
 sg13g2_decap_8 FILLER_40_544 ();
 sg13g2_decap_8 FILLER_40_551 ();
 sg13g2_decap_4 FILLER_40_558 ();
 sg13g2_fill_1 FILLER_40_562 ();
 sg13g2_decap_8 FILLER_40_614 ();
 sg13g2_fill_1 FILLER_40_631 ();
 sg13g2_decap_8 FILLER_40_640 ();
 sg13g2_decap_8 FILLER_40_647 ();
 sg13g2_fill_1 FILLER_40_654 ();
 sg13g2_fill_2 FILLER_40_675 ();
 sg13g2_fill_1 FILLER_40_677 ();
 sg13g2_decap_4 FILLER_40_682 ();
 sg13g2_fill_2 FILLER_40_703 ();
 sg13g2_fill_1 FILLER_40_705 ();
 sg13g2_decap_8 FILLER_40_718 ();
 sg13g2_decap_8 FILLER_40_725 ();
 sg13g2_decap_4 FILLER_40_732 ();
 sg13g2_fill_2 FILLER_40_736 ();
 sg13g2_fill_2 FILLER_40_753 ();
 sg13g2_fill_1 FILLER_40_755 ();
 sg13g2_decap_8 FILLER_40_759 ();
 sg13g2_fill_2 FILLER_40_766 ();
 sg13g2_decap_8 FILLER_40_773 ();
 sg13g2_decap_8 FILLER_40_785 ();
 sg13g2_decap_8 FILLER_40_792 ();
 sg13g2_decap_4 FILLER_40_799 ();
 sg13g2_fill_1 FILLER_40_803 ();
 sg13g2_fill_2 FILLER_40_838 ();
 sg13g2_decap_8 FILLER_40_874 ();
 sg13g2_fill_2 FILLER_40_881 ();
 sg13g2_fill_1 FILLER_40_883 ();
 sg13g2_fill_2 FILLER_40_888 ();
 sg13g2_fill_2 FILLER_40_893 ();
 sg13g2_fill_1 FILLER_40_895 ();
 sg13g2_decap_4 FILLER_40_900 ();
 sg13g2_fill_2 FILLER_40_908 ();
 sg13g2_fill_2 FILLER_40_937 ();
 sg13g2_fill_1 FILLER_40_939 ();
 sg13g2_decap_4 FILLER_40_953 ();
 sg13g2_fill_1 FILLER_40_957 ();
 sg13g2_decap_8 FILLER_40_962 ();
 sg13g2_fill_1 FILLER_40_999 ();
 sg13g2_fill_1 FILLER_40_1006 ();
 sg13g2_fill_1 FILLER_40_1033 ();
 sg13g2_decap_4 FILLER_40_1040 ();
 sg13g2_decap_8 FILLER_40_1070 ();
 sg13g2_fill_2 FILLER_40_1077 ();
 sg13g2_fill_2 FILLER_40_1088 ();
 sg13g2_fill_2 FILLER_40_1116 ();
 sg13g2_decap_8 FILLER_40_1122 ();
 sg13g2_decap_8 FILLER_40_1129 ();
 sg13g2_fill_1 FILLER_40_1136 ();
 sg13g2_fill_2 FILLER_40_1150 ();
 sg13g2_fill_1 FILLER_40_1152 ();
 sg13g2_decap_8 FILLER_40_1178 ();
 sg13g2_decap_8 FILLER_40_1185 ();
 sg13g2_decap_8 FILLER_40_1192 ();
 sg13g2_fill_2 FILLER_40_1199 ();
 sg13g2_decap_8 FILLER_40_1205 ();
 sg13g2_decap_4 FILLER_40_1212 ();
 sg13g2_fill_2 FILLER_40_1216 ();
 sg13g2_fill_1 FILLER_40_1223 ();
 sg13g2_decap_4 FILLER_40_1254 ();
 sg13g2_fill_1 FILLER_40_1258 ();
 sg13g2_fill_1 FILLER_40_1264 ();
 sg13g2_fill_1 FILLER_40_1271 ();
 sg13g2_fill_1 FILLER_40_1276 ();
 sg13g2_fill_2 FILLER_40_1312 ();
 sg13g2_fill_2 FILLER_40_1324 ();
 sg13g2_fill_1 FILLER_40_1334 ();
 sg13g2_decap_4 FILLER_40_1355 ();
 sg13g2_fill_2 FILLER_40_1359 ();
 sg13g2_decap_8 FILLER_40_1387 ();
 sg13g2_decap_8 FILLER_40_1394 ();
 sg13g2_decap_8 FILLER_40_1401 ();
 sg13g2_decap_8 FILLER_40_1408 ();
 sg13g2_fill_2 FILLER_40_1415 ();
 sg13g2_fill_1 FILLER_40_1422 ();
 sg13g2_decap_8 FILLER_40_1455 ();
 sg13g2_fill_1 FILLER_40_1462 ();
 sg13g2_decap_8 FILLER_40_1471 ();
 sg13g2_decap_4 FILLER_40_1478 ();
 sg13g2_fill_1 FILLER_40_1482 ();
 sg13g2_fill_1 FILLER_40_1517 ();
 sg13g2_decap_4 FILLER_40_1523 ();
 sg13g2_fill_2 FILLER_40_1527 ();
 sg13g2_decap_8 FILLER_40_1534 ();
 sg13g2_fill_1 FILLER_40_1564 ();
 sg13g2_decap_4 FILLER_40_1597 ();
 sg13g2_fill_2 FILLER_40_1601 ();
 sg13g2_decap_8 FILLER_40_1608 ();
 sg13g2_fill_2 FILLER_40_1615 ();
 sg13g2_fill_1 FILLER_40_1617 ();
 sg13g2_decap_8 FILLER_40_1623 ();
 sg13g2_decap_4 FILLER_40_1630 ();
 sg13g2_fill_1 FILLER_40_1643 ();
 sg13g2_fill_1 FILLER_40_1649 ();
 sg13g2_decap_8 FILLER_40_1676 ();
 sg13g2_fill_1 FILLER_40_1683 ();
 sg13g2_fill_2 FILLER_40_1726 ();
 sg13g2_decap_4 FILLER_40_1736 ();
 sg13g2_fill_2 FILLER_40_1740 ();
 sg13g2_decap_8 FILLER_40_1757 ();
 sg13g2_decap_8 FILLER_40_1764 ();
 sg13g2_fill_1 FILLER_40_1771 ();
 sg13g2_decap_8 FILLER_40_1778 ();
 sg13g2_decap_8 FILLER_40_1785 ();
 sg13g2_decap_8 FILLER_40_1792 ();
 sg13g2_decap_4 FILLER_40_1799 ();
 sg13g2_fill_2 FILLER_40_1803 ();
 sg13g2_fill_1 FILLER_40_1818 ();
 sg13g2_decap_8 FILLER_40_1859 ();
 sg13g2_decap_4 FILLER_40_1870 ();
 sg13g2_fill_2 FILLER_40_1874 ();
 sg13g2_fill_2 FILLER_40_1902 ();
 sg13g2_fill_1 FILLER_40_1904 ();
 sg13g2_decap_8 FILLER_40_1908 ();
 sg13g2_decap_8 FILLER_40_1915 ();
 sg13g2_decap_4 FILLER_40_1922 ();
 sg13g2_fill_2 FILLER_40_1926 ();
 sg13g2_decap_8 FILLER_40_1932 ();
 sg13g2_decap_8 FILLER_40_1939 ();
 sg13g2_decap_4 FILLER_40_1946 ();
 sg13g2_fill_2 FILLER_40_1950 ();
 sg13g2_decap_8 FILLER_40_1965 ();
 sg13g2_decap_8 FILLER_40_1972 ();
 sg13g2_fill_2 FILLER_40_1979 ();
 sg13g2_fill_1 FILLER_40_1981 ();
 sg13g2_decap_8 FILLER_40_1987 ();
 sg13g2_decap_8 FILLER_40_1994 ();
 sg13g2_decap_8 FILLER_40_2001 ();
 sg13g2_fill_1 FILLER_40_2008 ();
 sg13g2_fill_2 FILLER_40_2018 ();
 sg13g2_fill_1 FILLER_40_2020 ();
 sg13g2_fill_1 FILLER_40_2032 ();
 sg13g2_fill_1 FILLER_40_2037 ();
 sg13g2_fill_2 FILLER_40_2073 ();
 sg13g2_fill_1 FILLER_40_2075 ();
 sg13g2_fill_2 FILLER_40_2080 ();
 sg13g2_fill_1 FILLER_40_2108 ();
 sg13g2_fill_1 FILLER_40_2113 ();
 sg13g2_fill_2 FILLER_40_2120 ();
 sg13g2_fill_1 FILLER_40_2148 ();
 sg13g2_fill_2 FILLER_40_2180 ();
 sg13g2_fill_1 FILLER_40_2193 ();
 sg13g2_fill_2 FILLER_40_2198 ();
 sg13g2_fill_1 FILLER_40_2204 ();
 sg13g2_fill_2 FILLER_40_2211 ();
 sg13g2_decap_8 FILLER_40_2243 ();
 sg13g2_decap_8 FILLER_40_2250 ();
 sg13g2_fill_2 FILLER_40_2257 ();
 sg13g2_fill_1 FILLER_40_2272 ();
 sg13g2_decap_8 FILLER_40_2286 ();
 sg13g2_fill_2 FILLER_40_2293 ();
 sg13g2_fill_1 FILLER_40_2295 ();
 sg13g2_fill_2 FILLER_40_2301 ();
 sg13g2_decap_4 FILLER_40_2329 ();
 sg13g2_decap_4 FILLER_40_2359 ();
 sg13g2_decap_4 FILLER_40_2368 ();
 sg13g2_decap_8 FILLER_40_2381 ();
 sg13g2_fill_2 FILLER_40_2388 ();
 sg13g2_fill_1 FILLER_40_2390 ();
 sg13g2_fill_1 FILLER_40_2395 ();
 sg13g2_fill_2 FILLER_40_2406 ();
 sg13g2_fill_1 FILLER_40_2408 ();
 sg13g2_fill_2 FILLER_40_2415 ();
 sg13g2_fill_2 FILLER_40_2422 ();
 sg13g2_fill_1 FILLER_40_2432 ();
 sg13g2_decap_8 FILLER_40_2439 ();
 sg13g2_fill_1 FILLER_40_2451 ();
 sg13g2_fill_1 FILLER_40_2457 ();
 sg13g2_decap_8 FILLER_40_2489 ();
 sg13g2_fill_1 FILLER_40_2496 ();
 sg13g2_fill_2 FILLER_40_2502 ();
 sg13g2_decap_4 FILLER_40_2510 ();
 sg13g2_fill_1 FILLER_40_2514 ();
 sg13g2_decap_8 FILLER_40_2520 ();
 sg13g2_fill_2 FILLER_40_2527 ();
 sg13g2_decap_8 FILLER_40_2534 ();
 sg13g2_decap_4 FILLER_40_2541 ();
 sg13g2_fill_2 FILLER_40_2545 ();
 sg13g2_decap_4 FILLER_40_2556 ();
 sg13g2_fill_2 FILLER_40_2598 ();
 sg13g2_fill_1 FILLER_40_2600 ();
 sg13g2_decap_8 FILLER_40_2627 ();
 sg13g2_decap_8 FILLER_40_2634 ();
 sg13g2_decap_8 FILLER_40_2641 ();
 sg13g2_decap_8 FILLER_40_2648 ();
 sg13g2_decap_8 FILLER_40_2655 ();
 sg13g2_decap_8 FILLER_40_2662 ();
 sg13g2_fill_1 FILLER_40_2669 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_4 FILLER_41_14 ();
 sg13g2_fill_1 FILLER_41_18 ();
 sg13g2_decap_4 FILLER_41_23 ();
 sg13g2_fill_1 FILLER_41_27 ();
 sg13g2_decap_8 FILLER_41_41 ();
 sg13g2_decap_8 FILLER_41_48 ();
 sg13g2_fill_2 FILLER_41_55 ();
 sg13g2_fill_1 FILLER_41_57 ();
 sg13g2_decap_4 FILLER_41_62 ();
 sg13g2_fill_1 FILLER_41_66 ();
 sg13g2_fill_2 FILLER_41_79 ();
 sg13g2_fill_1 FILLER_41_81 ();
 sg13g2_decap_8 FILLER_41_152 ();
 sg13g2_decap_8 FILLER_41_159 ();
 sg13g2_decap_8 FILLER_41_166 ();
 sg13g2_fill_2 FILLER_41_173 ();
 sg13g2_fill_1 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_179 ();
 sg13g2_decap_4 FILLER_41_186 ();
 sg13g2_decap_8 FILLER_41_204 ();
 sg13g2_fill_2 FILLER_41_239 ();
 sg13g2_fill_2 FILLER_41_250 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_fill_2 FILLER_41_266 ();
 sg13g2_fill_1 FILLER_41_268 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_4 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_340 ();
 sg13g2_decap_8 FILLER_41_347 ();
 sg13g2_fill_1 FILLER_41_354 ();
 sg13g2_decap_4 FILLER_41_360 ();
 sg13g2_decap_8 FILLER_41_368 ();
 sg13g2_decap_8 FILLER_41_375 ();
 sg13g2_fill_2 FILLER_41_382 ();
 sg13g2_decap_4 FILLER_41_392 ();
 sg13g2_fill_1 FILLER_41_396 ();
 sg13g2_decap_8 FILLER_41_402 ();
 sg13g2_decap_4 FILLER_41_423 ();
 sg13g2_fill_2 FILLER_41_427 ();
 sg13g2_fill_2 FILLER_41_435 ();
 sg13g2_fill_1 FILLER_41_437 ();
 sg13g2_fill_2 FILLER_41_446 ();
 sg13g2_decap_8 FILLER_41_451 ();
 sg13g2_decap_8 FILLER_41_458 ();
 sg13g2_decap_8 FILLER_41_465 ();
 sg13g2_decap_8 FILLER_41_472 ();
 sg13g2_decap_4 FILLER_41_479 ();
 sg13g2_fill_1 FILLER_41_483 ();
 sg13g2_decap_8 FILLER_41_503 ();
 sg13g2_decap_4 FILLER_41_510 ();
 sg13g2_fill_1 FILLER_41_514 ();
 sg13g2_fill_2 FILLER_41_527 ();
 sg13g2_decap_8 FILLER_41_538 ();
 sg13g2_fill_2 FILLER_41_545 ();
 sg13g2_fill_1 FILLER_41_547 ();
 sg13g2_decap_8 FILLER_41_553 ();
 sg13g2_decap_4 FILLER_41_560 ();
 sg13g2_fill_1 FILLER_41_564 ();
 sg13g2_decap_4 FILLER_41_591 ();
 sg13g2_fill_1 FILLER_41_603 ();
 sg13g2_fill_2 FILLER_41_609 ();
 sg13g2_decap_8 FILLER_41_616 ();
 sg13g2_decap_8 FILLER_41_623 ();
 sg13g2_decap_8 FILLER_41_630 ();
 sg13g2_decap_8 FILLER_41_637 ();
 sg13g2_decap_8 FILLER_41_644 ();
 sg13g2_decap_4 FILLER_41_657 ();
 sg13g2_decap_8 FILLER_41_670 ();
 sg13g2_decap_4 FILLER_41_677 ();
 sg13g2_decap_4 FILLER_41_689 ();
 sg13g2_fill_2 FILLER_41_693 ();
 sg13g2_fill_2 FILLER_41_715 ();
 sg13g2_decap_4 FILLER_41_739 ();
 sg13g2_decap_8 FILLER_41_748 ();
 sg13g2_fill_2 FILLER_41_755 ();
 sg13g2_fill_2 FILLER_41_765 ();
 sg13g2_decap_8 FILLER_41_780 ();
 sg13g2_fill_2 FILLER_41_787 ();
 sg13g2_decap_8 FILLER_41_793 ();
 sg13g2_decap_4 FILLER_41_800 ();
 sg13g2_fill_1 FILLER_41_804 ();
 sg13g2_decap_4 FILLER_41_810 ();
 sg13g2_fill_1 FILLER_41_814 ();
 sg13g2_fill_1 FILLER_41_819 ();
 sg13g2_decap_8 FILLER_41_824 ();
 sg13g2_decap_4 FILLER_41_883 ();
 sg13g2_decap_4 FILLER_41_906 ();
 sg13g2_fill_1 FILLER_41_915 ();
 sg13g2_decap_4 FILLER_41_927 ();
 sg13g2_decap_8 FILLER_41_944 ();
 sg13g2_fill_2 FILLER_41_951 ();
 sg13g2_fill_2 FILLER_41_958 ();
 sg13g2_fill_1 FILLER_41_986 ();
 sg13g2_fill_2 FILLER_41_992 ();
 sg13g2_fill_2 FILLER_41_998 ();
 sg13g2_fill_2 FILLER_41_1005 ();
 sg13g2_fill_1 FILLER_41_1040 ();
 sg13g2_decap_8 FILLER_41_1047 ();
 sg13g2_decap_8 FILLER_41_1054 ();
 sg13g2_fill_2 FILLER_41_1061 ();
 sg13g2_fill_1 FILLER_41_1063 ();
 sg13g2_fill_2 FILLER_41_1068 ();
 sg13g2_fill_2 FILLER_41_1099 ();
 sg13g2_decap_4 FILLER_41_1109 ();
 sg13g2_fill_2 FILLER_41_1113 ();
 sg13g2_decap_4 FILLER_41_1120 ();
 sg13g2_fill_1 FILLER_41_1124 ();
 sg13g2_decap_8 FILLER_41_1130 ();
 sg13g2_decap_8 FILLER_41_1137 ();
 sg13g2_fill_2 FILLER_41_1149 ();
 sg13g2_fill_1 FILLER_41_1151 ();
 sg13g2_fill_1 FILLER_41_1160 ();
 sg13g2_decap_8 FILLER_41_1187 ();
 sg13g2_fill_2 FILLER_41_1194 ();
 sg13g2_fill_2 FILLER_41_1222 ();
 sg13g2_fill_1 FILLER_41_1224 ();
 sg13g2_fill_2 FILLER_41_1251 ();
 sg13g2_decap_4 FILLER_41_1265 ();
 sg13g2_fill_1 FILLER_41_1269 ();
 sg13g2_fill_2 FILLER_41_1306 ();
 sg13g2_fill_2 FILLER_41_1331 ();
 sg13g2_fill_1 FILLER_41_1333 ();
 sg13g2_fill_2 FILLER_41_1366 ();
 sg13g2_fill_1 FILLER_41_1368 ();
 sg13g2_decap_8 FILLER_41_1379 ();
 sg13g2_fill_2 FILLER_41_1386 ();
 sg13g2_fill_1 FILLER_41_1388 ();
 sg13g2_decap_8 FILLER_41_1393 ();
 sg13g2_decap_8 FILLER_41_1400 ();
 sg13g2_decap_8 FILLER_41_1407 ();
 sg13g2_decap_8 FILLER_41_1414 ();
 sg13g2_decap_4 FILLER_41_1421 ();
 sg13g2_decap_4 FILLER_41_1430 ();
 sg13g2_decap_8 FILLER_41_1452 ();
 sg13g2_decap_8 FILLER_41_1459 ();
 sg13g2_fill_2 FILLER_41_1466 ();
 sg13g2_decap_8 FILLER_41_1473 ();
 sg13g2_fill_2 FILLER_41_1486 ();
 sg13g2_fill_1 FILLER_41_1488 ();
 sg13g2_fill_2 FILLER_41_1493 ();
 sg13g2_decap_8 FILLER_41_1503 ();
 sg13g2_decap_4 FILLER_41_1510 ();
 sg13g2_fill_1 FILLER_41_1514 ();
 sg13g2_fill_2 FILLER_41_1546 ();
 sg13g2_fill_1 FILLER_41_1600 ();
 sg13g2_fill_2 FILLER_41_1605 ();
 sg13g2_fill_2 FILLER_41_1633 ();
 sg13g2_fill_1 FILLER_41_1635 ();
 sg13g2_decap_8 FILLER_41_1666 ();
 sg13g2_fill_2 FILLER_41_1673 ();
 sg13g2_decap_8 FILLER_41_1700 ();
 sg13g2_fill_2 FILLER_41_1707 ();
 sg13g2_fill_2 FILLER_41_1740 ();
 sg13g2_decap_8 FILLER_41_1799 ();
 sg13g2_decap_8 FILLER_41_1806 ();
 sg13g2_decap_4 FILLER_41_1813 ();
 sg13g2_fill_1 FILLER_41_1817 ();
 sg13g2_decap_8 FILLER_41_1822 ();
 sg13g2_fill_2 FILLER_41_1833 ();
 sg13g2_fill_1 FILLER_41_1840 ();
 sg13g2_fill_2 FILLER_41_1850 ();
 sg13g2_fill_1 FILLER_41_1852 ();
 sg13g2_fill_2 FILLER_41_1864 ();
 sg13g2_fill_1 FILLER_41_1866 ();
 sg13g2_decap_8 FILLER_41_1911 ();
 sg13g2_decap_4 FILLER_41_1918 ();
 sg13g2_decap_8 FILLER_41_1931 ();
 sg13g2_fill_2 FILLER_41_1938 ();
 sg13g2_decap_8 FILLER_41_1944 ();
 sg13g2_decap_8 FILLER_41_1951 ();
 sg13g2_fill_1 FILLER_41_1958 ();
 sg13g2_decap_8 FILLER_41_2028 ();
 sg13g2_fill_2 FILLER_41_2035 ();
 sg13g2_decap_8 FILLER_41_2042 ();
 sg13g2_fill_1 FILLER_41_2049 ();
 sg13g2_decap_4 FILLER_41_2055 ();
 sg13g2_fill_2 FILLER_41_2059 ();
 sg13g2_decap_4 FILLER_41_2069 ();
 sg13g2_fill_2 FILLER_41_2073 ();
 sg13g2_fill_1 FILLER_41_2089 ();
 sg13g2_fill_1 FILLER_41_2094 ();
 sg13g2_decap_8 FILLER_41_2126 ();
 sg13g2_fill_1 FILLER_41_2142 ();
 sg13g2_fill_2 FILLER_41_2151 ();
 sg13g2_fill_1 FILLER_41_2157 ();
 sg13g2_fill_1 FILLER_41_2167 ();
 sg13g2_decap_8 FILLER_41_2172 ();
 sg13g2_fill_1 FILLER_41_2179 ();
 sg13g2_decap_8 FILLER_41_2186 ();
 sg13g2_fill_2 FILLER_41_2193 ();
 sg13g2_fill_1 FILLER_41_2200 ();
 sg13g2_decap_4 FILLER_41_2206 ();
 sg13g2_fill_1 FILLER_41_2210 ();
 sg13g2_decap_8 FILLER_41_2215 ();
 sg13g2_decap_8 FILLER_41_2295 ();
 sg13g2_fill_2 FILLER_41_2307 ();
 sg13g2_fill_1 FILLER_41_2309 ();
 sg13g2_fill_2 FILLER_41_2323 ();
 sg13g2_fill_2 FILLER_41_2376 ();
 sg13g2_decap_8 FILLER_41_2404 ();
 sg13g2_fill_2 FILLER_41_2411 ();
 sg13g2_decap_4 FILLER_41_2428 ();
 sg13g2_fill_1 FILLER_41_2432 ();
 sg13g2_decap_4 FILLER_41_2439 ();
 sg13g2_fill_2 FILLER_41_2449 ();
 sg13g2_decap_4 FILLER_41_2477 ();
 sg13g2_fill_1 FILLER_41_2485 ();
 sg13g2_fill_1 FILLER_41_2517 ();
 sg13g2_fill_2 FILLER_41_2593 ();
 sg13g2_decap_8 FILLER_41_2608 ();
 sg13g2_decap_8 FILLER_41_2615 ();
 sg13g2_decap_8 FILLER_41_2622 ();
 sg13g2_decap_8 FILLER_41_2629 ();
 sg13g2_decap_8 FILLER_41_2636 ();
 sg13g2_decap_8 FILLER_41_2643 ();
 sg13g2_decap_8 FILLER_41_2650 ();
 sg13g2_decap_8 FILLER_41_2657 ();
 sg13g2_decap_4 FILLER_41_2664 ();
 sg13g2_fill_2 FILLER_41_2668 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_9 ();
 sg13g2_fill_2 FILLER_42_18 ();
 sg13g2_decap_8 FILLER_42_25 ();
 sg13g2_decap_8 FILLER_42_32 ();
 sg13g2_fill_2 FILLER_42_39 ();
 sg13g2_fill_1 FILLER_42_41 ();
 sg13g2_fill_2 FILLER_42_47 ();
 sg13g2_fill_1 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_fill_2 FILLER_42_84 ();
 sg13g2_fill_1 FILLER_42_86 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_4 FILLER_42_98 ();
 sg13g2_fill_1 FILLER_42_102 ();
 sg13g2_fill_2 FILLER_42_125 ();
 sg13g2_fill_1 FILLER_42_127 ();
 sg13g2_fill_1 FILLER_42_133 ();
 sg13g2_fill_1 FILLER_42_139 ();
 sg13g2_decap_4 FILLER_42_144 ();
 sg13g2_fill_1 FILLER_42_148 ();
 sg13g2_decap_8 FILLER_42_153 ();
 sg13g2_decap_8 FILLER_42_160 ();
 sg13g2_decap_4 FILLER_42_167 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_decap_4 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_236 ();
 sg13g2_decap_8 FILLER_42_246 ();
 sg13g2_decap_8 FILLER_42_253 ();
 sg13g2_decap_8 FILLER_42_260 ();
 sg13g2_decap_8 FILLER_42_267 ();
 sg13g2_decap_4 FILLER_42_274 ();
 sg13g2_fill_1 FILLER_42_283 ();
 sg13g2_decap_4 FILLER_42_288 ();
 sg13g2_fill_2 FILLER_42_292 ();
 sg13g2_fill_1 FILLER_42_301 ();
 sg13g2_fill_2 FILLER_42_307 ();
 sg13g2_fill_1 FILLER_42_309 ();
 sg13g2_fill_2 FILLER_42_320 ();
 sg13g2_fill_1 FILLER_42_331 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_389 ();
 sg13g2_decap_8 FILLER_42_396 ();
 sg13g2_fill_1 FILLER_42_403 ();
 sg13g2_decap_4 FILLER_42_434 ();
 sg13g2_fill_1 FILLER_42_438 ();
 sg13g2_decap_4 FILLER_42_445 ();
 sg13g2_fill_2 FILLER_42_449 ();
 sg13g2_decap_8 FILLER_42_455 ();
 sg13g2_decap_8 FILLER_42_462 ();
 sg13g2_decap_8 FILLER_42_469 ();
 sg13g2_fill_2 FILLER_42_476 ();
 sg13g2_fill_1 FILLER_42_483 ();
 sg13g2_fill_2 FILLER_42_487 ();
 sg13g2_fill_1 FILLER_42_489 ();
 sg13g2_decap_8 FILLER_42_493 ();
 sg13g2_decap_8 FILLER_42_500 ();
 sg13g2_decap_8 FILLER_42_507 ();
 sg13g2_decap_8 FILLER_42_514 ();
 sg13g2_decap_4 FILLER_42_521 ();
 sg13g2_fill_1 FILLER_42_525 ();
 sg13g2_decap_4 FILLER_42_539 ();
 sg13g2_decap_4 FILLER_42_548 ();
 sg13g2_decap_8 FILLER_42_557 ();
 sg13g2_fill_1 FILLER_42_564 ();
 sg13g2_decap_8 FILLER_42_569 ();
 sg13g2_fill_1 FILLER_42_576 ();
 sg13g2_decap_8 FILLER_42_592 ();
 sg13g2_decap_4 FILLER_42_599 ();
 sg13g2_fill_2 FILLER_42_603 ();
 sg13g2_decap_8 FILLER_42_619 ();
 sg13g2_fill_1 FILLER_42_626 ();
 sg13g2_fill_2 FILLER_42_633 ();
 sg13g2_fill_2 FILLER_42_645 ();
 sg13g2_fill_1 FILLER_42_647 ();
 sg13g2_fill_2 FILLER_42_653 ();
 sg13g2_fill_1 FILLER_42_655 ();
 sg13g2_decap_8 FILLER_42_671 ();
 sg13g2_fill_2 FILLER_42_678 ();
 sg13g2_fill_1 FILLER_42_680 ();
 sg13g2_fill_1 FILLER_42_707 ();
 sg13g2_fill_2 FILLER_42_713 ();
 sg13g2_fill_2 FILLER_42_718 ();
 sg13g2_fill_1 FILLER_42_723 ();
 sg13g2_decap_4 FILLER_42_750 ();
 sg13g2_fill_1 FILLER_42_767 ();
 sg13g2_decap_8 FILLER_42_794 ();
 sg13g2_decap_4 FILLER_42_801 ();
 sg13g2_fill_1 FILLER_42_805 ();
 sg13g2_decap_8 FILLER_42_832 ();
 sg13g2_decap_8 FILLER_42_839 ();
 sg13g2_decap_4 FILLER_42_846 ();
 sg13g2_fill_1 FILLER_42_850 ();
 sg13g2_decap_4 FILLER_42_869 ();
 sg13g2_decap_4 FILLER_42_893 ();
 sg13g2_decap_8 FILLER_42_902 ();
 sg13g2_fill_2 FILLER_42_909 ();
 sg13g2_fill_2 FILLER_42_925 ();
 sg13g2_fill_1 FILLER_42_927 ();
 sg13g2_decap_8 FILLER_42_932 ();
 sg13g2_decap_8 FILLER_42_939 ();
 sg13g2_decap_8 FILLER_42_946 ();
 sg13g2_decap_4 FILLER_42_953 ();
 sg13g2_fill_1 FILLER_42_957 ();
 sg13g2_fill_1 FILLER_42_973 ();
 sg13g2_fill_2 FILLER_42_978 ();
 sg13g2_fill_1 FILLER_42_980 ();
 sg13g2_decap_4 FILLER_42_986 ();
 sg13g2_fill_1 FILLER_42_990 ();
 sg13g2_decap_8 FILLER_42_994 ();
 sg13g2_decap_4 FILLER_42_1001 ();
 sg13g2_fill_2 FILLER_42_1005 ();
 sg13g2_fill_2 FILLER_42_1011 ();
 sg13g2_decap_8 FILLER_42_1017 ();
 sg13g2_fill_1 FILLER_42_1024 ();
 sg13g2_fill_1 FILLER_42_1033 ();
 sg13g2_fill_1 FILLER_42_1058 ();
 sg13g2_fill_2 FILLER_42_1064 ();
 sg13g2_decap_8 FILLER_42_1076 ();
 sg13g2_decap_8 FILLER_42_1083 ();
 sg13g2_fill_2 FILLER_42_1090 ();
 sg13g2_fill_2 FILLER_42_1097 ();
 sg13g2_decap_8 FILLER_42_1130 ();
 sg13g2_decap_8 FILLER_42_1137 ();
 sg13g2_decap_4 FILLER_42_1144 ();
 sg13g2_fill_1 FILLER_42_1148 ();
 sg13g2_decap_4 FILLER_42_1153 ();
 sg13g2_decap_8 FILLER_42_1161 ();
 sg13g2_decap_8 FILLER_42_1168 ();
 sg13g2_decap_8 FILLER_42_1175 ();
 sg13g2_decap_8 FILLER_42_1182 ();
 sg13g2_fill_2 FILLER_42_1189 ();
 sg13g2_fill_1 FILLER_42_1191 ();
 sg13g2_fill_1 FILLER_42_1196 ();
 sg13g2_fill_1 FILLER_42_1233 ();
 sg13g2_fill_2 FILLER_42_1275 ();
 sg13g2_fill_1 FILLER_42_1280 ();
 sg13g2_fill_1 FILLER_42_1287 ();
 sg13g2_fill_1 FILLER_42_1294 ();
 sg13g2_fill_2 FILLER_42_1335 ();
 sg13g2_fill_2 FILLER_42_1365 ();
 sg13g2_fill_1 FILLER_42_1367 ();
 sg13g2_decap_8 FILLER_42_1376 ();
 sg13g2_decap_8 FILLER_42_1383 ();
 sg13g2_fill_1 FILLER_42_1390 ();
 sg13g2_decap_4 FILLER_42_1435 ();
 sg13g2_fill_1 FILLER_42_1439 ();
 sg13g2_decap_8 FILLER_42_1444 ();
 sg13g2_decap_8 FILLER_42_1451 ();
 sg13g2_decap_4 FILLER_42_1467 ();
 sg13g2_decap_8 FILLER_42_1497 ();
 sg13g2_decap_4 FILLER_42_1504 ();
 sg13g2_fill_2 FILLER_42_1508 ();
 sg13g2_fill_2 FILLER_42_1513 ();
 sg13g2_decap_8 FILLER_42_1520 ();
 sg13g2_fill_1 FILLER_42_1531 ();
 sg13g2_decap_4 FILLER_42_1538 ();
 sg13g2_fill_1 FILLER_42_1542 ();
 sg13g2_decap_8 FILLER_42_1579 ();
 sg13g2_decap_4 FILLER_42_1586 ();
 sg13g2_fill_1 FILLER_42_1590 ();
 sg13g2_fill_2 FILLER_42_1617 ();
 sg13g2_fill_1 FILLER_42_1619 ();
 sg13g2_decap_4 FILLER_42_1624 ();
 sg13g2_fill_2 FILLER_42_1628 ();
 sg13g2_fill_1 FILLER_42_1647 ();
 sg13g2_decap_8 FILLER_42_1665 ();
 sg13g2_decap_4 FILLER_42_1672 ();
 sg13g2_fill_1 FILLER_42_1676 ();
 sg13g2_fill_1 FILLER_42_1708 ();
 sg13g2_decap_8 FILLER_42_1718 ();
 sg13g2_fill_1 FILLER_42_1756 ();
 sg13g2_decap_8 FILLER_42_1762 ();
 sg13g2_fill_2 FILLER_42_1769 ();
 sg13g2_fill_1 FILLER_42_1776 ();
 sg13g2_fill_1 FILLER_42_1781 ();
 sg13g2_decap_4 FILLER_42_1785 ();
 sg13g2_fill_2 FILLER_42_1789 ();
 sg13g2_decap_4 FILLER_42_1797 ();
 sg13g2_fill_1 FILLER_42_1801 ();
 sg13g2_fill_2 FILLER_42_1824 ();
 sg13g2_decap_8 FILLER_42_1833 ();
 sg13g2_decap_8 FILLER_42_1840 ();
 sg13g2_decap_8 FILLER_42_1860 ();
 sg13g2_fill_2 FILLER_42_1867 ();
 sg13g2_fill_1 FILLER_42_1869 ();
 sg13g2_decap_4 FILLER_42_1882 ();
 sg13g2_fill_1 FILLER_42_1886 ();
 sg13g2_fill_1 FILLER_42_1891 ();
 sg13g2_fill_1 FILLER_42_1918 ();
 sg13g2_fill_2 FILLER_42_1951 ();
 sg13g2_decap_4 FILLER_42_1960 ();
 sg13g2_fill_2 FILLER_42_1964 ();
 sg13g2_decap_8 FILLER_42_1980 ();
 sg13g2_decap_8 FILLER_42_1987 ();
 sg13g2_decap_8 FILLER_42_1994 ();
 sg13g2_decap_4 FILLER_42_2001 ();
 sg13g2_fill_1 FILLER_42_2005 ();
 sg13g2_fill_2 FILLER_42_2023 ();
 sg13g2_fill_1 FILLER_42_2039 ();
 sg13g2_fill_2 FILLER_42_2078 ();
 sg13g2_fill_1 FILLER_42_2080 ();
 sg13g2_fill_2 FILLER_42_2085 ();
 sg13g2_fill_1 FILLER_42_2087 ();
 sg13g2_decap_8 FILLER_42_2094 ();
 sg13g2_decap_8 FILLER_42_2101 ();
 sg13g2_decap_8 FILLER_42_2108 ();
 sg13g2_decap_8 FILLER_42_2115 ();
 sg13g2_decap_4 FILLER_42_2122 ();
 sg13g2_fill_1 FILLER_42_2126 ();
 sg13g2_decap_4 FILLER_42_2130 ();
 sg13g2_fill_1 FILLER_42_2134 ();
 sg13g2_fill_2 FILLER_42_2145 ();
 sg13g2_fill_1 FILLER_42_2147 ();
 sg13g2_fill_2 FILLER_42_2152 ();
 sg13g2_decap_4 FILLER_42_2197 ();
 sg13g2_fill_2 FILLER_42_2201 ();
 sg13g2_decap_8 FILLER_42_2212 ();
 sg13g2_fill_2 FILLER_42_2277 ();
 sg13g2_decap_8 FILLER_42_2283 ();
 sg13g2_decap_8 FILLER_42_2290 ();
 sg13g2_fill_2 FILLER_42_2297 ();
 sg13g2_fill_1 FILLER_42_2299 ();
 sg13g2_decap_8 FILLER_42_2304 ();
 sg13g2_fill_1 FILLER_42_2311 ();
 sg13g2_decap_4 FILLER_42_2318 ();
 sg13g2_fill_2 FILLER_42_2322 ();
 sg13g2_decap_4 FILLER_42_2350 ();
 sg13g2_fill_2 FILLER_42_2380 ();
 sg13g2_fill_1 FILLER_42_2382 ();
 sg13g2_decap_4 FILLER_42_2409 ();
 sg13g2_decap_8 FILLER_42_2468 ();
 sg13g2_decap_4 FILLER_42_2475 ();
 sg13g2_fill_2 FILLER_42_2479 ();
 sg13g2_decap_4 FILLER_42_2512 ();
 sg13g2_fill_1 FILLER_42_2516 ();
 sg13g2_decap_8 FILLER_42_2530 ();
 sg13g2_decap_8 FILLER_42_2537 ();
 sg13g2_fill_2 FILLER_42_2544 ();
 sg13g2_fill_1 FILLER_42_2555 ();
 sg13g2_decap_8 FILLER_42_2578 ();
 sg13g2_decap_4 FILLER_42_2585 ();
 sg13g2_fill_2 FILLER_42_2593 ();
 sg13g2_decap_8 FILLER_42_2598 ();
 sg13g2_decap_8 FILLER_42_2605 ();
 sg13g2_decap_8 FILLER_42_2612 ();
 sg13g2_decap_4 FILLER_42_2619 ();
 sg13g2_decap_4 FILLER_42_2627 ();
 sg13g2_fill_2 FILLER_42_2631 ();
 sg13g2_decap_8 FILLER_42_2637 ();
 sg13g2_decap_8 FILLER_42_2644 ();
 sg13g2_decap_8 FILLER_42_2651 ();
 sg13g2_decap_8 FILLER_42_2658 ();
 sg13g2_decap_4 FILLER_42_2665 ();
 sg13g2_fill_1 FILLER_42_2669 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_11 ();
 sg13g2_decap_8 FILLER_43_46 ();
 sg13g2_decap_8 FILLER_43_53 ();
 sg13g2_decap_8 FILLER_43_60 ();
 sg13g2_decap_8 FILLER_43_67 ();
 sg13g2_decap_8 FILLER_43_74 ();
 sg13g2_decap_8 FILLER_43_81 ();
 sg13g2_decap_8 FILLER_43_88 ();
 sg13g2_decap_8 FILLER_43_95 ();
 sg13g2_decap_8 FILLER_43_102 ();
 sg13g2_decap_4 FILLER_43_133 ();
 sg13g2_decap_4 FILLER_43_213 ();
 sg13g2_decap_4 FILLER_43_227 ();
 sg13g2_fill_2 FILLER_43_235 ();
 sg13g2_decap_8 FILLER_43_253 ();
 sg13g2_fill_1 FILLER_43_273 ();
 sg13g2_fill_2 FILLER_43_309 ();
 sg13g2_fill_1 FILLER_43_311 ();
 sg13g2_fill_2 FILLER_43_316 ();
 sg13g2_fill_1 FILLER_43_326 ();
 sg13g2_fill_2 FILLER_43_353 ();
 sg13g2_decap_8 FILLER_43_370 ();
 sg13g2_decap_4 FILLER_43_377 ();
 sg13g2_fill_1 FILLER_43_381 ();
 sg13g2_fill_1 FILLER_43_409 ();
 sg13g2_fill_2 FILLER_43_424 ();
 sg13g2_fill_1 FILLER_43_426 ();
 sg13g2_fill_1 FILLER_43_475 ();
 sg13g2_decap_8 FILLER_43_509 ();
 sg13g2_decap_8 FILLER_43_516 ();
 sg13g2_fill_2 FILLER_43_523 ();
 sg13g2_fill_2 FILLER_43_530 ();
 sg13g2_fill_2 FILLER_43_540 ();
 sg13g2_fill_1 FILLER_43_542 ();
 sg13g2_fill_1 FILLER_43_587 ();
 sg13g2_decap_8 FILLER_43_592 ();
 sg13g2_decap_8 FILLER_43_599 ();
 sg13g2_fill_1 FILLER_43_606 ();
 sg13g2_fill_2 FILLER_43_622 ();
 sg13g2_fill_1 FILLER_43_624 ();
 sg13g2_fill_2 FILLER_43_643 ();
 sg13g2_decap_8 FILLER_43_661 ();
 sg13g2_decap_8 FILLER_43_668 ();
 sg13g2_decap_8 FILLER_43_675 ();
 sg13g2_decap_8 FILLER_43_682 ();
 sg13g2_fill_2 FILLER_43_689 ();
 sg13g2_fill_1 FILLER_43_691 ();
 sg13g2_decap_8 FILLER_43_707 ();
 sg13g2_decap_8 FILLER_43_714 ();
 sg13g2_decap_4 FILLER_43_721 ();
 sg13g2_fill_2 FILLER_43_725 ();
 sg13g2_fill_2 FILLER_43_758 ();
 sg13g2_decap_8 FILLER_43_764 ();
 sg13g2_decap_8 FILLER_43_771 ();
 sg13g2_decap_8 FILLER_43_778 ();
 sg13g2_decap_8 FILLER_43_785 ();
 sg13g2_decap_4 FILLER_43_792 ();
 sg13g2_fill_2 FILLER_43_796 ();
 sg13g2_decap_8 FILLER_43_832 ();
 sg13g2_decap_8 FILLER_43_839 ();
 sg13g2_decap_8 FILLER_43_846 ();
 sg13g2_decap_8 FILLER_43_853 ();
 sg13g2_decap_8 FILLER_43_860 ();
 sg13g2_decap_8 FILLER_43_867 ();
 sg13g2_fill_2 FILLER_43_874 ();
 sg13g2_decap_8 FILLER_43_879 ();
 sg13g2_decap_8 FILLER_43_890 ();
 sg13g2_decap_8 FILLER_43_900 ();
 sg13g2_fill_2 FILLER_43_918 ();
 sg13g2_fill_1 FILLER_43_920 ();
 sg13g2_decap_8 FILLER_43_929 ();
 sg13g2_decap_8 FILLER_43_936 ();
 sg13g2_decap_8 FILLER_43_943 ();
 sg13g2_fill_2 FILLER_43_950 ();
 sg13g2_decap_8 FILLER_43_967 ();
 sg13g2_decap_8 FILLER_43_974 ();
 sg13g2_fill_2 FILLER_43_981 ();
 sg13g2_fill_1 FILLER_43_996 ();
 sg13g2_decap_8 FILLER_43_1001 ();
 sg13g2_decap_8 FILLER_43_1008 ();
 sg13g2_decap_8 FILLER_43_1015 ();
 sg13g2_decap_8 FILLER_43_1022 ();
 sg13g2_decap_4 FILLER_43_1029 ();
 sg13g2_fill_2 FILLER_43_1037 ();
 sg13g2_fill_1 FILLER_43_1039 ();
 sg13g2_decap_8 FILLER_43_1075 ();
 sg13g2_decap_4 FILLER_43_1082 ();
 sg13g2_decap_4 FILLER_43_1092 ();
 sg13g2_fill_2 FILLER_43_1096 ();
 sg13g2_fill_1 FILLER_43_1129 ();
 sg13g2_fill_2 FILLER_43_1140 ();
 sg13g2_fill_2 FILLER_43_1186 ();
 sg13g2_fill_2 FILLER_43_1227 ();
 sg13g2_fill_1 FILLER_43_1260 ();
 sg13g2_fill_1 FILLER_43_1267 ();
 sg13g2_fill_1 FILLER_43_1316 ();
 sg13g2_decap_8 FILLER_43_1325 ();
 sg13g2_decap_8 FILLER_43_1332 ();
 sg13g2_decap_4 FILLER_43_1339 ();
 sg13g2_decap_8 FILLER_43_1377 ();
 sg13g2_decap_8 FILLER_43_1384 ();
 sg13g2_fill_1 FILLER_43_1396 ();
 sg13g2_fill_1 FILLER_43_1401 ();
 sg13g2_decap_4 FILLER_43_1428 ();
 sg13g2_fill_2 FILLER_43_1432 ();
 sg13g2_fill_1 FILLER_43_1473 ();
 sg13g2_decap_4 FILLER_43_1480 ();
 sg13g2_decap_4 FILLER_43_1489 ();
 sg13g2_fill_2 FILLER_43_1497 ();
 sg13g2_fill_1 FILLER_43_1538 ();
 sg13g2_fill_2 FILLER_43_1551 ();
 sg13g2_decap_8 FILLER_43_1582 ();
 sg13g2_decap_8 FILLER_43_1589 ();
 sg13g2_fill_1 FILLER_43_1596 ();
 sg13g2_fill_1 FILLER_43_1602 ();
 sg13g2_fill_2 FILLER_43_1607 ();
 sg13g2_decap_8 FILLER_43_1613 ();
 sg13g2_decap_4 FILLER_43_1620 ();
 sg13g2_fill_1 FILLER_43_1624 ();
 sg13g2_fill_1 FILLER_43_1628 ();
 sg13g2_decap_4 FILLER_43_1638 ();
 sg13g2_fill_2 FILLER_43_1642 ();
 sg13g2_fill_2 FILLER_43_1647 ();
 sg13g2_fill_1 FILLER_43_1649 ();
 sg13g2_decap_8 FILLER_43_1656 ();
 sg13g2_decap_8 FILLER_43_1663 ();
 sg13g2_decap_8 FILLER_43_1670 ();
 sg13g2_decap_8 FILLER_43_1677 ();
 sg13g2_fill_2 FILLER_43_1684 ();
 sg13g2_fill_1 FILLER_43_1691 ();
 sg13g2_fill_2 FILLER_43_1725 ();
 sg13g2_fill_1 FILLER_43_1727 ();
 sg13g2_fill_1 FILLER_43_1741 ();
 sg13g2_fill_2 FILLER_43_1780 ();
 sg13g2_decap_8 FILLER_43_1795 ();
 sg13g2_decap_4 FILLER_43_1802 ();
 sg13g2_fill_1 FILLER_43_1806 ();
 sg13g2_decap_8 FILLER_43_1813 ();
 sg13g2_decap_8 FILLER_43_1820 ();
 sg13g2_decap_8 FILLER_43_1830 ();
 sg13g2_decap_4 FILLER_43_1846 ();
 sg13g2_fill_2 FILLER_43_1885 ();
 sg13g2_fill_1 FILLER_43_1910 ();
 sg13g2_fill_2 FILLER_43_1937 ();
 sg13g2_fill_2 FILLER_43_1953 ();
 sg13g2_fill_2 FILLER_43_1990 ();
 sg13g2_fill_1 FILLER_43_1992 ();
 sg13g2_fill_1 FILLER_43_1997 ();
 sg13g2_decap_4 FILLER_43_2029 ();
 sg13g2_fill_2 FILLER_43_2033 ();
 sg13g2_decap_4 FILLER_43_2040 ();
 sg13g2_fill_1 FILLER_43_2044 ();
 sg13g2_fill_1 FILLER_43_2071 ();
 sg13g2_decap_8 FILLER_43_2107 ();
 sg13g2_decap_4 FILLER_43_2114 ();
 sg13g2_fill_2 FILLER_43_2130 ();
 sg13g2_fill_1 FILLER_43_2141 ();
 sg13g2_decap_8 FILLER_43_2147 ();
 sg13g2_decap_8 FILLER_43_2154 ();
 sg13g2_decap_8 FILLER_43_2161 ();
 sg13g2_decap_8 FILLER_43_2168 ();
 sg13g2_decap_8 FILLER_43_2175 ();
 sg13g2_decap_8 FILLER_43_2182 ();
 sg13g2_fill_1 FILLER_43_2189 ();
 sg13g2_decap_4 FILLER_43_2199 ();
 sg13g2_fill_1 FILLER_43_2203 ();
 sg13g2_decap_4 FILLER_43_2230 ();
 sg13g2_fill_1 FILLER_43_2234 ();
 sg13g2_fill_2 FILLER_43_2244 ();
 sg13g2_decap_8 FILLER_43_2255 ();
 sg13g2_fill_1 FILLER_43_2262 ();
 sg13g2_decap_4 FILLER_43_2268 ();
 sg13g2_fill_1 FILLER_43_2272 ();
 sg13g2_decap_8 FILLER_43_2278 ();
 sg13g2_decap_8 FILLER_43_2285 ();
 sg13g2_decap_8 FILLER_43_2292 ();
 sg13g2_decap_4 FILLER_43_2335 ();
 sg13g2_fill_1 FILLER_43_2339 ();
 sg13g2_fill_2 FILLER_43_2350 ();
 sg13g2_fill_2 FILLER_43_2357 ();
 sg13g2_fill_2 FILLER_43_2363 ();
 sg13g2_fill_2 FILLER_43_2370 ();
 sg13g2_fill_1 FILLER_43_2377 ();
 sg13g2_fill_2 FILLER_43_2382 ();
 sg13g2_fill_1 FILLER_43_2384 ();
 sg13g2_fill_2 FILLER_43_2391 ();
 sg13g2_fill_1 FILLER_43_2393 ();
 sg13g2_fill_2 FILLER_43_2400 ();
 sg13g2_decap_4 FILLER_43_2419 ();
 sg13g2_fill_1 FILLER_43_2423 ();
 sg13g2_decap_8 FILLER_43_2429 ();
 sg13g2_decap_4 FILLER_43_2436 ();
 sg13g2_fill_2 FILLER_43_2445 ();
 sg13g2_fill_2 FILLER_43_2451 ();
 sg13g2_fill_1 FILLER_43_2453 ();
 sg13g2_decap_8 FILLER_43_2464 ();
 sg13g2_fill_2 FILLER_43_2471 ();
 sg13g2_fill_2 FILLER_43_2478 ();
 sg13g2_fill_1 FILLER_43_2480 ();
 sg13g2_fill_1 FILLER_43_2488 ();
 sg13g2_decap_8 FILLER_43_2493 ();
 sg13g2_decap_8 FILLER_43_2500 ();
 sg13g2_decap_8 FILLER_43_2507 ();
 sg13g2_decap_8 FILLER_43_2514 ();
 sg13g2_decap_4 FILLER_43_2521 ();
 sg13g2_fill_2 FILLER_43_2525 ();
 sg13g2_fill_2 FILLER_43_2592 ();
 sg13g2_fill_1 FILLER_43_2594 ();
 sg13g2_fill_1 FILLER_43_2600 ();
 sg13g2_decap_8 FILLER_43_2653 ();
 sg13g2_decap_8 FILLER_43_2660 ();
 sg13g2_fill_2 FILLER_43_2667 ();
 sg13g2_fill_1 FILLER_43_2669 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_decap_4 FILLER_44_47 ();
 sg13g2_decap_4 FILLER_44_128 ();
 sg13g2_decap_4 FILLER_44_136 ();
 sg13g2_fill_1 FILLER_44_140 ();
 sg13g2_fill_2 FILLER_44_159 ();
 sg13g2_fill_1 FILLER_44_177 ();
 sg13g2_fill_2 FILLER_44_207 ();
 sg13g2_decap_8 FILLER_44_213 ();
 sg13g2_decap_4 FILLER_44_220 ();
 sg13g2_fill_2 FILLER_44_228 ();
 sg13g2_fill_1 FILLER_44_230 ();
 sg13g2_fill_1 FILLER_44_235 ();
 sg13g2_decap_8 FILLER_44_244 ();
 sg13g2_decap_8 FILLER_44_251 ();
 sg13g2_fill_2 FILLER_44_258 ();
 sg13g2_fill_2 FILLER_44_268 ();
 sg13g2_fill_2 FILLER_44_296 ();
 sg13g2_decap_8 FILLER_44_303 ();
 sg13g2_fill_1 FILLER_44_314 ();
 sg13g2_fill_1 FILLER_44_319 ();
 sg13g2_fill_2 FILLER_44_324 ();
 sg13g2_fill_2 FILLER_44_330 ();
 sg13g2_decap_4 FILLER_44_335 ();
 sg13g2_fill_1 FILLER_44_339 ();
 sg13g2_fill_2 FILLER_44_352 ();
 sg13g2_fill_1 FILLER_44_359 ();
 sg13g2_decap_8 FILLER_44_369 ();
 sg13g2_decap_8 FILLER_44_376 ();
 sg13g2_decap_4 FILLER_44_387 ();
 sg13g2_fill_2 FILLER_44_395 ();
 sg13g2_fill_1 FILLER_44_397 ();
 sg13g2_decap_8 FILLER_44_452 ();
 sg13g2_fill_2 FILLER_44_459 ();
 sg13g2_fill_1 FILLER_44_461 ();
 sg13g2_fill_1 FILLER_44_472 ();
 sg13g2_decap_8 FILLER_44_504 ();
 sg13g2_decap_4 FILLER_44_511 ();
 sg13g2_fill_2 FILLER_44_515 ();
 sg13g2_fill_2 FILLER_44_521 ();
 sg13g2_fill_2 FILLER_44_541 ();
 sg13g2_fill_1 FILLER_44_547 ();
 sg13g2_decap_4 FILLER_44_556 ();
 sg13g2_fill_2 FILLER_44_560 ();
 sg13g2_fill_2 FILLER_44_567 ();
 sg13g2_fill_1 FILLER_44_569 ();
 sg13g2_decap_4 FILLER_44_574 ();
 sg13g2_fill_2 FILLER_44_578 ();
 sg13g2_fill_2 FILLER_44_586 ();
 sg13g2_fill_1 FILLER_44_588 ();
 sg13g2_decap_4 FILLER_44_594 ();
 sg13g2_fill_2 FILLER_44_598 ();
 sg13g2_fill_2 FILLER_44_610 ();
 sg13g2_fill_1 FILLER_44_621 ();
 sg13g2_fill_1 FILLER_44_645 ();
 sg13g2_decap_8 FILLER_44_659 ();
 sg13g2_fill_1 FILLER_44_666 ();
 sg13g2_decap_4 FILLER_44_684 ();
 sg13g2_fill_2 FILLER_44_688 ();
 sg13g2_decap_8 FILLER_44_705 ();
 sg13g2_decap_8 FILLER_44_712 ();
 sg13g2_decap_8 FILLER_44_719 ();
 sg13g2_decap_8 FILLER_44_726 ();
 sg13g2_decap_4 FILLER_44_733 ();
 sg13g2_decap_8 FILLER_44_781 ();
 sg13g2_decap_8 FILLER_44_788 ();
 sg13g2_decap_8 FILLER_44_795 ();
 sg13g2_decap_4 FILLER_44_802 ();
 sg13g2_fill_2 FILLER_44_806 ();
 sg13g2_decap_8 FILLER_44_816 ();
 sg13g2_fill_1 FILLER_44_823 ();
 sg13g2_decap_8 FILLER_44_830 ();
 sg13g2_fill_2 FILLER_44_837 ();
 sg13g2_fill_1 FILLER_44_839 ();
 sg13g2_fill_2 FILLER_44_845 ();
 sg13g2_fill_1 FILLER_44_847 ();
 sg13g2_decap_8 FILLER_44_861 ();
 sg13g2_fill_2 FILLER_44_868 ();
 sg13g2_fill_1 FILLER_44_870 ();
 sg13g2_fill_1 FILLER_44_876 ();
 sg13g2_fill_2 FILLER_44_916 ();
 sg13g2_decap_4 FILLER_44_935 ();
 sg13g2_fill_1 FILLER_44_952 ();
 sg13g2_fill_2 FILLER_44_1011 ();
 sg13g2_decap_8 FILLER_44_1023 ();
 sg13g2_decap_8 FILLER_44_1030 ();
 sg13g2_decap_8 FILLER_44_1037 ();
 sg13g2_decap_8 FILLER_44_1044 ();
 sg13g2_decap_4 FILLER_44_1051 ();
 sg13g2_fill_2 FILLER_44_1055 ();
 sg13g2_fill_2 FILLER_44_1088 ();
 sg13g2_fill_1 FILLER_44_1090 ();
 sg13g2_fill_2 FILLER_44_1117 ();
 sg13g2_fill_1 FILLER_44_1119 ();
 sg13g2_decap_8 FILLER_44_1150 ();
 sg13g2_fill_1 FILLER_44_1157 ();
 sg13g2_decap_8 FILLER_44_1162 ();
 sg13g2_decap_4 FILLER_44_1169 ();
 sg13g2_fill_2 FILLER_44_1173 ();
 sg13g2_decap_4 FILLER_44_1184 ();
 sg13g2_decap_8 FILLER_44_1192 ();
 sg13g2_fill_2 FILLER_44_1199 ();
 sg13g2_decap_8 FILLER_44_1205 ();
 sg13g2_decap_8 FILLER_44_1212 ();
 sg13g2_decap_8 FILLER_44_1219 ();
 sg13g2_fill_2 FILLER_44_1226 ();
 sg13g2_decap_8 FILLER_44_1233 ();
 sg13g2_decap_4 FILLER_44_1240 ();
 sg13g2_fill_1 FILLER_44_1244 ();
 sg13g2_decap_8 FILLER_44_1254 ();
 sg13g2_fill_2 FILLER_44_1261 ();
 sg13g2_fill_1 FILLER_44_1263 ();
 sg13g2_decap_8 FILLER_44_1301 ();
 sg13g2_decap_8 FILLER_44_1308 ();
 sg13g2_fill_2 FILLER_44_1315 ();
 sg13g2_fill_2 FILLER_44_1348 ();
 sg13g2_fill_2 FILLER_44_1359 ();
 sg13g2_fill_1 FILLER_44_1371 ();
 sg13g2_fill_2 FILLER_44_1398 ();
 sg13g2_fill_1 FILLER_44_1408 ();
 sg13g2_fill_2 FILLER_44_1414 ();
 sg13g2_fill_1 FILLER_44_1416 ();
 sg13g2_fill_2 FILLER_44_1425 ();
 sg13g2_decap_8 FILLER_44_1435 ();
 sg13g2_fill_2 FILLER_44_1442 ();
 sg13g2_fill_2 FILLER_44_1453 ();
 sg13g2_fill_1 FILLER_44_1455 ();
 sg13g2_decap_8 FILLER_44_1467 ();
 sg13g2_decap_8 FILLER_44_1474 ();
 sg13g2_fill_1 FILLER_44_1481 ();
 sg13g2_decap_4 FILLER_44_1516 ();
 sg13g2_fill_2 FILLER_44_1520 ();
 sg13g2_decap_4 FILLER_44_1528 ();
 sg13g2_fill_1 FILLER_44_1535 ();
 sg13g2_fill_2 FILLER_44_1551 ();
 sg13g2_fill_1 FILLER_44_1558 ();
 sg13g2_decap_8 FILLER_44_1573 ();
 sg13g2_decap_8 FILLER_44_1580 ();
 sg13g2_fill_2 FILLER_44_1613 ();
 sg13g2_fill_2 FILLER_44_1623 ();
 sg13g2_fill_2 FILLER_44_1628 ();
 sg13g2_decap_8 FILLER_44_1664 ();
 sg13g2_decap_8 FILLER_44_1671 ();
 sg13g2_decap_8 FILLER_44_1678 ();
 sg13g2_decap_4 FILLER_44_1685 ();
 sg13g2_decap_8 FILLER_44_1726 ();
 sg13g2_decap_4 FILLER_44_1733 ();
 sg13g2_fill_2 FILLER_44_1742 ();
 sg13g2_fill_1 FILLER_44_1775 ();
 sg13g2_fill_1 FILLER_44_1802 ();
 sg13g2_decap_4 FILLER_44_1810 ();
 sg13g2_fill_1 FILLER_44_1814 ();
 sg13g2_decap_8 FILLER_44_1853 ();
 sg13g2_decap_8 FILLER_44_1860 ();
 sg13g2_decap_8 FILLER_44_1867 ();
 sg13g2_decap_4 FILLER_44_1874 ();
 sg13g2_fill_1 FILLER_44_1878 ();
 sg13g2_fill_2 FILLER_44_1883 ();
 sg13g2_fill_1 FILLER_44_1894 ();
 sg13g2_fill_2 FILLER_44_1937 ();
 sg13g2_fill_1 FILLER_44_1943 ();
 sg13g2_decap_4 FILLER_44_1973 ();
 sg13g2_decap_8 FILLER_44_1986 ();
 sg13g2_decap_8 FILLER_44_1993 ();
 sg13g2_decap_8 FILLER_44_2000 ();
 sg13g2_fill_2 FILLER_44_2007 ();
 sg13g2_fill_1 FILLER_44_2022 ();
 sg13g2_fill_1 FILLER_44_2028 ();
 sg13g2_decap_8 FILLER_44_2033 ();
 sg13g2_decap_8 FILLER_44_2040 ();
 sg13g2_decap_8 FILLER_44_2047 ();
 sg13g2_decap_8 FILLER_44_2054 ();
 sg13g2_decap_8 FILLER_44_2061 ();
 sg13g2_decap_8 FILLER_44_2068 ();
 sg13g2_decap_4 FILLER_44_2075 ();
 sg13g2_fill_1 FILLER_44_2079 ();
 sg13g2_decap_8 FILLER_44_2101 ();
 sg13g2_decap_8 FILLER_44_2108 ();
 sg13g2_fill_2 FILLER_44_2115 ();
 sg13g2_fill_1 FILLER_44_2117 ();
 sg13g2_fill_1 FILLER_44_2127 ();
 sg13g2_decap_8 FILLER_44_2154 ();
 sg13g2_decap_8 FILLER_44_2161 ();
 sg13g2_decap_8 FILLER_44_2168 ();
 sg13g2_decap_8 FILLER_44_2175 ();
 sg13g2_decap_8 FILLER_44_2182 ();
 sg13g2_fill_1 FILLER_44_2189 ();
 sg13g2_decap_4 FILLER_44_2221 ();
 sg13g2_fill_1 FILLER_44_2231 ();
 sg13g2_decap_8 FILLER_44_2242 ();
 sg13g2_fill_1 FILLER_44_2249 ();
 sg13g2_fill_1 FILLER_44_2288 ();
 sg13g2_decap_4 FILLER_44_2295 ();
 sg13g2_fill_1 FILLER_44_2308 ();
 sg13g2_fill_1 FILLER_44_2315 ();
 sg13g2_fill_1 FILLER_44_2342 ();
 sg13g2_fill_1 FILLER_44_2348 ();
 sg13g2_fill_2 FILLER_44_2353 ();
 sg13g2_decap_8 FILLER_44_2361 ();
 sg13g2_decap_8 FILLER_44_2368 ();
 sg13g2_decap_8 FILLER_44_2375 ();
 sg13g2_decap_8 FILLER_44_2382 ();
 sg13g2_fill_2 FILLER_44_2389 ();
 sg13g2_fill_1 FILLER_44_2391 ();
 sg13g2_fill_1 FILLER_44_2397 ();
 sg13g2_decap_8 FILLER_44_2424 ();
 sg13g2_fill_2 FILLER_44_2435 ();
 sg13g2_fill_1 FILLER_44_2437 ();
 sg13g2_decap_8 FILLER_44_2527 ();
 sg13g2_decap_8 FILLER_44_2534 ();
 sg13g2_fill_2 FILLER_44_2544 ();
 sg13g2_decap_8 FILLER_44_2551 ();
 sg13g2_fill_2 FILLER_44_2558 ();
 sg13g2_fill_1 FILLER_44_2560 ();
 sg13g2_decap_4 FILLER_44_2565 ();
 sg13g2_decap_8 FILLER_44_2604 ();
 sg13g2_decap_8 FILLER_44_2611 ();
 sg13g2_decap_8 FILLER_44_2618 ();
 sg13g2_decap_8 FILLER_44_2625 ();
 sg13g2_decap_8 FILLER_44_2632 ();
 sg13g2_decap_8 FILLER_44_2639 ();
 sg13g2_decap_8 FILLER_44_2646 ();
 sg13g2_decap_8 FILLER_44_2653 ();
 sg13g2_decap_8 FILLER_44_2660 ();
 sg13g2_fill_2 FILLER_44_2667 ();
 sg13g2_fill_1 FILLER_44_2669 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_26 ();
 sg13g2_decap_8 FILLER_45_33 ();
 sg13g2_decap_8 FILLER_45_40 ();
 sg13g2_fill_1 FILLER_45_47 ();
 sg13g2_decap_4 FILLER_45_52 ();
 sg13g2_decap_8 FILLER_45_82 ();
 sg13g2_decap_8 FILLER_45_89 ();
 sg13g2_fill_2 FILLER_45_96 ();
 sg13g2_fill_2 FILLER_45_140 ();
 sg13g2_fill_1 FILLER_45_142 ();
 sg13g2_fill_2 FILLER_45_153 ();
 sg13g2_fill_1 FILLER_45_163 ();
 sg13g2_fill_2 FILLER_45_172 ();
 sg13g2_fill_1 FILLER_45_179 ();
 sg13g2_fill_1 FILLER_45_185 ();
 sg13g2_fill_2 FILLER_45_203 ();
 sg13g2_fill_2 FILLER_45_240 ();
 sg13g2_fill_1 FILLER_45_242 ();
 sg13g2_fill_2 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_fill_2 FILLER_45_308 ();
 sg13g2_fill_2 FILLER_45_315 ();
 sg13g2_fill_1 FILLER_45_325 ();
 sg13g2_decap_4 FILLER_45_329 ();
 sg13g2_fill_1 FILLER_45_333 ();
 sg13g2_decap_4 FILLER_45_340 ();
 sg13g2_fill_2 FILLER_45_344 ();
 sg13g2_decap_8 FILLER_45_352 ();
 sg13g2_decap_8 FILLER_45_359 ();
 sg13g2_fill_2 FILLER_45_366 ();
 sg13g2_fill_1 FILLER_45_368 ();
 sg13g2_decap_4 FILLER_45_372 ();
 sg13g2_fill_1 FILLER_45_402 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_decap_8 FILLER_45_422 ();
 sg13g2_decap_8 FILLER_45_429 ();
 sg13g2_decap_4 FILLER_45_436 ();
 sg13g2_fill_1 FILLER_45_440 ();
 sg13g2_fill_1 FILLER_45_444 ();
 sg13g2_decap_8 FILLER_45_450 ();
 sg13g2_fill_2 FILLER_45_457 ();
 sg13g2_fill_1 FILLER_45_509 ();
 sg13g2_decap_4 FILLER_45_515 ();
 sg13g2_fill_2 FILLER_45_519 ();
 sg13g2_decap_4 FILLER_45_551 ();
 sg13g2_fill_1 FILLER_45_555 ();
 sg13g2_decap_4 FILLER_45_559 ();
 sg13g2_fill_1 FILLER_45_563 ();
 sg13g2_decap_8 FILLER_45_594 ();
 sg13g2_decap_4 FILLER_45_601 ();
 sg13g2_decap_8 FILLER_45_617 ();
 sg13g2_fill_1 FILLER_45_624 ();
 sg13g2_fill_2 FILLER_45_634 ();
 sg13g2_fill_1 FILLER_45_636 ();
 sg13g2_decap_8 FILLER_45_651 ();
 sg13g2_decap_8 FILLER_45_658 ();
 sg13g2_decap_4 FILLER_45_665 ();
 sg13g2_fill_1 FILLER_45_669 ();
 sg13g2_fill_2 FILLER_45_676 ();
 sg13g2_fill_1 FILLER_45_678 ();
 sg13g2_decap_4 FILLER_45_684 ();
 sg13g2_fill_2 FILLER_45_688 ();
 sg13g2_fill_1 FILLER_45_695 ();
 sg13g2_fill_2 FILLER_45_701 ();
 sg13g2_fill_2 FILLER_45_708 ();
 sg13g2_decap_4 FILLER_45_727 ();
 sg13g2_fill_2 FILLER_45_734 ();
 sg13g2_decap_8 FILLER_45_739 ();
 sg13g2_decap_4 FILLER_45_750 ();
 sg13g2_decap_8 FILLER_45_758 ();
 sg13g2_fill_2 FILLER_45_765 ();
 sg13g2_fill_1 FILLER_45_767 ();
 sg13g2_decap_8 FILLER_45_773 ();
 sg13g2_fill_1 FILLER_45_780 ();
 sg13g2_fill_2 FILLER_45_786 ();
 sg13g2_decap_8 FILLER_45_795 ();
 sg13g2_decap_8 FILLER_45_802 ();
 sg13g2_decap_8 FILLER_45_809 ();
 sg13g2_decap_8 FILLER_45_816 ();
 sg13g2_decap_8 FILLER_45_823 ();
 sg13g2_fill_2 FILLER_45_830 ();
 sg13g2_fill_1 FILLER_45_832 ();
 sg13g2_decap_8 FILLER_45_838 ();
 sg13g2_fill_2 FILLER_45_845 ();
 sg13g2_fill_1 FILLER_45_847 ();
 sg13g2_fill_1 FILLER_45_854 ();
 sg13g2_fill_2 FILLER_45_861 ();
 sg13g2_fill_1 FILLER_45_863 ();
 sg13g2_fill_2 FILLER_45_879 ();
 sg13g2_fill_1 FILLER_45_881 ();
 sg13g2_decap_4 FILLER_45_887 ();
 sg13g2_fill_2 FILLER_45_891 ();
 sg13g2_fill_2 FILLER_45_905 ();
 sg13g2_fill_1 FILLER_45_907 ();
 sg13g2_decap_8 FILLER_45_924 ();
 sg13g2_decap_8 FILLER_45_931 ();
 sg13g2_fill_2 FILLER_45_938 ();
 sg13g2_fill_1 FILLER_45_940 ();
 sg13g2_decap_8 FILLER_45_946 ();
 sg13g2_fill_2 FILLER_45_953 ();
 sg13g2_decap_4 FILLER_45_964 ();
 sg13g2_fill_1 FILLER_45_968 ();
 sg13g2_decap_4 FILLER_45_979 ();
 sg13g2_decap_8 FILLER_45_988 ();
 sg13g2_fill_2 FILLER_45_1004 ();
 sg13g2_decap_8 FILLER_45_1032 ();
 sg13g2_decap_8 FILLER_45_1039 ();
 sg13g2_decap_8 FILLER_45_1046 ();
 sg13g2_decap_8 FILLER_45_1053 ();
 sg13g2_decap_8 FILLER_45_1060 ();
 sg13g2_decap_8 FILLER_45_1067 ();
 sg13g2_decap_8 FILLER_45_1074 ();
 sg13g2_decap_8 FILLER_45_1081 ();
 sg13g2_decap_8 FILLER_45_1088 ();
 sg13g2_decap_4 FILLER_45_1095 ();
 sg13g2_fill_2 FILLER_45_1099 ();
 sg13g2_fill_1 FILLER_45_1113 ();
 sg13g2_decap_8 FILLER_45_1127 ();
 sg13g2_decap_4 FILLER_45_1134 ();
 sg13g2_fill_1 FILLER_45_1138 ();
 sg13g2_decap_4 FILLER_45_1143 ();
 sg13g2_fill_1 FILLER_45_1147 ();
 sg13g2_decap_8 FILLER_45_1152 ();
 sg13g2_decap_4 FILLER_45_1159 ();
 sg13g2_fill_2 FILLER_45_1163 ();
 sg13g2_decap_4 FILLER_45_1173 ();
 sg13g2_fill_2 FILLER_45_1177 ();
 sg13g2_decap_8 FILLER_45_1199 ();
 sg13g2_decap_8 FILLER_45_1206 ();
 sg13g2_fill_2 FILLER_45_1213 ();
 sg13g2_fill_1 FILLER_45_1215 ();
 sg13g2_decap_8 FILLER_45_1229 ();
 sg13g2_fill_2 FILLER_45_1236 ();
 sg13g2_fill_1 FILLER_45_1238 ();
 sg13g2_decap_8 FILLER_45_1245 ();
 sg13g2_decap_8 FILLER_45_1252 ();
 sg13g2_decap_4 FILLER_45_1259 ();
 sg13g2_decap_8 FILLER_45_1307 ();
 sg13g2_fill_1 FILLER_45_1314 ();
 sg13g2_decap_8 FILLER_45_1319 ();
 sg13g2_decap_8 FILLER_45_1326 ();
 sg13g2_fill_2 FILLER_45_1350 ();
 sg13g2_decap_4 FILLER_45_1381 ();
 sg13g2_fill_2 FILLER_45_1407 ();
 sg13g2_fill_1 FILLER_45_1409 ();
 sg13g2_fill_2 FILLER_45_1418 ();
 sg13g2_fill_1 FILLER_45_1420 ();
 sg13g2_decap_4 FILLER_45_1425 ();
 sg13g2_fill_2 FILLER_45_1429 ();
 sg13g2_fill_2 FILLER_45_1467 ();
 sg13g2_decap_8 FILLER_45_1475 ();
 sg13g2_decap_4 FILLER_45_1482 ();
 sg13g2_fill_1 FILLER_45_1486 ();
 sg13g2_decap_8 FILLER_45_1493 ();
 sg13g2_decap_8 FILLER_45_1500 ();
 sg13g2_fill_2 FILLER_45_1507 ();
 sg13g2_fill_1 FILLER_45_1509 ();
 sg13g2_decap_8 FILLER_45_1515 ();
 sg13g2_decap_8 FILLER_45_1522 ();
 sg13g2_decap_4 FILLER_45_1529 ();
 sg13g2_fill_2 FILLER_45_1533 ();
 sg13g2_fill_2 FILLER_45_1561 ();
 sg13g2_fill_2 FILLER_45_1620 ();
 sg13g2_fill_1 FILLER_45_1637 ();
 sg13g2_decap_8 FILLER_45_1687 ();
 sg13g2_decap_8 FILLER_45_1694 ();
 sg13g2_decap_8 FILLER_45_1733 ();
 sg13g2_fill_1 FILLER_45_1740 ();
 sg13g2_decap_8 FILLER_45_1747 ();
 sg13g2_fill_1 FILLER_45_1754 ();
 sg13g2_decap_8 FILLER_45_1775 ();
 sg13g2_decap_4 FILLER_45_1782 ();
 sg13g2_fill_2 FILLER_45_1786 ();
 sg13g2_fill_2 FILLER_45_1792 ();
 sg13g2_fill_1 FILLER_45_1794 ();
 sg13g2_decap_4 FILLER_45_1800 ();
 sg13g2_fill_2 FILLER_45_1804 ();
 sg13g2_fill_2 FILLER_45_1825 ();
 sg13g2_decap_8 FILLER_45_1860 ();
 sg13g2_fill_2 FILLER_45_1867 ();
 sg13g2_fill_1 FILLER_45_1869 ();
 sg13g2_fill_2 FILLER_45_1875 ();
 sg13g2_fill_2 FILLER_45_1887 ();
 sg13g2_fill_2 FILLER_45_1902 ();
 sg13g2_decap_8 FILLER_45_1953 ();
 sg13g2_decap_8 FILLER_45_1960 ();
 sg13g2_decap_4 FILLER_45_1967 ();
 sg13g2_fill_1 FILLER_45_1971 ();
 sg13g2_decap_4 FILLER_45_1981 ();
 sg13g2_fill_1 FILLER_45_2019 ();
 sg13g2_decap_8 FILLER_45_2046 ();
 sg13g2_fill_2 FILLER_45_2053 ();
 sg13g2_fill_1 FILLER_45_2055 ();
 sg13g2_decap_8 FILLER_45_2061 ();
 sg13g2_fill_2 FILLER_45_2085 ();
 sg13g2_fill_1 FILLER_45_2087 ();
 sg13g2_fill_1 FILLER_45_2119 ();
 sg13g2_fill_1 FILLER_45_2146 ();
 sg13g2_fill_1 FILLER_45_2153 ();
 sg13g2_fill_1 FILLER_45_2158 ();
 sg13g2_fill_1 FILLER_45_2165 ();
 sg13g2_decap_4 FILLER_45_2171 ();
 sg13g2_fill_1 FILLER_45_2175 ();
 sg13g2_decap_8 FILLER_45_2202 ();
 sg13g2_decap_8 FILLER_45_2209 ();
 sg13g2_decap_8 FILLER_45_2216 ();
 sg13g2_decap_8 FILLER_45_2249 ();
 sg13g2_decap_8 FILLER_45_2256 ();
 sg13g2_decap_8 FILLER_45_2263 ();
 sg13g2_decap_4 FILLER_45_2270 ();
 sg13g2_fill_2 FILLER_45_2274 ();
 sg13g2_fill_1 FILLER_45_2302 ();
 sg13g2_decap_8 FILLER_45_2310 ();
 sg13g2_decap_8 FILLER_45_2317 ();
 sg13g2_fill_1 FILLER_45_2324 ();
 sg13g2_fill_2 FILLER_45_2337 ();
 sg13g2_fill_1 FILLER_45_2339 ();
 sg13g2_decap_8 FILLER_45_2371 ();
 sg13g2_decap_8 FILLER_45_2378 ();
 sg13g2_fill_1 FILLER_45_2385 ();
 sg13g2_decap_8 FILLER_45_2395 ();
 sg13g2_decap_8 FILLER_45_2408 ();
 sg13g2_fill_2 FILLER_45_2415 ();
 sg13g2_fill_1 FILLER_45_2417 ();
 sg13g2_fill_1 FILLER_45_2453 ();
 sg13g2_fill_2 FILLER_45_2458 ();
 sg13g2_fill_1 FILLER_45_2460 ();
 sg13g2_decap_8 FILLER_45_2478 ();
 sg13g2_decap_4 FILLER_45_2485 ();
 sg13g2_decap_8 FILLER_45_2492 ();
 sg13g2_fill_2 FILLER_45_2499 ();
 sg13g2_fill_2 FILLER_45_2506 ();
 sg13g2_decap_4 FILLER_45_2512 ();
 sg13g2_fill_1 FILLER_45_2516 ();
 sg13g2_decap_8 FILLER_45_2523 ();
 sg13g2_decap_8 FILLER_45_2530 ();
 sg13g2_decap_4 FILLER_45_2537 ();
 sg13g2_decap_4 FILLER_45_2554 ();
 sg13g2_fill_1 FILLER_45_2558 ();
 sg13g2_decap_8 FILLER_45_2563 ();
 sg13g2_fill_2 FILLER_45_2570 ();
 sg13g2_fill_1 FILLER_45_2572 ();
 sg13g2_decap_8 FILLER_45_2603 ();
 sg13g2_decap_4 FILLER_45_2610 ();
 sg13g2_fill_2 FILLER_45_2614 ();
 sg13g2_decap_8 FILLER_45_2646 ();
 sg13g2_decap_8 FILLER_45_2653 ();
 sg13g2_decap_8 FILLER_45_2660 ();
 sg13g2_fill_2 FILLER_45_2667 ();
 sg13g2_fill_1 FILLER_45_2669 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_30 ();
 sg13g2_decap_8 FILLER_46_37 ();
 sg13g2_fill_2 FILLER_46_44 ();
 sg13g2_fill_1 FILLER_46_46 ();
 sg13g2_fill_2 FILLER_46_59 ();
 sg13g2_decap_4 FILLER_46_91 ();
 sg13g2_fill_1 FILLER_46_95 ();
 sg13g2_decap_4 FILLER_46_132 ();
 sg13g2_fill_2 FILLER_46_136 ();
 sg13g2_decap_8 FILLER_46_222 ();
 sg13g2_decap_4 FILLER_46_229 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_fill_2 FILLER_46_245 ();
 sg13g2_fill_1 FILLER_46_247 ();
 sg13g2_fill_2 FILLER_46_251 ();
 sg13g2_fill_2 FILLER_46_265 ();
 sg13g2_decap_8 FILLER_46_270 ();
 sg13g2_fill_2 FILLER_46_277 ();
 sg13g2_decap_4 FILLER_46_308 ();
 sg13g2_decap_4 FILLER_46_316 ();
 sg13g2_fill_1 FILLER_46_320 ();
 sg13g2_decap_4 FILLER_46_352 ();
 sg13g2_fill_1 FILLER_46_359 ();
 sg13g2_decap_8 FILLER_46_398 ();
 sg13g2_fill_2 FILLER_46_410 ();
 sg13g2_fill_1 FILLER_46_412 ();
 sg13g2_decap_8 FILLER_46_416 ();
 sg13g2_decap_8 FILLER_46_423 ();
 sg13g2_fill_2 FILLER_46_430 ();
 sg13g2_fill_1 FILLER_46_471 ();
 sg13g2_fill_2 FILLER_46_482 ();
 sg13g2_fill_2 FILLER_46_489 ();
 sg13g2_fill_1 FILLER_46_496 ();
 sg13g2_fill_2 FILLER_46_508 ();
 sg13g2_decap_4 FILLER_46_515 ();
 sg13g2_decap_8 FILLER_46_550 ();
 sg13g2_decap_8 FILLER_46_557 ();
 sg13g2_fill_2 FILLER_46_569 ();
 sg13g2_decap_8 FILLER_46_575 ();
 sg13g2_decap_8 FILLER_46_582 ();
 sg13g2_decap_4 FILLER_46_589 ();
 sg13g2_fill_2 FILLER_46_593 ();
 sg13g2_decap_8 FILLER_46_600 ();
 sg13g2_decap_8 FILLER_46_607 ();
 sg13g2_decap_4 FILLER_46_614 ();
 sg13g2_decap_8 FILLER_46_623 ();
 sg13g2_decap_8 FILLER_46_630 ();
 sg13g2_decap_4 FILLER_46_637 ();
 sg13g2_fill_1 FILLER_46_641 ();
 sg13g2_decap_4 FILLER_46_661 ();
 sg13g2_fill_2 FILLER_46_712 ();
 sg13g2_fill_1 FILLER_46_714 ();
 sg13g2_decap_4 FILLER_46_719 ();
 sg13g2_fill_2 FILLER_46_731 ();
 sg13g2_decap_8 FILLER_46_742 ();
 sg13g2_decap_4 FILLER_46_749 ();
 sg13g2_fill_1 FILLER_46_792 ();
 sg13g2_fill_2 FILLER_46_811 ();
 sg13g2_fill_1 FILLER_46_827 ();
 sg13g2_fill_2 FILLER_46_832 ();
 sg13g2_decap_4 FILLER_46_844 ();
 sg13g2_decap_8 FILLER_46_865 ();
 sg13g2_fill_2 FILLER_46_872 ();
 sg13g2_fill_1 FILLER_46_874 ();
 sg13g2_decap_4 FILLER_46_888 ();
 sg13g2_decap_8 FILLER_46_906 ();
 sg13g2_decap_8 FILLER_46_913 ();
 sg13g2_fill_2 FILLER_46_930 ();
 sg13g2_fill_1 FILLER_46_932 ();
 sg13g2_decap_4 FILLER_46_945 ();
 sg13g2_fill_2 FILLER_46_949 ();
 sg13g2_fill_2 FILLER_46_965 ();
 sg13g2_fill_1 FILLER_46_967 ();
 sg13g2_decap_8 FILLER_46_980 ();
 sg13g2_decap_4 FILLER_46_987 ();
 sg13g2_fill_2 FILLER_46_996 ();
 sg13g2_fill_1 FILLER_46_998 ();
 sg13g2_fill_2 FILLER_46_1014 ();
 sg13g2_decap_4 FILLER_46_1020 ();
 sg13g2_decap_8 FILLER_46_1034 ();
 sg13g2_fill_2 FILLER_46_1041 ();
 sg13g2_fill_1 FILLER_46_1043 ();
 sg13g2_decap_4 FILLER_46_1048 ();
 sg13g2_decap_8 FILLER_46_1056 ();
 sg13g2_fill_2 FILLER_46_1068 ();
 sg13g2_fill_1 FILLER_46_1070 ();
 sg13g2_fill_2 FILLER_46_1081 ();
 sg13g2_fill_1 FILLER_46_1083 ();
 sg13g2_decap_8 FILLER_46_1088 ();
 sg13g2_decap_8 FILLER_46_1095 ();
 sg13g2_decap_4 FILLER_46_1102 ();
 sg13g2_fill_1 FILLER_46_1106 ();
 sg13g2_decap_8 FILLER_46_1220 ();
 sg13g2_fill_2 FILLER_46_1227 ();
 sg13g2_fill_1 FILLER_46_1229 ();
 sg13g2_decap_8 FILLER_46_1248 ();
 sg13g2_decap_8 FILLER_46_1255 ();
 sg13g2_decap_4 FILLER_46_1301 ();
 sg13g2_fill_2 FILLER_46_1315 ();
 sg13g2_fill_1 FILLER_46_1322 ();
 sg13g2_decap_8 FILLER_46_1329 ();
 sg13g2_decap_4 FILLER_46_1336 ();
 sg13g2_fill_1 FILLER_46_1340 ();
 sg13g2_fill_1 FILLER_46_1346 ();
 sg13g2_fill_1 FILLER_46_1351 ();
 sg13g2_fill_1 FILLER_46_1358 ();
 sg13g2_fill_1 FILLER_46_1385 ();
 sg13g2_fill_2 FILLER_46_1399 ();
 sg13g2_decap_8 FILLER_46_1413 ();
 sg13g2_decap_8 FILLER_46_1420 ();
 sg13g2_fill_2 FILLER_46_1427 ();
 sg13g2_decap_8 FILLER_46_1439 ();
 sg13g2_fill_2 FILLER_46_1446 ();
 sg13g2_fill_1 FILLER_46_1448 ();
 sg13g2_fill_1 FILLER_46_1459 ();
 sg13g2_decap_4 FILLER_46_1468 ();
 sg13g2_decap_8 FILLER_46_1502 ();
 sg13g2_decap_8 FILLER_46_1509 ();
 sg13g2_decap_4 FILLER_46_1516 ();
 sg13g2_fill_1 FILLER_46_1520 ();
 sg13g2_decap_8 FILLER_46_1527 ();
 sg13g2_decap_8 FILLER_46_1534 ();
 sg13g2_decap_4 FILLER_46_1541 ();
 sg13g2_fill_2 FILLER_46_1553 ();
 sg13g2_fill_1 FILLER_46_1559 ();
 sg13g2_fill_1 FILLER_46_1586 ();
 sg13g2_decap_4 FILLER_46_1593 ();
 sg13g2_fill_2 FILLER_46_1597 ();
 sg13g2_fill_2 FILLER_46_1611 ();
 sg13g2_fill_1 FILLER_46_1613 ();
 sg13g2_fill_1 FILLER_46_1640 ();
 sg13g2_fill_2 FILLER_46_1673 ();
 sg13g2_fill_2 FILLER_46_1699 ();
 sg13g2_fill_1 FILLER_46_1705 ();
 sg13g2_decap_4 FILLER_46_1732 ();
 sg13g2_decap_4 FILLER_46_1762 ();
 sg13g2_fill_1 FILLER_46_1798 ();
 sg13g2_decap_8 FILLER_46_1804 ();
 sg13g2_decap_8 FILLER_46_1811 ();
 sg13g2_fill_2 FILLER_46_1822 ();
 sg13g2_fill_2 FILLER_46_1841 ();
 sg13g2_fill_1 FILLER_46_1843 ();
 sg13g2_decap_8 FILLER_46_1848 ();
 sg13g2_decap_8 FILLER_46_1855 ();
 sg13g2_decap_8 FILLER_46_1862 ();
 sg13g2_decap_4 FILLER_46_1869 ();
 sg13g2_fill_1 FILLER_46_1873 ();
 sg13g2_decap_8 FILLER_46_1883 ();
 sg13g2_decap_4 FILLER_46_1890 ();
 sg13g2_fill_2 FILLER_46_1899 ();
 sg13g2_fill_2 FILLER_46_1940 ();
 sg13g2_fill_1 FILLER_46_1949 ();
 sg13g2_decap_8 FILLER_46_1954 ();
 sg13g2_decap_8 FILLER_46_1961 ();
 sg13g2_fill_2 FILLER_46_1968 ();
 sg13g2_fill_1 FILLER_46_1970 ();
 sg13g2_fill_2 FILLER_46_1976 ();
 sg13g2_fill_1 FILLER_46_1978 ();
 sg13g2_fill_2 FILLER_46_2016 ();
 sg13g2_fill_1 FILLER_46_2044 ();
 sg13g2_fill_1 FILLER_46_2130 ();
 sg13g2_fill_2 FILLER_46_2162 ();
 sg13g2_fill_1 FILLER_46_2164 ();
 sg13g2_decap_8 FILLER_46_2169 ();
 sg13g2_fill_1 FILLER_46_2176 ();
 sg13g2_decap_8 FILLER_46_2181 ();
 sg13g2_fill_2 FILLER_46_2188 ();
 sg13g2_fill_1 FILLER_46_2190 ();
 sg13g2_decap_8 FILLER_46_2195 ();
 sg13g2_decap_8 FILLER_46_2202 ();
 sg13g2_decap_8 FILLER_46_2209 ();
 sg13g2_fill_2 FILLER_46_2216 ();
 sg13g2_fill_1 FILLER_46_2218 ();
 sg13g2_decap_8 FILLER_46_2224 ();
 sg13g2_fill_1 FILLER_46_2231 ();
 sg13g2_decap_8 FILLER_46_2244 ();
 sg13g2_decap_4 FILLER_46_2251 ();
 sg13g2_fill_2 FILLER_46_2255 ();
 sg13g2_fill_2 FILLER_46_2300 ();
 sg13g2_decap_8 FILLER_46_2307 ();
 sg13g2_decap_8 FILLER_46_2314 ();
 sg13g2_decap_8 FILLER_46_2321 ();
 sg13g2_fill_1 FILLER_46_2328 ();
 sg13g2_fill_2 FILLER_46_2334 ();
 sg13g2_fill_2 FILLER_46_2340 ();
 sg13g2_fill_2 FILLER_46_2346 ();
 sg13g2_fill_1 FILLER_46_2348 ();
 sg13g2_decap_8 FILLER_46_2379 ();
 sg13g2_decap_8 FILLER_46_2412 ();
 sg13g2_fill_1 FILLER_46_2419 ();
 sg13g2_fill_1 FILLER_46_2446 ();
 sg13g2_fill_2 FILLER_46_2479 ();
 sg13g2_decap_8 FILLER_46_2495 ();
 sg13g2_fill_2 FILLER_46_2502 ();
 sg13g2_fill_1 FILLER_46_2504 ();
 sg13g2_fill_2 FILLER_46_2541 ();
 sg13g2_fill_1 FILLER_46_2543 ();
 sg13g2_decap_8 FILLER_46_2570 ();
 sg13g2_decap_8 FILLER_46_2577 ();
 sg13g2_decap_4 FILLER_46_2584 ();
 sg13g2_decap_8 FILLER_46_2593 ();
 sg13g2_decap_8 FILLER_46_2600 ();
 sg13g2_decap_8 FILLER_46_2607 ();
 sg13g2_decap_8 FILLER_46_2614 ();
 sg13g2_decap_8 FILLER_46_2621 ();
 sg13g2_fill_2 FILLER_46_2628 ();
 sg13g2_fill_1 FILLER_46_2630 ();
 sg13g2_decap_8 FILLER_46_2635 ();
 sg13g2_decap_8 FILLER_46_2642 ();
 sg13g2_decap_8 FILLER_46_2649 ();
 sg13g2_decap_8 FILLER_46_2656 ();
 sg13g2_decap_8 FILLER_46_2663 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_11 ();
 sg13g2_fill_2 FILLER_47_30 ();
 sg13g2_decap_4 FILLER_47_38 ();
 sg13g2_fill_1 FILLER_47_42 ();
 sg13g2_decap_4 FILLER_47_74 ();
 sg13g2_decap_8 FILLER_47_86 ();
 sg13g2_decap_8 FILLER_47_93 ();
 sg13g2_decap_8 FILLER_47_104 ();
 sg13g2_decap_4 FILLER_47_111 ();
 sg13g2_fill_2 FILLER_47_115 ();
 sg13g2_decap_8 FILLER_47_143 ();
 sg13g2_decap_8 FILLER_47_150 ();
 sg13g2_decap_8 FILLER_47_157 ();
 sg13g2_decap_8 FILLER_47_164 ();
 sg13g2_fill_2 FILLER_47_174 ();
 sg13g2_fill_1 FILLER_47_176 ();
 sg13g2_decap_4 FILLER_47_221 ();
 sg13g2_fill_2 FILLER_47_225 ();
 sg13g2_decap_4 FILLER_47_234 ();
 sg13g2_fill_1 FILLER_47_238 ();
 sg13g2_fill_1 FILLER_47_242 ();
 sg13g2_decap_8 FILLER_47_269 ();
 sg13g2_decap_8 FILLER_47_276 ();
 sg13g2_fill_1 FILLER_47_283 ();
 sg13g2_fill_1 FILLER_47_363 ();
 sg13g2_fill_1 FILLER_47_377 ();
 sg13g2_decap_8 FILLER_47_443 ();
 sg13g2_decap_4 FILLER_47_450 ();
 sg13g2_fill_1 FILLER_47_458 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_fill_1 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_482 ();
 sg13g2_decap_8 FILLER_47_489 ();
 sg13g2_decap_8 FILLER_47_496 ();
 sg13g2_decap_8 FILLER_47_503 ();
 sg13g2_decap_8 FILLER_47_510 ();
 sg13g2_fill_1 FILLER_47_517 ();
 sg13g2_fill_2 FILLER_47_527 ();
 sg13g2_fill_1 FILLER_47_529 ();
 sg13g2_fill_1 FILLER_47_535 ();
 sg13g2_decap_8 FILLER_47_540 ();
 sg13g2_fill_2 FILLER_47_547 ();
 sg13g2_fill_1 FILLER_47_554 ();
 sg13g2_fill_2 FILLER_47_559 ();
 sg13g2_fill_1 FILLER_47_566 ();
 sg13g2_decap_8 FILLER_47_574 ();
 sg13g2_fill_1 FILLER_47_581 ();
 sg13g2_decap_8 FILLER_47_587 ();
 sg13g2_fill_2 FILLER_47_594 ();
 sg13g2_decap_8 FILLER_47_606 ();
 sg13g2_decap_8 FILLER_47_613 ();
 sg13g2_fill_2 FILLER_47_620 ();
 sg13g2_fill_2 FILLER_47_661 ();
 sg13g2_fill_2 FILLER_47_687 ();
 sg13g2_fill_2 FILLER_47_694 ();
 sg13g2_fill_2 FILLER_47_701 ();
 sg13g2_fill_1 FILLER_47_703 ();
 sg13g2_decap_8 FILLER_47_712 ();
 sg13g2_fill_1 FILLER_47_724 ();
 sg13g2_decap_4 FILLER_47_730 ();
 sg13g2_decap_8 FILLER_47_738 ();
 sg13g2_decap_8 FILLER_47_745 ();
 sg13g2_fill_2 FILLER_47_752 ();
 sg13g2_fill_1 FILLER_47_754 ();
 sg13g2_decap_8 FILLER_47_760 ();
 sg13g2_decap_8 FILLER_47_767 ();
 sg13g2_decap_8 FILLER_47_779 ();
 sg13g2_fill_2 FILLER_47_786 ();
 sg13g2_fill_1 FILLER_47_788 ();
 sg13g2_fill_2 FILLER_47_799 ();
 sg13g2_decap_4 FILLER_47_806 ();
 sg13g2_fill_1 FILLER_47_810 ();
 sg13g2_decap_8 FILLER_47_821 ();
 sg13g2_fill_1 FILLER_47_828 ();
 sg13g2_decap_8 FILLER_47_838 ();
 sg13g2_decap_4 FILLER_47_845 ();
 sg13g2_decap_8 FILLER_47_853 ();
 sg13g2_decap_4 FILLER_47_860 ();
 sg13g2_fill_1 FILLER_47_869 ();
 sg13g2_fill_2 FILLER_47_897 ();
 sg13g2_fill_1 FILLER_47_899 ();
 sg13g2_decap_8 FILLER_47_921 ();
 sg13g2_fill_1 FILLER_47_928 ();
 sg13g2_fill_1 FILLER_47_949 ();
 sg13g2_fill_1 FILLER_47_967 ();
 sg13g2_fill_1 FILLER_47_973 ();
 sg13g2_fill_1 FILLER_47_978 ();
 sg13g2_fill_1 FILLER_47_983 ();
 sg13g2_fill_2 FILLER_47_997 ();
 sg13g2_fill_1 FILLER_47_1003 ();
 sg13g2_fill_2 FILLER_47_1009 ();
 sg13g2_fill_1 FILLER_47_1018 ();
 sg13g2_fill_2 FILLER_47_1033 ();
 sg13g2_fill_1 FILLER_47_1035 ();
 sg13g2_fill_2 FILLER_47_1062 ();
 sg13g2_decap_8 FILLER_47_1119 ();
 sg13g2_fill_1 FILLER_47_1126 ();
 sg13g2_fill_1 FILLER_47_1152 ();
 sg13g2_fill_2 FILLER_47_1160 ();
 sg13g2_fill_1 FILLER_47_1162 ();
 sg13g2_decap_8 FILLER_47_1167 ();
 sg13g2_decap_8 FILLER_47_1174 ();
 sg13g2_fill_2 FILLER_47_1181 ();
 sg13g2_fill_1 FILLER_47_1222 ();
 sg13g2_fill_2 FILLER_47_1230 ();
 sg13g2_fill_1 FILLER_47_1273 ();
 sg13g2_decap_4 FILLER_47_1314 ();
 sg13g2_fill_1 FILLER_47_1318 ();
 sg13g2_decap_4 FILLER_47_1345 ();
 sg13g2_decap_8 FILLER_47_1386 ();
 sg13g2_fill_1 FILLER_47_1393 ();
 sg13g2_decap_8 FILLER_47_1420 ();
 sg13g2_decap_8 FILLER_47_1427 ();
 sg13g2_fill_2 FILLER_47_1434 ();
 sg13g2_decap_4 FILLER_47_1450 ();
 sg13g2_fill_2 FILLER_47_1454 ();
 sg13g2_decap_4 FILLER_47_1460 ();
 sg13g2_fill_1 FILLER_47_1464 ();
 sg13g2_fill_2 FILLER_47_1506 ();
 sg13g2_fill_1 FILLER_47_1508 ();
 sg13g2_decap_4 FILLER_47_1535 ();
 sg13g2_fill_2 FILLER_47_1539 ();
 sg13g2_decap_4 FILLER_47_1545 ();
 sg13g2_decap_4 FILLER_47_1553 ();
 sg13g2_fill_2 FILLER_47_1557 ();
 sg13g2_fill_1 FILLER_47_1563 ();
 sg13g2_fill_1 FILLER_47_1568 ();
 sg13g2_fill_2 FILLER_47_1573 ();
 sg13g2_fill_2 FILLER_47_1619 ();
 sg13g2_fill_1 FILLER_47_1621 ();
 sg13g2_decap_4 FILLER_47_1638 ();
 sg13g2_fill_1 FILLER_47_1642 ();
 sg13g2_fill_1 FILLER_47_1651 ();
 sg13g2_fill_2 FILLER_47_1681 ();
 sg13g2_decap_8 FILLER_47_1725 ();
 sg13g2_decap_8 FILLER_47_1732 ();
 sg13g2_fill_2 FILLER_47_1739 ();
 sg13g2_fill_1 FILLER_47_1741 ();
 sg13g2_fill_2 FILLER_47_1747 ();
 sg13g2_decap_8 FILLER_47_1753 ();
 sg13g2_fill_1 FILLER_47_1760 ();
 sg13g2_decap_4 FILLER_47_1766 ();
 sg13g2_fill_2 FILLER_47_1770 ();
 sg13g2_fill_2 FILLER_47_1775 ();
 sg13g2_decap_4 FILLER_47_1786 ();
 sg13g2_fill_2 FILLER_47_1790 ();
 sg13g2_decap_8 FILLER_47_1796 ();
 sg13g2_decap_8 FILLER_47_1803 ();
 sg13g2_decap_8 FILLER_47_1810 ();
 sg13g2_fill_2 FILLER_47_1817 ();
 sg13g2_fill_1 FILLER_47_1819 ();
 sg13g2_decap_8 FILLER_47_1839 ();
 sg13g2_decap_4 FILLER_47_1846 ();
 sg13g2_fill_1 FILLER_47_1850 ();
 sg13g2_decap_8 FILLER_47_1860 ();
 sg13g2_decap_8 FILLER_47_1867 ();
 sg13g2_fill_1 FILLER_47_1874 ();
 sg13g2_fill_1 FILLER_47_1901 ();
 sg13g2_fill_1 FILLER_47_1915 ();
 sg13g2_fill_2 FILLER_47_1920 ();
 sg13g2_fill_1 FILLER_47_1922 ();
 sg13g2_fill_2 FILLER_47_1930 ();
 sg13g2_fill_1 FILLER_47_1954 ();
 sg13g2_decap_4 FILLER_47_1959 ();
 sg13g2_fill_1 FILLER_47_1963 ();
 sg13g2_fill_2 FILLER_47_1977 ();
 sg13g2_fill_1 FILLER_47_1983 ();
 sg13g2_fill_1 FILLER_47_1988 ();
 sg13g2_fill_1 FILLER_47_2011 ();
 sg13g2_decap_8 FILLER_47_2016 ();
 sg13g2_fill_2 FILLER_47_2027 ();
 sg13g2_fill_1 FILLER_47_2029 ();
 sg13g2_decap_4 FILLER_47_2049 ();
 sg13g2_fill_1 FILLER_47_2053 ();
 sg13g2_decap_8 FILLER_47_2062 ();
 sg13g2_fill_1 FILLER_47_2069 ();
 sg13g2_fill_2 FILLER_47_2099 ();
 sg13g2_fill_2 FILLER_47_2107 ();
 sg13g2_fill_2 FILLER_47_2112 ();
 sg13g2_decap_8 FILLER_47_2138 ();
 sg13g2_decap_8 FILLER_47_2145 ();
 sg13g2_fill_1 FILLER_47_2170 ();
 sg13g2_fill_2 FILLER_47_2232 ();
 sg13g2_decap_4 FILLER_47_2240 ();
 sg13g2_fill_2 FILLER_47_2252 ();
 sg13g2_decap_8 FILLER_47_2259 ();
 sg13g2_fill_2 FILLER_47_2266 ();
 sg13g2_fill_1 FILLER_47_2268 ();
 sg13g2_decap_8 FILLER_47_2295 ();
 sg13g2_fill_2 FILLER_47_2328 ();
 sg13g2_fill_1 FILLER_47_2401 ();
 sg13g2_decap_8 FILLER_47_2428 ();
 sg13g2_decap_8 FILLER_47_2439 ();
 sg13g2_decap_4 FILLER_47_2446 ();
 sg13g2_decap_8 FILLER_47_2456 ();
 sg13g2_decap_8 FILLER_47_2472 ();
 sg13g2_fill_1 FILLER_47_2479 ();
 sg13g2_decap_4 FILLER_47_2494 ();
 sg13g2_decap_8 FILLER_47_2555 ();
 sg13g2_decap_8 FILLER_47_2592 ();
 sg13g2_decap_8 FILLER_47_2599 ();
 sg13g2_decap_8 FILLER_47_2606 ();
 sg13g2_decap_8 FILLER_47_2613 ();
 sg13g2_decap_8 FILLER_47_2620 ();
 sg13g2_decap_8 FILLER_47_2631 ();
 sg13g2_decap_8 FILLER_47_2638 ();
 sg13g2_decap_8 FILLER_47_2645 ();
 sg13g2_decap_8 FILLER_47_2652 ();
 sg13g2_decap_8 FILLER_47_2659 ();
 sg13g2_decap_4 FILLER_47_2666 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_4 FILLER_48_35 ();
 sg13g2_fill_2 FILLER_48_39 ();
 sg13g2_fill_2 FILLER_48_62 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_fill_2 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_125 ();
 sg13g2_decap_8 FILLER_48_132 ();
 sg13g2_decap_8 FILLER_48_139 ();
 sg13g2_decap_8 FILLER_48_146 ();
 sg13g2_decap_8 FILLER_48_153 ();
 sg13g2_decap_4 FILLER_48_160 ();
 sg13g2_fill_2 FILLER_48_164 ();
 sg13g2_decap_8 FILLER_48_214 ();
 sg13g2_decap_8 FILLER_48_271 ();
 sg13g2_decap_4 FILLER_48_278 ();
 sg13g2_fill_2 FILLER_48_282 ();
 sg13g2_fill_1 FILLER_48_289 ();
 sg13g2_decap_4 FILLER_48_297 ();
 sg13g2_fill_1 FILLER_48_342 ();
 sg13g2_decap_8 FILLER_48_347 ();
 sg13g2_decap_8 FILLER_48_354 ();
 sg13g2_decap_8 FILLER_48_361 ();
 sg13g2_decap_8 FILLER_48_383 ();
 sg13g2_decap_4 FILLER_48_390 ();
 sg13g2_fill_2 FILLER_48_394 ();
 sg13g2_fill_2 FILLER_48_439 ();
 sg13g2_fill_2 FILLER_48_446 ();
 sg13g2_fill_1 FILLER_48_448 ();
 sg13g2_fill_2 FILLER_48_454 ();
 sg13g2_fill_1 FILLER_48_456 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_fill_1 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_520 ();
 sg13g2_fill_1 FILLER_48_536 ();
 sg13g2_fill_1 FILLER_48_542 ();
 sg13g2_fill_1 FILLER_48_548 ();
 sg13g2_fill_2 FILLER_48_566 ();
 sg13g2_fill_1 FILLER_48_568 ();
 sg13g2_fill_1 FILLER_48_573 ();
 sg13g2_decap_4 FILLER_48_587 ();
 sg13g2_fill_1 FILLER_48_591 ();
 sg13g2_fill_1 FILLER_48_619 ();
 sg13g2_fill_1 FILLER_48_633 ();
 sg13g2_decap_8 FILLER_48_661 ();
 sg13g2_decap_8 FILLER_48_668 ();
 sg13g2_decap_8 FILLER_48_680 ();
 sg13g2_decap_8 FILLER_48_687 ();
 sg13g2_fill_1 FILLER_48_694 ();
 sg13g2_decap_8 FILLER_48_702 ();
 sg13g2_decap_4 FILLER_48_709 ();
 sg13g2_fill_1 FILLER_48_713 ();
 sg13g2_decap_8 FILLER_48_731 ();
 sg13g2_decap_8 FILLER_48_738 ();
 sg13g2_decap_4 FILLER_48_770 ();
 sg13g2_decap_8 FILLER_48_779 ();
 sg13g2_decap_8 FILLER_48_786 ();
 sg13g2_decap_8 FILLER_48_793 ();
 sg13g2_decap_8 FILLER_48_800 ();
 sg13g2_decap_8 FILLER_48_807 ();
 sg13g2_decap_4 FILLER_48_814 ();
 sg13g2_fill_2 FILLER_48_818 ();
 sg13g2_fill_1 FILLER_48_824 ();
 sg13g2_fill_2 FILLER_48_830 ();
 sg13g2_decap_8 FILLER_48_850 ();
 sg13g2_decap_8 FILLER_48_857 ();
 sg13g2_fill_2 FILLER_48_864 ();
 sg13g2_fill_1 FILLER_48_893 ();
 sg13g2_decap_4 FILLER_48_920 ();
 sg13g2_fill_1 FILLER_48_924 ();
 sg13g2_decap_4 FILLER_48_940 ();
 sg13g2_fill_2 FILLER_48_944 ();
 sg13g2_decap_8 FILLER_48_951 ();
 sg13g2_decap_8 FILLER_48_958 ();
 sg13g2_fill_2 FILLER_48_965 ();
 sg13g2_decap_8 FILLER_48_973 ();
 sg13g2_fill_1 FILLER_48_980 ();
 sg13g2_decap_8 FILLER_48_985 ();
 sg13g2_decap_4 FILLER_48_992 ();
 sg13g2_fill_1 FILLER_48_996 ();
 sg13g2_decap_4 FILLER_48_1001 ();
 sg13g2_fill_1 FILLER_48_1053 ();
 sg13g2_fill_1 FILLER_48_1080 ();
 sg13g2_fill_1 FILLER_48_1140 ();
 sg13g2_fill_1 FILLER_48_1147 ();
 sg13g2_fill_1 FILLER_48_1159 ();
 sg13g2_decap_8 FILLER_48_1174 ();
 sg13g2_decap_8 FILLER_48_1181 ();
 sg13g2_decap_4 FILLER_48_1188 ();
 sg13g2_fill_1 FILLER_48_1235 ();
 sg13g2_fill_1 FILLER_48_1270 ();
 sg13g2_decap_8 FILLER_48_1312 ();
 sg13g2_decap_8 FILLER_48_1319 ();
 sg13g2_fill_1 FILLER_48_1326 ();
 sg13g2_decap_8 FILLER_48_1335 ();
 sg13g2_decap_8 FILLER_48_1342 ();
 sg13g2_fill_2 FILLER_48_1349 ();
 sg13g2_decap_8 FILLER_48_1386 ();
 sg13g2_decap_8 FILLER_48_1393 ();
 sg13g2_fill_1 FILLER_48_1400 ();
 sg13g2_decap_8 FILLER_48_1407 ();
 sg13g2_decap_8 FILLER_48_1414 ();
 sg13g2_decap_8 FILLER_48_1421 ();
 sg13g2_fill_2 FILLER_48_1467 ();
 sg13g2_fill_1 FILLER_48_1469 ();
 sg13g2_decap_8 FILLER_48_1474 ();
 sg13g2_decap_4 FILLER_48_1485 ();
 sg13g2_fill_2 FILLER_48_1489 ();
 sg13g2_fill_2 FILLER_48_1497 ();
 sg13g2_fill_1 FILLER_48_1503 ();
 sg13g2_fill_2 FILLER_48_1511 ();
 sg13g2_fill_2 FILLER_48_1539 ();
 sg13g2_fill_1 FILLER_48_1541 ();
 sg13g2_decap_8 FILLER_48_1568 ();
 sg13g2_fill_1 FILLER_48_1665 ();
 sg13g2_fill_1 FILLER_48_1674 ();
 sg13g2_fill_1 FILLER_48_1685 ();
 sg13g2_decap_8 FILLER_48_1717 ();
 sg13g2_decap_8 FILLER_48_1724 ();
 sg13g2_decap_8 FILLER_48_1731 ();
 sg13g2_decap_8 FILLER_48_1738 ();
 sg13g2_fill_2 FILLER_48_1745 ();
 sg13g2_fill_1 FILLER_48_1747 ();
 sg13g2_decap_8 FILLER_48_1816 ();
 sg13g2_decap_4 FILLER_48_1823 ();
 sg13g2_fill_2 FILLER_48_1827 ();
 sg13g2_decap_4 FILLER_48_1834 ();
 sg13g2_fill_2 FILLER_48_1838 ();
 sg13g2_fill_2 FILLER_48_1845 ();
 sg13g2_fill_1 FILLER_48_1847 ();
 sg13g2_decap_8 FILLER_48_1857 ();
 sg13g2_fill_1 FILLER_48_1864 ();
 sg13g2_decap_8 FILLER_48_1870 ();
 sg13g2_fill_2 FILLER_48_1877 ();
 sg13g2_fill_1 FILLER_48_1879 ();
 sg13g2_decap_8 FILLER_48_1890 ();
 sg13g2_fill_2 FILLER_48_1902 ();
 sg13g2_fill_1 FILLER_48_1904 ();
 sg13g2_decap_4 FILLER_48_1911 ();
 sg13g2_decap_4 FILLER_48_1919 ();
 sg13g2_decap_4 FILLER_48_1929 ();
 sg13g2_fill_1 FILLER_48_1937 ();
 sg13g2_decap_4 FILLER_48_1958 ();
 sg13g2_decap_4 FILLER_48_1966 ();
 sg13g2_decap_4 FILLER_48_1975 ();
 sg13g2_fill_1 FILLER_48_1979 ();
 sg13g2_fill_2 FILLER_48_1984 ();
 sg13g2_decap_8 FILLER_48_1990 ();
 sg13g2_decap_8 FILLER_48_1997 ();
 sg13g2_fill_1 FILLER_48_2004 ();
 sg13g2_fill_2 FILLER_48_2008 ();
 sg13g2_decap_8 FILLER_48_2014 ();
 sg13g2_decap_4 FILLER_48_2021 ();
 sg13g2_fill_2 FILLER_48_2034 ();
 sg13g2_decap_4 FILLER_48_2080 ();
 sg13g2_fill_1 FILLER_48_2084 ();
 sg13g2_fill_1 FILLER_48_2102 ();
 sg13g2_fill_2 FILLER_48_2123 ();
 sg13g2_decap_4 FILLER_48_2151 ();
 sg13g2_decap_8 FILLER_48_2194 ();
 sg13g2_fill_1 FILLER_48_2201 ();
 sg13g2_fill_1 FILLER_48_2279 ();
 sg13g2_decap_8 FILLER_48_2284 ();
 sg13g2_decap_8 FILLER_48_2291 ();
 sg13g2_fill_2 FILLER_48_2298 ();
 sg13g2_fill_1 FILLER_48_2300 ();
 sg13g2_decap_8 FILLER_48_2335 ();
 sg13g2_decap_8 FILLER_48_2342 ();
 sg13g2_decap_8 FILLER_48_2349 ();
 sg13g2_fill_2 FILLER_48_2356 ();
 sg13g2_fill_1 FILLER_48_2358 ();
 sg13g2_decap_8 FILLER_48_2365 ();
 sg13g2_fill_2 FILLER_48_2372 ();
 sg13g2_fill_1 FILLER_48_2374 ();
 sg13g2_decap_4 FILLER_48_2383 ();
 sg13g2_decap_8 FILLER_48_2406 ();
 sg13g2_fill_1 FILLER_48_2413 ();
 sg13g2_fill_1 FILLER_48_2420 ();
 sg13g2_decap_8 FILLER_48_2425 ();
 sg13g2_fill_2 FILLER_48_2432 ();
 sg13g2_fill_2 FILLER_48_2465 ();
 sg13g2_fill_2 FILLER_48_2493 ();
 sg13g2_fill_2 FILLER_48_2562 ();
 sg13g2_fill_1 FILLER_48_2577 ();
 sg13g2_decap_8 FILLER_48_2587 ();
 sg13g2_fill_1 FILLER_48_2594 ();
 sg13g2_decap_8 FILLER_48_2608 ();
 sg13g2_fill_1 FILLER_48_2619 ();
 sg13g2_decap_8 FILLER_48_2646 ();
 sg13g2_decap_8 FILLER_48_2653 ();
 sg13g2_decap_8 FILLER_48_2660 ();
 sg13g2_fill_2 FILLER_48_2667 ();
 sg13g2_fill_1 FILLER_48_2669 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_fill_1 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_23 ();
 sg13g2_decap_4 FILLER_49_30 ();
 sg13g2_fill_1 FILLER_49_34 ();
 sg13g2_fill_2 FILLER_49_39 ();
 sg13g2_fill_1 FILLER_49_58 ();
 sg13g2_decap_4 FILLER_49_68 ();
 sg13g2_fill_2 FILLER_49_72 ();
 sg13g2_decap_4 FILLER_49_99 ();
 sg13g2_decap_8 FILLER_49_117 ();
 sg13g2_decap_8 FILLER_49_124 ();
 sg13g2_decap_8 FILLER_49_131 ();
 sg13g2_decap_8 FILLER_49_138 ();
 sg13g2_decap_8 FILLER_49_145 ();
 sg13g2_decap_8 FILLER_49_152 ();
 sg13g2_decap_8 FILLER_49_159 ();
 sg13g2_decap_8 FILLER_49_166 ();
 sg13g2_decap_8 FILLER_49_173 ();
 sg13g2_decap_8 FILLER_49_180 ();
 sg13g2_decap_8 FILLER_49_187 ();
 sg13g2_decap_8 FILLER_49_194 ();
 sg13g2_decap_8 FILLER_49_201 ();
 sg13g2_decap_8 FILLER_49_208 ();
 sg13g2_decap_8 FILLER_49_215 ();
 sg13g2_fill_1 FILLER_49_266 ();
 sg13g2_fill_2 FILLER_49_272 ();
 sg13g2_decap_8 FILLER_49_303 ();
 sg13g2_decap_8 FILLER_49_310 ();
 sg13g2_decap_8 FILLER_49_317 ();
 sg13g2_fill_2 FILLER_49_324 ();
 sg13g2_decap_8 FILLER_49_330 ();
 sg13g2_decap_4 FILLER_49_337 ();
 sg13g2_fill_2 FILLER_49_341 ();
 sg13g2_decap_8 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_decap_4 FILLER_49_440 ();
 sg13g2_fill_2 FILLER_49_444 ();
 sg13g2_fill_1 FILLER_49_450 ();
 sg13g2_decap_4 FILLER_49_481 ();
 sg13g2_decap_8 FILLER_49_489 ();
 sg13g2_decap_4 FILLER_49_496 ();
 sg13g2_fill_2 FILLER_49_500 ();
 sg13g2_fill_1 FILLER_49_506 ();
 sg13g2_fill_1 FILLER_49_512 ();
 sg13g2_fill_1 FILLER_49_524 ();
 sg13g2_fill_1 FILLER_49_531 ();
 sg13g2_decap_8 FILLER_49_536 ();
 sg13g2_decap_8 FILLER_49_543 ();
 sg13g2_fill_2 FILLER_49_550 ();
 sg13g2_decap_4 FILLER_49_562 ();
 sg13g2_fill_1 FILLER_49_566 ();
 sg13g2_fill_2 FILLER_49_619 ();
 sg13g2_fill_1 FILLER_49_648 ();
 sg13g2_decap_8 FILLER_49_663 ();
 sg13g2_fill_1 FILLER_49_670 ();
 sg13g2_fill_2 FILLER_49_675 ();
 sg13g2_fill_2 FILLER_49_698 ();
 sg13g2_decap_4 FILLER_49_705 ();
 sg13g2_decap_4 FILLER_49_717 ();
 sg13g2_decap_8 FILLER_49_730 ();
 sg13g2_decap_4 FILLER_49_737 ();
 sg13g2_fill_1 FILLER_49_746 ();
 sg13g2_fill_2 FILLER_49_752 ();
 sg13g2_fill_1 FILLER_49_767 ();
 sg13g2_decap_4 FILLER_49_780 ();
 sg13g2_decap_8 FILLER_49_787 ();
 sg13g2_decap_8 FILLER_49_794 ();
 sg13g2_fill_1 FILLER_49_801 ();
 sg13g2_fill_1 FILLER_49_828 ();
 sg13g2_fill_1 FILLER_49_844 ();
 sg13g2_fill_2 FILLER_49_854 ();
 sg13g2_fill_1 FILLER_49_856 ();
 sg13g2_fill_2 FILLER_49_867 ();
 sg13g2_fill_1 FILLER_49_873 ();
 sg13g2_fill_1 FILLER_49_879 ();
 sg13g2_fill_2 FILLER_49_893 ();
 sg13g2_fill_2 FILLER_49_900 ();
 sg13g2_fill_2 FILLER_49_906 ();
 sg13g2_fill_1 FILLER_49_912 ();
 sg13g2_decap_4 FILLER_49_950 ();
 sg13g2_fill_1 FILLER_49_954 ();
 sg13g2_decap_4 FILLER_49_960 ();
 sg13g2_fill_1 FILLER_49_972 ();
 sg13g2_decap_4 FILLER_49_986 ();
 sg13g2_decap_8 FILLER_49_1020 ();
 sg13g2_decap_8 FILLER_49_1027 ();
 sg13g2_fill_2 FILLER_49_1034 ();
 sg13g2_decap_4 FILLER_49_1076 ();
 sg13g2_fill_1 FILLER_49_1080 ();
 sg13g2_fill_2 FILLER_49_1091 ();
 sg13g2_fill_1 FILLER_49_1093 ();
 sg13g2_fill_2 FILLER_49_1112 ();
 sg13g2_fill_1 FILLER_49_1157 ();
 sg13g2_fill_1 FILLER_49_1184 ();
 sg13g2_decap_8 FILLER_49_1188 ();
 sg13g2_fill_2 FILLER_49_1195 ();
 sg13g2_fill_1 FILLER_49_1212 ();
 sg13g2_fill_1 FILLER_49_1223 ();
 sg13g2_fill_1 FILLER_49_1300 ();
 sg13g2_fill_1 FILLER_49_1307 ();
 sg13g2_fill_1 FILLER_49_1321 ();
 sg13g2_decap_8 FILLER_49_1328 ();
 sg13g2_decap_8 FILLER_49_1335 ();
 sg13g2_decap_8 FILLER_49_1342 ();
 sg13g2_decap_8 FILLER_49_1349 ();
 sg13g2_decap_8 FILLER_49_1356 ();
 sg13g2_decap_8 FILLER_49_1363 ();
 sg13g2_decap_8 FILLER_49_1370 ();
 sg13g2_decap_8 FILLER_49_1377 ();
 sg13g2_decap_8 FILLER_49_1384 ();
 sg13g2_fill_2 FILLER_49_1391 ();
 sg13g2_fill_1 FILLER_49_1393 ();
 sg13g2_decap_4 FILLER_49_1433 ();
 sg13g2_fill_2 FILLER_49_1437 ();
 sg13g2_decap_4 FILLER_49_1454 ();
 sg13g2_decap_8 FILLER_49_1464 ();
 sg13g2_decap_4 FILLER_49_1471 ();
 sg13g2_fill_1 FILLER_49_1475 ();
 sg13g2_decap_8 FILLER_49_1480 ();
 sg13g2_decap_4 FILLER_49_1487 ();
 sg13g2_decap_8 FILLER_49_1494 ();
 sg13g2_fill_2 FILLER_49_1528 ();
 sg13g2_decap_8 FILLER_49_1564 ();
 sg13g2_decap_8 FILLER_49_1571 ();
 sg13g2_decap_8 FILLER_49_1578 ();
 sg13g2_fill_2 FILLER_49_1585 ();
 sg13g2_fill_2 FILLER_49_1591 ();
 sg13g2_fill_1 FILLER_49_1596 ();
 sg13g2_decap_8 FILLER_49_1607 ();
 sg13g2_fill_1 FILLER_49_1614 ();
 sg13g2_fill_2 FILLER_49_1619 ();
 sg13g2_fill_1 FILLER_49_1641 ();
 sg13g2_fill_2 FILLER_49_1646 ();
 sg13g2_fill_1 FILLER_49_1652 ();
 sg13g2_fill_2 FILLER_49_1661 ();
 sg13g2_fill_2 FILLER_49_1672 ();
 sg13g2_fill_1 FILLER_49_1681 ();
 sg13g2_decap_8 FILLER_49_1696 ();
 sg13g2_decap_4 FILLER_49_1703 ();
 sg13g2_fill_2 FILLER_49_1714 ();
 sg13g2_fill_1 FILLER_49_1759 ();
 sg13g2_fill_1 FILLER_49_1772 ();
 sg13g2_fill_2 FILLER_49_1842 ();
 sg13g2_fill_1 FILLER_49_1844 ();
 sg13g2_decap_8 FILLER_49_1850 ();
 sg13g2_decap_8 FILLER_49_1862 ();
 sg13g2_decap_8 FILLER_49_1869 ();
 sg13g2_decap_8 FILLER_49_1876 ();
 sg13g2_decap_8 FILLER_49_1883 ();
 sg13g2_decap_8 FILLER_49_1890 ();
 sg13g2_decap_8 FILLER_49_1897 ();
 sg13g2_decap_4 FILLER_49_1904 ();
 sg13g2_decap_8 FILLER_49_1914 ();
 sg13g2_decap_8 FILLER_49_1921 ();
 sg13g2_decap_8 FILLER_49_1928 ();
 sg13g2_fill_2 FILLER_49_1935 ();
 sg13g2_fill_1 FILLER_49_1937 ();
 sg13g2_fill_2 FILLER_49_1950 ();
 sg13g2_fill_1 FILLER_49_1952 ();
 sg13g2_fill_2 FILLER_49_1970 ();
 sg13g2_decap_8 FILLER_49_2023 ();
 sg13g2_decap_8 FILLER_49_2030 ();
 sg13g2_fill_2 FILLER_49_2037 ();
 sg13g2_fill_2 FILLER_49_2049 ();
 sg13g2_decap_4 FILLER_49_2063 ();
 sg13g2_fill_1 FILLER_49_2067 ();
 sg13g2_decap_4 FILLER_49_2072 ();
 sg13g2_fill_1 FILLER_49_2081 ();
 sg13g2_fill_1 FILLER_49_2111 ();
 sg13g2_fill_1 FILLER_49_2138 ();
 sg13g2_fill_1 FILLER_49_2169 ();
 sg13g2_fill_1 FILLER_49_2178 ();
 sg13g2_decap_8 FILLER_49_2183 ();
 sg13g2_decap_8 FILLER_49_2190 ();
 sg13g2_decap_8 FILLER_49_2197 ();
 sg13g2_fill_1 FILLER_49_2204 ();
 sg13g2_decap_8 FILLER_49_2210 ();
 sg13g2_decap_8 FILLER_49_2217 ();
 sg13g2_decap_8 FILLER_49_2263 ();
 sg13g2_decap_8 FILLER_49_2270 ();
 sg13g2_decap_8 FILLER_49_2281 ();
 sg13g2_decap_8 FILLER_49_2288 ();
 sg13g2_decap_8 FILLER_49_2295 ();
 sg13g2_decap_8 FILLER_49_2302 ();
 sg13g2_fill_2 FILLER_49_2309 ();
 sg13g2_decap_8 FILLER_49_2326 ();
 sg13g2_decap_8 FILLER_49_2333 ();
 sg13g2_decap_4 FILLER_49_2340 ();
 sg13g2_fill_1 FILLER_49_2344 ();
 sg13g2_fill_2 FILLER_49_2350 ();
 sg13g2_fill_1 FILLER_49_2352 ();
 sg13g2_decap_8 FILLER_49_2362 ();
 sg13g2_decap_8 FILLER_49_2369 ();
 sg13g2_decap_8 FILLER_49_2376 ();
 sg13g2_decap_8 FILLER_49_2383 ();
 sg13g2_decap_4 FILLER_49_2390 ();
 sg13g2_decap_8 FILLER_49_2402 ();
 sg13g2_decap_8 FILLER_49_2409 ();
 sg13g2_decap_8 FILLER_49_2416 ();
 sg13g2_fill_2 FILLER_49_2423 ();
 sg13g2_fill_2 FILLER_49_2451 ();
 sg13g2_fill_1 FILLER_49_2453 ();
 sg13g2_decap_8 FILLER_49_2463 ();
 sg13g2_decap_8 FILLER_49_2470 ();
 sg13g2_decap_8 FILLER_49_2477 ();
 sg13g2_fill_2 FILLER_49_2484 ();
 sg13g2_fill_1 FILLER_49_2486 ();
 sg13g2_decap_8 FILLER_49_2545 ();
 sg13g2_decap_8 FILLER_49_2552 ();
 sg13g2_decap_8 FILLER_49_2559 ();
 sg13g2_decap_8 FILLER_49_2566 ();
 sg13g2_decap_8 FILLER_49_2573 ();
 sg13g2_decap_8 FILLER_49_2580 ();
 sg13g2_decap_4 FILLER_49_2587 ();
 sg13g2_fill_1 FILLER_49_2598 ();
 sg13g2_decap_8 FILLER_49_2625 ();
 sg13g2_decap_8 FILLER_49_2632 ();
 sg13g2_decap_8 FILLER_49_2639 ();
 sg13g2_decap_8 FILLER_49_2646 ();
 sg13g2_decap_8 FILLER_49_2653 ();
 sg13g2_decap_8 FILLER_49_2660 ();
 sg13g2_fill_2 FILLER_49_2667 ();
 sg13g2_fill_1 FILLER_49_2669 ();
 sg13g2_decap_4 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_4 ();
 sg13g2_fill_1 FILLER_50_32 ();
 sg13g2_fill_1 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_62 ();
 sg13g2_decap_8 FILLER_50_69 ();
 sg13g2_decap_8 FILLER_50_76 ();
 sg13g2_decap_4 FILLER_50_83 ();
 sg13g2_decap_8 FILLER_50_117 ();
 sg13g2_fill_2 FILLER_50_124 ();
 sg13g2_decap_8 FILLER_50_181 ();
 sg13g2_decap_8 FILLER_50_188 ();
 sg13g2_decap_8 FILLER_50_195 ();
 sg13g2_decap_8 FILLER_50_202 ();
 sg13g2_decap_8 FILLER_50_209 ();
 sg13g2_decap_8 FILLER_50_216 ();
 sg13g2_fill_2 FILLER_50_223 ();
 sg13g2_fill_1 FILLER_50_241 ();
 sg13g2_fill_2 FILLER_50_245 ();
 sg13g2_fill_2 FILLER_50_256 ();
 sg13g2_fill_2 FILLER_50_277 ();
 sg13g2_decap_4 FILLER_50_282 ();
 sg13g2_fill_1 FILLER_50_286 ();
 sg13g2_decap_8 FILLER_50_306 ();
 sg13g2_decap_8 FILLER_50_313 ();
 sg13g2_fill_1 FILLER_50_320 ();
 sg13g2_fill_2 FILLER_50_327 ();
 sg13g2_decap_8 FILLER_50_342 ();
 sg13g2_decap_8 FILLER_50_349 ();
 sg13g2_decap_4 FILLER_50_359 ();
 sg13g2_fill_1 FILLER_50_363 ();
 sg13g2_decap_8 FILLER_50_388 ();
 sg13g2_decap_8 FILLER_50_395 ();
 sg13g2_fill_2 FILLER_50_402 ();
 sg13g2_fill_1 FILLER_50_404 ();
 sg13g2_fill_1 FILLER_50_418 ();
 sg13g2_fill_1 FILLER_50_423 ();
 sg13g2_decap_4 FILLER_50_439 ();
 sg13g2_fill_2 FILLER_50_466 ();
 sg13g2_fill_1 FILLER_50_468 ();
 sg13g2_decap_4 FILLER_50_473 ();
 sg13g2_decap_8 FILLER_50_482 ();
 sg13g2_fill_2 FILLER_50_489 ();
 sg13g2_decap_4 FILLER_50_496 ();
 sg13g2_fill_1 FILLER_50_500 ();
 sg13g2_decap_4 FILLER_50_508 ();
 sg13g2_fill_1 FILLER_50_518 ();
 sg13g2_fill_2 FILLER_50_528 ();
 sg13g2_fill_1 FILLER_50_530 ();
 sg13g2_decap_8 FILLER_50_558 ();
 sg13g2_decap_4 FILLER_50_565 ();
 sg13g2_fill_1 FILLER_50_569 ();
 sg13g2_fill_2 FILLER_50_574 ();
 sg13g2_fill_1 FILLER_50_576 ();
 sg13g2_decap_8 FILLER_50_582 ();
 sg13g2_decap_8 FILLER_50_589 ();
 sg13g2_decap_8 FILLER_50_596 ();
 sg13g2_fill_2 FILLER_50_623 ();
 sg13g2_fill_1 FILLER_50_639 ();
 sg13g2_fill_1 FILLER_50_645 ();
 sg13g2_decap_4 FILLER_50_655 ();
 sg13g2_decap_4 FILLER_50_663 ();
 sg13g2_decap_4 FILLER_50_671 ();
 sg13g2_decap_8 FILLER_50_700 ();
 sg13g2_fill_1 FILLER_50_707 ();
 sg13g2_fill_1 FILLER_50_727 ();
 sg13g2_decap_8 FILLER_50_732 ();
 sg13g2_decap_8 FILLER_50_739 ();
 sg13g2_fill_2 FILLER_50_746 ();
 sg13g2_fill_1 FILLER_50_782 ();
 sg13g2_fill_1 FILLER_50_787 ();
 sg13g2_fill_1 FILLER_50_820 ();
 sg13g2_fill_1 FILLER_50_848 ();
 sg13g2_decap_8 FILLER_50_854 ();
 sg13g2_decap_8 FILLER_50_861 ();
 sg13g2_fill_1 FILLER_50_868 ();
 sg13g2_fill_2 FILLER_50_908 ();
 sg13g2_fill_1 FILLER_50_919 ();
 sg13g2_fill_1 FILLER_50_925 ();
 sg13g2_decap_8 FILLER_50_938 ();
 sg13g2_decap_8 FILLER_50_945 ();
 sg13g2_fill_2 FILLER_50_952 ();
 sg13g2_fill_1 FILLER_50_954 ();
 sg13g2_fill_1 FILLER_50_961 ();
 sg13g2_fill_2 FILLER_50_970 ();
 sg13g2_fill_1 FILLER_50_998 ();
 sg13g2_decap_8 FILLER_50_1035 ();
 sg13g2_fill_1 FILLER_50_1042 ();
 sg13g2_decap_4 FILLER_50_1047 ();
 sg13g2_decap_8 FILLER_50_1056 ();
 sg13g2_decap_8 FILLER_50_1063 ();
 sg13g2_decap_8 FILLER_50_1070 ();
 sg13g2_decap_8 FILLER_50_1077 ();
 sg13g2_fill_2 FILLER_50_1104 ();
 sg13g2_fill_1 FILLER_50_1110 ();
 sg13g2_fill_1 FILLER_50_1152 ();
 sg13g2_fill_2 FILLER_50_1165 ();
 sg13g2_fill_2 FILLER_50_1180 ();
 sg13g2_fill_2 FILLER_50_1312 ();
 sg13g2_fill_1 FILLER_50_1318 ();
 sg13g2_fill_1 FILLER_50_1328 ();
 sg13g2_decap_4 FILLER_50_1363 ();
 sg13g2_fill_1 FILLER_50_1367 ();
 sg13g2_decap_8 FILLER_50_1372 ();
 sg13g2_decap_8 FILLER_50_1379 ();
 sg13g2_decap_8 FILLER_50_1386 ();
 sg13g2_decap_4 FILLER_50_1393 ();
 sg13g2_fill_1 FILLER_50_1397 ();
 sg13g2_fill_2 FILLER_50_1403 ();
 sg13g2_decap_4 FILLER_50_1410 ();
 sg13g2_decap_4 FILLER_50_1426 ();
 sg13g2_decap_4 FILLER_50_1442 ();
 sg13g2_fill_1 FILLER_50_1472 ();
 sg13g2_decap_8 FILLER_50_1486 ();
 sg13g2_decap_8 FILLER_50_1493 ();
 sg13g2_fill_2 FILLER_50_1500 ();
 sg13g2_fill_1 FILLER_50_1502 ();
 sg13g2_fill_2 FILLER_50_1508 ();
 sg13g2_fill_1 FILLER_50_1510 ();
 sg13g2_decap_4 FILLER_50_1515 ();
 sg13g2_fill_2 FILLER_50_1519 ();
 sg13g2_fill_1 FILLER_50_1526 ();
 sg13g2_decap_4 FILLER_50_1531 ();
 sg13g2_decap_8 FILLER_50_1538 ();
 sg13g2_decap_8 FILLER_50_1545 ();
 sg13g2_decap_4 FILLER_50_1552 ();
 sg13g2_fill_2 FILLER_50_1556 ();
 sg13g2_decap_8 FILLER_50_1580 ();
 sg13g2_fill_2 FILLER_50_1587 ();
 sg13g2_fill_1 FILLER_50_1589 ();
 sg13g2_fill_2 FILLER_50_1599 ();
 sg13g2_decap_4 FILLER_50_1605 ();
 sg13g2_fill_2 FILLER_50_1636 ();
 sg13g2_fill_1 FILLER_50_1684 ();
 sg13g2_decap_8 FILLER_50_1690 ();
 sg13g2_decap_8 FILLER_50_1697 ();
 sg13g2_fill_2 FILLER_50_1704 ();
 sg13g2_fill_1 FILLER_50_1706 ();
 sg13g2_decap_8 FILLER_50_1721 ();
 sg13g2_fill_2 FILLER_50_1728 ();
 sg13g2_decap_8 FILLER_50_1738 ();
 sg13g2_decap_4 FILLER_50_1745 ();
 sg13g2_fill_2 FILLER_50_1749 ();
 sg13g2_fill_2 FILLER_50_1761 ();
 sg13g2_fill_1 FILLER_50_1763 ();
 sg13g2_fill_1 FILLER_50_1777 ();
 sg13g2_fill_1 FILLER_50_1782 ();
 sg13g2_fill_1 FILLER_50_1789 ();
 sg13g2_fill_2 FILLER_50_1821 ();
 sg13g2_fill_1 FILLER_50_1823 ();
 sg13g2_fill_2 FILLER_50_1828 ();
 sg13g2_fill_1 FILLER_50_1830 ();
 sg13g2_decap_8 FILLER_50_1845 ();
 sg13g2_decap_4 FILLER_50_1852 ();
 sg13g2_decap_4 FILLER_50_1863 ();
 sg13g2_fill_2 FILLER_50_1881 ();
 sg13g2_decap_4 FILLER_50_1897 ();
 sg13g2_fill_1 FILLER_50_1901 ();
 sg13g2_fill_2 FILLER_50_1911 ();
 sg13g2_decap_8 FILLER_50_1928 ();
 sg13g2_decap_8 FILLER_50_1935 ();
 sg13g2_fill_2 FILLER_50_1946 ();
 sg13g2_fill_1 FILLER_50_1948 ();
 sg13g2_decap_8 FILLER_50_1954 ();
 sg13g2_decap_8 FILLER_50_1977 ();
 sg13g2_fill_1 FILLER_50_1984 ();
 sg13g2_decap_4 FILLER_50_1994 ();
 sg13g2_fill_1 FILLER_50_1998 ();
 sg13g2_decap_4 FILLER_50_2029 ();
 sg13g2_fill_1 FILLER_50_2033 ();
 sg13g2_decap_4 FILLER_50_2039 ();
 sg13g2_fill_2 FILLER_50_2101 ();
 sg13g2_fill_1 FILLER_50_2112 ();
 sg13g2_fill_1 FILLER_50_2126 ();
 sg13g2_decap_8 FILLER_50_2198 ();
 sg13g2_decap_8 FILLER_50_2205 ();
 sg13g2_fill_1 FILLER_50_2217 ();
 sg13g2_decap_8 FILLER_50_2239 ();
 sg13g2_decap_8 FILLER_50_2246 ();
 sg13g2_decap_8 FILLER_50_2253 ();
 sg13g2_fill_2 FILLER_50_2260 ();
 sg13g2_decap_4 FILLER_50_2267 ();
 sg13g2_fill_1 FILLER_50_2271 ();
 sg13g2_fill_2 FILLER_50_2276 ();
 sg13g2_decap_8 FILLER_50_2292 ();
 sg13g2_fill_2 FILLER_50_2299 ();
 sg13g2_fill_1 FILLER_50_2301 ();
 sg13g2_fill_2 FILLER_50_2316 ();
 sg13g2_decap_4 FILLER_50_2322 ();
 sg13g2_decap_4 FILLER_50_2332 ();
 sg13g2_fill_1 FILLER_50_2341 ();
 sg13g2_decap_8 FILLER_50_2372 ();
 sg13g2_decap_8 FILLER_50_2379 ();
 sg13g2_decap_8 FILLER_50_2386 ();
 sg13g2_decap_8 FILLER_50_2393 ();
 sg13g2_decap_8 FILLER_50_2400 ();
 sg13g2_decap_8 FILLER_50_2407 ();
 sg13g2_decap_8 FILLER_50_2414 ();
 sg13g2_decap_8 FILLER_50_2421 ();
 sg13g2_decap_8 FILLER_50_2428 ();
 sg13g2_decap_8 FILLER_50_2435 ();
 sg13g2_fill_1 FILLER_50_2442 ();
 sg13g2_decap_8 FILLER_50_2447 ();
 sg13g2_decap_8 FILLER_50_2454 ();
 sg13g2_decap_4 FILLER_50_2461 ();
 sg13g2_fill_2 FILLER_50_2465 ();
 sg13g2_decap_4 FILLER_50_2471 ();
 sg13g2_fill_1 FILLER_50_2475 ();
 sg13g2_decap_8 FILLER_50_2480 ();
 sg13g2_fill_2 FILLER_50_2487 ();
 sg13g2_fill_2 FILLER_50_2539 ();
 sg13g2_fill_2 FILLER_50_2567 ();
 sg13g2_decap_8 FILLER_50_2604 ();
 sg13g2_decap_8 FILLER_50_2611 ();
 sg13g2_decap_8 FILLER_50_2618 ();
 sg13g2_decap_8 FILLER_50_2625 ();
 sg13g2_decap_8 FILLER_50_2632 ();
 sg13g2_decap_8 FILLER_50_2639 ();
 sg13g2_decap_8 FILLER_50_2646 ();
 sg13g2_decap_8 FILLER_50_2653 ();
 sg13g2_decap_8 FILLER_50_2660 ();
 sg13g2_fill_2 FILLER_50_2667 ();
 sg13g2_fill_1 FILLER_50_2669 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_fill_1 FILLER_51_14 ();
 sg13g2_fill_2 FILLER_51_41 ();
 sg13g2_decap_8 FILLER_51_72 ();
 sg13g2_decap_8 FILLER_51_79 ();
 sg13g2_decap_4 FILLER_51_86 ();
 sg13g2_fill_1 FILLER_51_90 ();
 sg13g2_fill_1 FILLER_51_114 ();
 sg13g2_fill_1 FILLER_51_119 ();
 sg13g2_fill_2 FILLER_51_125 ();
 sg13g2_fill_2 FILLER_51_131 ();
 sg13g2_fill_2 FILLER_51_137 ();
 sg13g2_fill_1 FILLER_51_139 ();
 sg13g2_decap_8 FILLER_51_186 ();
 sg13g2_decap_8 FILLER_51_193 ();
 sg13g2_decap_8 FILLER_51_200 ();
 sg13g2_decap_8 FILLER_51_207 ();
 sg13g2_fill_2 FILLER_51_217 ();
 sg13g2_fill_1 FILLER_51_219 ();
 sg13g2_decap_8 FILLER_51_272 ();
 sg13g2_fill_1 FILLER_51_309 ();
 sg13g2_decap_4 FILLER_51_313 ();
 sg13g2_fill_2 FILLER_51_317 ();
 sg13g2_decap_4 FILLER_51_353 ();
 sg13g2_fill_1 FILLER_51_357 ();
 sg13g2_decap_4 FILLER_51_384 ();
 sg13g2_fill_2 FILLER_51_397 ();
 sg13g2_decap_8 FILLER_51_435 ();
 sg13g2_fill_2 FILLER_51_442 ();
 sg13g2_fill_1 FILLER_51_444 ();
 sg13g2_decap_8 FILLER_51_480 ();
 sg13g2_decap_4 FILLER_51_487 ();
 sg13g2_decap_4 FILLER_51_495 ();
 sg13g2_fill_1 FILLER_51_499 ();
 sg13g2_decap_4 FILLER_51_519 ();
 sg13g2_fill_2 FILLER_51_533 ();
 sg13g2_fill_1 FILLER_51_539 ();
 sg13g2_decap_8 FILLER_51_545 ();
 sg13g2_fill_2 FILLER_51_552 ();
 sg13g2_fill_1 FILLER_51_554 ();
 sg13g2_fill_2 FILLER_51_564 ();
 sg13g2_fill_1 FILLER_51_566 ();
 sg13g2_decap_8 FILLER_51_580 ();
 sg13g2_decap_8 FILLER_51_587 ();
 sg13g2_decap_4 FILLER_51_594 ();
 sg13g2_fill_2 FILLER_51_598 ();
 sg13g2_decap_8 FILLER_51_608 ();
 sg13g2_decap_4 FILLER_51_615 ();
 sg13g2_fill_2 FILLER_51_619 ();
 sg13g2_decap_4 FILLER_51_626 ();
 sg13g2_fill_2 FILLER_51_630 ();
 sg13g2_fill_1 FILLER_51_636 ();
 sg13g2_fill_1 FILLER_51_651 ();
 sg13g2_decap_8 FILLER_51_666 ();
 sg13g2_decap_8 FILLER_51_673 ();
 sg13g2_decap_4 FILLER_51_680 ();
 sg13g2_fill_2 FILLER_51_684 ();
 sg13g2_decap_8 FILLER_51_691 ();
 sg13g2_decap_4 FILLER_51_714 ();
 sg13g2_fill_1 FILLER_51_723 ();
 sg13g2_fill_1 FILLER_51_735 ();
 sg13g2_decap_8 FILLER_51_772 ();
 sg13g2_decap_8 FILLER_51_779 ();
 sg13g2_fill_2 FILLER_51_786 ();
 sg13g2_fill_1 FILLER_51_788 ();
 sg13g2_decap_8 FILLER_51_798 ();
 sg13g2_fill_1 FILLER_51_805 ();
 sg13g2_decap_4 FILLER_51_854 ();
 sg13g2_fill_2 FILLER_51_858 ();
 sg13g2_fill_2 FILLER_51_865 ();
 sg13g2_fill_1 FILLER_51_867 ();
 sg13g2_fill_1 FILLER_51_877 ();
 sg13g2_decap_4 FILLER_51_888 ();
 sg13g2_fill_1 FILLER_51_908 ();
 sg13g2_decap_4 FILLER_51_915 ();
 sg13g2_decap_4 FILLER_51_924 ();
 sg13g2_fill_1 FILLER_51_928 ();
 sg13g2_decap_8 FILLER_51_934 ();
 sg13g2_decap_8 FILLER_51_941 ();
 sg13g2_fill_1 FILLER_51_948 ();
 sg13g2_fill_2 FILLER_51_956 ();
 sg13g2_fill_2 FILLER_51_979 ();
 sg13g2_decap_4 FILLER_51_985 ();
 sg13g2_fill_2 FILLER_51_989 ();
 sg13g2_fill_2 FILLER_51_1001 ();
 sg13g2_decap_8 FILLER_51_1016 ();
 sg13g2_fill_2 FILLER_51_1023 ();
 sg13g2_fill_1 FILLER_51_1025 ();
 sg13g2_decap_4 FILLER_51_1030 ();
 sg13g2_fill_2 FILLER_51_1034 ();
 sg13g2_decap_8 FILLER_51_1040 ();
 sg13g2_decap_8 FILLER_51_1047 ();
 sg13g2_decap_8 FILLER_51_1054 ();
 sg13g2_decap_8 FILLER_51_1061 ();
 sg13g2_decap_8 FILLER_51_1068 ();
 sg13g2_fill_2 FILLER_51_1075 ();
 sg13g2_fill_2 FILLER_51_1101 ();
 sg13g2_fill_2 FILLER_51_1109 ();
 sg13g2_decap_8 FILLER_51_1126 ();
 sg13g2_decap_8 FILLER_51_1133 ();
 sg13g2_decap_4 FILLER_51_1140 ();
 sg13g2_fill_1 FILLER_51_1144 ();
 sg13g2_fill_2 FILLER_51_1148 ();
 sg13g2_decap_4 FILLER_51_1156 ();
 sg13g2_fill_2 FILLER_51_1160 ();
 sg13g2_decap_8 FILLER_51_1170 ();
 sg13g2_decap_4 FILLER_51_1177 ();
 sg13g2_fill_2 FILLER_51_1203 ();
 sg13g2_fill_1 FILLER_51_1231 ();
 sg13g2_fill_1 FILLER_51_1263 ();
 sg13g2_fill_2 FILLER_51_1308 ();
 sg13g2_decap_8 FILLER_51_1345 ();
 sg13g2_decap_8 FILLER_51_1352 ();
 sg13g2_decap_8 FILLER_51_1359 ();
 sg13g2_fill_2 FILLER_51_1366 ();
 sg13g2_decap_8 FILLER_51_1403 ();
 sg13g2_decap_4 FILLER_51_1410 ();
 sg13g2_fill_2 FILLER_51_1418 ();
 sg13g2_fill_1 FILLER_51_1420 ();
 sg13g2_decap_8 FILLER_51_1425 ();
 sg13g2_fill_1 FILLER_51_1432 ();
 sg13g2_fill_1 FILLER_51_1441 ();
 sg13g2_decap_8 FILLER_51_1446 ();
 sg13g2_decap_8 FILLER_51_1453 ();
 sg13g2_decap_8 FILLER_51_1466 ();
 sg13g2_fill_2 FILLER_51_1473 ();
 sg13g2_fill_2 FILLER_51_1501 ();
 sg13g2_fill_1 FILLER_51_1503 ();
 sg13g2_decap_8 FILLER_51_1509 ();
 sg13g2_decap_4 FILLER_51_1516 ();
 sg13g2_fill_2 FILLER_51_1520 ();
 sg13g2_fill_2 FILLER_51_1592 ();
 sg13g2_fill_2 FILLER_51_1606 ();
 sg13g2_fill_1 FILLER_51_1608 ();
 sg13g2_decap_8 FILLER_51_1613 ();
 sg13g2_fill_2 FILLER_51_1627 ();
 sg13g2_fill_2 FILLER_51_1638 ();
 sg13g2_fill_1 FILLER_51_1648 ();
 sg13g2_fill_1 FILLER_51_1654 ();
 sg13g2_decap_8 FILLER_51_1681 ();
 sg13g2_fill_2 FILLER_51_1688 ();
 sg13g2_fill_1 FILLER_51_1690 ();
 sg13g2_decap_8 FILLER_51_1699 ();
 sg13g2_decap_4 FILLER_51_1706 ();
 sg13g2_fill_1 FILLER_51_1710 ();
 sg13g2_fill_2 FILLER_51_1716 ();
 sg13g2_decap_4 FILLER_51_1724 ();
 sg13g2_fill_1 FILLER_51_1728 ();
 sg13g2_decap_8 FILLER_51_1733 ();
 sg13g2_decap_8 FILLER_51_1740 ();
 sg13g2_decap_8 FILLER_51_1747 ();
 sg13g2_fill_2 FILLER_51_1754 ();
 sg13g2_fill_2 FILLER_51_1761 ();
 sg13g2_fill_2 FILLER_51_1767 ();
 sg13g2_fill_1 FILLER_51_1778 ();
 sg13g2_fill_1 FILLER_51_1805 ();
 sg13g2_fill_1 FILLER_51_1832 ();
 sg13g2_decap_8 FILLER_51_1838 ();
 sg13g2_decap_4 FILLER_51_1845 ();
 sg13g2_fill_2 FILLER_51_1854 ();
 sg13g2_fill_2 FILLER_51_1861 ();
 sg13g2_fill_2 FILLER_51_1867 ();
 sg13g2_fill_2 FILLER_51_1874 ();
 sg13g2_fill_1 FILLER_51_1881 ();
 sg13g2_fill_1 FILLER_51_1895 ();
 sg13g2_fill_2 FILLER_51_1905 ();
 sg13g2_fill_1 FILLER_51_1922 ();
 sg13g2_decap_4 FILLER_51_1938 ();
 sg13g2_fill_2 FILLER_51_1982 ();
 sg13g2_fill_1 FILLER_51_1984 ();
 sg13g2_fill_2 FILLER_51_1994 ();
 sg13g2_fill_1 FILLER_51_1996 ();
 sg13g2_decap_8 FILLER_51_2006 ();
 sg13g2_decap_8 FILLER_51_2013 ();
 sg13g2_fill_2 FILLER_51_2020 ();
 sg13g2_decap_8 FILLER_51_2026 ();
 sg13g2_decap_8 FILLER_51_2033 ();
 sg13g2_decap_8 FILLER_51_2049 ();
 sg13g2_decap_4 FILLER_51_2056 ();
 sg13g2_fill_2 FILLER_51_2060 ();
 sg13g2_fill_2 FILLER_51_2075 ();
 sg13g2_decap_4 FILLER_51_2116 ();
 sg13g2_decap_8 FILLER_51_2123 ();
 sg13g2_decap_8 FILLER_51_2130 ();
 sg13g2_fill_2 FILLER_51_2137 ();
 sg13g2_fill_1 FILLER_51_2144 ();
 sg13g2_decap_8 FILLER_51_2157 ();
 sg13g2_fill_2 FILLER_51_2164 ();
 sg13g2_fill_1 FILLER_51_2166 ();
 sg13g2_decap_4 FILLER_51_2172 ();
 sg13g2_decap_8 FILLER_51_2181 ();
 sg13g2_fill_2 FILLER_51_2192 ();
 sg13g2_decap_4 FILLER_51_2198 ();
 sg13g2_fill_2 FILLER_51_2202 ();
 sg13g2_fill_2 FILLER_51_2252 ();
 sg13g2_fill_1 FILLER_51_2254 ();
 sg13g2_fill_2 FILLER_51_2259 ();
 sg13g2_fill_2 FILLER_51_2287 ();
 sg13g2_fill_1 FILLER_51_2289 ();
 sg13g2_decap_8 FILLER_51_2316 ();
 sg13g2_decap_4 FILLER_51_2381 ();
 sg13g2_fill_2 FILLER_51_2385 ();
 sg13g2_fill_1 FILLER_51_2392 ();
 sg13g2_fill_2 FILLER_51_2397 ();
 sg13g2_fill_1 FILLER_51_2399 ();
 sg13g2_decap_8 FILLER_51_2429 ();
 sg13g2_fill_2 FILLER_51_2436 ();
 sg13g2_decap_8 FILLER_51_2442 ();
 sg13g2_decap_4 FILLER_51_2449 ();
 sg13g2_fill_2 FILLER_51_2495 ();
 sg13g2_fill_1 FILLER_51_2497 ();
 sg13g2_fill_2 FILLER_51_2501 ();
 sg13g2_fill_2 FILLER_51_2518 ();
 sg13g2_decap_8 FILLER_51_2541 ();
 sg13g2_fill_1 FILLER_51_2553 ();
 sg13g2_fill_2 FILLER_51_2580 ();
 sg13g2_fill_2 FILLER_51_2587 ();
 sg13g2_fill_2 FILLER_51_2593 ();
 sg13g2_fill_1 FILLER_51_2595 ();
 sg13g2_fill_2 FILLER_51_2601 ();
 sg13g2_fill_1 FILLER_51_2603 ();
 sg13g2_decap_8 FILLER_51_2630 ();
 sg13g2_decap_8 FILLER_51_2637 ();
 sg13g2_decap_8 FILLER_51_2644 ();
 sg13g2_decap_8 FILLER_51_2651 ();
 sg13g2_decap_8 FILLER_51_2658 ();
 sg13g2_decap_4 FILLER_51_2665 ();
 sg13g2_fill_1 FILLER_51_2669 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_4 FILLER_52_21 ();
 sg13g2_fill_2 FILLER_52_25 ();
 sg13g2_fill_2 FILLER_52_57 ();
 sg13g2_decap_8 FILLER_52_62 ();
 sg13g2_decap_8 FILLER_52_69 ();
 sg13g2_decap_8 FILLER_52_76 ();
 sg13g2_decap_4 FILLER_52_83 ();
 sg13g2_fill_1 FILLER_52_91 ();
 sg13g2_fill_1 FILLER_52_107 ();
 sg13g2_decap_4 FILLER_52_128 ();
 sg13g2_fill_2 FILLER_52_132 ();
 sg13g2_fill_1 FILLER_52_152 ();
 sg13g2_fill_1 FILLER_52_180 ();
 sg13g2_fill_1 FILLER_52_186 ();
 sg13g2_decap_8 FILLER_52_201 ();
 sg13g2_decap_4 FILLER_52_208 ();
 sg13g2_decap_8 FILLER_52_276 ();
 sg13g2_fill_1 FILLER_52_283 ();
 sg13g2_decap_8 FILLER_52_347 ();
 sg13g2_decap_8 FILLER_52_354 ();
 sg13g2_fill_1 FILLER_52_370 ();
 sg13g2_fill_2 FILLER_52_376 ();
 sg13g2_fill_1 FILLER_52_378 ();
 sg13g2_decap_4 FILLER_52_388 ();
 sg13g2_fill_1 FILLER_52_396 ();
 sg13g2_decap_8 FILLER_52_438 ();
 sg13g2_decap_4 FILLER_52_445 ();
 sg13g2_fill_1 FILLER_52_449 ();
 sg13g2_decap_4 FILLER_52_453 ();
 sg13g2_fill_2 FILLER_52_457 ();
 sg13g2_decap_8 FILLER_52_465 ();
 sg13g2_decap_8 FILLER_52_472 ();
 sg13g2_fill_2 FILLER_52_479 ();
 sg13g2_fill_1 FILLER_52_481 ();
 sg13g2_fill_1 FILLER_52_495 ();
 sg13g2_fill_2 FILLER_52_544 ();
 sg13g2_fill_1 FILLER_52_546 ();
 sg13g2_fill_2 FILLER_52_551 ();
 sg13g2_decap_8 FILLER_52_558 ();
 sg13g2_fill_1 FILLER_52_565 ();
 sg13g2_decap_8 FILLER_52_606 ();
 sg13g2_decap_8 FILLER_52_613 ();
 sg13g2_decap_8 FILLER_52_620 ();
 sg13g2_decap_8 FILLER_52_627 ();
 sg13g2_decap_8 FILLER_52_644 ();
 sg13g2_fill_1 FILLER_52_655 ();
 sg13g2_decap_8 FILLER_52_670 ();
 sg13g2_decap_4 FILLER_52_677 ();
 sg13g2_fill_2 FILLER_52_681 ();
 sg13g2_fill_2 FILLER_52_715 ();
 sg13g2_fill_1 FILLER_52_717 ();
 sg13g2_decap_4 FILLER_52_723 ();
 sg13g2_fill_2 FILLER_52_727 ();
 sg13g2_decap_4 FILLER_52_733 ();
 sg13g2_fill_1 FILLER_52_737 ();
 sg13g2_decap_8 FILLER_52_743 ();
 sg13g2_fill_1 FILLER_52_750 ();
 sg13g2_fill_1 FILLER_52_756 ();
 sg13g2_fill_1 FILLER_52_761 ();
 sg13g2_fill_2 FILLER_52_765 ();
 sg13g2_decap_8 FILLER_52_774 ();
 sg13g2_decap_8 FILLER_52_781 ();
 sg13g2_decap_8 FILLER_52_788 ();
 sg13g2_fill_1 FILLER_52_795 ();
 sg13g2_fill_2 FILLER_52_804 ();
 sg13g2_fill_1 FILLER_52_806 ();
 sg13g2_fill_2 FILLER_52_832 ();
 sg13g2_decap_8 FILLER_52_845 ();
 sg13g2_decap_8 FILLER_52_852 ();
 sg13g2_decap_8 FILLER_52_866 ();
 sg13g2_decap_8 FILLER_52_873 ();
 sg13g2_fill_2 FILLER_52_880 ();
 sg13g2_fill_2 FILLER_52_887 ();
 sg13g2_decap_4 FILLER_52_894 ();
 sg13g2_decap_8 FILLER_52_908 ();
 sg13g2_decap_8 FILLER_52_915 ();
 sg13g2_decap_8 FILLER_52_922 ();
 sg13g2_decap_8 FILLER_52_929 ();
 sg13g2_decap_4 FILLER_52_936 ();
 sg13g2_fill_1 FILLER_52_940 ();
 sg13g2_decap_8 FILLER_52_990 ();
 sg13g2_fill_1 FILLER_52_997 ();
 sg13g2_decap_8 FILLER_52_1006 ();
 sg13g2_fill_2 FILLER_52_1018 ();
 sg13g2_fill_2 FILLER_52_1030 ();
 sg13g2_fill_2 FILLER_52_1058 ();
 sg13g2_fill_1 FILLER_52_1060 ();
 sg13g2_fill_2 FILLER_52_1069 ();
 sg13g2_fill_1 FILLER_52_1071 ();
 sg13g2_decap_8 FILLER_52_1135 ();
 sg13g2_fill_2 FILLER_52_1142 ();
 sg13g2_fill_1 FILLER_52_1144 ();
 sg13g2_fill_1 FILLER_52_1154 ();
 sg13g2_fill_2 FILLER_52_1181 ();
 sg13g2_fill_1 FILLER_52_1183 ();
 sg13g2_fill_2 FILLER_52_1209 ();
 sg13g2_fill_2 FILLER_52_1288 ();
 sg13g2_fill_1 FILLER_52_1300 ();
 sg13g2_fill_2 FILLER_52_1307 ();
 sg13g2_decap_8 FILLER_52_1335 ();
 sg13g2_fill_2 FILLER_52_1342 ();
 sg13g2_fill_1 FILLER_52_1344 ();
 sg13g2_fill_2 FILLER_52_1384 ();
 sg13g2_fill_2 FILLER_52_1401 ();
 sg13g2_decap_4 FILLER_52_1414 ();
 sg13g2_decap_4 FILLER_52_1422 ();
 sg13g2_decap_4 FILLER_52_1438 ();
 sg13g2_fill_1 FILLER_52_1442 ();
 sg13g2_fill_2 FILLER_52_1447 ();
 sg13g2_fill_1 FILLER_52_1449 ();
 sg13g2_fill_2 FILLER_52_1454 ();
 sg13g2_fill_1 FILLER_52_1456 ();
 sg13g2_decap_4 FILLER_52_1466 ();
 sg13g2_decap_8 FILLER_52_1488 ();
 sg13g2_fill_2 FILLER_52_1495 ();
 sg13g2_decap_4 FILLER_52_1509 ();
 sg13g2_decap_8 FILLER_52_1517 ();
 sg13g2_fill_1 FILLER_52_1524 ();
 sg13g2_decap_8 FILLER_52_1539 ();
 sg13g2_fill_2 FILLER_52_1546 ();
 sg13g2_fill_1 FILLER_52_1548 ();
 sg13g2_decap_4 FILLER_52_1623 ();
 sg13g2_fill_2 FILLER_52_1627 ();
 sg13g2_decap_8 FILLER_52_1666 ();
 sg13g2_decap_8 FILLER_52_1673 ();
 sg13g2_decap_8 FILLER_52_1680 ();
 sg13g2_decap_8 FILLER_52_1687 ();
 sg13g2_decap_8 FILLER_52_1694 ();
 sg13g2_decap_4 FILLER_52_1701 ();
 sg13g2_fill_1 FILLER_52_1705 ();
 sg13g2_fill_1 FILLER_52_1711 ();
 sg13g2_decap_8 FILLER_52_1748 ();
 sg13g2_decap_8 FILLER_52_1755 ();
 sg13g2_decap_4 FILLER_52_1762 ();
 sg13g2_fill_2 FILLER_52_1766 ();
 sg13g2_decap_4 FILLER_52_1771 ();
 sg13g2_fill_1 FILLER_52_1775 ();
 sg13g2_decap_8 FILLER_52_1779 ();
 sg13g2_fill_1 FILLER_52_1786 ();
 sg13g2_fill_1 FILLER_52_1792 ();
 sg13g2_decap_4 FILLER_52_1797 ();
 sg13g2_fill_1 FILLER_52_1801 ();
 sg13g2_decap_8 FILLER_52_1836 ();
 sg13g2_decap_8 FILLER_52_1843 ();
 sg13g2_decap_4 FILLER_52_1891 ();
 sg13g2_fill_2 FILLER_52_1905 ();
 sg13g2_fill_1 FILLER_52_1907 ();
 sg13g2_fill_2 FILLER_52_1912 ();
 sg13g2_fill_1 FILLER_52_1914 ();
 sg13g2_fill_1 FILLER_52_1925 ();
 sg13g2_fill_1 FILLER_52_1941 ();
 sg13g2_fill_1 FILLER_52_1981 ();
 sg13g2_fill_2 FILLER_52_1991 ();
 sg13g2_fill_1 FILLER_52_1993 ();
 sg13g2_fill_1 FILLER_52_2006 ();
 sg13g2_fill_1 FILLER_52_2036 ();
 sg13g2_fill_1 FILLER_52_2046 ();
 sg13g2_decap_8 FILLER_52_2052 ();
 sg13g2_decap_8 FILLER_52_2059 ();
 sg13g2_decap_8 FILLER_52_2066 ();
 sg13g2_decap_4 FILLER_52_2073 ();
 sg13g2_fill_1 FILLER_52_2077 ();
 sg13g2_decap_8 FILLER_52_2083 ();
 sg13g2_fill_2 FILLER_52_2090 ();
 sg13g2_fill_2 FILLER_52_2096 ();
 sg13g2_fill_1 FILLER_52_2098 ();
 sg13g2_decap_8 FILLER_52_2112 ();
 sg13g2_decap_8 FILLER_52_2119 ();
 sg13g2_decap_8 FILLER_52_2126 ();
 sg13g2_decap_8 FILLER_52_2133 ();
 sg13g2_fill_2 FILLER_52_2140 ();
 sg13g2_fill_2 FILLER_52_2150 ();
 sg13g2_decap_8 FILLER_52_2178 ();
 sg13g2_decap_8 FILLER_52_2185 ();
 sg13g2_decap_4 FILLER_52_2192 ();
 sg13g2_decap_4 FILLER_52_2237 ();
 sg13g2_fill_1 FILLER_52_2241 ();
 sg13g2_fill_2 FILLER_52_2246 ();
 sg13g2_fill_1 FILLER_52_2260 ();
 sg13g2_fill_2 FILLER_52_2290 ();
 sg13g2_decap_8 FILLER_52_2335 ();
 sg13g2_fill_2 FILLER_52_2342 ();
 sg13g2_fill_2 FILLER_52_2356 ();
 sg13g2_fill_1 FILLER_52_2364 ();
 sg13g2_fill_1 FILLER_52_2370 ();
 sg13g2_fill_2 FILLER_52_2384 ();
 sg13g2_fill_1 FILLER_52_2391 ();
 sg13g2_fill_2 FILLER_52_2395 ();
 sg13g2_fill_2 FILLER_52_2450 ();
 sg13g2_fill_1 FILLER_52_2452 ();
 sg13g2_decap_8 FILLER_52_2488 ();
 sg13g2_decap_8 FILLER_52_2495 ();
 sg13g2_decap_4 FILLER_52_2502 ();
 sg13g2_fill_1 FILLER_52_2575 ();
 sg13g2_decap_8 FILLER_52_2602 ();
 sg13g2_decap_8 FILLER_52_2609 ();
 sg13g2_decap_8 FILLER_52_2616 ();
 sg13g2_decap_8 FILLER_52_2623 ();
 sg13g2_decap_8 FILLER_52_2630 ();
 sg13g2_decap_8 FILLER_52_2637 ();
 sg13g2_decap_8 FILLER_52_2644 ();
 sg13g2_decap_8 FILLER_52_2651 ();
 sg13g2_decap_8 FILLER_52_2658 ();
 sg13g2_decap_4 FILLER_52_2665 ();
 sg13g2_fill_1 FILLER_52_2669 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_4 FILLER_53_7 ();
 sg13g2_fill_2 FILLER_53_11 ();
 sg13g2_fill_2 FILLER_53_18 ();
 sg13g2_fill_1 FILLER_53_20 ();
 sg13g2_decap_8 FILLER_53_29 ();
 sg13g2_decap_8 FILLER_53_36 ();
 sg13g2_fill_1 FILLER_53_43 ();
 sg13g2_fill_2 FILLER_53_52 ();
 sg13g2_fill_2 FILLER_53_92 ();
 sg13g2_fill_1 FILLER_53_97 ();
 sg13g2_fill_2 FILLER_53_111 ();
 sg13g2_fill_1 FILLER_53_113 ();
 sg13g2_fill_2 FILLER_53_120 ();
 sg13g2_decap_4 FILLER_53_131 ();
 sg13g2_fill_2 FILLER_53_166 ();
 sg13g2_fill_2 FILLER_53_189 ();
 sg13g2_fill_1 FILLER_53_191 ();
 sg13g2_fill_1 FILLER_53_197 ();
 sg13g2_fill_2 FILLER_53_234 ();
 sg13g2_fill_1 FILLER_53_236 ();
 sg13g2_decap_8 FILLER_53_242 ();
 sg13g2_decap_4 FILLER_53_249 ();
 sg13g2_fill_2 FILLER_53_253 ();
 sg13g2_decap_4 FILLER_53_258 ();
 sg13g2_decap_8 FILLER_53_265 ();
 sg13g2_decap_8 FILLER_53_272 ();
 sg13g2_decap_8 FILLER_53_279 ();
 sg13g2_decap_4 FILLER_53_286 ();
 sg13g2_fill_2 FILLER_53_290 ();
 sg13g2_decap_4 FILLER_53_295 ();
 sg13g2_fill_2 FILLER_53_317 ();
 sg13g2_fill_1 FILLER_53_319 ();
 sg13g2_decap_4 FILLER_53_326 ();
 sg13g2_fill_2 FILLER_53_330 ();
 sg13g2_fill_2 FILLER_53_335 ();
 sg13g2_decap_8 FILLER_53_346 ();
 sg13g2_fill_1 FILLER_53_353 ();
 sg13g2_fill_2 FILLER_53_382 ();
 sg13g2_fill_2 FILLER_53_389 ();
 sg13g2_fill_1 FILLER_53_391 ();
 sg13g2_fill_1 FILLER_53_400 ();
 sg13g2_fill_2 FILLER_53_427 ();
 sg13g2_fill_1 FILLER_53_429 ();
 sg13g2_fill_1 FILLER_53_440 ();
 sg13g2_decap_8 FILLER_53_444 ();
 sg13g2_decap_8 FILLER_53_451 ();
 sg13g2_decap_8 FILLER_53_458 ();
 sg13g2_fill_2 FILLER_53_469 ();
 sg13g2_fill_1 FILLER_53_471 ();
 sg13g2_decap_4 FILLER_53_480 ();
 sg13g2_decap_4 FILLER_53_488 ();
 sg13g2_fill_1 FILLER_53_496 ();
 sg13g2_fill_1 FILLER_53_516 ();
 sg13g2_fill_1 FILLER_53_522 ();
 sg13g2_fill_2 FILLER_53_532 ();
 sg13g2_decap_8 FILLER_53_539 ();
 sg13g2_decap_8 FILLER_53_546 ();
 sg13g2_fill_2 FILLER_53_553 ();
 sg13g2_decap_8 FILLER_53_564 ();
 sg13g2_fill_1 FILLER_53_571 ();
 sg13g2_decap_8 FILLER_53_576 ();
 sg13g2_fill_2 FILLER_53_583 ();
 sg13g2_fill_1 FILLER_53_629 ();
 sg13g2_fill_1 FILLER_53_640 ();
 sg13g2_fill_1 FILLER_53_663 ();
 sg13g2_decap_8 FILLER_53_668 ();
 sg13g2_decap_8 FILLER_53_675 ();
 sg13g2_decap_4 FILLER_53_682 ();
 sg13g2_fill_2 FILLER_53_686 ();
 sg13g2_decap_8 FILLER_53_696 ();
 sg13g2_fill_1 FILLER_53_703 ();
 sg13g2_decap_8 FILLER_53_709 ();
 sg13g2_decap_8 FILLER_53_716 ();
 sg13g2_decap_8 FILLER_53_723 ();
 sg13g2_decap_4 FILLER_53_730 ();
 sg13g2_fill_1 FILLER_53_734 ();
 sg13g2_decap_4 FILLER_53_742 ();
 sg13g2_fill_2 FILLER_53_746 ();
 sg13g2_decap_8 FILLER_53_765 ();
 sg13g2_decap_8 FILLER_53_772 ();
 sg13g2_decap_8 FILLER_53_779 ();
 sg13g2_decap_4 FILLER_53_786 ();
 sg13g2_fill_2 FILLER_53_812 ();
 sg13g2_fill_2 FILLER_53_831 ();
 sg13g2_fill_1 FILLER_53_833 ();
 sg13g2_decap_8 FILLER_53_851 ();
 sg13g2_decap_8 FILLER_53_858 ();
 sg13g2_decap_8 FILLER_53_865 ();
 sg13g2_decap_4 FILLER_53_872 ();
 sg13g2_fill_1 FILLER_53_876 ();
 sg13g2_fill_1 FILLER_53_882 ();
 sg13g2_fill_1 FILLER_53_888 ();
 sg13g2_decap_4 FILLER_53_893 ();
 sg13g2_fill_1 FILLER_53_901 ();
 sg13g2_decap_8 FILLER_53_905 ();
 sg13g2_decap_8 FILLER_53_912 ();
 sg13g2_fill_1 FILLER_53_919 ();
 sg13g2_decap_4 FILLER_53_924 ();
 sg13g2_decap_8 FILLER_53_934 ();
 sg13g2_decap_8 FILLER_53_941 ();
 sg13g2_fill_2 FILLER_53_948 ();
 sg13g2_fill_1 FILLER_53_950 ();
 sg13g2_fill_2 FILLER_53_955 ();
 sg13g2_fill_1 FILLER_53_957 ();
 sg13g2_decap_8 FILLER_53_974 ();
 sg13g2_decap_8 FILLER_53_981 ();
 sg13g2_fill_1 FILLER_53_988 ();
 sg13g2_decap_8 FILLER_53_1025 ();
 sg13g2_fill_1 FILLER_53_1032 ();
 sg13g2_fill_2 FILLER_53_1059 ();
 sg13g2_fill_1 FILLER_53_1061 ();
 sg13g2_decap_8 FILLER_53_1110 ();
 sg13g2_decap_8 FILLER_53_1117 ();
 sg13g2_decap_8 FILLER_53_1124 ();
 sg13g2_decap_8 FILLER_53_1131 ();
 sg13g2_decap_8 FILLER_53_1138 ();
 sg13g2_fill_1 FILLER_53_1145 ();
 sg13g2_fill_1 FILLER_53_1151 ();
 sg13g2_fill_2 FILLER_53_1156 ();
 sg13g2_fill_2 FILLER_53_1184 ();
 sg13g2_fill_1 FILLER_53_1239 ();
 sg13g2_decap_8 FILLER_53_1307 ();
 sg13g2_decap_8 FILLER_53_1314 ();
 sg13g2_decap_4 FILLER_53_1321 ();
 sg13g2_decap_8 FILLER_53_1331 ();
 sg13g2_decap_8 FILLER_53_1338 ();
 sg13g2_decap_8 FILLER_53_1345 ();
 sg13g2_decap_8 FILLER_53_1352 ();
 sg13g2_fill_2 FILLER_53_1359 ();
 sg13g2_decap_8 FILLER_53_1366 ();
 sg13g2_fill_1 FILLER_53_1373 ();
 sg13g2_fill_2 FILLER_53_1392 ();
 sg13g2_fill_2 FILLER_53_1402 ();
 sg13g2_fill_1 FILLER_53_1404 ();
 sg13g2_fill_1 FILLER_53_1415 ();
 sg13g2_fill_1 FILLER_53_1459 ();
 sg13g2_fill_2 FILLER_53_1475 ();
 sg13g2_fill_1 FILLER_53_1477 ();
 sg13g2_fill_2 FILLER_53_1486 ();
 sg13g2_fill_2 FILLER_53_1501 ();
 sg13g2_fill_1 FILLER_53_1503 ();
 sg13g2_fill_2 FILLER_53_1510 ();
 sg13g2_fill_1 FILLER_53_1512 ();
 sg13g2_fill_2 FILLER_53_1539 ();
 sg13g2_fill_1 FILLER_53_1592 ();
 sg13g2_fill_1 FILLER_53_1606 ();
 sg13g2_fill_1 FILLER_53_1638 ();
 sg13g2_decap_8 FILLER_53_1659 ();
 sg13g2_decap_8 FILLER_53_1666 ();
 sg13g2_decap_8 FILLER_53_1673 ();
 sg13g2_decap_4 FILLER_53_1680 ();
 sg13g2_decap_8 FILLER_53_1697 ();
 sg13g2_decap_4 FILLER_53_1704 ();
 sg13g2_fill_2 FILLER_53_1708 ();
 sg13g2_fill_2 FILLER_53_1729 ();
 sg13g2_decap_4 FILLER_53_1762 ();
 sg13g2_fill_2 FILLER_53_1766 ();
 sg13g2_decap_8 FILLER_53_1777 ();
 sg13g2_decap_8 FILLER_53_1784 ();
 sg13g2_decap_8 FILLER_53_1791 ();
 sg13g2_decap_8 FILLER_53_1798 ();
 sg13g2_decap_4 FILLER_53_1805 ();
 sg13g2_decap_8 FILLER_53_1821 ();
 sg13g2_decap_8 FILLER_53_1828 ();
 sg13g2_decap_8 FILLER_53_1835 ();
 sg13g2_decap_8 FILLER_53_1842 ();
 sg13g2_fill_2 FILLER_53_1849 ();
 sg13g2_fill_1 FILLER_53_1877 ();
 sg13g2_fill_2 FILLER_53_1887 ();
 sg13g2_fill_1 FILLER_53_1904 ();
 sg13g2_fill_2 FILLER_53_1940 ();
 sg13g2_fill_1 FILLER_53_1942 ();
 sg13g2_fill_2 FILLER_53_1968 ();
 sg13g2_fill_2 FILLER_53_1996 ();
 sg13g2_fill_1 FILLER_53_2026 ();
 sg13g2_decap_8 FILLER_53_2053 ();
 sg13g2_decap_8 FILLER_53_2068 ();
 sg13g2_fill_1 FILLER_53_2075 ();
 sg13g2_fill_1 FILLER_53_2106 ();
 sg13g2_decap_8 FILLER_53_2112 ();
 sg13g2_decap_8 FILLER_53_2119 ();
 sg13g2_decap_8 FILLER_53_2126 ();
 sg13g2_fill_2 FILLER_53_2133 ();
 sg13g2_fill_1 FILLER_53_2135 ();
 sg13g2_decap_4 FILLER_53_2141 ();
 sg13g2_fill_1 FILLER_53_2145 ();
 sg13g2_fill_2 FILLER_53_2150 ();
 sg13g2_fill_1 FILLER_53_2152 ();
 sg13g2_fill_1 FILLER_53_2157 ();
 sg13g2_decap_4 FILLER_53_2166 ();
 sg13g2_fill_2 FILLER_53_2170 ();
 sg13g2_fill_2 FILLER_53_2176 ();
 sg13g2_fill_1 FILLER_53_2178 ();
 sg13g2_fill_2 FILLER_53_2183 ();
 sg13g2_fill_1 FILLER_53_2201 ();
 sg13g2_decap_8 FILLER_53_2207 ();
 sg13g2_decap_4 FILLER_53_2214 ();
 sg13g2_decap_4 FILLER_53_2223 ();
 sg13g2_fill_2 FILLER_53_2227 ();
 sg13g2_fill_2 FILLER_53_2267 ();
 sg13g2_decap_8 FILLER_53_2295 ();
 sg13g2_fill_2 FILLER_53_2302 ();
 sg13g2_decap_8 FILLER_53_2308 ();
 sg13g2_decap_8 FILLER_53_2315 ();
 sg13g2_fill_2 FILLER_53_2322 ();
 sg13g2_fill_1 FILLER_53_2324 ();
 sg13g2_decap_4 FILLER_53_2333 ();
 sg13g2_fill_1 FILLER_53_2342 ();
 sg13g2_fill_1 FILLER_53_2363 ();
 sg13g2_fill_2 FILLER_53_2373 ();
 sg13g2_decap_8 FILLER_53_2405 ();
 sg13g2_fill_1 FILLER_53_2412 ();
 sg13g2_fill_1 FILLER_53_2419 ();
 sg13g2_fill_2 FILLER_53_2435 ();
 sg13g2_fill_2 FILLER_53_2499 ();
 sg13g2_fill_1 FILLER_53_2501 ();
 sg13g2_fill_1 FILLER_53_2507 ();
 sg13g2_fill_1 FILLER_53_2522 ();
 sg13g2_fill_1 FILLER_53_2535 ();
 sg13g2_fill_2 FILLER_53_2541 ();
 sg13g2_decap_8 FILLER_53_2608 ();
 sg13g2_decap_8 FILLER_53_2615 ();
 sg13g2_fill_2 FILLER_53_2622 ();
 sg13g2_decap_8 FILLER_53_2654 ();
 sg13g2_decap_8 FILLER_53_2661 ();
 sg13g2_fill_2 FILLER_53_2668 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_32 ();
 sg13g2_decap_4 FILLER_54_39 ();
 sg13g2_fill_1 FILLER_54_49 ();
 sg13g2_fill_1 FILLER_54_58 ();
 sg13g2_decap_4 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_75 ();
 sg13g2_fill_1 FILLER_54_82 ();
 sg13g2_fill_2 FILLER_54_114 ();
 sg13g2_fill_1 FILLER_54_116 ();
 sg13g2_decap_4 FILLER_54_122 ();
 sg13g2_fill_1 FILLER_54_126 ();
 sg13g2_decap_8 FILLER_54_131 ();
 sg13g2_fill_2 FILLER_54_160 ();
 sg13g2_decap_8 FILLER_54_216 ();
 sg13g2_decap_8 FILLER_54_223 ();
 sg13g2_decap_8 FILLER_54_230 ();
 sg13g2_decap_8 FILLER_54_237 ();
 sg13g2_decap_8 FILLER_54_244 ();
 sg13g2_decap_8 FILLER_54_251 ();
 sg13g2_decap_8 FILLER_54_258 ();
 sg13g2_decap_8 FILLER_54_265 ();
 sg13g2_decap_8 FILLER_54_272 ();
 sg13g2_decap_8 FILLER_54_279 ();
 sg13g2_decap_8 FILLER_54_286 ();
 sg13g2_decap_4 FILLER_54_293 ();
 sg13g2_fill_1 FILLER_54_297 ();
 sg13g2_decap_8 FILLER_54_312 ();
 sg13g2_decap_8 FILLER_54_319 ();
 sg13g2_decap_8 FILLER_54_326 ();
 sg13g2_fill_2 FILLER_54_337 ();
 sg13g2_fill_2 FILLER_54_344 ();
 sg13g2_fill_1 FILLER_54_346 ();
 sg13g2_decap_4 FILLER_54_356 ();
 sg13g2_fill_1 FILLER_54_396 ();
 sg13g2_fill_1 FILLER_54_415 ();
 sg13g2_fill_2 FILLER_54_426 ();
 sg13g2_decap_4 FILLER_54_432 ();
 sg13g2_fill_2 FILLER_54_471 ();
 sg13g2_decap_8 FILLER_54_477 ();
 sg13g2_fill_2 FILLER_54_484 ();
 sg13g2_fill_1 FILLER_54_486 ();
 sg13g2_decap_4 FILLER_54_491 ();
 sg13g2_decap_4 FILLER_54_500 ();
 sg13g2_decap_8 FILLER_54_538 ();
 sg13g2_fill_1 FILLER_54_545 ();
 sg13g2_fill_2 FILLER_54_551 ();
 sg13g2_fill_2 FILLER_54_557 ();
 sg13g2_decap_8 FILLER_54_564 ();
 sg13g2_decap_8 FILLER_54_571 ();
 sg13g2_decap_8 FILLER_54_578 ();
 sg13g2_decap_8 FILLER_54_585 ();
 sg13g2_decap_8 FILLER_54_592 ();
 sg13g2_decap_8 FILLER_54_607 ();
 sg13g2_decap_4 FILLER_54_614 ();
 sg13g2_fill_1 FILLER_54_618 ();
 sg13g2_fill_1 FILLER_54_623 ();
 sg13g2_fill_2 FILLER_54_629 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_fill_1 FILLER_54_652 ();
 sg13g2_fill_2 FILLER_54_658 ();
 sg13g2_fill_2 FILLER_54_672 ();
 sg13g2_fill_1 FILLER_54_674 ();
 sg13g2_decap_8 FILLER_54_679 ();
 sg13g2_decap_8 FILLER_54_694 ();
 sg13g2_decap_4 FILLER_54_701 ();
 sg13g2_fill_1 FILLER_54_705 ();
 sg13g2_decap_8 FILLER_54_709 ();
 sg13g2_decap_8 FILLER_54_716 ();
 sg13g2_decap_8 FILLER_54_723 ();
 sg13g2_fill_2 FILLER_54_746 ();
 sg13g2_fill_2 FILLER_54_795 ();
 sg13g2_fill_2 FILLER_54_839 ();
 sg13g2_fill_1 FILLER_54_841 ();
 sg13g2_fill_1 FILLER_54_868 ();
 sg13g2_fill_1 FILLER_54_873 ();
 sg13g2_fill_2 FILLER_54_900 ();
 sg13g2_fill_1 FILLER_54_902 ();
 sg13g2_decap_8 FILLER_54_946 ();
 sg13g2_decap_8 FILLER_54_953 ();
 sg13g2_decap_8 FILLER_54_960 ();
 sg13g2_decap_8 FILLER_54_967 ();
 sg13g2_decap_8 FILLER_54_974 ();
 sg13g2_decap_8 FILLER_54_1000 ();
 sg13g2_decap_8 FILLER_54_1007 ();
 sg13g2_decap_8 FILLER_54_1014 ();
 sg13g2_fill_2 FILLER_54_1021 ();
 sg13g2_fill_1 FILLER_54_1023 ();
 sg13g2_decap_4 FILLER_54_1034 ();
 sg13g2_fill_1 FILLER_54_1038 ();
 sg13g2_decap_8 FILLER_54_1043 ();
 sg13g2_decap_4 FILLER_54_1050 ();
 sg13g2_fill_1 FILLER_54_1054 ();
 sg13g2_decap_8 FILLER_54_1069 ();
 sg13g2_decap_4 FILLER_54_1076 ();
 sg13g2_fill_2 FILLER_54_1088 ();
 sg13g2_fill_1 FILLER_54_1090 ();
 sg13g2_fill_1 FILLER_54_1095 ();
 sg13g2_decap_8 FILLER_54_1108 ();
 sg13g2_decap_4 FILLER_54_1128 ();
 sg13g2_fill_2 FILLER_54_1132 ();
 sg13g2_decap_8 FILLER_54_1168 ();
 sg13g2_fill_1 FILLER_54_1175 ();
 sg13g2_fill_1 FILLER_54_1228 ();
 sg13g2_fill_2 FILLER_54_1263 ();
 sg13g2_decap_8 FILLER_54_1319 ();
 sg13g2_decap_8 FILLER_54_1326 ();
 sg13g2_decap_8 FILLER_54_1333 ();
 sg13g2_decap_8 FILLER_54_1340 ();
 sg13g2_fill_2 FILLER_54_1347 ();
 sg13g2_fill_1 FILLER_54_1349 ();
 sg13g2_fill_2 FILLER_54_1354 ();
 sg13g2_decap_8 FILLER_54_1366 ();
 sg13g2_decap_8 FILLER_54_1373 ();
 sg13g2_fill_2 FILLER_54_1380 ();
 sg13g2_fill_1 FILLER_54_1417 ();
 sg13g2_decap_4 FILLER_54_1455 ();
 sg13g2_fill_1 FILLER_54_1459 ();
 sg13g2_fill_2 FILLER_54_1468 ();
 sg13g2_fill_1 FILLER_54_1470 ();
 sg13g2_decap_4 FILLER_54_1536 ();
 sg13g2_fill_1 FILLER_54_1540 ();
 sg13g2_fill_2 FILLER_54_1559 ();
 sg13g2_decap_8 FILLER_54_1611 ();
 sg13g2_decap_4 FILLER_54_1618 ();
 sg13g2_fill_2 FILLER_54_1622 ();
 sg13g2_decap_8 FILLER_54_1627 ();
 sg13g2_fill_2 FILLER_54_1634 ();
 sg13g2_fill_1 FILLER_54_1652 ();
 sg13g2_decap_4 FILLER_54_1663 ();
 sg13g2_fill_1 FILLER_54_1667 ();
 sg13g2_decap_8 FILLER_54_1673 ();
 sg13g2_decap_8 FILLER_54_1680 ();
 sg13g2_fill_1 FILLER_54_1696 ();
 sg13g2_decap_4 FILLER_54_1701 ();
 sg13g2_fill_2 FILLER_54_1705 ();
 sg13g2_fill_2 FILLER_54_1724 ();
 sg13g2_fill_1 FILLER_54_1739 ();
 sg13g2_fill_2 FILLER_54_1745 ();
 sg13g2_fill_2 FILLER_54_1751 ();
 sg13g2_decap_4 FILLER_54_1784 ();
 sg13g2_decap_4 FILLER_54_1801 ();
 sg13g2_fill_1 FILLER_54_1805 ();
 sg13g2_fill_2 FILLER_54_1818 ();
 sg13g2_fill_1 FILLER_54_1820 ();
 sg13g2_decap_8 FILLER_54_1834 ();
 sg13g2_decap_4 FILLER_54_1841 ();
 sg13g2_fill_2 FILLER_54_1850 ();
 sg13g2_fill_1 FILLER_54_1865 ();
 sg13g2_fill_2 FILLER_54_1871 ();
 sg13g2_fill_2 FILLER_54_1878 ();
 sg13g2_fill_2 FILLER_54_1921 ();
 sg13g2_fill_1 FILLER_54_1923 ();
 sg13g2_decap_8 FILLER_54_1933 ();
 sg13g2_decap_4 FILLER_54_1940 ();
 sg13g2_fill_1 FILLER_54_1944 ();
 sg13g2_fill_1 FILLER_54_1950 ();
 sg13g2_fill_1 FILLER_54_1955 ();
 sg13g2_fill_2 FILLER_54_1965 ();
 sg13g2_fill_1 FILLER_54_1971 ();
 sg13g2_decap_4 FILLER_54_1976 ();
 sg13g2_fill_2 FILLER_54_1984 ();
 sg13g2_fill_2 FILLER_54_1989 ();
 sg13g2_decap_8 FILLER_54_2015 ();
 sg13g2_fill_2 FILLER_54_2040 ();
 sg13g2_decap_8 FILLER_54_2107 ();
 sg13g2_decap_8 FILLER_54_2114 ();
 sg13g2_fill_1 FILLER_54_2121 ();
 sg13g2_fill_2 FILLER_54_2138 ();
 sg13g2_decap_8 FILLER_54_2166 ();
 sg13g2_decap_8 FILLER_54_2173 ();
 sg13g2_decap_8 FILLER_54_2194 ();
 sg13g2_decap_8 FILLER_54_2201 ();
 sg13g2_decap_8 FILLER_54_2208 ();
 sg13g2_decap_8 FILLER_54_2215 ();
 sg13g2_decap_8 FILLER_54_2222 ();
 sg13g2_decap_8 FILLER_54_2229 ();
 sg13g2_decap_8 FILLER_54_2236 ();
 sg13g2_decap_4 FILLER_54_2243 ();
 sg13g2_fill_1 FILLER_54_2247 ();
 sg13g2_decap_8 FILLER_54_2283 ();
 sg13g2_decap_4 FILLER_54_2290 ();
 sg13g2_fill_2 FILLER_54_2294 ();
 sg13g2_fill_1 FILLER_54_2323 ();
 sg13g2_fill_2 FILLER_54_2327 ();
 sg13g2_fill_2 FILLER_54_2355 ();
 sg13g2_fill_1 FILLER_54_2357 ();
 sg13g2_fill_1 FILLER_54_2458 ();
 sg13g2_decap_4 FILLER_54_2497 ();
 sg13g2_fill_1 FILLER_54_2501 ();
 sg13g2_decap_4 FILLER_54_2511 ();
 sg13g2_decap_8 FILLER_54_2551 ();
 sg13g2_decap_8 FILLER_54_2558 ();
 sg13g2_decap_8 FILLER_54_2565 ();
 sg13g2_fill_1 FILLER_54_2576 ();
 sg13g2_fill_2 FILLER_54_2582 ();
 sg13g2_fill_1 FILLER_54_2594 ();
 sg13g2_decap_8 FILLER_54_2604 ();
 sg13g2_decap_4 FILLER_54_2611 ();
 sg13g2_decap_4 FILLER_54_2619 ();
 sg13g2_decap_8 FILLER_54_2649 ();
 sg13g2_decap_8 FILLER_54_2656 ();
 sg13g2_decap_8 FILLER_54_2663 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_9 ();
 sg13g2_decap_4 FILLER_55_14 ();
 sg13g2_fill_1 FILLER_55_31 ();
 sg13g2_fill_1 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_87 ();
 sg13g2_decap_8 FILLER_55_94 ();
 sg13g2_decap_4 FILLER_55_101 ();
 sg13g2_fill_1 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_136 ();
 sg13g2_decap_8 FILLER_55_143 ();
 sg13g2_decap_4 FILLER_55_150 ();
 sg13g2_fill_2 FILLER_55_154 ();
 sg13g2_fill_1 FILLER_55_185 ();
 sg13g2_fill_2 FILLER_55_195 ();
 sg13g2_decap_4 FILLER_55_201 ();
 sg13g2_fill_1 FILLER_55_205 ();
 sg13g2_fill_2 FILLER_55_262 ();
 sg13g2_decap_8 FILLER_55_277 ();
 sg13g2_decap_4 FILLER_55_284 ();
 sg13g2_fill_1 FILLER_55_295 ();
 sg13g2_fill_2 FILLER_55_339 ();
 sg13g2_fill_2 FILLER_55_345 ();
 sg13g2_fill_1 FILLER_55_347 ();
 sg13g2_decap_8 FILLER_55_353 ();
 sg13g2_fill_2 FILLER_55_360 ();
 sg13g2_fill_1 FILLER_55_374 ();
 sg13g2_decap_8 FILLER_55_379 ();
 sg13g2_decap_4 FILLER_55_386 ();
 sg13g2_fill_2 FILLER_55_390 ();
 sg13g2_fill_1 FILLER_55_427 ();
 sg13g2_fill_1 FILLER_55_433 ();
 sg13g2_decap_4 FILLER_55_478 ();
 sg13g2_fill_2 FILLER_55_487 ();
 sg13g2_fill_1 FILLER_55_489 ();
 sg13g2_fill_1 FILLER_55_499 ();
 sg13g2_fill_1 FILLER_55_507 ();
 sg13g2_fill_2 FILLER_55_526 ();
 sg13g2_fill_2 FILLER_55_535 ();
 sg13g2_fill_1 FILLER_55_537 ();
 sg13g2_fill_2 FILLER_55_545 ();
 sg13g2_fill_1 FILLER_55_547 ();
 sg13g2_decap_4 FILLER_55_556 ();
 sg13g2_fill_2 FILLER_55_560 ();
 sg13g2_decap_4 FILLER_55_566 ();
 sg13g2_decap_4 FILLER_55_574 ();
 sg13g2_fill_1 FILLER_55_578 ();
 sg13g2_fill_2 FILLER_55_605 ();
 sg13g2_fill_1 FILLER_55_617 ();
 sg13g2_fill_2 FILLER_55_626 ();
 sg13g2_fill_1 FILLER_55_628 ();
 sg13g2_fill_1 FILLER_55_638 ();
 sg13g2_fill_1 FILLER_55_654 ();
 sg13g2_decap_4 FILLER_55_662 ();
 sg13g2_fill_2 FILLER_55_666 ();
 sg13g2_fill_1 FILLER_55_674 ();
 sg13g2_decap_8 FILLER_55_680 ();
 sg13g2_decap_8 FILLER_55_687 ();
 sg13g2_decap_8 FILLER_55_694 ();
 sg13g2_decap_8 FILLER_55_701 ();
 sg13g2_fill_1 FILLER_55_708 ();
 sg13g2_fill_1 FILLER_55_727 ();
 sg13g2_fill_1 FILLER_55_736 ();
 sg13g2_fill_2 FILLER_55_741 ();
 sg13g2_fill_1 FILLER_55_743 ();
 sg13g2_decap_8 FILLER_55_757 ();
 sg13g2_decap_8 FILLER_55_764 ();
 sg13g2_fill_2 FILLER_55_771 ();
 sg13g2_fill_1 FILLER_55_800 ();
 sg13g2_fill_1 FILLER_55_817 ();
 sg13g2_fill_1 FILLER_55_828 ();
 sg13g2_decap_4 FILLER_55_834 ();
 sg13g2_fill_1 FILLER_55_872 ();
 sg13g2_fill_1 FILLER_55_903 ();
 sg13g2_decap_8 FILLER_55_913 ();
 sg13g2_decap_4 FILLER_55_920 ();
 sg13g2_fill_1 FILLER_55_932 ();
 sg13g2_decap_8 FILLER_55_944 ();
 sg13g2_fill_2 FILLER_55_951 ();
 sg13g2_fill_1 FILLER_55_953 ();
 sg13g2_fill_2 FILLER_55_984 ();
 sg13g2_fill_1 FILLER_55_986 ();
 sg13g2_fill_2 FILLER_55_1054 ();
 sg13g2_fill_1 FILLER_55_1056 ();
 sg13g2_fill_2 FILLER_55_1070 ();
 sg13g2_decap_4 FILLER_55_1076 ();
 sg13g2_decap_8 FILLER_55_1097 ();
 sg13g2_fill_2 FILLER_55_1104 ();
 sg13g2_fill_1 FILLER_55_1106 ();
 sg13g2_decap_4 FILLER_55_1137 ();
 sg13g2_fill_1 FILLER_55_1206 ();
 sg13g2_decap_4 FILLER_55_1239 ();
 sg13g2_decap_4 FILLER_55_1249 ();
 sg13g2_fill_2 FILLER_55_1253 ();
 sg13g2_fill_2 FILLER_55_1261 ();
 sg13g2_decap_4 FILLER_55_1293 ();
 sg13g2_fill_2 FILLER_55_1297 ();
 sg13g2_decap_8 FILLER_55_1304 ();
 sg13g2_decap_8 FILLER_55_1311 ();
 sg13g2_decap_8 FILLER_55_1318 ();
 sg13g2_decap_8 FILLER_55_1325 ();
 sg13g2_decap_4 FILLER_55_1332 ();
 sg13g2_fill_2 FILLER_55_1336 ();
 sg13g2_decap_4 FILLER_55_1375 ();
 sg13g2_fill_2 FILLER_55_1379 ();
 sg13g2_decap_8 FILLER_55_1385 ();
 sg13g2_decap_4 FILLER_55_1404 ();
 sg13g2_fill_1 FILLER_55_1408 ();
 sg13g2_fill_2 FILLER_55_1414 ();
 sg13g2_fill_1 FILLER_55_1445 ();
 sg13g2_decap_4 FILLER_55_1472 ();
 sg13g2_fill_1 FILLER_55_1476 ();
 sg13g2_decap_4 FILLER_55_1481 ();
 sg13g2_fill_1 FILLER_55_1485 ();
 sg13g2_fill_2 FILLER_55_1499 ();
 sg13g2_fill_1 FILLER_55_1501 ();
 sg13g2_decap_8 FILLER_55_1511 ();
 sg13g2_decap_8 FILLER_55_1518 ();
 sg13g2_fill_1 FILLER_55_1534 ();
 sg13g2_fill_1 FILLER_55_1539 ();
 sg13g2_fill_1 FILLER_55_1552 ();
 sg13g2_decap_8 FILLER_55_1589 ();
 sg13g2_decap_4 FILLER_55_1596 ();
 sg13g2_fill_2 FILLER_55_1600 ();
 sg13g2_decap_4 FILLER_55_1610 ();
 sg13g2_fill_1 FILLER_55_1623 ();
 sg13g2_fill_1 FILLER_55_1629 ();
 sg13g2_decap_8 FILLER_55_1639 ();
 sg13g2_decap_8 FILLER_55_1679 ();
 sg13g2_fill_2 FILLER_55_1686 ();
 sg13g2_fill_1 FILLER_55_1688 ();
 sg13g2_fill_1 FILLER_55_1699 ();
 sg13g2_fill_2 FILLER_55_1704 ();
 sg13g2_fill_1 FILLER_55_1709 ();
 sg13g2_decap_4 FILLER_55_1765 ();
 sg13g2_fill_2 FILLER_55_1769 ();
 sg13g2_decap_4 FILLER_55_1797 ();
 sg13g2_fill_2 FILLER_55_1807 ();
 sg13g2_fill_2 FILLER_55_1819 ();
 sg13g2_fill_1 FILLER_55_1821 ();
 sg13g2_decap_8 FILLER_55_1848 ();
 sg13g2_fill_2 FILLER_55_1869 ();
 sg13g2_fill_2 FILLER_55_1875 ();
 sg13g2_fill_1 FILLER_55_1881 ();
 sg13g2_fill_2 FILLER_55_1908 ();
 sg13g2_decap_8 FILLER_55_1914 ();
 sg13g2_decap_8 FILLER_55_1921 ();
 sg13g2_decap_8 FILLER_55_1928 ();
 sg13g2_decap_8 FILLER_55_1935 ();
 sg13g2_decap_8 FILLER_55_1942 ();
 sg13g2_fill_2 FILLER_55_1949 ();
 sg13g2_decap_8 FILLER_55_1956 ();
 sg13g2_decap_8 FILLER_55_1963 ();
 sg13g2_decap_4 FILLER_55_1970 ();
 sg13g2_fill_1 FILLER_55_1974 ();
 sg13g2_decap_4 FILLER_55_2011 ();
 sg13g2_fill_1 FILLER_55_2015 ();
 sg13g2_decap_8 FILLER_55_2021 ();
 sg13g2_decap_4 FILLER_55_2028 ();
 sg13g2_fill_2 FILLER_55_2032 ();
 sg13g2_decap_8 FILLER_55_2045 ();
 sg13g2_decap_4 FILLER_55_2052 ();
 sg13g2_fill_2 FILLER_55_2056 ();
 sg13g2_fill_2 FILLER_55_2065 ();
 sg13g2_fill_1 FILLER_55_2067 ();
 sg13g2_fill_1 FILLER_55_2072 ();
 sg13g2_decap_8 FILLER_55_2096 ();
 sg13g2_decap_8 FILLER_55_2103 ();
 sg13g2_decap_8 FILLER_55_2110 ();
 sg13g2_decap_8 FILLER_55_2117 ();
 sg13g2_decap_4 FILLER_55_2124 ();
 sg13g2_decap_8 FILLER_55_2211 ();
 sg13g2_decap_8 FILLER_55_2218 ();
 sg13g2_decap_4 FILLER_55_2225 ();
 sg13g2_fill_1 FILLER_55_2229 ();
 sg13g2_fill_1 FILLER_55_2237 ();
 sg13g2_decap_4 FILLER_55_2251 ();
 sg13g2_fill_1 FILLER_55_2255 ();
 sg13g2_decap_4 FILLER_55_2261 ();
 sg13g2_decap_4 FILLER_55_2269 ();
 sg13g2_fill_1 FILLER_55_2329 ();
 sg13g2_decap_8 FILLER_55_2362 ();
 sg13g2_decap_4 FILLER_55_2369 ();
 sg13g2_fill_1 FILLER_55_2385 ();
 sg13g2_decap_8 FILLER_55_2412 ();
 sg13g2_decap_4 FILLER_55_2419 ();
 sg13g2_fill_2 FILLER_55_2423 ();
 sg13g2_fill_2 FILLER_55_2429 ();
 sg13g2_fill_1 FILLER_55_2431 ();
 sg13g2_fill_1 FILLER_55_2442 ();
 sg13g2_fill_2 FILLER_55_2490 ();
 sg13g2_fill_1 FILLER_55_2492 ();
 sg13g2_fill_2 FILLER_55_2499 ();
 sg13g2_fill_1 FILLER_55_2501 ();
 sg13g2_decap_8 FILLER_55_2534 ();
 sg13g2_decap_8 FILLER_55_2545 ();
 sg13g2_decap_8 FILLER_55_2552 ();
 sg13g2_decap_8 FILLER_55_2559 ();
 sg13g2_decap_8 FILLER_55_2566 ();
 sg13g2_decap_4 FILLER_55_2573 ();
 sg13g2_fill_2 FILLER_55_2577 ();
 sg13g2_fill_2 FILLER_55_2619 ();
 sg13g2_fill_1 FILLER_55_2621 ();
 sg13g2_decap_8 FILLER_55_2652 ();
 sg13g2_decap_8 FILLER_55_2659 ();
 sg13g2_decap_4 FILLER_55_2666 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_52 ();
 sg13g2_fill_2 FILLER_56_59 ();
 sg13g2_decap_4 FILLER_56_66 ();
 sg13g2_decap_8 FILLER_56_78 ();
 sg13g2_decap_8 FILLER_56_85 ();
 sg13g2_decap_8 FILLER_56_92 ();
 sg13g2_decap_8 FILLER_56_99 ();
 sg13g2_decap_8 FILLER_56_106 ();
 sg13g2_decap_8 FILLER_56_113 ();
 sg13g2_decap_8 FILLER_56_120 ();
 sg13g2_decap_8 FILLER_56_127 ();
 sg13g2_decap_8 FILLER_56_134 ();
 sg13g2_decap_8 FILLER_56_141 ();
 sg13g2_decap_8 FILLER_56_148 ();
 sg13g2_decap_4 FILLER_56_155 ();
 sg13g2_fill_2 FILLER_56_159 ();
 sg13g2_decap_4 FILLER_56_228 ();
 sg13g2_fill_2 FILLER_56_232 ();
 sg13g2_decap_8 FILLER_56_260 ();
 sg13g2_fill_2 FILLER_56_267 ();
 sg13g2_fill_1 FILLER_56_269 ();
 sg13g2_decap_8 FILLER_56_303 ();
 sg13g2_decap_4 FILLER_56_310 ();
 sg13g2_fill_2 FILLER_56_314 ();
 sg13g2_decap_8 FILLER_56_324 ();
 sg13g2_decap_8 FILLER_56_331 ();
 sg13g2_fill_2 FILLER_56_338 ();
 sg13g2_fill_1 FILLER_56_354 ();
 sg13g2_decap_4 FILLER_56_372 ();
 sg13g2_fill_2 FILLER_56_376 ();
 sg13g2_fill_1 FILLER_56_392 ();
 sg13g2_fill_2 FILLER_56_398 ();
 sg13g2_fill_1 FILLER_56_405 ();
 sg13g2_fill_2 FILLER_56_410 ();
 sg13g2_fill_2 FILLER_56_416 ();
 sg13g2_fill_1 FILLER_56_418 ();
 sg13g2_fill_2 FILLER_56_423 ();
 sg13g2_fill_1 FILLER_56_425 ();
 sg13g2_fill_2 FILLER_56_430 ();
 sg13g2_decap_8 FILLER_56_455 ();
 sg13g2_fill_1 FILLER_56_462 ();
 sg13g2_decap_4 FILLER_56_468 ();
 sg13g2_fill_1 FILLER_56_472 ();
 sg13g2_decap_4 FILLER_56_481 ();
 sg13g2_fill_1 FILLER_56_485 ();
 sg13g2_fill_1 FILLER_56_491 ();
 sg13g2_fill_1 FILLER_56_500 ();
 sg13g2_fill_1 FILLER_56_519 ();
 sg13g2_fill_2 FILLER_56_529 ();
 sg13g2_fill_1 FILLER_56_542 ();
 sg13g2_fill_1 FILLER_56_548 ();
 sg13g2_decap_4 FILLER_56_557 ();
 sg13g2_fill_1 FILLER_56_571 ();
 sg13g2_decap_4 FILLER_56_578 ();
 sg13g2_fill_2 FILLER_56_582 ();
 sg13g2_decap_8 FILLER_56_594 ();
 sg13g2_decap_4 FILLER_56_601 ();
 sg13g2_fill_2 FILLER_56_605 ();
 sg13g2_fill_2 FILLER_56_611 ();
 sg13g2_decap_4 FILLER_56_623 ();
 sg13g2_fill_1 FILLER_56_627 ();
 sg13g2_fill_2 FILLER_56_643 ();
 sg13g2_fill_2 FILLER_56_650 ();
 sg13g2_decap_4 FILLER_56_670 ();
 sg13g2_decap_8 FILLER_56_696 ();
 sg13g2_decap_4 FILLER_56_703 ();
 sg13g2_fill_1 FILLER_56_707 ();
 sg13g2_fill_1 FILLER_56_716 ();
 sg13g2_decap_8 FILLER_56_761 ();
 sg13g2_decap_8 FILLER_56_768 ();
 sg13g2_decap_4 FILLER_56_775 ();
 sg13g2_fill_2 FILLER_56_795 ();
 sg13g2_fill_1 FILLER_56_803 ();
 sg13g2_decap_8 FILLER_56_820 ();
 sg13g2_decap_8 FILLER_56_827 ();
 sg13g2_decap_8 FILLER_56_834 ();
 sg13g2_fill_2 FILLER_56_841 ();
 sg13g2_fill_1 FILLER_56_843 ();
 sg13g2_decap_8 FILLER_56_852 ();
 sg13g2_fill_2 FILLER_56_859 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_decap_4 FILLER_56_872 ();
 sg13g2_fill_2 FILLER_56_880 ();
 sg13g2_fill_1 FILLER_56_882 ();
 sg13g2_fill_2 FILLER_56_945 ();
 sg13g2_decap_8 FILLER_56_951 ();
 sg13g2_decap_8 FILLER_56_958 ();
 sg13g2_decap_8 FILLER_56_965 ();
 sg13g2_decap_4 FILLER_56_977 ();
 sg13g2_fill_2 FILLER_56_1002 ();
 sg13g2_fill_1 FILLER_56_1030 ();
 sg13g2_fill_1 FILLER_56_1039 ();
 sg13g2_fill_2 FILLER_56_1046 ();
 sg13g2_fill_1 FILLER_56_1056 ();
 sg13g2_fill_1 FILLER_56_1061 ();
 sg13g2_fill_2 FILLER_56_1088 ();
 sg13g2_decap_8 FILLER_56_1102 ();
 sg13g2_decap_8 FILLER_56_1139 ();
 sg13g2_fill_1 FILLER_56_1146 ();
 sg13g2_decap_8 FILLER_56_1151 ();
 sg13g2_fill_2 FILLER_56_1158 ();
 sg13g2_fill_1 FILLER_56_1160 ();
 sg13g2_decap_8 FILLER_56_1166 ();
 sg13g2_decap_8 FILLER_56_1173 ();
 sg13g2_fill_2 FILLER_56_1180 ();
 sg13g2_decap_8 FILLER_56_1190 ();
 sg13g2_decap_8 FILLER_56_1197 ();
 sg13g2_decap_8 FILLER_56_1204 ();
 sg13g2_decap_4 FILLER_56_1215 ();
 sg13g2_decap_8 FILLER_56_1252 ();
 sg13g2_decap_8 FILLER_56_1259 ();
 sg13g2_decap_8 FILLER_56_1266 ();
 sg13g2_fill_1 FILLER_56_1273 ();
 sg13g2_fill_1 FILLER_56_1278 ();
 sg13g2_fill_1 FILLER_56_1290 ();
 sg13g2_decap_4 FILLER_56_1295 ();
 sg13g2_decap_4 FILLER_56_1308 ();
 sg13g2_fill_2 FILLER_56_1312 ();
 sg13g2_decap_8 FILLER_56_1327 ();
 sg13g2_fill_2 FILLER_56_1334 ();
 sg13g2_fill_2 FILLER_56_1340 ();
 sg13g2_fill_2 FILLER_56_1368 ();
 sg13g2_fill_1 FILLER_56_1391 ();
 sg13g2_decap_8 FILLER_56_1424 ();
 sg13g2_decap_4 FILLER_56_1431 ();
 sg13g2_decap_4 FILLER_56_1441 ();
 sg13g2_fill_2 FILLER_56_1445 ();
 sg13g2_fill_1 FILLER_56_1452 ();
 sg13g2_fill_2 FILLER_56_1459 ();
 sg13g2_decap_8 FILLER_56_1464 ();
 sg13g2_fill_1 FILLER_56_1471 ();
 sg13g2_decap_8 FILLER_56_1502 ();
 sg13g2_decap_8 FILLER_56_1509 ();
 sg13g2_decap_8 FILLER_56_1516 ();
 sg13g2_decap_4 FILLER_56_1523 ();
 sg13g2_fill_2 FILLER_56_1532 ();
 sg13g2_decap_4 FILLER_56_1563 ();
 sg13g2_fill_1 FILLER_56_1579 ();
 sg13g2_decap_4 FILLER_56_1593 ();
 sg13g2_fill_1 FILLER_56_1597 ();
 sg13g2_fill_2 FILLER_56_1606 ();
 sg13g2_fill_1 FILLER_56_1608 ();
 sg13g2_fill_1 FILLER_56_1661 ();
 sg13g2_decap_8 FILLER_56_1715 ();
 sg13g2_decap_8 FILLER_56_1722 ();
 sg13g2_decap_8 FILLER_56_1729 ();
 sg13g2_decap_4 FILLER_56_1736 ();
 sg13g2_fill_2 FILLER_56_1740 ();
 sg13g2_decap_8 FILLER_56_1747 ();
 sg13g2_decap_4 FILLER_56_1758 ();
 sg13g2_fill_1 FILLER_56_1762 ();
 sg13g2_decap_8 FILLER_56_1793 ();
 sg13g2_fill_2 FILLER_56_1800 ();
 sg13g2_fill_1 FILLER_56_1802 ();
 sg13g2_fill_2 FILLER_56_1824 ();
 sg13g2_fill_1 FILLER_56_1826 ();
 sg13g2_decap_4 FILLER_56_1834 ();
 sg13g2_fill_2 FILLER_56_1838 ();
 sg13g2_decap_4 FILLER_56_1844 ();
 sg13g2_fill_2 FILLER_56_1848 ();
 sg13g2_decap_8 FILLER_56_1863 ();
 sg13g2_decap_8 FILLER_56_1870 ();
 sg13g2_fill_2 FILLER_56_1877 ();
 sg13g2_fill_1 FILLER_56_1879 ();
 sg13g2_fill_2 FILLER_56_1884 ();
 sg13g2_fill_1 FILLER_56_1890 ();
 sg13g2_decap_4 FILLER_56_1896 ();
 sg13g2_fill_1 FILLER_56_1900 ();
 sg13g2_decap_8 FILLER_56_1905 ();
 sg13g2_fill_1 FILLER_56_1912 ();
 sg13g2_decap_8 FILLER_56_1922 ();
 sg13g2_fill_2 FILLER_56_1929 ();
 sg13g2_fill_1 FILLER_56_1931 ();
 sg13g2_fill_2 FILLER_56_1941 ();
 sg13g2_fill_2 FILLER_56_1948 ();
 sg13g2_fill_1 FILLER_56_1950 ();
 sg13g2_fill_1 FILLER_56_1956 ();
 sg13g2_decap_8 FILLER_56_1961 ();
 sg13g2_decap_4 FILLER_56_1968 ();
 sg13g2_fill_1 FILLER_56_1977 ();
 sg13g2_fill_1 FILLER_56_1988 ();
 sg13g2_decap_4 FILLER_56_2052 ();
 sg13g2_fill_2 FILLER_56_2056 ();
 sg13g2_fill_2 FILLER_56_2073 ();
 sg13g2_fill_1 FILLER_56_2075 ();
 sg13g2_decap_8 FILLER_56_2106 ();
 sg13g2_decap_8 FILLER_56_2113 ();
 sg13g2_fill_2 FILLER_56_2120 ();
 sg13g2_decap_8 FILLER_56_2126 ();
 sg13g2_fill_2 FILLER_56_2133 ();
 sg13g2_decap_4 FILLER_56_2139 ();
 sg13g2_fill_2 FILLER_56_2143 ();
 sg13g2_decap_4 FILLER_56_2162 ();
 sg13g2_fill_2 FILLER_56_2187 ();
 sg13g2_fill_1 FILLER_56_2189 ();
 sg13g2_fill_2 FILLER_56_2196 ();
 sg13g2_fill_1 FILLER_56_2198 ();
 sg13g2_fill_2 FILLER_56_2225 ();
 sg13g2_decap_4 FILLER_56_2245 ();
 sg13g2_decap_8 FILLER_56_2253 ();
 sg13g2_decap_8 FILLER_56_2260 ();
 sg13g2_decap_8 FILLER_56_2267 ();
 sg13g2_fill_1 FILLER_56_2274 ();
 sg13g2_decap_8 FILLER_56_2279 ();
 sg13g2_fill_1 FILLER_56_2286 ();
 sg13g2_decap_8 FILLER_56_2291 ();
 sg13g2_fill_1 FILLER_56_2298 ();
 sg13g2_fill_1 FILLER_56_2336 ();
 sg13g2_fill_1 FILLER_56_2342 ();
 sg13g2_fill_2 FILLER_56_2353 ();
 sg13g2_decap_8 FILLER_56_2406 ();
 sg13g2_decap_4 FILLER_56_2413 ();
 sg13g2_decap_8 FILLER_56_2422 ();
 sg13g2_decap_8 FILLER_56_2429 ();
 sg13g2_fill_1 FILLER_56_2436 ();
 sg13g2_fill_2 FILLER_56_2441 ();
 sg13g2_fill_1 FILLER_56_2448 ();
 sg13g2_fill_1 FILLER_56_2477 ();
 sg13g2_decap_8 FILLER_56_2507 ();
 sg13g2_fill_2 FILLER_56_2514 ();
 sg13g2_fill_2 FILLER_56_2528 ();
 sg13g2_fill_2 FILLER_56_2539 ();
 sg13g2_fill_1 FILLER_56_2541 ();
 sg13g2_fill_1 FILLER_56_2573 ();
 sg13g2_fill_2 FILLER_56_2587 ();
 sg13g2_decap_8 FILLER_56_2615 ();
 sg13g2_decap_8 FILLER_56_2622 ();
 sg13g2_fill_1 FILLER_56_2629 ();
 sg13g2_fill_1 FILLER_56_2638 ();
 sg13g2_decap_8 FILLER_56_2643 ();
 sg13g2_decap_8 FILLER_56_2650 ();
 sg13g2_decap_8 FILLER_56_2657 ();
 sg13g2_decap_4 FILLER_56_2664 ();
 sg13g2_fill_2 FILLER_56_2668 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_4 ();
 sg13g2_fill_2 FILLER_57_31 ();
 sg13g2_decap_4 FILLER_57_38 ();
 sg13g2_decap_8 FILLER_57_68 ();
 sg13g2_decap_8 FILLER_57_75 ();
 sg13g2_decap_8 FILLER_57_82 ();
 sg13g2_decap_8 FILLER_57_89 ();
 sg13g2_decap_8 FILLER_57_96 ();
 sg13g2_decap_8 FILLER_57_103 ();
 sg13g2_decap_8 FILLER_57_110 ();
 sg13g2_decap_8 FILLER_57_117 ();
 sg13g2_decap_8 FILLER_57_124 ();
 sg13g2_decap_8 FILLER_57_131 ();
 sg13g2_decap_8 FILLER_57_138 ();
 sg13g2_decap_8 FILLER_57_145 ();
 sg13g2_decap_8 FILLER_57_152 ();
 sg13g2_decap_8 FILLER_57_159 ();
 sg13g2_decap_8 FILLER_57_166 ();
 sg13g2_decap_8 FILLER_57_173 ();
 sg13g2_decap_8 FILLER_57_180 ();
 sg13g2_decap_8 FILLER_57_187 ();
 sg13g2_decap_8 FILLER_57_194 ();
 sg13g2_decap_8 FILLER_57_201 ();
 sg13g2_fill_1 FILLER_57_208 ();
 sg13g2_decap_8 FILLER_57_243 ();
 sg13g2_decap_8 FILLER_57_250 ();
 sg13g2_decap_8 FILLER_57_257 ();
 sg13g2_fill_2 FILLER_57_264 ();
 sg13g2_fill_1 FILLER_57_266 ();
 sg13g2_decap_4 FILLER_57_304 ();
 sg13g2_fill_1 FILLER_57_308 ();
 sg13g2_fill_2 FILLER_57_313 ();
 sg13g2_fill_1 FILLER_57_315 ();
 sg13g2_fill_2 FILLER_57_337 ();
 sg13g2_decap_8 FILLER_57_349 ();
 sg13g2_decap_8 FILLER_57_356 ();
 sg13g2_fill_2 FILLER_57_363 ();
 sg13g2_fill_1 FILLER_57_436 ();
 sg13g2_fill_1 FILLER_57_447 ();
 sg13g2_fill_2 FILLER_57_474 ();
 sg13g2_fill_2 FILLER_57_481 ();
 sg13g2_decap_8 FILLER_57_490 ();
 sg13g2_decap_8 FILLER_57_497 ();
 sg13g2_fill_1 FILLER_57_532 ();
 sg13g2_fill_2 FILLER_57_538 ();
 sg13g2_fill_1 FILLER_57_540 ();
 sg13g2_fill_2 FILLER_57_545 ();
 sg13g2_decap_8 FILLER_57_552 ();
 sg13g2_decap_4 FILLER_57_559 ();
 sg13g2_fill_2 FILLER_57_589 ();
 sg13g2_fill_1 FILLER_57_591 ();
 sg13g2_fill_1 FILLER_57_597 ();
 sg13g2_fill_2 FILLER_57_602 ();
 sg13g2_fill_1 FILLER_57_604 ();
 sg13g2_decap_4 FILLER_57_629 ();
 sg13g2_decap_4 FILLER_57_641 ();
 sg13g2_fill_1 FILLER_57_645 ();
 sg13g2_decap_8 FILLER_57_677 ();
 sg13g2_fill_2 FILLER_57_684 ();
 sg13g2_fill_2 FILLER_57_690 ();
 sg13g2_fill_1 FILLER_57_697 ();
 sg13g2_fill_2 FILLER_57_715 ();
 sg13g2_fill_1 FILLER_57_722 ();
 sg13g2_fill_1 FILLER_57_727 ();
 sg13g2_fill_2 FILLER_57_759 ();
 sg13g2_fill_1 FILLER_57_761 ();
 sg13g2_decap_8 FILLER_57_780 ();
 sg13g2_decap_8 FILLER_57_787 ();
 sg13g2_fill_2 FILLER_57_794 ();
 sg13g2_fill_1 FILLER_57_799 ();
 sg13g2_decap_8 FILLER_57_809 ();
 sg13g2_fill_2 FILLER_57_816 ();
 sg13g2_fill_1 FILLER_57_818 ();
 sg13g2_decap_8 FILLER_57_822 ();
 sg13g2_fill_2 FILLER_57_829 ();
 sg13g2_decap_8 FILLER_57_870 ();
 sg13g2_decap_8 FILLER_57_877 ();
 sg13g2_fill_2 FILLER_57_884 ();
 sg13g2_fill_1 FILLER_57_886 ();
 sg13g2_fill_1 FILLER_57_895 ();
 sg13g2_fill_2 FILLER_57_922 ();
 sg13g2_decap_4 FILLER_57_971 ();
 sg13g2_fill_1 FILLER_57_975 ();
 sg13g2_fill_2 FILLER_57_995 ();
 sg13g2_fill_1 FILLER_57_1009 ();
 sg13g2_decap_8 FILLER_57_1015 ();
 sg13g2_decap_8 FILLER_57_1022 ();
 sg13g2_decap_8 FILLER_57_1029 ();
 sg13g2_fill_2 FILLER_57_1036 ();
 sg13g2_decap_8 FILLER_57_1043 ();
 sg13g2_fill_2 FILLER_57_1050 ();
 sg13g2_decap_8 FILLER_57_1056 ();
 sg13g2_fill_1 FILLER_57_1067 ();
 sg13g2_fill_2 FILLER_57_1072 ();
 sg13g2_fill_1 FILLER_57_1079 ();
 sg13g2_fill_2 FILLER_57_1084 ();
 sg13g2_fill_2 FILLER_57_1092 ();
 sg13g2_fill_1 FILLER_57_1094 ();
 sg13g2_decap_8 FILLER_57_1132 ();
 sg13g2_fill_2 FILLER_57_1139 ();
 sg13g2_fill_1 FILLER_57_1141 ();
 sg13g2_decap_8 FILLER_57_1146 ();
 sg13g2_decap_8 FILLER_57_1153 ();
 sg13g2_decap_4 FILLER_57_1191 ();
 sg13g2_fill_2 FILLER_57_1207 ();
 sg13g2_fill_1 FILLER_57_1235 ();
 sg13g2_decap_4 FILLER_57_1250 ();
 sg13g2_fill_1 FILLER_57_1284 ();
 sg13g2_decap_8 FILLER_57_1315 ();
 sg13g2_fill_1 FILLER_57_1322 ();
 sg13g2_fill_2 FILLER_57_1327 ();
 sg13g2_fill_2 FILLER_57_1355 ();
 sg13g2_fill_1 FILLER_57_1407 ();
 sg13g2_decap_8 FILLER_57_1446 ();
 sg13g2_decap_4 FILLER_57_1453 ();
 sg13g2_fill_2 FILLER_57_1457 ();
 sg13g2_decap_8 FILLER_57_1464 ();
 sg13g2_decap_4 FILLER_57_1471 ();
 sg13g2_decap_4 FILLER_57_1479 ();
 sg13g2_decap_4 FILLER_57_1487 ();
 sg13g2_decap_8 FILLER_57_1506 ();
 sg13g2_decap_8 FILLER_57_1513 ();
 sg13g2_fill_1 FILLER_57_1520 ();
 sg13g2_decap_4 FILLER_57_1535 ();
 sg13g2_decap_8 FILLER_57_1543 ();
 sg13g2_decap_8 FILLER_57_1550 ();
 sg13g2_fill_1 FILLER_57_1557 ();
 sg13g2_fill_2 FILLER_57_1592 ();
 sg13g2_fill_1 FILLER_57_1594 ();
 sg13g2_fill_1 FILLER_57_1605 ();
 sg13g2_fill_2 FILLER_57_1611 ();
 sg13g2_decap_4 FILLER_57_1689 ();
 sg13g2_fill_2 FILLER_57_1693 ();
 sg13g2_fill_2 FILLER_57_1721 ();
 sg13g2_fill_1 FILLER_57_1723 ();
 sg13g2_decap_4 FILLER_57_1728 ();
 sg13g2_fill_1 FILLER_57_1732 ();
 sg13g2_fill_2 FILLER_57_1738 ();
 sg13g2_decap_8 FILLER_57_1766 ();
 sg13g2_decap_4 FILLER_57_1777 ();
 sg13g2_fill_2 FILLER_57_1781 ();
 sg13g2_fill_1 FILLER_57_1791 ();
 sg13g2_fill_1 FILLER_57_1823 ();
 sg13g2_decap_8 FILLER_57_1828 ();
 sg13g2_fill_2 FILLER_57_1835 ();
 sg13g2_fill_1 FILLER_57_1837 ();
 sg13g2_fill_1 FILLER_57_1859 ();
 sg13g2_decap_4 FILLER_57_1891 ();
 sg13g2_fill_2 FILLER_57_1895 ();
 sg13g2_decap_8 FILLER_57_1901 ();
 sg13g2_decap_8 FILLER_57_1908 ();
 sg13g2_decap_8 FILLER_57_1915 ();
 sg13g2_decap_4 FILLER_57_1922 ();
 sg13g2_fill_1 FILLER_57_1926 ();
 sg13g2_fill_1 FILLER_57_1997 ();
 sg13g2_fill_2 FILLER_57_2030 ();
 sg13g2_decap_4 FILLER_57_2042 ();
 sg13g2_fill_2 FILLER_57_2046 ();
 sg13g2_decap_4 FILLER_57_2052 ();
 sg13g2_fill_2 FILLER_57_2061 ();
 sg13g2_fill_2 FILLER_57_2067 ();
 sg13g2_decap_4 FILLER_57_2074 ();
 sg13g2_decap_4 FILLER_57_2086 ();
 sg13g2_fill_2 FILLER_57_2099 ();
 sg13g2_fill_1 FILLER_57_2101 ();
 sg13g2_decap_4 FILLER_57_2107 ();
 sg13g2_decap_8 FILLER_57_2137 ();
 sg13g2_decap_8 FILLER_57_2144 ();
 sg13g2_fill_2 FILLER_57_2151 ();
 sg13g2_fill_1 FILLER_57_2210 ();
 sg13g2_decap_4 FILLER_57_2215 ();
 sg13g2_fill_1 FILLER_57_2219 ();
 sg13g2_fill_2 FILLER_57_2238 ();
 sg13g2_fill_1 FILLER_57_2272 ();
 sg13g2_decap_8 FILLER_57_2277 ();
 sg13g2_decap_4 FILLER_57_2284 ();
 sg13g2_fill_2 FILLER_57_2288 ();
 sg13g2_decap_8 FILLER_57_2295 ();
 sg13g2_fill_2 FILLER_57_2302 ();
 sg13g2_fill_1 FILLER_57_2334 ();
 sg13g2_fill_1 FILLER_57_2340 ();
 sg13g2_fill_1 FILLER_57_2345 ();
 sg13g2_decap_4 FILLER_57_2351 ();
 sg13g2_decap_8 FILLER_57_2364 ();
 sg13g2_decap_8 FILLER_57_2371 ();
 sg13g2_fill_1 FILLER_57_2378 ();
 sg13g2_decap_8 FILLER_57_2384 ();
 sg13g2_fill_1 FILLER_57_2391 ();
 sg13g2_decap_4 FILLER_57_2422 ();
 sg13g2_fill_1 FILLER_57_2426 ();
 sg13g2_decap_4 FILLER_57_2431 ();
 sg13g2_fill_2 FILLER_57_2444 ();
 sg13g2_fill_2 FILLER_57_2450 ();
 sg13g2_fill_1 FILLER_57_2452 ();
 sg13g2_fill_2 FILLER_57_2461 ();
 sg13g2_fill_1 FILLER_57_2477 ();
 sg13g2_decap_8 FILLER_57_2499 ();
 sg13g2_decap_8 FILLER_57_2506 ();
 sg13g2_fill_1 FILLER_57_2513 ();
 sg13g2_decap_4 FILLER_57_2523 ();
 sg13g2_fill_2 FILLER_57_2571 ();
 sg13g2_fill_2 FILLER_57_2578 ();
 sg13g2_fill_2 FILLER_57_2584 ();
 sg13g2_fill_1 FILLER_57_2586 ();
 sg13g2_decap_8 FILLER_57_2592 ();
 sg13g2_decap_8 FILLER_57_2599 ();
 sg13g2_decap_8 FILLER_57_2606 ();
 sg13g2_decap_8 FILLER_57_2613 ();
 sg13g2_decap_8 FILLER_57_2620 ();
 sg13g2_decap_8 FILLER_57_2627 ();
 sg13g2_decap_8 FILLER_57_2634 ();
 sg13g2_decap_8 FILLER_57_2641 ();
 sg13g2_decap_8 FILLER_57_2648 ();
 sg13g2_decap_8 FILLER_57_2655 ();
 sg13g2_decap_8 FILLER_57_2662 ();
 sg13g2_fill_1 FILLER_57_2669 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_fill_2 FILLER_58_91 ();
 sg13g2_fill_1 FILLER_58_93 ();
 sg13g2_decap_8 FILLER_58_103 ();
 sg13g2_decap_8 FILLER_58_110 ();
 sg13g2_decap_8 FILLER_58_117 ();
 sg13g2_decap_8 FILLER_58_124 ();
 sg13g2_decap_8 FILLER_58_131 ();
 sg13g2_decap_8 FILLER_58_138 ();
 sg13g2_decap_8 FILLER_58_145 ();
 sg13g2_decap_8 FILLER_58_152 ();
 sg13g2_decap_8 FILLER_58_159 ();
 sg13g2_decap_8 FILLER_58_166 ();
 sg13g2_decap_8 FILLER_58_173 ();
 sg13g2_decap_8 FILLER_58_180 ();
 sg13g2_decap_8 FILLER_58_187 ();
 sg13g2_decap_8 FILLER_58_194 ();
 sg13g2_decap_8 FILLER_58_201 ();
 sg13g2_decap_8 FILLER_58_208 ();
 sg13g2_decap_4 FILLER_58_215 ();
 sg13g2_fill_2 FILLER_58_219 ();
 sg13g2_decap_4 FILLER_58_231 ();
 sg13g2_fill_1 FILLER_58_235 ();
 sg13g2_fill_2 FILLER_58_296 ();
 sg13g2_fill_2 FILLER_58_307 ();
 sg13g2_decap_8 FILLER_58_339 ();
 sg13g2_decap_8 FILLER_58_346 ();
 sg13g2_decap_8 FILLER_58_353 ();
 sg13g2_decap_8 FILLER_58_360 ();
 sg13g2_fill_1 FILLER_58_367 ();
 sg13g2_fill_2 FILLER_58_381 ();
 sg13g2_fill_2 FILLER_58_388 ();
 sg13g2_fill_1 FILLER_58_418 ();
 sg13g2_fill_1 FILLER_58_424 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_fill_1 FILLER_58_434 ();
 sg13g2_fill_2 FILLER_58_461 ();
 sg13g2_fill_2 FILLER_58_472 ();
 sg13g2_fill_2 FILLER_58_479 ();
 sg13g2_fill_1 FILLER_58_481 ();
 sg13g2_fill_1 FILLER_58_486 ();
 sg13g2_decap_4 FILLER_58_495 ();
 sg13g2_fill_1 FILLER_58_499 ();
 sg13g2_fill_1 FILLER_58_504 ();
 sg13g2_fill_1 FILLER_58_509 ();
 sg13g2_fill_2 FILLER_58_515 ();
 sg13g2_decap_8 FILLER_58_531 ();
 sg13g2_decap_8 FILLER_58_538 ();
 sg13g2_decap_8 FILLER_58_545 ();
 sg13g2_decap_8 FILLER_58_552 ();
 sg13g2_fill_2 FILLER_58_559 ();
 sg13g2_fill_1 FILLER_58_561 ();
 sg13g2_decap_4 FILLER_58_576 ();
 sg13g2_decap_4 FILLER_58_588 ();
 sg13g2_decap_8 FILLER_58_602 ();
 sg13g2_decap_8 FILLER_58_609 ();
 sg13g2_fill_2 FILLER_58_620 ();
 sg13g2_fill_1 FILLER_58_622 ();
 sg13g2_decap_4 FILLER_58_641 ();
 sg13g2_fill_2 FILLER_58_659 ();
 sg13g2_fill_1 FILLER_58_666 ();
 sg13g2_fill_1 FILLER_58_672 ();
 sg13g2_fill_2 FILLER_58_677 ();
 sg13g2_fill_1 FILLER_58_679 ();
 sg13g2_decap_4 FILLER_58_685 ();
 sg13g2_fill_2 FILLER_58_697 ();
 sg13g2_fill_2 FILLER_58_732 ();
 sg13g2_fill_1 FILLER_58_756 ();
 sg13g2_fill_1 FILLER_58_794 ();
 sg13g2_decap_8 FILLER_58_832 ();
 sg13g2_decap_8 FILLER_58_839 ();
 sg13g2_decap_8 FILLER_58_846 ();
 sg13g2_decap_8 FILLER_58_901 ();
 sg13g2_decap_8 FILLER_58_908 ();
 sg13g2_decap_8 FILLER_58_915 ();
 sg13g2_decap_8 FILLER_58_922 ();
 sg13g2_decap_8 FILLER_58_929 ();
 sg13g2_decap_8 FILLER_58_936 ();
 sg13g2_fill_2 FILLER_58_943 ();
 sg13g2_decap_4 FILLER_58_975 ();
 sg13g2_fill_1 FILLER_58_979 ();
 sg13g2_fill_1 FILLER_58_1028 ();
 sg13g2_decap_8 FILLER_58_1048 ();
 sg13g2_fill_2 FILLER_58_1059 ();
 sg13g2_fill_2 FILLER_58_1065 ();
 sg13g2_fill_1 FILLER_58_1067 ();
 sg13g2_fill_2 FILLER_58_1073 ();
 sg13g2_fill_1 FILLER_58_1075 ();
 sg13g2_fill_2 FILLER_58_1102 ();
 sg13g2_fill_1 FILLER_58_1121 ();
 sg13g2_decap_8 FILLER_58_1130 ();
 sg13g2_fill_1 FILLER_58_1137 ();
 sg13g2_fill_2 FILLER_58_1160 ();
 sg13g2_fill_1 FILLER_58_1162 ();
 sg13g2_fill_2 FILLER_58_1172 ();
 sg13g2_fill_1 FILLER_58_1200 ();
 sg13g2_fill_2 FILLER_58_1206 ();
 sg13g2_fill_2 FILLER_58_1228 ();
 sg13g2_fill_1 FILLER_58_1245 ();
 sg13g2_fill_2 FILLER_58_1292 ();
 sg13g2_decap_8 FILLER_58_1298 ();
 sg13g2_fill_2 FILLER_58_1305 ();
 sg13g2_fill_1 FILLER_58_1307 ();
 sg13g2_fill_2 FILLER_58_1363 ();
 sg13g2_fill_1 FILLER_58_1365 ();
 sg13g2_fill_1 FILLER_58_1401 ();
 sg13g2_decap_8 FILLER_58_1418 ();
 sg13g2_decap_8 FILLER_58_1425 ();
 sg13g2_decap_8 FILLER_58_1432 ();
 sg13g2_decap_8 FILLER_58_1439 ();
 sg13g2_fill_2 FILLER_58_1446 ();
 sg13g2_decap_8 FILLER_58_1451 ();
 sg13g2_decap_4 FILLER_58_1458 ();
 sg13g2_fill_2 FILLER_58_1467 ();
 sg13g2_fill_1 FILLER_58_1500 ();
 sg13g2_fill_1 FILLER_58_1534 ();
 sg13g2_decap_8 FILLER_58_1570 ();
 sg13g2_fill_2 FILLER_58_1577 ();
 sg13g2_fill_1 FILLER_58_1579 ();
 sg13g2_decap_8 FILLER_58_1586 ();
 sg13g2_decap_4 FILLER_58_1593 ();
 sg13g2_fill_1 FILLER_58_1597 ();
 sg13g2_decap_8 FILLER_58_1601 ();
 sg13g2_fill_1 FILLER_58_1626 ();
 sg13g2_fill_1 FILLER_58_1636 ();
 sg13g2_fill_1 FILLER_58_1650 ();
 sg13g2_fill_1 FILLER_58_1654 ();
 sg13g2_fill_1 FILLER_58_1666 ();
 sg13g2_fill_2 FILLER_58_1675 ();
 sg13g2_fill_2 FILLER_58_1703 ();
 sg13g2_fill_1 FILLER_58_1705 ();
 sg13g2_fill_2 FILLER_58_1725 ();
 sg13g2_fill_1 FILLER_58_1727 ();
 sg13g2_decap_4 FILLER_58_1747 ();
 sg13g2_fill_1 FILLER_58_1751 ();
 sg13g2_decap_8 FILLER_58_1761 ();
 sg13g2_decap_8 FILLER_58_1772 ();
 sg13g2_decap_4 FILLER_58_1779 ();
 sg13g2_fill_2 FILLER_58_1783 ();
 sg13g2_fill_2 FILLER_58_1793 ();
 sg13g2_fill_2 FILLER_58_1806 ();
 sg13g2_fill_2 FILLER_58_1813 ();
 sg13g2_fill_1 FILLER_58_1815 ();
 sg13g2_decap_8 FILLER_58_1821 ();
 sg13g2_fill_2 FILLER_58_1828 ();
 sg13g2_fill_2 FILLER_58_1853 ();
 sg13g2_fill_1 FILLER_58_1855 ();
 sg13g2_fill_2 FILLER_58_1865 ();
 sg13g2_fill_1 FILLER_58_1867 ();
 sg13g2_fill_2 FILLER_58_1886 ();
 sg13g2_fill_1 FILLER_58_1900 ();
 sg13g2_fill_2 FILLER_58_1976 ();
 sg13g2_fill_1 FILLER_58_1983 ();
 sg13g2_fill_1 FILLER_58_1994 ();
 sg13g2_fill_1 FILLER_58_2051 ();
 sg13g2_decap_8 FILLER_58_2084 ();
 sg13g2_fill_1 FILLER_58_2121 ();
 sg13g2_decap_8 FILLER_58_2149 ();
 sg13g2_decap_8 FILLER_58_2156 ();
 sg13g2_fill_1 FILLER_58_2163 ();
 sg13g2_decap_8 FILLER_58_2168 ();
 sg13g2_decap_4 FILLER_58_2175 ();
 sg13g2_decap_8 FILLER_58_2194 ();
 sg13g2_decap_8 FILLER_58_2201 ();
 sg13g2_fill_2 FILLER_58_2208 ();
 sg13g2_fill_1 FILLER_58_2210 ();
 sg13g2_decap_8 FILLER_58_2292 ();
 sg13g2_decap_8 FILLER_58_2299 ();
 sg13g2_decap_8 FILLER_58_2306 ();
 sg13g2_decap_8 FILLER_58_2313 ();
 sg13g2_fill_2 FILLER_58_2320 ();
 sg13g2_fill_1 FILLER_58_2322 ();
 sg13g2_decap_8 FILLER_58_2349 ();
 sg13g2_decap_8 FILLER_58_2356 ();
 sg13g2_decap_8 FILLER_58_2363 ();
 sg13g2_decap_8 FILLER_58_2370 ();
 sg13g2_decap_8 FILLER_58_2377 ();
 sg13g2_fill_1 FILLER_58_2431 ();
 sg13g2_fill_1 FILLER_58_2436 ();
 sg13g2_fill_1 FILLER_58_2510 ();
 sg13g2_fill_2 FILLER_58_2516 ();
 sg13g2_fill_1 FILLER_58_2531 ();
 sg13g2_fill_1 FILLER_58_2537 ();
 sg13g2_decap_8 FILLER_58_2567 ();
 sg13g2_fill_2 FILLER_58_2574 ();
 sg13g2_fill_2 FILLER_58_2602 ();
 sg13g2_fill_1 FILLER_58_2604 ();
 sg13g2_decap_8 FILLER_58_2635 ();
 sg13g2_decap_8 FILLER_58_2642 ();
 sg13g2_decap_8 FILLER_58_2649 ();
 sg13g2_decap_8 FILLER_58_2656 ();
 sg13g2_decap_8 FILLER_58_2663 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_fill_1 FILLER_59_35 ();
 sg13g2_decap_4 FILLER_59_48 ();
 sg13g2_fill_2 FILLER_59_52 ();
 sg13g2_fill_2 FILLER_59_75 ();
 sg13g2_decap_4 FILLER_59_82 ();
 sg13g2_fill_1 FILLER_59_86 ();
 sg13g2_fill_1 FILLER_59_91 ();
 sg13g2_fill_1 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_131 ();
 sg13g2_fill_1 FILLER_59_138 ();
 sg13g2_fill_2 FILLER_59_143 ();
 sg13g2_fill_1 FILLER_59_145 ();
 sg13g2_fill_1 FILLER_59_155 ();
 sg13g2_fill_2 FILLER_59_164 ();
 sg13g2_fill_1 FILLER_59_166 ();
 sg13g2_decap_4 FILLER_59_177 ();
 sg13g2_fill_2 FILLER_59_185 ();
 sg13g2_decap_8 FILLER_59_191 ();
 sg13g2_decap_8 FILLER_59_198 ();
 sg13g2_decap_8 FILLER_59_205 ();
 sg13g2_decap_8 FILLER_59_212 ();
 sg13g2_decap_8 FILLER_59_219 ();
 sg13g2_decap_4 FILLER_59_226 ();
 sg13g2_fill_2 FILLER_59_230 ();
 sg13g2_decap_8 FILLER_59_245 ();
 sg13g2_decap_8 FILLER_59_252 ();
 sg13g2_decap_8 FILLER_59_259 ();
 sg13g2_decap_8 FILLER_59_266 ();
 sg13g2_fill_1 FILLER_59_273 ();
 sg13g2_decap_8 FILLER_59_381 ();
 sg13g2_decap_8 FILLER_59_388 ();
 sg13g2_decap_8 FILLER_59_395 ();
 sg13g2_decap_4 FILLER_59_402 ();
 sg13g2_decap_8 FILLER_59_410 ();
 sg13g2_decap_4 FILLER_59_417 ();
 sg13g2_fill_2 FILLER_59_421 ();
 sg13g2_fill_2 FILLER_59_479 ();
 sg13g2_fill_1 FILLER_59_481 ();
 sg13g2_decap_8 FILLER_59_487 ();
 sg13g2_decap_8 FILLER_59_494 ();
 sg13g2_decap_8 FILLER_59_501 ();
 sg13g2_decap_8 FILLER_59_508 ();
 sg13g2_fill_2 FILLER_59_515 ();
 sg13g2_decap_8 FILLER_59_521 ();
 sg13g2_decap_8 FILLER_59_528 ();
 sg13g2_decap_8 FILLER_59_535 ();
 sg13g2_decap_8 FILLER_59_542 ();
 sg13g2_fill_1 FILLER_59_549 ();
 sg13g2_decap_8 FILLER_59_560 ();
 sg13g2_decap_4 FILLER_59_567 ();
 sg13g2_fill_2 FILLER_59_571 ();
 sg13g2_decap_8 FILLER_59_582 ();
 sg13g2_decap_4 FILLER_59_589 ();
 sg13g2_fill_2 FILLER_59_593 ();
 sg13g2_fill_2 FILLER_59_621 ();
 sg13g2_decap_4 FILLER_59_630 ();
 sg13g2_fill_2 FILLER_59_634 ();
 sg13g2_decap_4 FILLER_59_641 ();
 sg13g2_fill_1 FILLER_59_645 ();
 sg13g2_fill_2 FILLER_59_651 ();
 sg13g2_fill_2 FILLER_59_658 ();
 sg13g2_decap_8 FILLER_59_664 ();
 sg13g2_decap_8 FILLER_59_675 ();
 sg13g2_fill_1 FILLER_59_682 ();
 sg13g2_fill_2 FILLER_59_700 ();
 sg13g2_fill_1 FILLER_59_706 ();
 sg13g2_fill_1 FILLER_59_712 ();
 sg13g2_fill_1 FILLER_59_721 ();
 sg13g2_fill_2 FILLER_59_758 ();
 sg13g2_fill_1 FILLER_59_764 ();
 sg13g2_decap_8 FILLER_59_773 ();
 sg13g2_decap_8 FILLER_59_780 ();
 sg13g2_fill_1 FILLER_59_814 ();
 sg13g2_fill_1 FILLER_59_832 ();
 sg13g2_fill_2 FILLER_59_846 ();
 sg13g2_fill_1 FILLER_59_848 ();
 sg13g2_decap_4 FILLER_59_853 ();
 sg13g2_fill_1 FILLER_59_857 ();
 sg13g2_fill_2 FILLER_59_870 ();
 sg13g2_decap_8 FILLER_59_926 ();
 sg13g2_decap_8 FILLER_59_933 ();
 sg13g2_fill_1 FILLER_59_940 ();
 sg13g2_decap_4 FILLER_59_989 ();
 sg13g2_fill_2 FILLER_59_993 ();
 sg13g2_fill_2 FILLER_59_1000 ();
 sg13g2_fill_1 FILLER_59_1019 ();
 sg13g2_decap_8 FILLER_59_1046 ();
 sg13g2_decap_4 FILLER_59_1053 ();
 sg13g2_fill_2 FILLER_59_1057 ();
 sg13g2_fill_2 FILLER_59_1065 ();
 sg13g2_fill_1 FILLER_59_1071 ();
 sg13g2_decap_4 FILLER_59_1076 ();
 sg13g2_fill_1 FILLER_59_1080 ();
 sg13g2_decap_4 FILLER_59_1104 ();
 sg13g2_fill_1 FILLER_59_1108 ();
 sg13g2_decap_8 FILLER_59_1169 ();
 sg13g2_fill_2 FILLER_59_1176 ();
 sg13g2_decap_8 FILLER_59_1182 ();
 sg13g2_fill_1 FILLER_59_1189 ();
 sg13g2_fill_2 FILLER_59_1219 ();
 sg13g2_decap_4 FILLER_59_1279 ();
 sg13g2_fill_1 FILLER_59_1283 ();
 sg13g2_decap_4 FILLER_59_1288 ();
 sg13g2_fill_2 FILLER_59_1292 ();
 sg13g2_decap_4 FILLER_59_1339 ();
 sg13g2_decap_4 FILLER_59_1425 ();
 sg13g2_fill_1 FILLER_59_1429 ();
 sg13g2_fill_1 FILLER_59_1443 ();
 sg13g2_fill_2 FILLER_59_1463 ();
 sg13g2_fill_1 FILLER_59_1465 ();
 sg13g2_decap_8 FILLER_59_1477 ();
 sg13g2_decap_8 FILLER_59_1484 ();
 sg13g2_decap_8 FILLER_59_1491 ();
 sg13g2_fill_1 FILLER_59_1498 ();
 sg13g2_fill_2 FILLER_59_1516 ();
 sg13g2_decap_8 FILLER_59_1540 ();
 sg13g2_fill_1 FILLER_59_1547 ();
 sg13g2_fill_1 FILLER_59_1557 ();
 sg13g2_decap_4 FILLER_59_1566 ();
 sg13g2_fill_2 FILLER_59_1570 ();
 sg13g2_fill_2 FILLER_59_1608 ();
 sg13g2_decap_8 FILLER_59_1636 ();
 sg13g2_decap_8 FILLER_59_1643 ();
 sg13g2_fill_1 FILLER_59_1650 ();
 sg13g2_decap_8 FILLER_59_1657 ();
 sg13g2_fill_2 FILLER_59_1664 ();
 sg13g2_fill_1 FILLER_59_1666 ();
 sg13g2_decap_8 FILLER_59_1688 ();
 sg13g2_decap_8 FILLER_59_1695 ();
 sg13g2_fill_2 FILLER_59_1755 ();
 sg13g2_decap_8 FILLER_59_1788 ();
 sg13g2_fill_1 FILLER_59_1809 ();
 sg13g2_decap_8 FILLER_59_1815 ();
 sg13g2_fill_1 FILLER_59_1822 ();
 sg13g2_decap_8 FILLER_59_1827 ();
 sg13g2_decap_8 FILLER_59_1834 ();
 sg13g2_fill_2 FILLER_59_1841 ();
 sg13g2_fill_1 FILLER_59_1843 ();
 sg13g2_fill_1 FILLER_59_1850 ();
 sg13g2_decap_4 FILLER_59_1868 ();
 sg13g2_fill_2 FILLER_59_1872 ();
 sg13g2_fill_2 FILLER_59_1908 ();
 sg13g2_fill_1 FILLER_59_1917 ();
 sg13g2_fill_1 FILLER_59_2000 ();
 sg13g2_decap_8 FILLER_59_2006 ();
 sg13g2_decap_8 FILLER_59_2021 ();
 sg13g2_fill_2 FILLER_59_2028 ();
 sg13g2_fill_1 FILLER_59_2030 ();
 sg13g2_decap_4 FILLER_59_2040 ();
 sg13g2_fill_1 FILLER_59_2044 ();
 sg13g2_fill_2 FILLER_59_2075 ();
 sg13g2_fill_2 FILLER_59_2083 ();
 sg13g2_fill_1 FILLER_59_2090 ();
 sg13g2_fill_1 FILLER_59_2096 ();
 sg13g2_fill_2 FILLER_59_2123 ();
 sg13g2_decap_4 FILLER_59_2161 ();
 sg13g2_fill_1 FILLER_59_2165 ();
 sg13g2_decap_8 FILLER_59_2174 ();
 sg13g2_decap_8 FILLER_59_2181 ();
 sg13g2_fill_1 FILLER_59_2188 ();
 sg13g2_decap_8 FILLER_59_2198 ();
 sg13g2_fill_2 FILLER_59_2205 ();
 sg13g2_fill_1 FILLER_59_2207 ();
 sg13g2_fill_1 FILLER_59_2256 ();
 sg13g2_decap_4 FILLER_59_2261 ();
 sg13g2_fill_1 FILLER_59_2265 ();
 sg13g2_decap_8 FILLER_59_2298 ();
 sg13g2_decap_8 FILLER_59_2305 ();
 sg13g2_decap_8 FILLER_59_2312 ();
 sg13g2_decap_8 FILLER_59_2319 ();
 sg13g2_decap_8 FILLER_59_2326 ();
 sg13g2_decap_8 FILLER_59_2333 ();
 sg13g2_decap_8 FILLER_59_2340 ();
 sg13g2_decap_8 FILLER_59_2347 ();
 sg13g2_decap_8 FILLER_59_2354 ();
 sg13g2_fill_2 FILLER_59_2361 ();
 sg13g2_fill_1 FILLER_59_2363 ();
 sg13g2_decap_8 FILLER_59_2368 ();
 sg13g2_decap_8 FILLER_59_2375 ();
 sg13g2_decap_8 FILLER_59_2382 ();
 sg13g2_fill_2 FILLER_59_2389 ();
 sg13g2_fill_1 FILLER_59_2391 ();
 sg13g2_fill_2 FILLER_59_2402 ();
 sg13g2_decap_8 FILLER_59_2414 ();
 sg13g2_fill_1 FILLER_59_2426 ();
 sg13g2_decap_4 FILLER_59_2453 ();
 sg13g2_fill_2 FILLER_59_2457 ();
 sg13g2_decap_8 FILLER_59_2463 ();
 sg13g2_decap_4 FILLER_59_2470 ();
 sg13g2_decap_4 FILLER_59_2477 ();
 sg13g2_fill_1 FILLER_59_2481 ();
 sg13g2_decap_8 FILLER_59_2488 ();
 sg13g2_decap_8 FILLER_59_2495 ();
 sg13g2_fill_2 FILLER_59_2502 ();
 sg13g2_fill_2 FILLER_59_2512 ();
 sg13g2_decap_8 FILLER_59_2556 ();
 sg13g2_decap_8 FILLER_59_2563 ();
 sg13g2_decap_8 FILLER_59_2570 ();
 sg13g2_decap_8 FILLER_59_2577 ();
 sg13g2_decap_8 FILLER_59_2584 ();
 sg13g2_decap_8 FILLER_59_2591 ();
 sg13g2_decap_8 FILLER_59_2598 ();
 sg13g2_decap_8 FILLER_59_2635 ();
 sg13g2_decap_8 FILLER_59_2642 ();
 sg13g2_decap_8 FILLER_59_2649 ();
 sg13g2_decap_8 FILLER_59_2656 ();
 sg13g2_decap_8 FILLER_59_2663 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_4 FILLER_60_14 ();
 sg13g2_fill_2 FILLER_60_18 ();
 sg13g2_fill_1 FILLER_60_23 ();
 sg13g2_fill_1 FILLER_60_38 ();
 sg13g2_fill_1 FILLER_60_49 ();
 sg13g2_fill_1 FILLER_60_60 ();
 sg13g2_fill_2 FILLER_60_73 ();
 sg13g2_fill_1 FILLER_60_79 ();
 sg13g2_fill_1 FILLER_60_85 ();
 sg13g2_fill_2 FILLER_60_92 ();
 sg13g2_fill_1 FILLER_60_113 ();
 sg13g2_fill_1 FILLER_60_129 ();
 sg13g2_fill_1 FILLER_60_148 ();
 sg13g2_fill_2 FILLER_60_179 ();
 sg13g2_fill_2 FILLER_60_193 ();
 sg13g2_decap_8 FILLER_60_208 ();
 sg13g2_decap_8 FILLER_60_215 ();
 sg13g2_decap_8 FILLER_60_222 ();
 sg13g2_decap_8 FILLER_60_229 ();
 sg13g2_decap_8 FILLER_60_236 ();
 sg13g2_decap_4 FILLER_60_243 ();
 sg13g2_fill_1 FILLER_60_247 ();
 sg13g2_decap_8 FILLER_60_274 ();
 sg13g2_fill_2 FILLER_60_281 ();
 sg13g2_fill_2 FILLER_60_298 ();
 sg13g2_decap_8 FILLER_60_309 ();
 sg13g2_decap_8 FILLER_60_316 ();
 sg13g2_decap_4 FILLER_60_323 ();
 sg13g2_fill_1 FILLER_60_327 ();
 sg13g2_fill_2 FILLER_60_338 ();
 sg13g2_decap_8 FILLER_60_380 ();
 sg13g2_decap_8 FILLER_60_387 ();
 sg13g2_decap_8 FILLER_60_394 ();
 sg13g2_decap_8 FILLER_60_401 ();
 sg13g2_decap_8 FILLER_60_426 ();
 sg13g2_decap_8 FILLER_60_433 ();
 sg13g2_decap_8 FILLER_60_446 ();
 sg13g2_decap_4 FILLER_60_456 ();
 sg13g2_fill_2 FILLER_60_460 ();
 sg13g2_decap_8 FILLER_60_466 ();
 sg13g2_decap_4 FILLER_60_473 ();
 sg13g2_decap_8 FILLER_60_481 ();
 sg13g2_fill_2 FILLER_60_488 ();
 sg13g2_decap_8 FILLER_60_495 ();
 sg13g2_decap_8 FILLER_60_502 ();
 sg13g2_fill_2 FILLER_60_509 ();
 sg13g2_fill_1 FILLER_60_511 ();
 sg13g2_fill_1 FILLER_60_516 ();
 sg13g2_fill_1 FILLER_60_543 ();
 sg13g2_fill_2 FILLER_60_574 ();
 sg13g2_decap_8 FILLER_60_606 ();
 sg13g2_decap_4 FILLER_60_613 ();
 sg13g2_fill_1 FILLER_60_617 ();
 sg13g2_fill_2 FILLER_60_653 ();
 sg13g2_fill_2 FILLER_60_663 ();
 sg13g2_decap_8 FILLER_60_674 ();
 sg13g2_decap_8 FILLER_60_681 ();
 sg13g2_fill_2 FILLER_60_688 ();
 sg13g2_decap_8 FILLER_60_700 ();
 sg13g2_decap_8 FILLER_60_707 ();
 sg13g2_fill_1 FILLER_60_714 ();
 sg13g2_decap_4 FILLER_60_719 ();
 sg13g2_fill_1 FILLER_60_723 ();
 sg13g2_fill_1 FILLER_60_729 ();
 sg13g2_fill_2 FILLER_60_762 ();
 sg13g2_fill_1 FILLER_60_764 ();
 sg13g2_fill_1 FILLER_60_768 ();
 sg13g2_decap_4 FILLER_60_777 ();
 sg13g2_fill_1 FILLER_60_781 ();
 sg13g2_fill_2 FILLER_60_795 ();
 sg13g2_fill_2 FILLER_60_802 ();
 sg13g2_decap_8 FILLER_60_853 ();
 sg13g2_decap_8 FILLER_60_860 ();
 sg13g2_fill_1 FILLER_60_872 ();
 sg13g2_decap_8 FILLER_60_915 ();
 sg13g2_decap_8 FILLER_60_922 ();
 sg13g2_fill_2 FILLER_60_936 ();
 sg13g2_decap_4 FILLER_60_944 ();
 sg13g2_fill_1 FILLER_60_964 ();
 sg13g2_decap_8 FILLER_60_998 ();
 sg13g2_decap_8 FILLER_60_1005 ();
 sg13g2_decap_8 FILLER_60_1012 ();
 sg13g2_decap_4 FILLER_60_1019 ();
 sg13g2_fill_2 FILLER_60_1023 ();
 sg13g2_decap_4 FILLER_60_1042 ();
 sg13g2_fill_1 FILLER_60_1054 ();
 sg13g2_fill_2 FILLER_60_1061 ();
 sg13g2_fill_2 FILLER_60_1072 ();
 sg13g2_fill_1 FILLER_60_1074 ();
 sg13g2_fill_1 FILLER_60_1088 ();
 sg13g2_fill_2 FILLER_60_1093 ();
 sg13g2_fill_2 FILLER_60_1098 ();
 sg13g2_fill_1 FILLER_60_1100 ();
 sg13g2_fill_1 FILLER_60_1110 ();
 sg13g2_fill_1 FILLER_60_1117 ();
 sg13g2_fill_1 FILLER_60_1136 ();
 sg13g2_decap_8 FILLER_60_1167 ();
 sg13g2_fill_1 FILLER_60_1174 ();
 sg13g2_fill_1 FILLER_60_1198 ();
 sg13g2_fill_1 FILLER_60_1212 ();
 sg13g2_fill_1 FILLER_60_1246 ();
 sg13g2_fill_1 FILLER_60_1250 ();
 sg13g2_decap_8 FILLER_60_1261 ();
 sg13g2_fill_2 FILLER_60_1268 ();
 sg13g2_fill_2 FILLER_60_1290 ();
 sg13g2_fill_1 FILLER_60_1292 ();
 sg13g2_fill_2 FILLER_60_1305 ();
 sg13g2_fill_1 FILLER_60_1315 ();
 sg13g2_fill_2 FILLER_60_1335 ();
 sg13g2_fill_2 FILLER_60_1395 ();
 sg13g2_decap_8 FILLER_60_1427 ();
 sg13g2_fill_1 FILLER_60_1434 ();
 sg13g2_fill_1 FILLER_60_1441 ();
 sg13g2_fill_1 FILLER_60_1451 ();
 sg13g2_decap_4 FILLER_60_1504 ();
 sg13g2_decap_4 FILLER_60_1538 ();
 sg13g2_fill_1 FILLER_60_1542 ();
 sg13g2_fill_2 FILLER_60_1574 ();
 sg13g2_fill_1 FILLER_60_1576 ();
 sg13g2_decap_8 FILLER_60_1581 ();
 sg13g2_fill_2 FILLER_60_1588 ();
 sg13g2_decap_4 FILLER_60_1631 ();
 sg13g2_fill_1 FILLER_60_1635 ();
 sg13g2_fill_2 FILLER_60_1646 ();
 sg13g2_decap_8 FILLER_60_1678 ();
 sg13g2_fill_2 FILLER_60_1685 ();
 sg13g2_decap_8 FILLER_60_1692 ();
 sg13g2_decap_8 FILLER_60_1699 ();
 sg13g2_decap_4 FILLER_60_1706 ();
 sg13g2_fill_2 FILLER_60_1710 ();
 sg13g2_decap_4 FILLER_60_1720 ();
 sg13g2_decap_8 FILLER_60_1750 ();
 sg13g2_decap_8 FILLER_60_1757 ();
 sg13g2_fill_1 FILLER_60_1794 ();
 sg13g2_fill_1 FILLER_60_1798 ();
 sg13g2_decap_8 FILLER_60_1803 ();
 sg13g2_decap_8 FILLER_60_1810 ();
 sg13g2_fill_1 FILLER_60_1817 ();
 sg13g2_decap_8 FILLER_60_1848 ();
 sg13g2_decap_8 FILLER_60_1855 ();
 sg13g2_decap_4 FILLER_60_1862 ();
 sg13g2_decap_4 FILLER_60_1879 ();
 sg13g2_fill_1 FILLER_60_1883 ();
 sg13g2_fill_1 FILLER_60_1906 ();
 sg13g2_fill_1 FILLER_60_1924 ();
 sg13g2_fill_2 FILLER_60_1956 ();
 sg13g2_fill_2 FILLER_60_1984 ();
 sg13g2_fill_1 FILLER_60_1990 ();
 sg13g2_decap_4 FILLER_60_1995 ();
 sg13g2_fill_2 FILLER_60_1999 ();
 sg13g2_decap_8 FILLER_60_2019 ();
 sg13g2_decap_8 FILLER_60_2030 ();
 sg13g2_decap_4 FILLER_60_2037 ();
 sg13g2_fill_2 FILLER_60_2041 ();
 sg13g2_decap_4 FILLER_60_2083 ();
 sg13g2_decap_8 FILLER_60_2092 ();
 sg13g2_fill_1 FILLER_60_2099 ();
 sg13g2_fill_1 FILLER_60_2105 ();
 sg13g2_decap_4 FILLER_60_2115 ();
 sg13g2_fill_1 FILLER_60_2119 ();
 sg13g2_decap_8 FILLER_60_2155 ();
 sg13g2_fill_1 FILLER_60_2162 ();
 sg13g2_decap_4 FILLER_60_2168 ();
 sg13g2_decap_8 FILLER_60_2176 ();
 sg13g2_decap_8 FILLER_60_2208 ();
 sg13g2_decap_4 FILLER_60_2215 ();
 sg13g2_fill_2 FILLER_60_2250 ();
 sg13g2_fill_1 FILLER_60_2252 ();
 sg13g2_decap_8 FILLER_60_2288 ();
 sg13g2_decap_4 FILLER_60_2295 ();
 sg13g2_fill_1 FILLER_60_2299 ();
 sg13g2_decap_8 FILLER_60_2326 ();
 sg13g2_decap_4 FILLER_60_2333 ();
 sg13g2_decap_8 FILLER_60_2378 ();
 sg13g2_fill_2 FILLER_60_2385 ();
 sg13g2_fill_2 FILLER_60_2392 ();
 sg13g2_decap_4 FILLER_60_2398 ();
 sg13g2_fill_2 FILLER_60_2402 ();
 sg13g2_fill_2 FILLER_60_2428 ();
 sg13g2_decap_8 FILLER_60_2440 ();
 sg13g2_decap_8 FILLER_60_2447 ();
 sg13g2_fill_2 FILLER_60_2454 ();
 sg13g2_fill_2 FILLER_60_2464 ();
 sg13g2_fill_1 FILLER_60_2466 ();
 sg13g2_fill_2 FILLER_60_2511 ();
 sg13g2_fill_1 FILLER_60_2513 ();
 sg13g2_decap_8 FILLER_60_2522 ();
 sg13g2_decap_8 FILLER_60_2529 ();
 sg13g2_fill_1 FILLER_60_2536 ();
 sg13g2_decap_8 FILLER_60_2541 ();
 sg13g2_fill_2 FILLER_60_2548 ();
 sg13g2_fill_1 FILLER_60_2550 ();
 sg13g2_decap_8 FILLER_60_2554 ();
 sg13g2_fill_1 FILLER_60_2561 ();
 sg13g2_decap_8 FILLER_60_2567 ();
 sg13g2_decap_8 FILLER_60_2591 ();
 sg13g2_decap_8 FILLER_60_2598 ();
 sg13g2_decap_8 FILLER_60_2605 ();
 sg13g2_decap_8 FILLER_60_2620 ();
 sg13g2_decap_8 FILLER_60_2627 ();
 sg13g2_decap_8 FILLER_60_2634 ();
 sg13g2_decap_8 FILLER_60_2641 ();
 sg13g2_decap_8 FILLER_60_2648 ();
 sg13g2_decap_8 FILLER_60_2655 ();
 sg13g2_decap_8 FILLER_60_2662 ();
 sg13g2_fill_1 FILLER_60_2669 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_4 FILLER_61_14 ();
 sg13g2_fill_1 FILLER_61_18 ();
 sg13g2_fill_1 FILLER_61_54 ();
 sg13g2_fill_2 FILLER_61_99 ();
 sg13g2_fill_1 FILLER_61_111 ();
 sg13g2_fill_1 FILLER_61_121 ();
 sg13g2_fill_1 FILLER_61_183 ();
 sg13g2_fill_2 FILLER_61_189 ();
 sg13g2_fill_1 FILLER_61_196 ();
 sg13g2_fill_1 FILLER_61_202 ();
 sg13g2_fill_1 FILLER_61_208 ();
 sg13g2_fill_1 FILLER_61_213 ();
 sg13g2_fill_1 FILLER_61_219 ();
 sg13g2_fill_2 FILLER_61_225 ();
 sg13g2_fill_1 FILLER_61_227 ();
 sg13g2_decap_8 FILLER_61_231 ();
 sg13g2_decap_4 FILLER_61_238 ();
 sg13g2_decap_8 FILLER_61_247 ();
 sg13g2_fill_1 FILLER_61_254 ();
 sg13g2_decap_8 FILLER_61_308 ();
 sg13g2_decap_8 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_322 ();
 sg13g2_decap_4 FILLER_61_329 ();
 sg13g2_fill_2 FILLER_61_337 ();
 sg13g2_fill_1 FILLER_61_355 ();
 sg13g2_fill_2 FILLER_61_365 ();
 sg13g2_decap_8 FILLER_61_371 ();
 sg13g2_decap_8 FILLER_61_378 ();
 sg13g2_decap_8 FILLER_61_385 ();
 sg13g2_decap_4 FILLER_61_422 ();
 sg13g2_decap_8 FILLER_61_439 ();
 sg13g2_decap_8 FILLER_61_446 ();
 sg13g2_decap_8 FILLER_61_453 ();
 sg13g2_decap_8 FILLER_61_460 ();
 sg13g2_decap_8 FILLER_61_467 ();
 sg13g2_decap_8 FILLER_61_474 ();
 sg13g2_decap_4 FILLER_61_481 ();
 sg13g2_fill_1 FILLER_61_485 ();
 sg13g2_decap_8 FILLER_61_522 ();
 sg13g2_fill_2 FILLER_61_529 ();
 sg13g2_fill_1 FILLER_61_531 ();
 sg13g2_decap_4 FILLER_61_559 ();
 sg13g2_fill_1 FILLER_61_563 ();
 sg13g2_decap_8 FILLER_61_574 ();
 sg13g2_decap_8 FILLER_61_581 ();
 sg13g2_decap_8 FILLER_61_588 ();
 sg13g2_decap_8 FILLER_61_595 ();
 sg13g2_fill_2 FILLER_61_602 ();
 sg13g2_fill_1 FILLER_61_604 ();
 sg13g2_fill_1 FILLER_61_623 ();
 sg13g2_fill_2 FILLER_61_628 ();
 sg13g2_fill_1 FILLER_61_630 ();
 sg13g2_fill_1 FILLER_61_635 ();
 sg13g2_fill_1 FILLER_61_641 ();
 sg13g2_fill_2 FILLER_61_655 ();
 sg13g2_fill_1 FILLER_61_657 ();
 sg13g2_decap_8 FILLER_61_663 ();
 sg13g2_fill_2 FILLER_61_670 ();
 sg13g2_fill_1 FILLER_61_672 ();
 sg13g2_decap_8 FILLER_61_677 ();
 sg13g2_decap_4 FILLER_61_684 ();
 sg13g2_fill_2 FILLER_61_693 ();
 sg13g2_fill_1 FILLER_61_695 ();
 sg13g2_decap_8 FILLER_61_706 ();
 sg13g2_fill_2 FILLER_61_713 ();
 sg13g2_decap_8 FILLER_61_720 ();
 sg13g2_fill_2 FILLER_61_732 ();
 sg13g2_fill_1 FILLER_61_745 ();
 sg13g2_fill_2 FILLER_61_759 ();
 sg13g2_fill_2 FILLER_61_765 ();
 sg13g2_fill_1 FILLER_61_801 ();
 sg13g2_decap_4 FILLER_61_838 ();
 sg13g2_fill_2 FILLER_61_880 ();
 sg13g2_fill_1 FILLER_61_882 ();
 sg13g2_fill_2 FILLER_61_914 ();
 sg13g2_decap_4 FILLER_61_923 ();
 sg13g2_fill_2 FILLER_61_927 ();
 sg13g2_fill_1 FILLER_61_965 ();
 sg13g2_fill_2 FILLER_61_983 ();
 sg13g2_decap_8 FILLER_61_994 ();
 sg13g2_decap_8 FILLER_61_1001 ();
 sg13g2_decap_4 FILLER_61_1008 ();
 sg13g2_decap_4 FILLER_61_1022 ();
 sg13g2_fill_1 FILLER_61_1031 ();
 sg13g2_fill_1 FILLER_61_1037 ();
 sg13g2_fill_1 FILLER_61_1042 ();
 sg13g2_fill_1 FILLER_61_1047 ();
 sg13g2_fill_1 FILLER_61_1079 ();
 sg13g2_fill_2 FILLER_61_1124 ();
 sg13g2_decap_8 FILLER_61_1154 ();
 sg13g2_decap_4 FILLER_61_1161 ();
 sg13g2_fill_1 FILLER_61_1165 ();
 sg13g2_fill_2 FILLER_61_1171 ();
 sg13g2_fill_1 FILLER_61_1173 ();
 sg13g2_fill_2 FILLER_61_1184 ();
 sg13g2_fill_1 FILLER_61_1253 ();
 sg13g2_fill_2 FILLER_61_1313 ();
 sg13g2_decap_8 FILLER_61_1331 ();
 sg13g2_fill_2 FILLER_61_1338 ();
 sg13g2_decap_4 FILLER_61_1349 ();
 sg13g2_fill_1 FILLER_61_1353 ();
 sg13g2_fill_1 FILLER_61_1359 ();
 sg13g2_fill_2 FILLER_61_1397 ();
 sg13g2_fill_1 FILLER_61_1399 ();
 sg13g2_fill_2 FILLER_61_1409 ();
 sg13g2_fill_1 FILLER_61_1411 ();
 sg13g2_decap_8 FILLER_61_1417 ();
 sg13g2_decap_8 FILLER_61_1424 ();
 sg13g2_decap_8 FILLER_61_1440 ();
 sg13g2_fill_2 FILLER_61_1447 ();
 sg13g2_fill_2 FILLER_61_1457 ();
 sg13g2_fill_2 FILLER_61_1480 ();
 sg13g2_fill_2 FILLER_61_1486 ();
 sg13g2_fill_1 FILLER_61_1488 ();
 sg13g2_decap_4 FILLER_61_1493 ();
 sg13g2_fill_1 FILLER_61_1501 ();
 sg13g2_fill_2 FILLER_61_1515 ();
 sg13g2_fill_1 FILLER_61_1517 ();
 sg13g2_decap_8 FILLER_61_1522 ();
 sg13g2_decap_8 FILLER_61_1529 ();
 sg13g2_fill_1 FILLER_61_1536 ();
 sg13g2_decap_4 FILLER_61_1542 ();
 sg13g2_decap_4 FILLER_61_1550 ();
 sg13g2_fill_1 FILLER_61_1567 ();
 sg13g2_decap_8 FILLER_61_1573 ();
 sg13g2_fill_2 FILLER_61_1584 ();
 sg13g2_fill_1 FILLER_61_1586 ();
 sg13g2_fill_2 FILLER_61_1591 ();
 sg13g2_decap_4 FILLER_61_1601 ();
 sg13g2_fill_2 FILLER_61_1605 ();
 sg13g2_decap_8 FILLER_61_1615 ();
 sg13g2_decap_8 FILLER_61_1622 ();
 sg13g2_decap_8 FILLER_61_1629 ();
 sg13g2_decap_4 FILLER_61_1636 ();
 sg13g2_fill_1 FILLER_61_1640 ();
 sg13g2_decap_8 FILLER_61_1650 ();
 sg13g2_fill_2 FILLER_61_1657 ();
 sg13g2_fill_1 FILLER_61_1659 ();
 sg13g2_decap_8 FILLER_61_1664 ();
 sg13g2_fill_2 FILLER_61_1671 ();
 sg13g2_fill_1 FILLER_61_1673 ();
 sg13g2_decap_8 FILLER_61_1679 ();
 sg13g2_decap_4 FILLER_61_1686 ();
 sg13g2_decap_8 FILLER_61_1725 ();
 sg13g2_decap_8 FILLER_61_1732 ();
 sg13g2_decap_8 FILLER_61_1739 ();
 sg13g2_decap_8 FILLER_61_1807 ();
 sg13g2_fill_2 FILLER_61_1814 ();
 sg13g2_fill_1 FILLER_61_1816 ();
 sg13g2_fill_1 FILLER_61_1843 ();
 sg13g2_fill_2 FILLER_61_1849 ();
 sg13g2_fill_1 FILLER_61_1856 ();
 sg13g2_decap_8 FILLER_61_1861 ();
 sg13g2_decap_8 FILLER_61_1868 ();
 sg13g2_decap_8 FILLER_61_1875 ();
 sg13g2_decap_8 FILLER_61_1882 ();
 sg13g2_decap_8 FILLER_61_1889 ();
 sg13g2_fill_2 FILLER_61_1896 ();
 sg13g2_fill_1 FILLER_61_1904 ();
 sg13g2_fill_1 FILLER_61_1923 ();
 sg13g2_decap_4 FILLER_61_1929 ();
 sg13g2_fill_1 FILLER_61_1933 ();
 sg13g2_fill_1 FILLER_61_1948 ();
 sg13g2_fill_2 FILLER_61_1963 ();
 sg13g2_fill_1 FILLER_61_1965 ();
 sg13g2_decap_4 FILLER_61_1997 ();
 sg13g2_decap_8 FILLER_61_2041 ();
 sg13g2_decap_4 FILLER_61_2048 ();
 sg13g2_fill_1 FILLER_61_2052 ();
 sg13g2_decap_4 FILLER_61_2058 ();
 sg13g2_fill_2 FILLER_61_2072 ();
 sg13g2_fill_2 FILLER_61_2078 ();
 sg13g2_fill_1 FILLER_61_2087 ();
 sg13g2_decap_4 FILLER_61_2114 ();
 sg13g2_fill_2 FILLER_61_2127 ();
 sg13g2_fill_1 FILLER_61_2129 ();
 sg13g2_decap_8 FILLER_61_2148 ();
 sg13g2_decap_8 FILLER_61_2155 ();
 sg13g2_decap_4 FILLER_61_2162 ();
 sg13g2_decap_8 FILLER_61_2206 ();
 sg13g2_decap_8 FILLER_61_2213 ();
 sg13g2_fill_2 FILLER_61_2224 ();
 sg13g2_fill_1 FILLER_61_2231 ();
 sg13g2_fill_1 FILLER_61_2237 ();
 sg13g2_fill_2 FILLER_61_2242 ();
 sg13g2_fill_1 FILLER_61_2244 ();
 sg13g2_decap_8 FILLER_61_2269 ();
 sg13g2_decap_8 FILLER_61_2276 ();
 sg13g2_fill_2 FILLER_61_2283 ();
 sg13g2_decap_4 FILLER_61_2320 ();
 sg13g2_decap_8 FILLER_61_2330 ();
 sg13g2_fill_1 FILLER_61_2413 ();
 sg13g2_fill_2 FILLER_61_2444 ();
 sg13g2_fill_1 FILLER_61_2451 ();
 sg13g2_fill_2 FILLER_61_2478 ();
 sg13g2_fill_2 FILLER_61_2506 ();
 sg13g2_fill_2 FILLER_61_2513 ();
 sg13g2_fill_1 FILLER_61_2515 ();
 sg13g2_fill_2 FILLER_61_2564 ();
 sg13g2_fill_1 FILLER_61_2566 ();
 sg13g2_decap_4 FILLER_61_2571 ();
 sg13g2_fill_1 FILLER_61_2575 ();
 sg13g2_decap_4 FILLER_61_2606 ();
 sg13g2_fill_2 FILLER_61_2610 ();
 sg13g2_fill_2 FILLER_61_2616 ();
 sg13g2_fill_1 FILLER_61_2618 ();
 sg13g2_decap_8 FILLER_61_2645 ();
 sg13g2_decap_8 FILLER_61_2652 ();
 sg13g2_decap_8 FILLER_61_2659 ();
 sg13g2_decap_4 FILLER_61_2666 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_fill_1 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_27 ();
 sg13g2_fill_1 FILLER_62_34 ();
 sg13g2_fill_2 FILLER_62_45 ();
 sg13g2_fill_1 FILLER_62_52 ();
 sg13g2_fill_1 FILLER_62_58 ();
 sg13g2_decap_4 FILLER_62_101 ();
 sg13g2_fill_1 FILLER_62_105 ();
 sg13g2_fill_1 FILLER_62_120 ();
 sg13g2_fill_2 FILLER_62_134 ();
 sg13g2_fill_1 FILLER_62_160 ();
 sg13g2_fill_1 FILLER_62_165 ();
 sg13g2_decap_4 FILLER_62_181 ();
 sg13g2_fill_1 FILLER_62_190 ();
 sg13g2_decap_8 FILLER_62_196 ();
 sg13g2_fill_1 FILLER_62_208 ();
 sg13g2_fill_2 FILLER_62_217 ();
 sg13g2_fill_2 FILLER_62_223 ();
 sg13g2_fill_1 FILLER_62_225 ();
 sg13g2_fill_2 FILLER_62_235 ();
 sg13g2_fill_2 FILLER_62_241 ();
 sg13g2_decap_4 FILLER_62_248 ();
 sg13g2_fill_2 FILLER_62_268 ();
 sg13g2_fill_1 FILLER_62_270 ();
 sg13g2_decap_8 FILLER_62_275 ();
 sg13g2_decap_8 FILLER_62_282 ();
 sg13g2_fill_1 FILLER_62_289 ();
 sg13g2_decap_8 FILLER_62_330 ();
 sg13g2_decap_8 FILLER_62_337 ();
 sg13g2_decap_8 FILLER_62_344 ();
 sg13g2_fill_2 FILLER_62_351 ();
 sg13g2_decap_8 FILLER_62_360 ();
 sg13g2_fill_1 FILLER_62_367 ();
 sg13g2_fill_1 FILLER_62_373 ();
 sg13g2_fill_2 FILLER_62_379 ();
 sg13g2_fill_1 FILLER_62_419 ();
 sg13g2_decap_8 FILLER_62_425 ();
 sg13g2_decap_8 FILLER_62_432 ();
 sg13g2_decap_8 FILLER_62_439 ();
 sg13g2_decap_8 FILLER_62_446 ();
 sg13g2_decap_8 FILLER_62_453 ();
 sg13g2_fill_2 FILLER_62_460 ();
 sg13g2_fill_2 FILLER_62_472 ();
 sg13g2_fill_1 FILLER_62_474 ();
 sg13g2_decap_8 FILLER_62_493 ();
 sg13g2_fill_2 FILLER_62_504 ();
 sg13g2_fill_1 FILLER_62_506 ();
 sg13g2_decap_8 FILLER_62_512 ();
 sg13g2_decap_4 FILLER_62_519 ();
 sg13g2_decap_8 FILLER_62_559 ();
 sg13g2_decap_4 FILLER_62_566 ();
 sg13g2_decap_8 FILLER_62_600 ();
 sg13g2_fill_1 FILLER_62_607 ();
 sg13g2_fill_1 FILLER_62_612 ();
 sg13g2_decap_8 FILLER_62_635 ();
 sg13g2_fill_2 FILLER_62_642 ();
 sg13g2_fill_2 FILLER_62_688 ();
 sg13g2_decap_4 FILLER_62_693 ();
 sg13g2_decap_8 FILLER_62_701 ();
 sg13g2_decap_8 FILLER_62_714 ();
 sg13g2_fill_2 FILLER_62_721 ();
 sg13g2_fill_1 FILLER_62_723 ();
 sg13g2_decap_4 FILLER_62_728 ();
 sg13g2_fill_2 FILLER_62_732 ();
 sg13g2_fill_2 FILLER_62_811 ();
 sg13g2_fill_1 FILLER_62_813 ();
 sg13g2_fill_1 FILLER_62_825 ();
 sg13g2_decap_4 FILLER_62_837 ();
 sg13g2_fill_2 FILLER_62_841 ();
 sg13g2_fill_2 FILLER_62_859 ();
 sg13g2_decap_8 FILLER_62_865 ();
 sg13g2_decap_4 FILLER_62_872 ();
 sg13g2_fill_1 FILLER_62_876 ();
 sg13g2_decap_8 FILLER_62_936 ();
 sg13g2_decap_8 FILLER_62_943 ();
 sg13g2_decap_8 FILLER_62_950 ();
 sg13g2_fill_2 FILLER_62_957 ();
 sg13g2_fill_1 FILLER_62_959 ();
 sg13g2_fill_1 FILLER_62_973 ();
 sg13g2_decap_8 FILLER_62_978 ();
 sg13g2_decap_4 FILLER_62_985 ();
 sg13g2_fill_1 FILLER_62_989 ();
 sg13g2_fill_2 FILLER_62_1016 ();
 sg13g2_decap_4 FILLER_62_1023 ();
 sg13g2_fill_2 FILLER_62_1032 ();
 sg13g2_fill_2 FILLER_62_1053 ();
 sg13g2_fill_1 FILLER_62_1055 ();
 sg13g2_fill_1 FILLER_62_1065 ();
 sg13g2_fill_2 FILLER_62_1071 ();
 sg13g2_fill_1 FILLER_62_1078 ();
 sg13g2_fill_2 FILLER_62_1084 ();
 sg13g2_fill_1 FILLER_62_1091 ();
 sg13g2_fill_1 FILLER_62_1118 ();
 sg13g2_decap_8 FILLER_62_1153 ();
 sg13g2_decap_8 FILLER_62_1160 ();
 sg13g2_fill_1 FILLER_62_1167 ();
 sg13g2_decap_4 FILLER_62_1199 ();
 sg13g2_fill_1 FILLER_62_1203 ();
 sg13g2_fill_2 FILLER_62_1207 ();
 sg13g2_decap_4 FILLER_62_1226 ();
 sg13g2_fill_1 FILLER_62_1237 ();
 sg13g2_fill_2 FILLER_62_1245 ();
 sg13g2_fill_2 FILLER_62_1257 ();
 sg13g2_fill_2 FILLER_62_1281 ();
 sg13g2_fill_1 FILLER_62_1283 ();
 sg13g2_fill_2 FILLER_62_1288 ();
 sg13g2_fill_1 FILLER_62_1316 ();
 sg13g2_fill_2 FILLER_62_1343 ();
 sg13g2_fill_1 FILLER_62_1345 ();
 sg13g2_decap_4 FILLER_62_1363 ();
 sg13g2_fill_1 FILLER_62_1367 ();
 sg13g2_fill_2 FILLER_62_1374 ();
 sg13g2_fill_1 FILLER_62_1376 ();
 sg13g2_decap_8 FILLER_62_1383 ();
 sg13g2_fill_2 FILLER_62_1395 ();
 sg13g2_decap_4 FILLER_62_1411 ();
 sg13g2_fill_2 FILLER_62_1415 ();
 sg13g2_fill_2 FILLER_62_1457 ();
 sg13g2_fill_1 FILLER_62_1459 ();
 sg13g2_fill_2 FILLER_62_1475 ();
 sg13g2_fill_1 FILLER_62_1477 ();
 sg13g2_decap_4 FILLER_62_1483 ();
 sg13g2_decap_4 FILLER_62_1492 ();
 sg13g2_fill_1 FILLER_62_1496 ();
 sg13g2_decap_4 FILLER_62_1502 ();
 sg13g2_decap_4 FILLER_62_1532 ();
 sg13g2_fill_2 FILLER_62_1562 ();
 sg13g2_decap_4 FILLER_62_1597 ();
 sg13g2_fill_2 FILLER_62_1601 ();
 sg13g2_decap_8 FILLER_62_1638 ();
 sg13g2_decap_8 FILLER_62_1645 ();
 sg13g2_decap_8 FILLER_62_1652 ();
 sg13g2_fill_2 FILLER_62_1659 ();
 sg13g2_fill_1 FILLER_62_1661 ();
 sg13g2_decap_4 FILLER_62_1666 ();
 sg13g2_decap_4 FILLER_62_1696 ();
 sg13g2_fill_2 FILLER_62_1700 ();
 sg13g2_decap_8 FILLER_62_1706 ();
 sg13g2_decap_8 FILLER_62_1713 ();
 sg13g2_decap_8 FILLER_62_1720 ();
 sg13g2_decap_8 FILLER_62_1727 ();
 sg13g2_decap_8 FILLER_62_1734 ();
 sg13g2_decap_8 FILLER_62_1741 ();
 sg13g2_decap_8 FILLER_62_1748 ();
 sg13g2_decap_4 FILLER_62_1755 ();
 sg13g2_fill_2 FILLER_62_1773 ();
 sg13g2_fill_1 FILLER_62_1775 ();
 sg13g2_decap_8 FILLER_62_1782 ();
 sg13g2_fill_2 FILLER_62_1789 ();
 sg13g2_fill_2 FILLER_62_1809 ();
 sg13g2_fill_1 FILLER_62_1811 ();
 sg13g2_fill_2 FILLER_62_1817 ();
 sg13g2_decap_4 FILLER_62_1823 ();
 sg13g2_decap_8 FILLER_62_1836 ();
 sg13g2_fill_1 FILLER_62_1843 ();
 sg13g2_decap_4 FILLER_62_1870 ();
 sg13g2_fill_1 FILLER_62_1874 ();
 sg13g2_fill_2 FILLER_62_1880 ();
 sg13g2_fill_1 FILLER_62_1882 ();
 sg13g2_fill_2 FILLER_62_1888 ();
 sg13g2_fill_1 FILLER_62_1916 ();
 sg13g2_decap_8 FILLER_62_1948 ();
 sg13g2_decap_8 FILLER_62_1955 ();
 sg13g2_decap_8 FILLER_62_1962 ();
 sg13g2_decap_8 FILLER_62_1969 ();
 sg13g2_decap_4 FILLER_62_1976 ();
 sg13g2_decap_4 FILLER_62_1990 ();
 sg13g2_fill_1 FILLER_62_1994 ();
 sg13g2_fill_2 FILLER_62_2012 ();
 sg13g2_fill_1 FILLER_62_2014 ();
 sg13g2_decap_4 FILLER_62_2041 ();
 sg13g2_decap_4 FILLER_62_2071 ();
 sg13g2_fill_2 FILLER_62_2115 ();
 sg13g2_fill_1 FILLER_62_2117 ();
 sg13g2_fill_1 FILLER_62_2153 ();
 sg13g2_fill_2 FILLER_62_2215 ();
 sg13g2_fill_1 FILLER_62_2217 ();
 sg13g2_decap_8 FILLER_62_2244 ();
 sg13g2_fill_2 FILLER_62_2251 ();
 sg13g2_decap_8 FILLER_62_2258 ();
 sg13g2_fill_1 FILLER_62_2265 ();
 sg13g2_decap_8 FILLER_62_2287 ();
 sg13g2_fill_2 FILLER_62_2294 ();
 sg13g2_fill_1 FILLER_62_2296 ();
 sg13g2_decap_8 FILLER_62_2335 ();
 sg13g2_fill_2 FILLER_62_2342 ();
 sg13g2_fill_1 FILLER_62_2353 ();
 sg13g2_decap_8 FILLER_62_2385 ();
 sg13g2_decap_8 FILLER_62_2392 ();
 sg13g2_fill_2 FILLER_62_2399 ();
 sg13g2_fill_1 FILLER_62_2401 ();
 sg13g2_decap_8 FILLER_62_2405 ();
 sg13g2_fill_2 FILLER_62_2412 ();
 sg13g2_fill_1 FILLER_62_2440 ();
 sg13g2_fill_1 FILLER_62_2446 ();
 sg13g2_fill_2 FILLER_62_2457 ();
 sg13g2_decap_8 FILLER_62_2510 ();
 sg13g2_fill_1 FILLER_62_2517 ();
 sg13g2_decap_8 FILLER_62_2544 ();
 sg13g2_decap_8 FILLER_62_2551 ();
 sg13g2_decap_8 FILLER_62_2558 ();
 sg13g2_fill_1 FILLER_62_2565 ();
 sg13g2_fill_1 FILLER_62_2599 ();
 sg13g2_decap_8 FILLER_62_2634 ();
 sg13g2_decap_8 FILLER_62_2641 ();
 sg13g2_decap_8 FILLER_62_2648 ();
 sg13g2_decap_8 FILLER_62_2655 ();
 sg13g2_decap_8 FILLER_62_2662 ();
 sg13g2_fill_1 FILLER_62_2669 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_7 ();
 sg13g2_fill_1 FILLER_63_9 ();
 sg13g2_fill_1 FILLER_63_23 ();
 sg13g2_fill_1 FILLER_63_32 ();
 sg13g2_fill_1 FILLER_63_37 ();
 sg13g2_fill_1 FILLER_63_44 ();
 sg13g2_fill_2 FILLER_63_49 ();
 sg13g2_fill_1 FILLER_63_51 ();
 sg13g2_fill_1 FILLER_63_57 ();
 sg13g2_fill_2 FILLER_63_65 ();
 sg13g2_fill_2 FILLER_63_72 ();
 sg13g2_fill_2 FILLER_63_84 ();
 sg13g2_fill_1 FILLER_63_103 ();
 sg13g2_fill_1 FILLER_63_109 ();
 sg13g2_fill_1 FILLER_63_114 ();
 sg13g2_decap_4 FILLER_63_120 ();
 sg13g2_fill_1 FILLER_63_139 ();
 sg13g2_fill_2 FILLER_63_151 ();
 sg13g2_fill_1 FILLER_63_153 ();
 sg13g2_fill_2 FILLER_63_159 ();
 sg13g2_fill_1 FILLER_63_165 ();
 sg13g2_fill_1 FILLER_63_171 ();
 sg13g2_fill_1 FILLER_63_194 ();
 sg13g2_fill_2 FILLER_63_212 ();
 sg13g2_decap_4 FILLER_63_219 ();
 sg13g2_fill_2 FILLER_63_223 ();
 sg13g2_fill_2 FILLER_63_234 ();
 sg13g2_decap_8 FILLER_63_241 ();
 sg13g2_decap_8 FILLER_63_248 ();
 sg13g2_decap_8 FILLER_63_255 ();
 sg13g2_decap_8 FILLER_63_262 ();
 sg13g2_decap_8 FILLER_63_269 ();
 sg13g2_decap_8 FILLER_63_276 ();
 sg13g2_fill_2 FILLER_63_283 ();
 sg13g2_decap_8 FILLER_63_311 ();
 sg13g2_decap_8 FILLER_63_318 ();
 sg13g2_decap_8 FILLER_63_330 ();
 sg13g2_decap_8 FILLER_63_337 ();
 sg13g2_fill_2 FILLER_63_370 ();
 sg13g2_decap_8 FILLER_63_381 ();
 sg13g2_decap_8 FILLER_63_388 ();
 sg13g2_decap_8 FILLER_63_395 ();
 sg13g2_decap_8 FILLER_63_402 ();
 sg13g2_fill_1 FILLER_63_409 ();
 sg13g2_fill_2 FILLER_63_414 ();
 sg13g2_fill_2 FILLER_63_420 ();
 sg13g2_decap_8 FILLER_63_443 ();
 sg13g2_decap_4 FILLER_63_457 ();
 sg13g2_decap_8 FILLER_63_469 ();
 sg13g2_decap_8 FILLER_63_476 ();
 sg13g2_decap_8 FILLER_63_483 ();
 sg13g2_fill_2 FILLER_63_490 ();
 sg13g2_fill_2 FILLER_63_497 ();
 sg13g2_fill_1 FILLER_63_499 ();
 sg13g2_decap_8 FILLER_63_505 ();
 sg13g2_decap_4 FILLER_63_512 ();
 sg13g2_fill_2 FILLER_63_516 ();
 sg13g2_decap_4 FILLER_63_523 ();
 sg13g2_decap_8 FILLER_63_557 ();
 sg13g2_decap_8 FILLER_63_564 ();
 sg13g2_decap_8 FILLER_63_571 ();
 sg13g2_decap_8 FILLER_63_578 ();
 sg13g2_decap_8 FILLER_63_585 ();
 sg13g2_fill_1 FILLER_63_592 ();
 sg13g2_fill_1 FILLER_63_603 ();
 sg13g2_decap_8 FILLER_63_642 ();
 sg13g2_fill_1 FILLER_63_649 ();
 sg13g2_fill_2 FILLER_63_658 ();
 sg13g2_fill_1 FILLER_63_660 ();
 sg13g2_decap_4 FILLER_63_665 ();
 sg13g2_fill_1 FILLER_63_669 ();
 sg13g2_fill_2 FILLER_63_697 ();
 sg13g2_fill_2 FILLER_63_711 ();
 sg13g2_fill_1 FILLER_63_739 ();
 sg13g2_decap_4 FILLER_63_767 ();
 sg13g2_fill_2 FILLER_63_832 ();
 sg13g2_decap_8 FILLER_63_844 ();
 sg13g2_decap_4 FILLER_63_851 ();
 sg13g2_fill_1 FILLER_63_855 ();
 sg13g2_fill_1 FILLER_63_860 ();
 sg13g2_decap_8 FILLER_63_864 ();
 sg13g2_decap_8 FILLER_63_871 ();
 sg13g2_fill_2 FILLER_63_878 ();
 sg13g2_decap_8 FILLER_63_884 ();
 sg13g2_decap_8 FILLER_63_891 ();
 sg13g2_fill_2 FILLER_63_898 ();
 sg13g2_fill_1 FILLER_63_900 ();
 sg13g2_decap_8 FILLER_63_942 ();
 sg13g2_fill_1 FILLER_63_949 ();
 sg13g2_decap_4 FILLER_63_981 ();
 sg13g2_decap_4 FILLER_63_993 ();
 sg13g2_fill_2 FILLER_63_1002 ();
 sg13g2_fill_1 FILLER_63_1004 ();
 sg13g2_decap_8 FILLER_63_1009 ();
 sg13g2_fill_1 FILLER_63_1016 ();
 sg13g2_fill_2 FILLER_63_1022 ();
 sg13g2_fill_2 FILLER_63_1029 ();
 sg13g2_fill_1 FILLER_63_1031 ();
 sg13g2_fill_1 FILLER_63_1038 ();
 sg13g2_fill_2 FILLER_63_1049 ();
 sg13g2_decap_4 FILLER_63_1055 ();
 sg13g2_decap_8 FILLER_63_1063 ();
 sg13g2_fill_2 FILLER_63_1070 ();
 sg13g2_fill_1 FILLER_63_1072 ();
 sg13g2_decap_4 FILLER_63_1085 ();
 sg13g2_fill_2 FILLER_63_1089 ();
 sg13g2_decap_4 FILLER_63_1096 ();
 sg13g2_fill_1 FILLER_63_1100 ();
 sg13g2_decap_8 FILLER_63_1105 ();
 sg13g2_decap_4 FILLER_63_1112 ();
 sg13g2_fill_2 FILLER_63_1116 ();
 sg13g2_fill_2 FILLER_63_1121 ();
 sg13g2_fill_1 FILLER_63_1123 ();
 sg13g2_decap_4 FILLER_63_1128 ();
 sg13g2_fill_2 FILLER_63_1132 ();
 sg13g2_fill_2 FILLER_63_1141 ();
 sg13g2_fill_1 FILLER_63_1143 ();
 sg13g2_fill_2 FILLER_63_1157 ();
 sg13g2_fill_1 FILLER_63_1162 ();
 sg13g2_decap_8 FILLER_63_1168 ();
 sg13g2_decap_8 FILLER_63_1175 ();
 sg13g2_fill_1 FILLER_63_1212 ();
 sg13g2_fill_1 FILLER_63_1221 ();
 sg13g2_fill_1 FILLER_63_1229 ();
 sg13g2_fill_2 FILLER_63_1233 ();
 sg13g2_fill_1 FILLER_63_1235 ();
 sg13g2_fill_2 FILLER_63_1270 ();
 sg13g2_fill_1 FILLER_63_1272 ();
 sg13g2_fill_2 FILLER_63_1281 ();
 sg13g2_fill_2 FILLER_63_1288 ();
 sg13g2_fill_1 FILLER_63_1302 ();
 sg13g2_decap_8 FILLER_63_1335 ();
 sg13g2_fill_1 FILLER_63_1342 ();
 sg13g2_fill_2 FILLER_63_1347 ();
 sg13g2_fill_2 FILLER_63_1355 ();
 sg13g2_fill_1 FILLER_63_1357 ();
 sg13g2_fill_1 FILLER_63_1363 ();
 sg13g2_fill_2 FILLER_63_1370 ();
 sg13g2_decap_8 FILLER_63_1376 ();
 sg13g2_decap_4 FILLER_63_1383 ();
 sg13g2_fill_1 FILLER_63_1387 ();
 sg13g2_fill_2 FILLER_63_1402 ();
 sg13g2_fill_1 FILLER_63_1404 ();
 sg13g2_fill_2 FILLER_63_1422 ();
 sg13g2_fill_1 FILLER_63_1424 ();
 sg13g2_fill_2 FILLER_63_1429 ();
 sg13g2_fill_1 FILLER_63_1431 ();
 sg13g2_decap_4 FILLER_63_1436 ();
 sg13g2_fill_1 FILLER_63_1440 ();
 sg13g2_decap_4 FILLER_63_1454 ();
 sg13g2_fill_2 FILLER_63_1458 ();
 sg13g2_fill_1 FILLER_63_1468 ();
 sg13g2_decap_4 FILLER_63_1482 ();
 sg13g2_fill_1 FILLER_63_1486 ();
 sg13g2_fill_2 FILLER_63_1543 ();
 sg13g2_fill_2 FILLER_63_1569 ();
 sg13g2_decap_4 FILLER_63_1597 ();
 sg13g2_fill_2 FILLER_63_1606 ();
 sg13g2_fill_2 FILLER_63_1613 ();
 sg13g2_fill_2 FILLER_63_1620 ();
 sg13g2_fill_1 FILLER_63_1622 ();
 sg13g2_fill_1 FILLER_63_1627 ();
 sg13g2_fill_2 FILLER_63_1632 ();
 sg13g2_fill_1 FILLER_63_1634 ();
 sg13g2_decap_4 FILLER_63_1639 ();
 sg13g2_fill_2 FILLER_63_1643 ();
 sg13g2_decap_4 FILLER_63_1649 ();
 sg13g2_fill_2 FILLER_63_1653 ();
 sg13g2_decap_4 FILLER_63_1685 ();
 sg13g2_decap_8 FILLER_63_1697 ();
 sg13g2_decap_4 FILLER_63_1704 ();
 sg13g2_fill_2 FILLER_63_1708 ();
 sg13g2_decap_8 FILLER_63_1749 ();
 sg13g2_decap_8 FILLER_63_1756 ();
 sg13g2_fill_1 FILLER_63_1763 ();
 sg13g2_fill_1 FILLER_63_1769 ();
 sg13g2_fill_1 FILLER_63_1788 ();
 sg13g2_decap_4 FILLER_63_1800 ();
 sg13g2_decap_8 FILLER_63_1808 ();
 sg13g2_decap_8 FILLER_63_1819 ();
 sg13g2_decap_8 FILLER_63_1826 ();
 sg13g2_decap_8 FILLER_63_1833 ();
 sg13g2_decap_4 FILLER_63_1840 ();
 sg13g2_fill_1 FILLER_63_1844 ();
 sg13g2_decap_8 FILLER_63_1849 ();
 sg13g2_fill_1 FILLER_63_1856 ();
 sg13g2_decap_8 FILLER_63_1883 ();
 sg13g2_decap_4 FILLER_63_1890 ();
 sg13g2_fill_2 FILLER_63_1894 ();
 sg13g2_decap_4 FILLER_63_1906 ();
 sg13g2_fill_2 FILLER_63_1910 ();
 sg13g2_fill_2 FILLER_63_1941 ();
 sg13g2_fill_2 FILLER_63_1946 ();
 sg13g2_decap_4 FILLER_63_1955 ();
 sg13g2_fill_2 FILLER_63_1959 ();
 sg13g2_fill_2 FILLER_63_1970 ();
 sg13g2_decap_8 FILLER_63_1978 ();
 sg13g2_fill_1 FILLER_63_1985 ();
 sg13g2_decap_8 FILLER_63_1990 ();
 sg13g2_decap_4 FILLER_63_1997 ();
 sg13g2_decap_8 FILLER_63_2064 ();
 sg13g2_fill_1 FILLER_63_2071 ();
 sg13g2_decap_8 FILLER_63_2076 ();
 sg13g2_decap_8 FILLER_63_2083 ();
 sg13g2_decap_8 FILLER_63_2090 ();
 sg13g2_fill_1 FILLER_63_2097 ();
 sg13g2_fill_2 FILLER_63_2104 ();
 sg13g2_decap_8 FILLER_63_2115 ();
 sg13g2_decap_8 FILLER_63_2122 ();
 sg13g2_decap_4 FILLER_63_2129 ();
 sg13g2_decap_8 FILLER_63_2146 ();
 sg13g2_decap_8 FILLER_63_2153 ();
 sg13g2_decap_8 FILLER_63_2160 ();
 sg13g2_decap_8 FILLER_63_2167 ();
 sg13g2_decap_8 FILLER_63_2174 ();
 sg13g2_decap_4 FILLER_63_2181 ();
 sg13g2_fill_2 FILLER_63_2193 ();
 sg13g2_fill_1 FILLER_63_2195 ();
 sg13g2_fill_2 FILLER_63_2222 ();
 sg13g2_decap_4 FILLER_63_2250 ();
 sg13g2_fill_1 FILLER_63_2254 ();
 sg13g2_fill_1 FILLER_63_2291 ();
 sg13g2_fill_1 FILLER_63_2297 ();
 sg13g2_fill_1 FILLER_63_2302 ();
 sg13g2_fill_2 FILLER_63_2338 ();
 sg13g2_decap_8 FILLER_63_2346 ();
 sg13g2_decap_8 FILLER_63_2353 ();
 sg13g2_decap_8 FILLER_63_2360 ();
 sg13g2_fill_1 FILLER_63_2372 ();
 sg13g2_fill_2 FILLER_63_2408 ();
 sg13g2_decap_4 FILLER_63_2430 ();
 sg13g2_fill_2 FILLER_63_2434 ();
 sg13g2_decap_8 FILLER_63_2472 ();
 sg13g2_decap_8 FILLER_63_2479 ();
 sg13g2_fill_1 FILLER_63_2486 ();
 sg13g2_decap_8 FILLER_63_2493 ();
 sg13g2_decap_4 FILLER_63_2500 ();
 sg13g2_fill_1 FILLER_63_2539 ();
 sg13g2_decap_8 FILLER_63_2614 ();
 sg13g2_decap_8 FILLER_63_2621 ();
 sg13g2_decap_8 FILLER_63_2628 ();
 sg13g2_decap_8 FILLER_63_2635 ();
 sg13g2_decap_8 FILLER_63_2642 ();
 sg13g2_decap_8 FILLER_63_2649 ();
 sg13g2_decap_8 FILLER_63_2656 ();
 sg13g2_decap_8 FILLER_63_2663 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_fill_2 FILLER_64_14 ();
 sg13g2_fill_1 FILLER_64_16 ();
 sg13g2_fill_1 FILLER_64_21 ();
 sg13g2_fill_1 FILLER_64_31 ();
 sg13g2_fill_1 FILLER_64_37 ();
 sg13g2_fill_1 FILLER_64_44 ();
 sg13g2_fill_2 FILLER_64_51 ();
 sg13g2_fill_1 FILLER_64_58 ();
 sg13g2_fill_2 FILLER_64_64 ();
 sg13g2_fill_1 FILLER_64_75 ();
 sg13g2_fill_1 FILLER_64_80 ();
 sg13g2_fill_1 FILLER_64_85 ();
 sg13g2_fill_1 FILLER_64_96 ();
 sg13g2_fill_2 FILLER_64_108 ();
 sg13g2_fill_1 FILLER_64_110 ();
 sg13g2_fill_2 FILLER_64_141 ();
 sg13g2_fill_1 FILLER_64_147 ();
 sg13g2_fill_2 FILLER_64_168 ();
 sg13g2_fill_2 FILLER_64_174 ();
 sg13g2_fill_1 FILLER_64_176 ();
 sg13g2_fill_1 FILLER_64_191 ();
 sg13g2_fill_2 FILLER_64_207 ();
 sg13g2_decap_8 FILLER_64_227 ();
 sg13g2_decap_8 FILLER_64_234 ();
 sg13g2_decap_8 FILLER_64_241 ();
 sg13g2_decap_8 FILLER_64_248 ();
 sg13g2_decap_8 FILLER_64_255 ();
 sg13g2_decap_8 FILLER_64_262 ();
 sg13g2_decap_8 FILLER_64_269 ();
 sg13g2_decap_8 FILLER_64_276 ();
 sg13g2_decap_8 FILLER_64_323 ();
 sg13g2_decap_4 FILLER_64_330 ();
 sg13g2_fill_1 FILLER_64_334 ();
 sg13g2_decap_8 FILLER_64_379 ();
 sg13g2_decap_4 FILLER_64_386 ();
 sg13g2_fill_2 FILLER_64_390 ();
 sg13g2_fill_2 FILLER_64_419 ();
 sg13g2_fill_2 FILLER_64_428 ();
 sg13g2_decap_8 FILLER_64_435 ();
 sg13g2_decap_8 FILLER_64_442 ();
 sg13g2_decap_8 FILLER_64_449 ();
 sg13g2_decap_8 FILLER_64_456 ();
 sg13g2_decap_8 FILLER_64_463 ();
 sg13g2_fill_2 FILLER_64_470 ();
 sg13g2_decap_8 FILLER_64_485 ();
 sg13g2_fill_2 FILLER_64_492 ();
 sg13g2_fill_1 FILLER_64_494 ();
 sg13g2_fill_2 FILLER_64_499 ();
 sg13g2_decap_8 FILLER_64_506 ();
 sg13g2_decap_8 FILLER_64_513 ();
 sg13g2_fill_2 FILLER_64_520 ();
 sg13g2_decap_8 FILLER_64_526 ();
 sg13g2_decap_8 FILLER_64_533 ();
 sg13g2_decap_8 FILLER_64_540 ();
 sg13g2_decap_8 FILLER_64_547 ();
 sg13g2_fill_1 FILLER_64_564 ();
 sg13g2_fill_2 FILLER_64_573 ();
 sg13g2_decap_8 FILLER_64_580 ();
 sg13g2_decap_4 FILLER_64_587 ();
 sg13g2_fill_2 FILLER_64_591 ();
 sg13g2_fill_1 FILLER_64_628 ();
 sg13g2_decap_8 FILLER_64_638 ();
 sg13g2_decap_8 FILLER_64_645 ();
 sg13g2_decap_4 FILLER_64_652 ();
 sg13g2_fill_1 FILLER_64_656 ();
 sg13g2_decap_8 FILLER_64_662 ();
 sg13g2_decap_8 FILLER_64_669 ();
 sg13g2_decap_4 FILLER_64_676 ();
 sg13g2_fill_1 FILLER_64_680 ();
 sg13g2_decap_8 FILLER_64_701 ();
 sg13g2_decap_8 FILLER_64_708 ();
 sg13g2_decap_8 FILLER_64_720 ();
 sg13g2_decap_4 FILLER_64_727 ();
 sg13g2_decap_8 FILLER_64_757 ();
 sg13g2_decap_8 FILLER_64_764 ();
 sg13g2_fill_2 FILLER_64_771 ();
 sg13g2_decap_8 FILLER_64_776 ();
 sg13g2_decap_4 FILLER_64_783 ();
 sg13g2_fill_1 FILLER_64_787 ();
 sg13g2_fill_1 FILLER_64_812 ();
 sg13g2_fill_1 FILLER_64_834 ();
 sg13g2_fill_1 FILLER_64_864 ();
 sg13g2_fill_1 FILLER_64_873 ();
 sg13g2_decap_4 FILLER_64_904 ();
 sg13g2_fill_1 FILLER_64_908 ();
 sg13g2_fill_1 FILLER_64_972 ();
 sg13g2_fill_1 FILLER_64_1013 ();
 sg13g2_decap_4 FILLER_64_1020 ();
 sg13g2_fill_1 FILLER_64_1030 ();
 sg13g2_fill_1 FILLER_64_1059 ();
 sg13g2_fill_2 FILLER_64_1066 ();
 sg13g2_fill_2 FILLER_64_1102 ();
 sg13g2_fill_1 FILLER_64_1104 ();
 sg13g2_decap_8 FILLER_64_1111 ();
 sg13g2_fill_2 FILLER_64_1118 ();
 sg13g2_fill_2 FILLER_64_1125 ();
 sg13g2_fill_1 FILLER_64_1127 ();
 sg13g2_decap_8 FILLER_64_1141 ();
 sg13g2_fill_2 FILLER_64_1148 ();
 sg13g2_fill_1 FILLER_64_1150 ();
 sg13g2_fill_1 FILLER_64_1195 ();
 sg13g2_decap_8 FILLER_64_1233 ();
 sg13g2_fill_2 FILLER_64_1240 ();
 sg13g2_fill_1 FILLER_64_1242 ();
 sg13g2_fill_2 FILLER_64_1255 ();
 sg13g2_fill_2 FILLER_64_1380 ();
 sg13g2_fill_2 FILLER_64_1394 ();
 sg13g2_decap_4 FILLER_64_1457 ();
 sg13g2_decap_4 FILLER_64_1488 ();
 sg13g2_fill_2 FILLER_64_1492 ();
 sg13g2_fill_1 FILLER_64_1503 ();
 sg13g2_decap_8 FILLER_64_1510 ();
 sg13g2_decap_4 FILLER_64_1517 ();
 sg13g2_fill_1 FILLER_64_1521 ();
 sg13g2_fill_2 FILLER_64_1527 ();
 sg13g2_fill_1 FILLER_64_1533 ();
 sg13g2_decap_8 FILLER_64_1539 ();
 sg13g2_decap_8 FILLER_64_1546 ();
 sg13g2_fill_1 FILLER_64_1553 ();
 sg13g2_fill_1 FILLER_64_1562 ();
 sg13g2_fill_1 FILLER_64_1569 ();
 sg13g2_decap_4 FILLER_64_1575 ();
 sg13g2_fill_2 FILLER_64_1592 ();
 sg13g2_decap_4 FILLER_64_1599 ();
 sg13g2_decap_4 FILLER_64_1608 ();
 sg13g2_fill_1 FILLER_64_1664 ();
 sg13g2_decap_8 FILLER_64_1674 ();
 sg13g2_fill_2 FILLER_64_1681 ();
 sg13g2_decap_4 FILLER_64_1719 ();
 sg13g2_fill_2 FILLER_64_1723 ();
 sg13g2_decap_4 FILLER_64_1737 ();
 sg13g2_fill_1 FILLER_64_1741 ();
 sg13g2_fill_2 FILLER_64_1755 ();
 sg13g2_fill_2 FILLER_64_1814 ();
 sg13g2_decap_4 FILLER_64_1849 ();
 sg13g2_fill_1 FILLER_64_1853 ();
 sg13g2_decap_8 FILLER_64_1858 ();
 sg13g2_fill_1 FILLER_64_1865 ();
 sg13g2_decap_8 FILLER_64_1871 ();
 sg13g2_fill_1 FILLER_64_1878 ();
 sg13g2_fill_2 FILLER_64_1883 ();
 sg13g2_decap_8 FILLER_64_1896 ();
 sg13g2_decap_8 FILLER_64_1903 ();
 sg13g2_decap_8 FILLER_64_1910 ();
 sg13g2_fill_2 FILLER_64_1917 ();
 sg13g2_fill_2 FILLER_64_1936 ();
 sg13g2_fill_1 FILLER_64_1983 ();
 sg13g2_decap_4 FILLER_64_1988 ();
 sg13g2_decap_8 FILLER_64_1996 ();
 sg13g2_decap_4 FILLER_64_2003 ();
 sg13g2_fill_1 FILLER_64_2007 ();
 sg13g2_fill_2 FILLER_64_2016 ();
 sg13g2_fill_1 FILLER_64_2018 ();
 sg13g2_decap_4 FILLER_64_2048 ();
 sg13g2_fill_2 FILLER_64_2052 ();
 sg13g2_decap_4 FILLER_64_2063 ();
 sg13g2_fill_1 FILLER_64_2067 ();
 sg13g2_decap_8 FILLER_64_2099 ();
 sg13g2_fill_2 FILLER_64_2137 ();
 sg13g2_decap_8 FILLER_64_2142 ();
 sg13g2_fill_2 FILLER_64_2149 ();
 sg13g2_fill_1 FILLER_64_2151 ();
 sg13g2_decap_8 FILLER_64_2182 ();
 sg13g2_fill_2 FILLER_64_2189 ();
 sg13g2_fill_1 FILLER_64_2196 ();
 sg13g2_decap_4 FILLER_64_2201 ();
 sg13g2_fill_2 FILLER_64_2205 ();
 sg13g2_decap_8 FILLER_64_2210 ();
 sg13g2_fill_2 FILLER_64_2217 ();
 sg13g2_decap_4 FILLER_64_2242 ();
 sg13g2_fill_1 FILLER_64_2258 ();
 sg13g2_decap_4 FILLER_64_2290 ();
 sg13g2_fill_2 FILLER_64_2294 ();
 sg13g2_decap_4 FILLER_64_2327 ();
 sg13g2_fill_1 FILLER_64_2331 ();
 sg13g2_decap_8 FILLER_64_2339 ();
 sg13g2_decap_8 FILLER_64_2346 ();
 sg13g2_fill_1 FILLER_64_2353 ();
 sg13g2_decap_4 FILLER_64_2366 ();
 sg13g2_fill_2 FILLER_64_2370 ();
 sg13g2_decap_4 FILLER_64_2376 ();
 sg13g2_fill_2 FILLER_64_2386 ();
 sg13g2_fill_1 FILLER_64_2388 ();
 sg13g2_decap_8 FILLER_64_2402 ();
 sg13g2_fill_2 FILLER_64_2409 ();
 sg13g2_fill_1 FILLER_64_2411 ();
 sg13g2_decap_4 FILLER_64_2424 ();
 sg13g2_fill_1 FILLER_64_2428 ();
 sg13g2_decap_8 FILLER_64_2439 ();
 sg13g2_decap_8 FILLER_64_2446 ();
 sg13g2_decap_8 FILLER_64_2453 ();
 sg13g2_fill_2 FILLER_64_2470 ();
 sg13g2_decap_4 FILLER_64_2493 ();
 sg13g2_decap_8 FILLER_64_2523 ();
 sg13g2_decap_8 FILLER_64_2530 ();
 sg13g2_decap_8 FILLER_64_2537 ();
 sg13g2_decap_8 FILLER_64_2544 ();
 sg13g2_fill_2 FILLER_64_2551 ();
 sg13g2_fill_1 FILLER_64_2558 ();
 sg13g2_decap_8 FILLER_64_2563 ();
 sg13g2_fill_1 FILLER_64_2576 ();
 sg13g2_decap_8 FILLER_64_2582 ();
 sg13g2_decap_4 FILLER_64_2589 ();
 sg13g2_fill_1 FILLER_64_2593 ();
 sg13g2_decap_8 FILLER_64_2620 ();
 sg13g2_decap_8 FILLER_64_2627 ();
 sg13g2_decap_8 FILLER_64_2634 ();
 sg13g2_decap_8 FILLER_64_2641 ();
 sg13g2_decap_8 FILLER_64_2648 ();
 sg13g2_decap_8 FILLER_64_2655 ();
 sg13g2_decap_8 FILLER_64_2662 ();
 sg13g2_fill_1 FILLER_64_2669 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_11 ();
 sg13g2_fill_2 FILLER_65_25 ();
 sg13g2_fill_1 FILLER_65_34 ();
 sg13g2_decap_8 FILLER_65_54 ();
 sg13g2_fill_2 FILLER_65_69 ();
 sg13g2_fill_2 FILLER_65_75 ();
 sg13g2_fill_1 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_99 ();
 sg13g2_fill_1 FILLER_65_110 ();
 sg13g2_fill_1 FILLER_65_116 ();
 sg13g2_fill_1 FILLER_65_122 ();
 sg13g2_fill_2 FILLER_65_148 ();
 sg13g2_fill_1 FILLER_65_155 ();
 sg13g2_fill_1 FILLER_65_161 ();
 sg13g2_fill_1 FILLER_65_168 ();
 sg13g2_fill_1 FILLER_65_174 ();
 sg13g2_fill_2 FILLER_65_181 ();
 sg13g2_fill_2 FILLER_65_187 ();
 sg13g2_fill_2 FILLER_65_197 ();
 sg13g2_fill_1 FILLER_65_199 ();
 sg13g2_fill_2 FILLER_65_205 ();
 sg13g2_fill_2 FILLER_65_211 ();
 sg13g2_fill_1 FILLER_65_213 ();
 sg13g2_fill_2 FILLER_65_219 ();
 sg13g2_fill_1 FILLER_65_221 ();
 sg13g2_fill_2 FILLER_65_226 ();
 sg13g2_decap_8 FILLER_65_233 ();
 sg13g2_decap_8 FILLER_65_240 ();
 sg13g2_decap_4 FILLER_65_247 ();
 sg13g2_fill_1 FILLER_65_251 ();
 sg13g2_fill_1 FILLER_65_308 ();
 sg13g2_decap_8 FILLER_65_317 ();
 sg13g2_decap_8 FILLER_65_324 ();
 sg13g2_decap_4 FILLER_65_331 ();
 sg13g2_fill_2 FILLER_65_335 ();
 sg13g2_fill_1 FILLER_65_392 ();
 sg13g2_decap_4 FILLER_65_398 ();
 sg13g2_fill_1 FILLER_65_402 ();
 sg13g2_decap_4 FILLER_65_411 ();
 sg13g2_fill_2 FILLER_65_415 ();
 sg13g2_fill_2 FILLER_65_421 ();
 sg13g2_fill_1 FILLER_65_426 ();
 sg13g2_decap_8 FILLER_65_450 ();
 sg13g2_decap_8 FILLER_65_457 ();
 sg13g2_fill_1 FILLER_65_464 ();
 sg13g2_fill_1 FILLER_65_470 ();
 sg13g2_fill_1 FILLER_65_475 ();
 sg13g2_decap_4 FILLER_65_489 ();
 sg13g2_decap_4 FILLER_65_517 ();
 sg13g2_fill_1 FILLER_65_526 ();
 sg13g2_decap_4 FILLER_65_539 ();
 sg13g2_fill_2 FILLER_65_543 ();
 sg13g2_decap_8 FILLER_65_584 ();
 sg13g2_decap_8 FILLER_65_591 ();
 sg13g2_fill_2 FILLER_65_598 ();
 sg13g2_fill_1 FILLER_65_600 ();
 sg13g2_fill_1 FILLER_65_640 ();
 sg13g2_fill_2 FILLER_65_646 ();
 sg13g2_decap_4 FILLER_65_657 ();
 sg13g2_fill_1 FILLER_65_661 ();
 sg13g2_fill_1 FILLER_65_667 ();
 sg13g2_decap_8 FILLER_65_673 ();
 sg13g2_fill_2 FILLER_65_680 ();
 sg13g2_decap_8 FILLER_65_685 ();
 sg13g2_decap_8 FILLER_65_692 ();
 sg13g2_decap_8 FILLER_65_699 ();
 sg13g2_fill_2 FILLER_65_706 ();
 sg13g2_decap_8 FILLER_65_716 ();
 sg13g2_decap_8 FILLER_65_723 ();
 sg13g2_decap_8 FILLER_65_730 ();
 sg13g2_fill_2 FILLER_65_737 ();
 sg13g2_fill_1 FILLER_65_739 ();
 sg13g2_fill_2 FILLER_65_756 ();
 sg13g2_decap_8 FILLER_65_763 ();
 sg13g2_decap_8 FILLER_65_770 ();
 sg13g2_decap_4 FILLER_65_777 ();
 sg13g2_decap_4 FILLER_65_785 ();
 sg13g2_decap_4 FILLER_65_794 ();
 sg13g2_decap_8 FILLER_65_802 ();
 sg13g2_decap_4 FILLER_65_809 ();
 sg13g2_fill_1 FILLER_65_813 ();
 sg13g2_fill_2 FILLER_65_832 ();
 sg13g2_decap_8 FILLER_65_837 ();
 sg13g2_decap_4 FILLER_65_848 ();
 sg13g2_fill_1 FILLER_65_852 ();
 sg13g2_decap_4 FILLER_65_857 ();
 sg13g2_fill_1 FILLER_65_866 ();
 sg13g2_decap_8 FILLER_65_897 ();
 sg13g2_fill_2 FILLER_65_904 ();
 sg13g2_fill_2 FILLER_65_927 ();
 sg13g2_fill_1 FILLER_65_929 ();
 sg13g2_fill_2 FILLER_65_938 ();
 sg13g2_fill_1 FILLER_65_940 ();
 sg13g2_fill_2 FILLER_65_971 ();
 sg13g2_fill_2 FILLER_65_999 ();
 sg13g2_fill_1 FILLER_65_1022 ();
 sg13g2_fill_1 FILLER_65_1049 ();
 sg13g2_decap_4 FILLER_65_1056 ();
 sg13g2_fill_1 FILLER_65_1065 ();
 sg13g2_fill_2 FILLER_65_1072 ();
 sg13g2_decap_4 FILLER_65_1083 ();
 sg13g2_fill_2 FILLER_65_1091 ();
 sg13g2_decap_4 FILLER_65_1108 ();
 sg13g2_fill_1 FILLER_65_1112 ();
 sg13g2_decap_8 FILLER_65_1147 ();
 sg13g2_decap_4 FILLER_65_1154 ();
 sg13g2_fill_1 FILLER_65_1158 ();
 sg13g2_fill_1 FILLER_65_1188 ();
 sg13g2_decap_4 FILLER_65_1221 ();
 sg13g2_fill_2 FILLER_65_1225 ();
 sg13g2_fill_1 FILLER_65_1245 ();
 sg13g2_fill_2 FILLER_65_1278 ();
 sg13g2_fill_2 FILLER_65_1285 ();
 sg13g2_fill_1 FILLER_65_1328 ();
 sg13g2_fill_1 FILLER_65_1332 ();
 sg13g2_fill_2 FILLER_65_1343 ();
 sg13g2_fill_1 FILLER_65_1345 ();
 sg13g2_decap_4 FILLER_65_1355 ();
 sg13g2_fill_1 FILLER_65_1359 ();
 sg13g2_fill_1 FILLER_65_1365 ();
 sg13g2_fill_2 FILLER_65_1370 ();
 sg13g2_fill_1 FILLER_65_1378 ();
 sg13g2_fill_1 FILLER_65_1385 ();
 sg13g2_decap_8 FILLER_65_1391 ();
 sg13g2_fill_2 FILLER_65_1404 ();
 sg13g2_fill_2 FILLER_65_1416 ();
 sg13g2_fill_1 FILLER_65_1450 ();
 sg13g2_fill_1 FILLER_65_1493 ();
 sg13g2_fill_2 FILLER_65_1498 ();
 sg13g2_fill_1 FILLER_65_1500 ();
 sg13g2_decap_4 FILLER_65_1509 ();
 sg13g2_decap_4 FILLER_65_1525 ();
 sg13g2_fill_1 FILLER_65_1534 ();
 sg13g2_decap_4 FILLER_65_1552 ();
 sg13g2_fill_1 FILLER_65_1556 ();
 sg13g2_decap_8 FILLER_65_1562 ();
 sg13g2_decap_8 FILLER_65_1569 ();
 sg13g2_fill_1 FILLER_65_1576 ();
 sg13g2_fill_2 FILLER_65_1590 ();
 sg13g2_fill_1 FILLER_65_1592 ();
 sg13g2_decap_4 FILLER_65_1611 ();
 sg13g2_fill_1 FILLER_65_1615 ();
 sg13g2_decap_8 FILLER_65_1629 ();
 sg13g2_decap_8 FILLER_65_1636 ();
 sg13g2_decap_8 FILLER_65_1643 ();
 sg13g2_decap_8 FILLER_65_1650 ();
 sg13g2_fill_1 FILLER_65_1657 ();
 sg13g2_decap_4 FILLER_65_1675 ();
 sg13g2_fill_1 FILLER_65_1679 ();
 sg13g2_decap_8 FILLER_65_1706 ();
 sg13g2_decap_8 FILLER_65_1713 ();
 sg13g2_decap_8 FILLER_65_1720 ();
 sg13g2_decap_8 FILLER_65_1727 ();
 sg13g2_decap_8 FILLER_65_1789 ();
 sg13g2_decap_8 FILLER_65_1796 ();
 sg13g2_decap_8 FILLER_65_1803 ();
 sg13g2_decap_8 FILLER_65_1810 ();
 sg13g2_decap_4 FILLER_65_1817 ();
 sg13g2_fill_2 FILLER_65_1835 ();
 sg13g2_decap_8 FILLER_65_1869 ();
 sg13g2_decap_8 FILLER_65_1876 ();
 sg13g2_fill_2 FILLER_65_1891 ();
 sg13g2_fill_1 FILLER_65_1928 ();
 sg13g2_fill_1 FILLER_65_1932 ();
 sg13g2_fill_1 FILLER_65_1937 ();
 sg13g2_decap_4 FILLER_65_1941 ();
 sg13g2_fill_1 FILLER_65_1950 ();
 sg13g2_fill_2 FILLER_65_1955 ();
 sg13g2_decap_8 FILLER_65_1994 ();
 sg13g2_decap_8 FILLER_65_2001 ();
 sg13g2_decap_8 FILLER_65_2022 ();
 sg13g2_fill_1 FILLER_65_2029 ();
 sg13g2_decap_4 FILLER_65_2035 ();
 sg13g2_fill_1 FILLER_65_2039 ();
 sg13g2_decap_8 FILLER_65_2053 ();
 sg13g2_decap_8 FILLER_65_2060 ();
 sg13g2_decap_8 FILLER_65_2067 ();
 sg13g2_fill_1 FILLER_65_2074 ();
 sg13g2_fill_2 FILLER_65_2101 ();
 sg13g2_decap_4 FILLER_65_2107 ();
 sg13g2_fill_2 FILLER_65_2137 ();
 sg13g2_decap_4 FILLER_65_2145 ();
 sg13g2_fill_2 FILLER_65_2175 ();
 sg13g2_fill_1 FILLER_65_2177 ();
 sg13g2_decap_8 FILLER_65_2191 ();
 sg13g2_fill_1 FILLER_65_2198 ();
 sg13g2_decap_4 FILLER_65_2211 ();
 sg13g2_decap_8 FILLER_65_2270 ();
 sg13g2_decap_8 FILLER_65_2277 ();
 sg13g2_decap_8 FILLER_65_2289 ();
 sg13g2_decap_8 FILLER_65_2296 ();
 sg13g2_fill_2 FILLER_65_2312 ();
 sg13g2_decap_8 FILLER_65_2345 ();
 sg13g2_decap_8 FILLER_65_2352 ();
 sg13g2_decap_8 FILLER_65_2359 ();
 sg13g2_decap_4 FILLER_65_2366 ();
 sg13g2_fill_1 FILLER_65_2370 ();
 sg13g2_decap_8 FILLER_65_2375 ();
 sg13g2_decap_8 FILLER_65_2382 ();
 sg13g2_decap_8 FILLER_65_2389 ();
 sg13g2_decap_8 FILLER_65_2396 ();
 sg13g2_decap_8 FILLER_65_2403 ();
 sg13g2_decap_8 FILLER_65_2410 ();
 sg13g2_decap_8 FILLER_65_2417 ();
 sg13g2_fill_1 FILLER_65_2424 ();
 sg13g2_fill_2 FILLER_65_2451 ();
 sg13g2_decap_4 FILLER_65_2465 ();
 sg13g2_decap_8 FILLER_65_2507 ();
 sg13g2_decap_8 FILLER_65_2514 ();
 sg13g2_decap_4 FILLER_65_2521 ();
 sg13g2_fill_1 FILLER_65_2525 ();
 sg13g2_decap_4 FILLER_65_2532 ();
 sg13g2_fill_1 FILLER_65_2536 ();
 sg13g2_decap_8 FILLER_65_2542 ();
 sg13g2_decap_4 FILLER_65_2549 ();
 sg13g2_decap_8 FILLER_65_2558 ();
 sg13g2_decap_8 FILLER_65_2565 ();
 sg13g2_decap_4 FILLER_65_2572 ();
 sg13g2_fill_2 FILLER_65_2576 ();
 sg13g2_fill_2 FILLER_65_2613 ();
 sg13g2_fill_1 FILLER_65_2615 ();
 sg13g2_decap_8 FILLER_65_2646 ();
 sg13g2_decap_8 FILLER_65_2653 ();
 sg13g2_decap_8 FILLER_65_2660 ();
 sg13g2_fill_2 FILLER_65_2667 ();
 sg13g2_fill_1 FILLER_65_2669 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_fill_2 FILLER_66_14 ();
 sg13g2_fill_1 FILLER_66_16 ();
 sg13g2_fill_2 FILLER_66_47 ();
 sg13g2_fill_1 FILLER_66_49 ();
 sg13g2_fill_2 FILLER_66_54 ();
 sg13g2_fill_1 FILLER_66_56 ();
 sg13g2_fill_2 FILLER_66_62 ();
 sg13g2_fill_1 FILLER_66_64 ();
 sg13g2_fill_2 FILLER_66_71 ();
 sg13g2_fill_1 FILLER_66_73 ();
 sg13g2_fill_2 FILLER_66_83 ();
 sg13g2_fill_1 FILLER_66_85 ();
 sg13g2_fill_1 FILLER_66_101 ();
 sg13g2_decap_4 FILLER_66_119 ();
 sg13g2_fill_2 FILLER_66_123 ();
 sg13g2_fill_2 FILLER_66_130 ();
 sg13g2_decap_4 FILLER_66_139 ();
 sg13g2_decap_4 FILLER_66_151 ();
 sg13g2_fill_2 FILLER_66_162 ();
 sg13g2_fill_1 FILLER_66_164 ();
 sg13g2_fill_1 FILLER_66_169 ();
 sg13g2_fill_1 FILLER_66_174 ();
 sg13g2_fill_1 FILLER_66_179 ();
 sg13g2_fill_1 FILLER_66_185 ();
 sg13g2_fill_1 FILLER_66_192 ();
 sg13g2_fill_1 FILLER_66_197 ();
 sg13g2_fill_1 FILLER_66_203 ();
 sg13g2_fill_1 FILLER_66_209 ();
 sg13g2_fill_1 FILLER_66_216 ();
 sg13g2_fill_1 FILLER_66_222 ();
 sg13g2_fill_2 FILLER_66_228 ();
 sg13g2_decap_8 FILLER_66_235 ();
 sg13g2_decap_8 FILLER_66_242 ();
 sg13g2_fill_1 FILLER_66_249 ();
 sg13g2_fill_2 FILLER_66_281 ();
 sg13g2_decap_8 FILLER_66_337 ();
 sg13g2_fill_2 FILLER_66_344 ();
 sg13g2_fill_2 FILLER_66_362 ();
 sg13g2_fill_1 FILLER_66_364 ();
 sg13g2_decap_4 FILLER_66_414 ();
 sg13g2_decap_8 FILLER_66_444 ();
 sg13g2_decap_8 FILLER_66_451 ();
 sg13g2_decap_8 FILLER_66_458 ();
 sg13g2_decap_8 FILLER_66_465 ();
 sg13g2_fill_1 FILLER_66_493 ();
 sg13g2_fill_1 FILLER_66_499 ();
 sg13g2_fill_2 FILLER_66_521 ();
 sg13g2_decap_8 FILLER_66_563 ();
 sg13g2_fill_1 FILLER_66_570 ();
 sg13g2_decap_8 FILLER_66_581 ();
 sg13g2_decap_4 FILLER_66_588 ();
 sg13g2_fill_1 FILLER_66_592 ();
 sg13g2_fill_2 FILLER_66_601 ();
 sg13g2_fill_1 FILLER_66_603 ();
 sg13g2_fill_1 FILLER_66_630 ();
 sg13g2_decap_8 FILLER_66_640 ();
 sg13g2_fill_2 FILLER_66_669 ();
 sg13g2_fill_1 FILLER_66_671 ();
 sg13g2_fill_1 FILLER_66_687 ();
 sg13g2_decap_4 FILLER_66_696 ();
 sg13g2_fill_1 FILLER_66_714 ();
 sg13g2_decap_4 FILLER_66_739 ();
 sg13g2_decap_8 FILLER_66_778 ();
 sg13g2_decap_8 FILLER_66_785 ();
 sg13g2_fill_2 FILLER_66_792 ();
 sg13g2_fill_2 FILLER_66_820 ();
 sg13g2_fill_1 FILLER_66_858 ();
 sg13g2_decap_4 FILLER_66_863 ();
 sg13g2_fill_1 FILLER_66_867 ();
 sg13g2_fill_2 FILLER_66_882 ();
 sg13g2_decap_4 FILLER_66_910 ();
 sg13g2_decap_8 FILLER_66_940 ();
 sg13g2_decap_8 FILLER_66_947 ();
 sg13g2_fill_2 FILLER_66_954 ();
 sg13g2_fill_1 FILLER_66_956 ();
 sg13g2_decap_4 FILLER_66_962 ();
 sg13g2_fill_1 FILLER_66_966 ();
 sg13g2_fill_1 FILLER_66_975 ();
 sg13g2_fill_2 FILLER_66_1025 ();
 sg13g2_decap_4 FILLER_66_1062 ();
 sg13g2_fill_2 FILLER_66_1066 ();
 sg13g2_fill_1 FILLER_66_1074 ();
 sg13g2_fill_2 FILLER_66_1080 ();
 sg13g2_fill_1 FILLER_66_1082 ();
 sg13g2_decap_8 FILLER_66_1091 ();
 sg13g2_decap_4 FILLER_66_1114 ();
 sg13g2_fill_1 FILLER_66_1118 ();
 sg13g2_decap_4 FILLER_66_1123 ();
 sg13g2_fill_1 FILLER_66_1127 ();
 sg13g2_fill_1 FILLER_66_1133 ();
 sg13g2_fill_2 FILLER_66_1161 ();
 sg13g2_fill_1 FILLER_66_1210 ();
 sg13g2_fill_1 FILLER_66_1234 ();
 sg13g2_fill_1 FILLER_66_1298 ();
 sg13g2_fill_2 FILLER_66_1315 ();
 sg13g2_fill_1 FILLER_66_1321 ();
 sg13g2_decap_8 FILLER_66_1340 ();
 sg13g2_decap_8 FILLER_66_1347 ();
 sg13g2_decap_8 FILLER_66_1354 ();
 sg13g2_decap_8 FILLER_66_1387 ();
 sg13g2_fill_1 FILLER_66_1394 ();
 sg13g2_fill_2 FILLER_66_1401 ();
 sg13g2_decap_8 FILLER_66_1409 ();
 sg13g2_decap_4 FILLER_66_1416 ();
 sg13g2_fill_2 FILLER_66_1420 ();
 sg13g2_fill_2 FILLER_66_1432 ();
 sg13g2_fill_1 FILLER_66_1434 ();
 sg13g2_fill_2 FILLER_66_1442 ();
 sg13g2_fill_2 FILLER_66_1455 ();
 sg13g2_fill_2 FILLER_66_1476 ();
 sg13g2_fill_1 FILLER_66_1518 ();
 sg13g2_fill_1 FILLER_66_1532 ();
 sg13g2_fill_1 FILLER_66_1537 ();
 sg13g2_fill_2 FILLER_66_1564 ();
 sg13g2_fill_1 FILLER_66_1566 ();
 sg13g2_decap_8 FILLER_66_1579 ();
 sg13g2_decap_8 FILLER_66_1586 ();
 sg13g2_decap_4 FILLER_66_1593 ();
 sg13g2_fill_1 FILLER_66_1597 ();
 sg13g2_decap_8 FILLER_66_1603 ();
 sg13g2_fill_2 FILLER_66_1610 ();
 sg13g2_decap_8 FILLER_66_1616 ();
 sg13g2_decap_4 FILLER_66_1623 ();
 sg13g2_fill_1 FILLER_66_1627 ();
 sg13g2_decap_8 FILLER_66_1633 ();
 sg13g2_decap_4 FILLER_66_1640 ();
 sg13g2_fill_1 FILLER_66_1644 ();
 sg13g2_fill_1 FILLER_66_1699 ();
 sg13g2_decap_8 FILLER_66_1704 ();
 sg13g2_decap_4 FILLER_66_1711 ();
 sg13g2_fill_1 FILLER_66_1756 ();
 sg13g2_decap_4 FILLER_66_1791 ();
 sg13g2_fill_1 FILLER_66_1826 ();
 sg13g2_fill_2 FILLER_66_1841 ();
 sg13g2_decap_8 FILLER_66_1873 ();
 sg13g2_decap_8 FILLER_66_1880 ();
 sg13g2_decap_4 FILLER_66_1887 ();
 sg13g2_decap_8 FILLER_66_1920 ();
 sg13g2_fill_2 FILLER_66_1927 ();
 sg13g2_decap_8 FILLER_66_1947 ();
 sg13g2_decap_8 FILLER_66_1954 ();
 sg13g2_fill_1 FILLER_66_1961 ();
 sg13g2_decap_8 FILLER_66_1994 ();
 sg13g2_fill_2 FILLER_66_2001 ();
 sg13g2_fill_1 FILLER_66_2003 ();
 sg13g2_fill_2 FILLER_66_2013 ();
 sg13g2_decap_8 FILLER_66_2046 ();
 sg13g2_fill_2 FILLER_66_2053 ();
 sg13g2_fill_2 FILLER_66_2080 ();
 sg13g2_fill_2 FILLER_66_2112 ();
 sg13g2_decap_8 FILLER_66_2119 ();
 sg13g2_decap_4 FILLER_66_2126 ();
 sg13g2_decap_8 FILLER_66_2134 ();
 sg13g2_fill_2 FILLER_66_2141 ();
 sg13g2_decap_8 FILLER_66_2157 ();
 sg13g2_fill_2 FILLER_66_2164 ();
 sg13g2_fill_1 FILLER_66_2166 ();
 sg13g2_decap_8 FILLER_66_2216 ();
 sg13g2_decap_8 FILLER_66_2228 ();
 sg13g2_decap_4 FILLER_66_2235 ();
 sg13g2_fill_1 FILLER_66_2239 ();
 sg13g2_fill_1 FILLER_66_2258 ();
 sg13g2_fill_2 FILLER_66_2267 ();
 sg13g2_decap_8 FILLER_66_2281 ();
 sg13g2_decap_8 FILLER_66_2288 ();
 sg13g2_decap_8 FILLER_66_2295 ();
 sg13g2_decap_4 FILLER_66_2302 ();
 sg13g2_fill_1 FILLER_66_2306 ();
 sg13g2_fill_1 FILLER_66_2339 ();
 sg13g2_decap_8 FILLER_66_2344 ();
 sg13g2_decap_8 FILLER_66_2351 ();
 sg13g2_decap_8 FILLER_66_2358 ();
 sg13g2_decap_4 FILLER_66_2365 ();
 sg13g2_fill_1 FILLER_66_2369 ();
 sg13g2_fill_1 FILLER_66_2375 ();
 sg13g2_fill_1 FILLER_66_2385 ();
 sg13g2_decap_8 FILLER_66_2421 ();
 sg13g2_decap_8 FILLER_66_2433 ();
 sg13g2_fill_1 FILLER_66_2440 ();
 sg13g2_fill_1 FILLER_66_2446 ();
 sg13g2_fill_2 FILLER_66_2451 ();
 sg13g2_fill_2 FILLER_66_2458 ();
 sg13g2_fill_1 FILLER_66_2484 ();
 sg13g2_decap_4 FILLER_66_2582 ();
 sg13g2_fill_1 FILLER_66_2586 ();
 sg13g2_fill_2 FILLER_66_2592 ();
 sg13g2_decap_8 FILLER_66_2607 ();
 sg13g2_decap_8 FILLER_66_2614 ();
 sg13g2_decap_4 FILLER_66_2621 ();
 sg13g2_fill_2 FILLER_66_2625 ();
 sg13g2_decap_8 FILLER_66_2631 ();
 sg13g2_decap_8 FILLER_66_2638 ();
 sg13g2_decap_8 FILLER_66_2645 ();
 sg13g2_decap_8 FILLER_66_2652 ();
 sg13g2_decap_8 FILLER_66_2659 ();
 sg13g2_decap_4 FILLER_66_2666 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_27 ();
 sg13g2_fill_1 FILLER_67_64 ();
 sg13g2_fill_1 FILLER_67_75 ();
 sg13g2_fill_1 FILLER_67_81 ();
 sg13g2_fill_1 FILLER_67_90 ();
 sg13g2_decap_4 FILLER_67_101 ();
 sg13g2_fill_1 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_111 ();
 sg13g2_decap_8 FILLER_67_118 ();
 sg13g2_fill_1 FILLER_67_125 ();
 sg13g2_fill_1 FILLER_67_132 ();
 sg13g2_fill_2 FILLER_67_144 ();
 sg13g2_decap_8 FILLER_67_152 ();
 sg13g2_fill_1 FILLER_67_169 ();
 sg13g2_fill_1 FILLER_67_175 ();
 sg13g2_fill_2 FILLER_67_182 ();
 sg13g2_fill_1 FILLER_67_188 ();
 sg13g2_decap_8 FILLER_67_198 ();
 sg13g2_fill_2 FILLER_67_209 ();
 sg13g2_fill_1 FILLER_67_211 ();
 sg13g2_fill_1 FILLER_67_218 ();
 sg13g2_fill_2 FILLER_67_224 ();
 sg13g2_fill_1 FILLER_67_226 ();
 sg13g2_decap_8 FILLER_67_232 ();
 sg13g2_decap_8 FILLER_67_239 ();
 sg13g2_decap_4 FILLER_67_246 ();
 sg13g2_decap_8 FILLER_67_259 ();
 sg13g2_decap_8 FILLER_67_266 ();
 sg13g2_fill_1 FILLER_67_273 ();
 sg13g2_decap_8 FILLER_67_279 ();
 sg13g2_decap_4 FILLER_67_286 ();
 sg13g2_fill_2 FILLER_67_290 ();
 sg13g2_decap_8 FILLER_67_296 ();
 sg13g2_decap_8 FILLER_67_303 ();
 sg13g2_decap_8 FILLER_67_310 ();
 sg13g2_decap_8 FILLER_67_317 ();
 sg13g2_fill_2 FILLER_67_324 ();
 sg13g2_fill_1 FILLER_67_326 ();
 sg13g2_decap_8 FILLER_67_331 ();
 sg13g2_decap_4 FILLER_67_338 ();
 sg13g2_fill_2 FILLER_67_342 ();
 sg13g2_fill_1 FILLER_67_382 ();
 sg13g2_fill_1 FILLER_67_404 ();
 sg13g2_decap_8 FILLER_67_409 ();
 sg13g2_fill_1 FILLER_67_421 ();
 sg13g2_decap_8 FILLER_67_439 ();
 sg13g2_decap_8 FILLER_67_446 ();
 sg13g2_decap_8 FILLER_67_453 ();
 sg13g2_decap_8 FILLER_67_460 ();
 sg13g2_decap_8 FILLER_67_467 ();
 sg13g2_decap_4 FILLER_67_474 ();
 sg13g2_fill_2 FILLER_67_491 ();
 sg13g2_fill_1 FILLER_67_493 ();
 sg13g2_fill_1 FILLER_67_514 ();
 sg13g2_fill_1 FILLER_67_523 ();
 sg13g2_decap_8 FILLER_67_533 ();
 sg13g2_decap_4 FILLER_67_540 ();
 sg13g2_fill_2 FILLER_67_544 ();
 sg13g2_fill_1 FILLER_67_616 ();
 sg13g2_fill_2 FILLER_67_631 ();
 sg13g2_decap_8 FILLER_67_641 ();
 sg13g2_decap_4 FILLER_67_648 ();
 sg13g2_fill_1 FILLER_67_652 ();
 sg13g2_fill_2 FILLER_67_662 ();
 sg13g2_fill_1 FILLER_67_664 ();
 sg13g2_decap_4 FILLER_67_711 ();
 sg13g2_decap_4 FILLER_67_720 ();
 sg13g2_decap_8 FILLER_67_738 ();
 sg13g2_fill_1 FILLER_67_745 ();
 sg13g2_decap_4 FILLER_67_787 ();
 sg13g2_fill_1 FILLER_67_791 ();
 sg13g2_decap_8 FILLER_67_839 ();
 sg13g2_fill_2 FILLER_67_846 ();
 sg13g2_fill_1 FILLER_67_848 ();
 sg13g2_fill_2 FILLER_67_854 ();
 sg13g2_fill_1 FILLER_67_856 ();
 sg13g2_fill_2 FILLER_67_869 ();
 sg13g2_fill_1 FILLER_67_871 ();
 sg13g2_decap_4 FILLER_67_891 ();
 sg13g2_fill_2 FILLER_67_895 ();
 sg13g2_decap_8 FILLER_67_923 ();
 sg13g2_decap_8 FILLER_67_930 ();
 sg13g2_decap_4 FILLER_67_937 ();
 sg13g2_fill_2 FILLER_67_941 ();
 sg13g2_fill_1 FILLER_67_1013 ();
 sg13g2_fill_1 FILLER_67_1017 ();
 sg13g2_fill_1 FILLER_67_1052 ();
 sg13g2_decap_8 FILLER_67_1057 ();
 sg13g2_decap_8 FILLER_67_1064 ();
 sg13g2_decap_8 FILLER_67_1071 ();
 sg13g2_decap_8 FILLER_67_1078 ();
 sg13g2_decap_4 FILLER_67_1085 ();
 sg13g2_fill_2 FILLER_67_1089 ();
 sg13g2_fill_1 FILLER_67_1096 ();
 sg13g2_fill_2 FILLER_67_1121 ();
 sg13g2_fill_1 FILLER_67_1123 ();
 sg13g2_decap_4 FILLER_67_1141 ();
 sg13g2_decap_4 FILLER_67_1156 ();
 sg13g2_fill_1 FILLER_67_1160 ();
 sg13g2_decap_8 FILLER_67_1169 ();
 sg13g2_decap_8 FILLER_67_1181 ();
 sg13g2_fill_2 FILLER_67_1225 ();
 sg13g2_fill_1 FILLER_67_1243 ();
 sg13g2_decap_4 FILLER_67_1260 ();
 sg13g2_fill_2 FILLER_67_1264 ();
 sg13g2_fill_1 FILLER_67_1277 ();
 sg13g2_fill_1 FILLER_67_1292 ();
 sg13g2_fill_2 FILLER_67_1303 ();
 sg13g2_fill_1 FILLER_67_1322 ();
 sg13g2_decap_8 FILLER_67_1352 ();
 sg13g2_decap_8 FILLER_67_1359 ();
 sg13g2_decap_8 FILLER_67_1402 ();
 sg13g2_fill_2 FILLER_67_1409 ();
 sg13g2_decap_8 FILLER_67_1429 ();
 sg13g2_fill_2 FILLER_67_1436 ();
 sg13g2_fill_1 FILLER_67_1438 ();
 sg13g2_fill_2 FILLER_67_1447 ();
 sg13g2_fill_2 FILLER_67_1483 ();
 sg13g2_decap_8 FILLER_67_1511 ();
 sg13g2_fill_2 FILLER_67_1518 ();
 sg13g2_fill_2 FILLER_67_1524 ();
 sg13g2_fill_1 FILLER_67_1526 ();
 sg13g2_decap_8 FILLER_67_1537 ();
 sg13g2_decap_8 FILLER_67_1544 ();
 sg13g2_decap_8 FILLER_67_1560 ();
 sg13g2_decap_8 FILLER_67_1573 ();
 sg13g2_decap_8 FILLER_67_1580 ();
 sg13g2_decap_8 FILLER_67_1587 ();
 sg13g2_fill_1 FILLER_67_1594 ();
 sg13g2_decap_8 FILLER_67_1625 ();
 sg13g2_decap_4 FILLER_67_1632 ();
 sg13g2_fill_2 FILLER_67_1636 ();
 sg13g2_decap_8 FILLER_67_1683 ();
 sg13g2_decap_8 FILLER_67_1690 ();
 sg13g2_decap_8 FILLER_67_1697 ();
 sg13g2_decap_8 FILLER_67_1704 ();
 sg13g2_fill_2 FILLER_67_1711 ();
 sg13g2_decap_8 FILLER_67_1748 ();
 sg13g2_decap_8 FILLER_67_1755 ();
 sg13g2_decap_8 FILLER_67_1762 ();
 sg13g2_decap_8 FILLER_67_1793 ();
 sg13g2_fill_2 FILLER_67_1800 ();
 sg13g2_fill_1 FILLER_67_1802 ();
 sg13g2_decap_4 FILLER_67_1815 ();
 sg13g2_decap_4 FILLER_67_1849 ();
 sg13g2_fill_2 FILLER_67_1857 ();
 sg13g2_fill_1 FILLER_67_1859 ();
 sg13g2_fill_2 FILLER_67_1865 ();
 sg13g2_fill_1 FILLER_67_1867 ();
 sg13g2_decap_8 FILLER_67_1872 ();
 sg13g2_fill_2 FILLER_67_1879 ();
 sg13g2_fill_1 FILLER_67_1881 ();
 sg13g2_fill_2 FILLER_67_1891 ();
 sg13g2_decap_8 FILLER_67_1896 ();
 sg13g2_decap_4 FILLER_67_1903 ();
 sg13g2_fill_1 FILLER_67_1916 ();
 sg13g2_fill_2 FILLER_67_1923 ();
 sg13g2_fill_1 FILLER_67_1925 ();
 sg13g2_decap_8 FILLER_67_1971 ();
 sg13g2_fill_2 FILLER_67_1978 ();
 sg13g2_decap_4 FILLER_67_1988 ();
 sg13g2_decap_4 FILLER_67_2019 ();
 sg13g2_decap_4 FILLER_67_2033 ();
 sg13g2_decap_8 FILLER_67_2073 ();
 sg13g2_decap_8 FILLER_67_2090 ();
 sg13g2_decap_4 FILLER_67_2103 ();
 sg13g2_fill_2 FILLER_67_2107 ();
 sg13g2_decap_8 FILLER_67_2112 ();
 sg13g2_decap_8 FILLER_67_2119 ();
 sg13g2_decap_8 FILLER_67_2126 ();
 sg13g2_fill_2 FILLER_67_2133 ();
 sg13g2_fill_1 FILLER_67_2135 ();
 sg13g2_decap_8 FILLER_67_2139 ();
 sg13g2_decap_4 FILLER_67_2146 ();
 sg13g2_fill_2 FILLER_67_2150 ();
 sg13g2_fill_1 FILLER_67_2178 ();
 sg13g2_decap_8 FILLER_67_2225 ();
 sg13g2_decap_8 FILLER_67_2232 ();
 sg13g2_fill_2 FILLER_67_2239 ();
 sg13g2_fill_1 FILLER_67_2241 ();
 sg13g2_decap_4 FILLER_67_2260 ();
 sg13g2_fill_2 FILLER_67_2312 ();
 sg13g2_fill_1 FILLER_67_2314 ();
 sg13g2_fill_1 FILLER_67_2367 ();
 sg13g2_fill_2 FILLER_67_2411 ();
 sg13g2_fill_1 FILLER_67_2413 ();
 sg13g2_fill_2 FILLER_67_2492 ();
 sg13g2_decap_8 FILLER_67_2506 ();
 sg13g2_decap_8 FILLER_67_2513 ();
 sg13g2_fill_2 FILLER_67_2545 ();
 sg13g2_fill_1 FILLER_67_2547 ();
 sg13g2_decap_8 FILLER_67_2560 ();
 sg13g2_fill_2 FILLER_67_2572 ();
 sg13g2_decap_8 FILLER_67_2613 ();
 sg13g2_decap_8 FILLER_67_2620 ();
 sg13g2_decap_8 FILLER_67_2627 ();
 sg13g2_decap_8 FILLER_67_2634 ();
 sg13g2_decap_8 FILLER_67_2641 ();
 sg13g2_decap_8 FILLER_67_2648 ();
 sg13g2_decap_8 FILLER_67_2655 ();
 sg13g2_decap_8 FILLER_67_2662 ();
 sg13g2_fill_1 FILLER_67_2669 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_16 ();
 sg13g2_fill_1 FILLER_68_49 ();
 sg13g2_fill_1 FILLER_68_60 ();
 sg13g2_fill_1 FILLER_68_81 ();
 sg13g2_fill_2 FILLER_68_87 ();
 sg13g2_fill_1 FILLER_68_107 ();
 sg13g2_fill_1 FILLER_68_112 ();
 sg13g2_fill_1 FILLER_68_118 ();
 sg13g2_fill_1 FILLER_68_126 ();
 sg13g2_decap_4 FILLER_68_135 ();
 sg13g2_fill_1 FILLER_68_144 ();
 sg13g2_fill_1 FILLER_68_192 ();
 sg13g2_fill_1 FILLER_68_198 ();
 sg13g2_fill_2 FILLER_68_228 ();
 sg13g2_decap_8 FILLER_68_234 ();
 sg13g2_decap_4 FILLER_68_241 ();
 sg13g2_decap_8 FILLER_68_249 ();
 sg13g2_decap_8 FILLER_68_256 ();
 sg13g2_decap_8 FILLER_68_263 ();
 sg13g2_decap_8 FILLER_68_270 ();
 sg13g2_fill_2 FILLER_68_277 ();
 sg13g2_fill_2 FILLER_68_284 ();
 sg13g2_decap_8 FILLER_68_312 ();
 sg13g2_decap_8 FILLER_68_319 ();
 sg13g2_decap_8 FILLER_68_326 ();
 sg13g2_decap_8 FILLER_68_333 ();
 sg13g2_decap_4 FILLER_68_345 ();
 sg13g2_fill_1 FILLER_68_352 ();
 sg13g2_fill_1 FILLER_68_384 ();
 sg13g2_fill_1 FILLER_68_411 ();
 sg13g2_fill_1 FILLER_68_417 ();
 sg13g2_fill_1 FILLER_68_433 ();
 sg13g2_decap_8 FILLER_68_439 ();
 sg13g2_decap_8 FILLER_68_446 ();
 sg13g2_decap_8 FILLER_68_488 ();
 sg13g2_fill_2 FILLER_68_495 ();
 sg13g2_fill_1 FILLER_68_515 ();
 sg13g2_fill_2 FILLER_68_522 ();
 sg13g2_decap_8 FILLER_68_529 ();
 sg13g2_decap_8 FILLER_68_536 ();
 sg13g2_decap_4 FILLER_68_543 ();
 sg13g2_decap_8 FILLER_68_556 ();
 sg13g2_decap_8 FILLER_68_563 ();
 sg13g2_decap_8 FILLER_68_570 ();
 sg13g2_fill_2 FILLER_68_577 ();
 sg13g2_decap_8 FILLER_68_583 ();
 sg13g2_decap_4 FILLER_68_590 ();
 sg13g2_fill_1 FILLER_68_594 ();
 sg13g2_fill_2 FILLER_68_622 ();
 sg13g2_fill_1 FILLER_68_631 ();
 sg13g2_decap_8 FILLER_68_642 ();
 sg13g2_decap_8 FILLER_68_649 ();
 sg13g2_fill_1 FILLER_68_656 ();
 sg13g2_fill_1 FILLER_68_660 ();
 sg13g2_fill_1 FILLER_68_669 ();
 sg13g2_decap_4 FILLER_68_697 ();
 sg13g2_fill_1 FILLER_68_701 ();
 sg13g2_fill_1 FILLER_68_706 ();
 sg13g2_fill_2 FILLER_68_717 ();
 sg13g2_fill_1 FILLER_68_719 ();
 sg13g2_decap_4 FILLER_68_756 ();
 sg13g2_fill_1 FILLER_68_760 ();
 sg13g2_decap_8 FILLER_68_764 ();
 sg13g2_decap_4 FILLER_68_771 ();
 sg13g2_fill_1 FILLER_68_775 ();
 sg13g2_decap_8 FILLER_68_781 ();
 sg13g2_decap_8 FILLER_68_788 ();
 sg13g2_fill_2 FILLER_68_795 ();
 sg13g2_fill_2 FILLER_68_809 ();
 sg13g2_fill_1 FILLER_68_811 ();
 sg13g2_fill_2 FILLER_68_825 ();
 sg13g2_fill_2 FILLER_68_832 ();
 sg13g2_fill_1 FILLER_68_834 ();
 sg13g2_decap_8 FILLER_68_861 ();
 sg13g2_fill_1 FILLER_68_868 ();
 sg13g2_decap_4 FILLER_68_877 ();
 sg13g2_decap_8 FILLER_68_885 ();
 sg13g2_decap_8 FILLER_68_892 ();
 sg13g2_decap_4 FILLER_68_909 ();
 sg13g2_fill_2 FILLER_68_913 ();
 sg13g2_decap_8 FILLER_68_923 ();
 sg13g2_decap_8 FILLER_68_930 ();
 sg13g2_decap_8 FILLER_68_937 ();
 sg13g2_decap_4 FILLER_68_944 ();
 sg13g2_fill_1 FILLER_68_948 ();
 sg13g2_decap_4 FILLER_68_953 ();
 sg13g2_fill_1 FILLER_68_992 ();
 sg13g2_fill_2 FILLER_68_1003 ();
 sg13g2_decap_8 FILLER_68_1055 ();
 sg13g2_decap_8 FILLER_68_1067 ();
 sg13g2_fill_2 FILLER_68_1080 ();
 sg13g2_fill_1 FILLER_68_1082 ();
 sg13g2_fill_2 FILLER_68_1120 ();
 sg13g2_fill_1 FILLER_68_1122 ();
 sg13g2_fill_2 FILLER_68_1129 ();
 sg13g2_fill_1 FILLER_68_1137 ();
 sg13g2_fill_2 FILLER_68_1143 ();
 sg13g2_decap_4 FILLER_68_1155 ();
 sg13g2_fill_1 FILLER_68_1190 ();
 sg13g2_decap_8 FILLER_68_1197 ();
 sg13g2_fill_1 FILLER_68_1204 ();
 sg13g2_fill_2 FILLER_68_1224 ();
 sg13g2_fill_1 FILLER_68_1253 ();
 sg13g2_fill_1 FILLER_68_1289 ();
 sg13g2_fill_1 FILLER_68_1298 ();
 sg13g2_decap_8 FILLER_68_1338 ();
 sg13g2_fill_2 FILLER_68_1345 ();
 sg13g2_fill_1 FILLER_68_1347 ();
 sg13g2_fill_2 FILLER_68_1353 ();
 sg13g2_fill_1 FILLER_68_1355 ();
 sg13g2_fill_2 FILLER_68_1361 ();
 sg13g2_fill_1 FILLER_68_1363 ();
 sg13g2_decap_8 FILLER_68_1374 ();
 sg13g2_decap_8 FILLER_68_1381 ();
 sg13g2_fill_2 FILLER_68_1388 ();
 sg13g2_fill_2 FILLER_68_1405 ();
 sg13g2_decap_4 FILLER_68_1440 ();
 sg13g2_fill_2 FILLER_68_1478 ();
 sg13g2_decap_4 FILLER_68_1492 ();
 sg13g2_fill_1 FILLER_68_1496 ();
 sg13g2_decap_8 FILLER_68_1503 ();
 sg13g2_decap_4 FILLER_68_1510 ();
 sg13g2_fill_1 FILLER_68_1514 ();
 sg13g2_decap_8 FILLER_68_1545 ();
 sg13g2_decap_4 FILLER_68_1552 ();
 sg13g2_fill_2 FILLER_68_1556 ();
 sg13g2_fill_1 FILLER_68_1577 ();
 sg13g2_decap_4 FILLER_68_1591 ();
 sg13g2_decap_4 FILLER_68_1630 ();
 sg13g2_decap_8 FILLER_68_1694 ();
 sg13g2_decap_4 FILLER_68_1701 ();
 sg13g2_fill_2 FILLER_68_1705 ();
 sg13g2_decap_8 FILLER_68_1715 ();
 sg13g2_fill_1 FILLER_68_1722 ();
 sg13g2_fill_1 FILLER_68_1728 ();
 sg13g2_fill_2 FILLER_68_1733 ();
 sg13g2_fill_1 FILLER_68_1735 ();
 sg13g2_fill_2 FILLER_68_1748 ();
 sg13g2_fill_1 FILLER_68_1789 ();
 sg13g2_decap_8 FILLER_68_1796 ();
 sg13g2_fill_2 FILLER_68_1803 ();
 sg13g2_fill_2 FILLER_68_1810 ();
 sg13g2_decap_8 FILLER_68_1821 ();
 sg13g2_decap_4 FILLER_68_1828 ();
 sg13g2_decap_4 FILLER_68_1838 ();
 sg13g2_fill_2 FILLER_68_1842 ();
 sg13g2_fill_2 FILLER_68_1874 ();
 sg13g2_fill_2 FILLER_68_1907 ();
 sg13g2_fill_1 FILLER_68_1909 ();
 sg13g2_fill_1 FILLER_68_1925 ();
 sg13g2_fill_2 FILLER_68_1960 ();
 sg13g2_decap_8 FILLER_68_1967 ();
 sg13g2_fill_1 FILLER_68_1974 ();
 sg13g2_decap_8 FILLER_68_1979 ();
 sg13g2_fill_1 FILLER_68_1986 ();
 sg13g2_decap_4 FILLER_68_2022 ();
 sg13g2_fill_1 FILLER_68_2026 ();
 sg13g2_decap_4 FILLER_68_2032 ();
 sg13g2_fill_2 FILLER_68_2044 ();
 sg13g2_fill_2 FILLER_68_2052 ();
 sg13g2_fill_1 FILLER_68_2054 ();
 sg13g2_decap_8 FILLER_68_2091 ();
 sg13g2_decap_8 FILLER_68_2098 ();
 sg13g2_decap_8 FILLER_68_2105 ();
 sg13g2_decap_8 FILLER_68_2112 ();
 sg13g2_fill_2 FILLER_68_2119 ();
 sg13g2_decap_8 FILLER_68_2125 ();
 sg13g2_fill_1 FILLER_68_2132 ();
 sg13g2_decap_8 FILLER_68_2142 ();
 sg13g2_decap_4 FILLER_68_2149 ();
 sg13g2_fill_2 FILLER_68_2153 ();
 sg13g2_decap_4 FILLER_68_2167 ();
 sg13g2_fill_1 FILLER_68_2171 ();
 sg13g2_decap_4 FILLER_68_2201 ();
 sg13g2_decap_8 FILLER_68_2209 ();
 sg13g2_decap_8 FILLER_68_2216 ();
 sg13g2_fill_2 FILLER_68_2223 ();
 sg13g2_fill_1 FILLER_68_2225 ();
 sg13g2_fill_2 FILLER_68_2262 ();
 sg13g2_decap_8 FILLER_68_2269 ();
 sg13g2_decap_8 FILLER_68_2276 ();
 sg13g2_decap_4 FILLER_68_2283 ();
 sg13g2_decap_8 FILLER_68_2290 ();
 sg13g2_decap_8 FILLER_68_2302 ();
 sg13g2_fill_2 FILLER_68_2322 ();
 sg13g2_fill_1 FILLER_68_2367 ();
 sg13g2_decap_4 FILLER_68_2382 ();
 sg13g2_decap_8 FILLER_68_2396 ();
 sg13g2_fill_1 FILLER_68_2403 ();
 sg13g2_decap_8 FILLER_68_2434 ();
 sg13g2_decap_8 FILLER_68_2441 ();
 sg13g2_fill_2 FILLER_68_2448 ();
 sg13g2_fill_1 FILLER_68_2450 ();
 sg13g2_fill_1 FILLER_68_2454 ();
 sg13g2_fill_1 FILLER_68_2478 ();
 sg13g2_decap_4 FILLER_68_2485 ();
 sg13g2_decap_4 FILLER_68_2527 ();
 sg13g2_decap_8 FILLER_68_2566 ();
 sg13g2_fill_1 FILLER_68_2573 ();
 sg13g2_fill_1 FILLER_68_2585 ();
 sg13g2_decap_8 FILLER_68_2625 ();
 sg13g2_decap_8 FILLER_68_2632 ();
 sg13g2_decap_8 FILLER_68_2639 ();
 sg13g2_decap_8 FILLER_68_2646 ();
 sg13g2_decap_8 FILLER_68_2653 ();
 sg13g2_decap_8 FILLER_68_2660 ();
 sg13g2_fill_2 FILLER_68_2667 ();
 sg13g2_fill_1 FILLER_68_2669 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_9 ();
 sg13g2_decap_4 FILLER_69_15 ();
 sg13g2_fill_2 FILLER_69_47 ();
 sg13g2_fill_1 FILLER_69_60 ();
 sg13g2_fill_1 FILLER_69_89 ();
 sg13g2_fill_1 FILLER_69_100 ();
 sg13g2_fill_1 FILLER_69_105 ();
 sg13g2_fill_1 FILLER_69_111 ();
 sg13g2_fill_1 FILLER_69_123 ();
 sg13g2_fill_1 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_143 ();
 sg13g2_decap_8 FILLER_69_150 ();
 sg13g2_fill_1 FILLER_69_185 ();
 sg13g2_fill_1 FILLER_69_191 ();
 sg13g2_fill_1 FILLER_69_217 ();
 sg13g2_decap_8 FILLER_69_223 ();
 sg13g2_fill_1 FILLER_69_230 ();
 sg13g2_decap_4 FILLER_69_261 ();
 sg13g2_fill_1 FILLER_69_265 ();
 sg13g2_fill_2 FILLER_69_270 ();
 sg13g2_fill_1 FILLER_69_272 ();
 sg13g2_decap_8 FILLER_69_316 ();
 sg13g2_decap_8 FILLER_69_323 ();
 sg13g2_fill_2 FILLER_69_330 ();
 sg13g2_fill_1 FILLER_69_332 ();
 sg13g2_fill_2 FILLER_69_338 ();
 sg13g2_fill_1 FILLER_69_340 ();
 sg13g2_decap_4 FILLER_69_346 ();
 sg13g2_fill_2 FILLER_69_361 ();
 sg13g2_fill_1 FILLER_69_371 ();
 sg13g2_decap_8 FILLER_69_377 ();
 sg13g2_decap_4 FILLER_69_384 ();
 sg13g2_decap_4 FILLER_69_395 ();
 sg13g2_fill_2 FILLER_69_413 ();
 sg13g2_fill_2 FILLER_69_427 ();
 sg13g2_fill_1 FILLER_69_429 ();
 sg13g2_decap_8 FILLER_69_435 ();
 sg13g2_decap_8 FILLER_69_442 ();
 sg13g2_decap_8 FILLER_69_449 ();
 sg13g2_fill_1 FILLER_69_456 ();
 sg13g2_decap_4 FILLER_69_499 ();
 sg13g2_fill_2 FILLER_69_503 ();
 sg13g2_decap_4 FILLER_69_515 ();
 sg13g2_decap_8 FILLER_69_542 ();
 sg13g2_decap_4 FILLER_69_579 ();
 sg13g2_fill_2 FILLER_69_583 ();
 sg13g2_decap_4 FILLER_69_589 ();
 sg13g2_fill_2 FILLER_69_593 ();
 sg13g2_fill_1 FILLER_69_602 ();
 sg13g2_fill_2 FILLER_69_612 ();
 sg13g2_fill_1 FILLER_69_614 ();
 sg13g2_decap_8 FILLER_69_623 ();
 sg13g2_decap_4 FILLER_69_630 ();
 sg13g2_fill_1 FILLER_69_634 ();
 sg13g2_decap_8 FILLER_69_665 ();
 sg13g2_decap_8 FILLER_69_672 ();
 sg13g2_fill_1 FILLER_69_679 ();
 sg13g2_decap_4 FILLER_69_685 ();
 sg13g2_decap_8 FILLER_69_694 ();
 sg13g2_decap_8 FILLER_69_701 ();
 sg13g2_fill_2 FILLER_69_708 ();
 sg13g2_fill_1 FILLER_69_710 ();
 sg13g2_decap_4 FILLER_69_720 ();
 sg13g2_fill_1 FILLER_69_738 ();
 sg13g2_fill_2 FILLER_69_744 ();
 sg13g2_decap_8 FILLER_69_785 ();
 sg13g2_decap_8 FILLER_69_792 ();
 sg13g2_decap_8 FILLER_69_799 ();
 sg13g2_decap_8 FILLER_69_806 ();
 sg13g2_fill_2 FILLER_69_813 ();
 sg13g2_fill_1 FILLER_69_815 ();
 sg13g2_fill_2 FILLER_69_820 ();
 sg13g2_fill_1 FILLER_69_822 ();
 sg13g2_decap_8 FILLER_69_853 ();
 sg13g2_fill_2 FILLER_69_898 ();
 sg13g2_fill_1 FILLER_69_900 ();
 sg13g2_decap_8 FILLER_69_931 ();
 sg13g2_fill_2 FILLER_69_938 ();
 sg13g2_decap_8 FILLER_69_955 ();
 sg13g2_fill_2 FILLER_69_962 ();
 sg13g2_fill_2 FILLER_69_1007 ();
 sg13g2_fill_1 FILLER_69_1048 ();
 sg13g2_fill_1 FILLER_69_1079 ();
 sg13g2_fill_2 FILLER_69_1099 ();
 sg13g2_fill_2 FILLER_69_1112 ();
 sg13g2_fill_1 FILLER_69_1114 ();
 sg13g2_fill_2 FILLER_69_1126 ();
 sg13g2_fill_1 FILLER_69_1165 ();
 sg13g2_decap_4 FILLER_69_1201 ();
 sg13g2_fill_2 FILLER_69_1214 ();
 sg13g2_fill_1 FILLER_69_1271 ();
 sg13g2_fill_2 FILLER_69_1282 ();
 sg13g2_fill_1 FILLER_69_1288 ();
 sg13g2_fill_2 FILLER_69_1302 ();
 sg13g2_fill_1 FILLER_69_1304 ();
 sg13g2_fill_1 FILLER_69_1329 ();
 sg13g2_decap_4 FILLER_69_1335 ();
 sg13g2_fill_2 FILLER_69_1339 ();
 sg13g2_fill_2 FILLER_69_1357 ();
 sg13g2_fill_1 FILLER_69_1359 ();
 sg13g2_fill_1 FILLER_69_1392 ();
 sg13g2_fill_2 FILLER_69_1410 ();
 sg13g2_fill_2 FILLER_69_1454 ();
 sg13g2_fill_2 FILLER_69_1469 ();
 sg13g2_fill_2 FILLER_69_1482 ();
 sg13g2_fill_2 FILLER_69_1497 ();
 sg13g2_fill_1 FILLER_69_1499 ();
 sg13g2_decap_8 FILLER_69_1535 ();
 sg13g2_decap_8 FILLER_69_1542 ();
 sg13g2_decap_4 FILLER_69_1549 ();
 sg13g2_fill_1 FILLER_69_1553 ();
 sg13g2_decap_4 FILLER_69_1558 ();
 sg13g2_fill_1 FILLER_69_1562 ();
 sg13g2_fill_2 FILLER_69_1579 ();
 sg13g2_fill_2 FILLER_69_1595 ();
 sg13g2_decap_8 FILLER_69_1672 ();
 sg13g2_decap_8 FILLER_69_1679 ();
 sg13g2_decap_4 FILLER_69_1686 ();
 sg13g2_fill_2 FILLER_69_1690 ();
 sg13g2_decap_8 FILLER_69_1702 ();
 sg13g2_decap_8 FILLER_69_1709 ();
 sg13g2_decap_8 FILLER_69_1716 ();
 sg13g2_decap_8 FILLER_69_1723 ();
 sg13g2_decap_8 FILLER_69_1730 ();
 sg13g2_decap_8 FILLER_69_1737 ();
 sg13g2_decap_8 FILLER_69_1744 ();
 sg13g2_decap_4 FILLER_69_1751 ();
 sg13g2_fill_1 FILLER_69_1773 ();
 sg13g2_decap_8 FILLER_69_1824 ();
 sg13g2_decap_8 FILLER_69_1831 ();
 sg13g2_decap_4 FILLER_69_1838 ();
 sg13g2_fill_1 FILLER_69_1842 ();
 sg13g2_fill_2 FILLER_69_1875 ();
 sg13g2_decap_4 FILLER_69_1903 ();
 sg13g2_fill_2 FILLER_69_1919 ();
 sg13g2_decap_4 FILLER_69_1951 ();
 sg13g2_fill_2 FILLER_69_1961 ();
 sg13g2_decap_4 FILLER_69_1989 ();
 sg13g2_fill_2 FILLER_69_2025 ();
 sg13g2_fill_1 FILLER_69_2027 ();
 sg13g2_fill_2 FILLER_69_2067 ();
 sg13g2_fill_1 FILLER_69_2069 ();
 sg13g2_fill_2 FILLER_69_2096 ();
 sg13g2_fill_2 FILLER_69_2102 ();
 sg13g2_fill_1 FILLER_69_2104 ();
 sg13g2_fill_1 FILLER_69_2139 ();
 sg13g2_fill_1 FILLER_69_2144 ();
 sg13g2_decap_4 FILLER_69_2181 ();
 sg13g2_decap_8 FILLER_69_2215 ();
 sg13g2_fill_2 FILLER_69_2222 ();
 sg13g2_decap_8 FILLER_69_2234 ();
 sg13g2_fill_2 FILLER_69_2241 ();
 sg13g2_fill_1 FILLER_69_2243 ();
 sg13g2_fill_2 FILLER_69_2302 ();
 sg13g2_decap_8 FILLER_69_2361 ();
 sg13g2_fill_2 FILLER_69_2374 ();
 sg13g2_fill_1 FILLER_69_2402 ();
 sg13g2_decap_8 FILLER_69_2416 ();
 sg13g2_decap_8 FILLER_69_2431 ();
 sg13g2_decap_8 FILLER_69_2438 ();
 sg13g2_fill_2 FILLER_69_2445 ();
 sg13g2_fill_1 FILLER_69_2447 ();
 sg13g2_fill_1 FILLER_69_2457 ();
 sg13g2_decap_8 FILLER_69_2485 ();
 sg13g2_decap_8 FILLER_69_2492 ();
 sg13g2_decap_8 FILLER_69_2499 ();
 sg13g2_fill_2 FILLER_69_2506 ();
 sg13g2_fill_2 FILLER_69_2513 ();
 sg13g2_fill_1 FILLER_69_2515 ();
 sg13g2_fill_1 FILLER_69_2547 ();
 sg13g2_fill_2 FILLER_69_2574 ();
 sg13g2_fill_1 FILLER_69_2602 ();
 sg13g2_decap_8 FILLER_69_2608 ();
 sg13g2_decap_4 FILLER_69_2615 ();
 sg13g2_fill_1 FILLER_69_2619 ();
 sg13g2_decap_8 FILLER_69_2650 ();
 sg13g2_decap_8 FILLER_69_2657 ();
 sg13g2_decap_4 FILLER_69_2664 ();
 sg13g2_fill_2 FILLER_69_2668 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_7 ();
 sg13g2_fill_1 FILLER_70_9 ();
 sg13g2_decap_8 FILLER_70_62 ();
 sg13g2_fill_2 FILLER_70_69 ();
 sg13g2_decap_8 FILLER_70_75 ();
 sg13g2_decap_8 FILLER_70_82 ();
 sg13g2_decap_8 FILLER_70_89 ();
 sg13g2_decap_4 FILLER_70_96 ();
 sg13g2_fill_1 FILLER_70_114 ();
 sg13g2_fill_1 FILLER_70_119 ();
 sg13g2_fill_1 FILLER_70_132 ();
 sg13g2_fill_2 FILLER_70_153 ();
 sg13g2_fill_1 FILLER_70_155 ();
 sg13g2_fill_2 FILLER_70_194 ();
 sg13g2_decap_4 FILLER_70_215 ();
 sg13g2_decap_8 FILLER_70_222 ();
 sg13g2_decap_4 FILLER_70_229 ();
 sg13g2_fill_2 FILLER_70_233 ();
 sg13g2_fill_2 FILLER_70_240 ();
 sg13g2_decap_4 FILLER_70_246 ();
 sg13g2_decap_4 FILLER_70_254 ();
 sg13g2_fill_2 FILLER_70_284 ();
 sg13g2_fill_1 FILLER_70_286 ();
 sg13g2_decap_4 FILLER_70_312 ();
 sg13g2_decap_8 FILLER_70_325 ();
 sg13g2_decap_4 FILLER_70_332 ();
 sg13g2_decap_8 FILLER_70_351 ();
 sg13g2_decap_8 FILLER_70_362 ();
 sg13g2_fill_1 FILLER_70_369 ();
 sg13g2_decap_8 FILLER_70_377 ();
 sg13g2_decap_8 FILLER_70_384 ();
 sg13g2_fill_1 FILLER_70_391 ();
 sg13g2_decap_8 FILLER_70_427 ();
 sg13g2_decap_8 FILLER_70_434 ();
 sg13g2_decap_8 FILLER_70_441 ();
 sg13g2_decap_8 FILLER_70_448 ();
 sg13g2_decap_8 FILLER_70_455 ();
 sg13g2_fill_2 FILLER_70_462 ();
 sg13g2_fill_1 FILLER_70_464 ();
 sg13g2_fill_2 FILLER_70_513 ();
 sg13g2_decap_4 FILLER_70_529 ();
 sg13g2_decap_8 FILLER_70_539 ();
 sg13g2_decap_8 FILLER_70_546 ();
 sg13g2_decap_8 FILLER_70_557 ();
 sg13g2_fill_1 FILLER_70_564 ();
 sg13g2_fill_1 FILLER_70_570 ();
 sg13g2_fill_2 FILLER_70_613 ();
 sg13g2_fill_1 FILLER_70_615 ();
 sg13g2_decap_8 FILLER_70_633 ();
 sg13g2_decap_8 FILLER_70_640 ();
 sg13g2_decap_4 FILLER_70_647 ();
 sg13g2_fill_1 FILLER_70_651 ();
 sg13g2_decap_4 FILLER_70_656 ();
 sg13g2_decap_8 FILLER_70_668 ();
 sg13g2_decap_4 FILLER_70_675 ();
 sg13g2_fill_1 FILLER_70_683 ();
 sg13g2_fill_2 FILLER_70_724 ();
 sg13g2_decap_8 FILLER_70_752 ();
 sg13g2_decap_8 FILLER_70_759 ();
 sg13g2_decap_4 FILLER_70_766 ();
 sg13g2_decap_4 FILLER_70_781 ();
 sg13g2_fill_1 FILLER_70_785 ();
 sg13g2_decap_4 FILLER_70_790 ();
 sg13g2_decap_4 FILLER_70_798 ();
 sg13g2_fill_2 FILLER_70_802 ();
 sg13g2_decap_8 FILLER_70_838 ();
 sg13g2_fill_1 FILLER_70_845 ();
 sg13g2_decap_4 FILLER_70_850 ();
 sg13g2_decap_8 FILLER_70_864 ();
 sg13g2_decap_8 FILLER_70_871 ();
 sg13g2_decap_8 FILLER_70_886 ();
 sg13g2_decap_4 FILLER_70_893 ();
 sg13g2_fill_1 FILLER_70_897 ();
 sg13g2_decap_4 FILLER_70_915 ();
 sg13g2_fill_2 FILLER_70_919 ();
 sg13g2_decap_4 FILLER_70_926 ();
 sg13g2_decap_8 FILLER_70_960 ();
 sg13g2_fill_2 FILLER_70_967 ();
 sg13g2_fill_1 FILLER_70_969 ();
 sg13g2_fill_1 FILLER_70_975 ();
 sg13g2_fill_1 FILLER_70_1008 ();
 sg13g2_fill_2 FILLER_70_1027 ();
 sg13g2_fill_2 FILLER_70_1053 ();
 sg13g2_fill_1 FILLER_70_1055 ();
 sg13g2_fill_2 FILLER_70_1120 ();
 sg13g2_fill_1 FILLER_70_1140 ();
 sg13g2_fill_1 FILLER_70_1150 ();
 sg13g2_decap_8 FILLER_70_1161 ();
 sg13g2_fill_2 FILLER_70_1168 ();
 sg13g2_fill_2 FILLER_70_1244 ();
 sg13g2_fill_1 FILLER_70_1265 ();
 sg13g2_decap_4 FILLER_70_1303 ();
 sg13g2_decap_8 FILLER_70_1342 ();
 sg13g2_decap_8 FILLER_70_1349 ();
 sg13g2_fill_2 FILLER_70_1356 ();
 sg13g2_fill_1 FILLER_70_1358 ();
 sg13g2_fill_2 FILLER_70_1363 ();
 sg13g2_fill_2 FILLER_70_1375 ();
 sg13g2_fill_2 FILLER_70_1394 ();
 sg13g2_decap_4 FILLER_70_1404 ();
 sg13g2_fill_1 FILLER_70_1408 ();
 sg13g2_decap_4 FILLER_70_1419 ();
 sg13g2_decap_4 FILLER_70_1427 ();
 sg13g2_decap_8 FILLER_70_1444 ();
 sg13g2_decap_8 FILLER_70_1451 ();
 sg13g2_fill_2 FILLER_70_1468 ();
 sg13g2_fill_1 FILLER_70_1470 ();
 sg13g2_decap_8 FILLER_70_1474 ();
 sg13g2_decap_8 FILLER_70_1481 ();
 sg13g2_decap_8 FILLER_70_1488 ();
 sg13g2_decap_8 FILLER_70_1495 ();
 sg13g2_decap_8 FILLER_70_1502 ();
 sg13g2_decap_8 FILLER_70_1509 ();
 sg13g2_fill_2 FILLER_70_1516 ();
 sg13g2_fill_2 FILLER_70_1522 ();
 sg13g2_decap_8 FILLER_70_1528 ();
 sg13g2_decap_8 FILLER_70_1535 ();
 sg13g2_decap_8 FILLER_70_1542 ();
 sg13g2_decap_4 FILLER_70_1549 ();
 sg13g2_fill_1 FILLER_70_1553 ();
 sg13g2_decap_8 FILLER_70_1598 ();
 sg13g2_decap_4 FILLER_70_1605 ();
 sg13g2_fill_2 FILLER_70_1623 ();
 sg13g2_fill_1 FILLER_70_1625 ();
 sg13g2_decap_8 FILLER_70_1634 ();
 sg13g2_decap_4 FILLER_70_1641 ();
 sg13g2_fill_2 FILLER_70_1645 ();
 sg13g2_decap_4 FILLER_70_1681 ();
 sg13g2_fill_1 FILLER_70_1685 ();
 sg13g2_decap_8 FILLER_70_1721 ();
 sg13g2_decap_8 FILLER_70_1733 ();
 sg13g2_decap_8 FILLER_70_1740 ();
 sg13g2_fill_1 FILLER_70_1747 ();
 sg13g2_fill_2 FILLER_70_1823 ();
 sg13g2_fill_1 FILLER_70_1825 ();
 sg13g2_decap_4 FILLER_70_1887 ();
 sg13g2_fill_1 FILLER_70_1891 ();
 sg13g2_decap_4 FILLER_70_1897 ();
 sg13g2_fill_1 FILLER_70_1909 ();
 sg13g2_fill_1 FILLER_70_1923 ();
 sg13g2_fill_1 FILLER_70_1955 ();
 sg13g2_fill_1 FILLER_70_1985 ();
 sg13g2_fill_2 FILLER_70_1996 ();
 sg13g2_fill_2 FILLER_70_2003 ();
 sg13g2_decap_4 FILLER_70_2009 ();
 sg13g2_fill_1 FILLER_70_2013 ();
 sg13g2_fill_1 FILLER_70_2055 ();
 sg13g2_fill_2 FILLER_70_2061 ();
 sg13g2_fill_1 FILLER_70_2068 ();
 sg13g2_decap_8 FILLER_70_2100 ();
 sg13g2_decap_8 FILLER_70_2144 ();
 sg13g2_decap_4 FILLER_70_2151 ();
 sg13g2_fill_1 FILLER_70_2155 ();
 sg13g2_decap_8 FILLER_70_2165 ();
 sg13g2_decap_8 FILLER_70_2181 ();
 sg13g2_decap_8 FILLER_70_2188 ();
 sg13g2_decap_8 FILLER_70_2195 ();
 sg13g2_decap_8 FILLER_70_2202 ();
 sg13g2_decap_4 FILLER_70_2209 ();
 sg13g2_fill_2 FILLER_70_2213 ();
 sg13g2_fill_1 FILLER_70_2263 ();
 sg13g2_decap_4 FILLER_70_2268 ();
 sg13g2_fill_1 FILLER_70_2272 ();
 sg13g2_fill_1 FILLER_70_2278 ();
 sg13g2_fill_1 FILLER_70_2290 ();
 sg13g2_fill_2 FILLER_70_2307 ();
 sg13g2_fill_1 FILLER_70_2309 ();
 sg13g2_decap_4 FILLER_70_2340 ();
 sg13g2_fill_2 FILLER_70_2344 ();
 sg13g2_decap_8 FILLER_70_2352 ();
 sg13g2_decap_8 FILLER_70_2359 ();
 sg13g2_fill_1 FILLER_70_2366 ();
 sg13g2_decap_8 FILLER_70_2373 ();
 sg13g2_fill_1 FILLER_70_2380 ();
 sg13g2_fill_2 FILLER_70_2393 ();
 sg13g2_fill_1 FILLER_70_2395 ();
 sg13g2_decap_4 FILLER_70_2400 ();
 sg13g2_decap_4 FILLER_70_2430 ();
 sg13g2_fill_1 FILLER_70_2434 ();
 sg13g2_decap_8 FILLER_70_2441 ();
 sg13g2_decap_4 FILLER_70_2448 ();
 sg13g2_fill_2 FILLER_70_2467 ();
 sg13g2_decap_4 FILLER_70_2503 ();
 sg13g2_fill_1 FILLER_70_2507 ();
 sg13g2_fill_2 FILLER_70_2512 ();
 sg13g2_fill_1 FILLER_70_2514 ();
 sg13g2_decap_8 FILLER_70_2556 ();
 sg13g2_decap_4 FILLER_70_2563 ();
 sg13g2_decap_8 FILLER_70_2580 ();
 sg13g2_decap_4 FILLER_70_2587 ();
 sg13g2_fill_1 FILLER_70_2591 ();
 sg13g2_fill_1 FILLER_70_2597 ();
 sg13g2_decap_8 FILLER_70_2624 ();
 sg13g2_decap_8 FILLER_70_2635 ();
 sg13g2_decap_8 FILLER_70_2642 ();
 sg13g2_decap_8 FILLER_70_2649 ();
 sg13g2_decap_8 FILLER_70_2656 ();
 sg13g2_decap_8 FILLER_70_2663 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_4 FILLER_71_14 ();
 sg13g2_fill_1 FILLER_71_42 ();
 sg13g2_fill_1 FILLER_71_53 ();
 sg13g2_fill_2 FILLER_71_80 ();
 sg13g2_fill_2 FILLER_71_88 ();
 sg13g2_fill_1 FILLER_71_90 ();
 sg13g2_fill_2 FILLER_71_100 ();
 sg13g2_fill_1 FILLER_71_107 ();
 sg13g2_fill_1 FILLER_71_113 ();
 sg13g2_fill_1 FILLER_71_127 ();
 sg13g2_decap_4 FILLER_71_133 ();
 sg13g2_fill_1 FILLER_71_144 ();
 sg13g2_fill_1 FILLER_71_173 ();
 sg13g2_decap_4 FILLER_71_186 ();
 sg13g2_fill_1 FILLER_71_190 ();
 sg13g2_decap_8 FILLER_71_196 ();
 sg13g2_decap_8 FILLER_71_207 ();
 sg13g2_decap_8 FILLER_71_214 ();
 sg13g2_decap_4 FILLER_71_221 ();
 sg13g2_fill_1 FILLER_71_225 ();
 sg13g2_fill_2 FILLER_71_297 ();
 sg13g2_fill_1 FILLER_71_299 ();
 sg13g2_decap_4 FILLER_71_305 ();
 sg13g2_fill_1 FILLER_71_314 ();
 sg13g2_decap_8 FILLER_71_341 ();
 sg13g2_decap_4 FILLER_71_348 ();
 sg13g2_fill_1 FILLER_71_352 ();
 sg13g2_fill_2 FILLER_71_362 ();
 sg13g2_fill_1 FILLER_71_364 ();
 sg13g2_fill_1 FILLER_71_396 ();
 sg13g2_decap_8 FILLER_71_412 ();
 sg13g2_decap_4 FILLER_71_419 ();
 sg13g2_fill_1 FILLER_71_423 ();
 sg13g2_fill_1 FILLER_71_428 ();
 sg13g2_decap_8 FILLER_71_433 ();
 sg13g2_decap_8 FILLER_71_440 ();
 sg13g2_decap_8 FILLER_71_447 ();
 sg13g2_decap_4 FILLER_71_454 ();
 sg13g2_fill_2 FILLER_71_458 ();
 sg13g2_fill_2 FILLER_71_472 ();
 sg13g2_fill_2 FILLER_71_478 ();
 sg13g2_fill_2 FILLER_71_503 ();
 sg13g2_decap_8 FILLER_71_543 ();
 sg13g2_decap_8 FILLER_71_550 ();
 sg13g2_decap_8 FILLER_71_557 ();
 sg13g2_decap_8 FILLER_71_564 ();
 sg13g2_decap_8 FILLER_71_571 ();
 sg13g2_decap_8 FILLER_71_578 ();
 sg13g2_decap_4 FILLER_71_585 ();
 sg13g2_decap_8 FILLER_71_594 ();
 sg13g2_fill_2 FILLER_71_601 ();
 sg13g2_fill_1 FILLER_71_603 ();
 sg13g2_decap_4 FILLER_71_636 ();
 sg13g2_fill_1 FILLER_71_640 ();
 sg13g2_fill_1 FILLER_71_651 ();
 sg13g2_decap_4 FILLER_71_656 ();
 sg13g2_fill_2 FILLER_71_682 ();
 sg13g2_decap_8 FILLER_71_695 ();
 sg13g2_decap_4 FILLER_71_702 ();
 sg13g2_decap_8 FILLER_71_719 ();
 sg13g2_decap_8 FILLER_71_726 ();
 sg13g2_decap_8 FILLER_71_733 ();
 sg13g2_decap_8 FILLER_71_740 ();
 sg13g2_decap_8 FILLER_71_747 ();
 sg13g2_decap_8 FILLER_71_754 ();
 sg13g2_fill_1 FILLER_71_761 ();
 sg13g2_decap_4 FILLER_71_766 ();
 sg13g2_fill_1 FILLER_71_770 ();
 sg13g2_decap_8 FILLER_71_775 ();
 sg13g2_fill_2 FILLER_71_782 ();
 sg13g2_fill_2 FILLER_71_814 ();
 sg13g2_fill_1 FILLER_71_816 ();
 sg13g2_decap_4 FILLER_71_823 ();
 sg13g2_fill_2 FILLER_71_857 ();
 sg13g2_fill_1 FILLER_71_911 ();
 sg13g2_decap_4 FILLER_71_948 ();
 sg13g2_fill_1 FILLER_71_952 ();
 sg13g2_decap_8 FILLER_71_959 ();
 sg13g2_fill_1 FILLER_71_966 ();
 sg13g2_decap_8 FILLER_71_973 ();
 sg13g2_fill_2 FILLER_71_980 ();
 sg13g2_fill_1 FILLER_71_1017 ();
 sg13g2_fill_2 FILLER_71_1055 ();
 sg13g2_fill_1 FILLER_71_1062 ();
 sg13g2_fill_1 FILLER_71_1068 ();
 sg13g2_fill_1 FILLER_71_1073 ();
 sg13g2_fill_1 FILLER_71_1080 ();
 sg13g2_fill_2 FILLER_71_1085 ();
 sg13g2_fill_1 FILLER_71_1087 ();
 sg13g2_fill_2 FILLER_71_1094 ();
 sg13g2_fill_2 FILLER_71_1180 ();
 sg13g2_fill_2 FILLER_71_1260 ();
 sg13g2_fill_1 FILLER_71_1283 ();
 sg13g2_fill_1 FILLER_71_1307 ();
 sg13g2_fill_2 FILLER_71_1334 ();
 sg13g2_decap_8 FILLER_71_1341 ();
 sg13g2_fill_2 FILLER_71_1348 ();
 sg13g2_fill_1 FILLER_71_1359 ();
 sg13g2_fill_2 FILLER_71_1365 ();
 sg13g2_fill_1 FILLER_71_1375 ();
 sg13g2_fill_1 FILLER_71_1394 ();
 sg13g2_fill_1 FILLER_71_1399 ();
 sg13g2_fill_1 FILLER_71_1406 ();
 sg13g2_fill_2 FILLER_71_1412 ();
 sg13g2_decap_8 FILLER_71_1419 ();
 sg13g2_fill_1 FILLER_71_1426 ();
 sg13g2_decap_8 FILLER_71_1431 ();
 sg13g2_fill_2 FILLER_71_1438 ();
 sg13g2_decap_4 FILLER_71_1444 ();
 sg13g2_fill_2 FILLER_71_1448 ();
 sg13g2_decap_8 FILLER_71_1454 ();
 sg13g2_decap_8 FILLER_71_1461 ();
 sg13g2_fill_1 FILLER_71_1468 ();
 sg13g2_decap_4 FILLER_71_1488 ();
 sg13g2_decap_8 FILLER_71_1496 ();
 sg13g2_decap_8 FILLER_71_1503 ();
 sg13g2_decap_8 FILLER_71_1546 ();
 sg13g2_fill_2 FILLER_71_1590 ();
 sg13g2_decap_4 FILLER_71_1596 ();
 sg13g2_fill_1 FILLER_71_1600 ();
 sg13g2_decap_4 FILLER_71_1636 ();
 sg13g2_decap_8 FILLER_71_1670 ();
 sg13g2_fill_2 FILLER_71_1677 ();
 sg13g2_decap_8 FILLER_71_1713 ();
 sg13g2_decap_8 FILLER_71_1720 ();
 sg13g2_decap_8 FILLER_71_1727 ();
 sg13g2_decap_8 FILLER_71_1739 ();
 sg13g2_decap_8 FILLER_71_1746 ();
 sg13g2_decap_8 FILLER_71_1756 ();
 sg13g2_decap_8 FILLER_71_1763 ();
 sg13g2_fill_2 FILLER_71_1770 ();
 sg13g2_fill_1 FILLER_71_1814 ();
 sg13g2_fill_2 FILLER_71_1818 ();
 sg13g2_fill_2 FILLER_71_1846 ();
 sg13g2_fill_2 FILLER_71_1857 ();
 sg13g2_fill_2 FILLER_71_1863 ();
 sg13g2_fill_2 FILLER_71_1871 ();
 sg13g2_fill_2 FILLER_71_1904 ();
 sg13g2_fill_1 FILLER_71_1906 ();
 sg13g2_fill_2 FILLER_71_1948 ();
 sg13g2_fill_1 FILLER_71_1950 ();
 sg13g2_decap_8 FILLER_71_1956 ();
 sg13g2_decap_8 FILLER_71_1963 ();
 sg13g2_fill_2 FILLER_71_1986 ();
 sg13g2_decap_8 FILLER_71_2020 ();
 sg13g2_fill_2 FILLER_71_2032 ();
 sg13g2_fill_1 FILLER_71_2040 ();
 sg13g2_fill_1 FILLER_71_2045 ();
 sg13g2_fill_2 FILLER_71_2077 ();
 sg13g2_fill_1 FILLER_71_2079 ();
 sg13g2_fill_2 FILLER_71_2110 ();
 sg13g2_decap_8 FILLER_71_2142 ();
 sg13g2_fill_2 FILLER_71_2149 ();
 sg13g2_fill_1 FILLER_71_2151 ();
 sg13g2_fill_1 FILLER_71_2157 ();
 sg13g2_decap_8 FILLER_71_2210 ();
 sg13g2_decap_4 FILLER_71_2217 ();
 sg13g2_fill_2 FILLER_71_2221 ();
 sg13g2_decap_4 FILLER_71_2252 ();
 sg13g2_fill_1 FILLER_71_2256 ();
 sg13g2_decap_8 FILLER_71_2261 ();
 sg13g2_decap_4 FILLER_71_2268 ();
 sg13g2_fill_1 FILLER_71_2272 ();
 sg13g2_decap_8 FILLER_71_2311 ();
 sg13g2_fill_1 FILLER_71_2323 ();
 sg13g2_decap_8 FILLER_71_2331 ();
 sg13g2_fill_2 FILLER_71_2338 ();
 sg13g2_decap_8 FILLER_71_2352 ();
 sg13g2_fill_2 FILLER_71_2359 ();
 sg13g2_fill_1 FILLER_71_2365 ();
 sg13g2_decap_8 FILLER_71_2369 ();
 sg13g2_decap_8 FILLER_71_2376 ();
 sg13g2_fill_2 FILLER_71_2389 ();
 sg13g2_fill_1 FILLER_71_2391 ();
 sg13g2_fill_1 FILLER_71_2402 ();
 sg13g2_fill_1 FILLER_71_2429 ();
 sg13g2_fill_1 FILLER_71_2459 ();
 sg13g2_decap_4 FILLER_71_2464 ();
 sg13g2_decap_8 FILLER_71_2499 ();
 sg13g2_decap_4 FILLER_71_2506 ();
 sg13g2_decap_4 FILLER_71_2516 ();
 sg13g2_fill_2 FILLER_71_2520 ();
 sg13g2_decap_8 FILLER_71_2566 ();
 sg13g2_decap_8 FILLER_71_2573 ();
 sg13g2_decap_8 FILLER_71_2589 ();
 sg13g2_decap_8 FILLER_71_2596 ();
 sg13g2_decap_8 FILLER_71_2603 ();
 sg13g2_decap_8 FILLER_71_2610 ();
 sg13g2_decap_8 FILLER_71_2617 ();
 sg13g2_decap_8 FILLER_71_2624 ();
 sg13g2_decap_8 FILLER_71_2631 ();
 sg13g2_decap_8 FILLER_71_2638 ();
 sg13g2_decap_8 FILLER_71_2645 ();
 sg13g2_decap_8 FILLER_71_2652 ();
 sg13g2_decap_8 FILLER_71_2659 ();
 sg13g2_decap_4 FILLER_71_2666 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_4 FILLER_72_7 ();
 sg13g2_fill_1 FILLER_72_11 ();
 sg13g2_fill_1 FILLER_72_24 ();
 sg13g2_fill_2 FILLER_72_53 ();
 sg13g2_fill_1 FILLER_72_55 ();
 sg13g2_fill_1 FILLER_72_91 ();
 sg13g2_fill_2 FILLER_72_98 ();
 sg13g2_fill_1 FILLER_72_106 ();
 sg13g2_fill_1 FILLER_72_115 ();
 sg13g2_fill_2 FILLER_72_143 ();
 sg13g2_decap_4 FILLER_72_150 ();
 sg13g2_fill_2 FILLER_72_177 ();
 sg13g2_fill_1 FILLER_72_179 ();
 sg13g2_fill_1 FILLER_72_191 ();
 sg13g2_decap_4 FILLER_72_197 ();
 sg13g2_fill_2 FILLER_72_201 ();
 sg13g2_decap_8 FILLER_72_207 ();
 sg13g2_decap_4 FILLER_72_214 ();
 sg13g2_fill_1 FILLER_72_236 ();
 sg13g2_fill_1 FILLER_72_245 ();
 sg13g2_fill_2 FILLER_72_250 ();
 sg13g2_fill_2 FILLER_72_270 ();
 sg13g2_fill_2 FILLER_72_280 ();
 sg13g2_decap_4 FILLER_72_290 ();
 sg13g2_fill_2 FILLER_72_298 ();
 sg13g2_fill_1 FILLER_72_300 ();
 sg13g2_decap_8 FILLER_72_305 ();
 sg13g2_fill_2 FILLER_72_312 ();
 sg13g2_decap_8 FILLER_72_319 ();
 sg13g2_decap_8 FILLER_72_326 ();
 sg13g2_decap_8 FILLER_72_333 ();
 sg13g2_decap_8 FILLER_72_340 ();
 sg13g2_decap_4 FILLER_72_347 ();
 sg13g2_fill_2 FILLER_72_351 ();
 sg13g2_decap_4 FILLER_72_363 ();
 sg13g2_decap_8 FILLER_72_381 ();
 sg13g2_decap_4 FILLER_72_388 ();
 sg13g2_fill_2 FILLER_72_392 ();
 sg13g2_decap_8 FILLER_72_397 ();
 sg13g2_fill_1 FILLER_72_437 ();
 sg13g2_fill_2 FILLER_72_506 ();
 sg13g2_decap_4 FILLER_72_546 ();
 sg13g2_decap_8 FILLER_72_555 ();
 sg13g2_fill_2 FILLER_72_562 ();
 sg13g2_decap_8 FILLER_72_571 ();
 sg13g2_fill_2 FILLER_72_578 ();
 sg13g2_decap_8 FILLER_72_594 ();
 sg13g2_decap_4 FILLER_72_601 ();
 sg13g2_fill_2 FILLER_72_605 ();
 sg13g2_fill_2 FILLER_72_611 ();
 sg13g2_fill_1 FILLER_72_613 ();
 sg13g2_decap_4 FILLER_72_618 ();
 sg13g2_fill_1 FILLER_72_622 ();
 sg13g2_decap_8 FILLER_72_628 ();
 sg13g2_fill_1 FILLER_72_635 ();
 sg13g2_decap_4 FILLER_72_646 ();
 sg13g2_fill_1 FILLER_72_650 ();
 sg13g2_decap_4 FILLER_72_659 ();
 sg13g2_decap_8 FILLER_72_672 ();
 sg13g2_decap_8 FILLER_72_679 ();
 sg13g2_decap_4 FILLER_72_686 ();
 sg13g2_fill_1 FILLER_72_690 ();
 sg13g2_fill_2 FILLER_72_701 ();
 sg13g2_fill_1 FILLER_72_703 ();
 sg13g2_decap_8 FILLER_72_713 ();
 sg13g2_decap_4 FILLER_72_720 ();
 sg13g2_fill_2 FILLER_72_763 ();
 sg13g2_fill_1 FILLER_72_765 ();
 sg13g2_decap_8 FILLER_72_826 ();
 sg13g2_fill_2 FILLER_72_833 ();
 sg13g2_decap_4 FILLER_72_861 ();
 sg13g2_fill_2 FILLER_72_869 ();
 sg13g2_decap_8 FILLER_72_875 ();
 sg13g2_fill_2 FILLER_72_882 ();
 sg13g2_fill_1 FILLER_72_884 ();
 sg13g2_fill_2 FILLER_72_919 ();
 sg13g2_decap_4 FILLER_72_926 ();
 sg13g2_decap_8 FILLER_72_934 ();
 sg13g2_fill_1 FILLER_72_941 ();
 sg13g2_decap_8 FILLER_72_947 ();
 sg13g2_decap_8 FILLER_72_963 ();
 sg13g2_fill_1 FILLER_72_970 ();
 sg13g2_decap_4 FILLER_72_975 ();
 sg13g2_fill_2 FILLER_72_979 ();
 sg13g2_fill_1 FILLER_72_1052 ();
 sg13g2_decap_8 FILLER_72_1084 ();
 sg13g2_fill_2 FILLER_72_1096 ();
 sg13g2_fill_1 FILLER_72_1138 ();
 sg13g2_fill_2 FILLER_72_1143 ();
 sg13g2_fill_2 FILLER_72_1179 ();
 sg13g2_fill_1 FILLER_72_1181 ();
 sg13g2_fill_2 FILLER_72_1197 ();
 sg13g2_fill_2 FILLER_72_1220 ();
 sg13g2_fill_1 FILLER_72_1222 ();
 sg13g2_fill_1 FILLER_72_1291 ();
 sg13g2_fill_1 FILLER_72_1329 ();
 sg13g2_fill_2 FILLER_72_1335 ();
 sg13g2_fill_2 FILLER_72_1406 ();
 sg13g2_fill_1 FILLER_72_1408 ();
 sg13g2_fill_2 FILLER_72_1413 ();
 sg13g2_fill_1 FILLER_72_1415 ();
 sg13g2_fill_2 FILLER_72_1468 ();
 sg13g2_fill_1 FILLER_72_1476 ();
 sg13g2_decap_8 FILLER_72_1511 ();
 sg13g2_decap_4 FILLER_72_1518 ();
 sg13g2_fill_2 FILLER_72_1522 ();
 sg13g2_decap_8 FILLER_72_1533 ();
 sg13g2_decap_8 FILLER_72_1540 ();
 sg13g2_fill_1 FILLER_72_1547 ();
 sg13g2_fill_2 FILLER_72_1579 ();
 sg13g2_fill_1 FILLER_72_1581 ();
 sg13g2_decap_8 FILLER_72_1716 ();
 sg13g2_fill_2 FILLER_72_1723 ();
 sg13g2_decap_4 FILLER_72_1736 ();
 sg13g2_fill_1 FILLER_72_1740 ();
 sg13g2_fill_1 FILLER_72_1762 ();
 sg13g2_fill_1 FILLER_72_1777 ();
 sg13g2_fill_2 FILLER_72_1790 ();
 sg13g2_fill_2 FILLER_72_1810 ();
 sg13g2_decap_8 FILLER_72_1831 ();
 sg13g2_decap_4 FILLER_72_1838 ();
 sg13g2_decap_4 FILLER_72_1847 ();
 sg13g2_fill_1 FILLER_72_1851 ();
 sg13g2_fill_2 FILLER_72_1857 ();
 sg13g2_fill_1 FILLER_72_1859 ();
 sg13g2_fill_2 FILLER_72_1891 ();
 sg13g2_decap_8 FILLER_72_1899 ();
 sg13g2_decap_4 FILLER_72_1906 ();
 sg13g2_fill_2 FILLER_72_1913 ();
 sg13g2_fill_1 FILLER_72_1915 ();
 sg13g2_decap_8 FILLER_72_1921 ();
 sg13g2_decap_8 FILLER_72_1928 ();
 sg13g2_decap_8 FILLER_72_1935 ();
 sg13g2_fill_2 FILLER_72_1942 ();
 sg13g2_fill_1 FILLER_72_1944 ();
 sg13g2_decap_4 FILLER_72_1957 ();
 sg13g2_fill_2 FILLER_72_1979 ();
 sg13g2_decap_8 FILLER_72_1993 ();
 sg13g2_fill_2 FILLER_72_2000 ();
 sg13g2_fill_1 FILLER_72_2002 ();
 sg13g2_fill_2 FILLER_72_2032 ();
 sg13g2_decap_4 FILLER_72_2040 ();
 sg13g2_decap_4 FILLER_72_2048 ();
 sg13g2_fill_1 FILLER_72_2065 ();
 sg13g2_fill_2 FILLER_72_2101 ();
 sg13g2_fill_1 FILLER_72_2103 ();
 sg13g2_decap_8 FILLER_72_2116 ();
 sg13g2_fill_2 FILLER_72_2123 ();
 sg13g2_decap_8 FILLER_72_2139 ();
 sg13g2_decap_8 FILLER_72_2146 ();
 sg13g2_decap_4 FILLER_72_2153 ();
 sg13g2_fill_1 FILLER_72_2157 ();
 sg13g2_decap_4 FILLER_72_2164 ();
 sg13g2_decap_8 FILLER_72_2236 ();
 sg13g2_decap_4 FILLER_72_2243 ();
 sg13g2_fill_2 FILLER_72_2247 ();
 sg13g2_decap_8 FILLER_72_2280 ();
 sg13g2_decap_8 FILLER_72_2287 ();
 sg13g2_decap_8 FILLER_72_2294 ();
 sg13g2_decap_8 FILLER_72_2301 ();
 sg13g2_decap_4 FILLER_72_2308 ();
 sg13g2_decap_8 FILLER_72_2317 ();
 sg13g2_decap_4 FILLER_72_2324 ();
 sg13g2_fill_1 FILLER_72_2341 ();
 sg13g2_fill_1 FILLER_72_2348 ();
 sg13g2_fill_1 FILLER_72_2355 ();
 sg13g2_fill_2 FILLER_72_2361 ();
 sg13g2_fill_1 FILLER_72_2372 ();
 sg13g2_decap_4 FILLER_72_2377 ();
 sg13g2_fill_1 FILLER_72_2381 ();
 sg13g2_decap_8 FILLER_72_2412 ();
 sg13g2_decap_8 FILLER_72_2419 ();
 sg13g2_fill_2 FILLER_72_2432 ();
 sg13g2_fill_1 FILLER_72_2434 ();
 sg13g2_decap_4 FILLER_72_2470 ();
 sg13g2_fill_2 FILLER_72_2474 ();
 sg13g2_fill_2 FILLER_72_2485 ();
 sg13g2_decap_8 FILLER_72_2500 ();
 sg13g2_decap_8 FILLER_72_2507 ();
 sg13g2_decap_8 FILLER_72_2514 ();
 sg13g2_fill_2 FILLER_72_2521 ();
 sg13g2_decap_4 FILLER_72_2563 ();
 sg13g2_decap_8 FILLER_72_2571 ();
 sg13g2_fill_2 FILLER_72_2578 ();
 sg13g2_fill_1 FILLER_72_2580 ();
 sg13g2_fill_2 FILLER_72_2586 ();
 sg13g2_fill_1 FILLER_72_2588 ();
 sg13g2_decap_8 FILLER_72_2615 ();
 sg13g2_decap_8 FILLER_72_2622 ();
 sg13g2_decap_8 FILLER_72_2629 ();
 sg13g2_decap_8 FILLER_72_2636 ();
 sg13g2_decap_8 FILLER_72_2643 ();
 sg13g2_decap_8 FILLER_72_2650 ();
 sg13g2_decap_8 FILLER_72_2657 ();
 sg13g2_decap_4 FILLER_72_2664 ();
 sg13g2_fill_2 FILLER_72_2668 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_fill_1 FILLER_73_22 ();
 sg13g2_fill_1 FILLER_73_54 ();
 sg13g2_fill_2 FILLER_73_64 ();
 sg13g2_fill_1 FILLER_73_74 ();
 sg13g2_fill_2 FILLER_73_80 ();
 sg13g2_fill_1 FILLER_73_92 ();
 sg13g2_decap_8 FILLER_73_102 ();
 sg13g2_decap_4 FILLER_73_109 ();
 sg13g2_decap_4 FILLER_73_117 ();
 sg13g2_fill_1 FILLER_73_125 ();
 sg13g2_fill_2 FILLER_73_136 ();
 sg13g2_fill_1 FILLER_73_138 ();
 sg13g2_fill_1 FILLER_73_143 ();
 sg13g2_fill_1 FILLER_73_149 ();
 sg13g2_fill_1 FILLER_73_155 ();
 sg13g2_fill_1 FILLER_73_162 ();
 sg13g2_fill_2 FILLER_73_190 ();
 sg13g2_fill_1 FILLER_73_192 ();
 sg13g2_fill_1 FILLER_73_198 ();
 sg13g2_fill_1 FILLER_73_203 ();
 sg13g2_decap_4 FILLER_73_208 ();
 sg13g2_fill_2 FILLER_73_215 ();
 sg13g2_fill_1 FILLER_73_217 ();
 sg13g2_fill_1 FILLER_73_223 ();
 sg13g2_fill_2 FILLER_73_270 ();
 sg13g2_fill_1 FILLER_73_284 ();
 sg13g2_decap_8 FILLER_73_326 ();
 sg13g2_decap_8 FILLER_73_333 ();
 sg13g2_decap_4 FILLER_73_396 ();
 sg13g2_fill_2 FILLER_73_400 ();
 sg13g2_decap_8 FILLER_73_437 ();
 sg13g2_decap_8 FILLER_73_444 ();
 sg13g2_decap_8 FILLER_73_451 ();
 sg13g2_decap_8 FILLER_73_458 ();
 sg13g2_fill_2 FILLER_73_465 ();
 sg13g2_fill_1 FILLER_73_467 ();
 sg13g2_fill_2 FILLER_73_500 ();
 sg13g2_decap_8 FILLER_73_546 ();
 sg13g2_decap_8 FILLER_73_553 ();
 sg13g2_decap_8 FILLER_73_591 ();
 sg13g2_decap_8 FILLER_73_598 ();
 sg13g2_decap_4 FILLER_73_605 ();
 sg13g2_fill_1 FILLER_73_609 ();
 sg13g2_decap_8 FILLER_73_615 ();
 sg13g2_decap_8 FILLER_73_622 ();
 sg13g2_decap_4 FILLER_73_629 ();
 sg13g2_fill_1 FILLER_73_633 ();
 sg13g2_fill_1 FILLER_73_665 ();
 sg13g2_fill_2 FILLER_73_670 ();
 sg13g2_decap_4 FILLER_73_698 ();
 sg13g2_fill_2 FILLER_73_702 ();
 sg13g2_decap_4 FILLER_73_714 ();
 sg13g2_fill_2 FILLER_73_718 ();
 sg13g2_decap_8 FILLER_73_728 ();
 sg13g2_decap_8 FILLER_73_735 ();
 sg13g2_decap_4 FILLER_73_742 ();
 sg13g2_decap_4 FILLER_73_772 ();
 sg13g2_decap_4 FILLER_73_780 ();
 sg13g2_decap_8 FILLER_73_816 ();
 sg13g2_decap_8 FILLER_73_823 ();
 sg13g2_decap_8 FILLER_73_853 ();
 sg13g2_fill_2 FILLER_73_860 ();
 sg13g2_fill_1 FILLER_73_868 ();
 sg13g2_fill_1 FILLER_73_895 ();
 sg13g2_decap_4 FILLER_73_900 ();
 sg13g2_fill_2 FILLER_73_904 ();
 sg13g2_decap_8 FILLER_73_962 ();
 sg13g2_decap_8 FILLER_73_969 ();
 sg13g2_fill_2 FILLER_73_976 ();
 sg13g2_fill_1 FILLER_73_978 ();
 sg13g2_decap_8 FILLER_73_988 ();
 sg13g2_fill_2 FILLER_73_1025 ();
 sg13g2_decap_8 FILLER_73_1050 ();
 sg13g2_decap_8 FILLER_73_1057 ();
 sg13g2_decap_8 FILLER_73_1064 ();
 sg13g2_decap_8 FILLER_73_1071 ();
 sg13g2_decap_8 FILLER_73_1078 ();
 sg13g2_fill_2 FILLER_73_1085 ();
 sg13g2_fill_1 FILLER_73_1087 ();
 sg13g2_fill_2 FILLER_73_1118 ();
 sg13g2_decap_8 FILLER_73_1133 ();
 sg13g2_decap_4 FILLER_73_1140 ();
 sg13g2_fill_2 FILLER_73_1144 ();
 sg13g2_fill_2 FILLER_73_1175 ();
 sg13g2_fill_2 FILLER_73_1186 ();
 sg13g2_fill_1 FILLER_73_1188 ();
 sg13g2_decap_8 FILLER_73_1215 ();
 sg13g2_fill_1 FILLER_73_1222 ();
 sg13g2_fill_2 FILLER_73_1282 ();
 sg13g2_fill_2 FILLER_73_1299 ();
 sg13g2_fill_1 FILLER_73_1304 ();
 sg13g2_fill_1 FILLER_73_1314 ();
 sg13g2_fill_1 FILLER_73_1375 ();
 sg13g2_fill_2 FILLER_73_1386 ();
 sg13g2_decap_8 FILLER_73_1443 ();
 sg13g2_fill_1 FILLER_73_1469 ();
 sg13g2_fill_2 FILLER_73_1475 ();
 sg13g2_fill_1 FILLER_73_1477 ();
 sg13g2_fill_2 FILLER_73_1518 ();
 sg13g2_fill_1 FILLER_73_1520 ();
 sg13g2_decap_4 FILLER_73_1551 ();
 sg13g2_fill_2 FILLER_73_1555 ();
 sg13g2_fill_2 FILLER_73_1561 ();
 sg13g2_fill_1 FILLER_73_1563 ();
 sg13g2_decap_8 FILLER_73_1570 ();
 sg13g2_fill_2 FILLER_73_1577 ();
 sg13g2_fill_2 FILLER_73_1585 ();
 sg13g2_fill_2 FILLER_73_1613 ();
 sg13g2_fill_2 FILLER_73_1632 ();
 sg13g2_fill_1 FILLER_73_1652 ();
 sg13g2_fill_1 FILLER_73_1662 ();
 sg13g2_fill_2 FILLER_73_1667 ();
 sg13g2_decap_8 FILLER_73_1717 ();
 sg13g2_decap_4 FILLER_73_1750 ();
 sg13g2_fill_2 FILLER_73_1754 ();
 sg13g2_fill_1 FILLER_73_1789 ();
 sg13g2_fill_1 FILLER_73_1796 ();
 sg13g2_decap_4 FILLER_73_1810 ();
 sg13g2_fill_1 FILLER_73_1814 ();
 sg13g2_decap_8 FILLER_73_1821 ();
 sg13g2_decap_8 FILLER_73_1828 ();
 sg13g2_decap_4 FILLER_73_1840 ();
 sg13g2_fill_1 FILLER_73_1870 ();
 sg13g2_fill_2 FILLER_73_1878 ();
 sg13g2_decap_4 FILLER_73_1885 ();
 sg13g2_fill_2 FILLER_73_1889 ();
 sg13g2_decap_4 FILLER_73_1933 ();
 sg13g2_fill_2 FILLER_73_1941 ();
 sg13g2_decap_8 FILLER_73_1964 ();
 sg13g2_decap_4 FILLER_73_1971 ();
 sg13g2_decap_8 FILLER_73_1985 ();
 sg13g2_fill_2 FILLER_73_1992 ();
 sg13g2_fill_1 FILLER_73_1999 ();
 sg13g2_fill_1 FILLER_73_2013 ();
 sg13g2_decap_8 FILLER_73_2027 ();
 sg13g2_fill_2 FILLER_73_2034 ();
 sg13g2_fill_2 FILLER_73_2040 ();
 sg13g2_fill_1 FILLER_73_2042 ();
 sg13g2_decap_8 FILLER_73_2054 ();
 sg13g2_decap_8 FILLER_73_2061 ();
 sg13g2_fill_1 FILLER_73_2068 ();
 sg13g2_decap_4 FILLER_73_2098 ();
 sg13g2_decap_4 FILLER_73_2140 ();
 sg13g2_fill_1 FILLER_73_2148 ();
 sg13g2_fill_2 FILLER_73_2154 ();
 sg13g2_fill_1 FILLER_73_2156 ();
 sg13g2_fill_2 FILLER_73_2161 ();
 sg13g2_fill_1 FILLER_73_2163 ();
 sg13g2_decap_4 FILLER_73_2181 ();
 sg13g2_fill_2 FILLER_73_2185 ();
 sg13g2_decap_8 FILLER_73_2191 ();
 sg13g2_fill_2 FILLER_73_2209 ();
 sg13g2_fill_2 FILLER_73_2220 ();
 sg13g2_decap_8 FILLER_73_2239 ();
 sg13g2_fill_2 FILLER_73_2246 ();
 sg13g2_fill_1 FILLER_73_2248 ();
 sg13g2_fill_2 FILLER_73_2258 ();
 sg13g2_decap_8 FILLER_73_2264 ();
 sg13g2_decap_4 FILLER_73_2271 ();
 sg13g2_fill_1 FILLER_73_2275 ();
 sg13g2_fill_2 FILLER_73_2327 ();
 sg13g2_fill_1 FILLER_73_2393 ();
 sg13g2_fill_1 FILLER_73_2398 ();
 sg13g2_decap_8 FILLER_73_2425 ();
 sg13g2_fill_2 FILLER_73_2432 ();
 sg13g2_fill_1 FILLER_73_2434 ();
 sg13g2_fill_2 FILLER_73_2447 ();
 sg13g2_fill_1 FILLER_73_2454 ();
 sg13g2_fill_2 FILLER_73_2481 ();
 sg13g2_decap_8 FILLER_73_2509 ();
 sg13g2_fill_2 FILLER_73_2516 ();
 sg13g2_fill_1 FILLER_73_2518 ();
 sg13g2_decap_8 FILLER_73_2530 ();
 sg13g2_decap_8 FILLER_73_2537 ();
 sg13g2_decap_4 FILLER_73_2544 ();
 sg13g2_fill_1 FILLER_73_2548 ();
 sg13g2_fill_2 FILLER_73_2553 ();
 sg13g2_fill_1 FILLER_73_2555 ();
 sg13g2_fill_2 FILLER_73_2596 ();
 sg13g2_decap_8 FILLER_73_2624 ();
 sg13g2_decap_8 FILLER_73_2631 ();
 sg13g2_decap_8 FILLER_73_2638 ();
 sg13g2_decap_8 FILLER_73_2645 ();
 sg13g2_decap_8 FILLER_73_2652 ();
 sg13g2_decap_8 FILLER_73_2659 ();
 sg13g2_decap_4 FILLER_73_2666 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_7 ();
 sg13g2_fill_2 FILLER_74_11 ();
 sg13g2_fill_2 FILLER_74_37 ();
 sg13g2_fill_1 FILLER_74_39 ();
 sg13g2_fill_1 FILLER_74_44 ();
 sg13g2_fill_1 FILLER_74_59 ();
 sg13g2_fill_1 FILLER_74_64 ();
 sg13g2_fill_1 FILLER_74_69 ();
 sg13g2_fill_1 FILLER_74_74 ();
 sg13g2_fill_1 FILLER_74_80 ();
 sg13g2_fill_2 FILLER_74_90 ();
 sg13g2_decap_8 FILLER_74_97 ();
 sg13g2_fill_2 FILLER_74_117 ();
 sg13g2_fill_1 FILLER_74_125 ();
 sg13g2_fill_1 FILLER_74_131 ();
 sg13g2_fill_2 FILLER_74_145 ();
 sg13g2_fill_1 FILLER_74_154 ();
 sg13g2_fill_1 FILLER_74_160 ();
 sg13g2_fill_2 FILLER_74_174 ();
 sg13g2_fill_1 FILLER_74_176 ();
 sg13g2_fill_2 FILLER_74_193 ();
 sg13g2_fill_1 FILLER_74_195 ();
 sg13g2_decap_8 FILLER_74_201 ();
 sg13g2_fill_1 FILLER_74_208 ();
 sg13g2_fill_1 FILLER_74_213 ();
 sg13g2_decap_4 FILLER_74_222 ();
 sg13g2_fill_1 FILLER_74_237 ();
 sg13g2_decap_4 FILLER_74_243 ();
 sg13g2_fill_2 FILLER_74_247 ();
 sg13g2_decap_8 FILLER_74_268 ();
 sg13g2_fill_2 FILLER_74_275 ();
 sg13g2_fill_1 FILLER_74_277 ();
 sg13g2_decap_8 FILLER_74_281 ();
 sg13g2_decap_4 FILLER_74_288 ();
 sg13g2_fill_2 FILLER_74_310 ();
 sg13g2_decap_8 FILLER_74_343 ();
 sg13g2_decap_8 FILLER_74_350 ();
 sg13g2_decap_8 FILLER_74_357 ();
 sg13g2_fill_2 FILLER_74_364 ();
 sg13g2_decap_8 FILLER_74_382 ();
 sg13g2_decap_8 FILLER_74_389 ();
 sg13g2_fill_1 FILLER_74_396 ();
 sg13g2_decap_8 FILLER_74_446 ();
 sg13g2_decap_8 FILLER_74_453 ();
 sg13g2_decap_8 FILLER_74_460 ();
 sg13g2_decap_4 FILLER_74_467 ();
 sg13g2_fill_1 FILLER_74_475 ();
 sg13g2_fill_2 FILLER_74_491 ();
 sg13g2_fill_1 FILLER_74_503 ();
 sg13g2_decap_4 FILLER_74_527 ();
 sg13g2_decap_8 FILLER_74_541 ();
 sg13g2_decap_8 FILLER_74_548 ();
 sg13g2_decap_8 FILLER_74_555 ();
 sg13g2_decap_8 FILLER_74_566 ();
 sg13g2_decap_8 FILLER_74_609 ();
 sg13g2_decap_8 FILLER_74_616 ();
 sg13g2_decap_8 FILLER_74_623 ();
 sg13g2_fill_2 FILLER_74_630 ();
 sg13g2_fill_1 FILLER_74_662 ();
 sg13g2_decap_8 FILLER_74_668 ();
 sg13g2_fill_1 FILLER_74_675 ();
 sg13g2_decap_8 FILLER_74_686 ();
 sg13g2_decap_8 FILLER_74_693 ();
 sg13g2_decap_4 FILLER_74_700 ();
 sg13g2_decap_4 FILLER_74_709 ();
 sg13g2_decap_4 FILLER_74_744 ();
 sg13g2_fill_1 FILLER_74_748 ();
 sg13g2_decap_4 FILLER_74_785 ();
 sg13g2_fill_2 FILLER_74_789 ();
 sg13g2_decap_8 FILLER_74_795 ();
 sg13g2_decap_8 FILLER_74_806 ();
 sg13g2_fill_2 FILLER_74_813 ();
 sg13g2_fill_1 FILLER_74_815 ();
 sg13g2_decap_8 FILLER_74_882 ();
 sg13g2_decap_8 FILLER_74_889 ();
 sg13g2_decap_8 FILLER_74_896 ();
 sg13g2_decap_8 FILLER_74_903 ();
 sg13g2_decap_8 FILLER_74_910 ();
 sg13g2_decap_8 FILLER_74_917 ();
 sg13g2_fill_1 FILLER_74_924 ();
 sg13g2_decap_8 FILLER_74_1006 ();
 sg13g2_fill_2 FILLER_74_1045 ();
 sg13g2_fill_1 FILLER_74_1052 ();
 sg13g2_decap_8 FILLER_74_1057 ();
 sg13g2_decap_8 FILLER_74_1064 ();
 sg13g2_decap_4 FILLER_74_1071 ();
 sg13g2_fill_1 FILLER_74_1075 ();
 sg13g2_fill_2 FILLER_74_1102 ();
 sg13g2_decap_8 FILLER_74_1122 ();
 sg13g2_decap_8 FILLER_74_1129 ();
 sg13g2_decap_8 FILLER_74_1136 ();
 sg13g2_decap_8 FILLER_74_1143 ();
 sg13g2_decap_4 FILLER_74_1150 ();
 sg13g2_fill_1 FILLER_74_1154 ();
 sg13g2_fill_1 FILLER_74_1160 ();
 sg13g2_decap_8 FILLER_74_1165 ();
 sg13g2_decap_8 FILLER_74_1184 ();
 sg13g2_fill_2 FILLER_74_1191 ();
 sg13g2_fill_1 FILLER_74_1193 ();
 sg13g2_decap_4 FILLER_74_1207 ();
 sg13g2_decap_8 FILLER_74_1215 ();
 sg13g2_fill_1 FILLER_74_1235 ();
 sg13g2_fill_1 FILLER_74_1246 ();
 sg13g2_fill_1 FILLER_74_1253 ();
 sg13g2_fill_2 FILLER_74_1258 ();
 sg13g2_fill_1 FILLER_74_1260 ();
 sg13g2_fill_1 FILLER_74_1269 ();
 sg13g2_fill_2 FILLER_74_1291 ();
 sg13g2_fill_1 FILLER_74_1355 ();
 sg13g2_fill_1 FILLER_74_1365 ();
 sg13g2_fill_2 FILLER_74_1371 ();
 sg13g2_fill_1 FILLER_74_1387 ();
 sg13g2_fill_2 FILLER_74_1394 ();
 sg13g2_decap_8 FILLER_74_1407 ();
 sg13g2_decap_4 FILLER_74_1414 ();
 sg13g2_decap_8 FILLER_74_1435 ();
 sg13g2_fill_2 FILLER_74_1442 ();
 sg13g2_decap_8 FILLER_74_1448 ();
 sg13g2_decap_8 FILLER_74_1455 ();
 sg13g2_decap_4 FILLER_74_1462 ();
 sg13g2_fill_1 FILLER_74_1470 ();
 sg13g2_fill_2 FILLER_74_1476 ();
 sg13g2_fill_1 FILLER_74_1509 ();
 sg13g2_fill_2 FILLER_74_1516 ();
 sg13g2_decap_8 FILLER_74_1548 ();
 sg13g2_fill_2 FILLER_74_1555 ();
 sg13g2_fill_1 FILLER_74_1557 ();
 sg13g2_fill_2 FILLER_74_1562 ();
 sg13g2_decap_4 FILLER_74_1570 ();
 sg13g2_fill_1 FILLER_74_1585 ();
 sg13g2_fill_1 FILLER_74_1665 ();
 sg13g2_fill_2 FILLER_74_1695 ();
 sg13g2_decap_8 FILLER_74_1753 ();
 sg13g2_decap_4 FILLER_74_1760 ();
 sg13g2_fill_2 FILLER_74_1764 ();
 sg13g2_fill_2 FILLER_74_1771 ();
 sg13g2_fill_1 FILLER_74_1773 ();
 sg13g2_fill_1 FILLER_74_1778 ();
 sg13g2_fill_2 FILLER_74_1788 ();
 sg13g2_decap_8 FILLER_74_1804 ();
 sg13g2_decap_8 FILLER_74_1811 ();
 sg13g2_decap_8 FILLER_74_1818 ();
 sg13g2_decap_8 FILLER_74_1825 ();
 sg13g2_decap_8 FILLER_74_1832 ();
 sg13g2_decap_8 FILLER_74_1839 ();
 sg13g2_decap_8 FILLER_74_1846 ();
 sg13g2_decap_8 FILLER_74_1853 ();
 sg13g2_decap_4 FILLER_74_1860 ();
 sg13g2_fill_2 FILLER_74_1864 ();
 sg13g2_fill_2 FILLER_74_1875 ();
 sg13g2_fill_2 FILLER_74_1882 ();
 sg13g2_fill_1 FILLER_74_1884 ();
 sg13g2_decap_4 FILLER_74_1895 ();
 sg13g2_fill_2 FILLER_74_1918 ();
 sg13g2_fill_1 FILLER_74_1920 ();
 sg13g2_fill_1 FILLER_74_1951 ();
 sg13g2_fill_2 FILLER_74_1979 ();
 sg13g2_fill_1 FILLER_74_1981 ();
 sg13g2_fill_2 FILLER_74_1988 ();
 sg13g2_fill_1 FILLER_74_1990 ();
 sg13g2_decap_8 FILLER_74_2017 ();
 sg13g2_decap_4 FILLER_74_2024 ();
 sg13g2_fill_2 FILLER_74_2034 ();
 sg13g2_decap_8 FILLER_74_2072 ();
 sg13g2_fill_2 FILLER_74_2079 ();
 sg13g2_fill_1 FILLER_74_2081 ();
 sg13g2_decap_8 FILLER_74_2095 ();
 sg13g2_decap_8 FILLER_74_2108 ();
 sg13g2_decap_4 FILLER_74_2115 ();
 sg13g2_decap_8 FILLER_74_2124 ();
 sg13g2_decap_8 FILLER_74_2131 ();
 sg13g2_decap_8 FILLER_74_2138 ();
 sg13g2_decap_8 FILLER_74_2171 ();
 sg13g2_decap_4 FILLER_74_2178 ();
 sg13g2_fill_2 FILLER_74_2182 ();
 sg13g2_decap_8 FILLER_74_2189 ();
 sg13g2_fill_2 FILLER_74_2200 ();
 sg13g2_fill_2 FILLER_74_2228 ();
 sg13g2_fill_1 FILLER_74_2230 ();
 sg13g2_fill_2 FILLER_74_2236 ();
 sg13g2_fill_1 FILLER_74_2242 ();
 sg13g2_decap_8 FILLER_74_2248 ();
 sg13g2_decap_8 FILLER_74_2255 ();
 sg13g2_decap_8 FILLER_74_2262 ();
 sg13g2_fill_1 FILLER_74_2269 ();
 sg13g2_fill_1 FILLER_74_2275 ();
 sg13g2_fill_1 FILLER_74_2282 ();
 sg13g2_fill_1 FILLER_74_2289 ();
 sg13g2_fill_2 FILLER_74_2301 ();
 sg13g2_decap_4 FILLER_74_2310 ();
 sg13g2_fill_2 FILLER_74_2314 ();
 sg13g2_decap_8 FILLER_74_2363 ();
 sg13g2_decap_8 FILLER_74_2370 ();
 sg13g2_fill_1 FILLER_74_2377 ();
 sg13g2_fill_1 FILLER_74_2396 ();
 sg13g2_fill_1 FILLER_74_2403 ();
 sg13g2_fill_2 FILLER_74_2424 ();
 sg13g2_fill_1 FILLER_74_2426 ();
 sg13g2_decap_8 FILLER_74_2436 ();
 sg13g2_fill_1 FILLER_74_2443 ();
 sg13g2_fill_1 FILLER_74_2453 ();
 sg13g2_decap_4 FILLER_74_2458 ();
 sg13g2_fill_1 FILLER_74_2467 ();
 sg13g2_decap_4 FILLER_74_2500 ();
 sg13g2_fill_2 FILLER_74_2509 ();
 sg13g2_fill_1 FILLER_74_2511 ();
 sg13g2_decap_4 FILLER_74_2568 ();
 sg13g2_fill_2 FILLER_74_2585 ();
 sg13g2_decap_4 FILLER_74_2600 ();
 sg13g2_fill_1 FILLER_74_2604 ();
 sg13g2_decap_8 FILLER_74_2631 ();
 sg13g2_decap_8 FILLER_74_2638 ();
 sg13g2_decap_8 FILLER_74_2645 ();
 sg13g2_decap_8 FILLER_74_2652 ();
 sg13g2_decap_8 FILLER_74_2659 ();
 sg13g2_decap_4 FILLER_74_2666 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_7 ();
 sg13g2_fill_1 FILLER_75_14 ();
 sg13g2_fill_1 FILLER_75_43 ();
 sg13g2_fill_2 FILLER_75_56 ();
 sg13g2_fill_1 FILLER_75_58 ();
 sg13g2_fill_2 FILLER_75_74 ();
 sg13g2_fill_2 FILLER_75_118 ();
 sg13g2_fill_1 FILLER_75_120 ();
 sg13g2_fill_2 FILLER_75_140 ();
 sg13g2_fill_1 FILLER_75_155 ();
 sg13g2_fill_2 FILLER_75_173 ();
 sg13g2_decap_4 FILLER_75_180 ();
 sg13g2_decap_8 FILLER_75_197 ();
 sg13g2_decap_8 FILLER_75_204 ();
 sg13g2_fill_2 FILLER_75_211 ();
 sg13g2_fill_2 FILLER_75_238 ();
 sg13g2_decap_4 FILLER_75_245 ();
 sg13g2_decap_4 FILLER_75_271 ();
 sg13g2_fill_1 FILLER_75_275 ();
 sg13g2_fill_1 FILLER_75_283 ();
 sg13g2_fill_2 FILLER_75_323 ();
 sg13g2_fill_1 FILLER_75_325 ();
 sg13g2_decap_8 FILLER_75_333 ();
 sg13g2_decap_8 FILLER_75_340 ();
 sg13g2_decap_8 FILLER_75_347 ();
 sg13g2_fill_2 FILLER_75_354 ();
 sg13g2_fill_1 FILLER_75_364 ();
 sg13g2_fill_2 FILLER_75_379 ();
 sg13g2_fill_1 FILLER_75_381 ();
 sg13g2_fill_1 FILLER_75_403 ();
 sg13g2_fill_2 FILLER_75_417 ();
 sg13g2_fill_2 FILLER_75_424 ();
 sg13g2_decap_8 FILLER_75_443 ();
 sg13g2_decap_4 FILLER_75_450 ();
 sg13g2_fill_2 FILLER_75_454 ();
 sg13g2_fill_2 FILLER_75_498 ();
 sg13g2_fill_1 FILLER_75_505 ();
 sg13g2_fill_2 FILLER_75_543 ();
 sg13g2_decap_8 FILLER_75_553 ();
 sg13g2_decap_8 FILLER_75_560 ();
 sg13g2_decap_8 FILLER_75_577 ();
 sg13g2_decap_4 FILLER_75_584 ();
 sg13g2_fill_1 FILLER_75_588 ();
 sg13g2_decap_4 FILLER_75_615 ();
 sg13g2_fill_2 FILLER_75_619 ();
 sg13g2_fill_1 FILLER_75_627 ();
 sg13g2_fill_1 FILLER_75_684 ();
 sg13g2_decap_8 FILLER_75_691 ();
 sg13g2_fill_2 FILLER_75_698 ();
 sg13g2_fill_1 FILLER_75_700 ();
 sg13g2_decap_8 FILLER_75_710 ();
 sg13g2_decap_8 FILLER_75_717 ();
 sg13g2_decap_8 FILLER_75_724 ();
 sg13g2_fill_2 FILLER_75_736 ();
 sg13g2_decap_4 FILLER_75_742 ();
 sg13g2_fill_2 FILLER_75_746 ();
 sg13g2_fill_1 FILLER_75_778 ();
 sg13g2_decap_8 FILLER_75_785 ();
 sg13g2_decap_8 FILLER_75_792 ();
 sg13g2_decap_8 FILLER_75_799 ();
 sg13g2_decap_4 FILLER_75_806 ();
 sg13g2_fill_1 FILLER_75_810 ();
 sg13g2_decap_4 FILLER_75_847 ();
 sg13g2_fill_2 FILLER_75_851 ();
 sg13g2_decap_8 FILLER_75_857 ();
 sg13g2_decap_8 FILLER_75_864 ();
 sg13g2_decap_8 FILLER_75_871 ();
 sg13g2_decap_8 FILLER_75_878 ();
 sg13g2_decap_8 FILLER_75_885 ();
 sg13g2_decap_8 FILLER_75_892 ();
 sg13g2_decap_8 FILLER_75_899 ();
 sg13g2_fill_2 FILLER_75_906 ();
 sg13g2_fill_1 FILLER_75_908 ();
 sg13g2_decap_8 FILLER_75_969 ();
 sg13g2_decap_8 FILLER_75_976 ();
 sg13g2_fill_1 FILLER_75_983 ();
 sg13g2_decap_4 FILLER_75_990 ();
 sg13g2_decap_8 FILLER_75_1000 ();
 sg13g2_decap_8 FILLER_75_1007 ();
 sg13g2_decap_4 FILLER_75_1014 ();
 sg13g2_fill_2 FILLER_75_1036 ();
 sg13g2_decap_4 FILLER_75_1100 ();
 sg13g2_fill_2 FILLER_75_1113 ();
 sg13g2_decap_8 FILLER_75_1141 ();
 sg13g2_decap_8 FILLER_75_1148 ();
 sg13g2_decap_8 FILLER_75_1155 ();
 sg13g2_decap_8 FILLER_75_1162 ();
 sg13g2_decap_8 FILLER_75_1169 ();
 sg13g2_decap_8 FILLER_75_1176 ();
 sg13g2_decap_8 FILLER_75_1183 ();
 sg13g2_decap_4 FILLER_75_1190 ();
 sg13g2_decap_8 FILLER_75_1207 ();
 sg13g2_decap_8 FILLER_75_1214 ();
 sg13g2_decap_8 FILLER_75_1221 ();
 sg13g2_decap_8 FILLER_75_1228 ();
 sg13g2_decap_8 FILLER_75_1235 ();
 sg13g2_fill_2 FILLER_75_1258 ();
 sg13g2_fill_1 FILLER_75_1265 ();
 sg13g2_fill_2 FILLER_75_1335 ();
 sg13g2_fill_2 FILLER_75_1349 ();
 sg13g2_fill_2 FILLER_75_1413 ();
 sg13g2_fill_1 FILLER_75_1415 ();
 sg13g2_decap_4 FILLER_75_1502 ();
 sg13g2_fill_2 FILLER_75_1506 ();
 sg13g2_decap_8 FILLER_75_1516 ();
 sg13g2_decap_8 FILLER_75_1523 ();
 sg13g2_fill_2 FILLER_75_1530 ();
 sg13g2_fill_1 FILLER_75_1532 ();
 sg13g2_decap_8 FILLER_75_1543 ();
 sg13g2_decap_8 FILLER_75_1550 ();
 sg13g2_fill_2 FILLER_75_1557 ();
 sg13g2_fill_1 FILLER_75_1559 ();
 sg13g2_fill_1 FILLER_75_1564 ();
 sg13g2_decap_8 FILLER_75_1621 ();
 sg13g2_decap_8 FILLER_75_1646 ();
 sg13g2_decap_4 FILLER_75_1688 ();
 sg13g2_decap_8 FILLER_75_1705 ();
 sg13g2_decap_8 FILLER_75_1712 ();
 sg13g2_decap_8 FILLER_75_1719 ();
 sg13g2_decap_8 FILLER_75_1756 ();
 sg13g2_decap_4 FILLER_75_1763 ();
 sg13g2_fill_2 FILLER_75_1798 ();
 sg13g2_fill_1 FILLER_75_1800 ();
 sg13g2_decap_4 FILLER_75_1830 ();
 sg13g2_fill_1 FILLER_75_1834 ();
 sg13g2_decap_4 FILLER_75_1847 ();
 sg13g2_fill_2 FILLER_75_1906 ();
 sg13g2_fill_1 FILLER_75_1908 ();
 sg13g2_fill_2 FILLER_75_1918 ();
 sg13g2_fill_1 FILLER_75_1920 ();
 sg13g2_fill_1 FILLER_75_1965 ();
 sg13g2_decap_4 FILLER_75_1992 ();
 sg13g2_fill_2 FILLER_75_1996 ();
 sg13g2_fill_1 FILLER_75_2024 ();
 sg13g2_decap_8 FILLER_75_2064 ();
 sg13g2_decap_8 FILLER_75_2071 ();
 sg13g2_decap_4 FILLER_75_2078 ();
 sg13g2_fill_2 FILLER_75_2082 ();
 sg13g2_decap_8 FILLER_75_2110 ();
 sg13g2_decap_4 FILLER_75_2117 ();
 sg13g2_fill_2 FILLER_75_2121 ();
 sg13g2_decap_8 FILLER_75_2149 ();
 sg13g2_decap_8 FILLER_75_2156 ();
 sg13g2_decap_8 FILLER_75_2163 ();
 sg13g2_fill_2 FILLER_75_2175 ();
 sg13g2_fill_1 FILLER_75_2177 ();
 sg13g2_fill_2 FILLER_75_2182 ();
 sg13g2_fill_2 FILLER_75_2210 ();
 sg13g2_fill_1 FILLER_75_2212 ();
 sg13g2_fill_1 FILLER_75_2230 ();
 sg13g2_fill_2 FILLER_75_2261 ();
 sg13g2_fill_2 FILLER_75_2272 ();
 sg13g2_decap_8 FILLER_75_2312 ();
 sg13g2_decap_8 FILLER_75_2319 ();
 sg13g2_fill_1 FILLER_75_2326 ();
 sg13g2_decap_8 FILLER_75_2330 ();
 sg13g2_decap_8 FILLER_75_2337 ();
 sg13g2_decap_8 FILLER_75_2344 ();
 sg13g2_decap_4 FILLER_75_2351 ();
 sg13g2_fill_2 FILLER_75_2384 ();
 sg13g2_fill_1 FILLER_75_2386 ();
 sg13g2_fill_1 FILLER_75_2390 ();
 sg13g2_fill_2 FILLER_75_2416 ();
 sg13g2_fill_1 FILLER_75_2453 ();
 sg13g2_decap_8 FILLER_75_2465 ();
 sg13g2_decap_8 FILLER_75_2472 ();
 sg13g2_decap_4 FILLER_75_2479 ();
 sg13g2_fill_1 FILLER_75_2483 ();
 sg13g2_decap_8 FILLER_75_2492 ();
 sg13g2_fill_2 FILLER_75_2499 ();
 sg13g2_fill_2 FILLER_75_2527 ();
 sg13g2_fill_1 FILLER_75_2533 ();
 sg13g2_decap_4 FILLER_75_2546 ();
 sg13g2_fill_1 FILLER_75_2550 ();
 sg13g2_decap_8 FILLER_75_2585 ();
 sg13g2_decap_8 FILLER_75_2592 ();
 sg13g2_decap_8 FILLER_75_2599 ();
 sg13g2_decap_8 FILLER_75_2606 ();
 sg13g2_decap_8 FILLER_75_2613 ();
 sg13g2_decap_8 FILLER_75_2620 ();
 sg13g2_decap_8 FILLER_75_2627 ();
 sg13g2_decap_8 FILLER_75_2634 ();
 sg13g2_decap_8 FILLER_75_2641 ();
 sg13g2_decap_8 FILLER_75_2648 ();
 sg13g2_decap_8 FILLER_75_2655 ();
 sg13g2_decap_8 FILLER_75_2662 ();
 sg13g2_fill_1 FILLER_75_2669 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_7 ();
 sg13g2_fill_2 FILLER_76_13 ();
 sg13g2_fill_1 FILLER_76_15 ();
 sg13g2_fill_2 FILLER_76_30 ();
 sg13g2_fill_1 FILLER_76_58 ();
 sg13g2_fill_1 FILLER_76_68 ();
 sg13g2_fill_1 FILLER_76_78 ();
 sg13g2_fill_2 FILLER_76_83 ();
 sg13g2_fill_1 FILLER_76_96 ();
 sg13g2_fill_1 FILLER_76_103 ();
 sg13g2_decap_4 FILLER_76_114 ();
 sg13g2_fill_1 FILLER_76_129 ();
 sg13g2_fill_1 FILLER_76_158 ();
 sg13g2_fill_2 FILLER_76_165 ();
 sg13g2_fill_1 FILLER_76_176 ();
 sg13g2_decap_4 FILLER_76_182 ();
 sg13g2_fill_2 FILLER_76_191 ();
 sg13g2_fill_2 FILLER_76_201 ();
 sg13g2_decap_4 FILLER_76_215 ();
 sg13g2_fill_1 FILLER_76_238 ();
 sg13g2_fill_2 FILLER_76_243 ();
 sg13g2_decap_8 FILLER_76_288 ();
 sg13g2_decap_4 FILLER_76_295 ();
 sg13g2_decap_4 FILLER_76_340 ();
 sg13g2_fill_2 FILLER_76_344 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_fill_2 FILLER_76_357 ();
 sg13g2_decap_4 FILLER_76_414 ();
 sg13g2_decap_8 FILLER_76_425 ();
 sg13g2_fill_2 FILLER_76_442 ();
 sg13g2_fill_1 FILLER_76_444 ();
 sg13g2_decap_8 FILLER_76_451 ();
 sg13g2_decap_8 FILLER_76_458 ();
 sg13g2_decap_4 FILLER_76_465 ();
 sg13g2_fill_1 FILLER_76_469 ();
 sg13g2_fill_2 FILLER_76_515 ();
 sg13g2_fill_2 FILLER_76_521 ();
 sg13g2_fill_1 FILLER_76_567 ();
 sg13g2_decap_8 FILLER_76_575 ();
 sg13g2_fill_2 FILLER_76_582 ();
 sg13g2_fill_1 FILLER_76_584 ();
 sg13g2_decap_4 FILLER_76_590 ();
 sg13g2_fill_1 FILLER_76_607 ();
 sg13g2_decap_4 FILLER_76_621 ();
 sg13g2_fill_1 FILLER_76_625 ();
 sg13g2_fill_2 FILLER_76_631 ();
 sg13g2_fill_2 FILLER_76_664 ();
 sg13g2_fill_2 FILLER_76_676 ();
 sg13g2_fill_1 FILLER_76_689 ();
 sg13g2_decap_8 FILLER_76_694 ();
 sg13g2_decap_4 FILLER_76_701 ();
 sg13g2_fill_2 FILLER_76_705 ();
 sg13g2_decap_8 FILLER_76_711 ();
 sg13g2_decap_8 FILLER_76_718 ();
 sg13g2_decap_8 FILLER_76_725 ();
 sg13g2_fill_2 FILLER_76_732 ();
 sg13g2_fill_1 FILLER_76_734 ();
 sg13g2_decap_8 FILLER_76_752 ();
 sg13g2_fill_1 FILLER_76_759 ();
 sg13g2_decap_8 FILLER_76_772 ();
 sg13g2_decap_4 FILLER_76_779 ();
 sg13g2_decap_4 FILLER_76_817 ();
 sg13g2_fill_2 FILLER_76_821 ();
 sg13g2_decap_4 FILLER_76_831 ();
 sg13g2_fill_2 FILLER_76_835 ();
 sg13g2_decap_8 FILLER_76_853 ();
 sg13g2_decap_8 FILLER_76_860 ();
 sg13g2_decap_8 FILLER_76_867 ();
 sg13g2_decap_8 FILLER_76_874 ();
 sg13g2_decap_8 FILLER_76_881 ();
 sg13g2_decap_8 FILLER_76_888 ();
 sg13g2_decap_8 FILLER_76_895 ();
 sg13g2_fill_2 FILLER_76_902 ();
 sg13g2_fill_1 FILLER_76_908 ();
 sg13g2_fill_2 FILLER_76_935 ();
 sg13g2_fill_1 FILLER_76_937 ();
 sg13g2_decap_8 FILLER_76_964 ();
 sg13g2_fill_1 FILLER_76_971 ();
 sg13g2_decap_8 FILLER_76_976 ();
 sg13g2_decap_8 FILLER_76_983 ();
 sg13g2_decap_8 FILLER_76_990 ();
 sg13g2_decap_8 FILLER_76_997 ();
 sg13g2_decap_4 FILLER_76_1004 ();
 sg13g2_fill_1 FILLER_76_1008 ();
 sg13g2_fill_2 FILLER_76_1019 ();
 sg13g2_fill_1 FILLER_76_1021 ();
 sg13g2_decap_8 FILLER_76_1032 ();
 sg13g2_fill_1 FILLER_76_1039 ();
 sg13g2_decap_8 FILLER_76_1066 ();
 sg13g2_fill_2 FILLER_76_1073 ();
 sg13g2_fill_1 FILLER_76_1075 ();
 sg13g2_decap_8 FILLER_76_1138 ();
 sg13g2_decap_8 FILLER_76_1145 ();
 sg13g2_fill_1 FILLER_76_1152 ();
 sg13g2_fill_2 FILLER_76_1169 ();
 sg13g2_decap_4 FILLER_76_1179 ();
 sg13g2_fill_1 FILLER_76_1183 ();
 sg13g2_decap_8 FILLER_76_1193 ();
 sg13g2_decap_8 FILLER_76_1200 ();
 sg13g2_decap_8 FILLER_76_1207 ();
 sg13g2_decap_8 FILLER_76_1214 ();
 sg13g2_decap_8 FILLER_76_1221 ();
 sg13g2_fill_1 FILLER_76_1228 ();
 sg13g2_decap_8 FILLER_76_1259 ();
 sg13g2_fill_2 FILLER_76_1266 ();
 sg13g2_fill_2 FILLER_76_1300 ();
 sg13g2_fill_1 FILLER_76_1302 ();
 sg13g2_decap_4 FILLER_76_1323 ();
 sg13g2_fill_1 FILLER_76_1327 ();
 sg13g2_fill_1 FILLER_76_1334 ();
 sg13g2_decap_8 FILLER_76_1380 ();
 sg13g2_fill_1 FILLER_76_1387 ();
 sg13g2_decap_8 FILLER_76_1392 ();
 sg13g2_fill_2 FILLER_76_1399 ();
 sg13g2_fill_1 FILLER_76_1401 ();
 sg13g2_fill_1 FILLER_76_1428 ();
 sg13g2_fill_2 FILLER_76_1451 ();
 sg13g2_decap_8 FILLER_76_1460 ();
 sg13g2_decap_8 FILLER_76_1467 ();
 sg13g2_decap_8 FILLER_76_1474 ();
 sg13g2_fill_2 FILLER_76_1481 ();
 sg13g2_fill_1 FILLER_76_1483 ();
 sg13g2_decap_8 FILLER_76_1493 ();
 sg13g2_decap_4 FILLER_76_1500 ();
 sg13g2_fill_2 FILLER_76_1504 ();
 sg13g2_decap_4 FILLER_76_1541 ();
 sg13g2_fill_1 FILLER_76_1545 ();
 sg13g2_decap_8 FILLER_76_1551 ();
 sg13g2_decap_8 FILLER_76_1558 ();
 sg13g2_fill_2 FILLER_76_1565 ();
 sg13g2_fill_2 FILLER_76_1571 ();
 sg13g2_fill_1 FILLER_76_1573 ();
 sg13g2_fill_1 FILLER_76_1600 ();
 sg13g2_decap_8 FILLER_76_1627 ();
 sg13g2_decap_8 FILLER_76_1634 ();
 sg13g2_decap_4 FILLER_76_1641 ();
 sg13g2_fill_1 FILLER_76_1645 ();
 sg13g2_fill_1 FILLER_76_1656 ();
 sg13g2_decap_4 FILLER_76_1722 ();
 sg13g2_fill_2 FILLER_76_1732 ();
 sg13g2_fill_1 FILLER_76_1734 ();
 sg13g2_fill_1 FILLER_76_1739 ();
 sg13g2_decap_8 FILLER_76_1748 ();
 sg13g2_fill_2 FILLER_76_1755 ();
 sg13g2_fill_1 FILLER_76_1757 ();
 sg13g2_fill_2 FILLER_76_1763 ();
 sg13g2_fill_2 FILLER_76_1795 ();
 sg13g2_fill_1 FILLER_76_1797 ();
 sg13g2_decap_4 FILLER_76_1809 ();
 sg13g2_fill_1 FILLER_76_1813 ();
 sg13g2_decap_8 FILLER_76_1844 ();
 sg13g2_decap_8 FILLER_76_1857 ();
 sg13g2_fill_2 FILLER_76_1864 ();
 sg13g2_decap_8 FILLER_76_1874 ();
 sg13g2_decap_8 FILLER_76_1881 ();
 sg13g2_decap_8 FILLER_76_1888 ();
 sg13g2_decap_8 FILLER_76_1895 ();
 sg13g2_decap_4 FILLER_76_1928 ();
 sg13g2_fill_1 FILLER_76_1932 ();
 sg13g2_decap_8 FILLER_76_1996 ();
 sg13g2_decap_8 FILLER_76_2003 ();
 sg13g2_fill_2 FILLER_76_2010 ();
 sg13g2_fill_2 FILLER_76_2026 ();
 sg13g2_decap_8 FILLER_76_2075 ();
 sg13g2_decap_8 FILLER_76_2087 ();
 sg13g2_decap_4 FILLER_76_2094 ();
 sg13g2_decap_8 FILLER_76_2114 ();
 sg13g2_decap_8 FILLER_76_2121 ();
 sg13g2_decap_8 FILLER_76_2128 ();
 sg13g2_decap_8 FILLER_76_2135 ();
 sg13g2_decap_4 FILLER_76_2142 ();
 sg13g2_fill_2 FILLER_76_2161 ();
 sg13g2_fill_1 FILLER_76_2163 ();
 sg13g2_decap_4 FILLER_76_2190 ();
 sg13g2_fill_2 FILLER_76_2194 ();
 sg13g2_fill_1 FILLER_76_2227 ();
 sg13g2_fill_2 FILLER_76_2237 ();
 sg13g2_fill_1 FILLER_76_2239 ();
 sg13g2_decap_8 FILLER_76_2274 ();
 sg13g2_decap_8 FILLER_76_2287 ();
 sg13g2_decap_8 FILLER_76_2294 ();
 sg13g2_decap_8 FILLER_76_2333 ();
 sg13g2_fill_1 FILLER_76_2340 ();
 sg13g2_decap_4 FILLER_76_2374 ();
 sg13g2_fill_1 FILLER_76_2382 ();
 sg13g2_fill_1 FILLER_76_2387 ();
 sg13g2_fill_2 FILLER_76_2399 ();
 sg13g2_fill_1 FILLER_76_2401 ();
 sg13g2_fill_2 FILLER_76_2406 ();
 sg13g2_decap_8 FILLER_76_2442 ();
 sg13g2_decap_8 FILLER_76_2449 ();
 sg13g2_fill_2 FILLER_76_2456 ();
 sg13g2_fill_2 FILLER_76_2484 ();
 sg13g2_fill_1 FILLER_76_2486 ();
 sg13g2_decap_8 FILLER_76_2523 ();
 sg13g2_decap_8 FILLER_76_2530 ();
 sg13g2_decap_8 FILLER_76_2537 ();
 sg13g2_fill_1 FILLER_76_2544 ();
 sg13g2_decap_8 FILLER_76_2549 ();
 sg13g2_decap_8 FILLER_76_2556 ();
 sg13g2_decap_8 FILLER_76_2563 ();
 sg13g2_decap_4 FILLER_76_2570 ();
 sg13g2_decap_8 FILLER_76_2604 ();
 sg13g2_decap_8 FILLER_76_2611 ();
 sg13g2_decap_8 FILLER_76_2618 ();
 sg13g2_decap_8 FILLER_76_2625 ();
 sg13g2_decap_8 FILLER_76_2632 ();
 sg13g2_decap_8 FILLER_76_2639 ();
 sg13g2_decap_8 FILLER_76_2646 ();
 sg13g2_decap_8 FILLER_76_2653 ();
 sg13g2_decap_8 FILLER_76_2660 ();
 sg13g2_fill_2 FILLER_76_2667 ();
 sg13g2_fill_1 FILLER_76_2669 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_7 ();
 sg13g2_decap_4 FILLER_77_27 ();
 sg13g2_fill_2 FILLER_77_31 ();
 sg13g2_fill_1 FILLER_77_46 ();
 sg13g2_fill_2 FILLER_77_56 ();
 sg13g2_fill_1 FILLER_77_63 ();
 sg13g2_fill_1 FILLER_77_73 ();
 sg13g2_fill_1 FILLER_77_78 ();
 sg13g2_fill_1 FILLER_77_120 ();
 sg13g2_fill_1 FILLER_77_134 ();
 sg13g2_fill_2 FILLER_77_144 ();
 sg13g2_fill_2 FILLER_77_167 ();
 sg13g2_fill_1 FILLER_77_174 ();
 sg13g2_fill_1 FILLER_77_180 ();
 sg13g2_fill_2 FILLER_77_186 ();
 sg13g2_fill_2 FILLER_77_192 ();
 sg13g2_fill_1 FILLER_77_202 ();
 sg13g2_fill_1 FILLER_77_211 ();
 sg13g2_fill_1 FILLER_77_217 ();
 sg13g2_fill_2 FILLER_77_228 ();
 sg13g2_fill_1 FILLER_77_236 ();
 sg13g2_decap_4 FILLER_77_250 ();
 sg13g2_fill_1 FILLER_77_272 ();
 sg13g2_fill_1 FILLER_77_278 ();
 sg13g2_fill_1 FILLER_77_284 ();
 sg13g2_fill_1 FILLER_77_293 ();
 sg13g2_decap_8 FILLER_77_297 ();
 sg13g2_decap_8 FILLER_77_304 ();
 sg13g2_decap_4 FILLER_77_311 ();
 sg13g2_fill_1 FILLER_77_315 ();
 sg13g2_fill_2 FILLER_77_352 ();
 sg13g2_fill_2 FILLER_77_364 ();
 sg13g2_fill_1 FILLER_77_366 ();
 sg13g2_decap_8 FILLER_77_375 ();
 sg13g2_decap_8 FILLER_77_382 ();
 sg13g2_fill_2 FILLER_77_389 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_413 ();
 sg13g2_fill_1 FILLER_77_445 ();
 sg13g2_decap_8 FILLER_77_517 ();
 sg13g2_decap_8 FILLER_77_524 ();
 sg13g2_decap_4 FILLER_77_531 ();
 sg13g2_fill_1 FILLER_77_535 ();
 sg13g2_fill_1 FILLER_77_539 ();
 sg13g2_fill_2 FILLER_77_545 ();
 sg13g2_decap_8 FILLER_77_552 ();
 sg13g2_decap_4 FILLER_77_559 ();
 sg13g2_fill_2 FILLER_77_563 ();
 sg13g2_decap_4 FILLER_77_591 ();
 sg13g2_decap_8 FILLER_77_599 ();
 sg13g2_fill_2 FILLER_77_606 ();
 sg13g2_fill_2 FILLER_77_616 ();
 sg13g2_fill_2 FILLER_77_653 ();
 sg13g2_fill_1 FILLER_77_655 ();
 sg13g2_fill_2 FILLER_77_683 ();
 sg13g2_decap_8 FILLER_77_688 ();
 sg13g2_decap_8 FILLER_77_695 ();
 sg13g2_decap_8 FILLER_77_702 ();
 sg13g2_decap_8 FILLER_77_709 ();
 sg13g2_decap_8 FILLER_77_716 ();
 sg13g2_fill_2 FILLER_77_723 ();
 sg13g2_decap_4 FILLER_77_785 ();
 sg13g2_fill_1 FILLER_77_789 ();
 sg13g2_decap_8 FILLER_77_816 ();
 sg13g2_decap_8 FILLER_77_823 ();
 sg13g2_fill_2 FILLER_77_830 ();
 sg13g2_fill_1 FILLER_77_866 ();
 sg13g2_fill_1 FILLER_77_901 ();
 sg13g2_decap_8 FILLER_77_932 ();
 sg13g2_decap_8 FILLER_77_939 ();
 sg13g2_decap_8 FILLER_77_946 ();
 sg13g2_decap_8 FILLER_77_953 ();
 sg13g2_fill_2 FILLER_77_960 ();
 sg13g2_fill_1 FILLER_77_970 ();
 sg13g2_fill_2 FILLER_77_1023 ();
 sg13g2_fill_1 FILLER_77_1025 ();
 sg13g2_decap_4 FILLER_77_1052 ();
 sg13g2_fill_2 FILLER_77_1056 ();
 sg13g2_decap_8 FILLER_77_1084 ();
 sg13g2_decap_4 FILLER_77_1102 ();
 sg13g2_fill_2 FILLER_77_1106 ();
 sg13g2_decap_4 FILLER_77_1112 ();
 sg13g2_fill_1 FILLER_77_1116 ();
 sg13g2_decap_4 FILLER_77_1143 ();
 sg13g2_fill_1 FILLER_77_1156 ();
 sg13g2_fill_1 FILLER_77_1183 ();
 sg13g2_fill_1 FILLER_77_1210 ();
 sg13g2_fill_1 FILLER_77_1221 ();
 sg13g2_fill_2 FILLER_77_1227 ();
 sg13g2_decap_4 FILLER_77_1255 ();
 sg13g2_decap_8 FILLER_77_1271 ();
 sg13g2_decap_8 FILLER_77_1278 ();
 sg13g2_fill_2 FILLER_77_1285 ();
 sg13g2_decap_8 FILLER_77_1343 ();
 sg13g2_decap_8 FILLER_77_1350 ();
 sg13g2_decap_8 FILLER_77_1361 ();
 sg13g2_decap_8 FILLER_77_1398 ();
 sg13g2_fill_1 FILLER_77_1405 ();
 sg13g2_decap_4 FILLER_77_1414 ();
 sg13g2_fill_1 FILLER_77_1422 ();
 sg13g2_decap_8 FILLER_77_1449 ();
 sg13g2_decap_8 FILLER_77_1456 ();
 sg13g2_decap_4 FILLER_77_1463 ();
 sg13g2_fill_1 FILLER_77_1467 ();
 sg13g2_decap_8 FILLER_77_1512 ();
 sg13g2_decap_4 FILLER_77_1519 ();
 sg13g2_decap_8 FILLER_77_1527 ();
 sg13g2_decap_4 FILLER_77_1534 ();
 sg13g2_fill_1 FILLER_77_1542 ();
 sg13g2_decap_8 FILLER_77_1569 ();
 sg13g2_decap_8 FILLER_77_1576 ();
 sg13g2_decap_4 FILLER_77_1583 ();
 sg13g2_decap_8 FILLER_77_1590 ();
 sg13g2_decap_8 FILLER_77_1601 ();
 sg13g2_fill_2 FILLER_77_1608 ();
 sg13g2_fill_2 FILLER_77_1625 ();
 sg13g2_decap_8 FILLER_77_1637 ();
 sg13g2_decap_8 FILLER_77_1677 ();
 sg13g2_decap_4 FILLER_77_1684 ();
 sg13g2_fill_2 FILLER_77_1694 ();
 sg13g2_fill_1 FILLER_77_1747 ();
 sg13g2_fill_1 FILLER_77_1792 ();
 sg13g2_fill_1 FILLER_77_1804 ();
 sg13g2_fill_1 FILLER_77_1810 ();
 sg13g2_decap_8 FILLER_77_1846 ();
 sg13g2_fill_1 FILLER_77_1853 ();
 sg13g2_decap_4 FILLER_77_1863 ();
 sg13g2_fill_1 FILLER_77_1867 ();
 sg13g2_decap_4 FILLER_77_1872 ();
 sg13g2_fill_2 FILLER_77_1876 ();
 sg13g2_decap_8 FILLER_77_1882 ();
 sg13g2_fill_1 FILLER_77_1889 ();
 sg13g2_decap_4 FILLER_77_1920 ();
 sg13g2_decap_8 FILLER_77_1936 ();
 sg13g2_fill_2 FILLER_77_1943 ();
 sg13g2_fill_1 FILLER_77_1945 ();
 sg13g2_fill_2 FILLER_77_1964 ();
 sg13g2_fill_1 FILLER_77_1966 ();
 sg13g2_fill_1 FILLER_77_1971 ();
 sg13g2_fill_2 FILLER_77_2029 ();
 sg13g2_fill_1 FILLER_77_2060 ();
 sg13g2_decap_4 FILLER_77_2066 ();
 sg13g2_fill_1 FILLER_77_2070 ();
 sg13g2_decap_4 FILLER_77_2075 ();
 sg13g2_fill_1 FILLER_77_2079 ();
 sg13g2_fill_1 FILLER_77_2110 ();
 sg13g2_fill_2 FILLER_77_2115 ();
 sg13g2_fill_2 FILLER_77_2122 ();
 sg13g2_fill_2 FILLER_77_2150 ();
 sg13g2_fill_1 FILLER_77_2152 ();
 sg13g2_decap_8 FILLER_77_2179 ();
 sg13g2_fill_2 FILLER_77_2186 ();
 sg13g2_decap_4 FILLER_77_2193 ();
 sg13g2_fill_2 FILLER_77_2223 ();
 sg13g2_fill_1 FILLER_77_2225 ();
 sg13g2_decap_4 FILLER_77_2295 ();
 sg13g2_fill_2 FILLER_77_2304 ();
 sg13g2_fill_1 FILLER_77_2306 ();
 sg13g2_fill_2 FILLER_77_2333 ();
 sg13g2_fill_1 FILLER_77_2335 ();
 sg13g2_fill_1 FILLER_77_2367 ();
 sg13g2_decap_8 FILLER_77_2379 ();
 sg13g2_decap_4 FILLER_77_2386 ();
 sg13g2_fill_1 FILLER_77_2390 ();
 sg13g2_decap_4 FILLER_77_2394 ();
 sg13g2_fill_1 FILLER_77_2398 ();
 sg13g2_fill_1 FILLER_77_2404 ();
 sg13g2_decap_8 FILLER_77_2420 ();
 sg13g2_decap_4 FILLER_77_2427 ();
 sg13g2_fill_2 FILLER_77_2431 ();
 sg13g2_decap_8 FILLER_77_2489 ();
 sg13g2_fill_2 FILLER_77_2496 ();
 sg13g2_fill_1 FILLER_77_2498 ();
 sg13g2_decap_8 FILLER_77_2507 ();
 sg13g2_decap_8 FILLER_77_2514 ();
 sg13g2_decap_8 FILLER_77_2521 ();
 sg13g2_decap_8 FILLER_77_2528 ();
 sg13g2_fill_1 FILLER_77_2535 ();
 sg13g2_decap_8 FILLER_77_2575 ();
 sg13g2_fill_2 FILLER_77_2582 ();
 sg13g2_fill_1 FILLER_77_2584 ();
 sg13g2_decap_8 FILLER_77_2589 ();
 sg13g2_decap_8 FILLER_77_2596 ();
 sg13g2_decap_8 FILLER_77_2603 ();
 sg13g2_decap_8 FILLER_77_2610 ();
 sg13g2_decap_8 FILLER_77_2617 ();
 sg13g2_decap_8 FILLER_77_2624 ();
 sg13g2_decap_8 FILLER_77_2631 ();
 sg13g2_decap_8 FILLER_77_2638 ();
 sg13g2_decap_8 FILLER_77_2645 ();
 sg13g2_decap_8 FILLER_77_2652 ();
 sg13g2_decap_8 FILLER_77_2659 ();
 sg13g2_decap_4 FILLER_77_2666 ();
 sg13g2_decap_4 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_4 ();
 sg13g2_fill_1 FILLER_78_45 ();
 sg13g2_fill_1 FILLER_78_51 ();
 sg13g2_decap_8 FILLER_78_60 ();
 sg13g2_fill_2 FILLER_78_67 ();
 sg13g2_fill_1 FILLER_78_69 ();
 sg13g2_fill_2 FILLER_78_74 ();
 sg13g2_decap_4 FILLER_78_80 ();
 sg13g2_fill_1 FILLER_78_84 ();
 sg13g2_fill_1 FILLER_78_93 ();
 sg13g2_fill_1 FILLER_78_108 ();
 sg13g2_decap_8 FILLER_78_114 ();
 sg13g2_decap_8 FILLER_78_125 ();
 sg13g2_decap_8 FILLER_78_132 ();
 sg13g2_decap_8 FILLER_78_139 ();
 sg13g2_fill_1 FILLER_78_146 ();
 sg13g2_decap_8 FILLER_78_152 ();
 sg13g2_decap_8 FILLER_78_159 ();
 sg13g2_fill_2 FILLER_78_166 ();
 sg13g2_fill_1 FILLER_78_168 ();
 sg13g2_fill_1 FILLER_78_174 ();
 sg13g2_fill_1 FILLER_78_184 ();
 sg13g2_fill_1 FILLER_78_190 ();
 sg13g2_fill_2 FILLER_78_226 ();
 sg13g2_decap_4 FILLER_78_277 ();
 sg13g2_fill_1 FILLER_78_281 ();
 sg13g2_decap_8 FILLER_78_290 ();
 sg13g2_fill_2 FILLER_78_297 ();
 sg13g2_fill_2 FILLER_78_316 ();
 sg13g2_decap_4 FILLER_78_338 ();
 sg13g2_fill_1 FILLER_78_378 ();
 sg13g2_fill_1 FILLER_78_407 ();
 sg13g2_fill_1 FILLER_78_440 ();
 sg13g2_fill_1 FILLER_78_448 ();
 sg13g2_fill_2 FILLER_78_491 ();
 sg13g2_fill_1 FILLER_78_496 ();
 sg13g2_fill_2 FILLER_78_503 ();
 sg13g2_fill_1 FILLER_78_505 ();
 sg13g2_fill_2 FILLER_78_510 ();
 sg13g2_fill_1 FILLER_78_512 ();
 sg13g2_decap_8 FILLER_78_518 ();
 sg13g2_decap_8 FILLER_78_525 ();
 sg13g2_fill_2 FILLER_78_532 ();
 sg13g2_decap_4 FILLER_78_568 ();
 sg13g2_fill_1 FILLER_78_627 ();
 sg13g2_fill_1 FILLER_78_665 ();
 sg13g2_fill_2 FILLER_78_697 ();
 sg13g2_decap_8 FILLER_78_718 ();
 sg13g2_decap_8 FILLER_78_725 ();
 sg13g2_decap_4 FILLER_78_732 ();
 sg13g2_fill_2 FILLER_78_736 ();
 sg13g2_fill_2 FILLER_78_748 ();
 sg13g2_fill_2 FILLER_78_776 ();
 sg13g2_fill_1 FILLER_78_778 ();
 sg13g2_decap_4 FILLER_78_856 ();
 sg13g2_fill_2 FILLER_78_860 ();
 sg13g2_fill_1 FILLER_78_866 ();
 sg13g2_fill_1 FILLER_78_901 ();
 sg13g2_decap_8 FILLER_78_932 ();
 sg13g2_fill_2 FILLER_78_939 ();
 sg13g2_fill_1 FILLER_78_941 ();
 sg13g2_fill_2 FILLER_78_946 ();
 sg13g2_fill_1 FILLER_78_948 ();
 sg13g2_decap_8 FILLER_78_983 ();
 sg13g2_decap_4 FILLER_78_990 ();
 sg13g2_fill_1 FILLER_78_994 ();
 sg13g2_fill_1 FILLER_78_1005 ();
 sg13g2_fill_1 FILLER_78_1015 ();
 sg13g2_fill_1 FILLER_78_1046 ();
 sg13g2_fill_2 FILLER_78_1077 ();
 sg13g2_fill_2 FILLER_78_1091 ();
 sg13g2_fill_2 FILLER_78_1125 ();
 sg13g2_fill_1 FILLER_78_1127 ();
 sg13g2_fill_2 FILLER_78_1170 ();
 sg13g2_fill_1 FILLER_78_1172 ();
 sg13g2_decap_4 FILLER_78_1199 ();
 sg13g2_fill_1 FILLER_78_1203 ();
 sg13g2_decap_4 FILLER_78_1214 ();
 sg13g2_fill_2 FILLER_78_1218 ();
 sg13g2_fill_1 FILLER_78_1246 ();
 sg13g2_fill_2 FILLER_78_1251 ();
 sg13g2_fill_2 FILLER_78_1266 ();
 sg13g2_fill_1 FILLER_78_1268 ();
 sg13g2_decap_8 FILLER_78_1333 ();
 sg13g2_decap_4 FILLER_78_1370 ();
 sg13g2_decap_4 FILLER_78_1391 ();
 sg13g2_fill_1 FILLER_78_1395 ();
 sg13g2_decap_4 FILLER_78_1400 ();
 sg13g2_fill_1 FILLER_78_1404 ();
 sg13g2_decap_8 FILLER_78_1435 ();
 sg13g2_decap_8 FILLER_78_1442 ();
 sg13g2_decap_4 FILLER_78_1449 ();
 sg13g2_decap_8 FILLER_78_1457 ();
 sg13g2_fill_1 FILLER_78_1464 ();
 sg13g2_decap_8 FILLER_78_1513 ();
 sg13g2_decap_8 FILLER_78_1520 ();
 sg13g2_decap_8 FILLER_78_1527 ();
 sg13g2_fill_2 FILLER_78_1534 ();
 sg13g2_fill_1 FILLER_78_1536 ();
 sg13g2_fill_1 FILLER_78_1541 ();
 sg13g2_decap_8 FILLER_78_1568 ();
 sg13g2_fill_2 FILLER_78_1579 ();
 sg13g2_fill_2 FILLER_78_1585 ();
 sg13g2_fill_1 FILLER_78_1591 ();
 sg13g2_fill_1 FILLER_78_1605 ();
 sg13g2_fill_2 FILLER_78_1620 ();
 sg13g2_fill_1 FILLER_78_1652 ();
 sg13g2_decap_4 FILLER_78_1679 ();
 sg13g2_fill_2 FILLER_78_1683 ();
 sg13g2_decap_8 FILLER_78_1738 ();
 sg13g2_fill_2 FILLER_78_1745 ();
 sg13g2_decap_8 FILLER_78_1777 ();
 sg13g2_fill_2 FILLER_78_1784 ();
 sg13g2_decap_4 FILLER_78_1790 ();
 sg13g2_decap_4 FILLER_78_1829 ();
 sg13g2_decap_4 FILLER_78_1912 ();
 sg13g2_decap_4 FILLER_78_1921 ();
 sg13g2_decap_8 FILLER_78_1956 ();
 sg13g2_decap_8 FILLER_78_1963 ();
 sg13g2_decap_4 FILLER_78_1970 ();
 sg13g2_decap_4 FILLER_78_1998 ();
 sg13g2_fill_1 FILLER_78_2002 ();
 sg13g2_fill_2 FILLER_78_2057 ();
 sg13g2_fill_2 FILLER_78_2111 ();
 sg13g2_fill_1 FILLER_78_2113 ();
 sg13g2_decap_4 FILLER_78_2140 ();
 sg13g2_fill_1 FILLER_78_2144 ();
 sg13g2_decap_4 FILLER_78_2149 ();
 sg13g2_fill_1 FILLER_78_2153 ();
 sg13g2_fill_2 FILLER_78_2158 ();
 sg13g2_fill_1 FILLER_78_2160 ();
 sg13g2_decap_4 FILLER_78_2166 ();
 sg13g2_decap_4 FILLER_78_2174 ();
 sg13g2_fill_2 FILLER_78_2209 ();
 sg13g2_fill_1 FILLER_78_2211 ();
 sg13g2_fill_2 FILLER_78_2252 ();
 sg13g2_decap_8 FILLER_78_2297 ();
 sg13g2_decap_8 FILLER_78_2304 ();
 sg13g2_fill_1 FILLER_78_2311 ();
 sg13g2_fill_2 FILLER_78_2321 ();
 sg13g2_fill_1 FILLER_78_2336 ();
 sg13g2_fill_1 FILLER_78_2370 ();
 sg13g2_fill_2 FILLER_78_2405 ();
 sg13g2_fill_1 FILLER_78_2407 ();
 sg13g2_fill_2 FILLER_78_2411 ();
 sg13g2_fill_1 FILLER_78_2413 ();
 sg13g2_decap_8 FILLER_78_2440 ();
 sg13g2_decap_8 FILLER_78_2447 ();
 sg13g2_decap_8 FILLER_78_2454 ();
 sg13g2_decap_8 FILLER_78_2461 ();
 sg13g2_decap_8 FILLER_78_2468 ();
 sg13g2_decap_8 FILLER_78_2475 ();
 sg13g2_decap_8 FILLER_78_2572 ();
 sg13g2_decap_8 FILLER_78_2579 ();
 sg13g2_decap_8 FILLER_78_2586 ();
 sg13g2_decap_8 FILLER_78_2593 ();
 sg13g2_decap_8 FILLER_78_2600 ();
 sg13g2_decap_8 FILLER_78_2607 ();
 sg13g2_decap_8 FILLER_78_2614 ();
 sg13g2_decap_8 FILLER_78_2621 ();
 sg13g2_decap_8 FILLER_78_2628 ();
 sg13g2_decap_8 FILLER_78_2635 ();
 sg13g2_decap_8 FILLER_78_2642 ();
 sg13g2_decap_8 FILLER_78_2649 ();
 sg13g2_decap_8 FILLER_78_2656 ();
 sg13g2_decap_8 FILLER_78_2663 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_7 ();
 sg13g2_decap_4 FILLER_79_44 ();
 sg13g2_fill_1 FILLER_79_52 ();
 sg13g2_decap_8 FILLER_79_58 ();
 sg13g2_decap_8 FILLER_79_65 ();
 sg13g2_decap_8 FILLER_79_72 ();
 sg13g2_decap_8 FILLER_79_79 ();
 sg13g2_decap_4 FILLER_79_86 ();
 sg13g2_fill_1 FILLER_79_90 ();
 sg13g2_fill_2 FILLER_79_96 ();
 sg13g2_fill_1 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_103 ();
 sg13g2_decap_8 FILLER_79_110 ();
 sg13g2_decap_8 FILLER_79_117 ();
 sg13g2_decap_8 FILLER_79_124 ();
 sg13g2_decap_8 FILLER_79_131 ();
 sg13g2_decap_4 FILLER_79_138 ();
 sg13g2_fill_2 FILLER_79_142 ();
 sg13g2_decap_8 FILLER_79_148 ();
 sg13g2_decap_8 FILLER_79_155 ();
 sg13g2_decap_8 FILLER_79_162 ();
 sg13g2_decap_8 FILLER_79_169 ();
 sg13g2_decap_8 FILLER_79_176 ();
 sg13g2_decap_4 FILLER_79_183 ();
 sg13g2_fill_2 FILLER_79_187 ();
 sg13g2_fill_1 FILLER_79_238 ();
 sg13g2_fill_1 FILLER_79_243 ();
 sg13g2_decap_8 FILLER_79_263 ();
 sg13g2_decap_8 FILLER_79_270 ();
 sg13g2_fill_1 FILLER_79_285 ();
 sg13g2_fill_2 FILLER_79_316 ();
 sg13g2_fill_1 FILLER_79_318 ();
 sg13g2_fill_1 FILLER_79_323 ();
 sg13g2_fill_1 FILLER_79_343 ();
 sg13g2_fill_2 FILLER_79_368 ();
 sg13g2_fill_1 FILLER_79_370 ();
 sg13g2_fill_1 FILLER_79_397 ();
 sg13g2_fill_1 FILLER_79_411 ();
 sg13g2_fill_2 FILLER_79_436 ();
 sg13g2_fill_1 FILLER_79_438 ();
 sg13g2_fill_2 FILLER_79_444 ();
 sg13g2_fill_2 FILLER_79_452 ();
 sg13g2_decap_8 FILLER_79_483 ();
 sg13g2_decap_8 FILLER_79_490 ();
 sg13g2_decap_8 FILLER_79_497 ();
 sg13g2_decap_8 FILLER_79_504 ();
 sg13g2_fill_1 FILLER_79_511 ();
 sg13g2_fill_2 FILLER_79_538 ();
 sg13g2_fill_1 FILLER_79_540 ();
 sg13g2_decap_8 FILLER_79_580 ();
 sg13g2_fill_1 FILLER_79_587 ();
 sg13g2_decap_8 FILLER_79_601 ();
 sg13g2_fill_2 FILLER_79_608 ();
 sg13g2_fill_2 FILLER_79_631 ();
 sg13g2_fill_1 FILLER_79_633 ();
 sg13g2_fill_2 FILLER_79_638 ();
 sg13g2_fill_1 FILLER_79_640 ();
 sg13g2_decap_8 FILLER_79_646 ();
 sg13g2_fill_2 FILLER_79_653 ();
 sg13g2_decap_4 FILLER_79_690 ();
 sg13g2_fill_1 FILLER_79_694 ();
 sg13g2_fill_1 FILLER_79_707 ();
 sg13g2_fill_1 FILLER_79_713 ();
 sg13g2_fill_2 FILLER_79_753 ();
 sg13g2_fill_1 FILLER_79_755 ();
 sg13g2_decap_8 FILLER_79_760 ();
 sg13g2_fill_2 FILLER_79_767 ();
 sg13g2_fill_1 FILLER_79_769 ();
 sg13g2_fill_2 FILLER_79_774 ();
 sg13g2_decap_4 FILLER_79_786 ();
 sg13g2_fill_2 FILLER_79_790 ();
 sg13g2_decap_4 FILLER_79_800 ();
 sg13g2_decap_8 FILLER_79_808 ();
 sg13g2_fill_1 FILLER_79_815 ();
 sg13g2_fill_1 FILLER_79_820 ();
 sg13g2_fill_2 FILLER_79_847 ();
 sg13g2_fill_1 FILLER_79_853 ();
 sg13g2_decap_8 FILLER_79_884 ();
 sg13g2_decap_8 FILLER_79_891 ();
 sg13g2_fill_2 FILLER_79_898 ();
 sg13g2_fill_2 FILLER_79_904 ();
 sg13g2_fill_1 FILLER_79_936 ();
 sg13g2_fill_2 FILLER_79_980 ();
 sg13g2_fill_1 FILLER_79_982 ();
 sg13g2_decap_8 FILLER_79_1013 ();
 sg13g2_fill_2 FILLER_79_1020 ();
 sg13g2_fill_1 FILLER_79_1022 ();
 sg13g2_decap_4 FILLER_79_1027 ();
 sg13g2_fill_2 FILLER_79_1031 ();
 sg13g2_fill_1 FILLER_79_1068 ();
 sg13g2_decap_4 FILLER_79_1099 ();
 sg13g2_fill_1 FILLER_79_1103 ();
 sg13g2_decap_4 FILLER_79_1109 ();
 sg13g2_fill_1 FILLER_79_1124 ();
 sg13g2_decap_8 FILLER_79_1137 ();
 sg13g2_fill_1 FILLER_79_1144 ();
 sg13g2_decap_4 FILLER_79_1201 ();
 sg13g2_fill_1 FILLER_79_1205 ();
 sg13g2_decap_8 FILLER_79_1241 ();
 sg13g2_fill_1 FILLER_79_1248 ();
 sg13g2_fill_1 FILLER_79_1279 ();
 sg13g2_decap_8 FILLER_79_1306 ();
 sg13g2_fill_2 FILLER_79_1313 ();
 sg13g2_fill_2 FILLER_79_1345 ();
 sg13g2_fill_2 FILLER_79_1351 ();
 sg13g2_decap_4 FILLER_79_1379 ();
 sg13g2_fill_2 FILLER_79_1383 ();
 sg13g2_decap_8 FILLER_79_1505 ();
 sg13g2_fill_2 FILLER_79_1512 ();
 sg13g2_fill_1 FILLER_79_1518 ();
 sg13g2_fill_2 FILLER_79_1545 ();
 sg13g2_fill_2 FILLER_79_1551 ();
 sg13g2_fill_2 FILLER_79_1557 ();
 sg13g2_fill_1 FILLER_79_1559 ();
 sg13g2_fill_2 FILLER_79_1616 ();
 sg13g2_decap_8 FILLER_79_1644 ();
 sg13g2_fill_2 FILLER_79_1651 ();
 sg13g2_fill_1 FILLER_79_1653 ();
 sg13g2_fill_2 FILLER_79_1691 ();
 sg13g2_fill_1 FILLER_79_1693 ();
 sg13g2_fill_1 FILLER_79_1749 ();
 sg13g2_fill_2 FILLER_79_1780 ();
 sg13g2_fill_1 FILLER_79_1782 ();
 sg13g2_decap_8 FILLER_79_1809 ();
 sg13g2_fill_1 FILLER_79_1816 ();
 sg13g2_decap_8 FILLER_79_1825 ();
 sg13g2_decap_4 FILLER_79_1832 ();
 sg13g2_fill_2 FILLER_79_1836 ();
 sg13g2_fill_2 FILLER_79_1894 ();
 sg13g2_fill_1 FILLER_79_1896 ();
 sg13g2_decap_4 FILLER_79_1914 ();
 sg13g2_fill_1 FILLER_79_1918 ();
 sg13g2_decap_4 FILLER_79_1949 ();
 sg13g2_fill_2 FILLER_79_1953 ();
 sg13g2_fill_2 FILLER_79_1995 ();
 sg13g2_fill_1 FILLER_79_1997 ();
 sg13g2_decap_8 FILLER_79_2006 ();
 sg13g2_decap_4 FILLER_79_2013 ();
 sg13g2_decap_8 FILLER_79_2043 ();
 sg13g2_fill_1 FILLER_79_2050 ();
 sg13g2_fill_1 FILLER_79_2056 ();
 sg13g2_decap_8 FILLER_79_2070 ();
 sg13g2_fill_2 FILLER_79_2077 ();
 sg13g2_fill_1 FILLER_79_2079 ();
 sg13g2_fill_1 FILLER_79_2111 ();
 sg13g2_decap_4 FILLER_79_2129 ();
 sg13g2_fill_1 FILLER_79_2133 ();
 sg13g2_decap_4 FILLER_79_2139 ();
 sg13g2_fill_2 FILLER_79_2143 ();
 sg13g2_decap_4 FILLER_79_2197 ();
 sg13g2_decap_4 FILLER_79_2213 ();
 sg13g2_fill_1 FILLER_79_2217 ();
 sg13g2_decap_4 FILLER_79_2257 ();
 sg13g2_fill_1 FILLER_79_2261 ();
 sg13g2_decap_8 FILLER_79_2267 ();
 sg13g2_fill_2 FILLER_79_2274 ();
 sg13g2_fill_1 FILLER_79_2276 ();
 sg13g2_decap_8 FILLER_79_2281 ();
 sg13g2_decap_4 FILLER_79_2288 ();
 sg13g2_fill_2 FILLER_79_2292 ();
 sg13g2_fill_1 FILLER_79_2333 ();
 sg13g2_fill_2 FILLER_79_2339 ();
 sg13g2_fill_1 FILLER_79_2363 ();
 sg13g2_fill_1 FILLER_79_2368 ();
 sg13g2_fill_2 FILLER_79_2399 ();
 sg13g2_fill_1 FILLER_79_2401 ();
 sg13g2_fill_1 FILLER_79_2428 ();
 sg13g2_decap_8 FILLER_79_2442 ();
 sg13g2_fill_1 FILLER_79_2449 ();
 sg13g2_decap_8 FILLER_79_2454 ();
 sg13g2_fill_1 FILLER_79_2461 ();
 sg13g2_decap_4 FILLER_79_2492 ();
 sg13g2_decap_4 FILLER_79_2504 ();
 sg13g2_fill_1 FILLER_79_2508 ();
 sg13g2_decap_4 FILLER_79_2551 ();
 sg13g2_fill_1 FILLER_79_2555 ();
 sg13g2_decap_8 FILLER_79_2560 ();
 sg13g2_decap_8 FILLER_79_2567 ();
 sg13g2_decap_8 FILLER_79_2574 ();
 sg13g2_decap_8 FILLER_79_2581 ();
 sg13g2_decap_8 FILLER_79_2588 ();
 sg13g2_decap_8 FILLER_79_2595 ();
 sg13g2_decap_8 FILLER_79_2602 ();
 sg13g2_decap_8 FILLER_79_2609 ();
 sg13g2_decap_8 FILLER_79_2616 ();
 sg13g2_decap_8 FILLER_79_2623 ();
 sg13g2_decap_8 FILLER_79_2630 ();
 sg13g2_decap_8 FILLER_79_2637 ();
 sg13g2_decap_8 FILLER_79_2644 ();
 sg13g2_decap_8 FILLER_79_2651 ();
 sg13g2_decap_8 FILLER_79_2658 ();
 sg13g2_decap_4 FILLER_79_2665 ();
 sg13g2_fill_1 FILLER_79_2669 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_7 ();
 sg13g2_fill_1 FILLER_80_9 ();
 sg13g2_decap_4 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_22 ();
 sg13g2_decap_8 FILLER_80_29 ();
 sg13g2_decap_8 FILLER_80_36 ();
 sg13g2_decap_8 FILLER_80_43 ();
 sg13g2_decap_8 FILLER_80_50 ();
 sg13g2_decap_8 FILLER_80_57 ();
 sg13g2_decap_4 FILLER_80_64 ();
 sg13g2_fill_1 FILLER_80_68 ();
 sg13g2_fill_2 FILLER_80_93 ();
 sg13g2_fill_1 FILLER_80_95 ();
 sg13g2_fill_2 FILLER_80_112 ();
 sg13g2_fill_1 FILLER_80_114 ();
 sg13g2_decap_4 FILLER_80_139 ();
 sg13g2_fill_1 FILLER_80_143 ();
 sg13g2_decap_8 FILLER_80_148 ();
 sg13g2_decap_8 FILLER_80_155 ();
 sg13g2_decap_4 FILLER_80_162 ();
 sg13g2_fill_2 FILLER_80_170 ();
 sg13g2_fill_1 FILLER_80_172 ();
 sg13g2_decap_4 FILLER_80_177 ();
 sg13g2_fill_1 FILLER_80_181 ();
 sg13g2_fill_1 FILLER_80_189 ();
 sg13g2_fill_1 FILLER_80_198 ();
 sg13g2_fill_2 FILLER_80_228 ();
 sg13g2_fill_1 FILLER_80_238 ();
 sg13g2_decap_4 FILLER_80_246 ();
 sg13g2_fill_2 FILLER_80_250 ();
 sg13g2_fill_2 FILLER_80_260 ();
 sg13g2_decap_8 FILLER_80_265 ();
 sg13g2_decap_8 FILLER_80_272 ();
 sg13g2_decap_4 FILLER_80_279 ();
 sg13g2_fill_2 FILLER_80_283 ();
 sg13g2_decap_8 FILLER_80_289 ();
 sg13g2_decap_8 FILLER_80_296 ();
 sg13g2_decap_8 FILLER_80_303 ();
 sg13g2_decap_8 FILLER_80_310 ();
 sg13g2_decap_8 FILLER_80_317 ();
 sg13g2_decap_8 FILLER_80_324 ();
 sg13g2_decap_4 FILLER_80_331 ();
 sg13g2_fill_2 FILLER_80_335 ();
 sg13g2_fill_1 FILLER_80_341 ();
 sg13g2_decap_4 FILLER_80_346 ();
 sg13g2_decap_8 FILLER_80_358 ();
 sg13g2_decap_8 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_372 ();
 sg13g2_decap_4 FILLER_80_381 ();
 sg13g2_decap_4 FILLER_80_389 ();
 sg13g2_decap_4 FILLER_80_397 ();
 sg13g2_decap_8 FILLER_80_405 ();
 sg13g2_decap_8 FILLER_80_412 ();
 sg13g2_fill_2 FILLER_80_419 ();
 sg13g2_fill_2 FILLER_80_426 ();
 sg13g2_fill_1 FILLER_80_432 ();
 sg13g2_decap_8 FILLER_80_438 ();
 sg13g2_fill_1 FILLER_80_445 ();
 sg13g2_decap_8 FILLER_80_452 ();
 sg13g2_decap_8 FILLER_80_459 ();
 sg13g2_decap_8 FILLER_80_466 ();
 sg13g2_decap_8 FILLER_80_473 ();
 sg13g2_decap_8 FILLER_80_480 ();
 sg13g2_decap_8 FILLER_80_487 ();
 sg13g2_decap_8 FILLER_80_494 ();
 sg13g2_decap_8 FILLER_80_501 ();
 sg13g2_decap_8 FILLER_80_508 ();
 sg13g2_decap_8 FILLER_80_515 ();
 sg13g2_decap_8 FILLER_80_522 ();
 sg13g2_decap_8 FILLER_80_529 ();
 sg13g2_decap_4 FILLER_80_536 ();
 sg13g2_fill_2 FILLER_80_545 ();
 sg13g2_decap_8 FILLER_80_551 ();
 sg13g2_decap_8 FILLER_80_558 ();
 sg13g2_fill_2 FILLER_80_565 ();
 sg13g2_decap_8 FILLER_80_580 ();
 sg13g2_decap_8 FILLER_80_587 ();
 sg13g2_decap_8 FILLER_80_594 ();
 sg13g2_decap_8 FILLER_80_601 ();
 sg13g2_decap_8 FILLER_80_608 ();
 sg13g2_decap_8 FILLER_80_615 ();
 sg13g2_decap_8 FILLER_80_622 ();
 sg13g2_decap_8 FILLER_80_629 ();
 sg13g2_decap_8 FILLER_80_636 ();
 sg13g2_decap_8 FILLER_80_643 ();
 sg13g2_decap_8 FILLER_80_650 ();
 sg13g2_decap_8 FILLER_80_657 ();
 sg13g2_decap_8 FILLER_80_664 ();
 sg13g2_decap_8 FILLER_80_671 ();
 sg13g2_decap_8 FILLER_80_678 ();
 sg13g2_decap_8 FILLER_80_685 ();
 sg13g2_decap_8 FILLER_80_692 ();
 sg13g2_decap_8 FILLER_80_699 ();
 sg13g2_fill_1 FILLER_80_706 ();
 sg13g2_fill_2 FILLER_80_737 ();
 sg13g2_fill_1 FILLER_80_739 ();
 sg13g2_fill_2 FILLER_80_748 ();
 sg13g2_decap_4 FILLER_80_754 ();
 sg13g2_fill_1 FILLER_80_758 ();
 sg13g2_decap_8 FILLER_80_789 ();
 sg13g2_decap_8 FILLER_80_796 ();
 sg13g2_decap_8 FILLER_80_803 ();
 sg13g2_decap_8 FILLER_80_810 ();
 sg13g2_decap_8 FILLER_80_817 ();
 sg13g2_fill_2 FILLER_80_824 ();
 sg13g2_fill_1 FILLER_80_826 ();
 sg13g2_decap_8 FILLER_80_831 ();
 sg13g2_decap_8 FILLER_80_838 ();
 sg13g2_fill_2 FILLER_80_845 ();
 sg13g2_decap_8 FILLER_80_877 ();
 sg13g2_decap_8 FILLER_80_884 ();
 sg13g2_decap_8 FILLER_80_891 ();
 sg13g2_decap_8 FILLER_80_898 ();
 sg13g2_decap_4 FILLER_80_905 ();
 sg13g2_fill_1 FILLER_80_909 ();
 sg13g2_decap_8 FILLER_80_914 ();
 sg13g2_decap_8 FILLER_80_921 ();
 sg13g2_decap_8 FILLER_80_928 ();
 sg13g2_fill_1 FILLER_80_935 ();
 sg13g2_decap_8 FILLER_80_966 ();
 sg13g2_decap_8 FILLER_80_973 ();
 sg13g2_decap_8 FILLER_80_980 ();
 sg13g2_fill_2 FILLER_80_987 ();
 sg13g2_fill_1 FILLER_80_989 ();
 sg13g2_decap_8 FILLER_80_994 ();
 sg13g2_decap_8 FILLER_80_1001 ();
 sg13g2_decap_8 FILLER_80_1008 ();
 sg13g2_decap_8 FILLER_80_1015 ();
 sg13g2_fill_1 FILLER_80_1022 ();
 sg13g2_fill_2 FILLER_80_1031 ();
 sg13g2_fill_1 FILLER_80_1033 ();
 sg13g2_decap_4 FILLER_80_1059 ();
 sg13g2_decap_8 FILLER_80_1093 ();
 sg13g2_decap_8 FILLER_80_1100 ();
 sg13g2_decap_8 FILLER_80_1107 ();
 sg13g2_decap_4 FILLER_80_1114 ();
 sg13g2_fill_1 FILLER_80_1118 ();
 sg13g2_fill_2 FILLER_80_1122 ();
 sg13g2_decap_8 FILLER_80_1128 ();
 sg13g2_decap_8 FILLER_80_1135 ();
 sg13g2_decap_8 FILLER_80_1142 ();
 sg13g2_decap_8 FILLER_80_1149 ();
 sg13g2_decap_8 FILLER_80_1156 ();
 sg13g2_decap_4 FILLER_80_1163 ();
 sg13g2_fill_2 FILLER_80_1167 ();
 sg13g2_decap_4 FILLER_80_1173 ();
 sg13g2_decap_8 FILLER_80_1185 ();
 sg13g2_decap_8 FILLER_80_1192 ();
 sg13g2_decap_4 FILLER_80_1199 ();
 sg13g2_decap_8 FILLER_80_1233 ();
 sg13g2_decap_8 FILLER_80_1240 ();
 sg13g2_decap_8 FILLER_80_1247 ();
 sg13g2_decap_8 FILLER_80_1254 ();
 sg13g2_decap_8 FILLER_80_1261 ();
 sg13g2_decap_8 FILLER_80_1268 ();
 sg13g2_decap_4 FILLER_80_1275 ();
 sg13g2_fill_1 FILLER_80_1279 ();
 sg13g2_fill_2 FILLER_80_1284 ();
 sg13g2_fill_1 FILLER_80_1286 ();
 sg13g2_decap_8 FILLER_80_1291 ();
 sg13g2_decap_8 FILLER_80_1298 ();
 sg13g2_decap_8 FILLER_80_1305 ();
 sg13g2_decap_4 FILLER_80_1316 ();
 sg13g2_decap_8 FILLER_80_1328 ();
 sg13g2_decap_8 FILLER_80_1335 ();
 sg13g2_decap_8 FILLER_80_1342 ();
 sg13g2_decap_8 FILLER_80_1349 ();
 sg13g2_decap_4 FILLER_80_1356 ();
 sg13g2_fill_2 FILLER_80_1360 ();
 sg13g2_decap_8 FILLER_80_1366 ();
 sg13g2_decap_8 FILLER_80_1373 ();
 sg13g2_decap_8 FILLER_80_1380 ();
 sg13g2_decap_8 FILLER_80_1387 ();
 sg13g2_decap_8 FILLER_80_1394 ();
 sg13g2_decap_8 FILLER_80_1401 ();
 sg13g2_decap_4 FILLER_80_1408 ();
 sg13g2_decap_8 FILLER_80_1416 ();
 sg13g2_decap_8 FILLER_80_1427 ();
 sg13g2_decap_8 FILLER_80_1434 ();
 sg13g2_decap_8 FILLER_80_1441 ();
 sg13g2_decap_8 FILLER_80_1448 ();
 sg13g2_decap_8 FILLER_80_1455 ();
 sg13g2_decap_8 FILLER_80_1462 ();
 sg13g2_decap_8 FILLER_80_1469 ();
 sg13g2_fill_2 FILLER_80_1476 ();
 sg13g2_fill_1 FILLER_80_1478 ();
 sg13g2_fill_2 FILLER_80_1483 ();
 sg13g2_fill_1 FILLER_80_1485 ();
 sg13g2_decap_8 FILLER_80_1512 ();
 sg13g2_decap_4 FILLER_80_1519 ();
 sg13g2_fill_2 FILLER_80_1523 ();
 sg13g2_decap_8 FILLER_80_1529 ();
 sg13g2_decap_8 FILLER_80_1536 ();
 sg13g2_decap_8 FILLER_80_1543 ();
 sg13g2_decap_8 FILLER_80_1550 ();
 sg13g2_decap_8 FILLER_80_1557 ();
 sg13g2_decap_8 FILLER_80_1564 ();
 sg13g2_decap_8 FILLER_80_1575 ();
 sg13g2_decap_8 FILLER_80_1582 ();
 sg13g2_decap_4 FILLER_80_1589 ();
 sg13g2_decap_8 FILLER_80_1610 ();
 sg13g2_decap_8 FILLER_80_1617 ();
 sg13g2_decap_8 FILLER_80_1628 ();
 sg13g2_decap_8 FILLER_80_1635 ();
 sg13g2_decap_8 FILLER_80_1642 ();
 sg13g2_decap_8 FILLER_80_1649 ();
 sg13g2_decap_4 FILLER_80_1656 ();
 sg13g2_decap_8 FILLER_80_1664 ();
 sg13g2_decap_8 FILLER_80_1671 ();
 sg13g2_decap_8 FILLER_80_1678 ();
 sg13g2_fill_2 FILLER_80_1685 ();
 sg13g2_fill_1 FILLER_80_1687 ();
 sg13g2_decap_8 FILLER_80_1692 ();
 sg13g2_decap_8 FILLER_80_1699 ();
 sg13g2_decap_8 FILLER_80_1706 ();
 sg13g2_fill_2 FILLER_80_1713 ();
 sg13g2_decap_8 FILLER_80_1719 ();
 sg13g2_fill_1 FILLER_80_1726 ();
 sg13g2_decap_8 FILLER_80_1731 ();
 sg13g2_decap_4 FILLER_80_1738 ();
 sg13g2_fill_1 FILLER_80_1742 ();
 sg13g2_fill_1 FILLER_80_1756 ();
 sg13g2_decap_4 FILLER_80_1761 ();
 sg13g2_fill_1 FILLER_80_1765 ();
 sg13g2_decap_8 FILLER_80_1771 ();
 sg13g2_decap_4 FILLER_80_1778 ();
 sg13g2_fill_2 FILLER_80_1787 ();
 sg13g2_decap_8 FILLER_80_1793 ();
 sg13g2_decap_8 FILLER_80_1800 ();
 sg13g2_decap_8 FILLER_80_1807 ();
 sg13g2_decap_8 FILLER_80_1818 ();
 sg13g2_decap_8 FILLER_80_1825 ();
 sg13g2_decap_8 FILLER_80_1832 ();
 sg13g2_decap_8 FILLER_80_1839 ();
 sg13g2_decap_4 FILLER_80_1846 ();
 sg13g2_decap_8 FILLER_80_1855 ();
 sg13g2_decap_8 FILLER_80_1862 ();
 sg13g2_decap_8 FILLER_80_1869 ();
 sg13g2_decap_8 FILLER_80_1876 ();
 sg13g2_decap_8 FILLER_80_1883 ();
 sg13g2_decap_8 FILLER_80_1890 ();
 sg13g2_decap_8 FILLER_80_1897 ();
 sg13g2_decap_8 FILLER_80_1904 ();
 sg13g2_decap_8 FILLER_80_1911 ();
 sg13g2_decap_8 FILLER_80_1918 ();
 sg13g2_decap_8 FILLER_80_1925 ();
 sg13g2_decap_8 FILLER_80_1936 ();
 sg13g2_decap_8 FILLER_80_1943 ();
 sg13g2_decap_8 FILLER_80_1950 ();
 sg13g2_decap_8 FILLER_80_1957 ();
 sg13g2_decap_8 FILLER_80_1964 ();
 sg13g2_decap_8 FILLER_80_1971 ();
 sg13g2_decap_8 FILLER_80_1978 ();
 sg13g2_decap_8 FILLER_80_1985 ();
 sg13g2_fill_2 FILLER_80_1992 ();
 sg13g2_decap_8 FILLER_80_1998 ();
 sg13g2_decap_8 FILLER_80_2005 ();
 sg13g2_decap_8 FILLER_80_2012 ();
 sg13g2_decap_8 FILLER_80_2019 ();
 sg13g2_decap_8 FILLER_80_2026 ();
 sg13g2_decap_8 FILLER_80_2033 ();
 sg13g2_decap_8 FILLER_80_2040 ();
 sg13g2_decap_8 FILLER_80_2047 ();
 sg13g2_decap_8 FILLER_80_2054 ();
 sg13g2_decap_8 FILLER_80_2061 ();
 sg13g2_decap_8 FILLER_80_2068 ();
 sg13g2_decap_8 FILLER_80_2075 ();
 sg13g2_decap_8 FILLER_80_2087 ();
 sg13g2_decap_8 FILLER_80_2098 ();
 sg13g2_decap_4 FILLER_80_2105 ();
 sg13g2_fill_2 FILLER_80_2109 ();
 sg13g2_decap_8 FILLER_80_2119 ();
 sg13g2_decap_8 FILLER_80_2126 ();
 sg13g2_decap_8 FILLER_80_2133 ();
 sg13g2_fill_1 FILLER_80_2140 ();
 sg13g2_fill_2 FILLER_80_2149 ();
 sg13g2_fill_1 FILLER_80_2151 ();
 sg13g2_decap_4 FILLER_80_2156 ();
 sg13g2_fill_1 FILLER_80_2160 ();
 sg13g2_decap_8 FILLER_80_2169 ();
 sg13g2_decap_8 FILLER_80_2176 ();
 sg13g2_decap_8 FILLER_80_2183 ();
 sg13g2_decap_8 FILLER_80_2190 ();
 sg13g2_decap_8 FILLER_80_2197 ();
 sg13g2_decap_8 FILLER_80_2204 ();
 sg13g2_decap_8 FILLER_80_2211 ();
 sg13g2_decap_4 FILLER_80_2218 ();
 sg13g2_fill_1 FILLER_80_2222 ();
 sg13g2_decap_8 FILLER_80_2236 ();
 sg13g2_decap_8 FILLER_80_2243 ();
 sg13g2_decap_8 FILLER_80_2250 ();
 sg13g2_decap_8 FILLER_80_2257 ();
 sg13g2_decap_8 FILLER_80_2264 ();
 sg13g2_decap_8 FILLER_80_2271 ();
 sg13g2_decap_8 FILLER_80_2278 ();
 sg13g2_decap_8 FILLER_80_2285 ();
 sg13g2_decap_8 FILLER_80_2292 ();
 sg13g2_decap_8 FILLER_80_2299 ();
 sg13g2_decap_8 FILLER_80_2306 ();
 sg13g2_decap_8 FILLER_80_2313 ();
 sg13g2_decap_4 FILLER_80_2320 ();
 sg13g2_fill_2 FILLER_80_2324 ();
 sg13g2_decap_4 FILLER_80_2337 ();
 sg13g2_fill_1 FILLER_80_2344 ();
 sg13g2_decap_8 FILLER_80_2349 ();
 sg13g2_decap_8 FILLER_80_2356 ();
 sg13g2_decap_8 FILLER_80_2363 ();
 sg13g2_decap_4 FILLER_80_2370 ();
 sg13g2_decap_8 FILLER_80_2400 ();
 sg13g2_decap_8 FILLER_80_2407 ();
 sg13g2_decap_4 FILLER_80_2414 ();
 sg13g2_fill_1 FILLER_80_2418 ();
 sg13g2_fill_1 FILLER_80_2427 ();
 sg13g2_decap_8 FILLER_80_2438 ();
 sg13g2_decap_8 FILLER_80_2445 ();
 sg13g2_decap_8 FILLER_80_2452 ();
 sg13g2_decap_8 FILLER_80_2459 ();
 sg13g2_decap_8 FILLER_80_2466 ();
 sg13g2_decap_8 FILLER_80_2477 ();
 sg13g2_decap_8 FILLER_80_2484 ();
 sg13g2_decap_8 FILLER_80_2491 ();
 sg13g2_decap_8 FILLER_80_2498 ();
 sg13g2_decap_8 FILLER_80_2505 ();
 sg13g2_decap_8 FILLER_80_2512 ();
 sg13g2_fill_1 FILLER_80_2519 ();
 sg13g2_decap_8 FILLER_80_2528 ();
 sg13g2_fill_2 FILLER_80_2535 ();
 sg13g2_fill_1 FILLER_80_2537 ();
 sg13g2_decap_8 FILLER_80_2564 ();
 sg13g2_decap_8 FILLER_80_2571 ();
 sg13g2_decap_8 FILLER_80_2578 ();
 sg13g2_decap_8 FILLER_80_2585 ();
 sg13g2_decap_8 FILLER_80_2592 ();
 sg13g2_decap_8 FILLER_80_2599 ();
 sg13g2_decap_8 FILLER_80_2606 ();
 sg13g2_decap_8 FILLER_80_2613 ();
 sg13g2_decap_8 FILLER_80_2620 ();
 sg13g2_decap_8 FILLER_80_2627 ();
 sg13g2_decap_8 FILLER_80_2634 ();
 sg13g2_decap_8 FILLER_80_2641 ();
 sg13g2_decap_8 FILLER_80_2648 ();
 sg13g2_decap_8 FILLER_80_2655 ();
 sg13g2_decap_8 FILLER_80_2662 ();
 sg13g2_fill_1 FILLER_80_2669 ();
endmodule
