module tt_um_2048_vga_game (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire clknet_leaf_0_clk;
 wire net490;
 wire btn_down;
 wire \btn_down_debounce.button_sync_0 ;
 wire \btn_down_debounce.button_sync_1 ;
 wire \btn_down_debounce.debounce_counter[0] ;
 wire \btn_down_debounce.debounce_counter[10] ;
 wire \btn_down_debounce.debounce_counter[11] ;
 wire \btn_down_debounce.debounce_counter[12] ;
 wire \btn_down_debounce.debounce_counter[13] ;
 wire \btn_down_debounce.debounce_counter[14] ;
 wire \btn_down_debounce.debounce_counter[15] ;
 wire \btn_down_debounce.debounce_counter[16] ;
 wire \btn_down_debounce.debounce_counter[17] ;
 wire \btn_down_debounce.debounce_counter[1] ;
 wire \btn_down_debounce.debounce_counter[2] ;
 wire \btn_down_debounce.debounce_counter[3] ;
 wire \btn_down_debounce.debounce_counter[4] ;
 wire \btn_down_debounce.debounce_counter[5] ;
 wire \btn_down_debounce.debounce_counter[6] ;
 wire \btn_down_debounce.debounce_counter[7] ;
 wire \btn_down_debounce.debounce_counter[8] ;
 wire \btn_down_debounce.debounce_counter[9] ;
 wire btn_left;
 wire \btn_left_debounce.button_sync_0 ;
 wire \btn_left_debounce.button_sync_1 ;
 wire \btn_left_debounce.debounce_counter[0] ;
 wire \btn_left_debounce.debounce_counter[10] ;
 wire \btn_left_debounce.debounce_counter[11] ;
 wire \btn_left_debounce.debounce_counter[12] ;
 wire \btn_left_debounce.debounce_counter[13] ;
 wire \btn_left_debounce.debounce_counter[14] ;
 wire \btn_left_debounce.debounce_counter[15] ;
 wire \btn_left_debounce.debounce_counter[16] ;
 wire \btn_left_debounce.debounce_counter[17] ;
 wire \btn_left_debounce.debounce_counter[1] ;
 wire \btn_left_debounce.debounce_counter[2] ;
 wire \btn_left_debounce.debounce_counter[3] ;
 wire \btn_left_debounce.debounce_counter[4] ;
 wire \btn_left_debounce.debounce_counter[5] ;
 wire \btn_left_debounce.debounce_counter[6] ;
 wire \btn_left_debounce.debounce_counter[7] ;
 wire \btn_left_debounce.debounce_counter[8] ;
 wire \btn_left_debounce.debounce_counter[9] ;
 wire btn_right;
 wire \btn_right_debounce.button_sync_0 ;
 wire \btn_right_debounce.button_sync_1 ;
 wire \btn_right_debounce.debounce_counter[0] ;
 wire \btn_right_debounce.debounce_counter[10] ;
 wire \btn_right_debounce.debounce_counter[11] ;
 wire \btn_right_debounce.debounce_counter[12] ;
 wire \btn_right_debounce.debounce_counter[13] ;
 wire \btn_right_debounce.debounce_counter[14] ;
 wire \btn_right_debounce.debounce_counter[15] ;
 wire \btn_right_debounce.debounce_counter[16] ;
 wire \btn_right_debounce.debounce_counter[17] ;
 wire \btn_right_debounce.debounce_counter[1] ;
 wire \btn_right_debounce.debounce_counter[2] ;
 wire \btn_right_debounce.debounce_counter[3] ;
 wire \btn_right_debounce.debounce_counter[4] ;
 wire \btn_right_debounce.debounce_counter[5] ;
 wire \btn_right_debounce.debounce_counter[6] ;
 wire \btn_right_debounce.debounce_counter[7] ;
 wire \btn_right_debounce.debounce_counter[8] ;
 wire \btn_right_debounce.debounce_counter[9] ;
 wire btn_up;
 wire \btn_up_debounce.button_sync_0 ;
 wire \btn_up_debounce.button_sync_1 ;
 wire \btn_up_debounce.debounce_counter[0] ;
 wire \btn_up_debounce.debounce_counter[10] ;
 wire \btn_up_debounce.debounce_counter[11] ;
 wire \btn_up_debounce.debounce_counter[12] ;
 wire \btn_up_debounce.debounce_counter[13] ;
 wire \btn_up_debounce.debounce_counter[14] ;
 wire \btn_up_debounce.debounce_counter[15] ;
 wire \btn_up_debounce.debounce_counter[16] ;
 wire \btn_up_debounce.debounce_counter[17] ;
 wire \btn_up_debounce.debounce_counter[1] ;
 wire \btn_up_debounce.debounce_counter[2] ;
 wire \btn_up_debounce.debounce_counter[3] ;
 wire \btn_up_debounce.debounce_counter[4] ;
 wire \btn_up_debounce.debounce_counter[5] ;
 wire \btn_up_debounce.debounce_counter[6] ;
 wire \btn_up_debounce.debounce_counter[7] ;
 wire \btn_up_debounce.debounce_counter[8] ;
 wire \btn_up_debounce.debounce_counter[9] ;
 wire debug_btn_down;
 wire debug_btn_left;
 wire debug_btn_right;
 wire debug_btn_up;
 wire \debug_controller_inst.data_out_en ;
 wire \debug_controller_inst.grid_addr[0] ;
 wire \debug_controller_inst.grid_addr[1] ;
 wire \debug_controller_inst.grid_addr[2] ;
 wire \debug_controller_inst.grid_addr[3] ;
 wire \debug_controller_inst.grid_in[0] ;
 wire \debug_controller_inst.grid_in[10] ;
 wire \debug_controller_inst.grid_in[11] ;
 wire \debug_controller_inst.grid_in[12] ;
 wire \debug_controller_inst.grid_in[13] ;
 wire \debug_controller_inst.grid_in[14] ;
 wire \debug_controller_inst.grid_in[15] ;
 wire \debug_controller_inst.grid_in[16] ;
 wire \debug_controller_inst.grid_in[17] ;
 wire \debug_controller_inst.grid_in[18] ;
 wire \debug_controller_inst.grid_in[19] ;
 wire \debug_controller_inst.grid_in[1] ;
 wire \debug_controller_inst.grid_in[20] ;
 wire \debug_controller_inst.grid_in[21] ;
 wire \debug_controller_inst.grid_in[22] ;
 wire \debug_controller_inst.grid_in[23] ;
 wire \debug_controller_inst.grid_in[24] ;
 wire \debug_controller_inst.grid_in[25] ;
 wire \debug_controller_inst.grid_in[26] ;
 wire \debug_controller_inst.grid_in[27] ;
 wire \debug_controller_inst.grid_in[28] ;
 wire \debug_controller_inst.grid_in[29] ;
 wire \debug_controller_inst.grid_in[2] ;
 wire \debug_controller_inst.grid_in[30] ;
 wire \debug_controller_inst.grid_in[31] ;
 wire \debug_controller_inst.grid_in[32] ;
 wire \debug_controller_inst.grid_in[33] ;
 wire \debug_controller_inst.grid_in[34] ;
 wire \debug_controller_inst.grid_in[35] ;
 wire \debug_controller_inst.grid_in[36] ;
 wire \debug_controller_inst.grid_in[37] ;
 wire \debug_controller_inst.grid_in[38] ;
 wire \debug_controller_inst.grid_in[39] ;
 wire \debug_controller_inst.grid_in[3] ;
 wire \debug_controller_inst.grid_in[40] ;
 wire \debug_controller_inst.grid_in[41] ;
 wire \debug_controller_inst.grid_in[42] ;
 wire \debug_controller_inst.grid_in[43] ;
 wire \debug_controller_inst.grid_in[44] ;
 wire \debug_controller_inst.grid_in[45] ;
 wire \debug_controller_inst.grid_in[46] ;
 wire \debug_controller_inst.grid_in[47] ;
 wire \debug_controller_inst.grid_in[48] ;
 wire \debug_controller_inst.grid_in[49] ;
 wire \debug_controller_inst.grid_in[4] ;
 wire \debug_controller_inst.grid_in[50] ;
 wire \debug_controller_inst.grid_in[51] ;
 wire \debug_controller_inst.grid_in[52] ;
 wire \debug_controller_inst.grid_in[53] ;
 wire \debug_controller_inst.grid_in[54] ;
 wire \debug_controller_inst.grid_in[55] ;
 wire \debug_controller_inst.grid_in[56] ;
 wire \debug_controller_inst.grid_in[57] ;
 wire \debug_controller_inst.grid_in[58] ;
 wire \debug_controller_inst.grid_in[59] ;
 wire \debug_controller_inst.grid_in[5] ;
 wire \debug_controller_inst.grid_in[60] ;
 wire \debug_controller_inst.grid_in[61] ;
 wire \debug_controller_inst.grid_in[62] ;
 wire \debug_controller_inst.grid_in[63] ;
 wire \debug_controller_inst.grid_in[6] ;
 wire \debug_controller_inst.grid_in[7] ;
 wire \debug_controller_inst.grid_in[8] ;
 wire \debug_controller_inst.grid_in[9] ;
 wire \debug_controller_inst.grid_out_addr[0] ;
 wire \debug_controller_inst.grid_out_addr[1] ;
 wire \debug_controller_inst.grid_out_addr[2] ;
 wire \debug_controller_inst.grid_out_addr[3] ;
 wire \debug_controller_inst.grid_out_data[0] ;
 wire \debug_controller_inst.grid_out_data[1] ;
 wire \debug_controller_inst.grid_out_data[2] ;
 wire \debug_controller_inst.grid_out_data[3] ;
 wire \debug_controller_inst.grid_out_valid ;
 wire \draw_game_inst.board_x[0] ;
 wire \draw_game_inst.board_x[1] ;
 wire \draw_game_inst.board_x[2] ;
 wire \draw_game_inst.board_x[3] ;
 wire \draw_game_inst.board_x[4] ;
 wire \draw_game_inst.board_x[5] ;
 wire \draw_game_inst.board_y[0] ;
 wire \draw_game_inst.board_y[1] ;
 wire \draw_game_inst.board_y[2] ;
 wire \draw_game_inst.board_y[3] ;
 wire \draw_game_inst.board_y[4] ;
 wire \draw_game_inst.board_y[5] ;
 wire \draw_game_inst.board_y[6] ;
 wire \draw_game_inst.grid[0] ;
 wire \draw_game_inst.grid[10] ;
 wire \draw_game_inst.grid[11] ;
 wire \draw_game_inst.grid[12] ;
 wire \draw_game_inst.grid[13] ;
 wire \draw_game_inst.grid[14] ;
 wire \draw_game_inst.grid[15] ;
 wire \draw_game_inst.grid[16] ;
 wire \draw_game_inst.grid[17] ;
 wire \draw_game_inst.grid[18] ;
 wire \draw_game_inst.grid[19] ;
 wire \draw_game_inst.grid[1] ;
 wire \draw_game_inst.grid[20] ;
 wire \draw_game_inst.grid[21] ;
 wire \draw_game_inst.grid[22] ;
 wire \draw_game_inst.grid[23] ;
 wire \draw_game_inst.grid[24] ;
 wire \draw_game_inst.grid[25] ;
 wire \draw_game_inst.grid[26] ;
 wire \draw_game_inst.grid[27] ;
 wire \draw_game_inst.grid[28] ;
 wire \draw_game_inst.grid[29] ;
 wire \draw_game_inst.grid[2] ;
 wire \draw_game_inst.grid[30] ;
 wire \draw_game_inst.grid[31] ;
 wire \draw_game_inst.grid[32] ;
 wire \draw_game_inst.grid[33] ;
 wire \draw_game_inst.grid[34] ;
 wire \draw_game_inst.grid[35] ;
 wire \draw_game_inst.grid[36] ;
 wire \draw_game_inst.grid[37] ;
 wire \draw_game_inst.grid[38] ;
 wire \draw_game_inst.grid[39] ;
 wire \draw_game_inst.grid[3] ;
 wire \draw_game_inst.grid[40] ;
 wire \draw_game_inst.grid[41] ;
 wire \draw_game_inst.grid[42] ;
 wire \draw_game_inst.grid[43] ;
 wire \draw_game_inst.grid[44] ;
 wire \draw_game_inst.grid[45] ;
 wire \draw_game_inst.grid[46] ;
 wire \draw_game_inst.grid[47] ;
 wire \draw_game_inst.grid[48] ;
 wire \draw_game_inst.grid[49] ;
 wire \draw_game_inst.grid[4] ;
 wire \draw_game_inst.grid[50] ;
 wire \draw_game_inst.grid[51] ;
 wire \draw_game_inst.grid[52] ;
 wire \draw_game_inst.grid[53] ;
 wire \draw_game_inst.grid[54] ;
 wire \draw_game_inst.grid[55] ;
 wire \draw_game_inst.grid[56] ;
 wire \draw_game_inst.grid[57] ;
 wire \draw_game_inst.grid[58] ;
 wire \draw_game_inst.grid[59] ;
 wire \draw_game_inst.grid[5] ;
 wire \draw_game_inst.grid[60] ;
 wire \draw_game_inst.grid[61] ;
 wire \draw_game_inst.grid[62] ;
 wire \draw_game_inst.grid[63] ;
 wire \draw_game_inst.grid[6] ;
 wire \draw_game_inst.grid[7] ;
 wire \draw_game_inst.grid[8] ;
 wire \draw_game_inst.grid[9] ;
 wire \draw_game_inst.new_tiles[0] ;
 wire \draw_game_inst.new_tiles[10] ;
 wire \draw_game_inst.new_tiles[11] ;
 wire \draw_game_inst.new_tiles[12] ;
 wire \draw_game_inst.new_tiles[13] ;
 wire \draw_game_inst.new_tiles[14] ;
 wire \draw_game_inst.new_tiles[15] ;
 wire \draw_game_inst.new_tiles[1] ;
 wire \draw_game_inst.new_tiles[2] ;
 wire \draw_game_inst.new_tiles[3] ;
 wire \draw_game_inst.new_tiles[4] ;
 wire \draw_game_inst.new_tiles[5] ;
 wire \draw_game_inst.new_tiles[6] ;
 wire \draw_game_inst.new_tiles[7] ;
 wire \draw_game_inst.new_tiles[8] ;
 wire \draw_game_inst.new_tiles[9] ;
 wire \draw_game_inst.new_tiles_counter[0] ;
 wire \draw_game_inst.new_tiles_counter[1] ;
 wire \draw_game_inst.new_tiles_counter[2] ;
 wire \draw_game_inst.x[6] ;
 wire \draw_game_inst.x[7] ;
 wire \draw_game_inst.x[8] ;
 wire \draw_game_inst.x[9] ;
 wire \draw_game_inst.y[7] ;
 wire \draw_game_inst.y[8] ;
 wire \draw_game_inst.y[9] ;
 wire \game_logic_inst.add_new_tiles[0] ;
 wire \game_logic_inst.add_new_tiles[1] ;
 wire \game_logic_inst.added_tile_index[0] ;
 wire \game_logic_inst.added_tile_index[1] ;
 wire \game_logic_inst.added_tile_index[2] ;
 wire \game_logic_inst.added_tile_index[3] ;
 wire \game_logic_inst.calculate_move ;
 wire \game_logic_inst.current_direction[1] ;
 wire \game_logic_inst.current_direction[2] ;
 wire \game_logic_inst.current_direction[3] ;
 wire \game_logic_inst.current_row_index[0] ;
 wire \game_logic_inst.current_row_index[1] ;
 wire \game_logic_inst.debug_move_reg ;
 wire \game_logic_inst.game_started ;
 wire \game_logic_inst.lfsr_shift[0] ;
 wire \game_logic_inst.lfsr_shift[1] ;
 wire \game_logic_inst.lfsr_value[0] ;
 wire \game_logic_inst.lfsr_value[10] ;
 wire \game_logic_inst.lfsr_value[11] ;
 wire \game_logic_inst.lfsr_value[12] ;
 wire \game_logic_inst.lfsr_value[13] ;
 wire \game_logic_inst.lfsr_value[14] ;
 wire \game_logic_inst.lfsr_value[15] ;
 wire \game_logic_inst.lfsr_value[1] ;
 wire \game_logic_inst.lfsr_value[2] ;
 wire \game_logic_inst.lfsr_value[3] ;
 wire \game_logic_inst.lfsr_value[4] ;
 wire \game_logic_inst.lfsr_value[5] ;
 wire \game_logic_inst.lfsr_value[6] ;
 wire \game_logic_inst.lfsr_value[7] ;
 wire \game_logic_inst.lfsr_value[8] ;
 wire \game_logic_inst.lfsr_value[9] ;
 wire \game_logic_inst.prev_any_button_pressed ;
 wire \game_logic_inst.should_transpose ;
 wire \game_logic_inst.valid_move ;
 wire hsync;
 wire \lfsr_inst.lfsr[16] ;
 wire \lfsr_inst.lfsr[17] ;
 wire \lfsr_inst.lfsr[18] ;
 wire \lfsr_inst.lfsr[19] ;
 wire \lfsr_inst.lfsr[20] ;
 wire \lfsr_inst.lfsr[21] ;
 wire \lfsr_inst.lfsr[22] ;
 wire \lfsr_inst.lfsr[23] ;
 wire \lfsr_inst.lfsr[24] ;
 wire \lfsr_inst.lfsr[25] ;
 wire \lfsr_inst.lfsr[26] ;
 wire \lfsr_inst.lfsr[27] ;
 wire \lfsr_inst.lfsr[28] ;
 wire \lfsr_inst.lfsr[29] ;
 wire \lfsr_inst.lfsr[30] ;
 wire \lfsr_inst.lfsr[31] ;
 wire \new_tiles_counter[0] ;
 wire \new_tiles_counter[4] ;
 wire show_welcome_screen;
 wire \vga_sync_gen.vsync ;
 wire vsync_prev;
 wire \welcome_screen_grid[0] ;
 wire \welcome_screen_grid[11] ;
 wire \welcome_screen_grid[12] ;
 wire \welcome_screen_grid[16] ;
 wire \welcome_screen_grid[20] ;
 wire \welcome_screen_grid[24] ;
 wire \welcome_screen_grid[28] ;
 wire \welcome_screen_grid[32] ;
 wire \welcome_screen_grid[36] ;
 wire \welcome_screen_grid[40] ;
 wire \welcome_screen_grid[44] ;
 wire \welcome_screen_grid[48] ;
 wire \welcome_screen_grid[4] ;
 wire \welcome_screen_grid[52] ;
 wire \welcome_screen_grid[56] ;
 wire \welcome_screen_grid[60] ;
 wire \welcome_screen_inst.welcome_counter[0] ;
 wire \welcome_screen_inst.welcome_counter[1] ;
 wire \welcome_screen_inst.welcome_counter[2] ;
 wire \welcome_screen_inst.welcome_counter[3] ;
 wire \welcome_screen_inst.welcome_counter[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_dfrbp_1 \B[0]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net490),
    .D(_00171_),
    .Q_N(_05480_),
    .Q(net28));
 sg13g2_dfrbp_1 \B[1]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net491),
    .D(_00172_),
    .Q_N(_05479_),
    .Q(net24));
 sg13g2_dfrbp_1 \G[0]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net492),
    .D(_00173_),
    .Q_N(_05478_),
    .Q(net27));
 sg13g2_dfrbp_1 \G[1]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net493),
    .D(_00174_),
    .Q_N(_05477_),
    .Q(net23));
 sg13g2_dfrbp_1 \R[0]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net494),
    .D(_00175_),
    .Q_N(_05476_),
    .Q(net26));
 sg13g2_dfrbp_1 \R[1]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net495),
    .D(_00176_),
    .Q_N(_05475_),
    .Q(net22));
 sg13g2_buf_2 _05487_ (.A(rst_n),
    .X(_05057_));
 sg13g2_inv_1 _05488_ (.Y(_05058_),
    .A(_05057_));
 sg13g2_buf_1 _05489_ (.A(_05058_),
    .X(_05059_));
 sg13g2_buf_1 _05490_ (.A(_05059_),
    .X(_05060_));
 sg13g2_buf_1 _05491_ (.A(net413),
    .X(_05061_));
 sg13g2_buf_8 _05492_ (.A(\game_logic_inst.current_direction[3] ),
    .X(_05062_));
 sg13g2_buf_1 _05493_ (.A(\game_logic_inst.game_started ),
    .X(_05063_));
 sg13g2_buf_1 _05494_ (.A(show_welcome_screen),
    .X(_05064_));
 sg13g2_buf_1 _05495_ (.A(btn_right),
    .X(_05065_));
 sg13g2_buf_1 _05496_ (.A(btn_left),
    .X(_05066_));
 sg13g2_nor2_1 _05497_ (.A(_05065_),
    .B(_05066_),
    .Y(_05067_));
 sg13g2_nor2_1 _05498_ (.A(debug_btn_right),
    .B(debug_btn_left),
    .Y(_05068_));
 sg13g2_o21ai_1 _05499_ (.B1(_05068_),
    .Y(_05069_),
    .A1(_05064_),
    .A2(_05067_));
 sg13g2_buf_1 _05500_ (.A(btn_up),
    .X(_05070_));
 sg13g2_inv_1 _05501_ (.Y(_05071_),
    .A(show_welcome_screen));
 sg13g2_a21o_1 _05502_ (.A2(_05071_),
    .A1(_05070_),
    .B1(debug_btn_up),
    .X(_05072_));
 sg13g2_buf_1 _05503_ (.A(btn_down),
    .X(_05073_));
 sg13g2_a21oi_1 _05504_ (.A1(_05071_),
    .A2(_05073_),
    .Y(_05074_),
    .B1(debug_btn_down));
 sg13g2_nor2b_1 _05505_ (.A(_05072_),
    .B_N(_05074_),
    .Y(_05075_));
 sg13g2_nand2b_1 _05506_ (.Y(_05076_),
    .B(_05075_),
    .A_N(_05069_));
 sg13g2_nor2b_1 _05507_ (.A(\game_logic_inst.prev_any_button_pressed ),
    .B_N(_05076_),
    .Y(_05077_));
 sg13g2_buf_2 _05508_ (.A(_05077_),
    .X(_05078_));
 sg13g2_nand2_1 _05509_ (.Y(_05079_),
    .A(net480),
    .B(_05078_));
 sg13g2_buf_2 _05510_ (.A(_05079_),
    .X(_05080_));
 sg13g2_nor3_1 _05511_ (.A(_05069_),
    .B(_05072_),
    .C(_05080_),
    .Y(_05081_));
 sg13g2_a21oi_1 _05512_ (.A1(_05062_),
    .A2(_05080_),
    .Y(_05082_),
    .B1(_05081_));
 sg13g2_nor2_1 _05513_ (.A(net361),
    .B(_05082_),
    .Y(_00002_));
 sg13g2_buf_1 _05514_ (.A(\game_logic_inst.current_direction[2] ),
    .X(_05083_));
 sg13g2_nor2b_1 _05515_ (.A(_05064_),
    .B_N(_05066_),
    .Y(_05084_));
 sg13g2_a21oi_1 _05516_ (.A1(_05071_),
    .A2(_05065_),
    .Y(_05085_),
    .B1(debug_btn_right));
 sg13g2_nor4_1 _05517_ (.A(debug_btn_left),
    .B(_05080_),
    .C(_05084_),
    .D(_05085_),
    .Y(_05086_));
 sg13g2_a21oi_1 _05518_ (.A1(_05083_),
    .A2(_05080_),
    .Y(_05087_),
    .B1(_05086_));
 sg13g2_nor2_1 _05519_ (.A(net361),
    .B(_05087_),
    .Y(_00001_));
 sg13g2_nand2b_1 _05520_ (.Y(_05088_),
    .B(_05072_),
    .A_N(_05069_));
 sg13g2_nor2_1 _05521_ (.A(_05080_),
    .B(_05088_),
    .Y(_05089_));
 sg13g2_a21oi_1 _05522_ (.A1(\game_logic_inst.current_direction[1] ),
    .A2(_05080_),
    .Y(_05090_),
    .B1(_05089_));
 sg13g2_nor2_1 _05523_ (.A(net361),
    .B(_05090_),
    .Y(_00000_));
 sg13g2_buf_1 _05524_ (.A(\debug_controller_inst.grid_out_addr[3] ),
    .X(_05091_));
 sg13g2_inv_1 _05525_ (.Y(_05092_),
    .A(_05091_));
 sg13g2_buf_2 _05526_ (.A(\debug_controller_inst.grid_out_addr[2] ),
    .X(_05093_));
 sg13g2_buf_2 _05527_ (.A(\debug_controller_inst.grid_out_addr[1] ),
    .X(_05094_));
 sg13g2_buf_1 _05528_ (.A(\debug_controller_inst.grid_out_addr[0] ),
    .X(_05095_));
 sg13g2_nor3_1 _05529_ (.A(_05093_),
    .B(_05094_),
    .C(_05095_),
    .Y(_05096_));
 sg13g2_and4_1 _05530_ (.A(_05092_),
    .B(_00099_),
    .C(\debug_controller_inst.grid_out_valid ),
    .D(_05096_),
    .X(_05097_));
 sg13g2_buf_1 _05531_ (.A(_05097_),
    .X(_05098_));
 sg13g2_buf_1 _05532_ (.A(\game_logic_inst.calculate_move ),
    .X(_05099_));
 sg13g2_buf_1 _05533_ (.A(_05099_),
    .X(_05100_));
 sg13g2_buf_1 _05534_ (.A(net456),
    .X(_05101_));
 sg13g2_buf_1 _05535_ (.A(_05101_),
    .X(_05102_));
 sg13g2_buf_2 _05536_ (.A(\game_logic_inst.current_row_index[0] ),
    .X(_05103_));
 sg13g2_buf_8 _05537_ (.A(_05103_),
    .X(_05104_));
 sg13g2_buf_8 _05538_ (.A(net455),
    .X(_05105_));
 sg13g2_buf_8 _05539_ (.A(net411),
    .X(_05106_));
 sg13g2_buf_1 _05540_ (.A(net359),
    .X(_05107_));
 sg13g2_buf_8 _05541_ (.A(\game_logic_inst.current_row_index[1] ),
    .X(_05108_));
 sg13g2_buf_8 _05542_ (.A(_05108_),
    .X(_05109_));
 sg13g2_buf_8 _05543_ (.A(net454),
    .X(_05110_));
 sg13g2_buf_8 _05544_ (.A(net410),
    .X(_05111_));
 sg13g2_buf_8 _05545_ (.A(net358),
    .X(_05112_));
 sg13g2_buf_1 _05546_ (.A(_05112_),
    .X(_05113_));
 sg13g2_or2_1 _05547_ (.X(_05114_),
    .B(net161),
    .A(net262));
 sg13g2_buf_1 _05548_ (.A(_05114_),
    .X(_05115_));
 sg13g2_nor2_1 _05549_ (.A(_05062_),
    .B(_05083_),
    .Y(_05116_));
 sg13g2_buf_1 _05550_ (.A(_05116_),
    .X(_05117_));
 sg13g2_buf_1 _05551_ (.A(net409),
    .X(_05118_));
 sg13g2_buf_1 _05552_ (.A(_05118_),
    .X(_05119_));
 sg13g2_buf_1 _05553_ (.A(net260),
    .X(_05120_));
 sg13g2_buf_1 _05554_ (.A(_05120_),
    .X(_05121_));
 sg13g2_buf_2 _05555_ (.A(\debug_controller_inst.grid_in[17] ),
    .X(_05122_));
 sg13g2_buf_2 _05556_ (.A(\debug_controller_inst.grid_in[21] ),
    .X(_05123_));
 sg13g2_xor2_1 _05557_ (.B(_05123_),
    .A(_05122_),
    .X(_05124_));
 sg13g2_buf_2 _05558_ (.A(\debug_controller_inst.grid_in[29] ),
    .X(_05125_));
 sg13g2_buf_2 _05559_ (.A(\debug_controller_inst.grid_in[25] ),
    .X(_05126_));
 sg13g2_xor2_1 _05560_ (.B(_05126_),
    .A(_05125_),
    .X(_05127_));
 sg13g2_buf_2 _05561_ (.A(\debug_controller_inst.grid_in[49] ),
    .X(_05128_));
 sg13g2_buf_2 _05562_ (.A(\debug_controller_inst.grid_in[53] ),
    .X(_05129_));
 sg13g2_xor2_1 _05563_ (.B(_05129_),
    .A(_05128_),
    .X(_05130_));
 sg13g2_buf_2 _05564_ (.A(\debug_controller_inst.grid_in[61] ),
    .X(_05131_));
 sg13g2_buf_2 _05565_ (.A(\debug_controller_inst.grid_in[57] ),
    .X(_05132_));
 sg13g2_xor2_1 _05566_ (.B(_05132_),
    .A(_05131_),
    .X(_05133_));
 sg13g2_or2_1 _05567_ (.X(_05134_),
    .B(_05083_),
    .A(_05062_));
 sg13g2_buf_8 _05568_ (.A(_05134_),
    .X(_05135_));
 sg13g2_buf_8 _05569_ (.A(_05135_),
    .X(_05136_));
 sg13g2_mux4_1 _05570_ (.S0(net356),
    .A0(_05124_),
    .A1(_05127_),
    .A2(_05130_),
    .A3(_05133_),
    .S1(net358),
    .X(_05137_));
 sg13g2_inv_2 _05571_ (.Y(_05138_),
    .A(net455));
 sg13g2_buf_1 _05572_ (.A(_05138_),
    .X(_05139_));
 sg13g2_buf_8 _05573_ (.A(net410),
    .X(_05140_));
 sg13g2_buf_2 _05574_ (.A(\debug_controller_inst.grid_in[44] ),
    .X(_05141_));
 sg13g2_buf_2 _05575_ (.A(\debug_controller_inst.grid_in[40] ),
    .X(_05142_));
 sg13g2_xnor2_1 _05576_ (.Y(_05143_),
    .A(_05141_),
    .B(_05142_));
 sg13g2_buf_2 _05577_ (.A(\debug_controller_inst.grid_in[47] ),
    .X(_05144_));
 sg13g2_buf_2 _05578_ (.A(\debug_controller_inst.grid_in[43] ),
    .X(_05145_));
 sg13g2_xnor2_1 _05579_ (.Y(_05146_),
    .A(_05144_),
    .B(_05145_));
 sg13g2_nand4_1 _05580_ (.B(net356),
    .C(_05143_),
    .A(net354),
    .Y(_05147_),
    .D(_05146_));
 sg13g2_and2_1 _05581_ (.A(net355),
    .B(_05147_),
    .X(_05148_));
 sg13g2_buf_1 _05582_ (.A(\debug_controller_inst.grid_in[3] ),
    .X(_05149_));
 sg13g2_buf_2 _05583_ (.A(\debug_controller_inst.grid_in[7] ),
    .X(_05150_));
 sg13g2_xnor2_1 _05584_ (.Y(_05151_),
    .A(_05149_),
    .B(_05150_));
 sg13g2_buf_2 _05585_ (.A(\debug_controller_inst.grid_in[35] ),
    .X(_05152_));
 sg13g2_buf_2 _05586_ (.A(\debug_controller_inst.grid_in[39] ),
    .X(_05153_));
 sg13g2_xnor2_1 _05587_ (.Y(_05154_),
    .A(_05152_),
    .B(_05153_));
 sg13g2_buf_1 _05588_ (.A(net454),
    .X(_05155_));
 sg13g2_mux2_1 _05589_ (.A0(_05151_),
    .A1(_05154_),
    .S(_05155_),
    .X(_05156_));
 sg13g2_buf_2 _05590_ (.A(\debug_controller_inst.grid_in[15] ),
    .X(_05157_));
 sg13g2_buf_2 _05591_ (.A(\debug_controller_inst.grid_in[11] ),
    .X(_05158_));
 sg13g2_xnor2_1 _05592_ (.Y(_05159_),
    .A(_05157_),
    .B(_05158_));
 sg13g2_buf_2 _05593_ (.A(\debug_controller_inst.grid_in[12] ),
    .X(_05160_));
 sg13g2_buf_2 _05594_ (.A(\debug_controller_inst.grid_in[8] ),
    .X(_05161_));
 sg13g2_xor2_1 _05595_ (.B(_05161_),
    .A(_05160_),
    .X(_05162_));
 sg13g2_nor3_1 _05596_ (.A(net358),
    .B(net409),
    .C(_05162_),
    .Y(_05163_));
 sg13g2_a22oi_1 _05597_ (.Y(_05164_),
    .B1(_05159_),
    .B2(_05163_),
    .A2(_05156_),
    .A1(net409));
 sg13g2_buf_1 _05598_ (.A(\debug_controller_inst.grid_in[19] ),
    .X(_05165_));
 sg13g2_buf_2 _05599_ (.A(\debug_controller_inst.grid_in[23] ),
    .X(_05166_));
 sg13g2_xor2_1 _05600_ (.B(_05166_),
    .A(_05165_),
    .X(_05167_));
 sg13g2_buf_2 _05601_ (.A(\debug_controller_inst.grid_in[31] ),
    .X(_05168_));
 sg13g2_buf_2 _05602_ (.A(\debug_controller_inst.grid_in[27] ),
    .X(_05169_));
 sg13g2_xor2_1 _05603_ (.B(_05169_),
    .A(_05168_),
    .X(_05170_));
 sg13g2_buf_1 _05604_ (.A(\debug_controller_inst.grid_in[51] ),
    .X(_05171_));
 sg13g2_buf_2 _05605_ (.A(\debug_controller_inst.grid_in[55] ),
    .X(_05172_));
 sg13g2_xor2_1 _05606_ (.B(_05172_),
    .A(_05171_),
    .X(_05173_));
 sg13g2_buf_2 _05607_ (.A(\debug_controller_inst.grid_in[63] ),
    .X(_05174_));
 sg13g2_buf_2 _05608_ (.A(\debug_controller_inst.grid_in[59] ),
    .X(_05175_));
 sg13g2_xor2_1 _05609_ (.B(_05175_),
    .A(_05174_),
    .X(_05176_));
 sg13g2_mux4_1 _05610_ (.S0(_05135_),
    .A0(_05167_),
    .A1(_05170_),
    .A2(_05173_),
    .A3(_05176_),
    .S1(net354),
    .X(_05177_));
 sg13g2_buf_2 _05611_ (.A(\debug_controller_inst.grid_in[2] ),
    .X(_05178_));
 sg13g2_buf_2 _05612_ (.A(\debug_controller_inst.grid_in[6] ),
    .X(_05179_));
 sg13g2_xor2_1 _05613_ (.B(_05179_),
    .A(_05178_),
    .X(_05180_));
 sg13g2_buf_2 _05614_ (.A(\debug_controller_inst.grid_in[13] ),
    .X(_05181_));
 sg13g2_buf_2 _05615_ (.A(\debug_controller_inst.grid_in[9] ),
    .X(_05182_));
 sg13g2_xor2_1 _05616_ (.B(_05182_),
    .A(_05181_),
    .X(_05183_));
 sg13g2_buf_2 _05617_ (.A(\debug_controller_inst.grid_in[34] ),
    .X(_05184_));
 sg13g2_buf_2 _05618_ (.A(\debug_controller_inst.grid_in[38] ),
    .X(_05185_));
 sg13g2_xor2_1 _05619_ (.B(_05185_),
    .A(_05184_),
    .X(_05186_));
 sg13g2_buf_2 _05620_ (.A(\debug_controller_inst.grid_in[45] ),
    .X(_05187_));
 sg13g2_buf_2 _05621_ (.A(\debug_controller_inst.grid_in[41] ),
    .X(_05188_));
 sg13g2_xor2_1 _05622_ (.B(_05188_),
    .A(_05187_),
    .X(_05189_));
 sg13g2_mux4_1 _05623_ (.S0(_05135_),
    .A0(_05180_),
    .A1(_05183_),
    .A2(_05186_),
    .A3(_05189_),
    .S1(net354),
    .X(_05190_));
 sg13g2_mux2_1 _05624_ (.A0(_05177_),
    .A1(_05190_),
    .S(net355),
    .X(_05191_));
 sg13g2_a221oi_1 _05625_ (.B2(_05164_),
    .C1(_05191_),
    .B1(_05148_),
    .A1(net359),
    .Y(_05192_),
    .A2(_05137_));
 sg13g2_buf_8 _05626_ (.A(_05192_),
    .X(_05193_));
 sg13g2_buf_2 _05627_ (.A(\debug_controller_inst.grid_in[30] ),
    .X(_05194_));
 sg13g2_buf_2 _05628_ (.A(\debug_controller_inst.grid_in[26] ),
    .X(_05195_));
 sg13g2_xnor2_1 _05629_ (.Y(_05196_),
    .A(_05194_),
    .B(_05195_));
 sg13g2_buf_2 _05630_ (.A(\debug_controller_inst.grid_in[28] ),
    .X(_05197_));
 sg13g2_buf_2 _05631_ (.A(\debug_controller_inst.grid_in[24] ),
    .X(_05198_));
 sg13g2_xnor2_1 _05632_ (.Y(_05199_),
    .A(_05197_),
    .B(_05198_));
 sg13g2_nand2_1 _05633_ (.Y(_05200_),
    .A(_05196_),
    .B(_05199_));
 sg13g2_buf_2 _05634_ (.A(\debug_controller_inst.grid_in[18] ),
    .X(_05201_));
 sg13g2_buf_2 _05635_ (.A(\debug_controller_inst.grid_in[22] ),
    .X(_05202_));
 sg13g2_xor2_1 _05636_ (.B(_05202_),
    .A(_05201_),
    .X(_05203_));
 sg13g2_buf_2 _05637_ (.A(\debug_controller_inst.grid_in[62] ),
    .X(_05204_));
 sg13g2_buf_2 _05638_ (.A(\debug_controller_inst.grid_in[58] ),
    .X(_05205_));
 sg13g2_xnor2_1 _05639_ (.Y(_05206_),
    .A(_05204_),
    .B(_05205_));
 sg13g2_buf_2 _05640_ (.A(\debug_controller_inst.grid_in[60] ),
    .X(_05207_));
 sg13g2_buf_2 _05641_ (.A(\debug_controller_inst.grid_in[56] ),
    .X(_05208_));
 sg13g2_xnor2_1 _05642_ (.Y(_05209_),
    .A(_05207_),
    .B(_05208_));
 sg13g2_nand2_1 _05643_ (.Y(_05210_),
    .A(_05206_),
    .B(_05209_));
 sg13g2_buf_2 _05644_ (.A(\debug_controller_inst.grid_in[50] ),
    .X(_05211_));
 sg13g2_buf_2 _05645_ (.A(\debug_controller_inst.grid_in[54] ),
    .X(_05212_));
 sg13g2_xor2_1 _05646_ (.B(_05212_),
    .A(_05211_),
    .X(_05213_));
 sg13g2_mux4_1 _05647_ (.S0(_05117_),
    .A0(_05200_),
    .A1(_05203_),
    .A2(_05210_),
    .A3(_05213_),
    .S1(net358),
    .X(_05214_));
 sg13g2_buf_2 _05648_ (.A(\debug_controller_inst.grid_in[0] ),
    .X(_05215_));
 sg13g2_buf_2 _05649_ (.A(\debug_controller_inst.grid_in[4] ),
    .X(_05216_));
 sg13g2_xor2_1 _05650_ (.B(_05216_),
    .A(_05215_),
    .X(_05217_));
 sg13g2_buf_2 _05651_ (.A(\debug_controller_inst.grid_in[1] ),
    .X(_05218_));
 sg13g2_buf_2 _05652_ (.A(\debug_controller_inst.grid_in[5] ),
    .X(_05219_));
 sg13g2_xor2_1 _05653_ (.B(_05219_),
    .A(_05218_),
    .X(_05220_));
 sg13g2_nor3_1 _05654_ (.A(_05140_),
    .B(_05217_),
    .C(_05220_),
    .Y(_05221_));
 sg13g2_buf_2 _05655_ (.A(\debug_controller_inst.grid_in[32] ),
    .X(_05222_));
 sg13g2_buf_2 _05656_ (.A(\debug_controller_inst.grid_in[36] ),
    .X(_05223_));
 sg13g2_xnor2_1 _05657_ (.Y(_05224_),
    .A(_05222_),
    .B(_05223_));
 sg13g2_buf_2 _05658_ (.A(\debug_controller_inst.grid_in[33] ),
    .X(_05225_));
 sg13g2_buf_2 _05659_ (.A(\debug_controller_inst.grid_in[37] ),
    .X(_05226_));
 sg13g2_xnor2_1 _05660_ (.Y(_05227_),
    .A(_05225_),
    .B(_05226_));
 sg13g2_and3_1 _05661_ (.X(_05228_),
    .A(_05140_),
    .B(_05224_),
    .C(_05227_));
 sg13g2_o21ai_1 _05662_ (.B1(_05117_),
    .Y(_05229_),
    .A1(_05221_),
    .A2(_05228_));
 sg13g2_buf_2 _05663_ (.A(\debug_controller_inst.grid_in[14] ),
    .X(_00459_));
 sg13g2_buf_2 _05664_ (.A(\debug_controller_inst.grid_in[10] ),
    .X(_00460_));
 sg13g2_xnor2_1 _05665_ (.Y(_00461_),
    .A(_00459_),
    .B(_00460_));
 sg13g2_buf_2 _05666_ (.A(\debug_controller_inst.grid_in[46] ),
    .X(_00462_));
 sg13g2_buf_2 _05667_ (.A(\debug_controller_inst.grid_in[42] ),
    .X(_00463_));
 sg13g2_xnor2_1 _05668_ (.Y(_00464_),
    .A(_00462_),
    .B(_00463_));
 sg13g2_mux2_1 _05669_ (.A0(_00461_),
    .A1(_00464_),
    .S(_05155_),
    .X(_00465_));
 sg13g2_a21oi_1 _05670_ (.A1(net356),
    .A2(_00465_),
    .Y(_00466_),
    .B1(_05106_));
 sg13g2_nor2_1 _05671_ (.A(_05138_),
    .B(_05135_),
    .Y(_00467_));
 sg13g2_buf_2 _05672_ (.A(\debug_controller_inst.grid_in[16] ),
    .X(_00468_));
 sg13g2_buf_2 _05673_ (.A(\debug_controller_inst.grid_in[20] ),
    .X(_00469_));
 sg13g2_xor2_1 _05674_ (.B(_00469_),
    .A(_00468_),
    .X(_00470_));
 sg13g2_buf_2 _05675_ (.A(\debug_controller_inst.grid_in[48] ),
    .X(_00471_));
 sg13g2_buf_2 _05676_ (.A(\debug_controller_inst.grid_in[52] ),
    .X(_00472_));
 sg13g2_xor2_1 _05677_ (.B(_00472_),
    .A(_00471_),
    .X(_00473_));
 sg13g2_mux2_1 _05678_ (.A0(_00470_),
    .A1(_00473_),
    .S(net408),
    .X(_00474_));
 sg13g2_and2_1 _05679_ (.A(_00467_),
    .B(_00474_),
    .X(_00475_));
 sg13g2_a221oi_1 _05680_ (.B2(_00466_),
    .C1(_00475_),
    .B1(_05229_),
    .A1(net359),
    .Y(_00476_),
    .A2(_05214_));
 sg13g2_buf_1 _05681_ (.A(_00476_),
    .X(_00477_));
 sg13g2_mux4_1 _05682_ (.S0(net455),
    .A0(_05161_),
    .A1(_05198_),
    .A2(_05142_),
    .A3(_05208_),
    .S1(net354),
    .X(_00478_));
 sg13g2_buf_2 _05683_ (.A(_00478_),
    .X(_00479_));
 sg13g2_mux4_1 _05684_ (.S0(net411),
    .A0(_05216_),
    .A1(_00469_),
    .A2(_05223_),
    .A3(_00472_),
    .S1(net358),
    .X(_00480_));
 sg13g2_buf_2 _05685_ (.A(_00480_),
    .X(_00481_));
 sg13g2_buf_8 _05686_ (.A(net356),
    .X(_00482_));
 sg13g2_mux2_1 _05687_ (.A0(_00479_),
    .A1(_00481_),
    .S(net259),
    .X(_00483_));
 sg13g2_buf_1 _05688_ (.A(_00483_),
    .X(_00484_));
 sg13g2_nor2_1 _05689_ (.A(_00469_),
    .B(_05123_),
    .Y(_00485_));
 sg13g2_nor2_1 _05690_ (.A(_05198_),
    .B(_05126_),
    .Y(_00486_));
 sg13g2_nor2_1 _05691_ (.A(_00472_),
    .B(_05129_),
    .Y(_00487_));
 sg13g2_nor2_1 _05692_ (.A(_05208_),
    .B(_05132_),
    .Y(_00488_));
 sg13g2_mux4_1 _05693_ (.S0(net356),
    .A0(_00485_),
    .A1(_00486_),
    .A2(_00487_),
    .A3(_00488_),
    .S1(net358),
    .X(_00489_));
 sg13g2_nor2_1 _05694_ (.A(_05216_),
    .B(_05219_),
    .Y(_00490_));
 sg13g2_nor2_1 _05695_ (.A(_05161_),
    .B(_05182_),
    .Y(_00491_));
 sg13g2_nor2_1 _05696_ (.A(_05223_),
    .B(_05226_),
    .Y(_00492_));
 sg13g2_nor2_1 _05697_ (.A(_05142_),
    .B(_05188_),
    .Y(_00493_));
 sg13g2_mux4_1 _05698_ (.S0(net356),
    .A0(_00490_),
    .A1(_00491_),
    .A2(_00492_),
    .A3(_00493_),
    .S1(_05111_),
    .X(_00494_));
 sg13g2_mux2_1 _05699_ (.A0(_00489_),
    .A1(_00494_),
    .S(net355),
    .X(_00495_));
 sg13g2_mux4_1 _05700_ (.S0(_05103_),
    .A0(_05179_),
    .A1(_05202_),
    .A2(_05185_),
    .A3(_05212_),
    .S1(_05108_),
    .X(_00496_));
 sg13g2_buf_2 _05701_ (.A(_00496_),
    .X(_00497_));
 sg13g2_nor2_1 _05702_ (.A(_05135_),
    .B(_00497_),
    .Y(_00498_));
 sg13g2_mux2_1 _05703_ (.A0(_00460_),
    .A1(_00463_),
    .S(net454),
    .X(_00499_));
 sg13g2_buf_1 _05704_ (.A(_00499_),
    .X(_00500_));
 sg13g2_nor3_1 _05705_ (.A(net411),
    .B(net409),
    .C(_00500_),
    .Y(_00501_));
 sg13g2_o21ai_1 _05706_ (.B1(net455),
    .Y(_00502_),
    .A1(_05062_),
    .A2(_05083_));
 sg13g2_mux2_1 _05707_ (.A0(_05195_),
    .A1(_05205_),
    .S(net454),
    .X(_00503_));
 sg13g2_buf_1 _05708_ (.A(_00503_),
    .X(_00504_));
 sg13g2_nor2_1 _05709_ (.A(_00502_),
    .B(_00504_),
    .Y(_00505_));
 sg13g2_or3_1 _05710_ (.A(_00498_),
    .B(_00501_),
    .C(_00505_),
    .X(_00506_));
 sg13g2_buf_2 _05711_ (.A(_00506_),
    .X(_00507_));
 sg13g2_mux2_1 _05712_ (.A0(_05150_),
    .A1(_05153_),
    .S(_05108_),
    .X(_00508_));
 sg13g2_mux2_1 _05713_ (.A0(_05166_),
    .A1(_05172_),
    .S(_05109_),
    .X(_00509_));
 sg13g2_mux2_1 _05714_ (.A0(_00508_),
    .A1(_00509_),
    .S(net455),
    .X(_00510_));
 sg13g2_buf_2 _05715_ (.A(_00510_),
    .X(_00511_));
 sg13g2_mux4_1 _05716_ (.S0(net455),
    .A0(_05158_),
    .A1(_05169_),
    .A2(_05145_),
    .A3(_05175_),
    .S1(_05109_),
    .X(_00512_));
 sg13g2_or2_1 _05717_ (.X(_00513_),
    .B(_00512_),
    .A(_05116_));
 sg13g2_buf_1 _05718_ (.A(_00513_),
    .X(_00514_));
 sg13g2_o21ai_1 _05719_ (.B1(_00514_),
    .Y(_00515_),
    .A1(net356),
    .A2(_00511_));
 sg13g2_buf_2 _05720_ (.A(_00515_),
    .X(_00516_));
 sg13g2_nand3_1 _05721_ (.B(_00507_),
    .C(_00516_),
    .A(_00495_),
    .Y(_00517_));
 sg13g2_buf_1 _05722_ (.A(_00517_),
    .X(_00518_));
 sg13g2_and4_1 _05723_ (.A(net74),
    .B(net73),
    .C(net72),
    .D(_00518_),
    .X(_00519_));
 sg13g2_a21oi_1 _05724_ (.A1(net74),
    .A2(net73),
    .Y(_00520_),
    .B1(net72));
 sg13g2_mux2_1 _05725_ (.A0(_00468_),
    .A1(_05197_),
    .S(net259),
    .X(_00521_));
 sg13g2_mux2_1 _05726_ (.A0(_05215_),
    .A1(_05160_),
    .S(net259),
    .X(_00522_));
 sg13g2_mux2_1 _05727_ (.A0(_00471_),
    .A1(_05207_),
    .S(_00482_),
    .X(_00523_));
 sg13g2_mux2_1 _05728_ (.A0(_05222_),
    .A1(_05141_),
    .S(_00482_),
    .X(_00524_));
 sg13g2_mux4_1 _05729_ (.S0(net355),
    .A0(_00521_),
    .A1(_00522_),
    .A2(_00523_),
    .A3(_00524_),
    .S1(net261),
    .X(_00525_));
 sg13g2_buf_2 _05730_ (.A(_00525_),
    .X(_00526_));
 sg13g2_o21ai_1 _05731_ (.B1(_00526_),
    .Y(_00527_),
    .A1(_00519_),
    .A2(_00520_));
 sg13g2_nor2_1 _05732_ (.A(net355),
    .B(net409),
    .Y(_00528_));
 sg13g2_nor2_1 _05733_ (.A(_05207_),
    .B(_05204_),
    .Y(_00529_));
 sg13g2_nor3_1 _05734_ (.A(net410),
    .B(_05197_),
    .C(_05194_),
    .Y(_00530_));
 sg13g2_a21oi_1 _05735_ (.A1(net354),
    .A2(_00529_),
    .Y(_00531_),
    .B1(_00530_));
 sg13g2_nor2_1 _05736_ (.A(_05141_),
    .B(_00462_),
    .Y(_00532_));
 sg13g2_nor3_1 _05737_ (.A(net408),
    .B(_05160_),
    .C(_00459_),
    .Y(_00533_));
 sg13g2_a21oi_1 _05738_ (.A1(net358),
    .A2(_00532_),
    .Y(_00534_),
    .B1(_00533_));
 sg13g2_nor2_1 _05739_ (.A(net411),
    .B(net409),
    .Y(_00535_));
 sg13g2_a22oi_1 _05740_ (.Y(_00536_),
    .B1(_00534_),
    .B2(_00535_),
    .A2(_00531_),
    .A1(_00528_));
 sg13g2_buf_1 _05741_ (.A(_00536_),
    .X(_00537_));
 sg13g2_nor2_1 _05742_ (.A(_00471_),
    .B(_05211_),
    .Y(_00538_));
 sg13g2_nor3_1 _05743_ (.A(_00468_),
    .B(net410),
    .C(_05201_),
    .Y(_00539_));
 sg13g2_a21oi_1 _05744_ (.A1(net354),
    .A2(_00538_),
    .Y(_00540_),
    .B1(_00539_));
 sg13g2_nor2_1 _05745_ (.A(_05222_),
    .B(_05184_),
    .Y(_00541_));
 sg13g2_nor3_1 _05746_ (.A(_05215_),
    .B(net410),
    .C(_05178_),
    .Y(_00542_));
 sg13g2_a21oi_1 _05747_ (.A1(net358),
    .A2(_00541_),
    .Y(_00543_),
    .B1(_00542_));
 sg13g2_nor2_1 _05748_ (.A(net411),
    .B(_05136_),
    .Y(_00544_));
 sg13g2_a22oi_1 _05749_ (.Y(_00545_),
    .B1(_00543_),
    .B2(_00544_),
    .A2(_00540_),
    .A1(_00467_));
 sg13g2_buf_1 _05750_ (.A(_00545_),
    .X(_00546_));
 sg13g2_mux4_1 _05751_ (.S0(_05104_),
    .A0(_05149_),
    .A1(_05165_),
    .A2(_05152_),
    .A3(_05171_),
    .S1(net454),
    .X(_00547_));
 sg13g2_buf_2 _05752_ (.A(_00547_),
    .X(_00548_));
 sg13g2_nor2_1 _05753_ (.A(_05135_),
    .B(_00548_),
    .Y(_00549_));
 sg13g2_mux2_1 _05754_ (.A0(_05157_),
    .A1(_05144_),
    .S(net454),
    .X(_00550_));
 sg13g2_nor3_1 _05755_ (.A(net411),
    .B(_05116_),
    .C(_00550_),
    .Y(_00551_));
 sg13g2_mux2_1 _05756_ (.A0(_05168_),
    .A1(_05174_),
    .S(net454),
    .X(_00552_));
 sg13g2_nor2_1 _05757_ (.A(_00502_),
    .B(_00552_),
    .Y(_00553_));
 sg13g2_or3_1 _05758_ (.A(_00549_),
    .B(_00551_),
    .C(_00553_),
    .X(_00554_));
 sg13g2_buf_1 _05759_ (.A(_00554_),
    .X(_00555_));
 sg13g2_mux2_1 _05760_ (.A0(_05122_),
    .A1(_05128_),
    .S(net410),
    .X(_00556_));
 sg13g2_mux2_1 _05761_ (.A0(_05218_),
    .A1(_05225_),
    .S(net410),
    .X(_00557_));
 sg13g2_mux2_1 _05762_ (.A0(_05125_),
    .A1(_05131_),
    .S(net410),
    .X(_00558_));
 sg13g2_mux2_1 _05763_ (.A0(_05181_),
    .A1(_05187_),
    .S(net454),
    .X(_00559_));
 sg13g2_mux4_1 _05764_ (.S0(net355),
    .A0(_00556_),
    .A1(_00557_),
    .A2(_00558_),
    .A3(_00559_),
    .S1(_05136_),
    .X(_00560_));
 sg13g2_inv_1 _05765_ (.Y(_00561_),
    .A(_00560_));
 sg13g2_and4_1 _05766_ (.A(_00537_),
    .B(_00546_),
    .C(_00555_),
    .D(_00561_),
    .X(_00562_));
 sg13g2_buf_8 _05767_ (.A(_00562_),
    .X(_00563_));
 sg13g2_and2_1 _05768_ (.A(_00495_),
    .B(_00516_),
    .X(_00564_));
 sg13g2_mux2_1 _05769_ (.A0(_05179_),
    .A1(_05185_),
    .S(_05110_),
    .X(_00565_));
 sg13g2_mux2_1 _05770_ (.A0(_05202_),
    .A1(_05212_),
    .S(_05110_),
    .X(_00566_));
 sg13g2_mux4_1 _05771_ (.S0(net411),
    .A0(_00565_),
    .A1(_00566_),
    .A2(_00500_),
    .A3(_00504_),
    .S1(net409),
    .X(_00567_));
 sg13g2_buf_1 _05772_ (.A(_00567_),
    .X(_00568_));
 sg13g2_nand2_1 _05773_ (.Y(_00569_),
    .A(_00507_),
    .B(net159));
 sg13g2_nand2b_1 _05774_ (.Y(_00570_),
    .B(_00479_),
    .A_N(_00481_));
 sg13g2_nand2b_1 _05775_ (.Y(_00571_),
    .B(_00481_),
    .A_N(_00479_));
 sg13g2_nand2b_1 _05776_ (.Y(_00572_),
    .B(_00565_),
    .A_N(_00500_));
 sg13g2_nand2b_1 _05777_ (.Y(_00573_),
    .B(_00500_),
    .A_N(_00565_));
 sg13g2_nand2b_1 _05778_ (.Y(_00574_),
    .B(_00566_),
    .A_N(_00504_));
 sg13g2_nand2b_1 _05779_ (.Y(_00575_),
    .B(_00504_),
    .A_N(_00566_));
 sg13g2_mux4_1 _05780_ (.S0(net259),
    .A0(_00572_),
    .A1(_00573_),
    .A2(_00574_),
    .A3(_00575_),
    .S1(net359),
    .X(_00576_));
 sg13g2_and3_1 _05781_ (.X(_00577_),
    .A(_00570_),
    .B(_00571_),
    .C(_00576_));
 sg13g2_o21ai_1 _05782_ (.B1(_00577_),
    .Y(_00578_),
    .A1(_00564_),
    .A2(_00569_));
 sg13g2_and2_1 _05783_ (.A(net357),
    .B(_00479_),
    .X(_00579_));
 sg13g2_a21oi_1 _05784_ (.A1(net259),
    .A2(_00481_),
    .Y(_00580_),
    .B1(_00579_));
 sg13g2_buf_2 _05785_ (.A(_00580_),
    .X(_00581_));
 sg13g2_mux2_1 _05786_ (.A0(_05178_),
    .A1(_05184_),
    .S(net408),
    .X(_00582_));
 sg13g2_mux2_1 _05787_ (.A0(_00459_),
    .A1(_00462_),
    .S(net354),
    .X(_00583_));
 sg13g2_mux2_1 _05788_ (.A0(_05201_),
    .A1(_05211_),
    .S(net408),
    .X(_00584_));
 sg13g2_mux2_1 _05789_ (.A0(_05194_),
    .A1(_05204_),
    .S(net408),
    .X(_00585_));
 sg13g2_mux4_1 _05790_ (.S0(net356),
    .A0(_00582_),
    .A1(_00583_),
    .A2(_00584_),
    .A3(_00585_),
    .S1(_05106_),
    .X(_00586_));
 sg13g2_xor2_1 _05791_ (.B(_00586_),
    .A(_00568_),
    .X(_00587_));
 sg13g2_a21oi_1 _05792_ (.A1(_00526_),
    .A2(_00581_),
    .Y(_00588_),
    .B1(_00587_));
 sg13g2_nor2_1 _05793_ (.A(_00518_),
    .B(_00588_),
    .Y(_00589_));
 sg13g2_a21oi_1 _05794_ (.A1(net57),
    .A2(_00578_),
    .Y(_00590_),
    .B1(_00589_));
 sg13g2_nand2_1 _05795_ (.Y(_00591_),
    .A(net74),
    .B(net73));
 sg13g2_nor2_1 _05796_ (.A(_00526_),
    .B(net57),
    .Y(_00592_));
 sg13g2_nand3_1 _05797_ (.B(_00484_),
    .C(_00592_),
    .A(_00591_),
    .Y(_00593_));
 sg13g2_and2_1 _05798_ (.A(net74),
    .B(net73),
    .X(_00594_));
 sg13g2_buf_2 _05799_ (.A(_00594_),
    .X(_00595_));
 sg13g2_nand3_1 _05800_ (.B(_00581_),
    .C(_00592_),
    .A(_00595_),
    .Y(_00596_));
 sg13g2_nand4_1 _05801_ (.B(_00590_),
    .C(_00593_),
    .A(_00527_),
    .Y(_00597_),
    .D(_00596_));
 sg13g2_buf_1 _05802_ (.A(_00597_),
    .X(_00598_));
 sg13g2_mux2_1 _05803_ (.A0(_05158_),
    .A1(_05145_),
    .S(net261),
    .X(_00599_));
 sg13g2_mux2_1 _05804_ (.A0(_05169_),
    .A1(_05175_),
    .S(net261),
    .X(_00600_));
 sg13g2_mux4_1 _05805_ (.S0(net359),
    .A0(_00508_),
    .A1(_00509_),
    .A2(_00599_),
    .A3(_00600_),
    .S1(_05118_),
    .X(_00601_));
 sg13g2_buf_1 _05806_ (.A(_00601_),
    .X(_00602_));
 sg13g2_inv_1 _05807_ (.Y(_00603_),
    .A(_00555_));
 sg13g2_and2_1 _05808_ (.A(_00546_),
    .B(_00561_),
    .X(_00604_));
 sg13g2_nor2b_1 _05809_ (.A(_00516_),
    .B_N(_00537_),
    .Y(_00605_));
 sg13g2_a21oi_1 _05810_ (.A1(_00604_),
    .A2(_00605_),
    .Y(_00606_),
    .B1(_00603_));
 sg13g2_mux4_1 _05811_ (.S0(_05105_),
    .A0(_05215_),
    .A1(_00468_),
    .A2(_05222_),
    .A3(_00471_),
    .S1(net354),
    .X(_00607_));
 sg13g2_mux4_1 _05812_ (.S0(net455),
    .A0(_05218_),
    .A1(_05122_),
    .A2(_05225_),
    .A3(_05128_),
    .S1(net408),
    .X(_00608_));
 sg13g2_nand3_1 _05813_ (.B(_00607_),
    .C(_00608_),
    .A(net409),
    .Y(_00609_));
 sg13g2_mux4_1 _05814_ (.S0(_05104_),
    .A0(_05160_),
    .A1(_05197_),
    .A2(_05141_),
    .A3(_05207_),
    .S1(net408),
    .X(_00610_));
 sg13g2_mux4_1 _05815_ (.S0(net455),
    .A0(_05181_),
    .A1(_05125_),
    .A2(_05187_),
    .A3(_05131_),
    .S1(net408),
    .X(_00611_));
 sg13g2_nand3_1 _05816_ (.B(_00610_),
    .C(_00611_),
    .A(net259),
    .Y(_00612_));
 sg13g2_nand2_1 _05817_ (.Y(_00613_),
    .A(_00609_),
    .B(_00612_));
 sg13g2_and2_1 _05818_ (.A(_00586_),
    .B(_00613_),
    .X(_00614_));
 sg13g2_nand3_1 _05819_ (.B(_00477_),
    .C(_00614_),
    .A(net74),
    .Y(_00615_));
 sg13g2_mux2_1 _05820_ (.A0(_00603_),
    .A1(_00606_),
    .S(_00615_),
    .X(_00616_));
 sg13g2_buf_2 _05821_ (.A(_00616_),
    .X(_00617_));
 sg13g2_xnor2_1 _05822_ (.Y(_00618_),
    .A(net71),
    .B(_00617_));
 sg13g2_nand2b_1 _05823_ (.Y(_00619_),
    .B(_00518_),
    .A_N(_00587_));
 sg13g2_nand4_1 _05824_ (.B(_00546_),
    .C(_00555_),
    .A(_00537_),
    .Y(_00620_),
    .D(_00561_));
 sg13g2_buf_1 _05825_ (.A(_00620_),
    .X(_00621_));
 sg13g2_nand2_1 _05826_ (.Y(_00622_),
    .A(net56),
    .B(_00587_));
 sg13g2_nand3_1 _05827_ (.B(net73),
    .C(_00613_),
    .A(_05193_),
    .Y(_00623_));
 sg13g2_mux2_1 _05828_ (.A0(_00619_),
    .A1(_00622_),
    .S(_00623_),
    .X(_00624_));
 sg13g2_buf_1 _05829_ (.A(_00624_),
    .X(_00625_));
 sg13g2_nand3_1 _05830_ (.B(net74),
    .C(net73),
    .A(_00526_),
    .Y(_00626_));
 sg13g2_mux4_1 _05831_ (.S0(net411),
    .A0(_05219_),
    .A1(_05123_),
    .A2(_05226_),
    .A3(_05129_),
    .S1(net261),
    .X(_00627_));
 sg13g2_buf_2 _05832_ (.A(_00627_),
    .X(_00628_));
 sg13g2_mux4_1 _05833_ (.S0(_05105_),
    .A0(_05182_),
    .A1(_05126_),
    .A2(_05188_),
    .A3(_05132_),
    .S1(_05111_),
    .X(_00629_));
 sg13g2_buf_2 _05834_ (.A(_00629_),
    .X(_00630_));
 sg13g2_and2_1 _05835_ (.A(net259),
    .B(_00630_),
    .X(_00631_));
 sg13g2_a21o_1 _05836_ (.A2(_00628_),
    .A1(net357),
    .B1(_00631_),
    .X(_00632_));
 sg13g2_nand4_1 _05837_ (.B(_00546_),
    .C(_00555_),
    .A(_00537_),
    .Y(_00633_),
    .D(_00632_));
 sg13g2_and2_1 _05838_ (.A(_00561_),
    .B(_00633_),
    .X(_00634_));
 sg13g2_nand2b_1 _05839_ (.Y(_00635_),
    .B(net357),
    .A_N(_00630_));
 sg13g2_or2_1 _05840_ (.X(_00636_),
    .B(_00628_),
    .A(net357));
 sg13g2_nand2_2 _05841_ (.Y(_00637_),
    .A(_00635_),
    .B(_00636_));
 sg13g2_a221oi_1 _05842_ (.B2(_00634_),
    .C1(_00637_),
    .B1(_00626_),
    .A1(_00595_),
    .Y(_00638_),
    .A2(_00613_));
 sg13g2_inv_1 _05843_ (.Y(_00639_),
    .A(_00526_));
 sg13g2_a21oi_1 _05844_ (.A1(net74),
    .A2(net73),
    .Y(_00640_),
    .B1(_00639_));
 sg13g2_mux2_1 _05845_ (.A0(_00479_),
    .A1(_00481_),
    .S(net357),
    .X(_00641_));
 sg13g2_buf_1 _05846_ (.A(_00641_),
    .X(_00642_));
 sg13g2_nand2_1 _05847_ (.Y(_00643_),
    .A(net57),
    .B(_00642_));
 sg13g2_nand2b_1 _05848_ (.Y(_00644_),
    .B(_00643_),
    .A_N(_00640_));
 sg13g2_nand3_1 _05849_ (.B(_00638_),
    .C(_00644_),
    .A(_00625_),
    .Y(_00645_));
 sg13g2_buf_1 _05850_ (.A(_00645_),
    .X(_00646_));
 sg13g2_or3_1 _05851_ (.A(_00598_),
    .B(_00618_),
    .C(_00646_),
    .X(_00647_));
 sg13g2_buf_1 _05852_ (.A(_00647_),
    .X(_00648_));
 sg13g2_buf_1 _05853_ (.A(_00518_),
    .X(_00649_));
 sg13g2_and2_1 _05854_ (.A(_00649_),
    .B(net57),
    .X(_00650_));
 sg13g2_a21oi_1 _05855_ (.A1(net52),
    .A2(_00563_),
    .Y(_00651_),
    .B1(_00586_));
 sg13g2_and3_1 _05856_ (.X(_00652_),
    .A(_05193_),
    .B(_00477_),
    .C(_00614_));
 sg13g2_a221oi_1 _05857_ (.B2(_00623_),
    .C1(_00652_),
    .B1(_00651_),
    .A1(_00507_),
    .Y(_00653_),
    .A2(_00650_));
 sg13g2_buf_1 _05858_ (.A(_00653_),
    .X(_00654_));
 sg13g2_nor2_1 _05859_ (.A(_00518_),
    .B(net56),
    .Y(_00655_));
 sg13g2_buf_2 _05860_ (.A(_00655_),
    .X(_00656_));
 sg13g2_a221oi_1 _05861_ (.B2(_00564_),
    .C1(_00563_),
    .B1(_00507_),
    .A1(net74),
    .Y(_00657_),
    .A2(net73));
 sg13g2_buf_1 _05862_ (.A(_00657_),
    .X(_00658_));
 sg13g2_or2_1 _05863_ (.X(_00659_),
    .B(_00658_),
    .A(_00656_));
 sg13g2_buf_1 _05864_ (.A(_00659_),
    .X(_00660_));
 sg13g2_buf_1 _05865_ (.A(_00660_),
    .X(_00661_));
 sg13g2_buf_1 _05866_ (.A(net259),
    .X(_00662_));
 sg13g2_mux2_1 _05867_ (.A0(_00582_),
    .A1(_00584_),
    .S(net262),
    .X(_00663_));
 sg13g2_mux4_1 _05868_ (.S0(net359),
    .A0(_00459_),
    .A1(_05194_),
    .A2(_00462_),
    .A3(_05204_),
    .S1(net261),
    .X(_00664_));
 sg13g2_and2_1 _05869_ (.A(_05119_),
    .B(_00664_),
    .X(_00665_));
 sg13g2_a21o_1 _05870_ (.A2(_00663_),
    .A1(_00662_),
    .B1(_00665_),
    .X(_00666_));
 sg13g2_buf_1 _05871_ (.A(_00666_),
    .X(_00667_));
 sg13g2_nor3_1 _05872_ (.A(net37),
    .B(net35),
    .C(net55),
    .Y(_00668_));
 sg13g2_a21oi_1 _05873_ (.A1(_00662_),
    .A2(_00663_),
    .Y(_00669_),
    .B1(_00665_));
 sg13g2_buf_2 _05874_ (.A(_00669_),
    .X(_00670_));
 sg13g2_buf_8 _05875_ (.A(_00658_),
    .X(_00671_));
 sg13g2_or2_1 _05876_ (.X(_00672_),
    .B(net159),
    .A(net72));
 sg13g2_buf_1 _05877_ (.A(_00672_),
    .X(_00673_));
 sg13g2_mux2_1 _05878_ (.A0(_00628_),
    .A1(_00630_),
    .S(net357),
    .X(_00674_));
 sg13g2_buf_1 _05879_ (.A(_00674_),
    .X(_00675_));
 sg13g2_nor2_1 _05880_ (.A(net71),
    .B(net54),
    .Y(_00676_));
 sg13g2_nor2b_1 _05881_ (.A(_00673_),
    .B_N(_00676_),
    .Y(_00677_));
 sg13g2_nor3_2 _05882_ (.A(_00656_),
    .B(net44),
    .C(_00677_),
    .Y(_00678_));
 sg13g2_nand3_1 _05883_ (.B(_00670_),
    .C(_00678_),
    .A(net37),
    .Y(_00679_));
 sg13g2_nor2_1 _05884_ (.A(_00646_),
    .B(_00679_),
    .Y(_00680_));
 sg13g2_nor2_1 _05885_ (.A(_00598_),
    .B(_00618_),
    .Y(_00681_));
 sg13g2_buf_1 _05886_ (.A(_00677_),
    .X(_00682_));
 sg13g2_inv_1 _05887_ (.Y(_00683_),
    .A(_00586_));
 sg13g2_nand2b_1 _05888_ (.Y(_00684_),
    .B(_00676_),
    .A_N(_00673_));
 sg13g2_buf_1 _05889_ (.A(_00684_),
    .X(_00685_));
 sg13g2_o21ai_1 _05890_ (.B1(_00685_),
    .Y(_00686_),
    .A1(net52),
    .A2(net56));
 sg13g2_inv_1 _05891_ (.Y(_00687_),
    .A(net159));
 sg13g2_a22oi_1 _05892_ (.Y(_00688_),
    .B1(_00686_),
    .B2(_00687_),
    .A2(net44),
    .A1(_00683_));
 sg13g2_buf_1 _05893_ (.A(_00688_),
    .X(_00689_));
 sg13g2_a22oi_1 _05894_ (.Y(_00690_),
    .B1(_00689_),
    .B2(net35),
    .A2(net43),
    .A1(net37));
 sg13g2_or3_1 _05895_ (.A(net37),
    .B(net55),
    .C(_00689_),
    .X(_00691_));
 sg13g2_o21ai_1 _05896_ (.B1(_00691_),
    .Y(_00692_),
    .A1(_00670_),
    .A2(_00690_));
 sg13g2_a221oi_1 _05897_ (.B2(_00681_),
    .C1(_00692_),
    .B1(_00680_),
    .A1(_00648_),
    .Y(_00693_),
    .A2(_00668_));
 sg13g2_nand3b_1 _05898_ (.B(net55),
    .C(_00689_),
    .Y(_00694_),
    .A_N(net37));
 sg13g2_nand3_1 _05899_ (.B(net55),
    .C(_00689_),
    .A(net37),
    .Y(_00695_));
 sg13g2_mux2_1 _05900_ (.A0(_00694_),
    .A1(_00695_),
    .S(_00648_),
    .X(_00696_));
 sg13g2_nand2_1 _05901_ (.Y(_00697_),
    .A(net35),
    .B(net42));
 sg13g2_and4_1 _05902_ (.A(_00527_),
    .B(_00590_),
    .C(_00593_),
    .D(_00596_),
    .X(_00698_));
 sg13g2_buf_1 _05903_ (.A(_00698_),
    .X(_00699_));
 sg13g2_inv_1 _05904_ (.Y(_00700_),
    .A(net71));
 sg13g2_xnor2_1 _05905_ (.Y(_00701_),
    .A(_00700_),
    .B(_00617_));
 sg13g2_a22oi_1 _05906_ (.Y(_00702_),
    .B1(_00626_),
    .B2(_00634_),
    .A2(_00613_),
    .A1(_00595_));
 sg13g2_xnor2_1 _05907_ (.Y(_00703_),
    .A(net54),
    .B(_00702_));
 sg13g2_nand4_1 _05908_ (.B(_00701_),
    .C(_00625_),
    .A(_00699_),
    .Y(_00704_),
    .D(_00703_));
 sg13g2_buf_2 _05909_ (.A(_00704_),
    .X(_00705_));
 sg13g2_nand2_1 _05910_ (.Y(_00706_),
    .A(_00595_),
    .B(_00621_));
 sg13g2_o21ai_1 _05911_ (.B1(_00706_),
    .Y(_00707_),
    .A1(net43),
    .A2(_00705_));
 sg13g2_and2_1 _05912_ (.A(net357),
    .B(_00610_),
    .X(_00708_));
 sg13g2_buf_1 _05913_ (.A(_00708_),
    .X(_00709_));
 sg13g2_and2_1 _05914_ (.A(net158),
    .B(_00607_),
    .X(_00710_));
 sg13g2_buf_1 _05915_ (.A(_00710_),
    .X(_00711_));
 sg13g2_or2_1 _05916_ (.X(_00712_),
    .B(_00711_),
    .A(_00709_));
 sg13g2_buf_2 _05917_ (.A(_00712_),
    .X(_00713_));
 sg13g2_a221oi_1 _05918_ (.B2(net57),
    .C1(_00640_),
    .B1(_00642_),
    .A1(_00595_),
    .Y(_00714_),
    .A2(_00592_));
 sg13g2_buf_1 _05919_ (.A(_00714_),
    .X(_00715_));
 sg13g2_nand2_1 _05920_ (.Y(_00716_),
    .A(_00656_),
    .B(net42));
 sg13g2_buf_1 _05921_ (.A(_00716_),
    .X(_00717_));
 sg13g2_mux2_1 _05922_ (.A0(_00581_),
    .A1(_00715_),
    .S(_00717_),
    .X(_00718_));
 sg13g2_xnor2_1 _05923_ (.Y(_00719_),
    .A(_00713_),
    .B(_00718_));
 sg13g2_nor2_1 _05924_ (.A(_00709_),
    .B(_00711_),
    .Y(_00720_));
 sg13g2_buf_2 _05925_ (.A(_00720_),
    .X(_00721_));
 sg13g2_nand2b_1 _05926_ (.Y(_00722_),
    .B(net42),
    .A_N(net44));
 sg13g2_nor3_1 _05927_ (.A(net72),
    .B(net52),
    .C(net56),
    .Y(_00723_));
 sg13g2_nor3_1 _05928_ (.A(net44),
    .B(net43),
    .C(_00723_),
    .Y(_00724_));
 sg13g2_mux2_1 _05929_ (.A0(_00722_),
    .A1(_00724_),
    .S(_00715_),
    .X(_00725_));
 sg13g2_xnor2_1 _05930_ (.Y(_00726_),
    .A(_00721_),
    .B(_00725_));
 sg13g2_and2_1 _05931_ (.A(_00625_),
    .B(_00706_),
    .X(_00727_));
 sg13g2_and4_1 _05932_ (.A(_00699_),
    .B(_00701_),
    .C(_00703_),
    .D(_00727_),
    .X(_00728_));
 sg13g2_buf_1 _05933_ (.A(_00728_),
    .X(_00729_));
 sg13g2_mux2_1 _05934_ (.A0(_00719_),
    .A1(_00726_),
    .S(_00729_),
    .X(_00730_));
 sg13g2_a221oi_1 _05935_ (.B2(_00707_),
    .C1(_00730_),
    .B1(_00697_),
    .A1(_00693_),
    .Y(_00731_),
    .A2(_00696_));
 sg13g2_buf_2 _05936_ (.A(_00731_),
    .X(_00732_));
 sg13g2_mux4_1 _05937_ (.S0(net359),
    .A0(_05157_),
    .A1(_05168_),
    .A2(_05144_),
    .A3(_05174_),
    .S1(net261),
    .X(_00733_));
 sg13g2_and2_1 _05938_ (.A(net357),
    .B(_00733_),
    .X(_00734_));
 sg13g2_buf_1 _05939_ (.A(_00734_),
    .X(_00735_));
 sg13g2_a21oi_2 _05940_ (.B1(_00735_),
    .Y(_00736_),
    .A2(_00548_),
    .A1(net158));
 sg13g2_nand2_1 _05941_ (.Y(_00737_),
    .A(_00615_),
    .B(_00606_));
 sg13g2_nor3_1 _05942_ (.A(net52),
    .B(net56),
    .C(_00700_),
    .Y(_00738_));
 sg13g2_nand2_1 _05943_ (.Y(_00739_),
    .A(_00603_),
    .B(_00652_));
 sg13g2_o21ai_1 _05944_ (.B1(_00739_),
    .Y(_00740_),
    .A1(_00737_),
    .A2(_00738_));
 sg13g2_nor2_1 _05945_ (.A(net71),
    .B(_00717_),
    .Y(_00741_));
 sg13g2_mux2_1 _05946_ (.A0(_00678_),
    .A1(_00722_),
    .S(_00617_),
    .X(_00742_));
 sg13g2_or2_1 _05947_ (.X(_00743_),
    .B(_00742_),
    .A(_00741_));
 sg13g2_nand4_1 _05948_ (.B(_00638_),
    .C(_00644_),
    .A(_00625_),
    .Y(_00744_),
    .D(_00654_));
 sg13g2_nor3_1 _05949_ (.A(_00598_),
    .B(_00618_),
    .C(_00744_),
    .Y(_00745_));
 sg13g2_mux2_1 _05950_ (.A0(_00740_),
    .A1(_00743_),
    .S(_00745_),
    .X(_00746_));
 sg13g2_buf_1 _05951_ (.A(_00746_),
    .X(_00747_));
 sg13g2_xnor2_1 _05952_ (.Y(_00748_),
    .A(_00736_),
    .B(net33));
 sg13g2_buf_2 _05953_ (.A(_00748_),
    .X(_00749_));
 sg13g2_and2_1 _05954_ (.A(net158),
    .B(_00608_),
    .X(_00750_));
 sg13g2_buf_1 _05955_ (.A(_00750_),
    .X(_00751_));
 sg13g2_a21o_1 _05956_ (.A2(_00611_),
    .A1(net260),
    .B1(_00751_),
    .X(_00752_));
 sg13g2_buf_2 _05957_ (.A(_00752_),
    .X(_00753_));
 sg13g2_nor3_1 _05958_ (.A(_00598_),
    .B(_00618_),
    .C(_00646_),
    .Y(_00754_));
 sg13g2_nor2b_1 _05959_ (.A(_00702_),
    .B_N(_00717_),
    .Y(_00755_));
 sg13g2_or2_1 _05960_ (.X(_00756_),
    .B(_00640_),
    .A(net57));
 sg13g2_a21oi_1 _05961_ (.A1(_00649_),
    .A2(_00643_),
    .Y(_00757_),
    .B1(net43));
 sg13g2_a21o_1 _05962_ (.A2(_00757_),
    .A1(_00756_),
    .B1(_00702_),
    .X(_00758_));
 sg13g2_o21ai_1 _05963_ (.B1(_00758_),
    .Y(_00759_),
    .A1(_00675_),
    .A2(_00717_));
 sg13g2_a221oi_1 _05964_ (.B2(_00755_),
    .C1(_00759_),
    .B1(_00705_),
    .A1(_00754_),
    .Y(_00760_),
    .A2(_00678_));
 sg13g2_buf_2 _05965_ (.A(_00760_),
    .X(_00761_));
 sg13g2_xnor2_1 _05966_ (.Y(_00762_),
    .A(_00753_),
    .B(_00761_));
 sg13g2_nand2_1 _05967_ (.Y(_00763_),
    .A(_00670_),
    .B(_00721_));
 sg13g2_a21oi_1 _05968_ (.A1(net260),
    .A2(_00611_),
    .Y(_00764_),
    .B1(_00751_));
 sg13g2_buf_1 _05969_ (.A(_00764_),
    .X(_00765_));
 sg13g2_nand2_1 _05970_ (.Y(_00766_),
    .A(_00736_),
    .B(net51));
 sg13g2_nor2_1 _05971_ (.A(_00763_),
    .B(_00766_),
    .Y(_00767_));
 sg13g2_buf_2 _05972_ (.A(_00767_),
    .X(_00768_));
 sg13g2_nor4_2 _05973_ (.A(net52),
    .B(net56),
    .C(net42),
    .Y(_00769_),
    .D(_00768_));
 sg13g2_nand4_1 _05974_ (.B(_00701_),
    .C(_00703_),
    .A(_00699_),
    .Y(_00770_),
    .D(_00727_));
 sg13g2_buf_1 _05975_ (.A(_00770_),
    .X(_00771_));
 sg13g2_nand3_1 _05976_ (.B(net52),
    .C(net56),
    .A(_00591_),
    .Y(_00772_));
 sg13g2_buf_1 _05977_ (.A(_00772_),
    .X(_00773_));
 sg13g2_or2_1 _05978_ (.X(_00774_),
    .B(_00766_),
    .A(_00763_));
 sg13g2_buf_1 _05979_ (.A(_00774_),
    .X(_00775_));
 sg13g2_nand2_1 _05980_ (.Y(_00776_),
    .A(_00773_),
    .B(_00775_));
 sg13g2_a21o_1 _05981_ (.A2(net34),
    .A1(_00678_),
    .B1(_00776_),
    .X(_00777_));
 sg13g2_a21oi_1 _05982_ (.A1(_00721_),
    .A2(_00769_),
    .Y(_00778_),
    .B1(_00777_));
 sg13g2_nand4_1 _05983_ (.B(_00749_),
    .C(_00762_),
    .A(_00732_),
    .Y(_00779_),
    .D(_00778_));
 sg13g2_and2_1 _05984_ (.A(_00591_),
    .B(_00625_),
    .X(_00780_));
 sg13g2_nand4_1 _05985_ (.B(_00701_),
    .C(_00703_),
    .A(_00699_),
    .Y(_00781_),
    .D(_00780_));
 sg13g2_nor2_1 _05986_ (.A(net57),
    .B(net43),
    .Y(_00782_));
 sg13g2_and2_1 _05987_ (.A(net52),
    .B(net42),
    .X(_00783_));
 sg13g2_buf_1 _05988_ (.A(_00783_),
    .X(_00784_));
 sg13g2_buf_8 _05989_ (.A(net44),
    .X(_00785_));
 sg13g2_a21o_1 _05990_ (.A2(net43),
    .A1(_00656_),
    .B1(_00785_),
    .X(_00786_));
 sg13g2_a221oi_1 _05991_ (.B2(_00705_),
    .C1(_00786_),
    .B1(_00784_),
    .A1(_00781_),
    .Y(_00787_),
    .A2(_00782_));
 sg13g2_buf_1 _05992_ (.A(_00787_),
    .X(_00788_));
 sg13g2_nand2_2 _05993_ (.Y(_00789_),
    .A(_00775_),
    .B(_00788_));
 sg13g2_nor2_1 _05994_ (.A(net72),
    .B(_00717_),
    .Y(_00790_));
 sg13g2_a21oi_1 _05995_ (.A1(_00717_),
    .A2(_00715_),
    .Y(_00791_),
    .B1(_00790_));
 sg13g2_mux2_1 _05996_ (.A0(_00791_),
    .A1(_00725_),
    .S(_00729_),
    .X(_00792_));
 sg13g2_buf_2 _05997_ (.A(_00792_),
    .X(_00793_));
 sg13g2_a21oi_1 _05998_ (.A1(_00789_),
    .A2(_00778_),
    .Y(_00794_),
    .B1(_00793_));
 sg13g2_and4_1 _05999_ (.A(_00732_),
    .B(_00749_),
    .C(_00762_),
    .D(_00793_),
    .X(_00795_));
 sg13g2_a21oi_1 _06000_ (.A1(_00656_),
    .A2(net43),
    .Y(_00796_),
    .B1(_00768_));
 sg13g2_nand2_1 _06001_ (.Y(_00797_),
    .A(_00773_),
    .B(_00796_));
 sg13g2_a221oi_1 _06002_ (.B2(_00705_),
    .C1(_00797_),
    .B1(_00784_),
    .A1(_00781_),
    .Y(_00798_),
    .A2(_00782_));
 sg13g2_buf_2 _06003_ (.A(_00798_),
    .X(_00799_));
 sg13g2_a22oi_1 _06004_ (.Y(_00800_),
    .B1(_00795_),
    .B2(_00799_),
    .A2(_00794_),
    .A1(_00779_));
 sg13g2_xnor2_1 _06005_ (.Y(_00801_),
    .A(_05166_),
    .B(_05169_));
 sg13g2_xnor2_1 _06006_ (.Y(_00802_),
    .A(_05172_),
    .B(_05175_));
 sg13g2_mux2_1 _06007_ (.A0(_00801_),
    .A1(_00802_),
    .S(net261),
    .X(_00803_));
 sg13g2_xnor2_1 _06008_ (.Y(_00804_),
    .A(_00508_),
    .B(_00599_));
 sg13g2_mux2_1 _06009_ (.A0(_00803_),
    .A1(_00804_),
    .S(net355),
    .X(_00805_));
 sg13g2_mux4_1 _06010_ (.S0(net359),
    .A0(_00460_),
    .A1(_05195_),
    .A2(_00463_),
    .A3(_05205_),
    .S1(net261),
    .X(_00806_));
 sg13g2_buf_1 _06011_ (.A(_00806_),
    .X(_00807_));
 sg13g2_xor2_1 _06012_ (.B(_00807_),
    .A(_00497_),
    .X(_00808_));
 sg13g2_xor2_1 _06013_ (.B(_00630_),
    .A(_00628_),
    .X(_00809_));
 sg13g2_nor2_1 _06014_ (.A(_00808_),
    .B(_00809_),
    .Y(_00810_));
 sg13g2_nand4_1 _06015_ (.B(_00571_),
    .C(_00805_),
    .A(_00570_),
    .Y(_00811_),
    .D(_00810_));
 sg13g2_buf_2 _06016_ (.A(_00811_),
    .X(_00812_));
 sg13g2_buf_1 _06017_ (.A(_00812_),
    .X(_00813_));
 sg13g2_a21o_1 _06018_ (.A2(_00548_),
    .A1(net158),
    .B1(_00735_),
    .X(_00814_));
 sg13g2_buf_2 _06019_ (.A(_00814_),
    .X(_00815_));
 sg13g2_nor4_1 _06020_ (.A(net71),
    .B(_00637_),
    .C(_00815_),
    .D(net51),
    .Y(_00816_));
 sg13g2_nand3_1 _06021_ (.B(net41),
    .C(_00816_),
    .A(net36),
    .Y(_00817_));
 sg13g2_nand3_1 _06022_ (.B(_00736_),
    .C(net51),
    .A(_00676_),
    .Y(_00818_));
 sg13g2_xnor2_1 _06023_ (.Y(_00819_),
    .A(net54),
    .B(net51));
 sg13g2_nand2_1 _06024_ (.Y(_00820_),
    .A(net71),
    .B(_00815_));
 sg13g2_nor2_1 _06025_ (.A(_00819_),
    .B(_00820_),
    .Y(_00821_));
 sg13g2_nand3_1 _06026_ (.B(net41),
    .C(_00821_),
    .A(net44),
    .Y(_00822_));
 sg13g2_a21o_1 _06027_ (.A2(net41),
    .A1(net44),
    .B1(_00766_),
    .X(_00823_));
 sg13g2_nand4_1 _06028_ (.B(_00818_),
    .C(_00822_),
    .A(_00817_),
    .Y(_00824_),
    .D(_00823_));
 sg13g2_inv_1 _06029_ (.Y(_00825_),
    .A(_00763_));
 sg13g2_nand3_1 _06030_ (.B(_00673_),
    .C(net41),
    .A(net36),
    .Y(_00826_));
 sg13g2_xnor2_1 _06031_ (.Y(_00827_),
    .A(net159),
    .B(_00670_));
 sg13g2_nand2_1 _06032_ (.Y(_00828_),
    .A(net72),
    .B(_00713_));
 sg13g2_nand4_1 _06033_ (.B(net159),
    .C(net55),
    .A(_00581_),
    .Y(_00829_),
    .D(_00721_));
 sg13g2_o21ai_1 _06034_ (.B1(_00829_),
    .Y(_00830_),
    .A1(_00827_),
    .A2(_00828_));
 sg13g2_and3_1 _06035_ (.X(_00831_),
    .A(net36),
    .B(net41),
    .C(_00830_));
 sg13g2_a21o_1 _06036_ (.A2(_00826_),
    .A1(_00825_),
    .B1(_00831_),
    .X(_00832_));
 sg13g2_and2_1 _06037_ (.A(net36),
    .B(net41),
    .X(_00833_));
 sg13g2_buf_1 _06038_ (.A(_00833_),
    .X(_00834_));
 sg13g2_nand2_1 _06039_ (.Y(_00835_),
    .A(net42),
    .B(_00834_));
 sg13g2_a21oi_1 _06040_ (.A1(_00824_),
    .A2(_00832_),
    .Y(_00836_),
    .B1(_00835_));
 sg13g2_buf_1 _06041_ (.A(_00836_),
    .X(_00837_));
 sg13g2_and2_1 _06042_ (.A(_00711_),
    .B(net32),
    .X(_00838_));
 sg13g2_a21o_1 _06043_ (.A2(_00800_),
    .A1(net94),
    .B1(_00838_),
    .X(_00839_));
 sg13g2_buf_1 _06044_ (.A(_00839_),
    .X(_00840_));
 sg13g2_nand2_1 _06045_ (.Y(_00841_),
    .A(_00098_),
    .B(net75));
 sg13g2_o21ai_1 _06046_ (.B1(_00841_),
    .Y(_00842_),
    .A1(net75),
    .A2(_00840_));
 sg13g2_buf_2 _06047_ (.A(\game_logic_inst.should_transpose ),
    .X(_00843_));
 sg13g2_inv_1 _06048_ (.Y(_00844_),
    .A(_05078_));
 sg13g2_nand2_1 _06049_ (.Y(_00845_),
    .A(net480),
    .B(_00844_));
 sg13g2_buf_1 _06050_ (.A(_00845_),
    .X(_00846_));
 sg13g2_nor2_1 _06051_ (.A(_00843_),
    .B(_00846_),
    .Y(_00847_));
 sg13g2_buf_2 _06052_ (.A(_00847_),
    .X(_00848_));
 sg13g2_nand3_1 _06053_ (.B(_00842_),
    .C(_00848_),
    .A(net360),
    .Y(_00849_));
 sg13g2_buf_4 _06054_ (.X(_00850_),
    .A(\game_logic_inst.lfsr_shift[0] ));
 sg13g2_buf_2 _06055_ (.A(\game_logic_inst.lfsr_shift[1] ),
    .X(_00851_));
 sg13g2_mux4_1 _06056_ (.S0(_00850_),
    .A0(\game_logic_inst.lfsr_value[2] ),
    .A1(\game_logic_inst.lfsr_value[6] ),
    .A2(\game_logic_inst.lfsr_value[10] ),
    .A3(\game_logic_inst.lfsr_value[14] ),
    .S1(_00851_),
    .X(_00852_));
 sg13g2_buf_2 _06057_ (.A(_00852_),
    .X(_00853_));
 sg13g2_mux4_1 _06058_ (.S0(_00850_),
    .A0(\game_logic_inst.lfsr_value[1] ),
    .A1(\game_logic_inst.lfsr_value[5] ),
    .A2(\game_logic_inst.lfsr_value[9] ),
    .A3(\game_logic_inst.lfsr_value[13] ),
    .S1(_00851_),
    .X(_00854_));
 sg13g2_buf_2 _06059_ (.A(_00854_),
    .X(_00855_));
 sg13g2_inv_1 _06060_ (.Y(_00856_),
    .A(_00855_));
 sg13g2_mux4_1 _06061_ (.S0(_00850_),
    .A0(\game_logic_inst.lfsr_value[0] ),
    .A1(\game_logic_inst.lfsr_value[4] ),
    .A2(\game_logic_inst.lfsr_value[8] ),
    .A3(\game_logic_inst.lfsr_value[12] ),
    .S1(_00851_),
    .X(_00857_));
 sg13g2_buf_4 _06062_ (.X(_00858_),
    .A(_00857_));
 sg13g2_inv_1 _06063_ (.Y(_00859_),
    .A(_00858_));
 sg13g2_nand2_1 _06064_ (.Y(_00860_),
    .A(_00856_),
    .B(_00859_));
 sg13g2_buf_2 _06065_ (.A(_00860_),
    .X(_00861_));
 sg13g2_mux4_1 _06066_ (.S0(_00850_),
    .A0(\game_logic_inst.lfsr_value[3] ),
    .A1(\game_logic_inst.lfsr_value[7] ),
    .A2(\game_logic_inst.lfsr_value[11] ),
    .A3(\game_logic_inst.lfsr_value[15] ),
    .S1(_00851_),
    .X(_00862_));
 sg13g2_buf_1 _06067_ (.A(_00862_),
    .X(_00863_));
 sg13g2_nor2_1 _06068_ (.A(\game_logic_inst.add_new_tiles[0] ),
    .B(\game_logic_inst.add_new_tiles[1] ),
    .Y(_00864_));
 sg13g2_nor4_1 _06069_ (.A(_00471_),
    .B(_05128_),
    .C(_05211_),
    .D(_05171_),
    .Y(_00865_));
 sg13g2_nor4_1 _06070_ (.A(_00472_),
    .B(_05129_),
    .C(_05212_),
    .D(_05172_),
    .Y(_00866_));
 sg13g2_nor4_1 _06071_ (.A(_05208_),
    .B(_05132_),
    .C(_05205_),
    .D(_05175_),
    .Y(_00867_));
 sg13g2_nor4_1 _06072_ (.A(_05207_),
    .B(_05131_),
    .C(_05204_),
    .D(_05174_),
    .Y(_00868_));
 sg13g2_mux4_1 _06073_ (.S0(_00858_),
    .A0(_00865_),
    .A1(_00866_),
    .A2(_00867_),
    .A3(_00868_),
    .S1(_00855_),
    .X(_00869_));
 sg13g2_nor4_1 _06074_ (.A(_05222_),
    .B(_05225_),
    .C(_05184_),
    .D(_05152_),
    .Y(_00870_));
 sg13g2_nor4_1 _06075_ (.A(_05223_),
    .B(_05226_),
    .C(_05185_),
    .D(_05153_),
    .Y(_00871_));
 sg13g2_nor4_1 _06076_ (.A(_05142_),
    .B(_05188_),
    .C(_00463_),
    .D(_05145_),
    .Y(_00872_));
 sg13g2_nor4_1 _06077_ (.A(_05141_),
    .B(_05187_),
    .C(_00462_),
    .D(_05144_),
    .Y(_00873_));
 sg13g2_mux4_1 _06078_ (.S0(_00858_),
    .A0(_00870_),
    .A1(_00871_),
    .A2(_00872_),
    .A3(_00873_),
    .S1(_00855_),
    .X(_00874_));
 sg13g2_nor4_1 _06079_ (.A(_00468_),
    .B(_05122_),
    .C(_05201_),
    .D(_05165_),
    .Y(_00875_));
 sg13g2_nor4_1 _06080_ (.A(_00469_),
    .B(_05123_),
    .C(_05202_),
    .D(_05166_),
    .Y(_00876_));
 sg13g2_nor4_1 _06081_ (.A(_05198_),
    .B(_05126_),
    .C(_05195_),
    .D(_05169_),
    .Y(_00877_));
 sg13g2_nor4_1 _06082_ (.A(_05197_),
    .B(_05125_),
    .C(_05194_),
    .D(_05168_),
    .Y(_00878_));
 sg13g2_mux4_1 _06083_ (.S0(_00858_),
    .A0(_00875_),
    .A1(_00876_),
    .A2(_00877_),
    .A3(_00878_),
    .S1(_00855_),
    .X(_00879_));
 sg13g2_nor4_1 _06084_ (.A(_05215_),
    .B(_05218_),
    .C(_05178_),
    .D(_05149_),
    .Y(_00880_));
 sg13g2_nor4_1 _06085_ (.A(_05216_),
    .B(_05219_),
    .C(_05179_),
    .D(_05150_),
    .Y(_00881_));
 sg13g2_nor4_1 _06086_ (.A(_05161_),
    .B(_05182_),
    .C(_00460_),
    .D(_05158_),
    .Y(_00882_));
 sg13g2_nor4_1 _06087_ (.A(_05160_),
    .B(_05181_),
    .C(_00459_),
    .D(_05157_),
    .Y(_00883_));
 sg13g2_mux4_1 _06088_ (.S0(_00858_),
    .A0(_00880_),
    .A1(_00881_),
    .A2(_00882_),
    .A3(_00883_),
    .S1(_00855_),
    .X(_00884_));
 sg13g2_inv_1 _06089_ (.Y(_00885_),
    .A(_00853_));
 sg13g2_inv_1 _06090_ (.Y(_00886_),
    .A(_00863_));
 sg13g2_mux4_1 _06091_ (.S0(_00885_),
    .A0(_00869_),
    .A1(_00874_),
    .A2(_00879_),
    .A3(_00884_),
    .S1(_00886_),
    .X(_00887_));
 sg13g2_nand2b_1 _06092_ (.Y(_00888_),
    .B(_00887_),
    .A_N(_00864_));
 sg13g2_buf_1 _06093_ (.A(_00888_),
    .X(_00889_));
 sg13g2_nor4_1 _06094_ (.A(_00853_),
    .B(_00861_),
    .C(_00863_),
    .D(_00889_),
    .Y(_00890_));
 sg13g2_o21ai_1 _06095_ (.B1(_00848_),
    .Y(_00891_),
    .A1(_05100_),
    .A2(_00890_));
 sg13g2_buf_1 _06096_ (.A(_00891_),
    .X(_00892_));
 sg13g2_a21oi_1 _06097_ (.A1(_00098_),
    .A2(_00892_),
    .Y(_00893_),
    .B1(net457));
 sg13g2_nand2_1 _06098_ (.Y(_00894_),
    .A(_00849_),
    .B(_00893_));
 sg13g2_buf_1 _06099_ (.A(\debug_controller_inst.grid_out_data[0] ),
    .X(_00895_));
 sg13g2_buf_1 _06100_ (.A(_00895_),
    .X(_00896_));
 sg13g2_nand2_1 _06101_ (.Y(_00897_),
    .A(_00896_),
    .B(_05098_));
 sg13g2_o21ai_1 _06102_ (.B1(_00897_),
    .Y(_00003_),
    .A1(_05098_),
    .A2(_00894_));
 sg13g2_inv_1 _06103_ (.Y(_00898_),
    .A(_00100_));
 sg13g2_nor2_1 _06104_ (.A(net262),
    .B(net161),
    .Y(_00899_));
 sg13g2_buf_1 _06105_ (.A(_00899_),
    .X(_00900_));
 sg13g2_nand2b_1 _06106_ (.Y(_00901_),
    .B(_00799_),
    .A_N(_00761_));
 sg13g2_a21o_1 _06107_ (.A2(_00749_),
    .A1(_00732_),
    .B1(_00901_),
    .X(_00902_));
 sg13g2_and4_1 _06108_ (.A(_00753_),
    .B(_00761_),
    .C(_00793_),
    .D(_00799_),
    .X(_00903_));
 sg13g2_nand3_1 _06109_ (.B(_00749_),
    .C(_00903_),
    .A(_00732_),
    .Y(_00904_));
 sg13g2_or2_1 _06110_ (.X(_00905_),
    .B(_00901_),
    .A(_00762_));
 sg13g2_nor2_1 _06111_ (.A(_00761_),
    .B(_00793_),
    .Y(_00906_));
 sg13g2_a21oi_2 _06112_ (.B1(_00776_),
    .Y(_00907_),
    .A2(net34),
    .A1(_00678_));
 sg13g2_nor2_1 _06113_ (.A(_00761_),
    .B(_00907_),
    .Y(_00908_));
 sg13g2_a221oi_1 _06114_ (.B2(_00799_),
    .C1(_00908_),
    .B1(_00906_),
    .A1(net51),
    .Y(_00909_),
    .A2(_00769_));
 sg13g2_and4_1 _06115_ (.A(_00902_),
    .B(_00904_),
    .C(_00905_),
    .D(_00909_),
    .X(_00910_));
 sg13g2_buf_1 _06116_ (.A(_00910_),
    .X(_00911_));
 sg13g2_a22oi_1 _06117_ (.Y(_00912_),
    .B1(_00911_),
    .B2(net160),
    .A2(net32),
    .A1(_00751_));
 sg13g2_buf_2 _06118_ (.A(_00912_),
    .X(_00913_));
 sg13g2_nand3b_1 _06119_ (.B(_00848_),
    .C(net70),
    .Y(_00914_),
    .A_N(_00913_));
 sg13g2_o21ai_1 _06120_ (.B1(_00914_),
    .Y(_00915_),
    .A1(_00100_),
    .A2(net70));
 sg13g2_a22oi_1 _06121_ (.Y(_00916_),
    .B1(_00915_),
    .B2(net360),
    .A2(_00892_),
    .A1(_00898_));
 sg13g2_buf_1 _06122_ (.A(_05057_),
    .X(_00917_));
 sg13g2_buf_1 _06123_ (.A(_00917_),
    .X(_00918_));
 sg13g2_buf_1 _06124_ (.A(net452),
    .X(_00919_));
 sg13g2_nand2b_1 _06125_ (.Y(_00920_),
    .B(net407),
    .A_N(_05098_));
 sg13g2_buf_1 _06126_ (.A(\debug_controller_inst.grid_out_data[1] ),
    .X(_00921_));
 sg13g2_buf_1 _06127_ (.A(_00921_),
    .X(_00922_));
 sg13g2_nand2_1 _06128_ (.Y(_00923_),
    .A(net451),
    .B(_05098_));
 sg13g2_o21ai_1 _06129_ (.B1(_00923_),
    .Y(_00014_),
    .A1(_00916_),
    .A2(_00920_));
 sg13g2_inv_1 _06130_ (.Y(_00924_),
    .A(_00101_));
 sg13g2_and2_1 _06131_ (.A(_00761_),
    .B(_00793_),
    .X(_00925_));
 sg13g2_buf_1 _06132_ (.A(_00925_),
    .X(_00926_));
 sg13g2_nand4_1 _06133_ (.B(_00749_),
    .C(_00753_),
    .A(_00732_),
    .Y(_00927_),
    .D(_00926_));
 sg13g2_buf_2 _06134_ (.A(_00927_),
    .X(_00928_));
 sg13g2_inv_1 _06135_ (.Y(_00929_),
    .A(_00689_));
 sg13g2_nor3_1 _06136_ (.A(_00646_),
    .B(net37),
    .C(_00929_),
    .Y(_00930_));
 sg13g2_and2_1 _06137_ (.A(net37),
    .B(_00689_),
    .X(_00931_));
 sg13g2_inv_1 _06138_ (.Y(_00932_),
    .A(_00690_));
 sg13g2_a221oi_1 _06139_ (.B2(_00648_),
    .C1(_00932_),
    .B1(_00931_),
    .A1(_00681_),
    .Y(_00933_),
    .A2(_00930_));
 sg13g2_buf_2 _06140_ (.A(_00933_),
    .X(_00934_));
 sg13g2_xnor2_1 _06141_ (.Y(_00935_),
    .A(_00928_),
    .B(_00934_));
 sg13g2_buf_1 _06142_ (.A(net158),
    .X(_00936_));
 sg13g2_nor2_1 _06143_ (.A(net93),
    .B(_00789_),
    .Y(_00937_));
 sg13g2_and2_1 _06144_ (.A(_00670_),
    .B(_00769_),
    .X(_00938_));
 sg13g2_a21o_1 _06145_ (.A2(_00934_),
    .A1(_00777_),
    .B1(_00938_),
    .X(_00939_));
 sg13g2_nand2_1 _06146_ (.Y(_00940_),
    .A(_00667_),
    .B(net32));
 sg13g2_mux2_1 _06147_ (.A0(_00939_),
    .A1(_00940_),
    .S(net93),
    .X(_00941_));
 sg13g2_a21oi_2 _06148_ (.B1(_00941_),
    .Y(_00942_),
    .A2(_00937_),
    .A1(_00935_));
 sg13g2_nand3_1 _06149_ (.B(_00848_),
    .C(_00942_),
    .A(net70),
    .Y(_00943_));
 sg13g2_o21ai_1 _06150_ (.B1(_00943_),
    .Y(_00944_),
    .A1(_00101_),
    .A2(_00900_));
 sg13g2_a22oi_1 _06151_ (.Y(_00945_),
    .B1(_00944_),
    .B2(net360),
    .A2(_00892_),
    .A1(_00924_));
 sg13g2_buf_1 _06152_ (.A(\debug_controller_inst.grid_out_data[2] ),
    .X(_00946_));
 sg13g2_nand2_1 _06153_ (.Y(_00947_),
    .A(net477),
    .B(_05098_));
 sg13g2_o21ai_1 _06154_ (.B1(_00947_),
    .Y(_00025_),
    .A1(_00920_),
    .A2(_00945_));
 sg13g2_buf_1 _06155_ (.A(\debug_controller_inst.grid_out_data[3] ),
    .X(_00948_));
 sg13g2_buf_1 _06156_ (.A(net93),
    .X(_00949_));
 sg13g2_nand3_1 _06157_ (.B(_00788_),
    .C(_00934_),
    .A(net33),
    .Y(_00950_));
 sg13g2_and2_1 _06158_ (.A(_00736_),
    .B(_00769_),
    .X(_00951_));
 sg13g2_a21oi_1 _06159_ (.A1(net33),
    .A2(_00777_),
    .Y(_00952_),
    .B1(_00951_));
 sg13g2_nand2_1 _06160_ (.Y(_00953_),
    .A(_00950_),
    .B(_00952_));
 sg13g2_inv_1 _06161_ (.Y(_00954_),
    .A(_00934_));
 sg13g2_nand3b_1 _06162_ (.B(_00799_),
    .C(_00954_),
    .Y(_00955_),
    .A_N(net33));
 sg13g2_nand2_1 _06163_ (.Y(_00956_),
    .A(net33),
    .B(_00799_));
 sg13g2_mux2_1 _06164_ (.A0(_00955_),
    .A1(_00956_),
    .S(_00928_),
    .X(_00957_));
 sg13g2_buf_2 _06165_ (.A(_00957_),
    .X(_00958_));
 sg13g2_nand2b_1 _06166_ (.Y(_00959_),
    .B(_00958_),
    .A_N(_00953_));
 sg13g2_nand3_1 _06167_ (.B(_00548_),
    .C(net32),
    .A(net69),
    .Y(_00960_));
 sg13g2_o21ai_1 _06168_ (.B1(_00960_),
    .Y(_00961_),
    .A1(net69),
    .A2(_00959_));
 sg13g2_buf_1 _06169_ (.A(_00961_),
    .X(_00962_));
 sg13g2_nand4_1 _06170_ (.B(_00900_),
    .C(_00848_),
    .A(net360),
    .Y(_00963_),
    .D(_00962_));
 sg13g2_inv_1 _06171_ (.Y(_00964_),
    .A(_00102_));
 sg13g2_nor2b_1 _06172_ (.A(_00102_),
    .B_N(_05101_),
    .Y(_00965_));
 sg13g2_a22oi_1 _06173_ (.Y(_00966_),
    .B1(_00965_),
    .B2(_05115_),
    .A2(_00892_),
    .A1(_00964_));
 sg13g2_a21oi_1 _06174_ (.A1(_00963_),
    .A2(_00966_),
    .Y(_00967_),
    .B1(_00920_));
 sg13g2_a21o_1 _06175_ (.A2(_05098_),
    .A1(_00948_),
    .B1(_00967_),
    .X(_00036_));
 sg13g2_buf_1 _06176_ (.A(_05095_),
    .X(_00968_));
 sg13g2_nor2_2 _06177_ (.A(_05093_),
    .B(_05094_),
    .Y(_00969_));
 sg13g2_nand2_2 _06178_ (.Y(_00970_),
    .A(_00968_),
    .B(_00969_));
 sg13g2_inv_1 _06179_ (.Y(_00971_),
    .A(\debug_controller_inst.grid_out_valid ));
 sg13g2_inv_2 _06180_ (.Y(_00972_),
    .A(_05095_));
 sg13g2_o21ai_1 _06181_ (.B1(_00969_),
    .Y(_00973_),
    .A1(_00972_),
    .A2(_00099_));
 sg13g2_a21o_1 _06182_ (.A2(_00969_),
    .A1(_00099_),
    .B1(_05092_),
    .X(_00974_));
 sg13g2_o21ai_1 _06183_ (.B1(_00974_),
    .Y(_00975_),
    .A1(_05091_),
    .A2(_00973_));
 sg13g2_nor2_1 _06184_ (.A(_00971_),
    .B(_00975_),
    .Y(_00976_));
 sg13g2_buf_1 _06185_ (.A(_00976_),
    .X(_00977_));
 sg13g2_buf_1 _06186_ (.A(_00977_),
    .X(_00978_));
 sg13g2_nand2_2 _06187_ (.Y(_00979_),
    .A(_00895_),
    .B(_00978_));
 sg13g2_buf_1 _06188_ (.A(_00846_),
    .X(_00980_));
 sg13g2_buf_1 _06189_ (.A(net50),
    .X(_00981_));
 sg13g2_buf_1 _06190_ (.A(net46),
    .X(_00982_));
 sg13g2_buf_1 _06191_ (.A(_00843_),
    .X(_00983_));
 sg13g2_buf_1 _06192_ (.A(net449),
    .X(_00984_));
 sg13g2_nand2b_1 _06193_ (.Y(_00985_),
    .B(_05099_),
    .A_N(_00843_));
 sg13g2_buf_1 _06194_ (.A(_00985_),
    .X(_00986_));
 sg13g2_buf_1 _06195_ (.A(_00986_),
    .X(_00987_));
 sg13g2_nor2_2 _06196_ (.A(net75),
    .B(net353),
    .Y(_00988_));
 sg13g2_xnor2_1 _06197_ (.Y(_00989_),
    .A(_00642_),
    .B(_00812_));
 sg13g2_nor2_1 _06198_ (.A(_00581_),
    .B(net35),
    .Y(_00990_));
 sg13g2_a22oi_1 _06199_ (.Y(_00991_),
    .B1(_00990_),
    .B2(net34),
    .A2(_00989_),
    .A1(net44));
 sg13g2_buf_1 _06200_ (.A(_00991_),
    .X(_00992_));
 sg13g2_a21oi_1 _06201_ (.A1(_05119_),
    .A2(_00628_),
    .Y(_00993_),
    .B1(_00631_));
 sg13g2_inv_1 _06202_ (.Y(_00994_),
    .A(_00642_));
 sg13g2_nor4_1 _06203_ (.A(_00507_),
    .B(_00993_),
    .C(_00994_),
    .D(_00812_),
    .Y(_00995_));
 sg13g2_xnor2_1 _06204_ (.Y(_00996_),
    .A(_00516_),
    .B(_00995_));
 sg13g2_and2_1 _06205_ (.A(_00671_),
    .B(_00996_),
    .X(_00997_));
 sg13g2_buf_1 _06206_ (.A(_00997_),
    .X(_00998_));
 sg13g2_nor2_1 _06207_ (.A(_00815_),
    .B(_00998_),
    .Y(_00999_));
 sg13g2_nor2_1 _06208_ (.A(_00656_),
    .B(_00671_),
    .Y(_01000_));
 sg13g2_a221oi_1 _06209_ (.B2(net36),
    .C1(_00815_),
    .B1(_00996_),
    .A1(net71),
    .Y(_01001_),
    .A2(_01000_));
 sg13g2_a21oi_1 _06210_ (.A1(_00729_),
    .A2(_00999_),
    .Y(_01002_),
    .B1(_01001_));
 sg13g2_nor2_1 _06211_ (.A(net35),
    .B(_00820_),
    .Y(_01003_));
 sg13g2_a22oi_1 _06212_ (.Y(_01004_),
    .B1(_01003_),
    .B2(net34),
    .A2(_00998_),
    .A1(_00815_));
 sg13g2_a22oi_1 _06213_ (.Y(_01005_),
    .B1(_00721_),
    .B2(net72),
    .A2(_00670_),
    .A1(net159));
 sg13g2_nor2_1 _06214_ (.A(_00661_),
    .B(_01005_),
    .Y(_01006_));
 sg13g2_nor2_1 _06215_ (.A(_00507_),
    .B(_00667_),
    .Y(_01007_));
 sg13g2_a21oi_1 _06216_ (.A1(_00642_),
    .A2(_00721_),
    .Y(_01008_),
    .B1(_01007_));
 sg13g2_a21oi_1 _06217_ (.A1(_00813_),
    .A2(_01008_),
    .Y(_01009_),
    .B1(_00773_));
 sg13g2_a21o_1 _06218_ (.A2(_01006_),
    .A1(net34),
    .B1(_01009_),
    .X(_01010_));
 sg13g2_a221oi_1 _06219_ (.B2(_01004_),
    .C1(_01010_),
    .B1(_01002_),
    .A1(_00713_),
    .Y(_01011_),
    .A2(_00992_));
 sg13g2_buf_1 _06220_ (.A(_01011_),
    .X(_01012_));
 sg13g2_buf_1 _06221_ (.A(_01012_),
    .X(_01013_));
 sg13g2_nor2_1 _06222_ (.A(_00687_),
    .B(_00660_),
    .Y(_01014_));
 sg13g2_nor3_1 _06223_ (.A(_00993_),
    .B(_00994_),
    .C(_00812_),
    .Y(_01015_));
 sg13g2_xor2_1 _06224_ (.B(_01015_),
    .A(_00507_),
    .X(_01016_));
 sg13g2_nor2_1 _06225_ (.A(_00773_),
    .B(_01016_),
    .Y(_01017_));
 sg13g2_a21oi_2 _06226_ (.B1(_01017_),
    .Y(_01018_),
    .A2(_01014_),
    .A1(net34));
 sg13g2_nor2_1 _06227_ (.A(_00994_),
    .B(_00812_),
    .Y(_01019_));
 sg13g2_nor2_1 _06228_ (.A(_00632_),
    .B(_01019_),
    .Y(_01020_));
 sg13g2_nor4_2 _06229_ (.A(_00595_),
    .B(net57),
    .C(_01015_),
    .Y(_01021_),
    .D(_01020_));
 sg13g2_nand2b_1 _06230_ (.Y(_01022_),
    .B(net51),
    .A_N(_01021_));
 sg13g2_nand3b_1 _06231_ (.B(_00753_),
    .C(net54),
    .Y(_01023_),
    .A_N(net35));
 sg13g2_mux2_1 _06232_ (.A0(_01022_),
    .A1(_01023_),
    .S(net34),
    .X(_01024_));
 sg13g2_nand2_1 _06233_ (.Y(_01025_),
    .A(_00637_),
    .B(net51));
 sg13g2_nand2_1 _06234_ (.Y(_01026_),
    .A(_00660_),
    .B(net51));
 sg13g2_a21oi_1 _06235_ (.A1(_01025_),
    .A2(_01026_),
    .Y(_01027_),
    .B1(_01021_));
 sg13g2_a21oi_1 _06236_ (.A1(_00753_),
    .A2(_01021_),
    .Y(_01028_),
    .B1(_01027_));
 sg13g2_a22oi_1 _06237_ (.Y(_01029_),
    .B1(_01024_),
    .B2(_01028_),
    .A2(_01018_),
    .A1(net55));
 sg13g2_buf_2 _06238_ (.A(_01029_),
    .X(_01030_));
 sg13g2_xnor2_1 _06239_ (.Y(_01031_),
    .A(net52),
    .B(net56));
 sg13g2_nor2_1 _06240_ (.A(_00682_),
    .B(_01031_),
    .Y(_01032_));
 sg13g2_a21o_1 _06241_ (.A2(_00813_),
    .A1(_00685_),
    .B1(_00773_),
    .X(_01033_));
 sg13g2_o21ai_1 _06242_ (.B1(_01033_),
    .Y(_01034_),
    .A1(_00682_),
    .A2(_00706_));
 sg13g2_a21o_1 _06243_ (.A2(_01032_),
    .A1(_00705_),
    .B1(_01034_),
    .X(_01035_));
 sg13g2_buf_1 _06244_ (.A(_01035_),
    .X(_01036_));
 sg13g2_nand2_1 _06245_ (.Y(_01037_),
    .A(_00713_),
    .B(net31));
 sg13g2_a21oi_1 _06246_ (.A1(net30),
    .A2(_01030_),
    .Y(_01038_),
    .B1(_01037_));
 sg13g2_and4_1 _06247_ (.A(_00817_),
    .B(_00818_),
    .C(_00822_),
    .D(_00823_),
    .X(_01039_));
 sg13g2_buf_1 _06248_ (.A(_01039_),
    .X(_01040_));
 sg13g2_a21oi_1 _06249_ (.A1(_00825_),
    .A2(_00826_),
    .Y(_01041_),
    .B1(_00831_));
 sg13g2_nor3_2 _06250_ (.A(_00581_),
    .B(_01040_),
    .C(_01041_),
    .Y(_01042_));
 sg13g2_o21ai_1 _06251_ (.B1(_00581_),
    .Y(_01043_),
    .A1(_01040_),
    .A2(_01041_));
 sg13g2_nand2_2 _06252_ (.Y(_01044_),
    .A(net36),
    .B(net41));
 sg13g2_nor2_1 _06253_ (.A(net43),
    .B(_01044_),
    .Y(_01045_));
 sg13g2_nand3b_1 _06254_ (.B(_01043_),
    .C(_01045_),
    .Y(_01046_),
    .A_N(_01042_));
 sg13g2_nand2b_1 _06255_ (.Y(_01047_),
    .B(_01046_),
    .A_N(_01038_));
 sg13g2_buf_1 _06256_ (.A(_01047_),
    .X(_01048_));
 sg13g2_nand3_1 _06257_ (.B(_00749_),
    .C(_00762_),
    .A(_00732_),
    .Y(_01049_));
 sg13g2_buf_2 _06258_ (.A(_01049_),
    .X(_01050_));
 sg13g2_a22oi_1 _06259_ (.Y(_01051_),
    .B1(_00784_),
    .B2(_00705_),
    .A2(_00782_),
    .A1(_00781_));
 sg13g2_nand2b_1 _06260_ (.Y(_01052_),
    .B(_01051_),
    .A_N(_00786_));
 sg13g2_nor2_1 _06261_ (.A(_00721_),
    .B(_01052_),
    .Y(_01053_));
 sg13g2_inv_1 _06262_ (.Y(_01054_),
    .A(_00992_));
 sg13g2_a21o_1 _06263_ (.A2(_01030_),
    .A1(_01012_),
    .B1(_01054_),
    .X(_01055_));
 sg13g2_a221oi_1 _06264_ (.B2(_01028_),
    .C1(_00992_),
    .B1(_01024_),
    .A1(net55),
    .Y(_01056_),
    .A2(_01018_));
 sg13g2_buf_2 _06265_ (.A(_01056_),
    .X(_01057_));
 sg13g2_a21oi_2 _06266_ (.B1(_01034_),
    .Y(_01058_),
    .A2(_01032_),
    .A1(_00705_));
 sg13g2_a21oi_1 _06267_ (.A1(_01013_),
    .A2(_01057_),
    .Y(_01059_),
    .B1(_01058_));
 sg13g2_and2_1 _06268_ (.A(_00796_),
    .B(_00835_),
    .X(_01060_));
 sg13g2_buf_1 _06269_ (.A(_01060_),
    .X(_01061_));
 sg13g2_nor2_1 _06270_ (.A(_01061_),
    .B(_00992_),
    .Y(_01062_));
 sg13g2_a221oi_1 _06271_ (.B2(_01059_),
    .C1(_01062_),
    .B1(_01055_),
    .A1(_01050_),
    .Y(_01063_),
    .A2(_01053_));
 sg13g2_buf_2 _06272_ (.A(_01063_),
    .X(_01064_));
 sg13g2_nand2_1 _06273_ (.Y(_01065_),
    .A(net94),
    .B(_01064_));
 sg13g2_o21ai_1 _06274_ (.B1(_01065_),
    .Y(_01066_),
    .A1(_05121_),
    .A2(_01048_));
 sg13g2_buf_2 _06275_ (.A(_01066_),
    .X(_01067_));
 sg13g2_nand2_2 _06276_ (.Y(_01068_),
    .A(_00856_),
    .B(_00858_));
 sg13g2_xnor2_1 _06277_ (.Y(_01069_),
    .A(_00861_),
    .B(_00863_));
 sg13g2_nor3_2 _06278_ (.A(_00853_),
    .B(_00889_),
    .C(_01069_),
    .Y(_01070_));
 sg13g2_nand2b_1 _06279_ (.Y(_01071_),
    .B(_01070_),
    .A_N(_01068_));
 sg13g2_nor2_1 _06280_ (.A(_00843_),
    .B(_05099_),
    .Y(_01072_));
 sg13g2_buf_2 _06281_ (.A(_01072_),
    .X(_01073_));
 sg13g2_buf_1 _06282_ (.A(_01073_),
    .X(_01074_));
 sg13g2_and3_1 _06283_ (.X(_01075_),
    .A(_00103_),
    .B(_01071_),
    .C(net352));
 sg13g2_a221oi_1 _06284_ (.B2(_01067_),
    .C1(_01075_),
    .B1(_00988_),
    .A1(net406),
    .Y(_01076_),
    .A2(_00104_));
 sg13g2_inv_1 _06285_ (.Y(_01077_),
    .A(_05063_));
 sg13g2_nor2_1 _06286_ (.A(_01077_),
    .B(_05078_),
    .Y(_01078_));
 sg13g2_buf_2 _06287_ (.A(_01078_),
    .X(_01079_));
 sg13g2_o21ai_1 _06288_ (.B1(_01079_),
    .Y(_01080_),
    .A1(_00899_),
    .A2(_00986_));
 sg13g2_buf_2 _06289_ (.A(_01080_),
    .X(_01081_));
 sg13g2_and2_1 _06290_ (.A(_05095_),
    .B(_00969_),
    .X(_01082_));
 sg13g2_buf_1 _06291_ (.A(_01082_),
    .X(_01083_));
 sg13g2_nand2_1 _06292_ (.Y(_01084_),
    .A(_01083_),
    .B(_00977_));
 sg13g2_nand2_1 _06293_ (.Y(_01085_),
    .A(net452),
    .B(_01084_));
 sg13g2_a21oi_1 _06294_ (.A1(_00103_),
    .A2(_01081_),
    .Y(_01086_),
    .B1(_01085_));
 sg13g2_o21ai_1 _06295_ (.B1(_01086_),
    .Y(_01087_),
    .A1(net40),
    .A2(_01076_));
 sg13g2_o21ai_1 _06296_ (.B1(_01087_),
    .Y(_00047_),
    .A1(_00970_),
    .A2(_00979_));
 sg13g2_nor2b_1 _06297_ (.A(_00843_),
    .B_N(net456),
    .Y(_01088_));
 sg13g2_buf_1 _06298_ (.A(_01088_),
    .X(_01089_));
 sg13g2_nand2_1 _06299_ (.Y(_01090_),
    .A(_00899_),
    .B(net351));
 sg13g2_nor2_1 _06300_ (.A(_00637_),
    .B(net35),
    .Y(_01091_));
 sg13g2_a21oi_2 _06301_ (.B1(_01021_),
    .Y(_01092_),
    .A2(_01091_),
    .A1(_00771_));
 sg13g2_nor2_1 _06302_ (.A(_00768_),
    .B(_01092_),
    .Y(_01093_));
 sg13g2_and4_1 _06303_ (.A(_01036_),
    .B(net30),
    .C(_01057_),
    .D(_01093_),
    .X(_01094_));
 sg13g2_nand2_1 _06304_ (.Y(_01095_),
    .A(net31),
    .B(_01092_));
 sg13g2_a21oi_1 _06305_ (.A1(net30),
    .A2(_01057_),
    .Y(_01096_),
    .B1(_01095_));
 sg13g2_and4_1 _06306_ (.A(_00732_),
    .B(_00749_),
    .C(_00761_),
    .D(_00799_),
    .X(_01097_));
 sg13g2_nand2_1 _06307_ (.Y(_01098_),
    .A(_00796_),
    .B(_00835_));
 sg13g2_nand2_1 _06308_ (.Y(_01099_),
    .A(_01098_),
    .B(_01092_));
 sg13g2_o21ai_1 _06309_ (.B1(_01099_),
    .Y(_01100_),
    .A1(_00753_),
    .A2(_00789_));
 sg13g2_nor4_2 _06310_ (.A(_01094_),
    .B(_01096_),
    .C(_01097_),
    .Y(_01101_),
    .D(_01100_));
 sg13g2_a21o_1 _06311_ (.A2(_01030_),
    .A1(net30),
    .B1(_00765_),
    .X(_01102_));
 sg13g2_nand3b_1 _06312_ (.B(net42),
    .C(_00775_),
    .Y(_01103_),
    .A_N(net35));
 sg13g2_nand2_1 _06313_ (.Y(_01104_),
    .A(_00785_),
    .B(_00775_));
 sg13g2_o21ai_1 _06314_ (.B1(_01104_),
    .Y(_01105_),
    .A1(_00729_),
    .A2(_01103_));
 sg13g2_a21o_1 _06315_ (.A2(_01042_),
    .A1(_00637_),
    .B1(_01044_),
    .X(_01106_));
 sg13g2_nor2_1 _06316_ (.A(net42),
    .B(_00768_),
    .Y(_01107_));
 sg13g2_a22oi_1 _06317_ (.Y(_01108_),
    .B1(_00834_),
    .B2(net54),
    .A2(_01107_),
    .A1(net36));
 sg13g2_nor2_1 _06318_ (.A(_01042_),
    .B(_01108_),
    .Y(_01109_));
 sg13g2_a21oi_2 _06319_ (.B1(_01109_),
    .Y(_01110_),
    .A2(_01106_),
    .A1(_01105_));
 sg13g2_or2_1 _06320_ (.X(_01111_),
    .B(_01110_),
    .A(net260));
 sg13g2_a21oi_1 _06321_ (.A1(net31),
    .A2(_01102_),
    .Y(_01112_),
    .B1(_01111_));
 sg13g2_a21o_1 _06322_ (.A2(_01101_),
    .A1(net94),
    .B1(_01112_),
    .X(_01113_));
 sg13g2_buf_1 _06323_ (.A(_01113_),
    .X(_01114_));
 sg13g2_nand2b_1 _06324_ (.Y(_01115_),
    .B(_01071_),
    .A_N(_00105_));
 sg13g2_a22oi_1 _06325_ (.Y(_01116_),
    .B1(net352),
    .B2(_01115_),
    .A2(_00106_),
    .A1(net449));
 sg13g2_o21ai_1 _06326_ (.B1(_01116_),
    .Y(_01117_),
    .A1(_01090_),
    .A2(_01114_));
 sg13g2_buf_1 _06327_ (.A(_01079_),
    .X(_01118_));
 sg13g2_buf_1 _06328_ (.A(net53),
    .X(_01119_));
 sg13g2_buf_1 _06329_ (.A(net457),
    .X(_01120_));
 sg13g2_a221oi_1 _06330_ (.B2(net49),
    .C1(net405),
    .B1(_01117_),
    .A1(_00105_),
    .Y(_01121_),
    .A2(_01081_));
 sg13g2_mux2_1 _06331_ (.A0(net451),
    .A1(_01121_),
    .S(_01084_),
    .X(_00058_));
 sg13g2_nand2_1 _06332_ (.Y(_01122_),
    .A(net477),
    .B(net92));
 sg13g2_and2_1 _06333_ (.A(_01012_),
    .B(_01057_),
    .X(_01123_));
 sg13g2_a21o_1 _06334_ (.A2(_01014_),
    .A1(net34),
    .B1(_01017_),
    .X(_01124_));
 sg13g2_a21o_1 _06335_ (.A2(_01093_),
    .A1(_01123_),
    .B1(_01124_),
    .X(_01125_));
 sg13g2_nor3_1 _06336_ (.A(_00768_),
    .B(_01018_),
    .C(_01092_),
    .Y(_01126_));
 sg13g2_nand3_1 _06337_ (.B(_01057_),
    .C(_01126_),
    .A(_01012_),
    .Y(_01127_));
 sg13g2_buf_1 _06338_ (.A(_01127_),
    .X(_01128_));
 sg13g2_and2_1 _06339_ (.A(net31),
    .B(_01128_),
    .X(_01129_));
 sg13g2_buf_1 _06340_ (.A(_01129_),
    .X(_01130_));
 sg13g2_nor2_1 _06341_ (.A(_00670_),
    .B(_01052_),
    .Y(_01131_));
 sg13g2_nor2_1 _06342_ (.A(_01061_),
    .B(_01018_),
    .Y(_01132_));
 sg13g2_a221oi_1 _06343_ (.B2(_01050_),
    .C1(_01132_),
    .B1(_01131_),
    .A1(_01125_),
    .Y(_01133_),
    .A2(_01130_));
 sg13g2_and2_1 _06344_ (.A(net30),
    .B(_01030_),
    .X(_01134_));
 sg13g2_nor2_1 _06345_ (.A(_00768_),
    .B(_01058_),
    .Y(_01135_));
 sg13g2_a21o_1 _06346_ (.A2(_00834_),
    .A1(net159),
    .B1(_01105_),
    .X(_01136_));
 sg13g2_nand2_1 _06347_ (.Y(_01137_),
    .A(net54),
    .B(_01042_));
 sg13g2_nand3_1 _06348_ (.B(_01045_),
    .C(_01137_),
    .A(_00687_),
    .Y(_01138_));
 sg13g2_and3_1 _06349_ (.X(_01139_),
    .A(net36),
    .B(net55),
    .C(net41));
 sg13g2_a22oi_1 _06350_ (.Y(_01140_),
    .B1(_01139_),
    .B2(_00713_),
    .A2(_01044_),
    .A1(_00825_));
 sg13g2_nand3_1 _06351_ (.B(net159),
    .C(net54),
    .A(net72),
    .Y(_01141_));
 sg13g2_nor3_2 _06352_ (.A(_01040_),
    .B(_01140_),
    .C(_01141_),
    .Y(_01142_));
 sg13g2_nand2_1 _06353_ (.Y(_01143_),
    .A(_00834_),
    .B(_01142_));
 sg13g2_nand3_1 _06354_ (.B(_00775_),
    .C(net31),
    .A(_00670_),
    .Y(_01144_));
 sg13g2_nand4_1 _06355_ (.B(_01138_),
    .C(_01143_),
    .A(_01136_),
    .Y(_01145_),
    .D(_01144_));
 sg13g2_a21oi_2 _06356_ (.B1(_01145_),
    .Y(_01146_),
    .A2(_01135_),
    .A1(_01134_));
 sg13g2_inv_1 _06357_ (.Y(_01147_),
    .A(_01146_));
 sg13g2_mux2_1 _06358_ (.A0(_01133_),
    .A1(_01147_),
    .S(_00949_),
    .X(_01148_));
 sg13g2_buf_2 _06359_ (.A(_01148_),
    .X(_01149_));
 sg13g2_inv_1 _06360_ (.Y(_01150_),
    .A(_00107_));
 sg13g2_or2_1 _06361_ (.X(_01151_),
    .B(_05099_),
    .A(_00843_));
 sg13g2_buf_2 _06362_ (.A(_01151_),
    .X(_01152_));
 sg13g2_buf_1 _06363_ (.A(_01152_),
    .X(_01153_));
 sg13g2_a21oi_1 _06364_ (.A1(_01150_),
    .A2(_01071_),
    .Y(_01154_),
    .B1(net350));
 sg13g2_a221oi_1 _06365_ (.B2(_01149_),
    .C1(_01154_),
    .B1(_00988_),
    .A1(net406),
    .Y(_01155_),
    .A2(_00108_));
 sg13g2_a21oi_1 _06366_ (.A1(_00107_),
    .A2(_01081_),
    .Y(_01156_),
    .B1(_01085_));
 sg13g2_o21ai_1 _06367_ (.B1(_01156_),
    .Y(_01157_),
    .A1(net40),
    .A2(_01155_));
 sg13g2_o21ai_1 _06368_ (.B1(_01157_),
    .Y(_00063_),
    .A1(_00970_),
    .A2(_01122_));
 sg13g2_nand4_1 _06369_ (.B(_00747_),
    .C(_00762_),
    .A(_00732_),
    .Y(_01158_),
    .D(_00788_));
 sg13g2_nand2_1 _06370_ (.Y(_01159_),
    .A(_00815_),
    .B(_00788_));
 sg13g2_nand4_1 _06371_ (.B(_01013_),
    .C(_01057_),
    .A(_01036_),
    .Y(_01160_),
    .D(_01126_));
 sg13g2_nand3_1 _06372_ (.B(_01159_),
    .C(_01160_),
    .A(_01158_),
    .Y(_01161_));
 sg13g2_nor2_1 _06373_ (.A(_00661_),
    .B(_00729_),
    .Y(_01162_));
 sg13g2_a21oi_1 _06374_ (.A1(_00602_),
    .A2(_01162_),
    .Y(_01163_),
    .B1(_00998_));
 sg13g2_nand2_1 _06375_ (.Y(_01164_),
    .A(_01061_),
    .B(_01163_));
 sg13g2_nor2b_1 _06376_ (.A(_01164_),
    .B_N(_01050_),
    .Y(_01165_));
 sg13g2_a21o_1 _06377_ (.A2(_01128_),
    .A1(net31),
    .B1(_01098_),
    .X(_01166_));
 sg13g2_inv_1 _06378_ (.Y(_01167_),
    .A(_01163_));
 sg13g2_a22oi_1 _06379_ (.Y(_01168_),
    .B1(_01166_),
    .B2(_01167_),
    .A2(_01165_),
    .A1(_01161_));
 sg13g2_buf_1 _06380_ (.A(_01168_),
    .X(_01169_));
 sg13g2_nor2_1 _06381_ (.A(_00700_),
    .B(_00768_),
    .Y(_01170_));
 sg13g2_mux2_1 _06382_ (.A0(_00700_),
    .A1(_01170_),
    .S(_01142_),
    .X(_01171_));
 sg13g2_nor2_1 _06383_ (.A(_01044_),
    .B(_01171_),
    .Y(_01172_));
 sg13g2_a21o_1 _06384_ (.A2(_01030_),
    .A1(net30),
    .B1(_01058_),
    .X(_01173_));
 sg13g2_nor2_1 _06385_ (.A(_00736_),
    .B(_01173_),
    .Y(_01174_));
 sg13g2_nor2_1 _06386_ (.A(_01172_),
    .B(_01174_),
    .Y(_01175_));
 sg13g2_and2_1 _06387_ (.A(net69),
    .B(_01175_),
    .X(_01176_));
 sg13g2_a21oi_2 _06388_ (.B1(_01176_),
    .Y(_01177_),
    .A2(_01169_),
    .A1(net94));
 sg13g2_nor2_1 _06389_ (.A(_01090_),
    .B(_01177_),
    .Y(_01178_));
 sg13g2_nor2b_1 _06390_ (.A(_00109_),
    .B_N(_01071_),
    .Y(_01179_));
 sg13g2_buf_1 _06391_ (.A(_00843_),
    .X(_01180_));
 sg13g2_buf_1 _06392_ (.A(net448),
    .X(_01181_));
 sg13g2_a221oi_1 _06393_ (.B2(_00109_),
    .C1(_01085_),
    .B1(_01081_),
    .A1(net404),
    .Y(_01182_),
    .A2(_00110_));
 sg13g2_o21ai_1 _06394_ (.B1(_01182_),
    .Y(_01183_),
    .A1(net350),
    .A2(_01179_));
 sg13g2_and2_1 _06395_ (.A(net476),
    .B(net92),
    .X(_01184_));
 sg13g2_buf_1 _06396_ (.A(_01184_),
    .X(_01185_));
 sg13g2_buf_1 _06397_ (.A(net53),
    .X(_01186_));
 sg13g2_nor3_1 _06398_ (.A(_00109_),
    .B(net48),
    .C(_01085_),
    .Y(_01187_));
 sg13g2_a21oi_1 _06399_ (.A1(_01083_),
    .A2(_01185_),
    .Y(_01188_),
    .B1(_01187_));
 sg13g2_o21ai_1 _06400_ (.B1(_01188_),
    .Y(_00064_),
    .A1(_01178_),
    .A2(_01183_));
 sg13g2_nor2b_1 _06401_ (.A(_05093_),
    .B_N(_05094_),
    .Y(_01189_));
 sg13g2_nand2_1 _06402_ (.Y(_01190_),
    .A(_00972_),
    .B(_01189_));
 sg13g2_inv_1 _06403_ (.Y(_01191_),
    .A(_01046_));
 sg13g2_nor3_1 _06404_ (.A(net93),
    .B(_01038_),
    .C(_01191_),
    .Y(_01192_));
 sg13g2_a21o_1 _06405_ (.A2(_01064_),
    .A1(net69),
    .B1(_01192_),
    .X(_01193_));
 sg13g2_buf_2 _06406_ (.A(_01193_),
    .X(_01194_));
 sg13g2_nand3_1 _06407_ (.B(_00859_),
    .C(_01070_),
    .A(_00855_),
    .Y(_01195_));
 sg13g2_buf_1 _06408_ (.A(_01195_),
    .X(_01196_));
 sg13g2_and3_1 _06409_ (.X(_01197_),
    .A(_00111_),
    .B(net352),
    .C(_01196_));
 sg13g2_a221oi_1 _06410_ (.B2(_01194_),
    .C1(_01197_),
    .B1(_00988_),
    .A1(net406),
    .Y(_01198_),
    .A2(_00112_));
 sg13g2_nand2b_1 _06411_ (.Y(_01199_),
    .B(_05094_),
    .A_N(_05093_));
 sg13g2_buf_1 _06412_ (.A(_01199_),
    .X(_01200_));
 sg13g2_nor2_2 _06413_ (.A(_00968_),
    .B(_01200_),
    .Y(_01201_));
 sg13g2_nand2_1 _06414_ (.Y(_01202_),
    .A(_00977_),
    .B(_01201_));
 sg13g2_nand2_1 _06415_ (.Y(_01203_),
    .A(net452),
    .B(_01202_));
 sg13g2_a21oi_1 _06416_ (.A1(_00111_),
    .A2(_01081_),
    .Y(_01204_),
    .B1(_01203_));
 sg13g2_o21ai_1 _06417_ (.B1(_01204_),
    .Y(_01205_),
    .A1(net40),
    .A2(_01198_));
 sg13g2_o21ai_1 _06418_ (.B1(_01205_),
    .Y(_00065_),
    .A1(_00979_),
    .A2(_01190_));
 sg13g2_nand2b_1 _06419_ (.Y(_01206_),
    .B(_01196_),
    .A_N(_00113_));
 sg13g2_a22oi_1 _06420_ (.Y(_01207_),
    .B1(_01074_),
    .B2(_01206_),
    .A2(_00114_),
    .A1(_01181_));
 sg13g2_or2_1 _06421_ (.X(_01208_),
    .B(_00558_),
    .A(net355));
 sg13g2_o21ai_1 _06422_ (.B1(_01208_),
    .Y(_01209_),
    .A1(net262),
    .A2(_00559_));
 sg13g2_buf_1 _06423_ (.A(_01209_),
    .X(_01210_));
 sg13g2_a21o_1 _06424_ (.A2(_01030_),
    .A1(net30),
    .B1(_01210_),
    .X(_01211_));
 sg13g2_nand2_1 _06425_ (.Y(_01212_),
    .A(net31),
    .B(_01211_));
 sg13g2_nor2_1 _06426_ (.A(_00936_),
    .B(_01110_),
    .Y(_01213_));
 sg13g2_a22oi_1 _06427_ (.Y(_01214_),
    .B1(_01212_),
    .B2(_01213_),
    .A2(_01101_),
    .A1(_00936_));
 sg13g2_buf_1 _06428_ (.A(_01214_),
    .X(_01215_));
 sg13g2_nand2_1 _06429_ (.Y(_01216_),
    .A(_00988_),
    .B(_01215_));
 sg13g2_nand2_1 _06430_ (.Y(_01217_),
    .A(_01207_),
    .B(_01216_));
 sg13g2_a221oi_1 _06431_ (.B2(net49),
    .C1(_01120_),
    .B1(_01217_),
    .A1(_00113_),
    .Y(_01218_),
    .A2(_01081_));
 sg13g2_mux2_1 _06432_ (.A0(net451),
    .A1(_01218_),
    .S(_01202_),
    .X(_00066_));
 sg13g2_mux2_1 _06433_ (.A0(_01133_),
    .A1(_01147_),
    .S(net94),
    .X(_01219_));
 sg13g2_buf_2 _06434_ (.A(_01219_),
    .X(_01220_));
 sg13g2_inv_1 _06435_ (.Y(_01221_),
    .A(_00115_));
 sg13g2_a21oi_1 _06436_ (.A1(_01221_),
    .A2(_01196_),
    .Y(_01222_),
    .B1(_01153_));
 sg13g2_a221oi_1 _06437_ (.B2(_01220_),
    .C1(_01222_),
    .B1(_00988_),
    .A1(net406),
    .Y(_01223_),
    .A2(_00116_));
 sg13g2_a21oi_1 _06438_ (.A1(_00115_),
    .A2(_01081_),
    .Y(_01224_),
    .B1(_01203_));
 sg13g2_o21ai_1 _06439_ (.B1(_01224_),
    .Y(_01225_),
    .A1(net40),
    .A2(_01223_));
 sg13g2_o21ai_1 _06440_ (.B1(_01225_),
    .Y(_00004_),
    .A1(_01122_),
    .A2(_01190_));
 sg13g2_mux2_1 _06441_ (.A0(_01169_),
    .A1(_01175_),
    .S(_05121_),
    .X(_01226_));
 sg13g2_inv_1 _06442_ (.Y(_01227_),
    .A(_01226_));
 sg13g2_buf_1 _06443_ (.A(net353),
    .X(_01228_));
 sg13g2_a21oi_1 _06444_ (.A1(net70),
    .A2(_01227_),
    .Y(_01229_),
    .B1(_01228_));
 sg13g2_nand2b_1 _06445_ (.Y(_01230_),
    .B(_01196_),
    .A_N(_00117_));
 sg13g2_a221oi_1 _06446_ (.B2(_01230_),
    .C1(net50),
    .B1(_01073_),
    .A1(net448),
    .Y(_01231_),
    .A2(_00118_));
 sg13g2_nand2b_1 _06447_ (.Y(_01232_),
    .B(_01231_),
    .A_N(_01203_));
 sg13g2_buf_1 _06448_ (.A(net50),
    .X(_01233_));
 sg13g2_a21oi_1 _06449_ (.A1(net75),
    .A2(_01231_),
    .Y(_01234_),
    .B1(net45));
 sg13g2_nor3_1 _06450_ (.A(_00117_),
    .B(_01203_),
    .C(_01234_),
    .Y(_01235_));
 sg13g2_a21oi_1 _06451_ (.A1(_01185_),
    .A2(_01201_),
    .Y(_01236_),
    .B1(_01235_));
 sg13g2_o21ai_1 _06452_ (.B1(_01236_),
    .Y(_00005_),
    .A1(_01229_),
    .A2(_01232_));
 sg13g2_nand2b_1 _06453_ (.Y(_01237_),
    .B(\debug_controller_inst.grid_out_valid ),
    .A_N(_00975_));
 sg13g2_buf_1 _06454_ (.A(_01237_),
    .X(_01238_));
 sg13g2_nor3_2 _06455_ (.A(_00972_),
    .B(_01238_),
    .C(_01200_),
    .Y(_01239_));
 sg13g2_buf_1 _06456_ (.A(net45),
    .X(_01240_));
 sg13g2_a22oi_1 _06457_ (.Y(_01241_),
    .B1(net32),
    .B2(_00709_),
    .A2(_00800_),
    .A1(net69));
 sg13g2_buf_1 _06458_ (.A(_01241_),
    .X(_01242_));
 sg13g2_nand2_1 _06459_ (.Y(_01243_),
    .A(net70),
    .B(_01242_));
 sg13g2_a21oi_1 _06460_ (.A1(_00119_),
    .A2(net75),
    .Y(_01244_),
    .B1(net353));
 sg13g2_nand2_1 _06461_ (.Y(_01245_),
    .A(_01243_),
    .B(_01244_));
 sg13g2_inv_1 _06462_ (.Y(_01246_),
    .A(_00120_));
 sg13g2_buf_1 _06463_ (.A(net352),
    .X(_01247_));
 sg13g2_nand2_1 _06464_ (.Y(_01248_),
    .A(_00855_),
    .B(_00858_));
 sg13g2_inv_1 _06465_ (.Y(_01249_),
    .A(_01248_));
 sg13g2_nand2_2 _06466_ (.Y(_01250_),
    .A(_01070_),
    .B(_01249_));
 sg13g2_nand2_1 _06467_ (.Y(_01251_),
    .A(_00119_),
    .B(_01250_));
 sg13g2_a221oi_1 _06468_ (.B2(_01251_),
    .C1(net45),
    .B1(net257),
    .A1(net404),
    .Y(_01252_),
    .A2(_01246_));
 sg13g2_buf_1 _06469_ (.A(_00917_),
    .X(_01253_));
 sg13g2_nand3_1 _06470_ (.B(_00977_),
    .C(_01189_),
    .A(net450),
    .Y(_01254_));
 sg13g2_buf_1 _06471_ (.A(_01254_),
    .X(_01255_));
 sg13g2_nand2_1 _06472_ (.Y(_01256_),
    .A(net447),
    .B(_01255_));
 sg13g2_a221oi_1 _06473_ (.B2(_01252_),
    .C1(_01256_),
    .B1(_01245_),
    .A1(_00119_),
    .Y(_01257_),
    .A2(net39));
 sg13g2_a21o_1 _06474_ (.A2(_01239_),
    .A1(net453),
    .B1(_01257_),
    .X(_00006_));
 sg13g2_nand2b_1 _06475_ (.Y(_01258_),
    .B(_01250_),
    .A_N(_00121_));
 sg13g2_a221oi_1 _06476_ (.B2(_01258_),
    .C1(net50),
    .B1(_01073_),
    .A1(net448),
    .Y(_01259_),
    .A2(_00122_));
 sg13g2_and2_1 _06477_ (.A(net260),
    .B(net32),
    .X(_01260_));
 sg13g2_and2_1 _06478_ (.A(_00611_),
    .B(_01260_),
    .X(_01261_));
 sg13g2_a21o_1 _06479_ (.A2(_00911_),
    .A1(net93),
    .B1(_01261_),
    .X(_01262_));
 sg13g2_buf_1 _06480_ (.A(_01262_),
    .X(_01263_));
 sg13g2_a21o_1 _06481_ (.A2(_01263_),
    .A1(net70),
    .B1(net258),
    .X(_01264_));
 sg13g2_a21oi_1 _06482_ (.A1(net75),
    .A2(_01259_),
    .Y(_01265_),
    .B1(net45));
 sg13g2_nor2_1 _06483_ (.A(_00121_),
    .B(_01265_),
    .Y(_01266_));
 sg13g2_a21oi_1 _06484_ (.A1(_01259_),
    .A2(_01264_),
    .Y(_01267_),
    .B1(_01266_));
 sg13g2_nand2_1 _06485_ (.Y(_01268_),
    .A(net451),
    .B(_01239_));
 sg13g2_o21ai_1 _06486_ (.B1(_01268_),
    .Y(_00007_),
    .A1(_01256_),
    .A2(_01267_));
 sg13g2_nand2b_1 _06487_ (.Y(_01269_),
    .B(_01250_),
    .A_N(_00123_));
 sg13g2_a221oi_1 _06488_ (.B2(_01269_),
    .C1(net50),
    .B1(_01073_),
    .A1(net448),
    .Y(_01270_),
    .A2(_00124_));
 sg13g2_nor3_1 _06489_ (.A(net160),
    .B(_00789_),
    .C(_00934_),
    .Y(_01271_));
 sg13g2_nor3_1 _06490_ (.A(net160),
    .B(_00789_),
    .C(_00954_),
    .Y(_01272_));
 sg13g2_mux2_1 _06491_ (.A0(_01271_),
    .A1(_01272_),
    .S(_00928_),
    .X(_01273_));
 sg13g2_mux2_1 _06492_ (.A0(_00939_),
    .A1(_00940_),
    .S(net160),
    .X(_01274_));
 sg13g2_nor2_2 _06493_ (.A(_01273_),
    .B(_01274_),
    .Y(_01275_));
 sg13g2_a21o_1 _06494_ (.A2(_01275_),
    .A1(net70),
    .B1(net258),
    .X(_01276_));
 sg13g2_a21oi_1 _06495_ (.A1(net75),
    .A2(_01270_),
    .Y(_01277_),
    .B1(net45));
 sg13g2_nor2_1 _06496_ (.A(_00123_),
    .B(_01277_),
    .Y(_01278_));
 sg13g2_a21oi_1 _06497_ (.A1(_01270_),
    .A2(_01276_),
    .Y(_01279_),
    .B1(_01278_));
 sg13g2_nand2_1 _06498_ (.Y(_01280_),
    .A(net477),
    .B(_01239_));
 sg13g2_o21ai_1 _06499_ (.B1(_01280_),
    .Y(_00008_),
    .A1(_01256_),
    .A2(_01279_));
 sg13g2_nor2_1 _06500_ (.A(net160),
    .B(_00953_),
    .Y(_01281_));
 sg13g2_a22oi_1 _06501_ (.Y(_01282_),
    .B1(_00958_),
    .B2(_01281_),
    .A2(_00837_),
    .A1(_00735_));
 sg13g2_buf_1 _06502_ (.A(_01282_),
    .X(_01283_));
 sg13g2_and2_1 _06503_ (.A(_00125_),
    .B(net75),
    .X(_01284_));
 sg13g2_a21oi_1 _06504_ (.A1(net70),
    .A2(_01283_),
    .Y(_01285_),
    .B1(_01284_));
 sg13g2_buf_1 _06505_ (.A(net404),
    .X(_01286_));
 sg13g2_buf_1 _06506_ (.A(net257),
    .X(_01287_));
 sg13g2_nand2b_1 _06507_ (.Y(_01288_),
    .B(_01250_),
    .A_N(_00125_));
 sg13g2_nand3_1 _06508_ (.B(net53),
    .C(_01255_),
    .A(net447),
    .Y(_01289_));
 sg13g2_a221oi_1 _06509_ (.B2(_01288_),
    .C1(_01289_),
    .B1(net157),
    .A1(net349),
    .Y(_01290_),
    .A2(_00126_));
 sg13g2_o21ai_1 _06510_ (.B1(_01290_),
    .Y(_01291_),
    .A1(net258),
    .A2(_01285_));
 sg13g2_nand2_2 _06511_ (.Y(_01292_),
    .A(net478),
    .B(_00846_));
 sg13g2_o21ai_1 _06512_ (.B1(_01255_),
    .Y(_01293_),
    .A1(_00125_),
    .A2(_01292_));
 sg13g2_o21ai_1 _06513_ (.B1(_01293_),
    .Y(_01294_),
    .A1(net476),
    .A2(_01255_));
 sg13g2_nand2_1 _06514_ (.Y(_00009_),
    .A(_01291_),
    .B(_01294_));
 sg13g2_nor2b_1 _06515_ (.A(_05094_),
    .B_N(_05093_),
    .Y(_01295_));
 sg13g2_buf_1 _06516_ (.A(_01295_),
    .X(_01296_));
 sg13g2_nand2_1 _06517_ (.Y(_01297_),
    .A(_00972_),
    .B(_01296_));
 sg13g2_buf_1 _06518_ (.A(net404),
    .X(_01298_));
 sg13g2_nand2b_1 _06519_ (.Y(_01299_),
    .B(net262),
    .A_N(net161));
 sg13g2_buf_2 _06520_ (.A(_01299_),
    .X(_01300_));
 sg13g2_nand2_1 _06521_ (.Y(_01301_),
    .A(_05139_),
    .B(net161));
 sg13g2_buf_2 _06522_ (.A(_00097_),
    .X(_01302_));
 sg13g2_a21oi_1 _06523_ (.A1(_01300_),
    .A2(_01301_),
    .Y(_01303_),
    .B1(_01302_));
 sg13g2_buf_1 _06524_ (.A(_01303_),
    .X(_01304_));
 sg13g2_nor2_1 _06525_ (.A(_05139_),
    .B(net161),
    .Y(_01305_));
 sg13g2_buf_1 _06526_ (.A(_01305_),
    .X(_01306_));
 sg13g2_o21ai_1 _06527_ (.B1(net351),
    .Y(_01307_),
    .A1(_00104_),
    .A2(_01306_));
 sg13g2_a21oi_1 _06528_ (.A1(_00840_),
    .A2(net47),
    .Y(_01308_),
    .B1(_01307_));
 sg13g2_a21oi_1 _06529_ (.A1(net348),
    .A2(_00103_),
    .Y(_01309_),
    .B1(_01308_));
 sg13g2_inv_1 _06530_ (.Y(_01310_),
    .A(_00889_));
 sg13g2_nand3_1 _06531_ (.B(_00886_),
    .C(_01310_),
    .A(_00853_),
    .Y(_01311_));
 sg13g2_buf_1 _06532_ (.A(_01311_),
    .X(_01312_));
 sg13g2_nor2_2 _06533_ (.A(_00861_),
    .B(_01312_),
    .Y(_01313_));
 sg13g2_o21ai_1 _06534_ (.B1(net53),
    .Y(_01314_),
    .A1(net350),
    .A2(_01313_));
 sg13g2_o21ai_1 _06535_ (.B1(net478),
    .Y(_01315_),
    .A1(_01238_),
    .A2(_01297_));
 sg13g2_buf_1 _06536_ (.A(_01315_),
    .X(_01316_));
 sg13g2_a21oi_1 _06537_ (.A1(_00104_),
    .A2(_01314_),
    .Y(_01317_),
    .B1(_01316_));
 sg13g2_o21ai_1 _06538_ (.B1(_01317_),
    .Y(_01318_),
    .A1(net40),
    .A2(_01309_));
 sg13g2_o21ai_1 _06539_ (.B1(_01318_),
    .Y(_00010_),
    .A1(_00979_),
    .A2(_01297_));
 sg13g2_nand2_2 _06540_ (.Y(_01319_),
    .A(_01079_),
    .B(_01152_));
 sg13g2_or2_1 _06541_ (.X(_01320_),
    .B(_01313_),
    .A(_00106_));
 sg13g2_a22oi_1 _06542_ (.Y(_01321_),
    .B1(_01319_),
    .B2(_01320_),
    .A2(_00105_),
    .A1(net449));
 sg13g2_a21o_1 _06543_ (.A2(_01301_),
    .A1(_01300_),
    .B1(_01302_),
    .X(_01322_));
 sg13g2_buf_2 _06544_ (.A(_01322_),
    .X(_01323_));
 sg13g2_buf_1 _06545_ (.A(net351),
    .X(_01324_));
 sg13g2_o21ai_1 _06546_ (.B1(net256),
    .Y(_01325_),
    .A1(_00913_),
    .A2(_01323_));
 sg13g2_a21oi_1 _06547_ (.A1(_01300_),
    .A2(_01321_),
    .Y(_01326_),
    .B1(net45));
 sg13g2_nor2_1 _06548_ (.A(_00106_),
    .B(_01326_),
    .Y(_01327_));
 sg13g2_a21oi_1 _06549_ (.A1(_01321_),
    .A2(_01325_),
    .Y(_01328_),
    .B1(_01327_));
 sg13g2_and2_1 _06550_ (.A(_00972_),
    .B(_01296_),
    .X(_01329_));
 sg13g2_buf_2 _06551_ (.A(_01329_),
    .X(_01330_));
 sg13g2_nand3_1 _06552_ (.B(net92),
    .C(_01330_),
    .A(net451),
    .Y(_01331_));
 sg13g2_o21ai_1 _06553_ (.B1(_01331_),
    .Y(_00011_),
    .A1(_01316_),
    .A2(_01328_));
 sg13g2_nor2_1 _06554_ (.A(net46),
    .B(_01316_),
    .Y(_01332_));
 sg13g2_o21ai_1 _06555_ (.B1(net157),
    .Y(_01333_),
    .A1(_00108_),
    .A2(_01313_));
 sg13g2_nand2_1 _06556_ (.Y(_01334_),
    .A(net348),
    .B(_00107_));
 sg13g2_nand3_1 _06557_ (.B(_01333_),
    .C(_01334_),
    .A(_01332_),
    .Y(_01335_));
 sg13g2_inv_1 _06558_ (.Y(_01336_),
    .A(_00108_));
 sg13g2_a221oi_1 _06559_ (.B2(net47),
    .C1(net258),
    .B1(_00942_),
    .A1(_01336_),
    .Y(_01337_),
    .A2(_01300_));
 sg13g2_inv_1 _06560_ (.Y(_01338_),
    .A(net477));
 sg13g2_nor2_1 _06561_ (.A(_01338_),
    .B(_01238_),
    .Y(_01339_));
 sg13g2_nor2_1 _06562_ (.A(net48),
    .B(_01316_),
    .Y(_01340_));
 sg13g2_a22oi_1 _06563_ (.Y(_01341_),
    .B1(_01340_),
    .B2(_01336_),
    .A2(_01330_),
    .A1(_01339_));
 sg13g2_o21ai_1 _06564_ (.B1(_01341_),
    .Y(_00012_),
    .A1(_01335_),
    .A2(_01337_));
 sg13g2_o21ai_1 _06565_ (.B1(net157),
    .Y(_01342_),
    .A1(_00110_),
    .A2(_01313_));
 sg13g2_nand2_1 _06566_ (.Y(_01343_),
    .A(net348),
    .B(_00109_));
 sg13g2_nand3_1 _06567_ (.B(_01342_),
    .C(_01343_),
    .A(_01332_),
    .Y(_01344_));
 sg13g2_inv_1 _06568_ (.Y(_01345_),
    .A(_00110_));
 sg13g2_a221oi_1 _06569_ (.B2(net47),
    .C1(net258),
    .B1(_00962_),
    .A1(_01345_),
    .Y(_01346_),
    .A2(_01300_));
 sg13g2_a22oi_1 _06570_ (.Y(_01347_),
    .B1(_01340_),
    .B2(_01345_),
    .A2(_01330_),
    .A1(_01185_));
 sg13g2_o21ai_1 _06571_ (.B1(_01347_),
    .Y(_00013_),
    .A1(_01344_),
    .A2(_01346_));
 sg13g2_o21ai_1 _06572_ (.B1(net351),
    .Y(_01348_),
    .A1(_00127_),
    .A2(net68));
 sg13g2_inv_1 _06573_ (.Y(_01349_),
    .A(_01348_));
 sg13g2_o21ai_1 _06574_ (.B1(_01349_),
    .Y(_01350_),
    .A1(_01067_),
    .A2(_01323_));
 sg13g2_or2_1 _06575_ (.X(_01351_),
    .B(_01312_),
    .A(_01068_));
 sg13g2_nand3_1 _06576_ (.B(_01247_),
    .C(_01351_),
    .A(_00127_),
    .Y(_01352_));
 sg13g2_a21oi_1 _06577_ (.A1(_01350_),
    .A2(_01352_),
    .Y(_01353_),
    .B1(net39));
 sg13g2_nand3_1 _06578_ (.B(net92),
    .C(_01296_),
    .A(net450),
    .Y(_01354_));
 sg13g2_nand2b_1 _06579_ (.Y(_01355_),
    .B(_01079_),
    .A_N(net448));
 sg13g2_buf_2 _06580_ (.A(_01355_),
    .X(_01356_));
 sg13g2_a21oi_1 _06581_ (.A1(_00127_),
    .A2(_01356_),
    .Y(_01357_),
    .B1(net457));
 sg13g2_nand2_1 _06582_ (.Y(_01358_),
    .A(_01354_),
    .B(_01357_));
 sg13g2_and3_1 _06583_ (.X(_01359_),
    .A(net450),
    .B(_00977_),
    .C(_01296_));
 sg13g2_buf_1 _06584_ (.A(_01359_),
    .X(_01360_));
 sg13g2_nand2_1 _06585_ (.Y(_01361_),
    .A(net453),
    .B(_01360_));
 sg13g2_o21ai_1 _06586_ (.B1(_01361_),
    .Y(_00015_),
    .A1(_01353_),
    .A2(_01358_));
 sg13g2_nor2_1 _06587_ (.A(_01068_),
    .B(_01312_),
    .Y(_01362_));
 sg13g2_nand2b_1 _06588_ (.Y(_01363_),
    .B(_01114_),
    .A_N(_01302_));
 sg13g2_nor2_1 _06589_ (.A(_01300_),
    .B(net353),
    .Y(_01364_));
 sg13g2_a22oi_1 _06590_ (.Y(_01365_),
    .B1(_01363_),
    .B2(_01364_),
    .A2(_01362_),
    .A1(net257));
 sg13g2_nor2_1 _06591_ (.A(net39),
    .B(_01365_),
    .Y(_01366_));
 sg13g2_buf_1 _06592_ (.A(_01253_),
    .X(_01367_));
 sg13g2_a21oi_1 _06593_ (.A1(net94),
    .A2(_01101_),
    .Y(_01368_),
    .B1(_01112_));
 sg13g2_nand3_1 _06594_ (.B(net256),
    .C(net47),
    .A(net53),
    .Y(_01369_));
 sg13g2_o21ai_1 _06595_ (.B1(_00128_),
    .Y(_01370_),
    .A1(_01368_),
    .A2(_01369_));
 sg13g2_nand3_1 _06596_ (.B(_01354_),
    .C(_01370_),
    .A(net403),
    .Y(_01371_));
 sg13g2_nand2_1 _06597_ (.Y(_01372_),
    .A(net451),
    .B(_01360_));
 sg13g2_o21ai_1 _06598_ (.B1(_01372_),
    .Y(_00016_),
    .A1(_01366_),
    .A2(_01371_));
 sg13g2_nor2_1 _06599_ (.A(_01149_),
    .B(_01323_),
    .Y(_01373_));
 sg13g2_o21ai_1 _06600_ (.B1(_01324_),
    .Y(_01374_),
    .A1(_00129_),
    .A2(net68));
 sg13g2_o21ai_1 _06601_ (.B1(net257),
    .Y(_01375_),
    .A1(_00129_),
    .A2(_01362_));
 sg13g2_o21ai_1 _06602_ (.B1(_01375_),
    .Y(_01376_),
    .A1(_01373_),
    .A2(_01374_));
 sg13g2_nor2_1 _06603_ (.A(net39),
    .B(_01360_),
    .Y(_01377_));
 sg13g2_a21oi_1 _06604_ (.A1(_00129_),
    .A2(_01356_),
    .Y(_01378_),
    .B1(net457));
 sg13g2_nor2_1 _06605_ (.A(_01360_),
    .B(_01378_),
    .Y(_01379_));
 sg13g2_a221oi_1 _06606_ (.B2(_01377_),
    .C1(_01379_),
    .B1(_01376_),
    .A1(_01338_),
    .Y(_00017_),
    .A2(_01360_));
 sg13g2_and2_1 _06607_ (.A(net412),
    .B(net47),
    .X(_01380_));
 sg13g2_nand2_1 _06608_ (.Y(_01381_),
    .A(net456),
    .B(_01305_));
 sg13g2_o21ai_1 _06609_ (.B1(_01381_),
    .Y(_01382_),
    .A1(net456),
    .A2(_01351_));
 sg13g2_a21oi_1 _06610_ (.A1(_01292_),
    .A2(_01382_),
    .Y(_01383_),
    .B1(_00130_));
 sg13g2_or2_1 _06611_ (.X(_01384_),
    .B(_01383_),
    .A(net406));
 sg13g2_a21oi_1 _06612_ (.A1(_01177_),
    .A2(_01380_),
    .Y(_01385_),
    .B1(_01384_));
 sg13g2_a21oi_1 _06613_ (.A1(_00130_),
    .A2(_01356_),
    .Y(_01386_),
    .B1(net457));
 sg13g2_nand2_1 _06614_ (.Y(_01387_),
    .A(_01354_),
    .B(_01386_));
 sg13g2_nand2_1 _06615_ (.Y(_01388_),
    .A(net476),
    .B(_01360_));
 sg13g2_o21ai_1 _06616_ (.B1(_01388_),
    .Y(_00018_),
    .A1(_01385_),
    .A2(_01387_));
 sg13g2_nand2_1 _06617_ (.Y(_01389_),
    .A(_00855_),
    .B(_00859_));
 sg13g2_nor2_1 _06618_ (.A(_01389_),
    .B(_01312_),
    .Y(_01390_));
 sg13g2_o21ai_1 _06619_ (.B1(_01118_),
    .Y(_01391_),
    .A1(net350),
    .A2(_01390_));
 sg13g2_nor2_1 _06620_ (.A(_01194_),
    .B(_01323_),
    .Y(_01392_));
 sg13g2_o21ai_1 _06621_ (.B1(net256),
    .Y(_01393_),
    .A1(_00131_),
    .A2(_01306_));
 sg13g2_nand2_1 _06622_ (.Y(_01394_),
    .A(_01181_),
    .B(_00132_));
 sg13g2_o21ai_1 _06623_ (.B1(_01394_),
    .Y(_01395_),
    .A1(_01392_),
    .A2(_01393_));
 sg13g2_nand2_1 _06624_ (.Y(_01396_),
    .A(_05093_),
    .B(_05094_));
 sg13g2_nor2_1 _06625_ (.A(_05095_),
    .B(_01396_),
    .Y(_01397_));
 sg13g2_buf_1 _06626_ (.A(_01397_),
    .X(_01398_));
 sg13g2_a21oi_2 _06627_ (.B1(net457),
    .Y(_01399_),
    .A2(net347),
    .A1(net92));
 sg13g2_inv_1 _06628_ (.Y(_01400_),
    .A(_01399_));
 sg13g2_a221oi_1 _06629_ (.B2(net49),
    .C1(_01400_),
    .B1(_01395_),
    .A1(_00131_),
    .Y(_01401_),
    .A2(_01391_));
 sg13g2_nand3_1 _06630_ (.B(net92),
    .C(net347),
    .A(net453),
    .Y(_01402_));
 sg13g2_nand2b_1 _06631_ (.Y(_00019_),
    .B(_01402_),
    .A_N(_01401_));
 sg13g2_nand2_1 _06632_ (.Y(_01403_),
    .A(net92),
    .B(net347));
 sg13g2_or2_1 _06633_ (.X(_01404_),
    .B(_01390_),
    .A(_00133_));
 sg13g2_a22oi_1 _06634_ (.Y(_01405_),
    .B1(net352),
    .B2(_01404_),
    .A2(_00134_),
    .A1(net448));
 sg13g2_a21oi_1 _06635_ (.A1(_01300_),
    .A2(_01405_),
    .Y(_01406_),
    .B1(net50));
 sg13g2_nor3_1 _06636_ (.A(net457),
    .B(_00133_),
    .C(_01406_),
    .Y(_01407_));
 sg13g2_o21ai_1 _06637_ (.B1(net256),
    .Y(_01408_),
    .A1(_01215_),
    .A2(_01323_));
 sg13g2_nand4_1 _06638_ (.B(net48),
    .C(_01405_),
    .A(net447),
    .Y(_01409_),
    .D(_01408_));
 sg13g2_nor2b_1 _06639_ (.A(_01407_),
    .B_N(_01409_),
    .Y(_01410_));
 sg13g2_nor2_1 _06640_ (.A(net451),
    .B(_01403_),
    .Y(_01411_));
 sg13g2_a21oi_1 _06641_ (.A1(_01403_),
    .A2(_01410_),
    .Y(_00020_),
    .B1(_01411_));
 sg13g2_or2_1 _06642_ (.X(_01412_),
    .B(_01390_),
    .A(_00135_));
 sg13g2_a22oi_1 _06643_ (.Y(_01413_),
    .B1(_01287_),
    .B2(_01412_),
    .A2(_00136_),
    .A1(_01298_));
 sg13g2_o21ai_1 _06644_ (.B1(_01324_),
    .Y(_01414_),
    .A1(_00135_),
    .A2(net68));
 sg13g2_inv_1 _06645_ (.Y(_01415_),
    .A(_01414_));
 sg13g2_o21ai_1 _06646_ (.B1(_01415_),
    .Y(_01416_),
    .A1(_01220_),
    .A2(_01323_));
 sg13g2_nand4_1 _06647_ (.B(_01399_),
    .C(_01413_),
    .A(net49),
    .Y(_01417_),
    .D(_01416_));
 sg13g2_nor2_1 _06648_ (.A(_00135_),
    .B(net49),
    .Y(_01418_));
 sg13g2_a22oi_1 _06649_ (.Y(_01419_),
    .B1(_01399_),
    .B2(_01418_),
    .A2(net347),
    .A1(_01339_));
 sg13g2_nand2_1 _06650_ (.Y(_00021_),
    .A(_01417_),
    .B(_01419_));
 sg13g2_buf_1 _06651_ (.A(_00137_),
    .X(_01420_));
 sg13g2_o21ai_1 _06652_ (.B1(_01247_),
    .Y(_01421_),
    .A1(_01420_),
    .A2(_01390_));
 sg13g2_a21oi_1 _06653_ (.A1(net349),
    .A2(_00138_),
    .Y(_01422_),
    .B1(_00981_));
 sg13g2_nand3_1 _06654_ (.B(_01421_),
    .C(_01422_),
    .A(_01399_),
    .Y(_01423_));
 sg13g2_buf_1 _06655_ (.A(net256),
    .X(_01424_));
 sg13g2_o21ai_1 _06656_ (.B1(net156),
    .Y(_01425_),
    .A1(_01420_),
    .A2(net68));
 sg13g2_a21oi_1 _06657_ (.A1(_01227_),
    .A2(_01304_),
    .Y(_01426_),
    .B1(_01425_));
 sg13g2_nor2_1 _06658_ (.A(_01420_),
    .B(net49),
    .Y(_01427_));
 sg13g2_a22oi_1 _06659_ (.Y(_01428_),
    .B1(_01399_),
    .B2(_01427_),
    .A2(net347),
    .A1(_01185_));
 sg13g2_o21ai_1 _06660_ (.B1(_01428_),
    .Y(_00022_),
    .A1(_01423_),
    .A2(_01426_));
 sg13g2_nand3_1 _06661_ (.B(_05094_),
    .C(net450),
    .A(_05093_),
    .Y(_01429_));
 sg13g2_buf_2 _06662_ (.A(_01429_),
    .X(_01430_));
 sg13g2_nand2b_1 _06663_ (.Y(_01431_),
    .B(net47),
    .A_N(_01242_));
 sg13g2_o21ai_1 _06664_ (.B1(net256),
    .Y(_01432_),
    .A1(_00139_),
    .A2(net68));
 sg13g2_inv_1 _06665_ (.Y(_01433_),
    .A(_01432_));
 sg13g2_a22oi_1 _06666_ (.Y(_01434_),
    .B1(_01431_),
    .B2(_01433_),
    .A2(_00140_),
    .A1(net348));
 sg13g2_nor2_1 _06667_ (.A(_01248_),
    .B(_01312_),
    .Y(_01435_));
 sg13g2_o21ai_1 _06668_ (.B1(net53),
    .Y(_01436_),
    .A1(net350),
    .A2(_01435_));
 sg13g2_o21ai_1 _06669_ (.B1(net478),
    .Y(_01437_),
    .A1(_01238_),
    .A2(_01430_));
 sg13g2_buf_1 _06670_ (.A(_01437_),
    .X(_01438_));
 sg13g2_a21oi_1 _06671_ (.A1(_00139_),
    .A2(_01436_),
    .Y(_01439_),
    .B1(_01438_));
 sg13g2_o21ai_1 _06672_ (.B1(_01439_),
    .Y(_01440_),
    .A1(net40),
    .A2(_01434_));
 sg13g2_o21ai_1 _06673_ (.B1(_01440_),
    .Y(_00023_),
    .A1(_00979_),
    .A2(_01430_));
 sg13g2_buf_1 _06674_ (.A(_00141_),
    .X(_01441_));
 sg13g2_o21ai_1 _06675_ (.B1(net156),
    .Y(_01442_),
    .A1(_01441_),
    .A2(net68));
 sg13g2_a21oi_1 _06676_ (.A1(_01263_),
    .A2(net47),
    .Y(_01443_),
    .B1(_01442_));
 sg13g2_a21oi_1 _06677_ (.A1(net349),
    .A2(_00142_),
    .Y(_01444_),
    .B1(net46));
 sg13g2_o21ai_1 _06678_ (.B1(net157),
    .Y(_01445_),
    .A1(_01441_),
    .A2(_01435_));
 sg13g2_nand3b_1 _06679_ (.B(_01444_),
    .C(_01445_),
    .Y(_01446_),
    .A_N(_01438_));
 sg13g2_nor2_1 _06680_ (.A(_01238_),
    .B(_01430_),
    .Y(_01447_));
 sg13g2_nor3_1 _06681_ (.A(_01441_),
    .B(net48),
    .C(_01438_),
    .Y(_01448_));
 sg13g2_a21oi_1 _06682_ (.A1(_00921_),
    .A2(_01447_),
    .Y(_01449_),
    .B1(_01448_));
 sg13g2_o21ai_1 _06683_ (.B1(_01449_),
    .Y(_00024_),
    .A1(_01443_),
    .A2(_01446_));
 sg13g2_or2_1 _06684_ (.X(_01450_),
    .B(_01435_),
    .A(_00143_));
 sg13g2_o21ai_1 _06685_ (.B1(net351),
    .Y(_01451_),
    .A1(_00143_),
    .A2(net68));
 sg13g2_a21oi_1 _06686_ (.A1(_01275_),
    .A2(net47),
    .Y(_01452_),
    .B1(_01451_));
 sg13g2_a221oi_1 _06687_ (.B2(_01450_),
    .C1(_01452_),
    .B1(net257),
    .A1(net404),
    .Y(_01453_),
    .A2(_00144_));
 sg13g2_nor2_1 _06688_ (.A(_00143_),
    .B(net48),
    .Y(_01454_));
 sg13g2_a21oi_1 _06689_ (.A1(net49),
    .A2(_01453_),
    .Y(_01455_),
    .B1(_01454_));
 sg13g2_nor2_1 _06690_ (.A(_00972_),
    .B(_01396_),
    .Y(_01456_));
 sg13g2_nand2_1 _06691_ (.Y(_01457_),
    .A(_01339_),
    .B(_01456_));
 sg13g2_o21ai_1 _06692_ (.B1(_01457_),
    .Y(_00026_),
    .A1(_01438_),
    .A2(_01455_));
 sg13g2_nor2_1 _06693_ (.A(_01283_),
    .B(_01323_),
    .Y(_01458_));
 sg13g2_o21ai_1 _06694_ (.B1(net156),
    .Y(_01459_),
    .A1(_00145_),
    .A2(net68));
 sg13g2_buf_1 _06695_ (.A(_00146_),
    .X(_01460_));
 sg13g2_or2_1 _06696_ (.X(_01461_),
    .B(_01435_),
    .A(_00145_));
 sg13g2_a221oi_1 _06697_ (.B2(_01461_),
    .C1(_01438_),
    .B1(_01319_),
    .A1(_01286_),
    .Y(_01462_),
    .A2(_01460_));
 sg13g2_o21ai_1 _06698_ (.B1(_01462_),
    .Y(_01463_),
    .A1(_01458_),
    .A2(_01459_));
 sg13g2_nor3_1 _06699_ (.A(_00145_),
    .B(net48),
    .C(_01438_),
    .Y(_01464_));
 sg13g2_a21oi_1 _06700_ (.A1(_01185_),
    .A2(_01456_),
    .Y(_01465_),
    .B1(_01464_));
 sg13g2_nand2_1 _06701_ (.Y(_00027_),
    .A(_01463_),
    .B(_01465_));
 sg13g2_nand3_1 _06702_ (.B(_05096_),
    .C(_00978_),
    .A(_05091_),
    .Y(_01466_));
 sg13g2_buf_1 _06703_ (.A(_01466_),
    .X(_01467_));
 sg13g2_nand2_1 _06704_ (.Y(_01468_),
    .A(_00112_),
    .B(_00981_));
 sg13g2_nand3_1 _06705_ (.B(_00111_),
    .C(_01118_),
    .A(_00984_),
    .Y(_01469_));
 sg13g2_nand4_1 _06706_ (.B(_01467_),
    .C(_01468_),
    .A(net403),
    .Y(_01470_),
    .D(_01469_));
 sg13g2_buf_1 _06707_ (.A(_01301_),
    .X(_01471_));
 sg13g2_nand2_1 _06708_ (.Y(_01472_),
    .A(_00112_),
    .B(_01471_));
 sg13g2_o21ai_1 _06709_ (.B1(_01472_),
    .Y(_01473_),
    .A1(_01471_),
    .A2(_00840_));
 sg13g2_inv_1 _06710_ (.Y(_01474_),
    .A(_00112_));
 sg13g2_nand2_1 _06711_ (.Y(_01475_),
    .A(_00863_),
    .B(_01310_));
 sg13g2_nor3_2 _06712_ (.A(_00853_),
    .B(_00861_),
    .C(_01475_),
    .Y(_01476_));
 sg13g2_nor3_1 _06713_ (.A(net412),
    .B(_01474_),
    .C(_01476_),
    .Y(_01477_));
 sg13g2_a21oi_1 _06714_ (.A1(_05102_),
    .A2(_01473_),
    .Y(_01478_),
    .B1(_01477_));
 sg13g2_nor2_1 _06715_ (.A(_01356_),
    .B(_01478_),
    .Y(_01479_));
 sg13g2_nand4_1 _06716_ (.B(_00895_),
    .C(_05096_),
    .A(_05091_),
    .Y(_01480_),
    .D(net92));
 sg13g2_o21ai_1 _06717_ (.B1(_01480_),
    .Y(_00028_),
    .A1(_01470_),
    .A2(_01479_));
 sg13g2_nand2_1 _06718_ (.Y(_01481_),
    .A(net449),
    .B(_00113_));
 sg13g2_o21ai_1 _06719_ (.B1(net352),
    .Y(_01482_),
    .A1(_00114_),
    .A2(_01476_));
 sg13g2_nor2_2 _06720_ (.A(_01301_),
    .B(_00987_),
    .Y(_01483_));
 sg13g2_nand2_1 _06721_ (.Y(_01484_),
    .A(_00913_),
    .B(_01483_));
 sg13g2_nand3_1 _06722_ (.B(_01482_),
    .C(_01484_),
    .A(_01481_),
    .Y(_01485_));
 sg13g2_nor2b_1 _06723_ (.A(net262),
    .B_N(net161),
    .Y(_01486_));
 sg13g2_buf_2 _06724_ (.A(_01486_),
    .X(_01487_));
 sg13g2_o21ai_1 _06725_ (.B1(_01079_),
    .Y(_01488_),
    .A1(_01487_),
    .A2(_00986_));
 sg13g2_buf_2 _06726_ (.A(_01488_),
    .X(_01489_));
 sg13g2_a221oi_1 _06727_ (.B2(_00114_),
    .C1(net405),
    .B1(_01489_),
    .A1(_01186_),
    .Y(_01490_),
    .A2(_01485_));
 sg13g2_mux2_1 _06728_ (.A0(_00922_),
    .A1(_01490_),
    .S(_01467_),
    .X(_00029_));
 sg13g2_nand2_1 _06729_ (.Y(_01491_),
    .A(_01487_),
    .B(_01089_));
 sg13g2_nor2_1 _06730_ (.A(_00116_),
    .B(_01476_),
    .Y(_01492_));
 sg13g2_nor3_1 _06731_ (.A(net449),
    .B(net456),
    .C(_01492_),
    .Y(_01493_));
 sg13g2_a21oi_1 _06732_ (.A1(net449),
    .A2(_00115_),
    .Y(_01494_),
    .B1(_01493_));
 sg13g2_o21ai_1 _06733_ (.B1(_01494_),
    .Y(_01495_),
    .A1(_00942_),
    .A2(_01491_));
 sg13g2_a221oi_1 _06734_ (.B2(_01119_),
    .C1(net405),
    .B1(_01495_),
    .A1(_00116_),
    .Y(_01496_),
    .A2(_01489_));
 sg13g2_mux2_1 _06735_ (.A0(net477),
    .A1(_01496_),
    .S(_01467_),
    .X(_00030_));
 sg13g2_nor2_1 _06736_ (.A(_00118_),
    .B(_01476_),
    .Y(_01497_));
 sg13g2_nor3_1 _06737_ (.A(_00983_),
    .B(net456),
    .C(_01497_),
    .Y(_01498_));
 sg13g2_a21oi_1 _06738_ (.A1(_00983_),
    .A2(_00117_),
    .Y(_01499_),
    .B1(_01498_));
 sg13g2_o21ai_1 _06739_ (.B1(_01499_),
    .Y(_01500_),
    .A1(_00962_),
    .A2(_01491_));
 sg13g2_a221oi_1 _06740_ (.B2(_01119_),
    .C1(net405),
    .B1(_01500_),
    .A1(_00118_),
    .Y(_01501_),
    .A2(_01489_));
 sg13g2_mux2_1 _06741_ (.A0(net476),
    .A1(_01501_),
    .S(_01467_),
    .X(_00031_));
 sg13g2_nand4_1 _06742_ (.B(_05095_),
    .C(_00099_),
    .A(_05092_),
    .Y(_01502_),
    .D(_00969_));
 sg13g2_a21oi_1 _06743_ (.A1(_00974_),
    .A2(_01502_),
    .Y(_01503_),
    .B1(_00971_));
 sg13g2_buf_1 _06744_ (.A(_01503_),
    .X(_01504_));
 sg13g2_nand3_1 _06745_ (.B(_01083_),
    .C(net255),
    .A(net453),
    .Y(_01505_));
 sg13g2_inv_1 _06746_ (.Y(_01506_),
    .A(_00132_));
 sg13g2_inv_1 _06747_ (.Y(_01507_),
    .A(_01475_));
 sg13g2_nand3_1 _06748_ (.B(_00861_),
    .C(_01507_),
    .A(_00885_),
    .Y(_01508_));
 sg13g2_buf_1 _06749_ (.A(_01508_),
    .X(_01509_));
 sg13g2_nor2_1 _06750_ (.A(_01068_),
    .B(_01509_),
    .Y(_01510_));
 sg13g2_nor3_1 _06751_ (.A(_01506_),
    .B(net350),
    .C(_01510_),
    .Y(_01511_));
 sg13g2_a221oi_1 _06752_ (.B2(_01483_),
    .C1(_01511_),
    .B1(_01067_),
    .A1(net406),
    .Y(_01512_),
    .A2(_00131_));
 sg13g2_inv_2 _06753_ (.Y(_01513_),
    .A(_01503_));
 sg13g2_o21ai_1 _06754_ (.B1(_05057_),
    .Y(_01514_),
    .A1(_00970_),
    .A2(_01513_));
 sg13g2_buf_1 _06755_ (.A(_01514_),
    .X(_01515_));
 sg13g2_a21oi_1 _06756_ (.A1(_00132_),
    .A2(_01489_),
    .Y(_01516_),
    .B1(_01515_));
 sg13g2_o21ai_1 _06757_ (.B1(_01516_),
    .Y(_01517_),
    .A1(_00982_),
    .A2(_01512_));
 sg13g2_nand2_1 _06758_ (.Y(_00032_),
    .A(_01505_),
    .B(_01517_));
 sg13g2_a21o_1 _06759_ (.A2(_01489_),
    .A1(_00134_),
    .B1(_01515_),
    .X(_01518_));
 sg13g2_nor2b_1 _06760_ (.A(_00133_),
    .B_N(_00984_),
    .Y(_01519_));
 sg13g2_or3_1 _06761_ (.A(net412),
    .B(_00134_),
    .C(_01510_),
    .X(_01520_));
 sg13g2_o21ai_1 _06762_ (.B1(net412),
    .Y(_01521_),
    .A1(net67),
    .A2(_01114_));
 sg13g2_a21oi_1 _06763_ (.A1(_01520_),
    .A2(_01521_),
    .Y(_01522_),
    .B1(net348));
 sg13g2_nor3_1 _06764_ (.A(_01240_),
    .B(_01519_),
    .C(_01522_),
    .Y(_01523_));
 sg13g2_and2_1 _06765_ (.A(_00921_),
    .B(net255),
    .X(_01524_));
 sg13g2_buf_1 _06766_ (.A(_01524_),
    .X(_01525_));
 sg13g2_nand2_1 _06767_ (.Y(_01526_),
    .A(_01083_),
    .B(_01525_));
 sg13g2_o21ai_1 _06768_ (.B1(_01526_),
    .Y(_00033_),
    .A1(_01518_),
    .A2(_01523_));
 sg13g2_nand2_1 _06769_ (.Y(_01527_),
    .A(_00946_),
    .B(net255));
 sg13g2_o21ai_1 _06770_ (.B1(net352),
    .Y(_01528_),
    .A1(_00136_),
    .A2(_01510_));
 sg13g2_inv_1 _06771_ (.Y(_01529_),
    .A(_01528_));
 sg13g2_a221oi_1 _06772_ (.B2(_01483_),
    .C1(_01529_),
    .B1(_01149_),
    .A1(net406),
    .Y(_01530_),
    .A2(_00135_));
 sg13g2_a21oi_1 _06773_ (.A1(_00136_),
    .A2(_01489_),
    .Y(_01531_),
    .B1(_01515_));
 sg13g2_o21ai_1 _06774_ (.B1(_01531_),
    .Y(_01532_),
    .A1(_00982_),
    .A2(_01530_));
 sg13g2_o21ai_1 _06775_ (.B1(_01532_),
    .Y(_00034_),
    .A1(_00970_),
    .A2(_01527_));
 sg13g2_a21o_1 _06776_ (.A2(_01489_),
    .A1(_00138_),
    .B1(_01515_),
    .X(_01533_));
 sg13g2_or2_1 _06777_ (.X(_01534_),
    .B(_01510_),
    .A(_00138_));
 sg13g2_a22oi_1 _06778_ (.Y(_01535_),
    .B1(_01287_),
    .B2(_01534_),
    .A2(_01420_),
    .A1(_01286_));
 sg13g2_o21ai_1 _06779_ (.B1(_01535_),
    .Y(_01536_),
    .A1(_01177_),
    .A2(_01491_));
 sg13g2_and2_1 _06780_ (.A(net476),
    .B(_01504_),
    .X(_01537_));
 sg13g2_buf_1 _06781_ (.A(_01537_),
    .X(_01538_));
 sg13g2_nor2_1 _06782_ (.A(net48),
    .B(_01533_),
    .Y(_01539_));
 sg13g2_a21oi_1 _06783_ (.A1(_01083_),
    .A2(_01538_),
    .Y(_01540_),
    .B1(_01539_));
 sg13g2_o21ai_1 _06784_ (.B1(_01540_),
    .Y(_00035_),
    .A1(_01533_),
    .A2(_01536_));
 sg13g2_nand2_1 _06785_ (.Y(_01541_),
    .A(_01201_),
    .B(net255));
 sg13g2_nor2_1 _06786_ (.A(_01389_),
    .B(_01509_),
    .Y(_01542_));
 sg13g2_nor2_1 _06787_ (.A(_00843_),
    .B(_05078_),
    .Y(_01543_));
 sg13g2_o21ai_1 _06788_ (.B1(_01543_),
    .Y(_01544_),
    .A1(_01152_),
    .A2(_01542_));
 sg13g2_nand2_1 _06789_ (.Y(_01545_),
    .A(net480),
    .B(_05057_));
 sg13g2_a21oi_1 _06790_ (.A1(_00147_),
    .A2(_01544_),
    .Y(_01546_),
    .B1(_01545_));
 sg13g2_o21ai_1 _06791_ (.B1(net156),
    .Y(_01547_),
    .A1(net67),
    .A2(_01194_));
 sg13g2_nand2_1 _06792_ (.Y(_01548_),
    .A(net67),
    .B(_01546_));
 sg13g2_a21oi_1 _06793_ (.A1(_01292_),
    .A2(_01548_),
    .Y(_01549_),
    .B1(_00147_));
 sg13g2_a21oi_1 _06794_ (.A1(_01546_),
    .A2(_01547_),
    .Y(_01550_),
    .B1(_01549_));
 sg13g2_nor2_1 _06795_ (.A(net453),
    .B(_01541_),
    .Y(_01551_));
 sg13g2_a21oi_1 _06796_ (.A1(_01541_),
    .A2(_01550_),
    .Y(_00037_),
    .B1(_01551_));
 sg13g2_nand2_1 _06797_ (.Y(_01552_),
    .A(net452),
    .B(_01541_));
 sg13g2_nand2_1 _06798_ (.Y(_01553_),
    .A(_01487_),
    .B(_00848_));
 sg13g2_inv_1 _06799_ (.Y(_01554_),
    .A(_00148_));
 sg13g2_nand2_1 _06800_ (.Y(_01555_),
    .A(_01554_),
    .B(net67));
 sg13g2_o21ai_1 _06801_ (.B1(_01555_),
    .Y(_01556_),
    .A1(_01215_),
    .A2(_01553_));
 sg13g2_o21ai_1 _06802_ (.B1(_00848_),
    .Y(_01557_),
    .A1(net412),
    .A2(_01542_));
 sg13g2_a22oi_1 _06803_ (.Y(_01558_),
    .B1(_01557_),
    .B2(_01554_),
    .A2(_01556_),
    .A1(net360));
 sg13g2_nand2_1 _06804_ (.Y(_01559_),
    .A(_01201_),
    .B(_01525_));
 sg13g2_o21ai_1 _06805_ (.B1(_01559_),
    .Y(_00038_),
    .A1(_01552_),
    .A2(_01558_));
 sg13g2_a21oi_1 _06806_ (.A1(net456),
    .A2(_01487_),
    .Y(_01560_),
    .B1(net449));
 sg13g2_and2_1 _06807_ (.A(_00149_),
    .B(_01560_),
    .X(_01561_));
 sg13g2_a221oi_1 _06808_ (.B2(net257),
    .C1(_01561_),
    .B1(_01542_),
    .A1(_01220_),
    .Y(_01562_),
    .A2(_01483_));
 sg13g2_a21oi_1 _06809_ (.A1(_00149_),
    .A2(_01356_),
    .Y(_01563_),
    .B1(_01552_));
 sg13g2_o21ai_1 _06810_ (.B1(_01563_),
    .Y(_01564_),
    .A1(net40),
    .A2(_01562_));
 sg13g2_o21ai_1 _06811_ (.B1(_01564_),
    .Y(_00039_),
    .A1(_01190_),
    .A2(_01527_));
 sg13g2_buf_1 _06812_ (.A(net447),
    .X(_01565_));
 sg13g2_or2_1 _06813_ (.X(_01566_),
    .B(_01487_),
    .A(_00150_));
 sg13g2_o21ai_1 _06814_ (.B1(_01566_),
    .Y(_01567_),
    .A1(_01226_),
    .A2(_01553_));
 sg13g2_nand4_1 _06815_ (.B(net360),
    .C(_01541_),
    .A(net402),
    .Y(_01568_),
    .D(_01567_));
 sg13g2_nor2_1 _06816_ (.A(_00150_),
    .B(_01552_),
    .Y(_01569_));
 sg13g2_a22oi_1 _06817_ (.Y(_01570_),
    .B1(_01557_),
    .B2(_01569_),
    .A2(_01538_),
    .A1(_01201_));
 sg13g2_nand2_1 _06818_ (.Y(_00040_),
    .A(_01568_),
    .B(_01570_));
 sg13g2_nand2_1 _06819_ (.Y(_01571_),
    .A(net450),
    .B(net255));
 sg13g2_o21ai_1 _06820_ (.B1(net452),
    .Y(_01572_),
    .A1(_01200_),
    .A2(_01571_));
 sg13g2_buf_1 _06821_ (.A(_01572_),
    .X(_01573_));
 sg13g2_nand3_1 _06822_ (.B(_00152_),
    .C(_01186_),
    .A(net349),
    .Y(_01574_));
 sg13g2_nand2_1 _06823_ (.Y(_01575_),
    .A(_00151_),
    .B(net46));
 sg13g2_nand3b_1 _06824_ (.B(_01574_),
    .C(_01575_),
    .Y(_01576_),
    .A_N(_01573_));
 sg13g2_mux2_1 _06825_ (.A0(_00151_),
    .A1(_01242_),
    .S(_01487_),
    .X(_01577_));
 sg13g2_inv_1 _06826_ (.Y(_01578_),
    .A(_00151_));
 sg13g2_nor2_1 _06827_ (.A(_01248_),
    .B(_01509_),
    .Y(_01579_));
 sg13g2_nor3_1 _06828_ (.A(net412),
    .B(_01578_),
    .C(_01579_),
    .Y(_01580_));
 sg13g2_a21oi_1 _06829_ (.A1(_05102_),
    .A2(_01577_),
    .Y(_01581_),
    .B1(_01580_));
 sg13g2_nor2_1 _06830_ (.A(_01356_),
    .B(_01581_),
    .Y(_01582_));
 sg13g2_nor2_1 _06831_ (.A(_01200_),
    .B(_01571_),
    .Y(_01583_));
 sg13g2_nand2_1 _06832_ (.Y(_01584_),
    .A(net453),
    .B(_01583_));
 sg13g2_o21ai_1 _06833_ (.B1(_01584_),
    .Y(_00041_),
    .A1(_01576_),
    .A2(_01582_));
 sg13g2_or2_1 _06834_ (.X(_01585_),
    .B(_01579_),
    .A(_00153_));
 sg13g2_a221oi_1 _06835_ (.B2(_01585_),
    .C1(_00980_),
    .B1(_01073_),
    .A1(_01180_),
    .Y(_01586_),
    .A2(_00154_));
 sg13g2_a21o_1 _06836_ (.A2(_01263_),
    .A1(_01487_),
    .B1(net353),
    .X(_01587_));
 sg13g2_a21oi_1 _06837_ (.A1(net67),
    .A2(_01586_),
    .Y(_01588_),
    .B1(net45));
 sg13g2_nor2_1 _06838_ (.A(_00153_),
    .B(_01588_),
    .Y(_01589_));
 sg13g2_a21oi_1 _06839_ (.A1(_01586_),
    .A2(_01587_),
    .Y(_01590_),
    .B1(_01589_));
 sg13g2_nand2_1 _06840_ (.Y(_01591_),
    .A(net451),
    .B(_01583_));
 sg13g2_o21ai_1 _06841_ (.B1(_01591_),
    .Y(_00042_),
    .A1(_01573_),
    .A2(_01590_));
 sg13g2_or2_1 _06842_ (.X(_01592_),
    .B(_01579_),
    .A(_00155_));
 sg13g2_a221oi_1 _06843_ (.B2(_01592_),
    .C1(_00980_),
    .B1(_01073_),
    .A1(net448),
    .Y(_01593_),
    .A2(_00156_));
 sg13g2_a21o_1 _06844_ (.A2(_01275_),
    .A1(_01487_),
    .B1(net353),
    .X(_01594_));
 sg13g2_a21oi_1 _06845_ (.A1(net67),
    .A2(_01593_),
    .Y(_01595_),
    .B1(_01233_));
 sg13g2_nor2_1 _06846_ (.A(_00155_),
    .B(_01595_),
    .Y(_01596_));
 sg13g2_a21oi_1 _06847_ (.A1(_01593_),
    .A2(_01594_),
    .Y(_01597_),
    .B1(_01596_));
 sg13g2_nand2_1 _06848_ (.Y(_01598_),
    .A(net477),
    .B(_01583_));
 sg13g2_o21ai_1 _06849_ (.B1(_01598_),
    .Y(_00043_),
    .A1(_01573_),
    .A2(_01597_));
 sg13g2_or2_1 _06850_ (.X(_01599_),
    .B(_01579_),
    .A(_00157_));
 sg13g2_a221oi_1 _06851_ (.B2(_01599_),
    .C1(_00846_),
    .B1(_01073_),
    .A1(_01180_),
    .Y(_01600_),
    .A2(_00158_));
 sg13g2_o21ai_1 _06852_ (.B1(net256),
    .Y(_01601_),
    .A1(net67),
    .A2(_01283_));
 sg13g2_a21oi_1 _06853_ (.A1(net67),
    .A2(_01600_),
    .Y(_01602_),
    .B1(_01233_));
 sg13g2_nor2_1 _06854_ (.A(_00157_),
    .B(_01602_),
    .Y(_01603_));
 sg13g2_a21oi_1 _06855_ (.A1(_01600_),
    .A2(_01601_),
    .Y(_01604_),
    .B1(_01603_));
 sg13g2_nand2_1 _06856_ (.Y(_01605_),
    .A(net476),
    .B(_01583_));
 sg13g2_o21ai_1 _06857_ (.B1(_01605_),
    .Y(_00044_),
    .A1(_01573_),
    .A2(_01604_));
 sg13g2_o21ai_1 _06858_ (.B1(net478),
    .Y(_01606_),
    .A1(_01297_),
    .A2(_01513_));
 sg13g2_buf_1 _06859_ (.A(_01606_),
    .X(_01607_));
 sg13g2_nand2_1 _06860_ (.Y(_01608_),
    .A(_00853_),
    .B(_01507_));
 sg13g2_nor2_2 _06861_ (.A(_00861_),
    .B(_01608_),
    .Y(_01609_));
 sg13g2_nand2_1 _06862_ (.Y(_01610_),
    .A(_00120_),
    .B(net352));
 sg13g2_a21oi_1 _06863_ (.A1(net449),
    .A2(_00119_),
    .Y(_01611_),
    .B1(net50));
 sg13g2_o21ai_1 _06864_ (.B1(_01611_),
    .Y(_01612_),
    .A1(_01609_),
    .A2(_01610_));
 sg13g2_nand2_1 _06865_ (.Y(_01613_),
    .A(net262),
    .B(net161));
 sg13g2_buf_1 _06866_ (.A(_01613_),
    .X(_01614_));
 sg13g2_nor2_2 _06867_ (.A(_01302_),
    .B(_01613_),
    .Y(_01615_));
 sg13g2_a221oi_1 _06868_ (.B2(_01615_),
    .C1(net353),
    .B1(_00840_),
    .A1(_01246_),
    .Y(_01616_),
    .A2(net66));
 sg13g2_nor2_1 _06869_ (.A(_01612_),
    .B(_01616_),
    .Y(_01617_));
 sg13g2_a21oi_1 _06870_ (.A1(_01246_),
    .A2(net39),
    .Y(_01618_),
    .B1(_01617_));
 sg13g2_nand3_1 _06871_ (.B(_01330_),
    .C(net255),
    .A(net453),
    .Y(_01619_));
 sg13g2_o21ai_1 _06872_ (.B1(_01619_),
    .Y(_00045_),
    .A1(_01607_),
    .A2(_01618_));
 sg13g2_o21ai_1 _06873_ (.B1(_01319_),
    .Y(_01620_),
    .A1(_00122_),
    .A2(_01609_));
 sg13g2_a21oi_1 _06874_ (.A1(net348),
    .A2(_00121_),
    .Y(_01621_),
    .B1(_01607_));
 sg13g2_and2_1 _06875_ (.A(net262),
    .B(_05112_),
    .X(_01622_));
 sg13g2_buf_1 _06876_ (.A(_01622_),
    .X(_01623_));
 sg13g2_buf_1 _06877_ (.A(_01623_),
    .X(_01624_));
 sg13g2_nand2b_1 _06878_ (.Y(_01625_),
    .B(net65),
    .A_N(_01302_));
 sg13g2_buf_2 _06879_ (.A(_01625_),
    .X(_01626_));
 sg13g2_inv_1 _06880_ (.Y(_01627_),
    .A(_00122_));
 sg13g2_a21oi_1 _06881_ (.A1(_01627_),
    .A2(net66),
    .Y(_01628_),
    .B1(net353));
 sg13g2_o21ai_1 _06882_ (.B1(_01628_),
    .Y(_01629_),
    .A1(_00913_),
    .A2(_01626_));
 sg13g2_nand3_1 _06883_ (.B(_01621_),
    .C(_01629_),
    .A(_01620_),
    .Y(_01630_));
 sg13g2_nor2_1 _06884_ (.A(net53),
    .B(_01607_),
    .Y(_01631_));
 sg13g2_a22oi_1 _06885_ (.Y(_01632_),
    .B1(_01631_),
    .B2(_01627_),
    .A2(_01525_),
    .A1(_01330_));
 sg13g2_nand2_1 _06886_ (.Y(_00046_),
    .A(_01630_),
    .B(_01632_));
 sg13g2_o21ai_1 _06887_ (.B1(net157),
    .Y(_01633_),
    .A1(_00124_),
    .A2(_01609_));
 sg13g2_nand2_1 _06888_ (.Y(_01634_),
    .A(net348),
    .B(_00123_));
 sg13g2_nor2_1 _06889_ (.A(net45),
    .B(_01607_),
    .Y(_01635_));
 sg13g2_nand3_1 _06890_ (.B(_01634_),
    .C(_01635_),
    .A(_01633_),
    .Y(_01636_));
 sg13g2_inv_1 _06891_ (.Y(_01637_),
    .A(_00124_));
 sg13g2_a221oi_1 _06892_ (.B2(_01615_),
    .C1(net258),
    .B1(_00942_),
    .A1(_01637_),
    .Y(_01638_),
    .A2(net66));
 sg13g2_nor2_1 _06893_ (.A(_01338_),
    .B(_01513_),
    .Y(_01639_));
 sg13g2_a22oi_1 _06894_ (.Y(_01640_),
    .B1(_01631_),
    .B2(_01637_),
    .A2(_01639_),
    .A1(_01330_));
 sg13g2_o21ai_1 _06895_ (.B1(_01640_),
    .Y(_00048_),
    .A1(_01636_),
    .A2(_01638_));
 sg13g2_inv_1 _06896_ (.Y(_01641_),
    .A(_00126_));
 sg13g2_a221oi_1 _06897_ (.B2(_01615_),
    .C1(net258),
    .B1(_00962_),
    .A1(_01641_),
    .Y(_01642_),
    .A2(net66));
 sg13g2_o21ai_1 _06898_ (.B1(net157),
    .Y(_01643_),
    .A1(_00126_),
    .A2(_01609_));
 sg13g2_nand2_1 _06899_ (.Y(_01644_),
    .A(net348),
    .B(_00125_));
 sg13g2_nand3_1 _06900_ (.B(_01643_),
    .C(_01644_),
    .A(_01635_),
    .Y(_01645_));
 sg13g2_a22oi_1 _06901_ (.Y(_01646_),
    .B1(_01631_),
    .B2(_01641_),
    .A2(_01538_),
    .A1(_01330_));
 sg13g2_o21ai_1 _06902_ (.B1(_01646_),
    .Y(_00049_),
    .A1(_01642_),
    .A2(_01645_));
 sg13g2_inv_1 _06903_ (.Y(_01647_),
    .A(_00140_));
 sg13g2_nor2_1 _06904_ (.A(_01068_),
    .B(_01608_),
    .Y(_01648_));
 sg13g2_inv_1 _06905_ (.Y(_01649_),
    .A(_01648_));
 sg13g2_nor2_1 _06906_ (.A(_01647_),
    .B(_01152_),
    .Y(_01650_));
 sg13g2_a221oi_1 _06907_ (.B2(_01650_),
    .C1(net46),
    .B1(_01649_),
    .A1(net404),
    .Y(_01651_),
    .A2(_00139_));
 sg13g2_o21ai_1 _06908_ (.B1(net351),
    .Y(_01652_),
    .A1(_00140_),
    .A2(net65));
 sg13g2_inv_1 _06909_ (.Y(_01653_),
    .A(_01652_));
 sg13g2_o21ai_1 _06910_ (.B1(_01653_),
    .Y(_01654_),
    .A1(_01067_),
    .A2(_01626_));
 sg13g2_a22oi_1 _06911_ (.Y(_01655_),
    .B1(_01651_),
    .B2(_01654_),
    .A2(net39),
    .A1(_01647_));
 sg13g2_nand3_1 _06912_ (.B(_01296_),
    .C(net255),
    .A(net450),
    .Y(_01656_));
 sg13g2_buf_1 _06913_ (.A(_01656_),
    .X(_01657_));
 sg13g2_nand2_1 _06914_ (.Y(_01658_),
    .A(net452),
    .B(_01657_));
 sg13g2_and3_1 _06915_ (.X(_01659_),
    .A(net450),
    .B(_01296_),
    .C(net255));
 sg13g2_buf_1 _06916_ (.A(_01659_),
    .X(_01660_));
 sg13g2_nand2_1 _06917_ (.Y(_01661_),
    .A(net453),
    .B(_01660_));
 sg13g2_o21ai_1 _06918_ (.B1(_01661_),
    .Y(_00050_),
    .A1(_01655_),
    .A2(_01658_));
 sg13g2_or2_1 _06919_ (.X(_01662_),
    .B(_01648_),
    .A(_00142_));
 sg13g2_a221oi_1 _06920_ (.B2(_01662_),
    .C1(_00846_),
    .B1(_01073_),
    .A1(net448),
    .Y(_01663_),
    .A2(_01441_));
 sg13g2_o21ai_1 _06921_ (.B1(net156),
    .Y(_01664_),
    .A1(net66),
    .A2(_01363_));
 sg13g2_a21oi_1 _06922_ (.A1(net66),
    .A2(_01663_),
    .Y(_01665_),
    .B1(net50));
 sg13g2_o21ai_1 _06923_ (.B1(_01657_),
    .Y(_01666_),
    .A1(_00142_),
    .A2(_01665_));
 sg13g2_a21oi_1 _06924_ (.A1(_01663_),
    .A2(_01664_),
    .Y(_01667_),
    .B1(_01666_));
 sg13g2_nand2_1 _06925_ (.Y(_01668_),
    .A(net405),
    .B(_01657_));
 sg13g2_o21ai_1 _06926_ (.B1(_01668_),
    .Y(_01669_),
    .A1(_00921_),
    .A2(_01657_));
 sg13g2_nor2_1 _06927_ (.A(_01667_),
    .B(_01669_),
    .Y(_00051_));
 sg13g2_inv_1 _06928_ (.Y(_01670_),
    .A(_00144_));
 sg13g2_nand2_1 _06929_ (.Y(_01671_),
    .A(_01670_),
    .B(_01649_));
 sg13g2_a221oi_1 _06930_ (.B2(_01671_),
    .C1(net46),
    .B1(net257),
    .A1(net404),
    .Y(_01672_),
    .A2(_00143_));
 sg13g2_o21ai_1 _06931_ (.B1(net256),
    .Y(_01673_),
    .A1(_00144_),
    .A2(net65));
 sg13g2_inv_1 _06932_ (.Y(_01674_),
    .A(_01673_));
 sg13g2_o21ai_1 _06933_ (.B1(_01674_),
    .Y(_01675_),
    .A1(_01149_),
    .A2(_01626_));
 sg13g2_a22oi_1 _06934_ (.Y(_01676_),
    .B1(_01672_),
    .B2(_01675_),
    .A2(net39),
    .A1(_01670_));
 sg13g2_nand2_1 _06935_ (.Y(_01677_),
    .A(net477),
    .B(_01660_));
 sg13g2_o21ai_1 _06936_ (.B1(_01677_),
    .Y(_00052_),
    .A1(_01658_),
    .A2(_01676_));
 sg13g2_o21ai_1 _06937_ (.B1(net257),
    .Y(_01678_),
    .A1(_01460_),
    .A2(_01648_));
 sg13g2_a21oi_1 _06938_ (.A1(net406),
    .A2(_00145_),
    .Y(_01679_),
    .B1(net46));
 sg13g2_nand4_1 _06939_ (.B(_01657_),
    .C(_01678_),
    .A(net403),
    .Y(_01680_),
    .D(_01679_));
 sg13g2_o21ai_1 _06940_ (.B1(net156),
    .Y(_01681_),
    .A1(_01460_),
    .A2(net65));
 sg13g2_a21oi_1 _06941_ (.A1(_01177_),
    .A2(_01615_),
    .Y(_01682_),
    .B1(_01681_));
 sg13g2_nor3_1 _06942_ (.A(_01460_),
    .B(net48),
    .C(_01658_),
    .Y(_01683_));
 sg13g2_a21oi_1 _06943_ (.A1(net476),
    .A2(_01660_),
    .Y(_01684_),
    .B1(_01683_));
 sg13g2_o21ai_1 _06944_ (.B1(_01684_),
    .Y(_00053_),
    .A1(_01680_),
    .A2(_01682_));
 sg13g2_nand2_1 _06945_ (.Y(_01685_),
    .A(_01398_),
    .B(_01503_));
 sg13g2_nand2_1 _06946_ (.Y(_01686_),
    .A(_05057_),
    .B(_01685_));
 sg13g2_inv_1 _06947_ (.Y(_01687_),
    .A(_00152_));
 sg13g2_nor2_1 _06948_ (.A(_01389_),
    .B(_01608_),
    .Y(_01688_));
 sg13g2_inv_1 _06949_ (.Y(_01689_),
    .A(_01688_));
 sg13g2_nor2_1 _06950_ (.A(_01687_),
    .B(net350),
    .Y(_01690_));
 sg13g2_a221oi_1 _06951_ (.B2(_01690_),
    .C1(net46),
    .B1(_01689_),
    .A1(net404),
    .Y(_01691_),
    .A2(_00151_));
 sg13g2_o21ai_1 _06952_ (.B1(net351),
    .Y(_01692_),
    .A1(_00152_),
    .A2(net65));
 sg13g2_inv_1 _06953_ (.Y(_01693_),
    .A(_01692_));
 sg13g2_o21ai_1 _06954_ (.B1(_01693_),
    .Y(_01694_),
    .A1(_01194_),
    .A2(_01626_));
 sg13g2_a22oi_1 _06955_ (.Y(_01695_),
    .B1(_01691_),
    .B2(_01694_),
    .A2(_01240_),
    .A1(_01687_));
 sg13g2_nand3_1 _06956_ (.B(_01398_),
    .C(_01504_),
    .A(_00895_),
    .Y(_01696_));
 sg13g2_o21ai_1 _06957_ (.B1(_01696_),
    .Y(_00054_),
    .A1(_01686_),
    .A2(_01695_));
 sg13g2_nor2_1 _06958_ (.A(_01215_),
    .B(_01626_),
    .Y(_01697_));
 sg13g2_o21ai_1 _06959_ (.B1(_01424_),
    .Y(_01698_),
    .A1(_00154_),
    .A2(_01624_));
 sg13g2_or2_1 _06960_ (.X(_01699_),
    .B(_01688_),
    .A(_00154_));
 sg13g2_a221oi_1 _06961_ (.B2(_01699_),
    .C1(_01686_),
    .B1(_01319_),
    .A1(net349),
    .Y(_01700_),
    .A2(_00153_));
 sg13g2_o21ai_1 _06962_ (.B1(_01700_),
    .Y(_01701_),
    .A1(_01697_),
    .A2(_01698_));
 sg13g2_or2_1 _06963_ (.X(_01702_),
    .B(_01686_),
    .A(_01079_));
 sg13g2_buf_1 _06964_ (.A(_01702_),
    .X(_01703_));
 sg13g2_nor2_1 _06965_ (.A(_00154_),
    .B(_01703_),
    .Y(_01704_));
 sg13g2_a21oi_1 _06966_ (.A1(net347),
    .A2(_01525_),
    .Y(_01705_),
    .B1(_01704_));
 sg13g2_nand2_1 _06967_ (.Y(_00055_),
    .A(_01701_),
    .B(_01705_));
 sg13g2_nand2b_1 _06968_ (.Y(_01706_),
    .B(net66),
    .A_N(_00156_));
 sg13g2_o21ai_1 _06969_ (.B1(_01706_),
    .Y(_01707_),
    .A1(_01220_),
    .A2(_01626_));
 sg13g2_or2_1 _06970_ (.X(_01708_),
    .B(_01688_),
    .A(_00156_));
 sg13g2_nand3_1 _06971_ (.B(net53),
    .C(_01685_),
    .A(net452),
    .Y(_01709_));
 sg13g2_a221oi_1 _06972_ (.B2(_01708_),
    .C1(_01709_),
    .B1(net157),
    .A1(net349),
    .Y(_01710_),
    .A2(_00155_));
 sg13g2_o21ai_1 _06973_ (.B1(_01710_),
    .Y(_01711_),
    .A1(net258),
    .A2(_01707_));
 sg13g2_nor2_1 _06974_ (.A(_00156_),
    .B(_01703_),
    .Y(_01712_));
 sg13g2_a21oi_1 _06975_ (.A1(net347),
    .A2(_01639_),
    .Y(_01713_),
    .B1(_01712_));
 sg13g2_nand2_1 _06976_ (.Y(_00056_),
    .A(_01711_),
    .B(_01713_));
 sg13g2_nor2_1 _06977_ (.A(_01226_),
    .B(_01626_),
    .Y(_01714_));
 sg13g2_o21ai_1 _06978_ (.B1(net156),
    .Y(_01715_),
    .A1(_00158_),
    .A2(_01624_));
 sg13g2_or2_1 _06979_ (.X(_01716_),
    .B(_01688_),
    .A(_00158_));
 sg13g2_a221oi_1 _06980_ (.B2(_01716_),
    .C1(_01709_),
    .B1(net157),
    .A1(net349),
    .Y(_01717_),
    .A2(_00157_));
 sg13g2_o21ai_1 _06981_ (.B1(_01717_),
    .Y(_01718_),
    .A1(_01714_),
    .A2(_01715_));
 sg13g2_nor2_1 _06982_ (.A(_00158_),
    .B(_01703_),
    .Y(_01719_));
 sg13g2_a21oi_1 _06983_ (.A1(net347),
    .A2(_01538_),
    .Y(_01720_),
    .B1(_01719_));
 sg13g2_nand2_1 _06984_ (.Y(_00057_),
    .A(_01718_),
    .B(_01720_));
 sg13g2_inv_1 _06985_ (.Y(_01721_),
    .A(_00159_));
 sg13g2_nand3_1 _06986_ (.B(_01249_),
    .C(_01507_),
    .A(_00853_),
    .Y(_01722_));
 sg13g2_nor2_1 _06987_ (.A(net456),
    .B(_01722_),
    .Y(_01723_));
 sg13g2_a21oi_1 _06988_ (.A1(net412),
    .A2(net65),
    .Y(_01724_),
    .B1(_01723_));
 sg13g2_nand2b_1 _06989_ (.Y(_01725_),
    .B(_01543_),
    .A_N(_01545_));
 sg13g2_o21ai_1 _06990_ (.B1(_00159_),
    .Y(_01726_),
    .A1(_01724_),
    .A2(_01725_));
 sg13g2_nor2_1 _06991_ (.A(net66),
    .B(_00987_),
    .Y(_01727_));
 sg13g2_o21ai_1 _06992_ (.B1(_01727_),
    .Y(_01728_),
    .A1(_01302_),
    .A2(_01242_));
 sg13g2_a22oi_1 _06993_ (.Y(_01729_),
    .B1(_01726_),
    .B2(_01728_),
    .A2(net39),
    .A1(_01721_));
 sg13g2_o21ai_1 _06994_ (.B1(net452),
    .Y(_01730_),
    .A1(_01430_),
    .A2(_01513_));
 sg13g2_nor2_2 _06995_ (.A(_01430_),
    .B(_01513_),
    .Y(_01731_));
 sg13g2_nand2_1 _06996_ (.Y(_01732_),
    .A(_00896_),
    .B(_01731_));
 sg13g2_o21ai_1 _06997_ (.B1(_01732_),
    .Y(_00059_),
    .A1(_01729_),
    .A2(_01730_));
 sg13g2_o21ai_1 _06998_ (.B1(net351),
    .Y(_01733_),
    .A1(_00160_),
    .A2(net65));
 sg13g2_a21o_1 _06999_ (.A2(_01615_),
    .A1(_01263_),
    .B1(_01733_),
    .X(_01734_));
 sg13g2_nor2_1 _07000_ (.A(_01152_),
    .B(_01722_),
    .Y(_01735_));
 sg13g2_nand2_1 _07001_ (.Y(_01736_),
    .A(_01152_),
    .B(_01543_));
 sg13g2_o21ai_1 _07002_ (.B1(_01736_),
    .Y(_01737_),
    .A1(_00160_),
    .A2(_01735_));
 sg13g2_nand4_1 _07003_ (.B(net447),
    .C(_01734_),
    .A(net480),
    .Y(_01738_),
    .D(_01737_));
 sg13g2_o21ai_1 _07004_ (.B1(_01738_),
    .Y(_01739_),
    .A1(_00160_),
    .A2(_01292_));
 sg13g2_mux2_1 _07005_ (.A0(_01739_),
    .A1(_00922_),
    .S(_01731_),
    .X(_00060_));
 sg13g2_inv_1 _07006_ (.Y(_01740_),
    .A(_00161_));
 sg13g2_a22oi_1 _07007_ (.Y(_01741_),
    .B1(_01275_),
    .B2(_01615_),
    .A2(_01614_),
    .A1(_01740_));
 sg13g2_a21oi_1 _07008_ (.A1(_01740_),
    .A2(_01722_),
    .Y(_01742_),
    .B1(net350));
 sg13g2_a21oi_1 _07009_ (.A1(net156),
    .A2(_01741_),
    .Y(_01743_),
    .B1(_01742_));
 sg13g2_a21oi_1 _07010_ (.A1(_00161_),
    .A2(_01356_),
    .Y(_01744_),
    .B1(_01730_));
 sg13g2_o21ai_1 _07011_ (.B1(_01744_),
    .Y(_01745_),
    .A1(net40),
    .A2(_01743_));
 sg13g2_o21ai_1 _07012_ (.B1(_01745_),
    .Y(_00061_),
    .A1(_01430_),
    .A2(_01527_));
 sg13g2_o21ai_1 _07013_ (.B1(_01736_),
    .Y(_01746_),
    .A1(_00162_),
    .A2(_01735_));
 sg13g2_o21ai_1 _07014_ (.B1(_01088_),
    .Y(_01747_),
    .A1(_00162_),
    .A2(net65));
 sg13g2_inv_1 _07015_ (.Y(_01748_),
    .A(_01747_));
 sg13g2_o21ai_1 _07016_ (.B1(_01748_),
    .Y(_01749_),
    .A1(_01283_),
    .A2(_01626_));
 sg13g2_nand4_1 _07017_ (.B(net447),
    .C(_01746_),
    .A(net480),
    .Y(_01750_),
    .D(_01749_));
 sg13g2_o21ai_1 _07018_ (.B1(_01750_),
    .Y(_01751_),
    .A1(_00162_),
    .A2(_01292_));
 sg13g2_mux2_1 _07019_ (.A0(_01751_),
    .A1(_00948_),
    .S(_01731_),
    .X(_00062_));
 sg13g2_buf_2 _07020_ (.A(\draw_game_inst.y[9] ),
    .X(_01752_));
 sg13g2_buf_1 _07021_ (.A(\draw_game_inst.board_y[4] ),
    .X(_01753_));
 sg13g2_buf_1 _07022_ (.A(_01753_),
    .X(_01754_));
 sg13g2_buf_1 _07023_ (.A(net446),
    .X(_01755_));
 sg13g2_buf_1 _07024_ (.A(_01755_),
    .X(_01756_));
 sg13g2_buf_1 _07025_ (.A(\draw_game_inst.y[8] ),
    .X(_01757_));
 sg13g2_buf_2 _07026_ (.A(\draw_game_inst.y[7] ),
    .X(_01758_));
 sg13g2_buf_1 _07027_ (.A(_01758_),
    .X(_01759_));
 sg13g2_buf_1 _07028_ (.A(\draw_game_inst.board_y[6] ),
    .X(_01760_));
 sg13g2_buf_1 _07029_ (.A(\draw_game_inst.board_y[5] ),
    .X(_01761_));
 sg13g2_buf_1 _07030_ (.A(net474),
    .X(_01762_));
 sg13g2_buf_1 _07031_ (.A(net444),
    .X(_01763_));
 sg13g2_nand4_1 _07032_ (.B(net445),
    .C(net475),
    .A(_01757_),
    .Y(_01764_),
    .D(net400));
 sg13g2_buf_2 _07033_ (.A(\draw_game_inst.board_y[1] ),
    .X(_01765_));
 sg13g2_buf_1 _07034_ (.A(_01765_),
    .X(_01766_));
 sg13g2_buf_1 _07035_ (.A(\draw_game_inst.board_y[2] ),
    .X(_01767_));
 sg13g2_nor2b_1 _07036_ (.A(_01767_),
    .B_N(\draw_game_inst.board_y[3] ),
    .Y(_01768_));
 sg13g2_buf_1 _07037_ (.A(_01768_),
    .X(_01769_));
 sg13g2_nand2_1 _07038_ (.Y(_01770_),
    .A(net443),
    .B(net399));
 sg13g2_buf_2 _07039_ (.A(_01770_),
    .X(_01771_));
 sg13g2_or4_1 _07040_ (.A(_01752_),
    .B(net346),
    .C(_01764_),
    .D(_01771_),
    .X(_00068_));
 sg13g2_buf_1 _07041_ (.A(\draw_game_inst.x[8] ),
    .X(_01772_));
 sg13g2_inv_1 _07042_ (.Y(_01773_),
    .A(_01772_));
 sg13g2_buf_2 _07043_ (.A(\draw_game_inst.x[9] ),
    .X(_01774_));
 sg13g2_buf_1 _07044_ (.A(\draw_game_inst.x[7] ),
    .X(_01775_));
 sg13g2_buf_2 _07045_ (.A(net473),
    .X(_01776_));
 sg13g2_buf_1 _07046_ (.A(_01776_),
    .X(_01777_));
 sg13g2_buf_1 _07047_ (.A(\draw_game_inst.x[6] ),
    .X(_01778_));
 sg13g2_buf_1 _07048_ (.A(net472),
    .X(_01779_));
 sg13g2_buf_1 _07049_ (.A(net441),
    .X(_01780_));
 sg13g2_buf_1 _07050_ (.A(\draw_game_inst.board_x[5] ),
    .X(_01781_));
 sg13g2_buf_1 _07051_ (.A(net471),
    .X(_01782_));
 sg13g2_buf_1 _07052_ (.A(\draw_game_inst.board_x[4] ),
    .X(_01783_));
 sg13g2_buf_1 _07053_ (.A(net470),
    .X(_01784_));
 sg13g2_and2_1 _07054_ (.A(_01782_),
    .B(net439),
    .X(_01785_));
 sg13g2_buf_2 _07055_ (.A(_01785_),
    .X(_01786_));
 sg13g2_or2_1 _07056_ (.X(_01787_),
    .B(net470),
    .A(net471));
 sg13g2_buf_1 _07057_ (.A(_01787_),
    .X(_01788_));
 sg13g2_buf_1 _07058_ (.A(_01788_),
    .X(_01789_));
 sg13g2_nor2_1 _07059_ (.A(net397),
    .B(net345),
    .Y(_01790_));
 sg13g2_a21oi_1 _07060_ (.A1(_01780_),
    .A2(_01786_),
    .Y(_01791_),
    .B1(_01790_));
 sg13g2_nand4_1 _07061_ (.B(_01774_),
    .C(net398),
    .A(_01773_),
    .Y(_00067_),
    .D(_01791_));
 sg13g2_nor2b_1 _07062_ (.A(vsync_prev),
    .B_N(\vga_sync_gen.vsync ),
    .Y(_01792_));
 sg13g2_buf_2 _07063_ (.A(_01792_),
    .X(_01793_));
 sg13g2_buf_1 _07064_ (.A(_01793_),
    .X(_01794_));
 sg13g2_buf_1 _07065_ (.A(\draw_game_inst.new_tiles_counter[1] ),
    .X(_01795_));
 sg13g2_buf_1 _07066_ (.A(\draw_game_inst.new_tiles_counter[2] ),
    .X(_01796_));
 sg13g2_or2_1 _07067_ (.X(_01797_),
    .B(\new_tiles_counter[0] ),
    .A(\draw_game_inst.new_tiles_counter[0] ));
 sg13g2_buf_1 _07068_ (.A(_01797_),
    .X(_01798_));
 sg13g2_nor3_1 _07069_ (.A(_01795_),
    .B(_01796_),
    .C(_01798_),
    .Y(_01799_));
 sg13g2_nor2b_1 _07070_ (.A(\new_tiles_counter[4] ),
    .B_N(_01799_),
    .Y(_01800_));
 sg13g2_nand3_1 _07071_ (.B(net396),
    .C(_01800_),
    .A(net403),
    .Y(_01801_));
 sg13g2_and2_1 _07072_ (.A(\draw_game_inst.new_tiles[0] ),
    .B(_01801_),
    .X(_00395_));
 sg13g2_buf_1 _07073_ (.A(net405),
    .X(_01802_));
 sg13g2_buf_1 _07074_ (.A(\game_logic_inst.added_tile_index[2] ),
    .X(_01803_));
 sg13g2_buf_1 _07075_ (.A(\game_logic_inst.added_tile_index[3] ),
    .X(_01804_));
 sg13g2_nor2b_1 _07076_ (.A(_01803_),
    .B_N(_01804_),
    .Y(_01805_));
 sg13g2_buf_1 _07077_ (.A(\game_logic_inst.added_tile_index[0] ),
    .X(_01806_));
 sg13g2_buf_1 _07078_ (.A(\game_logic_inst.added_tile_index[1] ),
    .X(_01807_));
 sg13g2_nor2b_1 _07079_ (.A(_01806_),
    .B_N(_01807_),
    .Y(_01808_));
 sg13g2_nand2_1 _07080_ (.Y(_01809_),
    .A(_01805_),
    .B(_01808_));
 sg13g2_a21o_1 _07081_ (.A2(_01800_),
    .A1(_01793_),
    .B1(_05058_),
    .X(_01810_));
 sg13g2_buf_1 _07082_ (.A(_01810_),
    .X(_01811_));
 sg13g2_buf_1 _07083_ (.A(_01811_),
    .X(_01812_));
 sg13g2_a21oi_1 _07084_ (.A1(_00080_),
    .A2(_01809_),
    .Y(_01813_),
    .B1(net91));
 sg13g2_a21o_1 _07085_ (.A2(\draw_game_inst.new_tiles[10] ),
    .A1(net344),
    .B1(_01813_),
    .X(_00396_));
 sg13g2_and2_1 _07086_ (.A(_01807_),
    .B(_01806_),
    .X(_01814_));
 sg13g2_buf_1 _07087_ (.A(_01814_),
    .X(_01815_));
 sg13g2_inv_1 _07088_ (.Y(_01816_),
    .A(_00081_));
 sg13g2_a21oi_1 _07089_ (.A1(_01805_),
    .A2(_01815_),
    .Y(_01817_),
    .B1(_01816_));
 sg13g2_nand2_1 _07090_ (.Y(_01818_),
    .A(net413),
    .B(\draw_game_inst.new_tiles[11] ));
 sg13g2_o21ai_1 _07091_ (.B1(_01818_),
    .Y(_00397_),
    .A1(net91),
    .A2(_01817_));
 sg13g2_nor2_1 _07092_ (.A(_01807_),
    .B(_01806_),
    .Y(_01819_));
 sg13g2_and2_1 _07093_ (.A(_01804_),
    .B(_01803_),
    .X(_01820_));
 sg13g2_buf_1 _07094_ (.A(_01820_),
    .X(_01821_));
 sg13g2_inv_1 _07095_ (.Y(_01822_),
    .A(_00082_));
 sg13g2_a21oi_1 _07096_ (.A1(_01819_),
    .A2(_01821_),
    .Y(_01823_),
    .B1(_01822_));
 sg13g2_nand2_1 _07097_ (.Y(_01824_),
    .A(net413),
    .B(\draw_game_inst.new_tiles[12] ));
 sg13g2_o21ai_1 _07098_ (.B1(_01824_),
    .Y(_00398_),
    .A1(net91),
    .A2(_01823_));
 sg13g2_nor2b_1 _07099_ (.A(_01807_),
    .B_N(_01806_),
    .Y(_01825_));
 sg13g2_inv_1 _07100_ (.Y(_01826_),
    .A(_00083_));
 sg13g2_a21oi_1 _07101_ (.A1(_01821_),
    .A2(_01825_),
    .Y(_01827_),
    .B1(_01826_));
 sg13g2_nand2_1 _07102_ (.Y(_01828_),
    .A(net413),
    .B(\draw_game_inst.new_tiles[13] ));
 sg13g2_o21ai_1 _07103_ (.B1(_01828_),
    .Y(_00399_),
    .A1(net91),
    .A2(_01827_));
 sg13g2_inv_1 _07104_ (.Y(_01829_),
    .A(_00084_));
 sg13g2_a21oi_1 _07105_ (.A1(_01808_),
    .A2(_01821_),
    .Y(_01830_),
    .B1(_01829_));
 sg13g2_nand2_1 _07106_ (.Y(_01831_),
    .A(net413),
    .B(\draw_game_inst.new_tiles[14] ));
 sg13g2_o21ai_1 _07107_ (.B1(_01831_),
    .Y(_00400_),
    .A1(_01812_),
    .A2(_01830_));
 sg13g2_inv_1 _07108_ (.Y(_01832_),
    .A(_00085_));
 sg13g2_a21oi_1 _07109_ (.A1(_01815_),
    .A2(_01821_),
    .Y(_01833_),
    .B1(_01832_));
 sg13g2_nand2_1 _07110_ (.Y(_01834_),
    .A(net413),
    .B(\draw_game_inst.new_tiles[15] ));
 sg13g2_o21ai_1 _07111_ (.B1(_01834_),
    .Y(_00401_),
    .A1(_01812_),
    .A2(_01833_));
 sg13g2_nor2_1 _07112_ (.A(_01804_),
    .B(_01803_),
    .Y(_01835_));
 sg13g2_nand2_1 _07113_ (.Y(_01836_),
    .A(_01825_),
    .B(_01835_));
 sg13g2_a21oi_1 _07114_ (.A1(_00071_),
    .A2(_01836_),
    .Y(_01837_),
    .B1(net91));
 sg13g2_a21o_1 _07115_ (.A2(\draw_game_inst.new_tiles[1] ),
    .A1(_01802_),
    .B1(_01837_),
    .X(_00402_));
 sg13g2_nand2_1 _07116_ (.Y(_01838_),
    .A(_01808_),
    .B(_01835_));
 sg13g2_a21oi_1 _07117_ (.A1(_00072_),
    .A2(_01838_),
    .Y(_01839_),
    .B1(net91));
 sg13g2_a21o_1 _07118_ (.A2(\draw_game_inst.new_tiles[2] ),
    .A1(net344),
    .B1(_01839_),
    .X(_00403_));
 sg13g2_inv_1 _07119_ (.Y(_01840_),
    .A(_00073_));
 sg13g2_a21oi_1 _07120_ (.A1(_01815_),
    .A2(_01835_),
    .Y(_01841_),
    .B1(_01840_));
 sg13g2_nand2_1 _07121_ (.Y(_01842_),
    .A(_05060_),
    .B(\draw_game_inst.new_tiles[3] ));
 sg13g2_o21ai_1 _07122_ (.B1(_01842_),
    .Y(_00404_),
    .A1(net91),
    .A2(_01841_));
 sg13g2_nor2b_1 _07123_ (.A(_01804_),
    .B_N(_01803_),
    .Y(_01843_));
 sg13g2_nand2_1 _07124_ (.Y(_01844_),
    .A(_01819_),
    .B(_01843_));
 sg13g2_a21oi_1 _07125_ (.A1(_00074_),
    .A2(_01844_),
    .Y(_01845_),
    .B1(_01811_));
 sg13g2_a21o_1 _07126_ (.A2(\draw_game_inst.new_tiles[4] ),
    .A1(net344),
    .B1(_01845_),
    .X(_00405_));
 sg13g2_nand2_1 _07127_ (.Y(_01846_),
    .A(_01825_),
    .B(_01843_));
 sg13g2_a21oi_1 _07128_ (.A1(_00075_),
    .A2(_01846_),
    .Y(_01847_),
    .B1(_01811_));
 sg13g2_a21o_1 _07129_ (.A2(\draw_game_inst.new_tiles[5] ),
    .A1(_01802_),
    .B1(_01847_),
    .X(_00406_));
 sg13g2_nand2_1 _07130_ (.Y(_01848_),
    .A(_01808_),
    .B(_01843_));
 sg13g2_a21oi_1 _07131_ (.A1(_00076_),
    .A2(_01848_),
    .Y(_01849_),
    .B1(_01811_));
 sg13g2_a21o_1 _07132_ (.A2(\draw_game_inst.new_tiles[6] ),
    .A1(net344),
    .B1(_01849_),
    .X(_00407_));
 sg13g2_inv_1 _07133_ (.Y(_01850_),
    .A(_00077_));
 sg13g2_a21oi_1 _07134_ (.A1(_01815_),
    .A2(_01843_),
    .Y(_01851_),
    .B1(_01850_));
 sg13g2_nand2_1 _07135_ (.Y(_01852_),
    .A(_05060_),
    .B(\draw_game_inst.new_tiles[7] ));
 sg13g2_o21ai_1 _07136_ (.B1(_01852_),
    .Y(_00408_),
    .A1(net91),
    .A2(_01851_));
 sg13g2_nand2_1 _07137_ (.Y(_01853_),
    .A(_01805_),
    .B(_01819_));
 sg13g2_a21oi_1 _07138_ (.A1(_00078_),
    .A2(_01853_),
    .Y(_01854_),
    .B1(_01811_));
 sg13g2_a21o_1 _07139_ (.A2(\draw_game_inst.new_tiles[8] ),
    .A1(net344),
    .B1(_01854_),
    .X(_00409_));
 sg13g2_nand2_1 _07140_ (.Y(_01855_),
    .A(_01805_),
    .B(_01825_));
 sg13g2_a21oi_1 _07141_ (.A1(_00079_),
    .A2(_01855_),
    .Y(_01856_),
    .B1(_01811_));
 sg13g2_a21o_1 _07142_ (.A2(\draw_game_inst.new_tiles[9] ),
    .A1(net344),
    .B1(_01856_),
    .X(_00410_));
 sg13g2_and2_1 _07143_ (.A(_01819_),
    .B(_01835_),
    .X(_01857_));
 sg13g2_buf_1 _07144_ (.A(_01857_),
    .X(_01858_));
 sg13g2_nand2_1 _07145_ (.Y(_01859_),
    .A(_00086_),
    .B(_01858_));
 sg13g2_nand2b_1 _07146_ (.Y(_01860_),
    .B(\vga_sync_gen.vsync ),
    .A_N(vsync_prev));
 sg13g2_buf_1 _07147_ (.A(_01860_),
    .X(_01861_));
 sg13g2_nor2_2 _07148_ (.A(net438),
    .B(_01800_),
    .Y(_01862_));
 sg13g2_mux2_1 _07149_ (.A0(_01859_),
    .A1(_00086_),
    .S(_01862_),
    .X(_01863_));
 sg13g2_buf_1 _07150_ (.A(net407),
    .X(_01864_));
 sg13g2_mux2_1 _07151_ (.A0(\new_tiles_counter[0] ),
    .A1(_01863_),
    .S(net343),
    .X(_00411_));
 sg13g2_nor2b_1 _07152_ (.A(_01862_),
    .B_N(_01858_),
    .Y(_01865_));
 sg13g2_inv_1 _07153_ (.Y(_01866_),
    .A(_01865_));
 sg13g2_nand2b_1 _07154_ (.Y(_01867_),
    .B(_01862_),
    .A_N(_01798_));
 sg13g2_o21ai_1 _07155_ (.B1(_01867_),
    .Y(_01868_),
    .A1(_00087_),
    .A2(_01866_));
 sg13g2_a21o_1 _07156_ (.A2(net396),
    .A1(\new_tiles_counter[0] ),
    .B1(_05059_),
    .X(_01869_));
 sg13g2_a22oi_1 _07157_ (.Y(_01870_),
    .B1(_01869_),
    .B2(\draw_game_inst.new_tiles_counter[0] ),
    .A2(_01868_),
    .A1(net402));
 sg13g2_inv_1 _07158_ (.Y(_00412_),
    .A(_01870_));
 sg13g2_or3_1 _07159_ (.A(_05058_),
    .B(_01795_),
    .C(_01798_),
    .X(_01871_));
 sg13g2_buf_1 _07160_ (.A(_01871_),
    .X(_01872_));
 sg13g2_nand2_1 _07161_ (.Y(_01873_),
    .A(_01795_),
    .B(_01798_));
 sg13g2_nand2_1 _07162_ (.Y(_01874_),
    .A(_01872_),
    .B(_01873_));
 sg13g2_nand2_1 _07163_ (.Y(_01875_),
    .A(net407),
    .B(_01866_));
 sg13g2_a22oi_1 _07164_ (.Y(_01876_),
    .B1(_01875_),
    .B2(_01795_),
    .A2(_01874_),
    .A1(_01862_));
 sg13g2_inv_1 _07165_ (.Y(_00413_),
    .A(_01876_));
 sg13g2_o21ai_1 _07166_ (.B1(_01253_),
    .Y(_01877_),
    .A1(_01861_),
    .A2(_01799_));
 sg13g2_buf_1 _07167_ (.A(_01861_),
    .X(_01878_));
 sg13g2_o21ai_1 _07168_ (.B1(_01796_),
    .Y(_01879_),
    .A1(_01878_),
    .A2(_01872_));
 sg13g2_o21ai_1 _07169_ (.B1(_01879_),
    .Y(_00414_),
    .A1(_01865_),
    .A2(_01877_));
 sg13g2_nor2_1 _07170_ (.A(_01796_),
    .B(_01872_),
    .Y(_01880_));
 sg13g2_nor2_1 _07171_ (.A(_01858_),
    .B(_01877_),
    .Y(_01881_));
 sg13g2_nor2_1 _07172_ (.A(\new_tiles_counter[4] ),
    .B(_01881_),
    .Y(_01882_));
 sg13g2_a21oi_1 _07173_ (.A1(_01862_),
    .A2(_01880_),
    .Y(_00415_),
    .B1(_01882_));
 sg13g2_buf_1 _07174_ (.A(\draw_game_inst.board_y[0] ),
    .X(_01883_));
 sg13g2_buf_1 _07175_ (.A(_01883_),
    .X(_01884_));
 sg13g2_buf_1 _07176_ (.A(net437),
    .X(_01885_));
 sg13g2_buf_1 _07177_ (.A(net394),
    .X(_01886_));
 sg13g2_buf_2 _07178_ (.A(net342),
    .X(_01887_));
 sg13g2_buf_1 _07179_ (.A(net254),
    .X(_01888_));
 sg13g2_buf_1 _07180_ (.A(net155),
    .X(_01889_));
 sg13g2_buf_1 _07181_ (.A(\draw_game_inst.board_x[1] ),
    .X(_01890_));
 sg13g2_buf_1 _07182_ (.A(\draw_game_inst.board_x[0] ),
    .X(_01891_));
 sg13g2_buf_2 _07183_ (.A(\draw_game_inst.board_x[2] ),
    .X(_01892_));
 sg13g2_nand3_1 _07184_ (.B(net469),
    .C(_01892_),
    .A(_01890_),
    .Y(_01893_));
 sg13g2_buf_1 _07185_ (.A(_01893_),
    .X(_01894_));
 sg13g2_buf_1 _07186_ (.A(net471),
    .X(_01895_));
 sg13g2_buf_1 _07187_ (.A(\draw_game_inst.board_x[3] ),
    .X(_01896_));
 sg13g2_buf_1 _07188_ (.A(_01896_),
    .X(_01897_));
 sg13g2_nand3b_1 _07189_ (.B(_01784_),
    .C(_01897_),
    .Y(_01898_),
    .A_N(net436));
 sg13g2_buf_2 _07190_ (.A(_01898_),
    .X(_01899_));
 sg13g2_buf_1 _07191_ (.A(_01899_),
    .X(_01900_));
 sg13g2_buf_1 _07192_ (.A(net253),
    .X(_01901_));
 sg13g2_or2_1 _07193_ (.X(_01902_),
    .B(net154),
    .A(_01894_));
 sg13g2_nand2_1 _07194_ (.Y(_01903_),
    .A(_01772_),
    .B(_01774_));
 sg13g2_nor4_2 _07195_ (.A(net398),
    .B(_01779_),
    .C(_01902_),
    .Y(_01904_),
    .D(_01903_));
 sg13g2_nor2_1 _07196_ (.A(_05058_),
    .B(_01904_),
    .Y(_01905_));
 sg13g2_buf_2 _07197_ (.A(_01905_),
    .X(_01906_));
 sg13g2_inv_1 _07198_ (.Y(_01907_),
    .A(_01904_));
 sg13g2_buf_1 _07199_ (.A(\draw_game_inst.board_y[3] ),
    .X(_01908_));
 sg13g2_buf_1 _07200_ (.A(_01767_),
    .X(_01909_));
 sg13g2_nand2_1 _07201_ (.Y(_01910_),
    .A(_01908_),
    .B(net434));
 sg13g2_buf_1 _07202_ (.A(_01910_),
    .X(_01911_));
 sg13g2_buf_1 _07203_ (.A(net341),
    .X(_01912_));
 sg13g2_inv_2 _07204_ (.Y(_01913_),
    .A(_01753_));
 sg13g2_nor4_1 _07205_ (.A(_01757_),
    .B(net445),
    .C(net475),
    .D(net400),
    .Y(_01914_));
 sg13g2_nor2_1 _07206_ (.A(_01765_),
    .B(net437),
    .Y(_01915_));
 sg13g2_buf_1 _07207_ (.A(_01915_),
    .X(_01916_));
 sg13g2_buf_1 _07208_ (.A(_01916_),
    .X(_01917_));
 sg13g2_buf_1 _07209_ (.A(net251),
    .X(_01918_));
 sg13g2_buf_1 _07210_ (.A(net153),
    .X(_01919_));
 sg13g2_nand4_1 _07211_ (.B(_01913_),
    .C(_01914_),
    .A(_01752_),
    .Y(_01920_),
    .D(net89));
 sg13g2_o21ai_1 _07212_ (.B1(_05057_),
    .Y(_01921_),
    .A1(net252),
    .A2(_01920_));
 sg13g2_buf_2 _07213_ (.A(_01921_),
    .X(_01922_));
 sg13g2_nor2_1 _07214_ (.A(_01907_),
    .B(_01922_),
    .Y(_01923_));
 sg13g2_buf_1 _07215_ (.A(_01923_),
    .X(_01924_));
 sg13g2_buf_1 _07216_ (.A(_00164_),
    .X(_01925_));
 sg13g2_buf_1 _07217_ (.A(_01925_),
    .X(_01926_));
 sg13g2_a22oi_1 _07218_ (.Y(_01927_),
    .B1(net38),
    .B2(net433),
    .A2(_01906_),
    .A1(net90));
 sg13g2_inv_1 _07219_ (.Y(_00427_),
    .A(_01927_));
 sg13g2_inv_1 _07220_ (.Y(_01928_),
    .A(_01765_));
 sg13g2_buf_1 _07221_ (.A(_01928_),
    .X(_01929_));
 sg13g2_buf_1 _07222_ (.A(net393),
    .X(_01930_));
 sg13g2_buf_1 _07223_ (.A(_01930_),
    .X(_01931_));
 sg13g2_buf_1 _07224_ (.A(net250),
    .X(_01932_));
 sg13g2_nand2_1 _07225_ (.Y(_01933_),
    .A(net90),
    .B(_01904_));
 sg13g2_xnor2_1 _07226_ (.Y(_01934_),
    .A(net152),
    .B(_01933_));
 sg13g2_nor2_1 _07227_ (.A(net361),
    .B(_01934_),
    .Y(_00428_));
 sg13g2_buf_1 _07228_ (.A(net434),
    .X(_01935_));
 sg13g2_buf_1 _07229_ (.A(net392),
    .X(_01936_));
 sg13g2_buf_1 _07230_ (.A(net339),
    .X(_01937_));
 sg13g2_buf_1 _07231_ (.A(net249),
    .X(_01938_));
 sg13g2_and2_1 _07232_ (.A(_01765_),
    .B(net437),
    .X(_01939_));
 sg13g2_buf_1 _07233_ (.A(_01939_),
    .X(_01940_));
 sg13g2_buf_2 _07234_ (.A(net338),
    .X(_01941_));
 sg13g2_buf_1 _07235_ (.A(net248),
    .X(_01942_));
 sg13g2_buf_1 _07236_ (.A(net150),
    .X(_01943_));
 sg13g2_nand2_1 _07237_ (.Y(_01944_),
    .A(net478),
    .B(_01907_));
 sg13g2_buf_2 _07238_ (.A(_01944_),
    .X(_01945_));
 sg13g2_o21ai_1 _07239_ (.B1(_01945_),
    .Y(_01946_),
    .A1(_01922_),
    .A2(net88));
 sg13g2_nand2_1 _07240_ (.Y(_01947_),
    .A(_01765_),
    .B(_01883_));
 sg13g2_buf_1 _07241_ (.A(_01947_),
    .X(_01948_));
 sg13g2_buf_1 _07242_ (.A(_01948_),
    .X(_01949_));
 sg13g2_nor2_1 _07243_ (.A(net392),
    .B(net337),
    .Y(_01950_));
 sg13g2_a22oi_1 _07244_ (.Y(_01951_),
    .B1(_01950_),
    .B2(net38),
    .A2(_01946_),
    .A1(net151));
 sg13g2_inv_1 _07245_ (.Y(_00429_),
    .A(_01951_));
 sg13g2_buf_1 _07246_ (.A(net434),
    .X(_01952_));
 sg13g2_buf_1 _07247_ (.A(net443),
    .X(_01953_));
 sg13g2_buf_1 _07248_ (.A(_01883_),
    .X(_01954_));
 sg13g2_buf_1 _07249_ (.A(net432),
    .X(_01955_));
 sg13g2_nand3_1 _07250_ (.B(net390),
    .C(net389),
    .A(net391),
    .Y(_01956_));
 sg13g2_buf_1 _07251_ (.A(_01956_),
    .X(_01957_));
 sg13g2_nor2b_1 _07252_ (.A(_01922_),
    .B_N(_01957_),
    .Y(_01958_));
 sg13g2_buf_1 _07253_ (.A(net468),
    .X(_01959_));
 sg13g2_buf_2 _07254_ (.A(net431),
    .X(_01960_));
 sg13g2_buf_1 _07255_ (.A(net388),
    .X(_01961_));
 sg13g2_buf_1 _07256_ (.A(net336),
    .X(_01962_));
 sg13g2_buf_1 _07257_ (.A(_01962_),
    .X(_01963_));
 sg13g2_buf_1 _07258_ (.A(net149),
    .X(_01964_));
 sg13g2_o21ai_1 _07259_ (.B1(net87),
    .Y(_01965_),
    .A1(_01906_),
    .A2(_01958_));
 sg13g2_inv_1 _07260_ (.Y(_01966_),
    .A(_01767_));
 sg13g2_buf_1 _07261_ (.A(_01966_),
    .X(_01967_));
 sg13g2_nor2_1 _07262_ (.A(_01908_),
    .B(net387),
    .Y(_01968_));
 sg13g2_buf_1 _07263_ (.A(_01968_),
    .X(_01969_));
 sg13g2_nand3_1 _07264_ (.B(net88),
    .C(net246),
    .A(net38),
    .Y(_01970_));
 sg13g2_nand2_1 _07265_ (.Y(_00430_),
    .A(_01965_),
    .B(_01970_));
 sg13g2_buf_1 _07266_ (.A(_01948_),
    .X(_01971_));
 sg13g2_nor2_2 _07267_ (.A(_01910_),
    .B(net335),
    .Y(_01972_));
 sg13g2_o21ai_1 _07268_ (.B1(_01945_),
    .Y(_01973_),
    .A1(_01922_),
    .A2(_01972_));
 sg13g2_inv_1 _07269_ (.Y(_01974_),
    .A(net38));
 sg13g2_and2_1 _07270_ (.A(net468),
    .B(_01767_),
    .X(_01975_));
 sg13g2_buf_2 _07271_ (.A(_01975_),
    .X(_01976_));
 sg13g2_nand2_1 _07272_ (.Y(_01977_),
    .A(_01976_),
    .B(_01940_));
 sg13g2_buf_2 _07273_ (.A(_01977_),
    .X(_01978_));
 sg13g2_nor3_1 _07274_ (.A(net346),
    .B(_01974_),
    .C(_01978_),
    .Y(_01979_));
 sg13g2_a21o_1 _07275_ (.A2(_01973_),
    .A1(net346),
    .B1(_01979_),
    .X(_00431_));
 sg13g2_nand3_1 _07276_ (.B(net38),
    .C(_01972_),
    .A(net346),
    .Y(_01980_));
 sg13g2_a21oi_1 _07277_ (.A1(net346),
    .A2(_01972_),
    .Y(_01981_),
    .B1(_01922_));
 sg13g2_o21ai_1 _07278_ (.B1(net400),
    .Y(_01982_),
    .A1(_01906_),
    .A2(_01981_));
 sg13g2_o21ai_1 _07279_ (.B1(_01982_),
    .Y(_00432_),
    .A1(net400),
    .A2(_01980_));
 sg13g2_nand2_1 _07280_ (.Y(_01983_),
    .A(net474),
    .B(_01753_));
 sg13g2_buf_1 _07281_ (.A(_01983_),
    .X(_01984_));
 sg13g2_nor2_1 _07282_ (.A(_01978_),
    .B(net386),
    .Y(_01985_));
 sg13g2_nand2_1 _07283_ (.Y(_01986_),
    .A(net38),
    .B(_01985_));
 sg13g2_nor2_1 _07284_ (.A(_01922_),
    .B(_01985_),
    .Y(_01987_));
 sg13g2_o21ai_1 _07285_ (.B1(_01760_),
    .Y(_01988_),
    .A1(_01906_),
    .A2(_01987_));
 sg13g2_o21ai_1 _07286_ (.B1(_01988_),
    .Y(_00433_),
    .A1(_01760_),
    .A2(_01986_));
 sg13g2_and2_1 _07287_ (.A(net475),
    .B(_01985_),
    .X(_01989_));
 sg13g2_buf_1 _07288_ (.A(_01989_),
    .X(_01990_));
 sg13g2_nand2_1 _07289_ (.Y(_01991_),
    .A(net38),
    .B(_01990_));
 sg13g2_nor2_1 _07290_ (.A(_01922_),
    .B(_01990_),
    .Y(_01992_));
 sg13g2_o21ai_1 _07291_ (.B1(net445),
    .Y(_01993_),
    .A1(_01906_),
    .A2(_01992_));
 sg13g2_o21ai_1 _07292_ (.B1(_01993_),
    .Y(_00434_),
    .A1(net445),
    .A2(_01991_));
 sg13g2_nand3_1 _07293_ (.B(net38),
    .C(_01990_),
    .A(net445),
    .Y(_01994_));
 sg13g2_a21oi_1 _07294_ (.A1(_01759_),
    .A2(_01990_),
    .Y(_01995_),
    .B1(_01974_));
 sg13g2_o21ai_1 _07295_ (.B1(_01757_),
    .Y(_01996_),
    .A1(_01906_),
    .A2(_01995_));
 sg13g2_o21ai_1 _07296_ (.B1(_01996_),
    .Y(_00435_),
    .A1(_01757_),
    .A2(_01994_));
 sg13g2_nand2_1 _07297_ (.Y(_01997_),
    .A(_01757_),
    .B(net445));
 sg13g2_nand2b_1 _07298_ (.Y(_01998_),
    .B(_01990_),
    .A_N(_01997_));
 sg13g2_a21o_1 _07299_ (.A2(_01998_),
    .A1(_01924_),
    .B1(_01906_),
    .X(_01999_));
 sg13g2_nor3_1 _07300_ (.A(_01752_),
    .B(_01997_),
    .C(_01991_),
    .Y(_02000_));
 sg13g2_a21o_1 _07301_ (.A2(_01999_),
    .A1(_01752_),
    .B1(_02000_),
    .X(_00436_));
 sg13g2_buf_1 _07302_ (.A(\welcome_screen_inst.welcome_counter[0] ),
    .X(_02001_));
 sg13g2_buf_1 _07303_ (.A(\lfsr_inst.lfsr[28] ),
    .X(_02002_));
 sg13g2_buf_1 _07304_ (.A(_02002_),
    .X(_02003_));
 sg13g2_buf_1 _07305_ (.A(\lfsr_inst.lfsr[29] ),
    .X(_02004_));
 sg13g2_mux4_1 _07306_ (.S0(net430),
    .A0(\welcome_screen_grid[0] ),
    .A1(\welcome_screen_grid[4] ),
    .A2(\welcome_screen_grid[11] ),
    .A3(\welcome_screen_grid[12] ),
    .S1(net466),
    .X(_02005_));
 sg13g2_mux4_1 _07307_ (.S0(net430),
    .A0(\welcome_screen_grid[16] ),
    .A1(\welcome_screen_grid[20] ),
    .A2(\welcome_screen_grid[24] ),
    .A3(\welcome_screen_grid[28] ),
    .S1(net466),
    .X(_02006_));
 sg13g2_mux4_1 _07308_ (.S0(_02002_),
    .A0(\welcome_screen_grid[32] ),
    .A1(\welcome_screen_grid[36] ),
    .A2(\welcome_screen_grid[40] ),
    .A3(\welcome_screen_grid[44] ),
    .S1(\lfsr_inst.lfsr[29] ),
    .X(_02007_));
 sg13g2_mux4_1 _07309_ (.S0(net430),
    .A0(\welcome_screen_grid[48] ),
    .A1(\welcome_screen_grid[52] ),
    .A2(\welcome_screen_grid[56] ),
    .A3(\welcome_screen_grid[60] ),
    .S1(net466),
    .X(_02008_));
 sg13g2_buf_1 _07310_ (.A(\lfsr_inst.lfsr[30] ),
    .X(_02009_));
 sg13g2_buf_1 _07311_ (.A(\lfsr_inst.lfsr[31] ),
    .X(_02010_));
 sg13g2_mux4_1 _07312_ (.S0(net465),
    .A0(_02005_),
    .A1(_02006_),
    .A2(_02007_),
    .A3(_02008_),
    .S1(net464),
    .X(_02011_));
 sg13g2_buf_1 _07313_ (.A(\welcome_screen_inst.welcome_counter[1] ),
    .X(_02012_));
 sg13g2_buf_1 _07314_ (.A(\welcome_screen_inst.welcome_counter[3] ),
    .X(_02013_));
 sg13g2_buf_1 _07315_ (.A(\welcome_screen_inst.welcome_counter[2] ),
    .X(_02014_));
 sg13g2_nand4_1 _07316_ (.B(_02013_),
    .C(_02014_),
    .A(_02012_),
    .Y(_02015_),
    .D(\welcome_screen_inst.welcome_counter[4] ));
 sg13g2_nor3_2 _07317_ (.A(_02001_),
    .B(_02011_),
    .C(_02015_),
    .Y(_02016_));
 sg13g2_nand2_1 _07318_ (.Y(_02017_),
    .A(net478),
    .B(_02016_));
 sg13g2_buf_1 _07319_ (.A(_02017_),
    .X(_02018_));
 sg13g2_buf_1 _07320_ (.A(_02018_),
    .X(_02019_));
 sg13g2_buf_1 _07321_ (.A(_02018_),
    .X(_02020_));
 sg13g2_nand2b_1 _07322_ (.Y(_02021_),
    .B(net466),
    .A_N(net430));
 sg13g2_nor4_1 _07323_ (.A(net465),
    .B(net464),
    .C(_02020_),
    .D(_02021_),
    .Y(_02022_));
 sg13g2_a21o_1 _07324_ (.A2(net64),
    .A1(\welcome_screen_grid[11] ),
    .B1(_02022_),
    .X(_00438_));
 sg13g2_nand2_1 _07325_ (.Y(_02023_),
    .A(net430),
    .B(net466));
 sg13g2_nor4_1 _07326_ (.A(net465),
    .B(net464),
    .C(net63),
    .D(_02023_),
    .Y(_02024_));
 sg13g2_a21o_1 _07327_ (.A2(net64),
    .A1(\welcome_screen_grid[12] ),
    .B1(_02024_),
    .X(_00439_));
 sg13g2_nand2b_1 _07328_ (.Y(_02025_),
    .B(net465),
    .A_N(net464));
 sg13g2_nor4_1 _07329_ (.A(net430),
    .B(net466),
    .C(net63),
    .D(_02025_),
    .Y(_02026_));
 sg13g2_a21o_1 _07330_ (.A2(net64),
    .A1(\welcome_screen_grid[16] ),
    .B1(_02026_),
    .X(_00440_));
 sg13g2_buf_1 _07331_ (.A(_02018_),
    .X(_02027_));
 sg13g2_nand2b_1 _07332_ (.Y(_02028_),
    .B(net430),
    .A_N(_02004_));
 sg13g2_nor3_1 _07333_ (.A(net62),
    .B(_02025_),
    .C(_02028_),
    .Y(_02029_));
 sg13g2_a21o_1 _07334_ (.A2(net64),
    .A1(\welcome_screen_grid[20] ),
    .B1(_02029_),
    .X(_00441_));
 sg13g2_nor3_1 _07335_ (.A(net62),
    .B(_02021_),
    .C(_02025_),
    .Y(_02030_));
 sg13g2_a21o_1 _07336_ (.A2(net64),
    .A1(\welcome_screen_grid[24] ),
    .B1(_02030_),
    .X(_00442_));
 sg13g2_nor3_1 _07337_ (.A(net62),
    .B(_02023_),
    .C(_02025_),
    .Y(_02031_));
 sg13g2_a21o_1 _07338_ (.A2(net64),
    .A1(\welcome_screen_grid[28] ),
    .B1(_02031_),
    .X(_00443_));
 sg13g2_nand2b_1 _07339_ (.Y(_02032_),
    .B(net464),
    .A_N(net465));
 sg13g2_nor2_1 _07340_ (.A(_02003_),
    .B(net466),
    .Y(_02033_));
 sg13g2_nand2_1 _07341_ (.Y(_02034_),
    .A(_00070_),
    .B(_02033_));
 sg13g2_nor3_1 _07342_ (.A(net62),
    .B(_02032_),
    .C(_02034_),
    .Y(_02035_));
 sg13g2_a21o_1 _07343_ (.A2(_02019_),
    .A1(\welcome_screen_grid[32] ),
    .B1(_02035_),
    .X(_00444_));
 sg13g2_xnor2_1 _07344_ (.Y(_02036_),
    .A(net464),
    .B(_00070_));
 sg13g2_nor4_1 _07345_ (.A(_02009_),
    .B(_02018_),
    .C(_02028_),
    .D(_02036_),
    .Y(_02037_));
 sg13g2_a21o_1 _07346_ (.A2(_02019_),
    .A1(\welcome_screen_grid[36] ),
    .B1(_02037_),
    .X(_00445_));
 sg13g2_nor4_1 _07347_ (.A(net465),
    .B(net464),
    .C(net63),
    .D(_02034_),
    .Y(_02038_));
 sg13g2_a21o_1 _07348_ (.A2(net64),
    .A1(\welcome_screen_grid[0] ),
    .B1(_02038_),
    .X(_00446_));
 sg13g2_nor3_1 _07349_ (.A(net63),
    .B(_02021_),
    .C(_02032_),
    .Y(_02039_));
 sg13g2_a21o_1 _07350_ (.A2(net64),
    .A1(\welcome_screen_grid[40] ),
    .B1(_02039_),
    .X(_00447_));
 sg13g2_nor3_1 _07351_ (.A(net63),
    .B(_02023_),
    .C(_02032_),
    .Y(_02040_));
 sg13g2_a21o_1 _07352_ (.A2(net62),
    .A1(\welcome_screen_grid[44] ),
    .B1(_02040_),
    .X(_00448_));
 sg13g2_nand2_1 _07353_ (.Y(_02041_),
    .A(net465),
    .B(net464));
 sg13g2_nor4_1 _07354_ (.A(net430),
    .B(_02004_),
    .C(net63),
    .D(_02041_),
    .Y(_02042_));
 sg13g2_a21o_1 _07355_ (.A2(_02027_),
    .A1(\welcome_screen_grid[48] ),
    .B1(_02042_),
    .X(_00449_));
 sg13g2_nor3_1 _07356_ (.A(net63),
    .B(_02028_),
    .C(_02041_),
    .Y(_02043_));
 sg13g2_a21o_1 _07357_ (.A2(_02027_),
    .A1(\welcome_screen_grid[52] ),
    .B1(_02043_),
    .X(_00450_));
 sg13g2_nor3_1 _07358_ (.A(net63),
    .B(_02021_),
    .C(_02041_),
    .Y(_02044_));
 sg13g2_a21o_1 _07359_ (.A2(net62),
    .A1(\welcome_screen_grid[56] ),
    .B1(_02044_),
    .X(_00451_));
 sg13g2_nor3_1 _07360_ (.A(_02020_),
    .B(_02023_),
    .C(_02041_),
    .Y(_02045_));
 sg13g2_a21o_1 _07361_ (.A2(net62),
    .A1(\welcome_screen_grid[60] ),
    .B1(_02045_),
    .X(_00452_));
 sg13g2_nor2_1 _07362_ (.A(_02009_),
    .B(_02028_),
    .Y(_02046_));
 sg13g2_and4_1 _07363_ (.A(net407),
    .B(_02016_),
    .C(_02036_),
    .D(_02046_),
    .X(_02047_));
 sg13g2_a21o_1 _07364_ (.A2(net62),
    .A1(\welcome_screen_grid[4] ),
    .B1(_02047_),
    .X(_00453_));
 sg13g2_inv_1 _07365_ (.Y(_02048_),
    .A(_00166_));
 sg13g2_xor2_1 _07366_ (.B(\btn_down_debounce.button_sync_1 ),
    .A(_05073_),
    .X(_02049_));
 sg13g2_buf_1 _07367_ (.A(\btn_down_debounce.debounce_counter[0] ),
    .X(_02050_));
 sg13g2_inv_1 _07368_ (.Y(_02051_),
    .A(\btn_down_debounce.debounce_counter[7] ));
 sg13g2_nor4_1 _07369_ (.A(_02050_),
    .B(\btn_down_debounce.debounce_counter[3] ),
    .C(\btn_down_debounce.debounce_counter[2] ),
    .D(_02051_),
    .Y(_02052_));
 sg13g2_buf_1 _07370_ (.A(\btn_down_debounce.debounce_counter[1] ),
    .X(_02053_));
 sg13g2_buf_1 _07371_ (.A(\btn_down_debounce.debounce_counter[5] ),
    .X(_02054_));
 sg13g2_buf_1 _07372_ (.A(\btn_down_debounce.debounce_counter[4] ),
    .X(_02055_));
 sg13g2_inv_1 _07373_ (.Y(_02056_),
    .A(_02055_));
 sg13g2_nor4_1 _07374_ (.A(_02053_),
    .B(_02054_),
    .C(_02056_),
    .D(\btn_down_debounce.debounce_counter[6] ),
    .Y(_02057_));
 sg13g2_buf_1 _07375_ (.A(\btn_down_debounce.debounce_counter[14] ),
    .X(_02058_));
 sg13g2_nand3_1 _07376_ (.B(_02058_),
    .C(\btn_down_debounce.debounce_counter[16] ),
    .A(\btn_down_debounce.debounce_counter[15] ),
    .Y(_02059_));
 sg13g2_inv_1 _07377_ (.Y(_02060_),
    .A(\btn_down_debounce.debounce_counter[13] ));
 sg13g2_buf_1 _07378_ (.A(\btn_down_debounce.debounce_counter[8] ),
    .X(_02061_));
 sg13g2_buf_1 _07379_ (.A(\btn_down_debounce.debounce_counter[11] ),
    .X(_02062_));
 sg13g2_nor4_1 _07380_ (.A(\btn_down_debounce.debounce_counter[9] ),
    .B(_02061_),
    .C(_02062_),
    .D(\btn_down_debounce.debounce_counter[10] ),
    .Y(_02063_));
 sg13g2_nand4_1 _07381_ (.B(\btn_down_debounce.debounce_counter[12] ),
    .C(\btn_down_debounce.debounce_counter[17] ),
    .A(_02060_),
    .Y(_02064_),
    .D(_02063_));
 sg13g2_nor2_1 _07382_ (.A(_02059_),
    .B(_02064_),
    .Y(_02065_));
 sg13g2_nand3_1 _07383_ (.B(_02057_),
    .C(_02065_),
    .A(_02052_),
    .Y(_02066_));
 sg13g2_nand3_1 _07384_ (.B(_02049_),
    .C(_02066_),
    .A(_00918_),
    .Y(_02067_));
 sg13g2_buf_1 _07385_ (.A(_02067_),
    .X(_02068_));
 sg13g2_buf_1 _07386_ (.A(net86),
    .X(_02069_));
 sg13g2_nor2_1 _07387_ (.A(_02048_),
    .B(net61),
    .Y(_00179_));
 sg13g2_inv_1 _07388_ (.Y(_02070_),
    .A(\btn_down_debounce.debounce_counter[10] ));
 sg13g2_inv_1 _07389_ (.Y(_02071_),
    .A(\btn_down_debounce.debounce_counter[3] ));
 sg13g2_nand3_1 _07390_ (.B(_02050_),
    .C(\btn_down_debounce.debounce_counter[2] ),
    .A(_02053_),
    .Y(_02072_));
 sg13g2_nor2_2 _07391_ (.A(_02071_),
    .B(_02072_),
    .Y(_02073_));
 sg13g2_nand4_1 _07392_ (.B(_02055_),
    .C(\btn_down_debounce.debounce_counter[6] ),
    .A(_02054_),
    .Y(_02074_),
    .D(_02073_));
 sg13g2_nor2_1 _07393_ (.A(_02051_),
    .B(_02074_),
    .Y(_02075_));
 sg13g2_nand3_1 _07394_ (.B(_02061_),
    .C(_02075_),
    .A(\btn_down_debounce.debounce_counter[9] ),
    .Y(_02076_));
 sg13g2_xnor2_1 _07395_ (.Y(_02077_),
    .A(_02070_),
    .B(_02076_));
 sg13g2_nor2_1 _07396_ (.A(net61),
    .B(_02077_),
    .Y(_00180_));
 sg13g2_nor2_1 _07397_ (.A(_02070_),
    .B(_02076_),
    .Y(_02078_));
 sg13g2_xnor2_1 _07398_ (.Y(_02079_),
    .A(_02062_),
    .B(_02078_));
 sg13g2_nor2_1 _07399_ (.A(net61),
    .B(_02079_),
    .Y(_00181_));
 sg13g2_nand2_1 _07400_ (.Y(_02080_),
    .A(_02062_),
    .B(_02078_));
 sg13g2_xor2_1 _07401_ (.B(_02080_),
    .A(\btn_down_debounce.debounce_counter[12] ),
    .X(_02081_));
 sg13g2_nor2_1 _07402_ (.A(net61),
    .B(_02081_),
    .Y(_00182_));
 sg13g2_nand3_1 _07403_ (.B(\btn_down_debounce.debounce_counter[12] ),
    .C(_02078_),
    .A(_02062_),
    .Y(_02082_));
 sg13g2_xnor2_1 _07404_ (.Y(_02083_),
    .A(_02060_),
    .B(_02082_));
 sg13g2_nor2_1 _07405_ (.A(net61),
    .B(_02083_),
    .Y(_00183_));
 sg13g2_nor2_2 _07406_ (.A(_02060_),
    .B(_02082_),
    .Y(_02084_));
 sg13g2_xnor2_1 _07407_ (.Y(_02085_),
    .A(_02058_),
    .B(_02084_));
 sg13g2_nor2_1 _07408_ (.A(net61),
    .B(_02085_),
    .Y(_00184_));
 sg13g2_nand2_1 _07409_ (.Y(_02086_),
    .A(_02058_),
    .B(_02084_));
 sg13g2_xor2_1 _07410_ (.B(_02086_),
    .A(\btn_down_debounce.debounce_counter[15] ),
    .X(_02087_));
 sg13g2_nor2_1 _07411_ (.A(net61),
    .B(_02087_),
    .Y(_00185_));
 sg13g2_nand3_1 _07412_ (.B(_02058_),
    .C(_02084_),
    .A(\btn_down_debounce.debounce_counter[15] ),
    .Y(_02088_));
 sg13g2_xor2_1 _07413_ (.B(_02088_),
    .A(\btn_down_debounce.debounce_counter[16] ),
    .X(_02089_));
 sg13g2_nor2_1 _07414_ (.A(_02069_),
    .B(_02089_),
    .Y(_00186_));
 sg13g2_nand2b_1 _07415_ (.Y(_02090_),
    .B(_02084_),
    .A_N(_02059_));
 sg13g2_xor2_1 _07416_ (.B(_02090_),
    .A(\btn_down_debounce.debounce_counter[17] ),
    .X(_02091_));
 sg13g2_nor2_1 _07417_ (.A(_02069_),
    .B(_02091_),
    .Y(_00187_));
 sg13g2_xnor2_1 _07418_ (.Y(_02092_),
    .A(_02053_),
    .B(_02050_));
 sg13g2_nor2_1 _07419_ (.A(net61),
    .B(_02092_),
    .Y(_00188_));
 sg13g2_nand2_1 _07420_ (.Y(_02093_),
    .A(_02053_),
    .B(_02050_));
 sg13g2_xor2_1 _07421_ (.B(_02093_),
    .A(\btn_down_debounce.debounce_counter[2] ),
    .X(_02094_));
 sg13g2_nor2_1 _07422_ (.A(net86),
    .B(_02094_),
    .Y(_00189_));
 sg13g2_xnor2_1 _07423_ (.Y(_02095_),
    .A(_02071_),
    .B(_02072_));
 sg13g2_nor2_1 _07424_ (.A(net86),
    .B(_02095_),
    .Y(_00190_));
 sg13g2_xnor2_1 _07425_ (.Y(_02096_),
    .A(_02055_),
    .B(_02073_));
 sg13g2_nor2_1 _07426_ (.A(net86),
    .B(_02096_),
    .Y(_00191_));
 sg13g2_nand2_1 _07427_ (.Y(_02097_),
    .A(_02055_),
    .B(_02073_));
 sg13g2_xor2_1 _07428_ (.B(_02097_),
    .A(_02054_),
    .X(_02098_));
 sg13g2_nor2_1 _07429_ (.A(net86),
    .B(_02098_),
    .Y(_00192_));
 sg13g2_nand3_1 _07430_ (.B(_02055_),
    .C(_02073_),
    .A(_02054_),
    .Y(_02099_));
 sg13g2_xor2_1 _07431_ (.B(_02099_),
    .A(\btn_down_debounce.debounce_counter[6] ),
    .X(_02100_));
 sg13g2_nor2_1 _07432_ (.A(net86),
    .B(_02100_),
    .Y(_00193_));
 sg13g2_xnor2_1 _07433_ (.Y(_02101_),
    .A(_02051_),
    .B(_02074_));
 sg13g2_nor2_1 _07434_ (.A(_02068_),
    .B(_02101_),
    .Y(_00194_));
 sg13g2_xnor2_1 _07435_ (.Y(_02102_),
    .A(_02061_),
    .B(_02075_));
 sg13g2_nor2_1 _07436_ (.A(net86),
    .B(_02102_),
    .Y(_00195_));
 sg13g2_nand2_1 _07437_ (.Y(_02103_),
    .A(_02061_),
    .B(_02075_));
 sg13g2_xor2_1 _07438_ (.B(_02103_),
    .A(\btn_down_debounce.debounce_counter[9] ),
    .X(_02104_));
 sg13g2_nor2_1 _07439_ (.A(net86),
    .B(_02104_),
    .Y(_00196_));
 sg13g2_inv_1 _07440_ (.Y(_02105_),
    .A(_00167_));
 sg13g2_inv_1 _07441_ (.Y(_02106_),
    .A(\btn_left_debounce.debounce_counter[6] ));
 sg13g2_buf_1 _07442_ (.A(\btn_left_debounce.debounce_counter[4] ),
    .X(_02107_));
 sg13g2_nor2b_1 _07443_ (.A(\btn_left_debounce.debounce_counter[5] ),
    .B_N(_02107_),
    .Y(_02108_));
 sg13g2_buf_1 _07444_ (.A(\btn_left_debounce.debounce_counter[1] ),
    .X(_02109_));
 sg13g2_buf_1 _07445_ (.A(\btn_left_debounce.debounce_counter[8] ),
    .X(_02110_));
 sg13g2_buf_1 _07446_ (.A(\btn_left_debounce.debounce_counter[11] ),
    .X(_02111_));
 sg13g2_nor4_1 _07447_ (.A(_02109_),
    .B(_02110_),
    .C(_02111_),
    .D(\btn_left_debounce.debounce_counter[10] ),
    .Y(_02112_));
 sg13g2_nand4_1 _07448_ (.B(\btn_left_debounce.debounce_counter[7] ),
    .C(_02108_),
    .A(_02106_),
    .Y(_02113_),
    .D(_02112_));
 sg13g2_inv_1 _07449_ (.Y(_02114_),
    .A(\btn_left_debounce.debounce_counter[13] ));
 sg13g2_nand4_1 _07450_ (.B(\btn_left_debounce.debounce_counter[12] ),
    .C(\btn_left_debounce.debounce_counter[14] ),
    .A(_02114_),
    .Y(_02115_),
    .D(\btn_left_debounce.debounce_counter[17] ));
 sg13g2_buf_1 _07451_ (.A(\btn_left_debounce.debounce_counter[15] ),
    .X(_02116_));
 sg13g2_buf_1 _07452_ (.A(\btn_left_debounce.debounce_counter[0] ),
    .X(_02117_));
 sg13g2_nor4_1 _07453_ (.A(_02117_),
    .B(\btn_left_debounce.debounce_counter[3] ),
    .C(\btn_left_debounce.debounce_counter[2] ),
    .D(\btn_left_debounce.debounce_counter[9] ),
    .Y(_02118_));
 sg13g2_nand3_1 _07454_ (.B(\btn_left_debounce.debounce_counter[16] ),
    .C(_02118_),
    .A(_02116_),
    .Y(_02119_));
 sg13g2_nor3_2 _07455_ (.A(_02113_),
    .B(_02115_),
    .C(_02119_),
    .Y(_02120_));
 sg13g2_xor2_1 _07456_ (.B(\btn_left_debounce.button_sync_1 ),
    .A(_05066_),
    .X(_02121_));
 sg13g2_nand3b_1 _07457_ (.B(_02121_),
    .C(_00918_),
    .Y(_02122_),
    .A_N(_02120_));
 sg13g2_buf_1 _07458_ (.A(_02122_),
    .X(_02123_));
 sg13g2_buf_1 _07459_ (.A(net148),
    .X(_02124_));
 sg13g2_nor2_1 _07460_ (.A(_02105_),
    .B(net85),
    .Y(_00200_));
 sg13g2_inv_1 _07461_ (.Y(_02125_),
    .A(\btn_left_debounce.debounce_counter[10] ));
 sg13g2_inv_1 _07462_ (.Y(_02126_),
    .A(\btn_left_debounce.debounce_counter[7] ));
 sg13g2_inv_1 _07463_ (.Y(_02127_),
    .A(\btn_left_debounce.debounce_counter[3] ));
 sg13g2_nand3_1 _07464_ (.B(_02117_),
    .C(\btn_left_debounce.debounce_counter[2] ),
    .A(_02109_),
    .Y(_02128_));
 sg13g2_nor2_1 _07465_ (.A(_02127_),
    .B(_02128_),
    .Y(_02129_));
 sg13g2_nand3_1 _07466_ (.B(_02107_),
    .C(_02129_),
    .A(\btn_left_debounce.debounce_counter[5] ),
    .Y(_02130_));
 sg13g2_or2_1 _07467_ (.X(_02131_),
    .B(_02130_),
    .A(_02106_));
 sg13g2_nor2_1 _07468_ (.A(_02126_),
    .B(_02131_),
    .Y(_02132_));
 sg13g2_nand3_1 _07469_ (.B(_02110_),
    .C(_02132_),
    .A(\btn_left_debounce.debounce_counter[9] ),
    .Y(_02133_));
 sg13g2_xnor2_1 _07470_ (.Y(_02134_),
    .A(_02125_),
    .B(_02133_));
 sg13g2_nor2_1 _07471_ (.A(net85),
    .B(_02134_),
    .Y(_00201_));
 sg13g2_nor2_1 _07472_ (.A(_02125_),
    .B(_02133_),
    .Y(_02135_));
 sg13g2_xnor2_1 _07473_ (.Y(_02136_),
    .A(_02111_),
    .B(_02135_));
 sg13g2_nor2_1 _07474_ (.A(net85),
    .B(_02136_),
    .Y(_00202_));
 sg13g2_nand2_1 _07475_ (.Y(_02137_),
    .A(_02111_),
    .B(_02135_));
 sg13g2_xor2_1 _07476_ (.B(_02137_),
    .A(\btn_left_debounce.debounce_counter[12] ),
    .X(_02138_));
 sg13g2_nor2_1 _07477_ (.A(net85),
    .B(_02138_),
    .Y(_00203_));
 sg13g2_nand3_1 _07478_ (.B(\btn_left_debounce.debounce_counter[12] ),
    .C(_02135_),
    .A(_02111_),
    .Y(_02139_));
 sg13g2_xnor2_1 _07479_ (.Y(_02140_),
    .A(_02114_),
    .B(_02139_));
 sg13g2_nor2_1 _07480_ (.A(net85),
    .B(_02140_),
    .Y(_00204_));
 sg13g2_nor2_1 _07481_ (.A(_02114_),
    .B(_02139_),
    .Y(_02141_));
 sg13g2_xnor2_1 _07482_ (.Y(_02142_),
    .A(\btn_left_debounce.debounce_counter[14] ),
    .B(_02141_));
 sg13g2_nor2_1 _07483_ (.A(net85),
    .B(_02142_),
    .Y(_00205_));
 sg13g2_and2_1 _07484_ (.A(\btn_left_debounce.debounce_counter[14] ),
    .B(_02141_),
    .X(_02143_));
 sg13g2_buf_1 _07485_ (.A(_02143_),
    .X(_02144_));
 sg13g2_xnor2_1 _07486_ (.Y(_02145_),
    .A(_02116_),
    .B(_02144_));
 sg13g2_nor2_1 _07487_ (.A(_02124_),
    .B(_02145_),
    .Y(_00206_));
 sg13g2_nand2_1 _07488_ (.Y(_02146_),
    .A(_02116_),
    .B(_02144_));
 sg13g2_xor2_1 _07489_ (.B(_02146_),
    .A(\btn_left_debounce.debounce_counter[16] ),
    .X(_02147_));
 sg13g2_nor2_1 _07490_ (.A(net85),
    .B(_02147_),
    .Y(_00207_));
 sg13g2_nand3_1 _07491_ (.B(\btn_left_debounce.debounce_counter[16] ),
    .C(_02144_),
    .A(_02116_),
    .Y(_02148_));
 sg13g2_xor2_1 _07492_ (.B(_02148_),
    .A(\btn_left_debounce.debounce_counter[17] ),
    .X(_02149_));
 sg13g2_nor2_1 _07493_ (.A(_02124_),
    .B(_02149_),
    .Y(_00208_));
 sg13g2_xnor2_1 _07494_ (.Y(_02150_),
    .A(_02109_),
    .B(_02117_));
 sg13g2_nor2_1 _07495_ (.A(net85),
    .B(_02150_),
    .Y(_00209_));
 sg13g2_nand2_1 _07496_ (.Y(_02151_),
    .A(_02109_),
    .B(_02117_));
 sg13g2_xor2_1 _07497_ (.B(_02151_),
    .A(\btn_left_debounce.debounce_counter[2] ),
    .X(_02152_));
 sg13g2_nor2_1 _07498_ (.A(net148),
    .B(_02152_),
    .Y(_00210_));
 sg13g2_xnor2_1 _07499_ (.Y(_02153_),
    .A(_02127_),
    .B(_02128_));
 sg13g2_nor2_1 _07500_ (.A(net148),
    .B(_02153_),
    .Y(_00211_));
 sg13g2_xnor2_1 _07501_ (.Y(_02154_),
    .A(_02107_),
    .B(_02129_));
 sg13g2_nor2_1 _07502_ (.A(net148),
    .B(_02154_),
    .Y(_00212_));
 sg13g2_nand2_1 _07503_ (.Y(_02155_),
    .A(_02107_),
    .B(_02129_));
 sg13g2_xor2_1 _07504_ (.B(_02155_),
    .A(\btn_left_debounce.debounce_counter[5] ),
    .X(_02156_));
 sg13g2_nor2_1 _07505_ (.A(net148),
    .B(_02156_),
    .Y(_00213_));
 sg13g2_xnor2_1 _07506_ (.Y(_02157_),
    .A(_02106_),
    .B(_02130_));
 sg13g2_nor2_1 _07507_ (.A(net148),
    .B(_02157_),
    .Y(_00214_));
 sg13g2_xnor2_1 _07508_ (.Y(_02158_),
    .A(_02126_),
    .B(_02131_));
 sg13g2_nor2_1 _07509_ (.A(net148),
    .B(_02158_),
    .Y(_00215_));
 sg13g2_xnor2_1 _07510_ (.Y(_02159_),
    .A(_02110_),
    .B(_02132_));
 sg13g2_nor2_1 _07511_ (.A(net148),
    .B(_02159_),
    .Y(_00216_));
 sg13g2_nand2_1 _07512_ (.Y(_02160_),
    .A(_02110_),
    .B(_02132_));
 sg13g2_xor2_1 _07513_ (.B(_02160_),
    .A(\btn_left_debounce.debounce_counter[9] ),
    .X(_02161_));
 sg13g2_nor2_1 _07514_ (.A(_02123_),
    .B(_02161_),
    .Y(_00217_));
 sg13g2_inv_1 _07515_ (.Y(_02162_),
    .A(_00168_));
 sg13g2_inv_1 _07516_ (.Y(_02163_),
    .A(\btn_right_debounce.debounce_counter[6] ));
 sg13g2_buf_1 _07517_ (.A(\btn_right_debounce.debounce_counter[4] ),
    .X(_02164_));
 sg13g2_nor2b_1 _07518_ (.A(\btn_right_debounce.debounce_counter[5] ),
    .B_N(_02164_),
    .Y(_02165_));
 sg13g2_buf_1 _07519_ (.A(\btn_right_debounce.debounce_counter[1] ),
    .X(_02166_));
 sg13g2_buf_1 _07520_ (.A(\btn_right_debounce.debounce_counter[8] ),
    .X(_02167_));
 sg13g2_buf_1 _07521_ (.A(\btn_right_debounce.debounce_counter[11] ),
    .X(_02168_));
 sg13g2_nor4_1 _07522_ (.A(_02166_),
    .B(_02167_),
    .C(_02168_),
    .D(\btn_right_debounce.debounce_counter[10] ),
    .Y(_02169_));
 sg13g2_nand4_1 _07523_ (.B(\btn_right_debounce.debounce_counter[7] ),
    .C(_02165_),
    .A(_02163_),
    .Y(_02170_),
    .D(_02169_));
 sg13g2_inv_1 _07524_ (.Y(_02171_),
    .A(\btn_right_debounce.debounce_counter[13] ));
 sg13g2_nand4_1 _07525_ (.B(\btn_right_debounce.debounce_counter[12] ),
    .C(\btn_right_debounce.debounce_counter[14] ),
    .A(_02171_),
    .Y(_02172_),
    .D(\btn_right_debounce.debounce_counter[17] ));
 sg13g2_buf_1 _07526_ (.A(\btn_right_debounce.debounce_counter[15] ),
    .X(_02173_));
 sg13g2_buf_1 _07527_ (.A(\btn_right_debounce.debounce_counter[0] ),
    .X(_02174_));
 sg13g2_nor4_1 _07528_ (.A(_02174_),
    .B(\btn_right_debounce.debounce_counter[3] ),
    .C(\btn_right_debounce.debounce_counter[2] ),
    .D(\btn_right_debounce.debounce_counter[9] ),
    .Y(_02175_));
 sg13g2_nand3_1 _07529_ (.B(\btn_right_debounce.debounce_counter[16] ),
    .C(_02175_),
    .A(_02173_),
    .Y(_02176_));
 sg13g2_nor3_2 _07530_ (.A(_02170_),
    .B(_02172_),
    .C(_02176_),
    .Y(_02177_));
 sg13g2_xor2_1 _07531_ (.B(\btn_right_debounce.button_sync_1 ),
    .A(_05065_),
    .X(_02178_));
 sg13g2_nand3b_1 _07532_ (.B(_02178_),
    .C(net478),
    .Y(_02179_),
    .A_N(_02177_));
 sg13g2_buf_1 _07533_ (.A(_02179_),
    .X(_02180_));
 sg13g2_buf_1 _07534_ (.A(net147),
    .X(_02181_));
 sg13g2_nor2_1 _07535_ (.A(_02162_),
    .B(net84),
    .Y(_00221_));
 sg13g2_inv_1 _07536_ (.Y(_02182_),
    .A(\btn_right_debounce.debounce_counter[10] ));
 sg13g2_inv_1 _07537_ (.Y(_02183_),
    .A(\btn_right_debounce.debounce_counter[7] ));
 sg13g2_inv_1 _07538_ (.Y(_02184_),
    .A(\btn_right_debounce.debounce_counter[3] ));
 sg13g2_nand3_1 _07539_ (.B(_02174_),
    .C(\btn_right_debounce.debounce_counter[2] ),
    .A(_02166_),
    .Y(_02185_));
 sg13g2_nor2_1 _07540_ (.A(_02184_),
    .B(_02185_),
    .Y(_02186_));
 sg13g2_nand3_1 _07541_ (.B(_02164_),
    .C(_02186_),
    .A(\btn_right_debounce.debounce_counter[5] ),
    .Y(_02187_));
 sg13g2_or2_1 _07542_ (.X(_02188_),
    .B(_02187_),
    .A(_02163_));
 sg13g2_nor2_1 _07543_ (.A(_02183_),
    .B(_02188_),
    .Y(_02189_));
 sg13g2_nand3_1 _07544_ (.B(_02167_),
    .C(_02189_),
    .A(\btn_right_debounce.debounce_counter[9] ),
    .Y(_02190_));
 sg13g2_xnor2_1 _07545_ (.Y(_02191_),
    .A(_02182_),
    .B(_02190_));
 sg13g2_nor2_1 _07546_ (.A(net84),
    .B(_02191_),
    .Y(_00222_));
 sg13g2_nor2_1 _07547_ (.A(_02182_),
    .B(_02190_),
    .Y(_02192_));
 sg13g2_xnor2_1 _07548_ (.Y(_02193_),
    .A(_02168_),
    .B(_02192_));
 sg13g2_nor2_1 _07549_ (.A(net84),
    .B(_02193_),
    .Y(_00223_));
 sg13g2_nand2_1 _07550_ (.Y(_02194_),
    .A(_02168_),
    .B(_02192_));
 sg13g2_xor2_1 _07551_ (.B(_02194_),
    .A(\btn_right_debounce.debounce_counter[12] ),
    .X(_02195_));
 sg13g2_nor2_1 _07552_ (.A(net84),
    .B(_02195_),
    .Y(_00224_));
 sg13g2_nand3_1 _07553_ (.B(\btn_right_debounce.debounce_counter[12] ),
    .C(_02192_),
    .A(_02168_),
    .Y(_02196_));
 sg13g2_xnor2_1 _07554_ (.Y(_02197_),
    .A(_02171_),
    .B(_02196_));
 sg13g2_nor2_1 _07555_ (.A(net84),
    .B(_02197_),
    .Y(_00225_));
 sg13g2_nor2_1 _07556_ (.A(_02171_),
    .B(_02196_),
    .Y(_02198_));
 sg13g2_xnor2_1 _07557_ (.Y(_02199_),
    .A(\btn_right_debounce.debounce_counter[14] ),
    .B(_02198_));
 sg13g2_nor2_1 _07558_ (.A(net84),
    .B(_02199_),
    .Y(_00226_));
 sg13g2_and2_1 _07559_ (.A(\btn_right_debounce.debounce_counter[14] ),
    .B(_02198_),
    .X(_02200_));
 sg13g2_buf_1 _07560_ (.A(_02200_),
    .X(_02201_));
 sg13g2_xnor2_1 _07561_ (.Y(_02202_),
    .A(_02173_),
    .B(_02201_));
 sg13g2_nor2_1 _07562_ (.A(net84),
    .B(_02202_),
    .Y(_00227_));
 sg13g2_nand2_1 _07563_ (.Y(_02203_),
    .A(_02173_),
    .B(_02201_));
 sg13g2_xor2_1 _07564_ (.B(_02203_),
    .A(\btn_right_debounce.debounce_counter[16] ),
    .X(_02204_));
 sg13g2_nor2_1 _07565_ (.A(_02181_),
    .B(_02204_),
    .Y(_00228_));
 sg13g2_nand3_1 _07566_ (.B(\btn_right_debounce.debounce_counter[16] ),
    .C(_02201_),
    .A(_02173_),
    .Y(_02205_));
 sg13g2_xor2_1 _07567_ (.B(_02205_),
    .A(\btn_right_debounce.debounce_counter[17] ),
    .X(_02206_));
 sg13g2_nor2_1 _07568_ (.A(_02181_),
    .B(_02206_),
    .Y(_00229_));
 sg13g2_xnor2_1 _07569_ (.Y(_02207_),
    .A(_02166_),
    .B(_02174_));
 sg13g2_nor2_1 _07570_ (.A(net84),
    .B(_02207_),
    .Y(_00230_));
 sg13g2_nand2_1 _07571_ (.Y(_02208_),
    .A(_02166_),
    .B(_02174_));
 sg13g2_xor2_1 _07572_ (.B(_02208_),
    .A(\btn_right_debounce.debounce_counter[2] ),
    .X(_02209_));
 sg13g2_nor2_1 _07573_ (.A(net147),
    .B(_02209_),
    .Y(_00231_));
 sg13g2_xnor2_1 _07574_ (.Y(_02210_),
    .A(_02184_),
    .B(_02185_));
 sg13g2_nor2_1 _07575_ (.A(net147),
    .B(_02210_),
    .Y(_00232_));
 sg13g2_xnor2_1 _07576_ (.Y(_02211_),
    .A(_02164_),
    .B(_02186_));
 sg13g2_nor2_1 _07577_ (.A(net147),
    .B(_02211_),
    .Y(_00233_));
 sg13g2_nand2_1 _07578_ (.Y(_02212_),
    .A(_02164_),
    .B(_02186_));
 sg13g2_xor2_1 _07579_ (.B(_02212_),
    .A(\btn_right_debounce.debounce_counter[5] ),
    .X(_02213_));
 sg13g2_nor2_1 _07580_ (.A(net147),
    .B(_02213_),
    .Y(_00234_));
 sg13g2_xnor2_1 _07581_ (.Y(_02214_),
    .A(_02163_),
    .B(_02187_));
 sg13g2_nor2_1 _07582_ (.A(net147),
    .B(_02214_),
    .Y(_00235_));
 sg13g2_xnor2_1 _07583_ (.Y(_02215_),
    .A(_02183_),
    .B(_02188_));
 sg13g2_nor2_1 _07584_ (.A(_02180_),
    .B(_02215_),
    .Y(_00236_));
 sg13g2_xnor2_1 _07585_ (.Y(_02216_),
    .A(_02167_),
    .B(_02189_));
 sg13g2_nor2_1 _07586_ (.A(net147),
    .B(_02216_),
    .Y(_00237_));
 sg13g2_nand2_1 _07587_ (.Y(_02217_),
    .A(_02167_),
    .B(_02189_));
 sg13g2_xor2_1 _07588_ (.B(_02217_),
    .A(\btn_right_debounce.debounce_counter[9] ),
    .X(_02218_));
 sg13g2_nor2_1 _07589_ (.A(net147),
    .B(_02218_),
    .Y(_00238_));
 sg13g2_inv_1 _07590_ (.Y(_02219_),
    .A(_00169_));
 sg13g2_inv_1 _07591_ (.Y(_02220_),
    .A(\btn_up_debounce.debounce_counter[6] ));
 sg13g2_buf_1 _07592_ (.A(\btn_up_debounce.debounce_counter[4] ),
    .X(_02221_));
 sg13g2_nor2b_1 _07593_ (.A(\btn_up_debounce.debounce_counter[5] ),
    .B_N(_02221_),
    .Y(_02222_));
 sg13g2_buf_1 _07594_ (.A(\btn_up_debounce.debounce_counter[1] ),
    .X(_02223_));
 sg13g2_buf_1 _07595_ (.A(\btn_up_debounce.debounce_counter[8] ),
    .X(_02224_));
 sg13g2_buf_1 _07596_ (.A(\btn_up_debounce.debounce_counter[11] ),
    .X(_02225_));
 sg13g2_nor4_1 _07597_ (.A(_02223_),
    .B(_02224_),
    .C(_02225_),
    .D(\btn_up_debounce.debounce_counter[10] ),
    .Y(_02226_));
 sg13g2_nand4_1 _07598_ (.B(\btn_up_debounce.debounce_counter[7] ),
    .C(_02222_),
    .A(_02220_),
    .Y(_02227_),
    .D(_02226_));
 sg13g2_inv_1 _07599_ (.Y(_02228_),
    .A(\btn_up_debounce.debounce_counter[13] ));
 sg13g2_nand4_1 _07600_ (.B(\btn_up_debounce.debounce_counter[12] ),
    .C(\btn_up_debounce.debounce_counter[14] ),
    .A(_02228_),
    .Y(_02229_),
    .D(\btn_up_debounce.debounce_counter[17] ));
 sg13g2_buf_1 _07601_ (.A(\btn_up_debounce.debounce_counter[15] ),
    .X(_02230_));
 sg13g2_buf_1 _07602_ (.A(\btn_up_debounce.debounce_counter[0] ),
    .X(_02231_));
 sg13g2_nor4_1 _07603_ (.A(_02231_),
    .B(\btn_up_debounce.debounce_counter[3] ),
    .C(\btn_up_debounce.debounce_counter[2] ),
    .D(\btn_up_debounce.debounce_counter[9] ),
    .Y(_02232_));
 sg13g2_nand3_1 _07604_ (.B(\btn_up_debounce.debounce_counter[16] ),
    .C(_02232_),
    .A(_02230_),
    .Y(_02233_));
 sg13g2_nor3_2 _07605_ (.A(_02227_),
    .B(_02229_),
    .C(_02233_),
    .Y(_02234_));
 sg13g2_xor2_1 _07606_ (.B(\btn_up_debounce.button_sync_1 ),
    .A(_05070_),
    .X(_02235_));
 sg13g2_nand3b_1 _07607_ (.B(_02235_),
    .C(net478),
    .Y(_02236_),
    .A_N(_02234_));
 sg13g2_buf_1 _07608_ (.A(_02236_),
    .X(_02237_));
 sg13g2_buf_1 _07609_ (.A(net146),
    .X(_02238_));
 sg13g2_nor2_1 _07610_ (.A(_02219_),
    .B(net83),
    .Y(_00242_));
 sg13g2_inv_1 _07611_ (.Y(_02239_),
    .A(\btn_up_debounce.debounce_counter[10] ));
 sg13g2_inv_1 _07612_ (.Y(_02240_),
    .A(\btn_up_debounce.debounce_counter[7] ));
 sg13g2_inv_1 _07613_ (.Y(_02241_),
    .A(\btn_up_debounce.debounce_counter[3] ));
 sg13g2_nand3_1 _07614_ (.B(_02231_),
    .C(\btn_up_debounce.debounce_counter[2] ),
    .A(_02223_),
    .Y(_02242_));
 sg13g2_nor2_1 _07615_ (.A(_02241_),
    .B(_02242_),
    .Y(_02243_));
 sg13g2_nand3_1 _07616_ (.B(_02221_),
    .C(_02243_),
    .A(\btn_up_debounce.debounce_counter[5] ),
    .Y(_02244_));
 sg13g2_or2_1 _07617_ (.X(_02245_),
    .B(_02244_),
    .A(_02220_));
 sg13g2_nor2_1 _07618_ (.A(_02240_),
    .B(_02245_),
    .Y(_02246_));
 sg13g2_nand3_1 _07619_ (.B(_02224_),
    .C(_02246_),
    .A(\btn_up_debounce.debounce_counter[9] ),
    .Y(_02247_));
 sg13g2_xnor2_1 _07620_ (.Y(_02248_),
    .A(_02239_),
    .B(_02247_));
 sg13g2_nor2_1 _07621_ (.A(net83),
    .B(_02248_),
    .Y(_00243_));
 sg13g2_nor2_1 _07622_ (.A(_02239_),
    .B(_02247_),
    .Y(_02249_));
 sg13g2_xnor2_1 _07623_ (.Y(_02250_),
    .A(_02225_),
    .B(_02249_));
 sg13g2_nor2_1 _07624_ (.A(net83),
    .B(_02250_),
    .Y(_00244_));
 sg13g2_nand2_1 _07625_ (.Y(_02251_),
    .A(_02225_),
    .B(_02249_));
 sg13g2_xor2_1 _07626_ (.B(_02251_),
    .A(\btn_up_debounce.debounce_counter[12] ),
    .X(_02252_));
 sg13g2_nor2_1 _07627_ (.A(net83),
    .B(_02252_),
    .Y(_00245_));
 sg13g2_nand3_1 _07628_ (.B(\btn_up_debounce.debounce_counter[12] ),
    .C(_02249_),
    .A(_02225_),
    .Y(_02253_));
 sg13g2_xnor2_1 _07629_ (.Y(_02254_),
    .A(_02228_),
    .B(_02253_));
 sg13g2_nor2_1 _07630_ (.A(net83),
    .B(_02254_),
    .Y(_00246_));
 sg13g2_nor2_1 _07631_ (.A(_02228_),
    .B(_02253_),
    .Y(_02255_));
 sg13g2_xnor2_1 _07632_ (.Y(_02256_),
    .A(\btn_up_debounce.debounce_counter[14] ),
    .B(_02255_));
 sg13g2_nor2_1 _07633_ (.A(net83),
    .B(_02256_),
    .Y(_00247_));
 sg13g2_and2_1 _07634_ (.A(\btn_up_debounce.debounce_counter[14] ),
    .B(_02255_),
    .X(_02257_));
 sg13g2_buf_1 _07635_ (.A(_02257_),
    .X(_02258_));
 sg13g2_xnor2_1 _07636_ (.Y(_02259_),
    .A(_02230_),
    .B(_02258_));
 sg13g2_nor2_1 _07637_ (.A(_02238_),
    .B(_02259_),
    .Y(_00248_));
 sg13g2_nand2_1 _07638_ (.Y(_02260_),
    .A(_02230_),
    .B(_02258_));
 sg13g2_xor2_1 _07639_ (.B(_02260_),
    .A(\btn_up_debounce.debounce_counter[16] ),
    .X(_02261_));
 sg13g2_nor2_1 _07640_ (.A(net83),
    .B(_02261_),
    .Y(_00249_));
 sg13g2_nand3_1 _07641_ (.B(\btn_up_debounce.debounce_counter[16] ),
    .C(_02258_),
    .A(_02230_),
    .Y(_02262_));
 sg13g2_xor2_1 _07642_ (.B(_02262_),
    .A(\btn_up_debounce.debounce_counter[17] ),
    .X(_02263_));
 sg13g2_nor2_1 _07643_ (.A(_02238_),
    .B(_02263_),
    .Y(_00250_));
 sg13g2_xnor2_1 _07644_ (.Y(_02264_),
    .A(_02223_),
    .B(_02231_));
 sg13g2_nor2_1 _07645_ (.A(net83),
    .B(_02264_),
    .Y(_00251_));
 sg13g2_nand2_1 _07646_ (.Y(_02265_),
    .A(_02223_),
    .B(_02231_));
 sg13g2_xor2_1 _07647_ (.B(_02265_),
    .A(\btn_up_debounce.debounce_counter[2] ),
    .X(_02266_));
 sg13g2_nor2_1 _07648_ (.A(net146),
    .B(_02266_),
    .Y(_00252_));
 sg13g2_xnor2_1 _07649_ (.Y(_02267_),
    .A(_02241_),
    .B(_02242_));
 sg13g2_nor2_1 _07650_ (.A(net146),
    .B(_02267_),
    .Y(_00253_));
 sg13g2_xnor2_1 _07651_ (.Y(_02268_),
    .A(_02221_),
    .B(_02243_));
 sg13g2_nor2_1 _07652_ (.A(net146),
    .B(_02268_),
    .Y(_00254_));
 sg13g2_nand2_1 _07653_ (.Y(_02269_),
    .A(_02221_),
    .B(_02243_));
 sg13g2_xor2_1 _07654_ (.B(_02269_),
    .A(\btn_up_debounce.debounce_counter[5] ),
    .X(_02270_));
 sg13g2_nor2_1 _07655_ (.A(net146),
    .B(_02270_),
    .Y(_00255_));
 sg13g2_xnor2_1 _07656_ (.Y(_02271_),
    .A(_02220_),
    .B(_02244_));
 sg13g2_nor2_1 _07657_ (.A(net146),
    .B(_02271_),
    .Y(_00256_));
 sg13g2_xnor2_1 _07658_ (.Y(_02272_),
    .A(_02240_),
    .B(_02245_));
 sg13g2_nor2_1 _07659_ (.A(net146),
    .B(_02272_),
    .Y(_00257_));
 sg13g2_xnor2_1 _07660_ (.Y(_02273_),
    .A(_02224_),
    .B(_02246_));
 sg13g2_nor2_1 _07661_ (.A(net146),
    .B(_02273_),
    .Y(_00258_));
 sg13g2_nand2_1 _07662_ (.Y(_02274_),
    .A(_02224_),
    .B(_02246_));
 sg13g2_xor2_1 _07663_ (.B(_02274_),
    .A(\btn_up_debounce.debounce_counter[9] ),
    .X(_02275_));
 sg13g2_nor2_1 _07664_ (.A(_02237_),
    .B(_02275_),
    .Y(_00259_));
 sg13g2_buf_2 _07665_ (.A(_00163_),
    .X(_02276_));
 sg13g2_nor3_1 _07666_ (.A(net457),
    .B(_02276_),
    .C(_01153_),
    .Y(_02277_));
 sg13g2_nand3_1 _07667_ (.B(_01310_),
    .C(_02277_),
    .A(_00844_),
    .Y(_02278_));
 sg13g2_buf_1 _07668_ (.A(_02278_),
    .X(_02279_));
 sg13g2_nor2_1 _07669_ (.A(_00859_),
    .B(_02279_),
    .Y(_00285_));
 sg13g2_nor2_1 _07670_ (.A(_00856_),
    .B(_02279_),
    .Y(_00286_));
 sg13g2_nor2_1 _07671_ (.A(_00885_),
    .B(_02279_),
    .Y(_00287_));
 sg13g2_nor2_1 _07672_ (.A(_00886_),
    .B(_02279_),
    .Y(_00288_));
 sg13g2_and2_1 _07673_ (.A(_00165_),
    .B(_01906_),
    .X(_00417_));
 sg13g2_xnor2_1 _07674_ (.Y(_02280_),
    .A(_01890_),
    .B(net469));
 sg13g2_nor2_1 _07675_ (.A(net361),
    .B(_02280_),
    .Y(_00418_));
 sg13g2_nand2_1 _07676_ (.Y(_02281_),
    .A(_01890_),
    .B(net469));
 sg13g2_xor2_1 _07677_ (.B(_02281_),
    .A(_01892_),
    .X(_02282_));
 sg13g2_nor2_1 _07678_ (.A(net361),
    .B(_02282_),
    .Y(_00419_));
 sg13g2_inv_1 _07679_ (.Y(_02283_),
    .A(_01896_));
 sg13g2_buf_1 _07680_ (.A(net429),
    .X(_02284_));
 sg13g2_buf_1 _07681_ (.A(net385),
    .X(_02285_));
 sg13g2_buf_1 _07682_ (.A(net334),
    .X(_02286_));
 sg13g2_xnor2_1 _07683_ (.Y(_02287_),
    .A(net245),
    .B(_01894_));
 sg13g2_nor2_1 _07684_ (.A(_05061_),
    .B(_02287_),
    .Y(_00420_));
 sg13g2_inv_2 _07685_ (.Y(_02288_),
    .A(net439));
 sg13g2_buf_1 _07686_ (.A(_02288_),
    .X(_02289_));
 sg13g2_buf_1 _07687_ (.A(net333),
    .X(_02290_));
 sg13g2_buf_1 _07688_ (.A(_02290_),
    .X(_02291_));
 sg13g2_or2_1 _07689_ (.X(_02292_),
    .B(_01894_),
    .A(net245));
 sg13g2_xnor2_1 _07690_ (.Y(_02293_),
    .A(net145),
    .B(_02292_));
 sg13g2_nor2_1 _07691_ (.A(_05061_),
    .B(_02293_),
    .Y(_00421_));
 sg13g2_buf_1 _07692_ (.A(_01896_),
    .X(_02294_));
 sg13g2_buf_1 _07693_ (.A(net428),
    .X(_02295_));
 sg13g2_nand2_1 _07694_ (.Y(_02296_),
    .A(net384),
    .B(net439));
 sg13g2_buf_1 _07695_ (.A(_02296_),
    .X(_02297_));
 sg13g2_buf_1 _07696_ (.A(net440),
    .X(_02298_));
 sg13g2_buf_1 _07697_ (.A(net383),
    .X(_02299_));
 sg13g2_buf_1 _07698_ (.A(net332),
    .X(_02300_));
 sg13g2_buf_1 _07699_ (.A(net242),
    .X(_02301_));
 sg13g2_o21ai_1 _07700_ (.B1(net144),
    .Y(_02302_),
    .A1(_01894_),
    .A2(net243));
 sg13g2_a21oi_1 _07701_ (.A1(_01902_),
    .A2(_02302_),
    .Y(_00422_),
    .B1(_01945_));
 sg13g2_nand3_1 _07702_ (.B(net440),
    .C(_01784_),
    .A(net435),
    .Y(_02303_));
 sg13g2_buf_2 _07703_ (.A(_02303_),
    .X(_02304_));
 sg13g2_nor2_2 _07704_ (.A(_01894_),
    .B(_02304_),
    .Y(_02305_));
 sg13g2_xnor2_1 _07705_ (.Y(_02306_),
    .A(net397),
    .B(_02305_));
 sg13g2_nor2_1 _07706_ (.A(_01945_),
    .B(_02306_),
    .Y(_00423_));
 sg13g2_nand2_1 _07707_ (.Y(_02307_),
    .A(net397),
    .B(_02305_));
 sg13g2_xor2_1 _07708_ (.B(_02307_),
    .A(net398),
    .X(_02308_));
 sg13g2_nor2_1 _07709_ (.A(_01945_),
    .B(_02308_),
    .Y(_00424_));
 sg13g2_nand3_1 _07710_ (.B(net397),
    .C(_02305_),
    .A(_01777_),
    .Y(_02309_));
 sg13g2_xnor2_1 _07711_ (.Y(_02310_),
    .A(_01773_),
    .B(_02309_));
 sg13g2_nor2_1 _07712_ (.A(_01945_),
    .B(_02310_),
    .Y(_00425_));
 sg13g2_or2_1 _07713_ (.X(_02311_),
    .B(_02309_),
    .A(_01773_));
 sg13g2_xor2_1 _07714_ (.B(_02311_),
    .A(_01774_),
    .X(_02312_));
 sg13g2_nor2_1 _07715_ (.A(_01945_),
    .B(_02312_),
    .Y(_00426_));
 sg13g2_inv_1 _07716_ (.Y(_02313_),
    .A(_01752_));
 sg13g2_or2_1 _07717_ (.X(_02314_),
    .B(net398),
    .A(_01772_));
 sg13g2_nand2_1 _07718_ (.Y(_02315_),
    .A(_01774_),
    .B(_02314_));
 sg13g2_nand4_1 _07719_ (.B(_02313_),
    .C(_01764_),
    .A(net447),
    .Y(_02316_),
    .D(_02315_));
 sg13g2_buf_1 _07720_ (.A(_02316_),
    .X(_02317_));
 sg13g2_inv_1 _07721_ (.Y(_02318_),
    .A(net468));
 sg13g2_buf_1 _07722_ (.A(_02318_),
    .X(_02319_));
 sg13g2_nor2_2 _07723_ (.A(_01767_),
    .B(net443),
    .Y(_02320_));
 sg13g2_nand2_1 _07724_ (.Y(_02321_),
    .A(net382),
    .B(_02320_));
 sg13g2_buf_2 _07725_ (.A(_02321_),
    .X(_02322_));
 sg13g2_nor4_1 _07726_ (.A(net400),
    .B(net346),
    .C(net90),
    .D(_02322_),
    .Y(_02323_));
 sg13g2_nand3b_1 _07727_ (.B(_02323_),
    .C(net445),
    .Y(_02324_),
    .A_N(net475));
 sg13g2_nor2_1 _07728_ (.A(_01752_),
    .B(_01757_),
    .Y(_02325_));
 sg13g2_nand3_1 _07729_ (.B(_02324_),
    .C(_02325_),
    .A(_00089_),
    .Y(_02326_));
 sg13g2_nor2_1 _07730_ (.A(_01774_),
    .B(_01752_),
    .Y(_02327_));
 sg13g2_nand2_1 _07731_ (.Y(_02328_),
    .A(_01776_),
    .B(_01779_));
 sg13g2_xnor2_1 _07732_ (.Y(_02329_),
    .A(_01772_),
    .B(_02328_));
 sg13g2_nand4_1 _07733_ (.B(_02326_),
    .C(_02327_),
    .A(_01997_),
    .Y(_02330_),
    .D(_02329_));
 sg13g2_buf_1 _07734_ (.A(_02330_),
    .X(_02331_));
 sg13g2_buf_1 _07735_ (.A(_02295_),
    .X(_02332_));
 sg13g2_nor2_2 _07736_ (.A(net331),
    .B(net338),
    .Y(_02333_));
 sg13g2_buf_1 _07737_ (.A(net393),
    .X(_02334_));
 sg13g2_buf_1 _07738_ (.A(net439),
    .X(_02335_));
 sg13g2_buf_1 _07739_ (.A(net381),
    .X(_02336_));
 sg13g2_nor2_1 _07740_ (.A(_02334_),
    .B(net329),
    .Y(_02337_));
 sg13g2_nor3_1 _07741_ (.A(net144),
    .B(_02333_),
    .C(_02337_),
    .Y(_02338_));
 sg13g2_buf_1 _07742_ (.A(net443),
    .X(_02339_));
 sg13g2_buf_1 _07743_ (.A(net380),
    .X(_02340_));
 sg13g2_buf_1 _07744_ (.A(net328),
    .X(_02341_));
 sg13g2_buf_1 _07745_ (.A(net241),
    .X(_02342_));
 sg13g2_buf_1 _07746_ (.A(_02342_),
    .X(_02343_));
 sg13g2_buf_1 _07747_ (.A(net381),
    .X(_02344_));
 sg13g2_buf_1 _07748_ (.A(_00095_),
    .X(_02345_));
 sg13g2_inv_1 _07749_ (.Y(_02346_),
    .A(net463));
 sg13g2_buf_1 _07750_ (.A(_00094_),
    .X(_02347_));
 sg13g2_buf_1 _07751_ (.A(net462),
    .X(_02348_));
 sg13g2_nand2_1 _07752_ (.Y(_02349_),
    .A(net327),
    .B(net427));
 sg13g2_o21ai_1 _07753_ (.B1(_02349_),
    .Y(_02350_),
    .A1(net327),
    .A2(_02346_));
 sg13g2_buf_1 _07754_ (.A(net390),
    .X(_02351_));
 sg13g2_buf_1 _07755_ (.A(net326),
    .X(_02352_));
 sg13g2_buf_1 _07756_ (.A(net240),
    .X(_02353_));
 sg13g2_nor2b_1 _07757_ (.A(net440),
    .B_N(net435),
    .Y(_02354_));
 sg13g2_buf_1 _07758_ (.A(_02354_),
    .X(_02355_));
 sg13g2_buf_1 _07759_ (.A(_02355_),
    .X(_02356_));
 sg13g2_buf_1 _07760_ (.A(net239),
    .X(_02357_));
 sg13g2_nand2b_1 _07761_ (.Y(_02358_),
    .B(net468),
    .A_N(_01767_));
 sg13g2_buf_1 _07762_ (.A(_02358_),
    .X(_02359_));
 sg13g2_buf_1 _07763_ (.A(_02359_),
    .X(_02360_));
 sg13g2_buf_1 _07764_ (.A(_02360_),
    .X(_02361_));
 sg13g2_a21oi_1 _07765_ (.A1(net142),
    .A2(net141),
    .Y(_02362_),
    .B1(net238));
 sg13g2_o21ai_1 _07766_ (.B1(_02362_),
    .Y(_02363_),
    .A1(net82),
    .A2(_02350_));
 sg13g2_o21ai_1 _07767_ (.B1(_02363_),
    .Y(_02364_),
    .A1(net252),
    .A2(_02338_));
 sg13g2_buf_1 _07768_ (.A(net388),
    .X(_02365_));
 sg13g2_buf_1 _07769_ (.A(net324),
    .X(_02366_));
 sg13g2_buf_1 _07770_ (.A(net237),
    .X(_02367_));
 sg13g2_buf_1 _07771_ (.A(net387),
    .X(_02368_));
 sg13g2_buf_1 _07772_ (.A(net323),
    .X(_02369_));
 sg13g2_buf_1 _07773_ (.A(net236),
    .X(_02370_));
 sg13g2_buf_1 _07774_ (.A(net470),
    .X(_02371_));
 sg13g2_nand3b_1 _07775_ (.B(net436),
    .C(net428),
    .Y(_02372_),
    .A_N(net426));
 sg13g2_buf_2 _07776_ (.A(_02372_),
    .X(_02373_));
 sg13g2_or2_1 _07777_ (.X(_02374_),
    .B(_00095_),
    .A(net436));
 sg13g2_buf_2 _07778_ (.A(_02374_),
    .X(_02375_));
 sg13g2_and2_1 _07779_ (.A(_02373_),
    .B(_02375_),
    .X(_02376_));
 sg13g2_buf_1 _07780_ (.A(_02376_),
    .X(_02377_));
 sg13g2_buf_1 _07781_ (.A(_01971_),
    .X(_02378_));
 sg13g2_buf_1 _07782_ (.A(net235),
    .X(_02379_));
 sg13g2_nor2_1 _07783_ (.A(net138),
    .B(_02350_),
    .Y(_02380_));
 sg13g2_buf_1 _07784_ (.A(net330),
    .X(_02381_));
 sg13g2_buf_1 _07785_ (.A(net436),
    .X(_02382_));
 sg13g2_nand2_2 _07786_ (.Y(_02383_),
    .A(net432),
    .B(net379));
 sg13g2_nand2_1 _07787_ (.Y(_02384_),
    .A(_02381_),
    .B(_02383_));
 sg13g2_or2_1 _07788_ (.X(_02385_),
    .B(net379),
    .A(net432));
 sg13g2_buf_1 _07789_ (.A(_02385_),
    .X(_02386_));
 sg13g2_nand2b_1 _07790_ (.Y(_02387_),
    .B(net435),
    .A_N(_02371_));
 sg13g2_buf_2 _07791_ (.A(_02387_),
    .X(_02388_));
 sg13g2_buf_1 _07792_ (.A(_02388_),
    .X(_02389_));
 sg13g2_buf_1 _07793_ (.A(net233),
    .X(_02390_));
 sg13g2_a21oi_1 _07794_ (.A1(_02384_),
    .A2(_02386_),
    .Y(_02391_),
    .B1(_02390_));
 sg13g2_nor3_1 _07795_ (.A(net236),
    .B(_02380_),
    .C(_02391_),
    .Y(_02392_));
 sg13g2_a21oi_1 _07796_ (.A1(net139),
    .A2(_02377_),
    .Y(_02393_),
    .B1(_02392_));
 sg13g2_nor2_1 _07797_ (.A(_02367_),
    .B(_02393_),
    .Y(_02394_));
 sg13g2_nor3_1 _07798_ (.A(_01756_),
    .B(_02364_),
    .C(_02394_),
    .Y(_02395_));
 sg13g2_nor2b_1 _07799_ (.A(net471),
    .B_N(net470),
    .Y(_02396_));
 sg13g2_buf_1 _07800_ (.A(_02396_),
    .X(_02397_));
 sg13g2_buf_1 _07801_ (.A(_02397_),
    .X(_02398_));
 sg13g2_nand2_1 _07802_ (.Y(_02399_),
    .A(net387),
    .B(_01928_));
 sg13g2_buf_1 _07803_ (.A(_02399_),
    .X(_02400_));
 sg13g2_nor2_1 _07804_ (.A(net468),
    .B(net232),
    .Y(_02401_));
 sg13g2_buf_2 _07805_ (.A(_02401_),
    .X(_02402_));
 sg13g2_buf_1 _07806_ (.A(_02402_),
    .X(_02403_));
 sg13g2_nand2_1 _07807_ (.Y(_02404_),
    .A(net394),
    .B(net331));
 sg13g2_and4_1 _07808_ (.A(_01756_),
    .B(net322),
    .C(net60),
    .D(_02404_),
    .X(_02405_));
 sg13g2_o21ai_1 _07809_ (.B1(net400),
    .Y(_02406_),
    .A1(_02395_),
    .A2(_02405_));
 sg13g2_nand2_1 _07810_ (.Y(_02407_),
    .A(net382),
    .B(net387));
 sg13g2_buf_1 _07811_ (.A(_02407_),
    .X(_02408_));
 sg13g2_buf_1 _07812_ (.A(_02408_),
    .X(_02409_));
 sg13g2_buf_1 _07813_ (.A(_00096_),
    .X(_02410_));
 sg13g2_nand3b_1 _07814_ (.B(net436),
    .C(net426),
    .Y(_02411_),
    .A_N(_01896_));
 sg13g2_buf_1 _07815_ (.A(_02411_),
    .X(_02412_));
 sg13g2_buf_1 _07816_ (.A(_02412_),
    .X(_02413_));
 sg13g2_o21ai_1 _07817_ (.B1(net231),
    .Y(_02414_),
    .A1(net383),
    .A2(net461));
 sg13g2_nor2_1 _07818_ (.A(net337),
    .B(_02414_),
    .Y(_02415_));
 sg13g2_nand2_1 _07819_ (.Y(_02416_),
    .A(net429),
    .B(net378));
 sg13g2_buf_2 _07820_ (.A(_02416_),
    .X(_02417_));
 sg13g2_o21ai_1 _07821_ (.B1(net393),
    .Y(_02418_),
    .A1(net467),
    .A2(_02417_));
 sg13g2_nor2b_1 _07822_ (.A(_02415_),
    .B_N(_02418_),
    .Y(_02419_));
 sg13g2_nand2b_1 _07823_ (.Y(_02420_),
    .B(net426),
    .A_N(net471));
 sg13g2_buf_1 _07824_ (.A(_02420_),
    .X(_02421_));
 sg13g2_buf_1 _07825_ (.A(_02421_),
    .X(_02422_));
 sg13g2_buf_1 _07826_ (.A(net230),
    .X(_02423_));
 sg13g2_nor2b_1 _07827_ (.A(net432),
    .B_N(_01766_),
    .Y(_02424_));
 sg13g2_buf_1 _07828_ (.A(_02424_),
    .X(_02425_));
 sg13g2_nand2_1 _07829_ (.Y(_02426_),
    .A(net135),
    .B(_02425_));
 sg13g2_and2_1 _07830_ (.A(_02419_),
    .B(_02426_),
    .X(_02427_));
 sg13g2_inv_1 _07831_ (.Y(_02428_),
    .A(net474));
 sg13g2_buf_1 _07832_ (.A(_00090_),
    .X(_02429_));
 sg13g2_inv_2 _07833_ (.Y(_02430_),
    .A(net460));
 sg13g2_nand2_1 _07834_ (.Y(_02431_),
    .A(_02428_),
    .B(_02430_));
 sg13g2_buf_2 _07835_ (.A(_02431_),
    .X(_02432_));
 sg13g2_buf_1 _07836_ (.A(_02432_),
    .X(_02433_));
 sg13g2_buf_1 _07837_ (.A(_02433_),
    .X(_02434_));
 sg13g2_buf_1 _07838_ (.A(net399),
    .X(_02435_));
 sg13g2_buf_1 _07839_ (.A(net320),
    .X(_02436_));
 sg13g2_nor2_1 _07840_ (.A(net436),
    .B(net426),
    .Y(_02437_));
 sg13g2_nand2_1 _07841_ (.Y(_02438_),
    .A(net384),
    .B(_02437_));
 sg13g2_buf_1 _07842_ (.A(_02438_),
    .X(_02439_));
 sg13g2_or2_1 _07843_ (.X(_02440_),
    .B(_01883_),
    .A(_01765_));
 sg13g2_buf_2 _07844_ (.A(_02440_),
    .X(_02441_));
 sg13g2_or2_1 _07845_ (.X(_02442_),
    .B(_02412_),
    .A(_02441_));
 sg13g2_buf_1 _07846_ (.A(_02442_),
    .X(_02443_));
 sg13g2_and3_1 _07847_ (.X(_02444_),
    .A(net228),
    .B(net227),
    .C(_02443_));
 sg13g2_nand2_1 _07848_ (.Y(_02445_),
    .A(net382),
    .B(net434));
 sg13g2_buf_1 _07849_ (.A(_02445_),
    .X(_02446_));
 sg13g2_nor2_2 _07850_ (.A(net383),
    .B(net463),
    .Y(_02447_));
 sg13g2_inv_1 _07851_ (.Y(_02448_),
    .A(net436));
 sg13g2_nand2b_1 _07852_ (.Y(_02449_),
    .B(net470),
    .A_N(_01896_));
 sg13g2_buf_1 _07853_ (.A(_02449_),
    .X(_02450_));
 sg13g2_nor2_1 _07854_ (.A(_02448_),
    .B(net377),
    .Y(_02451_));
 sg13g2_buf_1 _07855_ (.A(_02451_),
    .X(_02452_));
 sg13g2_nor2_2 _07856_ (.A(_02447_),
    .B(net225),
    .Y(_02453_));
 sg13g2_buf_1 _07857_ (.A(net335),
    .X(_02454_));
 sg13g2_xnor2_1 _07858_ (.Y(_02455_),
    .A(net428),
    .B(net436));
 sg13g2_nor2_2 _07859_ (.A(_02288_),
    .B(_02455_),
    .Y(_02456_));
 sg13g2_nand2_1 _07860_ (.Y(_02457_),
    .A(net224),
    .B(_02456_));
 sg13g2_o21ai_1 _07861_ (.B1(_02457_),
    .Y(_02458_),
    .A1(net138),
    .A2(_02453_));
 sg13g2_nor2_1 _07862_ (.A(net226),
    .B(_02458_),
    .Y(_02459_));
 sg13g2_buf_1 _07863_ (.A(_02448_),
    .X(_02460_));
 sg13g2_nor2_2 _07864_ (.A(net319),
    .B(_02388_),
    .Y(_02461_));
 sg13g2_or2_1 _07865_ (.X(_02462_),
    .B(net426),
    .A(_01896_));
 sg13g2_buf_1 _07866_ (.A(_02462_),
    .X(_02463_));
 sg13g2_o21ai_1 _07867_ (.B1(_02463_),
    .Y(_02464_),
    .A1(net394),
    .A2(_02296_));
 sg13g2_nand2_1 _07868_ (.Y(_02465_),
    .A(net152),
    .B(_02464_));
 sg13g2_buf_1 _07869_ (.A(_02463_),
    .X(_02466_));
 sg13g2_nor2_1 _07870_ (.A(net389),
    .B(net223),
    .Y(_02467_));
 sg13g2_buf_1 _07871_ (.A(net393),
    .X(_02468_));
 sg13g2_inv_1 _07872_ (.Y(_02469_),
    .A(net437));
 sg13g2_buf_1 _07873_ (.A(_02469_),
    .X(_02470_));
 sg13g2_buf_1 _07874_ (.A(net317),
    .X(_02471_));
 sg13g2_buf_1 _07875_ (.A(_02346_),
    .X(_02472_));
 sg13g2_nor3_1 _07876_ (.A(net318),
    .B(net222),
    .C(net376),
    .Y(_02473_));
 sg13g2_nor3_1 _07877_ (.A(net144),
    .B(_02467_),
    .C(_02473_),
    .Y(_02474_));
 sg13g2_a221oi_1 _07878_ (.B2(_02474_),
    .C1(net252),
    .B1(_02465_),
    .A1(net88),
    .Y(_02475_),
    .A2(_02461_));
 sg13g2_nor4_1 _07879_ (.A(net134),
    .B(_02444_),
    .C(_02459_),
    .D(_02475_),
    .Y(_02476_));
 sg13g2_o21ai_1 _07880_ (.B1(_02476_),
    .Y(_02477_),
    .A1(net136),
    .A2(_02427_));
 sg13g2_mux4_1 _07881_ (.S0(net442),
    .A0(\draw_game_inst.grid[39] ),
    .A1(\draw_game_inst.grid[47] ),
    .A2(\draw_game_inst.grid[43] ),
    .A3(\draw_game_inst.grid[35] ),
    .S1(net472),
    .X(_02478_));
 sg13g2_mux4_1 _07882_ (.S0(net442),
    .A0(\draw_game_inst.grid[7] ),
    .A1(\draw_game_inst.grid[15] ),
    .A2(\draw_game_inst.grid[11] ),
    .A3(\draw_game_inst.grid[3] ),
    .S1(net441),
    .X(_02479_));
 sg13g2_mux4_1 _07883_ (.S0(net473),
    .A0(\draw_game_inst.grid[55] ),
    .A1(\draw_game_inst.grid[63] ),
    .A2(\draw_game_inst.grid[59] ),
    .A3(\draw_game_inst.grid[51] ),
    .S1(net472),
    .X(_02480_));
 sg13g2_mux4_1 _07884_ (.S0(net473),
    .A0(\draw_game_inst.grid[23] ),
    .A1(\draw_game_inst.grid[31] ),
    .A2(\draw_game_inst.grid[27] ),
    .A3(\draw_game_inst.grid[19] ),
    .S1(net472),
    .X(_02481_));
 sg13g2_mux4_1 _07885_ (.S0(_01758_),
    .A0(_02478_),
    .A1(_02479_),
    .A2(_02480_),
    .A3(_02481_),
    .S1(net475),
    .X(_02482_));
 sg13g2_mux4_1 _07886_ (.S0(_01775_),
    .A0(\draw_game_inst.grid[38] ),
    .A1(\draw_game_inst.grid[46] ),
    .A2(\draw_game_inst.grid[42] ),
    .A3(\draw_game_inst.grid[34] ),
    .S1(_01778_),
    .X(_02483_));
 sg13g2_mux4_1 _07887_ (.S0(net473),
    .A0(\draw_game_inst.grid[6] ),
    .A1(\draw_game_inst.grid[14] ),
    .A2(\draw_game_inst.grid[10] ),
    .A3(\draw_game_inst.grid[2] ),
    .S1(net472),
    .X(_02484_));
 sg13g2_mux4_1 _07888_ (.S0(net473),
    .A0(\draw_game_inst.grid[54] ),
    .A1(\draw_game_inst.grid[62] ),
    .A2(\draw_game_inst.grid[58] ),
    .A3(\draw_game_inst.grid[50] ),
    .S1(_01778_),
    .X(_02485_));
 sg13g2_mux4_1 _07889_ (.S0(net473),
    .A0(\draw_game_inst.grid[22] ),
    .A1(\draw_game_inst.grid[30] ),
    .A2(\draw_game_inst.grid[26] ),
    .A3(\draw_game_inst.grid[18] ),
    .S1(net472),
    .X(_02486_));
 sg13g2_mux4_1 _07890_ (.S0(_01758_),
    .A0(_02483_),
    .A1(_02484_),
    .A2(_02485_),
    .A3(_02486_),
    .S1(\draw_game_inst.board_y[6] ),
    .X(_02487_));
 sg13g2_nor2b_1 _07891_ (.A(_02482_),
    .B_N(_02487_),
    .Y(_02488_));
 sg13g2_buf_1 _07892_ (.A(_02488_),
    .X(_02489_));
 sg13g2_mux4_1 _07893_ (.S0(net442),
    .A0(\draw_game_inst.grid[37] ),
    .A1(\draw_game_inst.grid[45] ),
    .A2(\draw_game_inst.grid[41] ),
    .A3(\draw_game_inst.grid[33] ),
    .S1(net441),
    .X(_02490_));
 sg13g2_mux4_1 _07894_ (.S0(net442),
    .A0(\draw_game_inst.grid[5] ),
    .A1(\draw_game_inst.grid[13] ),
    .A2(\draw_game_inst.grid[9] ),
    .A3(\draw_game_inst.grid[1] ),
    .S1(net441),
    .X(_02491_));
 sg13g2_mux4_1 _07895_ (.S0(net442),
    .A0(\draw_game_inst.grid[53] ),
    .A1(\draw_game_inst.grid[61] ),
    .A2(\draw_game_inst.grid[57] ),
    .A3(\draw_game_inst.grid[49] ),
    .S1(net441),
    .X(_02492_));
 sg13g2_mux4_1 _07896_ (.S0(net442),
    .A0(\draw_game_inst.grid[21] ),
    .A1(\draw_game_inst.grid[29] ),
    .A2(\draw_game_inst.grid[25] ),
    .A3(\draw_game_inst.grid[17] ),
    .S1(net441),
    .X(_02493_));
 sg13g2_mux4_1 _07897_ (.S0(_01759_),
    .A0(_02490_),
    .A1(_02491_),
    .A2(_02492_),
    .A3(_02493_),
    .S1(net475),
    .X(_02494_));
 sg13g2_buf_1 _07898_ (.A(_02494_),
    .X(_02495_));
 sg13g2_inv_1 _07899_ (.Y(_02496_),
    .A(_02495_));
 sg13g2_mux4_1 _07900_ (.S0(net442),
    .A0(\draw_game_inst.grid[36] ),
    .A1(\draw_game_inst.grid[44] ),
    .A2(\draw_game_inst.grid[40] ),
    .A3(\draw_game_inst.grid[32] ),
    .S1(net441),
    .X(_02497_));
 sg13g2_mux4_1 _07901_ (.S0(net442),
    .A0(\draw_game_inst.grid[4] ),
    .A1(\draw_game_inst.grid[12] ),
    .A2(\draw_game_inst.grid[8] ),
    .A3(\draw_game_inst.grid[0] ),
    .S1(net441),
    .X(_02498_));
 sg13g2_mux4_1 _07902_ (.S0(net473),
    .A0(\draw_game_inst.grid[52] ),
    .A1(\draw_game_inst.grid[60] ),
    .A2(\draw_game_inst.grid[56] ),
    .A3(\draw_game_inst.grid[48] ),
    .S1(net472),
    .X(_02499_));
 sg13g2_mux4_1 _07903_ (.S0(net473),
    .A0(\draw_game_inst.grid[20] ),
    .A1(\draw_game_inst.grid[28] ),
    .A2(\draw_game_inst.grid[24] ),
    .A3(\draw_game_inst.grid[16] ),
    .S1(net472),
    .X(_02500_));
 sg13g2_mux4_1 _07904_ (.S0(_01758_),
    .A0(_02497_),
    .A1(_02498_),
    .A2(_02499_),
    .A3(_02500_),
    .S1(net475),
    .X(_02501_));
 sg13g2_buf_2 _07905_ (.A(_02501_),
    .X(_02502_));
 sg13g2_nor2_2 _07906_ (.A(_02496_),
    .B(_02502_),
    .Y(_02503_));
 sg13g2_nand2_2 _07907_ (.Y(_02504_),
    .A(_02489_),
    .B(_02503_));
 sg13g2_a21oi_1 _07908_ (.A1(_02406_),
    .A2(_02477_),
    .Y(_02505_),
    .B1(_02504_));
 sg13g2_buf_1 _07909_ (.A(_02428_),
    .X(_02506_));
 sg13g2_buf_1 _07910_ (.A(net375),
    .X(_02507_));
 sg13g2_nand2b_1 _07911_ (.Y(_02508_),
    .B(net471),
    .A_N(_01783_));
 sg13g2_buf_1 _07912_ (.A(_02508_),
    .X(_02509_));
 sg13g2_o21ai_1 _07913_ (.B1(net230),
    .Y(_02510_),
    .A1(net342),
    .A2(_02509_));
 sg13g2_nor2_2 _07914_ (.A(net380),
    .B(net429),
    .Y(_02511_));
 sg13g2_a22oi_1 _07915_ (.Y(_02512_),
    .B1(_02510_),
    .B2(_02511_),
    .A2(_02384_),
    .A1(net376));
 sg13g2_buf_1 _07916_ (.A(net461),
    .X(_02513_));
 sg13g2_nor2_1 _07917_ (.A(_02299_),
    .B(_02513_),
    .Y(_02514_));
 sg13g2_o21ai_1 _07918_ (.B1(net82),
    .Y(_02515_),
    .A1(_02461_),
    .A2(_02514_));
 sg13g2_nor2b_1 _07919_ (.A(net428),
    .B_N(net426),
    .Y(_02516_));
 sg13g2_buf_1 _07920_ (.A(_02516_),
    .X(_02517_));
 sg13g2_buf_1 _07921_ (.A(_02517_),
    .X(_02518_));
 sg13g2_buf_1 _07922_ (.A(net221),
    .X(_02519_));
 sg13g2_buf_1 _07923_ (.A(_01953_),
    .X(_02520_));
 sg13g2_nor2_2 _07924_ (.A(net315),
    .B(net433),
    .Y(_02521_));
 sg13g2_buf_1 _07925_ (.A(net332),
    .X(_02522_));
 sg13g2_nand2_1 _07926_ (.Y(_02523_),
    .A(net315),
    .B(net220));
 sg13g2_nand2b_1 _07927_ (.Y(_02524_),
    .B(_02523_),
    .A_N(_02521_));
 sg13g2_buf_1 _07928_ (.A(net392),
    .X(_02525_));
 sg13g2_buf_1 _07929_ (.A(_02525_),
    .X(_02526_));
 sg13g2_buf_1 _07930_ (.A(net219),
    .X(_02527_));
 sg13g2_a21oi_1 _07931_ (.A1(_02519_),
    .A2(_02524_),
    .Y(_02528_),
    .B1(net132));
 sg13g2_a22oi_1 _07932_ (.Y(_02529_),
    .B1(_02515_),
    .B2(_02528_),
    .A2(_02512_),
    .A1(net151));
 sg13g2_buf_1 _07933_ (.A(net460),
    .X(_02530_));
 sg13g2_buf_1 _07934_ (.A(net380),
    .X(_02531_));
 sg13g2_buf_1 _07935_ (.A(_02531_),
    .X(_02532_));
 sg13g2_buf_1 _07936_ (.A(_02532_),
    .X(_02533_));
 sg13g2_buf_1 _07937_ (.A(net389),
    .X(_02534_));
 sg13g2_nand2_2 _07938_ (.Y(_02535_),
    .A(_02304_),
    .B(_02375_));
 sg13g2_nor2_1 _07939_ (.A(net312),
    .B(_02535_),
    .Y(_02536_));
 sg13g2_buf_1 _07940_ (.A(net315),
    .X(_02537_));
 sg13g2_buf_1 _07941_ (.A(net389),
    .X(_02538_));
 sg13g2_mux2_1 _07942_ (.A0(net376),
    .A1(_02535_),
    .S(_02538_),
    .X(_02539_));
 sg13g2_nor2_1 _07943_ (.A(net217),
    .B(_02539_),
    .Y(_02540_));
 sg13g2_a21oi_1 _07944_ (.A1(net131),
    .A2(_02536_),
    .Y(_02541_),
    .B1(_02540_));
 sg13g2_nor2_1 _07945_ (.A(net238),
    .B(_02541_),
    .Y(_02542_));
 sg13g2_nor2_1 _07946_ (.A(_02348_),
    .B(_02296_),
    .Y(_02543_));
 sg13g2_buf_2 _07947_ (.A(_02543_),
    .X(_02544_));
 sg13g2_nand2_1 _07948_ (.Y(_02545_),
    .A(net254),
    .B(net253));
 sg13g2_nor3_1 _07949_ (.A(_01771_),
    .B(_02544_),
    .C(_02545_),
    .Y(_02546_));
 sg13g2_and2_1 _07950_ (.A(net428),
    .B(net426),
    .X(_02547_));
 sg13g2_buf_1 _07951_ (.A(_02547_),
    .X(_02548_));
 sg13g2_buf_1 _07952_ (.A(net310),
    .X(_02549_));
 sg13g2_a21oi_1 _07953_ (.A1(net216),
    .A2(_02523_),
    .Y(_02550_),
    .B1(net252));
 sg13g2_nor4_1 _07954_ (.A(_02530_),
    .B(_02542_),
    .C(_02546_),
    .D(_02550_),
    .Y(_02551_));
 sg13g2_o21ai_1 _07955_ (.B1(_02551_),
    .Y(_02552_),
    .A1(_01964_),
    .A2(_02529_));
 sg13g2_nor2_1 _07956_ (.A(net468),
    .B(net434),
    .Y(_02553_));
 sg13g2_buf_1 _07957_ (.A(_02553_),
    .X(_02554_));
 sg13g2_buf_1 _07958_ (.A(_02554_),
    .X(_02555_));
 sg13g2_nand3_1 _07959_ (.B(net435),
    .C(net439),
    .A(net437),
    .Y(_02556_));
 sg13g2_or2_1 _07960_ (.X(_02557_),
    .B(net461),
    .A(_01883_));
 sg13g2_buf_1 _07961_ (.A(_02557_),
    .X(_02558_));
 sg13g2_a21oi_1 _07962_ (.A1(_02556_),
    .A2(_02558_),
    .Y(_02559_),
    .B1(net383));
 sg13g2_nor3_1 _07963_ (.A(net393),
    .B(net225),
    .C(_02559_),
    .Y(_02560_));
 sg13g2_buf_1 _07964_ (.A(net338),
    .X(_02561_));
 sg13g2_buf_1 _07965_ (.A(net214),
    .X(_02562_));
 sg13g2_nor2_1 _07966_ (.A(net462),
    .B(net377),
    .Y(_02563_));
 sg13g2_buf_2 _07967_ (.A(_02563_),
    .X(_02564_));
 sg13g2_buf_1 _07968_ (.A(_02564_),
    .X(_02565_));
 sg13g2_a21oi_1 _07969_ (.A1(net130),
    .A2(net129),
    .Y(_02566_),
    .B1(net226));
 sg13g2_nor2b_1 _07970_ (.A(net432),
    .B_N(_02295_),
    .Y(_02567_));
 sg13g2_buf_1 _07971_ (.A(_02567_),
    .X(_02568_));
 sg13g2_o21ai_1 _07972_ (.B1(_02402_),
    .Y(_02569_),
    .A1(net135),
    .A2(net213));
 sg13g2_nor2_2 _07973_ (.A(net380),
    .B(net319),
    .Y(_02570_));
 sg13g2_o21ai_1 _07974_ (.B1(_01769_),
    .Y(_02571_),
    .A1(net137),
    .A2(_02570_));
 sg13g2_nand3_1 _07975_ (.B(_02569_),
    .C(_02571_),
    .A(_01913_),
    .Y(_02572_));
 sg13g2_a221oi_1 _07976_ (.B2(_02566_),
    .C1(_02572_),
    .B1(_02457_),
    .A1(net215),
    .Y(_02573_),
    .A2(_02560_));
 sg13g2_nand3_1 _07977_ (.B(_02373_),
    .C(_02375_),
    .A(net335),
    .Y(_02574_));
 sg13g2_nor2b_1 _07978_ (.A(net470),
    .B_N(net471),
    .Y(_02575_));
 sg13g2_buf_2 _07979_ (.A(_02575_),
    .X(_02576_));
 sg13g2_nand2_1 _07980_ (.Y(_02577_),
    .A(net429),
    .B(_02576_));
 sg13g2_buf_1 _07981_ (.A(_02577_),
    .X(_02578_));
 sg13g2_nand2_1 _07982_ (.Y(_02579_),
    .A(net319),
    .B(net425));
 sg13g2_nand2_1 _07983_ (.Y(_02580_),
    .A(net212),
    .B(_02579_));
 sg13g2_nand2_1 _07984_ (.Y(_02581_),
    .A(net150),
    .B(_02580_));
 sg13g2_a21o_1 _07985_ (.A2(_02581_),
    .A1(_02574_),
    .B1(net252),
    .X(_02582_));
 sg13g2_buf_1 _07986_ (.A(net312),
    .X(_02583_));
 sg13g2_buf_1 _07987_ (.A(net211),
    .X(_02584_));
 sg13g2_buf_1 _07988_ (.A(net385),
    .X(_02585_));
 sg13g2_inv_1 _07989_ (.Y(_02586_),
    .A(net462));
 sg13g2_buf_1 _07990_ (.A(net423),
    .X(_02587_));
 sg13g2_nor2_1 _07991_ (.A(_02585_),
    .B(net374),
    .Y(_02588_));
 sg13g2_a21oi_1 _07992_ (.A1(_02585_),
    .A2(_02513_),
    .Y(_02589_),
    .B1(_02588_));
 sg13g2_nand2_1 _07993_ (.Y(_02590_),
    .A(net128),
    .B(_02589_));
 sg13g2_o21ai_1 _07994_ (.B1(_02590_),
    .Y(_02591_),
    .A1(net90),
    .A2(_02580_));
 sg13g2_nor2_1 _07995_ (.A(_01913_),
    .B(_02322_),
    .Y(_02592_));
 sg13g2_buf_2 _07996_ (.A(_02592_),
    .X(_02593_));
 sg13g2_a22oi_1 _07997_ (.Y(_02594_),
    .B1(_02591_),
    .B2(_02593_),
    .A2(_02582_),
    .A1(_02573_));
 sg13g2_nor2b_1 _07998_ (.A(_02495_),
    .B_N(_02502_),
    .Y(_02595_));
 sg13g2_nand2_1 _07999_ (.Y(_02596_),
    .A(_02489_),
    .B(_02595_));
 sg13g2_a21o_1 _08000_ (.A2(_02594_),
    .A1(net444),
    .B1(_02596_),
    .X(_02597_));
 sg13g2_a21o_1 _08001_ (.A2(_02552_),
    .A1(_02507_),
    .B1(_02597_),
    .X(_02598_));
 sg13g2_xor2_1 _08002_ (.B(_02371_),
    .A(net428),
    .X(_02599_));
 sg13g2_buf_1 _08003_ (.A(_02599_),
    .X(_02600_));
 sg13g2_nand2_2 _08004_ (.Y(_02601_),
    .A(net423),
    .B(net308));
 sg13g2_nor2_1 _08005_ (.A(_02322_),
    .B(_02601_),
    .Y(_02602_));
 sg13g2_nor2_2 _08006_ (.A(_02495_),
    .B(_02502_),
    .Y(_02603_));
 sg13g2_and2_1 _08007_ (.A(_02489_),
    .B(_02603_),
    .X(_02604_));
 sg13g2_o21ai_1 _08008_ (.B1(_02604_),
    .Y(_02605_),
    .A1(net386),
    .A2(_02602_));
 sg13g2_inv_1 _08009_ (.Y(_02606_),
    .A(_02605_));
 sg13g2_buf_1 _08010_ (.A(net377),
    .X(_02607_));
 sg13g2_a21oi_1 _08011_ (.A1(net307),
    .A2(_02373_),
    .Y(_02608_),
    .B1(net234));
 sg13g2_a21oi_1 _08012_ (.A1(net129),
    .A2(_02521_),
    .Y(_02609_),
    .B1(_02608_));
 sg13g2_a21oi_1 _08013_ (.A1(net215),
    .A2(_02609_),
    .Y(_02610_),
    .B1(net460));
 sg13g2_xor2_1 _08014_ (.B(net426),
    .A(_01895_),
    .X(_02611_));
 sg13g2_buf_2 _08015_ (.A(_02611_),
    .X(_02612_));
 sg13g2_buf_1 _08016_ (.A(_02455_),
    .X(_02613_));
 sg13g2_nand2_2 _08017_ (.Y(_02614_),
    .A(_02612_),
    .B(net306));
 sg13g2_nand2_1 _08018_ (.Y(_02615_),
    .A(net138),
    .B(_02614_));
 sg13g2_o21ai_1 _08019_ (.B1(_02615_),
    .Y(_02616_),
    .A1(net138),
    .A2(_02544_));
 sg13g2_nand2_1 _08020_ (.Y(_02617_),
    .A(net246),
    .B(_02616_));
 sg13g2_buf_1 _08021_ (.A(net462),
    .X(_02618_));
 sg13g2_buf_1 _08022_ (.A(net422),
    .X(_02619_));
 sg13g2_and2_1 _08023_ (.A(net434),
    .B(net443),
    .X(_02620_));
 sg13g2_buf_1 _08024_ (.A(_02620_),
    .X(_02621_));
 sg13g2_buf_1 _08025_ (.A(_02621_),
    .X(_02622_));
 sg13g2_nor2b_1 _08026_ (.A(net470),
    .B_N(_01896_),
    .Y(_02623_));
 sg13g2_buf_1 _08027_ (.A(_02623_),
    .X(_02624_));
 sg13g2_buf_1 _08028_ (.A(_02624_),
    .X(_02625_));
 sg13g2_buf_1 _08029_ (.A(_02625_),
    .X(_02626_));
 sg13g2_buf_1 _08030_ (.A(_02332_),
    .X(_02627_));
 sg13g2_buf_1 _08031_ (.A(net208),
    .X(_02628_));
 sg13g2_buf_1 _08032_ (.A(_02320_),
    .X(_02629_));
 sg13g2_buf_1 _08033_ (.A(net392),
    .X(_02630_));
 sg13g2_a22oi_1 _08034_ (.Y(_02631_),
    .B1(_02333_),
    .B2(net302),
    .A2(net303),
    .A1(net127));
 sg13g2_inv_1 _08035_ (.Y(_02632_),
    .A(_02631_));
 sg13g2_buf_1 _08036_ (.A(_02336_),
    .X(_02633_));
 sg13g2_buf_1 _08037_ (.A(net207),
    .X(_02634_));
 sg13g2_a22oi_1 _08038_ (.Y(_02635_),
    .B1(_02632_),
    .B2(net126),
    .A2(net209),
    .A1(net210));
 sg13g2_buf_1 _08039_ (.A(net431),
    .X(_02636_));
 sg13g2_buf_1 _08040_ (.A(net372),
    .X(_02637_));
 sg13g2_buf_1 _08041_ (.A(net301),
    .X(_02638_));
 sg13g2_o21ai_1 _08042_ (.B1(net206),
    .Y(_02639_),
    .A1(net373),
    .A2(_02635_));
 sg13g2_nand3_1 _08043_ (.B(_02617_),
    .C(_02639_),
    .A(_02610_),
    .Y(_02640_));
 sg13g2_nand2_1 _08044_ (.Y(_02641_),
    .A(net423),
    .B(_02517_));
 sg13g2_buf_2 _08045_ (.A(_02641_),
    .X(_02642_));
 sg13g2_a21oi_1 _08046_ (.A1(net90),
    .A2(_02642_),
    .Y(_02643_),
    .B1(_01913_));
 sg13g2_nor2_2 _08047_ (.A(net427),
    .B(_02388_),
    .Y(_02644_));
 sg13g2_buf_1 _08048_ (.A(_02644_),
    .X(_02645_));
 sg13g2_nand2_1 _08049_ (.Y(_02646_),
    .A(_01928_),
    .B(net467));
 sg13g2_buf_2 _08050_ (.A(_02646_),
    .X(_02647_));
 sg13g2_a221oi_1 _08051_ (.B2(net150),
    .C1(net252),
    .B1(net129),
    .A1(net125),
    .Y(_02648_),
    .A2(_02647_));
 sg13g2_nor3_1 _08052_ (.A(net324),
    .B(net303),
    .C(_02544_),
    .Y(_02649_));
 sg13g2_buf_1 _08053_ (.A(net392),
    .X(_02650_));
 sg13g2_buf_1 _08054_ (.A(_02650_),
    .X(_02651_));
 sg13g2_nand2_1 _08055_ (.Y(_02652_),
    .A(net423),
    .B(net310));
 sg13g2_buf_2 _08056_ (.A(_02652_),
    .X(_02653_));
 sg13g2_nor2_1 _08057_ (.A(net388),
    .B(net241),
    .Y(_02654_));
 sg13g2_nor2_2 _08058_ (.A(_02344_),
    .B(net422),
    .Y(_02655_));
 sg13g2_nand2_2 _08059_ (.Y(_02656_),
    .A(_02655_),
    .B(net213));
 sg13g2_a22oi_1 _08060_ (.Y(_02657_),
    .B1(_02654_),
    .B2(_02656_),
    .A2(_02653_),
    .A1(net372));
 sg13g2_nor2_1 _08061_ (.A(net205),
    .B(_02657_),
    .Y(_02658_));
 sg13g2_nor4_1 _08062_ (.A(net401),
    .B(_02648_),
    .C(_02649_),
    .D(_02658_),
    .Y(_02659_));
 sg13g2_buf_1 _08063_ (.A(net474),
    .X(_02660_));
 sg13g2_o21ai_1 _08064_ (.B1(net421),
    .Y(_02661_),
    .A1(_02643_),
    .A2(_02659_));
 sg13g2_o21ai_1 _08065_ (.B1(_02661_),
    .Y(_02662_),
    .A1(net444),
    .A2(_02640_));
 sg13g2_nor2_2 _08066_ (.A(_02482_),
    .B(_02487_),
    .Y(_02663_));
 sg13g2_nand2_2 _08067_ (.Y(_02664_),
    .A(_02663_),
    .B(_02503_));
 sg13g2_nand2_1 _08068_ (.Y(_02665_),
    .A(net234),
    .B(net125));
 sg13g2_buf_1 _08069_ (.A(_02576_),
    .X(_02666_));
 sg13g2_buf_1 _08070_ (.A(net299),
    .X(_02667_));
 sg13g2_a21oi_1 _08071_ (.A1(net142),
    .A2(net204),
    .Y(_02668_),
    .B1(net226));
 sg13g2_a21oi_1 _08072_ (.A1(_02665_),
    .A2(_02668_),
    .Y(_02669_),
    .B1(net424));
 sg13g2_a21oi_1 _08073_ (.A1(net125),
    .A2(_02647_),
    .Y(_02670_),
    .B1(net249));
 sg13g2_buf_1 _08074_ (.A(net399),
    .X(_02671_));
 sg13g2_buf_1 _08075_ (.A(net323),
    .X(_02672_));
 sg13g2_nand2_1 _08076_ (.Y(_02673_),
    .A(net423),
    .B(net304));
 sg13g2_buf_1 _08077_ (.A(_02673_),
    .X(_02674_));
 sg13g2_nor2_1 _08078_ (.A(_02672_),
    .B(net124),
    .Y(_02675_));
 sg13g2_a21oi_1 _08079_ (.A1(net298),
    .A2(net204),
    .Y(_02676_),
    .B1(_02675_));
 sg13g2_o21ai_1 _08080_ (.B1(_02676_),
    .Y(_02677_),
    .A1(net206),
    .A2(_02670_));
 sg13g2_a21oi_1 _08081_ (.A1(_02669_),
    .A2(_02677_),
    .Y(_02678_),
    .B1(net421));
 sg13g2_buf_1 _08082_ (.A(net382),
    .X(_02679_));
 sg13g2_buf_1 _08083_ (.A(_02679_),
    .X(_02680_));
 sg13g2_buf_1 _08084_ (.A(net202),
    .X(_02681_));
 sg13g2_nand2_2 _08085_ (.Y(_02682_),
    .A(net214),
    .B(net299));
 sg13g2_xnor2_1 _08086_ (.Y(_02683_),
    .A(net471),
    .B(net470));
 sg13g2_buf_2 _08087_ (.A(_02683_),
    .X(_02684_));
 sg13g2_nor2_1 _08088_ (.A(net429),
    .B(_02684_),
    .Y(_02685_));
 sg13g2_buf_1 _08089_ (.A(_02685_),
    .X(_02686_));
 sg13g2_nor2_1 _08090_ (.A(_02445_),
    .B(net201),
    .Y(_02687_));
 sg13g2_buf_1 _08091_ (.A(net380),
    .X(_02688_));
 sg13g2_buf_1 _08092_ (.A(net296),
    .X(_02689_));
 sg13g2_nor2_1 _08093_ (.A(net328),
    .B(_02673_),
    .Y(_02690_));
 sg13g2_a21oi_1 _08094_ (.A1(net200),
    .A2(net201),
    .Y(_02691_),
    .B1(_02690_));
 sg13g2_a221oi_1 _08095_ (.B2(_02554_),
    .C1(net446),
    .B1(_02691_),
    .A1(_02682_),
    .Y(_02692_),
    .A2(_02687_));
 sg13g2_buf_1 _08096_ (.A(net303),
    .X(_02693_));
 sg13g2_nand3_1 _08097_ (.B(net199),
    .C(net125),
    .A(_01754_),
    .Y(_02694_));
 sg13g2_nand2b_1 _08098_ (.Y(_02695_),
    .B(_02694_),
    .A_N(_02692_));
 sg13g2_nand2_2 _08099_ (.Y(_02696_),
    .A(_01899_),
    .B(_02509_));
 sg13g2_nand2_1 _08100_ (.Y(_02697_),
    .A(_02320_),
    .B(_02696_));
 sg13g2_o21ai_1 _08101_ (.B1(_02697_),
    .Y(_02698_),
    .A1(net199),
    .A2(net124));
 sg13g2_a221oi_1 _08102_ (.B2(_02692_),
    .C1(net375),
    .B1(_02698_),
    .A1(net123),
    .Y(_02699_),
    .A2(_02695_));
 sg13g2_nor3_1 _08103_ (.A(_02664_),
    .B(_02678_),
    .C(_02699_),
    .Y(_02700_));
 sg13g2_a21oi_1 _08104_ (.A1(_02606_),
    .A2(_02662_),
    .Y(_02701_),
    .B1(_02700_));
 sg13g2_nand2_1 _08105_ (.Y(_02702_),
    .A(net474),
    .B(_01913_));
 sg13g2_buf_2 _08106_ (.A(_02702_),
    .X(_02703_));
 sg13g2_buf_1 _08107_ (.A(_02703_),
    .X(_02704_));
 sg13g2_buf_1 _08108_ (.A(net198),
    .X(_02705_));
 sg13g2_buf_1 _08109_ (.A(_02672_),
    .X(_02706_));
 sg13g2_nand2_1 _08110_ (.Y(_02707_),
    .A(net379),
    .B(_02335_));
 sg13g2_buf_1 _08111_ (.A(_02707_),
    .X(_02708_));
 sg13g2_nor2_1 _08112_ (.A(net429),
    .B(_01788_),
    .Y(_02709_));
 sg13g2_buf_1 _08113_ (.A(_02709_),
    .X(_02710_));
 sg13g2_buf_2 _08114_ (.A(_02627_),
    .X(_02711_));
 sg13g2_buf_1 _08115_ (.A(_02437_),
    .X(_02712_));
 sg13g2_nor2_1 _08116_ (.A(net120),
    .B(net295),
    .Y(_02713_));
 sg13g2_buf_1 _08117_ (.A(net311),
    .X(_02714_));
 sg13g2_o21ai_1 _08118_ (.B1(net195),
    .Y(_02715_),
    .A1(net196),
    .A2(_02713_));
 sg13g2_nand3_1 _08119_ (.B(net197),
    .C(_02715_),
    .A(net143),
    .Y(_02716_));
 sg13g2_buf_1 _08120_ (.A(net330),
    .X(_02717_));
 sg13g2_buf_1 _08121_ (.A(net194),
    .X(_02718_));
 sg13g2_nand2b_2 _08122_ (.Y(_02719_),
    .B(net389),
    .A_N(net381));
 sg13g2_buf_1 _08123_ (.A(net319),
    .X(_02720_));
 sg13g2_nor2_1 _08124_ (.A(net193),
    .B(net425),
    .Y(_02721_));
 sg13g2_a22oi_1 _08125_ (.Y(_02722_),
    .B1(_02721_),
    .B2(net195),
    .A2(_02719_),
    .A1(net239));
 sg13g2_nand2_1 _08126_ (.Y(_02723_),
    .A(net119),
    .B(_02722_));
 sg13g2_nand3_1 _08127_ (.B(_02716_),
    .C(_02723_),
    .A(net121),
    .Y(_02724_));
 sg13g2_buf_1 _08128_ (.A(net302),
    .X(_02725_));
 sg13g2_buf_1 _08129_ (.A(net192),
    .X(_02726_));
 sg13g2_nor2_2 _08130_ (.A(net331),
    .B(_01788_),
    .Y(_02727_));
 sg13g2_nor2_1 _08131_ (.A(net201),
    .B(_02727_),
    .Y(_02728_));
 sg13g2_nand3_1 _08132_ (.B(net89),
    .C(_02728_),
    .A(net118),
    .Y(_02729_));
 sg13g2_and3_1 _08133_ (.X(_02730_),
    .A(_01963_),
    .B(_02724_),
    .C(_02729_));
 sg13g2_nor2_1 _08134_ (.A(_02534_),
    .B(net232),
    .Y(_02731_));
 sg13g2_nand2_1 _08135_ (.Y(_02732_),
    .A(net393),
    .B(net327));
 sg13g2_nand2b_1 _08136_ (.Y(_02733_),
    .B(_01909_),
    .A_N(net380));
 sg13g2_nor2_1 _08137_ (.A(net327),
    .B(net467),
    .Y(_02734_));
 sg13g2_nor2_1 _08138_ (.A(_02733_),
    .B(_02734_),
    .Y(_02735_));
 sg13g2_a21oi_1 _08139_ (.A1(net121),
    .A2(_02732_),
    .Y(_02736_),
    .B1(_02735_));
 sg13g2_buf_1 _08140_ (.A(net237),
    .X(_02737_));
 sg13g2_a221oi_1 _08141_ (.B2(net141),
    .C1(net117),
    .B1(_02736_),
    .A1(_02456_),
    .Y(_02738_),
    .A2(_02731_));
 sg13g2_nor3_1 _08142_ (.A(net122),
    .B(_02730_),
    .C(_02738_),
    .Y(_02739_));
 sg13g2_nor2_1 _08143_ (.A(_02538_),
    .B(_02607_),
    .Y(_02740_));
 sg13g2_buf_1 _08144_ (.A(_02471_),
    .X(_02741_));
 sg13g2_nor2_1 _08145_ (.A(net116),
    .B(_02417_),
    .Y(_02742_));
 sg13g2_nor4_1 _08146_ (.A(net82),
    .B(net238),
    .C(_02740_),
    .D(_02742_),
    .Y(_02743_));
 sg13g2_buf_1 _08147_ (.A(_02469_),
    .X(_02744_));
 sg13g2_buf_1 _08148_ (.A(net294),
    .X(_02745_));
 sg13g2_nand2_1 _08149_ (.Y(_02746_),
    .A(net191),
    .B(net127));
 sg13g2_a21oi_1 _08150_ (.A1(net322),
    .A2(_02746_),
    .Y(_02747_),
    .B1(_01771_));
 sg13g2_buf_1 _08151_ (.A(_00092_),
    .X(_02748_));
 sg13g2_buf_1 _08152_ (.A(net459),
    .X(_02749_));
 sg13g2_buf_1 _08153_ (.A(net307),
    .X(_02750_));
 sg13g2_nor2b_1 _08154_ (.A(_01954_),
    .B_N(net379),
    .Y(_02751_));
 sg13g2_buf_1 _08155_ (.A(_02751_),
    .X(_02752_));
 sg13g2_a22oi_1 _08156_ (.Y(_02753_),
    .B1(net189),
    .B2(net425),
    .A2(net190),
    .A1(net211));
 sg13g2_nor3_1 _08157_ (.A(_02352_),
    .B(_02461_),
    .C(_02740_),
    .Y(_02754_));
 sg13g2_a21oi_1 _08158_ (.A1(net143),
    .A2(_02753_),
    .Y(_02755_),
    .B1(_02754_));
 sg13g2_buf_1 _08159_ (.A(net379),
    .X(_02756_));
 sg13g2_nor2_2 _08160_ (.A(net293),
    .B(net308),
    .Y(_02757_));
 sg13g2_nor3_1 _08161_ (.A(net420),
    .B(_02755_),
    .C(_02757_),
    .Y(_02758_));
 sg13g2_buf_1 _08162_ (.A(_01976_),
    .X(_02759_));
 sg13g2_buf_1 _08163_ (.A(net292),
    .X(_02760_));
 sg13g2_buf_1 _08164_ (.A(net212),
    .X(_02761_));
 sg13g2_o21ai_1 _08165_ (.B1(_02761_),
    .Y(_02762_),
    .A1(net195),
    .A2(_02423_));
 sg13g2_buf_1 _08166_ (.A(net200),
    .X(_02763_));
 sg13g2_nand2_1 _08167_ (.Y(_02764_),
    .A(net114),
    .B(net425));
 sg13g2_o21ai_1 _08168_ (.B1(_02764_),
    .Y(_02765_),
    .A1(net131),
    .A2(_02762_));
 sg13g2_nor2_1 _08169_ (.A(net315),
    .B(_02304_),
    .Y(_02766_));
 sg13g2_o21ai_1 _08170_ (.B1(net128),
    .Y(_02767_),
    .A1(_02514_),
    .A2(_02766_));
 sg13g2_nand3_1 _08171_ (.B(_02765_),
    .C(_02767_),
    .A(_02760_),
    .Y(_02768_));
 sg13g2_o21ai_1 _08172_ (.B1(_02768_),
    .Y(_02769_),
    .A1(net117),
    .A2(_02758_));
 sg13g2_nor4_1 _08173_ (.A(net134),
    .B(_02743_),
    .C(_02747_),
    .D(_02769_),
    .Y(_02770_));
 sg13g2_nor2b_1 _08174_ (.A(_02487_),
    .B_N(_02482_),
    .Y(_02771_));
 sg13g2_buf_1 _08175_ (.A(_02771_),
    .X(_02772_));
 sg13g2_nand2_2 _08176_ (.Y(_02773_),
    .A(_02603_),
    .B(_02772_));
 sg13g2_inv_1 _08177_ (.Y(_02774_),
    .A(_02773_));
 sg13g2_o21ai_1 _08178_ (.B1(_02774_),
    .Y(_02775_),
    .A1(_02739_),
    .A2(_02770_));
 sg13g2_and2_1 _08179_ (.A(_02495_),
    .B(_02502_),
    .X(_02776_));
 sg13g2_buf_1 _08180_ (.A(_02776_),
    .X(_02777_));
 sg13g2_and2_1 _08181_ (.A(_02777_),
    .B(_02772_),
    .X(_02778_));
 sg13g2_buf_2 _08182_ (.A(_02778_),
    .X(_02779_));
 sg13g2_nor2b_1 _08183_ (.A(_01765_),
    .B_N(net467),
    .Y(_02780_));
 sg13g2_buf_1 _08184_ (.A(_02780_),
    .X(_02781_));
 sg13g2_nor2_2 _08185_ (.A(net391),
    .B(_02781_),
    .Y(_02782_));
 sg13g2_nand3_1 _08186_ (.B(_02535_),
    .C(_02782_),
    .A(net235),
    .Y(_02783_));
 sg13g2_a21oi_1 _08187_ (.A1(_02636_),
    .A2(_02783_),
    .Y(_02784_),
    .B1(_02703_));
 sg13g2_nand2_1 _08188_ (.Y(_02785_),
    .A(_02289_),
    .B(_02511_));
 sg13g2_nand2_1 _08189_ (.Y(_02786_),
    .A(net340),
    .B(_02544_));
 sg13g2_nor2_1 _08190_ (.A(_01929_),
    .B(net467),
    .Y(_02787_));
 sg13g2_buf_1 _08191_ (.A(_02787_),
    .X(_02788_));
 sg13g2_a21oi_1 _08192_ (.A1(net187),
    .A2(net196),
    .Y(_02789_),
    .B1(_02408_));
 sg13g2_a22oi_1 _08193_ (.Y(_02790_),
    .B1(_02786_),
    .B2(_02789_),
    .A2(_02785_),
    .A1(net246));
 sg13g2_buf_1 _08194_ (.A(net391),
    .X(_02791_));
 sg13g2_buf_1 _08195_ (.A(net291),
    .X(_02792_));
 sg13g2_a221oi_1 _08196_ (.B2(net234),
    .C1(net314),
    .B1(_02535_),
    .A1(_02644_),
    .Y(_02793_),
    .A2(net187));
 sg13g2_a21oi_1 _08197_ (.A1(net186),
    .A2(_02665_),
    .Y(_02794_),
    .B1(_02793_));
 sg13g2_nor2_2 _08198_ (.A(_00091_),
    .B(_02432_),
    .Y(_02795_));
 sg13g2_a22oi_1 _08199_ (.Y(_02796_),
    .B1(_02794_),
    .B2(_02795_),
    .A2(_02790_),
    .A1(_02784_));
 sg13g2_inv_1 _08200_ (.Y(_02797_),
    .A(_02796_));
 sg13g2_nor2_1 _08201_ (.A(net474),
    .B(net460),
    .Y(_02798_));
 sg13g2_buf_2 _08202_ (.A(_02798_),
    .X(_02799_));
 sg13g2_nand2b_1 _08203_ (.Y(_02800_),
    .B(_02799_),
    .A_N(_00091_));
 sg13g2_buf_1 _08204_ (.A(_02800_),
    .X(_02801_));
 sg13g2_a22oi_1 _08205_ (.Y(_02802_),
    .B1(_02544_),
    .B2(_01887_),
    .A2(net213),
    .A1(net295));
 sg13g2_buf_1 _08206_ (.A(net296),
    .X(_02803_));
 sg13g2_nand2_1 _08207_ (.Y(_02804_),
    .A(_02373_),
    .B(_02375_));
 sg13g2_nor2_1 _08208_ (.A(net184),
    .B(_02804_),
    .Y(_02805_));
 sg13g2_a21oi_1 _08209_ (.A1(net217),
    .A2(_02802_),
    .Y(_02806_),
    .B1(_02805_));
 sg13g2_nand2_1 _08210_ (.Y(_02807_),
    .A(net192),
    .B(_02786_));
 sg13g2_o21ai_1 _08211_ (.B1(_02807_),
    .Y(_02808_),
    .A1(net219),
    .A2(_02806_));
 sg13g2_nand2_1 _08212_ (.Y(_02809_),
    .A(net384),
    .B(net440));
 sg13g2_buf_1 _08213_ (.A(_02809_),
    .X(_02810_));
 sg13g2_nor2_1 _08214_ (.A(net296),
    .B(net183),
    .Y(_02811_));
 sg13g2_buf_2 _08215_ (.A(_00093_),
    .X(_02812_));
 sg13g2_nor3_1 _08216_ (.A(_01935_),
    .B(net433),
    .C(_02812_),
    .Y(_02813_));
 sg13g2_a22oi_1 _08217_ (.Y(_02814_),
    .B1(_02813_),
    .B2(net125),
    .A2(_02811_),
    .A1(net302));
 sg13g2_nor2_1 _08218_ (.A(net336),
    .B(_02814_),
    .Y(_02815_));
 sg13g2_buf_1 _08219_ (.A(_01916_),
    .X(_02816_));
 sg13g2_nand2_1 _08220_ (.Y(_02817_),
    .A(_02332_),
    .B(_02612_));
 sg13g2_buf_1 _08221_ (.A(_02817_),
    .X(_02818_));
 sg13g2_nor2_1 _08222_ (.A(net182),
    .B(net113),
    .Y(_02819_));
 sg13g2_nor2_1 _08223_ (.A(_02360_),
    .B(net248),
    .Y(_02820_));
 sg13g2_and2_1 _08224_ (.A(_02819_),
    .B(_02820_),
    .X(_02821_));
 sg13g2_nor2_1 _08225_ (.A(_02428_),
    .B(_01753_),
    .Y(_02822_));
 sg13g2_buf_1 _08226_ (.A(_02822_),
    .X(_02823_));
 sg13g2_buf_1 _08227_ (.A(_02823_),
    .X(_02824_));
 sg13g2_o21ai_1 _08228_ (.B1(net181),
    .Y(_02825_),
    .A1(_02815_),
    .A2(_02821_));
 sg13g2_o21ai_1 _08229_ (.B1(_02825_),
    .Y(_02826_),
    .A1(_02801_),
    .A2(_02808_));
 sg13g2_and2_1 _08230_ (.A(_02503_),
    .B(_02772_),
    .X(_02827_));
 sg13g2_buf_2 _08231_ (.A(_02827_),
    .X(_02828_));
 sg13g2_a22oi_1 _08232_ (.Y(_02829_),
    .B1(_02826_),
    .B2(_02828_),
    .A2(_02797_),
    .A1(_02779_));
 sg13g2_buf_1 _08233_ (.A(_02799_),
    .X(_02830_));
 sg13g2_nand3b_1 _08234_ (.B(net439),
    .C(net437),
    .Y(_02831_),
    .A_N(net435));
 sg13g2_buf_1 _08235_ (.A(_02831_),
    .X(_02832_));
 sg13g2_a21oi_1 _08236_ (.A1(_02832_),
    .A2(_02558_),
    .Y(_02833_),
    .B1(net193));
 sg13g2_nor3_1 _08237_ (.A(net234),
    .B(net196),
    .C(_02833_),
    .Y(_02834_));
 sg13g2_nor2_1 _08238_ (.A(net422),
    .B(net304),
    .Y(_02835_));
 sg13g2_inv_1 _08239_ (.Y(_02836_),
    .A(net459));
 sg13g2_o21ai_1 _08240_ (.B1(_02836_),
    .Y(_02837_),
    .A1(net241),
    .A2(_02835_));
 sg13g2_o21ai_1 _08241_ (.B1(net202),
    .Y(_02838_),
    .A1(_02834_),
    .A2(_02837_));
 sg13g2_buf_1 _08242_ (.A(net182),
    .X(_02839_));
 sg13g2_a21oi_1 _08243_ (.A1(net182),
    .A2(_02564_),
    .Y(_02840_),
    .B1(net341));
 sg13g2_o21ai_1 _08244_ (.B1(_02840_),
    .Y(_02841_),
    .A1(net197),
    .A2(net112));
 sg13g2_buf_1 _08245_ (.A(_01955_),
    .X(_02842_));
 sg13g2_nand2b_1 _08246_ (.Y(_02843_),
    .B(net428),
    .A_N(_01781_));
 sg13g2_buf_1 _08247_ (.A(_02843_),
    .X(_02844_));
 sg13g2_buf_1 _08248_ (.A(_02844_),
    .X(_02845_));
 sg13g2_nand3b_1 _08249_ (.B(net440),
    .C(net437),
    .Y(_02846_),
    .A_N(net435));
 sg13g2_buf_2 _08250_ (.A(_02846_),
    .X(_02847_));
 sg13g2_nand2_1 _08251_ (.Y(_02848_),
    .A(net180),
    .B(_02847_));
 sg13g2_buf_1 _08252_ (.A(_02441_),
    .X(_02849_));
 sg13g2_nand2b_1 _08253_ (.Y(_02850_),
    .B(net440),
    .A_N(_02294_));
 sg13g2_buf_1 _08254_ (.A(_02850_),
    .X(_02851_));
 sg13g2_buf_1 _08255_ (.A(_02851_),
    .X(_02852_));
 sg13g2_nor2_1 _08256_ (.A(net288),
    .B(net179),
    .Y(_02853_));
 sg13g2_a221oi_1 _08257_ (.B2(_02803_),
    .C1(_02853_),
    .B1(_02848_),
    .A1(net289),
    .Y(_02854_),
    .A2(_02356_));
 sg13g2_a21oi_1 _08258_ (.A1(net153),
    .A2(_02447_),
    .Y(_02855_),
    .B1(net325));
 sg13g2_o21ai_1 _08259_ (.B1(_02855_),
    .Y(_02856_),
    .A1(net145),
    .A2(_02854_));
 sg13g2_and4_1 _08260_ (.A(net290),
    .B(_02838_),
    .C(_02841_),
    .D(_02856_),
    .X(_02857_));
 sg13g2_nor2_1 _08261_ (.A(_01765_),
    .B(net428),
    .Y(_02858_));
 sg13g2_and2_1 _08262_ (.A(_02576_),
    .B(_02858_),
    .X(_02859_));
 sg13g2_buf_1 _08263_ (.A(_02859_),
    .X(_02860_));
 sg13g2_nor2_1 _08264_ (.A(_02445_),
    .B(_02860_),
    .Y(_02861_));
 sg13g2_nor2b_1 _08265_ (.A(_01897_),
    .B_N(_01895_),
    .Y(_02862_));
 sg13g2_buf_2 _08266_ (.A(_02862_),
    .X(_02863_));
 sg13g2_nand2_2 _08267_ (.Y(_02864_),
    .A(net394),
    .B(_02335_));
 sg13g2_nand3_1 _08268_ (.B(_02863_),
    .C(_02864_),
    .A(net184),
    .Y(_02865_));
 sg13g2_o21ai_1 _08269_ (.B1(_02865_),
    .Y(_02866_),
    .A1(net218),
    .A2(net197));
 sg13g2_buf_1 _08270_ (.A(_01976_),
    .X(_02867_));
 sg13g2_buf_1 _08271_ (.A(_02781_),
    .X(_02868_));
 sg13g2_or2_1 _08272_ (.X(_02869_),
    .B(net440),
    .A(net435));
 sg13g2_buf_1 _08273_ (.A(_02869_),
    .X(_02870_));
 sg13g2_buf_1 _08274_ (.A(_02870_),
    .X(_02871_));
 sg13g2_nand3_1 _08275_ (.B(net286),
    .C(net178),
    .A(net137),
    .Y(_02872_));
 sg13g2_nand2_1 _08276_ (.Y(_02873_),
    .A(net287),
    .B(_02872_));
 sg13g2_o21ai_1 _08277_ (.B1(_02873_),
    .Y(_02874_),
    .A1(net136),
    .A2(_02866_));
 sg13g2_nand2b_1 _08278_ (.Y(_02875_),
    .B(_02298_),
    .A_N(net461));
 sg13g2_and3_1 _08279_ (.X(_02876_),
    .A(net294),
    .B(_01899_),
    .C(_02875_));
 sg13g2_mux2_1 _08280_ (.A0(net462),
    .A1(net461),
    .S(net384),
    .X(_02877_));
 sg13g2_and2_1 _08281_ (.A(net342),
    .B(_02877_),
    .X(_02878_));
 sg13g2_nor2_1 _08282_ (.A(_02876_),
    .B(_02878_),
    .Y(_02879_));
 sg13g2_a221oi_1 _08283_ (.B2(_02342_),
    .C1(_02361_),
    .B1(_02879_),
    .A1(net129),
    .Y(_02880_),
    .A2(_02521_));
 sg13g2_nor4_1 _08284_ (.A(net198),
    .B(_02861_),
    .C(_02874_),
    .D(_02880_),
    .Y(_02881_));
 sg13g2_and2_1 _08285_ (.A(_02777_),
    .B(_02489_),
    .X(_02882_));
 sg13g2_buf_2 _08286_ (.A(_02882_),
    .X(_02883_));
 sg13g2_o21ai_1 _08287_ (.B1(_02883_),
    .Y(_02884_),
    .A1(_02857_),
    .A2(_02881_));
 sg13g2_nand2_1 _08288_ (.Y(_02885_),
    .A(_02829_),
    .B(_02884_));
 sg13g2_nand2_1 _08289_ (.Y(_02886_),
    .A(_02772_),
    .B(_02595_));
 sg13g2_buf_2 _08290_ (.A(_02886_),
    .X(_02887_));
 sg13g2_nand2_1 _08291_ (.Y(_02888_),
    .A(net112),
    .B(net129));
 sg13g2_buf_1 _08292_ (.A(net329),
    .X(_02889_));
 sg13g2_nor2_1 _08293_ (.A(net177),
    .B(net130),
    .Y(_02890_));
 sg13g2_and2_1 _08294_ (.A(net443),
    .B(net381),
    .X(_02891_));
 sg13g2_buf_1 _08295_ (.A(_02891_),
    .X(_02892_));
 sg13g2_a22oi_1 _08296_ (.Y(_02893_),
    .B1(net306),
    .B2(_02892_),
    .A2(_02890_),
    .A1(net239));
 sg13g2_a221oi_1 _08297_ (.B2(_02759_),
    .C1(net229),
    .B1(_02893_),
    .A1(_02671_),
    .Y(_02894_),
    .A2(_02888_));
 sg13g2_buf_1 _08298_ (.A(_02863_),
    .X(_02895_));
 sg13g2_nand2_1 _08299_ (.Y(_02896_),
    .A(net208),
    .B(_02684_));
 sg13g2_nand2_1 _08300_ (.Y(_02897_),
    .A(_02284_),
    .B(_02612_));
 sg13g2_a21oi_1 _08301_ (.A1(_02896_),
    .A2(_02897_),
    .Y(_02898_),
    .B1(net240));
 sg13g2_a221oi_1 _08302_ (.B2(_02835_),
    .C1(_02898_),
    .B1(net321),
    .A1(net155),
    .Y(_02899_),
    .A2(_02895_));
 sg13g2_buf_1 _08303_ (.A(net382),
    .X(_02900_));
 sg13g2_buf_1 _08304_ (.A(_02900_),
    .X(_02901_));
 sg13g2_o21ai_1 _08305_ (.B1(net175),
    .Y(_02902_),
    .A1(net420),
    .A2(_02899_));
 sg13g2_buf_1 _08306_ (.A(_02417_),
    .X(_02903_));
 sg13g2_o21ai_1 _08307_ (.B1(net89),
    .Y(_02904_),
    .A1(net196),
    .A2(_02721_));
 sg13g2_a21oi_1 _08308_ (.A1(net227),
    .A2(_02875_),
    .Y(_02905_),
    .B1(net224));
 sg13g2_o21ai_1 _08309_ (.B1(net320),
    .Y(_02906_),
    .A1(net130),
    .A2(net190));
 sg13g2_and2_1 _08310_ (.A(net384),
    .B(net379),
    .X(_02907_));
 sg13g2_buf_1 _08311_ (.A(_02907_),
    .X(_02908_));
 sg13g2_buf_1 _08312_ (.A(_02908_),
    .X(_02909_));
 sg13g2_nor2_1 _08313_ (.A(_02294_),
    .B(net440),
    .Y(_02910_));
 sg13g2_buf_1 _08314_ (.A(_02910_),
    .X(_02911_));
 sg13g2_a21oi_1 _08315_ (.A1(net235),
    .A2(net110),
    .Y(_02912_),
    .B1(net284));
 sg13g2_o21ai_1 _08316_ (.B1(net215),
    .Y(_02913_),
    .A1(net244),
    .A2(_02912_));
 sg13g2_o21ai_1 _08317_ (.B1(_02913_),
    .Y(_02914_),
    .A1(_02905_),
    .A2(_02906_));
 sg13g2_a221oi_1 _08318_ (.B2(net188),
    .C1(_02914_),
    .B1(_02904_),
    .A1(net111),
    .Y(_02915_),
    .A2(_02566_));
 sg13g2_buf_1 _08319_ (.A(net181),
    .X(_02916_));
 sg13g2_a22oi_1 _08320_ (.Y(_02917_),
    .B1(_02915_),
    .B2(net109),
    .A2(_02902_),
    .A1(_02894_));
 sg13g2_and2_1 _08321_ (.A(_02482_),
    .B(_02487_),
    .X(_02918_));
 sg13g2_a21oi_2 _08322_ (.B1(_02918_),
    .Y(_02919_),
    .A2(_02663_),
    .A1(_02496_));
 sg13g2_buf_1 _08323_ (.A(_02919_),
    .X(_02920_));
 sg13g2_o21ai_1 _08324_ (.B1(net59),
    .Y(_02921_),
    .A1(_02887_),
    .A2(_02917_));
 sg13g2_buf_1 _08325_ (.A(_02824_),
    .X(_02922_));
 sg13g2_buf_1 _08326_ (.A(_02509_),
    .X(_02923_));
 sg13g2_buf_1 _08327_ (.A(net283),
    .X(_02924_));
 sg13g2_o21ai_1 _08328_ (.B1(net113),
    .Y(_02925_),
    .A1(_01957_),
    .A2(_02924_));
 sg13g2_nor2_1 _08329_ (.A(_02288_),
    .B(_02844_),
    .Y(_02926_));
 sg13g2_nor2_1 _08330_ (.A(net384),
    .B(_02509_),
    .Y(_02927_));
 sg13g2_buf_1 _08331_ (.A(_02927_),
    .X(_02928_));
 sg13g2_a21oi_2 _08332_ (.B1(_02928_),
    .Y(_02929_),
    .A2(_02926_),
    .A1(_01886_));
 sg13g2_nand2_1 _08333_ (.Y(_02930_),
    .A(net303),
    .B(_02929_));
 sg13g2_o21ai_1 _08334_ (.B1(_02930_),
    .Y(_02931_),
    .A1(net199),
    .A2(net201));
 sg13g2_nor2_1 _08335_ (.A(_02366_),
    .B(_02931_),
    .Y(_02932_));
 sg13g2_a21oi_1 _08336_ (.A1(net149),
    .A2(_02925_),
    .Y(_02933_),
    .B1(_02932_));
 sg13g2_nand3_1 _08337_ (.B(_01957_),
    .C(net113),
    .A(net237),
    .Y(_02934_));
 sg13g2_nor2_1 _08338_ (.A(net372),
    .B(net201),
    .Y(_02935_));
 sg13g2_nand2_1 _08339_ (.Y(_02936_),
    .A(net431),
    .B(net212));
 sg13g2_nor2_1 _08340_ (.A(_02379_),
    .B(_02936_),
    .Y(_02937_));
 sg13g2_o21ai_1 _08341_ (.B1(_02726_),
    .Y(_02938_),
    .A1(_02935_),
    .A2(_02937_));
 sg13g2_buf_1 _08342_ (.A(_02928_),
    .X(_02939_));
 sg13g2_a21oi_1 _08343_ (.A1(net155),
    .A2(_02696_),
    .Y(_02940_),
    .B1(net107));
 sg13g2_a21oi_1 _08344_ (.A1(net107),
    .A2(_02521_),
    .Y(_02941_),
    .B1(net136));
 sg13g2_o21ai_1 _08345_ (.B1(_02941_),
    .Y(_02942_),
    .A1(net152),
    .A2(_02940_));
 sg13g2_nand4_1 _08346_ (.B(_02934_),
    .C(_02938_),
    .A(_02430_),
    .Y(_02943_),
    .D(_02942_));
 sg13g2_buf_1 _08347_ (.A(net115),
    .X(_02944_));
 sg13g2_nand2_2 _08348_ (.Y(_02945_),
    .A(net378),
    .B(net213));
 sg13g2_a21oi_1 _08349_ (.A1(net81),
    .A2(_02945_),
    .Y(_02946_),
    .B1(_02322_));
 sg13g2_nand2_1 _08350_ (.Y(_02947_),
    .A(_02663_),
    .B(_02777_));
 sg13g2_inv_1 _08351_ (.Y(_02948_),
    .A(_02947_));
 sg13g2_o21ai_1 _08352_ (.B1(_02948_),
    .Y(_02949_),
    .A1(net386),
    .A2(_02946_));
 sg13g2_a221oi_1 _08353_ (.B2(net316),
    .C1(_02949_),
    .B1(_02943_),
    .A1(net108),
    .Y(_02950_),
    .A2(_02933_));
 sg13g2_nor3_1 _08354_ (.A(_02885_),
    .B(_02921_),
    .C(_02950_),
    .Y(_02951_));
 sg13g2_nand4_1 _08355_ (.B(_02701_),
    .C(_02775_),
    .A(_02598_),
    .Y(_02952_),
    .D(_02951_));
 sg13g2_a21oi_2 _08356_ (.B1(net386),
    .Y(_02953_),
    .A2(_02696_),
    .A1(net60));
 sg13g2_nor2_1 _08357_ (.A(net391),
    .B(net338),
    .Y(_02954_));
 sg13g2_buf_1 _08358_ (.A(_02954_),
    .X(_02955_));
 sg13g2_a22oi_1 _08359_ (.Y(_02956_),
    .B1(_02818_),
    .B2(net106),
    .A2(net124),
    .A1(net150));
 sg13g2_inv_1 _08360_ (.Y(_02957_),
    .A(_02956_));
 sg13g2_a21o_1 _08361_ (.A2(net124),
    .A1(_02365_),
    .B1(_02935_),
    .X(_02958_));
 sg13g2_a221oi_1 _08362_ (.B2(net132),
    .C1(_02530_),
    .B1(_02958_),
    .A1(net237),
    .Y(_02959_),
    .A2(_02957_));
 sg13g2_nand2_1 _08363_ (.Y(_02960_),
    .A(net217),
    .B(_02746_));
 sg13g2_o21ai_1 _08364_ (.B1(_02941_),
    .Y(_02961_),
    .A1(net174),
    .A2(_02960_));
 sg13g2_a21oi_1 _08365_ (.A1(_02959_),
    .A2(_02961_),
    .Y(_02962_),
    .B1(net444));
 sg13g2_buf_1 _08366_ (.A(net387),
    .X(_02963_));
 sg13g2_a21o_1 _08367_ (.A2(_02682_),
    .A1(net253),
    .B1(_02963_),
    .X(_02964_));
 sg13g2_inv_1 _08368_ (.Y(_02965_),
    .A(_02964_));
 sg13g2_a21oi_1 _08369_ (.A1(net139),
    .A2(_02860_),
    .Y(_02966_),
    .B1(_02965_));
 sg13g2_buf_1 _08370_ (.A(net107),
    .X(_02967_));
 sg13g2_nand2_1 _08371_ (.Y(_02968_),
    .A(net249),
    .B(net80));
 sg13g2_nand3_1 _08372_ (.B(_02655_),
    .C(_02568_),
    .A(_02693_),
    .Y(_02969_));
 sg13g2_and3_1 _08373_ (.X(_02970_),
    .A(net123),
    .B(_02968_),
    .C(_02969_));
 sg13g2_a21oi_1 _08374_ (.A1(net140),
    .A2(_02966_),
    .Y(_02971_),
    .B1(_02970_));
 sg13g2_nor2_1 _08375_ (.A(net122),
    .B(_02971_),
    .Y(_02972_));
 sg13g2_nor3_1 _08376_ (.A(_02953_),
    .B(_02962_),
    .C(_02972_),
    .Y(_02973_));
 sg13g2_or2_1 _08377_ (.X(_02974_),
    .B(_02973_),
    .A(net59));
 sg13g2_o21ai_1 _08378_ (.B1(_02974_),
    .Y(_02975_),
    .A1(_02505_),
    .A2(_02952_));
 sg13g2_nor2_1 _08379_ (.A(net310),
    .B(_02727_),
    .Y(_02976_));
 sg13g2_a21oi_1 _08380_ (.A1(_02402_),
    .A2(_02976_),
    .Y(_02977_),
    .B1(_01983_));
 sg13g2_nor2_1 _08381_ (.A(_02596_),
    .B(_02977_),
    .Y(_02978_));
 sg13g2_nand2_1 _08382_ (.Y(_02979_),
    .A(net333),
    .B(net178));
 sg13g2_o21ai_1 _08383_ (.B1(net313),
    .Y(_02980_),
    .A1(net342),
    .A2(net183));
 sg13g2_a21oi_1 _08384_ (.A1(_02832_),
    .A2(_02979_),
    .Y(_02981_),
    .B1(_02980_));
 sg13g2_nor2_1 _08385_ (.A(net341),
    .B(_02981_),
    .Y(_02982_));
 sg13g2_buf_1 _08386_ (.A(net208),
    .X(_02983_));
 sg13g2_nand2_1 _08387_ (.Y(_02984_),
    .A(_02650_),
    .B(_02983_));
 sg13g2_nor2_1 _08388_ (.A(net230),
    .B(net251),
    .Y(_02985_));
 sg13g2_a21oi_1 _08389_ (.A1(net218),
    .A2(net204),
    .Y(_02986_),
    .B1(_02985_));
 sg13g2_o21ai_1 _08390_ (.B1(_02680_),
    .Y(_02987_),
    .A1(_02984_),
    .A2(_02986_));
 sg13g2_buf_1 _08391_ (.A(net220),
    .X(_02988_));
 sg13g2_nor2_2 _08392_ (.A(net294),
    .B(_02587_),
    .Y(_02989_));
 sg13g2_nor2_1 _08393_ (.A(net384),
    .B(_02421_),
    .Y(_02990_));
 sg13g2_buf_2 _08394_ (.A(_02990_),
    .X(_02991_));
 sg13g2_buf_1 _08395_ (.A(_02991_),
    .X(_02992_));
 sg13g2_o21ai_1 _08396_ (.B1(net116),
    .Y(_02993_),
    .A1(net374),
    .A2(net79));
 sg13g2_buf_1 _08397_ (.A(_02341_),
    .X(_02994_));
 sg13g2_nand2_1 _08398_ (.Y(_02995_),
    .A(net282),
    .B(net133));
 sg13g2_a221oi_1 _08399_ (.B2(net103),
    .C1(_02995_),
    .B1(_02993_),
    .A1(net104),
    .Y(_02996_),
    .A2(_02989_));
 sg13g2_nor2_1 _08400_ (.A(_02987_),
    .B(_02996_),
    .Y(_02997_));
 sg13g2_a221oi_1 _08401_ (.B2(_02945_),
    .C1(_02997_),
    .B1(_02982_),
    .A1(_02818_),
    .Y(_02998_),
    .A2(_02820_));
 sg13g2_nor2_1 _08402_ (.A(_02361_),
    .B(_02545_),
    .Y(_02999_));
 sg13g2_o21ai_1 _08403_ (.B1(net82),
    .Y(_03000_),
    .A1(_02982_),
    .A2(_02999_));
 sg13g2_a21o_1 _08404_ (.A2(_03000_),
    .A1(_02998_),
    .B1(net122),
    .X(_03001_));
 sg13g2_o21ai_1 _08405_ (.B1(net377),
    .Y(_03002_),
    .A1(net381),
    .A2(_02844_));
 sg13g2_buf_1 _08406_ (.A(_03002_),
    .X(_03003_));
 sg13g2_a21oi_1 _08407_ (.A1(net383),
    .A2(net462),
    .Y(_03004_),
    .B1(net377));
 sg13g2_buf_2 _08408_ (.A(_03004_),
    .X(_03005_));
 sg13g2_a21oi_1 _08409_ (.A1(net116),
    .A2(net102),
    .Y(_03006_),
    .B1(_03005_));
 sg13g2_nor2_1 _08410_ (.A(_02322_),
    .B(_03006_),
    .Y(_03007_));
 sg13g2_nor2_1 _08411_ (.A(_01984_),
    .B(_03007_),
    .Y(_03008_));
 sg13g2_nor2_1 _08412_ (.A(_02504_),
    .B(_03008_),
    .Y(_03009_));
 sg13g2_buf_1 _08413_ (.A(_02637_),
    .X(_03010_));
 sg13g2_nor2_1 _08414_ (.A(net394),
    .B(_02347_),
    .Y(_03011_));
 sg13g2_buf_2 _08415_ (.A(_03011_),
    .X(_03012_));
 sg13g2_nand2b_1 _08416_ (.Y(_03013_),
    .B(net437),
    .A_N(_01782_));
 sg13g2_buf_2 _08417_ (.A(_03013_),
    .X(_03014_));
 sg13g2_nor2_1 _08418_ (.A(_02389_),
    .B(_03014_),
    .Y(_03015_));
 sg13g2_a21oi_1 _08419_ (.A1(net133),
    .A2(_03012_),
    .Y(_03016_),
    .B1(_03015_));
 sg13g2_nand2_1 _08420_ (.Y(_03017_),
    .A(net172),
    .B(_03016_));
 sg13g2_nand3_1 _08421_ (.B(net154),
    .C(_02852_),
    .A(net175),
    .Y(_03018_));
 sg13g2_nand2b_1 _08422_ (.Y(_03019_),
    .B(_01884_),
    .A_N(net435));
 sg13g2_buf_1 _08423_ (.A(_03019_),
    .X(_03020_));
 sg13g2_nor2b_1 _08424_ (.A(net443),
    .B_N(net434),
    .Y(_03021_));
 sg13g2_buf_1 _08425_ (.A(_03021_),
    .X(_03022_));
 sg13g2_buf_1 _08426_ (.A(_03022_),
    .X(_03023_));
 sg13g2_o21ai_1 _08427_ (.B1(net171),
    .Y(_03024_),
    .A1(net197),
    .A2(net281));
 sg13g2_a21oi_1 _08428_ (.A1(_03017_),
    .A2(_03018_),
    .Y(_03025_),
    .B1(_03024_));
 sg13g2_nand2_1 _08429_ (.Y(_03026_),
    .A(net153),
    .B(net196));
 sg13g2_nor2_1 _08430_ (.A(net340),
    .B(net306),
    .Y(_03027_));
 sg13g2_buf_1 _08431_ (.A(_02628_),
    .X(_03028_));
 sg13g2_nor2_1 _08432_ (.A(net317),
    .B(net427),
    .Y(_03029_));
 sg13g2_a21oi_1 _08433_ (.A1(net194),
    .A2(_03029_),
    .Y(_03030_),
    .B1(net189));
 sg13g2_nor2_1 _08434_ (.A(net78),
    .B(_03030_),
    .Y(_03031_));
 sg13g2_o21ai_1 _08435_ (.B1(net126),
    .Y(_03032_),
    .A1(_03027_),
    .A2(_03031_));
 sg13g2_nand3_1 _08436_ (.B(_03026_),
    .C(_03032_),
    .A(net215),
    .Y(_03033_));
 sg13g2_nand2_1 _08437_ (.Y(_03034_),
    .A(net227),
    .B(_02832_));
 sg13g2_nor2_1 _08438_ (.A(net468),
    .B(net385),
    .Y(_03035_));
 sg13g2_nand2_1 _08439_ (.Y(_03036_),
    .A(net434),
    .B(net443));
 sg13g2_buf_1 _08440_ (.A(_03036_),
    .X(_03037_));
 sg13g2_a221oi_1 _08441_ (.B2(net378),
    .C1(_03037_),
    .B1(_03035_),
    .A1(net431),
    .Y(_03038_),
    .A2(_03034_));
 sg13g2_a21oi_1 _08442_ (.A1(net208),
    .A2(_02719_),
    .Y(_03039_),
    .B1(net431));
 sg13g2_o21ai_1 _08443_ (.B1(net220),
    .Y(_03040_),
    .A1(net221),
    .A2(_03039_));
 sg13g2_o21ai_1 _08444_ (.B1(net377),
    .Y(_03041_),
    .A1(net296),
    .A2(net329));
 sg13g2_a221oi_1 _08445_ (.B2(net220),
    .C1(net325),
    .B1(_03041_),
    .A1(net127),
    .Y(_03042_),
    .A2(net378));
 sg13g2_a21oi_1 _08446_ (.A1(_03038_),
    .A2(_03040_),
    .Y(_03043_),
    .B1(_03042_));
 sg13g2_nand2_1 _08447_ (.Y(_03044_),
    .A(_03033_),
    .B(_03043_));
 sg13g2_o21ai_1 _08448_ (.B1(_01913_),
    .Y(_03045_),
    .A1(_03025_),
    .A2(_03044_));
 sg13g2_a22oi_1 _08449_ (.Y(_03046_),
    .B1(_03009_),
    .B2(_03045_),
    .A2(_03001_),
    .A1(_02978_));
 sg13g2_nand2_1 _08450_ (.Y(_03047_),
    .A(_02369_),
    .B(_02570_));
 sg13g2_o21ai_1 _08451_ (.B1(_03047_),
    .Y(_03048_),
    .A1(_02369_),
    .A2(net104));
 sg13g2_nand2_1 _08452_ (.Y(_03049_),
    .A(net245),
    .B(_03048_));
 sg13g2_o21ai_1 _08453_ (.B1(net199),
    .Y(_03050_),
    .A1(_01926_),
    .A2(net141));
 sg13g2_nor2_1 _08454_ (.A(_02624_),
    .B(_02517_),
    .Y(_03051_));
 sg13g2_buf_1 _08455_ (.A(_03051_),
    .X(_03052_));
 sg13g2_nor2_1 _08456_ (.A(_02638_),
    .B(net101),
    .Y(_03053_));
 sg13g2_o21ai_1 _08457_ (.B1(net132),
    .Y(_03054_),
    .A1(_02909_),
    .A2(net187));
 sg13g2_nand4_1 _08458_ (.B(_03050_),
    .C(_03053_),
    .A(_03049_),
    .Y(_03055_),
    .D(_03054_));
 sg13g2_nor3_1 _08459_ (.A(net339),
    .B(net115),
    .C(net187),
    .Y(_03056_));
 sg13g2_a22oi_1 _08460_ (.Y(_03057_),
    .B1(_02742_),
    .B2(_02353_),
    .A2(_02565_),
    .A1(_02647_));
 sg13g2_nor2_1 _08461_ (.A(net121),
    .B(_03057_),
    .Y(_03058_));
 sg13g2_o21ai_1 _08462_ (.B1(_02367_),
    .Y(_03059_),
    .A1(_03056_),
    .A2(_03058_));
 sg13g2_a21oi_1 _08463_ (.A1(_03055_),
    .A2(_03059_),
    .Y(_03060_),
    .B1(net424));
 sg13g2_a21oi_1 _08464_ (.A1(_02978_),
    .A2(_03060_),
    .Y(_03061_),
    .B1(net400));
 sg13g2_nand2_1 _08465_ (.Y(_03062_),
    .A(net295),
    .B(net335));
 sg13g2_nor2_1 _08466_ (.A(net333),
    .B(_02441_),
    .Y(_03063_));
 sg13g2_nand2_1 _08467_ (.Y(_03064_),
    .A(net110),
    .B(_03063_));
 sg13g2_nor2_1 _08468_ (.A(_02586_),
    .B(_02463_),
    .Y(_03065_));
 sg13g2_buf_2 _08469_ (.A(_03065_),
    .X(_03066_));
 sg13g2_nand2_1 _08470_ (.Y(_03067_),
    .A(net214),
    .B(_03066_));
 sg13g2_nand4_1 _08471_ (.B(_03062_),
    .C(_03064_),
    .A(net287),
    .Y(_03068_),
    .D(_03067_));
 sg13g2_nand2_1 _08472_ (.Y(_03069_),
    .A(net296),
    .B(_03066_));
 sg13g2_o21ai_1 _08473_ (.B1(net243),
    .Y(_03070_),
    .A1(net327),
    .A2(_02870_));
 sg13g2_nand2_1 _08474_ (.Y(_03071_),
    .A(net318),
    .B(_03070_));
 sg13g2_nand4_1 _08475_ (.B(_02653_),
    .C(_03069_),
    .A(net399),
    .Y(_03072_),
    .D(_03071_));
 sg13g2_nand3_1 _08476_ (.B(_03068_),
    .C(_03072_),
    .A(_02799_),
    .Y(_03073_));
 sg13g2_inv_1 _08477_ (.Y(_03074_),
    .A(_03073_));
 sg13g2_nor2_1 _08478_ (.A(net384),
    .B(net439),
    .Y(_03075_));
 sg13g2_buf_1 _08479_ (.A(_03075_),
    .X(_03076_));
 sg13g2_nand2_2 _08480_ (.Y(_03077_),
    .A(net422),
    .B(net170));
 sg13g2_nor2_1 _08481_ (.A(net254),
    .B(_03077_),
    .Y(_03078_));
 sg13g2_a21oi_1 _08482_ (.A1(net195),
    .A2(_02757_),
    .Y(_03079_),
    .B1(_03078_));
 sg13g2_nor2_1 _08483_ (.A(net390),
    .B(net295),
    .Y(_03080_));
 sg13g2_a221oi_1 _08484_ (.B2(net231),
    .C1(net420),
    .B1(_03080_),
    .A1(net142),
    .Y(_03081_),
    .A2(_03079_));
 sg13g2_a22oi_1 _08485_ (.Y(_03082_),
    .B1(_02333_),
    .B2(_02618_),
    .A2(net214),
    .A1(net376));
 sg13g2_nor2_2 _08486_ (.A(_02288_),
    .B(net427),
    .Y(_03083_));
 sg13g2_a21oi_1 _08487_ (.A1(net214),
    .A2(_03083_),
    .Y(_03084_),
    .B1(net325));
 sg13g2_o21ai_1 _08488_ (.B1(_03084_),
    .Y(_03085_),
    .A1(net177),
    .A2(_03082_));
 sg13g2_buf_1 _08489_ (.A(net288),
    .X(_03086_));
 sg13g2_o21ai_1 _08490_ (.B1(net287),
    .Y(_03087_),
    .A1(net169),
    .A2(_02350_));
 sg13g2_nand3_1 _08491_ (.B(_03085_),
    .C(_03087_),
    .A(_02823_),
    .Y(_03088_));
 sg13g2_nand2_1 _08492_ (.Y(_03089_),
    .A(net340),
    .B(_03066_));
 sg13g2_nand2_1 _08493_ (.Y(_03090_),
    .A(_02564_),
    .B(net187));
 sg13g2_nand2_1 _08494_ (.Y(_03091_),
    .A(_03089_),
    .B(_03090_));
 sg13g2_nand2_1 _08495_ (.Y(_03092_),
    .A(net337),
    .B(_02564_));
 sg13g2_nand3_1 _08496_ (.B(_03092_),
    .C(_03069_),
    .A(net339),
    .Y(_03093_));
 sg13g2_o21ai_1 _08497_ (.B1(_03093_),
    .Y(_03094_),
    .A1(net192),
    .A2(_03091_));
 sg13g2_o21ai_1 _08498_ (.B1(_02502_),
    .Y(_03095_),
    .A1(_03088_),
    .A2(_03094_));
 sg13g2_a21oi_1 _08499_ (.A1(_03074_),
    .A2(_03081_),
    .Y(_03096_),
    .B1(_03095_));
 sg13g2_a21o_1 _08500_ (.A2(_03073_),
    .A1(_03088_),
    .B1(net123),
    .X(_03097_));
 sg13g2_o21ai_1 _08501_ (.B1(_02847_),
    .Y(_03098_),
    .A1(net312),
    .A2(_02601_));
 sg13g2_a221oi_1 _08502_ (.B2(net234),
    .C1(_01911_),
    .B1(_03098_),
    .A1(net169),
    .Y(_03099_),
    .A2(_02696_));
 sg13g2_a21oi_1 _08503_ (.A1(net462),
    .A2(_03075_),
    .Y(_03100_),
    .B1(_02359_));
 sg13g2_buf_2 _08504_ (.A(_03100_),
    .X(_03101_));
 sg13g2_o21ai_1 _08505_ (.B1(_03101_),
    .Y(_03102_),
    .A1(net248),
    .A2(_02653_));
 sg13g2_nand2_1 _08506_ (.Y(_03103_),
    .A(_02799_),
    .B(_03102_));
 sg13g2_nor2_1 _08507_ (.A(_03099_),
    .B(_03103_),
    .Y(_03104_));
 sg13g2_buf_1 _08508_ (.A(_02537_),
    .X(_03105_));
 sg13g2_nand2_2 _08509_ (.Y(_03106_),
    .A(_02844_),
    .B(_02851_));
 sg13g2_o21ai_1 _08510_ (.B1(_02836_),
    .Y(_03107_),
    .A1(net240),
    .A2(_03106_));
 sg13g2_a21oi_1 _08511_ (.A1(net100),
    .A2(_03077_),
    .Y(_03108_),
    .B1(_03107_));
 sg13g2_a21oi_1 _08512_ (.A1(_03104_),
    .A2(_03108_),
    .Y(_03109_),
    .B1(_02502_));
 sg13g2_nor2_1 _08513_ (.A(_02460_),
    .B(net463),
    .Y(_03110_));
 sg13g2_nor3_1 _08514_ (.A(net311),
    .B(net196),
    .C(_03110_),
    .Y(_03111_));
 sg13g2_a21oi_1 _08515_ (.A1(net211),
    .A2(net183),
    .Y(_03112_),
    .B1(_03111_));
 sg13g2_a21o_1 _08516_ (.A2(_02544_),
    .A1(net211),
    .B1(_02980_),
    .X(_03113_));
 sg13g2_o21ai_1 _08517_ (.B1(_03113_),
    .Y(_03114_),
    .A1(net103),
    .A2(_03112_));
 sg13g2_nand2_2 _08518_ (.Y(_03115_),
    .A(net383),
    .B(net377));
 sg13g2_nand3_1 _08519_ (.B(_02417_),
    .C(_03115_),
    .A(_01917_),
    .Y(_03116_));
 sg13g2_a21oi_1 _08520_ (.A1(_01976_),
    .A2(_03116_),
    .Y(_03117_),
    .B1(_02703_));
 sg13g2_o21ai_1 _08521_ (.B1(_02351_),
    .Y(_03118_),
    .A1(net196),
    .A2(_03110_));
 sg13g2_nand2_2 _08522_ (.Y(_03119_),
    .A(net317),
    .B(net427));
 sg13g2_nor2b_1 _08523_ (.A(net379),
    .B_N(_01884_),
    .Y(_03120_));
 sg13g2_buf_2 _08524_ (.A(_03120_),
    .X(_03121_));
 sg13g2_nand2_1 _08525_ (.Y(_03122_),
    .A(_02388_),
    .B(_03121_));
 sg13g2_nand4_1 _08526_ (.B(net307),
    .C(_03119_),
    .A(net330),
    .Y(_03123_),
    .D(_03122_));
 sg13g2_nand3_1 _08527_ (.B(_03118_),
    .C(_03123_),
    .A(_02554_),
    .Y(_03124_));
 sg13g2_nand2_1 _08528_ (.Y(_03125_),
    .A(_01899_),
    .B(_02847_));
 sg13g2_a21oi_1 _08529_ (.A1(net331),
    .A2(_03014_),
    .Y(_03126_),
    .B1(net327));
 sg13g2_o21ai_1 _08530_ (.B1(_02340_),
    .Y(_03127_),
    .A1(_03125_),
    .A2(_03126_));
 sg13g2_nand3_1 _08531_ (.B(_03119_),
    .C(_02464_),
    .A(net318),
    .Y(_03128_));
 sg13g2_nand3_1 _08532_ (.B(_03127_),
    .C(_03128_),
    .A(_01769_),
    .Y(_03129_));
 sg13g2_nand3_1 _08533_ (.B(_03124_),
    .C(_03129_),
    .A(_03117_),
    .Y(_03130_));
 sg13g2_a21oi_1 _08534_ (.A1(net118),
    .A2(_03114_),
    .Y(_03131_),
    .B1(_03130_));
 sg13g2_nand2b_1 _08535_ (.Y(_03132_),
    .B(_03130_),
    .A_N(_03104_));
 sg13g2_o21ai_1 _08536_ (.B1(_03132_),
    .Y(_03133_),
    .A1(net149),
    .A2(_03131_));
 sg13g2_a221oi_1 _08537_ (.B2(_03133_),
    .C1(_02495_),
    .B1(_03109_),
    .A1(_03096_),
    .Y(_03134_),
    .A2(_03097_));
 sg13g2_nor2_1 _08538_ (.A(net327),
    .B(net423),
    .Y(_03135_));
 sg13g2_a21o_1 _08539_ (.A2(net463),
    .A1(net329),
    .B1(_03135_),
    .X(_03136_));
 sg13g2_nand2_1 _08540_ (.Y(_03137_),
    .A(net332),
    .B(net305));
 sg13g2_o21ai_1 _08541_ (.B1(_03137_),
    .Y(_03138_),
    .A1(net220),
    .A2(net232));
 sg13g2_buf_1 _08542_ (.A(_02345_),
    .X(_03139_));
 sg13g2_a221oi_1 _08543_ (.B2(_03139_),
    .C1(net336),
    .B1(_03138_),
    .A1(_03022_),
    .Y(_03140_),
    .A2(_03136_));
 sg13g2_o21ai_1 _08544_ (.B1(_03140_),
    .Y(_03141_),
    .A1(_02304_),
    .A2(net232));
 sg13g2_buf_1 _08545_ (.A(_02926_),
    .X(_03142_));
 sg13g2_nor2_1 _08546_ (.A(net99),
    .B(_03110_),
    .Y(_03143_));
 sg13g2_nand2_1 _08547_ (.Y(_03144_),
    .A(net243),
    .B(net281));
 sg13g2_nand2_1 _08548_ (.Y(_03145_),
    .A(net323),
    .B(net289));
 sg13g2_o21ai_1 _08549_ (.B1(_03145_),
    .Y(_03146_),
    .A1(net242),
    .A2(_03144_));
 sg13g2_o21ai_1 _08550_ (.B1(_03146_),
    .Y(_03147_),
    .A1(net339),
    .A2(_03143_));
 sg13g2_nor2_1 _08551_ (.A(net152),
    .B(_03147_),
    .Y(_03148_));
 sg13g2_nor2_2 _08552_ (.A(net317),
    .B(_02288_),
    .Y(_03149_));
 sg13g2_buf_1 _08553_ (.A(_02344_),
    .X(_03150_));
 sg13g2_nor2_1 _08554_ (.A(net168),
    .B(net169),
    .Y(_03151_));
 sg13g2_o21ai_1 _08555_ (.B1(net239),
    .Y(_03152_),
    .A1(_03149_),
    .A2(_03151_));
 sg13g2_o21ai_1 _08556_ (.B1(net217),
    .Y(_03153_),
    .A1(net211),
    .A2(net207));
 sg13g2_nand4_1 _08557_ (.B(_02944_),
    .C(_03152_),
    .A(net298),
    .Y(_03154_),
    .D(_03153_));
 sg13g2_o21ai_1 _08558_ (.B1(_03154_),
    .Y(_03155_),
    .A1(_03141_),
    .A2(_03148_));
 sg13g2_nand2_1 _08559_ (.Y(_03156_),
    .A(_02289_),
    .B(net374));
 sg13g2_a221oi_1 _08560_ (.B2(net128),
    .C1(_02645_),
    .B1(net308),
    .A1(net131),
    .Y(_03157_),
    .A2(_03156_));
 sg13g2_nor2b_1 _08561_ (.A(_02382_),
    .B_N(net463),
    .Y(_03158_));
 sg13g2_buf_2 _08562_ (.A(_03158_),
    .X(_03159_));
 sg13g2_nand2_1 _08563_ (.Y(_03160_),
    .A(net318),
    .B(net378));
 sg13g2_buf_1 _08564_ (.A(net120),
    .X(_03161_));
 sg13g2_a21oi_1 _08565_ (.A1(net283),
    .A2(_03160_),
    .Y(_03162_),
    .B1(net77));
 sg13g2_a21oi_1 _08566_ (.A1(net131),
    .A2(_03159_),
    .Y(_03163_),
    .B1(_03162_));
 sg13g2_nand2_1 _08567_ (.Y(_03164_),
    .A(net118),
    .B(_03163_));
 sg13g2_o21ai_1 _08568_ (.B1(_03164_),
    .Y(_03165_),
    .A1(net151),
    .A2(_03157_));
 sg13g2_a22oi_1 _08569_ (.Y(_03166_),
    .B1(_03165_),
    .B2(_02795_),
    .A2(_03155_),
    .A1(net109));
 sg13g2_nor2b_1 _08570_ (.A(_03166_),
    .B_N(_02777_),
    .Y(_03167_));
 sg13g2_o21ai_1 _08571_ (.B1(_02772_),
    .Y(_03168_),
    .A1(_03134_),
    .A2(_03167_));
 sg13g2_o21ai_1 _08572_ (.B1(_03168_),
    .Y(_03169_),
    .A1(_03046_),
    .A2(_03061_));
 sg13g2_mux2_1 _08573_ (.A0(_03136_),
    .A1(net102),
    .S(net116),
    .X(_03170_));
 sg13g2_nor2b_1 _08574_ (.A(net389),
    .B_N(net461),
    .Y(_03171_));
 sg13g2_a21oi_1 _08575_ (.A1(net155),
    .A2(net209),
    .Y(_03172_),
    .B1(_03171_));
 sg13g2_o21ai_1 _08576_ (.B1(net231),
    .Y(_03173_),
    .A1(net144),
    .A2(_03172_));
 sg13g2_nand2_1 _08577_ (.Y(_03174_),
    .A(net191),
    .B(_02653_));
 sg13g2_nand2_2 _08578_ (.Y(_03175_),
    .A(_02756_),
    .B(net376));
 sg13g2_nand3_1 _08579_ (.B(net111),
    .C(_03175_),
    .A(_01888_),
    .Y(_03176_));
 sg13g2_nand2_1 _08580_ (.Y(_03177_),
    .A(_03174_),
    .B(_03176_));
 sg13g2_mux4_1 _08581_ (.S0(net152),
    .A0(_03143_),
    .A1(_03170_),
    .A2(_03173_),
    .A3(_03177_),
    .S1(net139),
    .X(_03178_));
 sg13g2_nor2_1 _08582_ (.A(net185),
    .B(_03178_),
    .Y(_03179_));
 sg13g2_a21oi_1 _08583_ (.A1(_02810_),
    .A2(net111),
    .Y(_03180_),
    .B1(_02741_));
 sg13g2_a221oi_1 _08584_ (.B2(_02741_),
    .C1(_03180_),
    .B1(_02514_),
    .A1(net104),
    .Y(_03181_),
    .A2(_03052_));
 sg13g2_nand3_1 _08585_ (.B(_02750_),
    .C(_03012_),
    .A(_03105_),
    .Y(_03182_));
 sg13g2_o21ai_1 _08586_ (.B1(_03182_),
    .Y(_03183_),
    .A1(net82),
    .A2(_03181_));
 sg13g2_nand2_1 _08587_ (.Y(_03184_),
    .A(_01900_),
    .B(_02875_));
 sg13g2_nand2_1 _08588_ (.Y(_03185_),
    .A(_02548_),
    .B(_03014_));
 sg13g2_o21ai_1 _08589_ (.B1(_02583_),
    .Y(_03186_),
    .A1(net173),
    .A2(_02514_));
 sg13g2_nand3_1 _08590_ (.B(_03185_),
    .C(_03186_),
    .A(net103),
    .Y(_03187_));
 sg13g2_o21ai_1 _08591_ (.B1(_03187_),
    .Y(_03188_),
    .A1(net142),
    .A2(_03184_));
 sg13g2_nand2_1 _08592_ (.Y(_03189_),
    .A(_02469_),
    .B(_02382_));
 sg13g2_buf_1 _08593_ (.A(_03189_),
    .X(_03190_));
 sg13g2_nor2_1 _08594_ (.A(net218),
    .B(net223),
    .Y(_03191_));
 sg13g2_a21oi_1 _08595_ (.A1(net217),
    .A2(_02558_),
    .Y(_03192_),
    .B1(_03191_));
 sg13g2_buf_1 _08596_ (.A(net186),
    .X(_03193_));
 sg13g2_a221oi_1 _08597_ (.B2(net144),
    .C1(net98),
    .B1(_03192_),
    .A1(net216),
    .Y(_03194_),
    .A2(net167));
 sg13g2_a21oi_1 _08598_ (.A1(net151),
    .A2(_03188_),
    .Y(_03195_),
    .B1(_03194_));
 sg13g2_a22oi_1 _08599_ (.Y(_03196_),
    .B1(_03195_),
    .B2(net123),
    .A2(_03183_),
    .A1(net228));
 sg13g2_nor2_1 _08600_ (.A(net122),
    .B(_03196_),
    .Y(_03197_));
 sg13g2_o21ai_1 _08601_ (.B1(_02828_),
    .Y(_03198_),
    .A1(_03179_),
    .A2(_03197_));
 sg13g2_nor4_1 _08602_ (.A(net114),
    .B(_02446_),
    .C(_02710_),
    .D(net225),
    .Y(_03199_));
 sg13g2_nor2_1 _08603_ (.A(net424),
    .B(_03199_),
    .Y(_03200_));
 sg13g2_o21ai_1 _08604_ (.B1(_02422_),
    .Y(_03201_),
    .A1(net294),
    .A2(_02923_));
 sg13g2_and2_1 _08605_ (.A(_03161_),
    .B(_03201_),
    .X(_03202_));
 sg13g2_nand2_1 _08606_ (.Y(_03203_),
    .A(net330),
    .B(net231));
 sg13g2_nand2_1 _08607_ (.Y(_03204_),
    .A(net328),
    .B(_02601_));
 sg13g2_o21ai_1 _08608_ (.B1(_03204_),
    .Y(_03205_),
    .A1(_03202_),
    .A2(_03203_));
 sg13g2_nand2_1 _08609_ (.Y(_03206_),
    .A(_01942_),
    .B(net306));
 sg13g2_nor2_1 _08610_ (.A(net390),
    .B(net293),
    .Y(_03207_));
 sg13g2_o21ai_1 _08611_ (.B1(net127),
    .Y(_03208_),
    .A1(net168),
    .A2(_03207_));
 sg13g2_nand4_1 _08612_ (.B(_02466_),
    .C(_03206_),
    .A(net249),
    .Y(_03209_),
    .D(_03208_));
 sg13g2_o21ai_1 _08613_ (.B1(_03209_),
    .Y(_03210_),
    .A1(net132),
    .A2(_03205_));
 sg13g2_buf_1 _08614_ (.A(_03037_),
    .X(_03211_));
 sg13g2_nor2_1 _08615_ (.A(net166),
    .B(net225),
    .Y(_03212_));
 sg13g2_nor2_1 _08616_ (.A(_01954_),
    .B(net439),
    .Y(_03213_));
 sg13g2_buf_2 _08617_ (.A(_03213_),
    .X(_03214_));
 sg13g2_o21ai_1 _08618_ (.B1(net141),
    .Y(_03215_),
    .A1(_03214_),
    .A2(_03149_));
 sg13g2_a21oi_1 _08619_ (.A1(_03212_),
    .A2(_03215_),
    .Y(_03216_),
    .B1(_01963_));
 sg13g2_nand2_1 _08620_ (.Y(_03217_),
    .A(net184),
    .B(net102));
 sg13g2_inv_1 _08621_ (.Y(_03218_),
    .A(net467));
 sg13g2_nand3_1 _08622_ (.B(_03218_),
    .C(_03005_),
    .A(net340),
    .Y(_03219_));
 sg13g2_nand3_1 _08623_ (.B(_03217_),
    .C(_03219_),
    .A(net282),
    .Y(_03220_));
 sg13g2_a22oi_1 _08624_ (.Y(_03221_),
    .B1(_03216_),
    .B2(_03220_),
    .A2(_03210_),
    .A1(net140));
 sg13g2_nor2_1 _08625_ (.A(_02504_),
    .B(_03221_),
    .Y(_03222_));
 sg13g2_nand3_1 _08626_ (.B(_03200_),
    .C(_03222_),
    .A(net316),
    .Y(_03223_));
 sg13g2_nand2_1 _08627_ (.Y(_03224_),
    .A(_01899_),
    .B(net212));
 sg13g2_buf_2 _08628_ (.A(_03224_),
    .X(_03225_));
 sg13g2_a21oi_1 _08629_ (.A1(_02402_),
    .A2(_03225_),
    .Y(_03226_),
    .B1(_01983_));
 sg13g2_nor2_1 _08630_ (.A(_02947_),
    .B(_03226_),
    .Y(_03227_));
 sg13g2_o21ai_1 _08631_ (.B1(_02578_),
    .Y(_03228_),
    .A1(net191),
    .A2(net253));
 sg13g2_nor2_1 _08632_ (.A(_01967_),
    .B(_02812_),
    .Y(_03229_));
 sg13g2_nor2_1 _08633_ (.A(net392),
    .B(_02711_),
    .Y(_03230_));
 sg13g2_and2_1 _08634_ (.A(net322),
    .B(_03230_),
    .X(_03231_));
 sg13g2_a21oi_1 _08635_ (.A1(_03228_),
    .A2(_03229_),
    .Y(_03232_),
    .B1(_03231_));
 sg13g2_nand2_1 _08636_ (.Y(_03233_),
    .A(net391),
    .B(net385));
 sg13g2_nor2_1 _08637_ (.A(net135),
    .B(_03233_),
    .Y(_03234_));
 sg13g2_inv_1 _08638_ (.Y(_03235_),
    .A(_02812_));
 sg13g2_a221oi_1 _08639_ (.B2(_03235_),
    .C1(net237),
    .B1(_03234_),
    .A1(net106),
    .Y(_03236_),
    .A2(_03225_));
 sg13g2_a21o_1 _08640_ (.A2(_03232_),
    .A1(net149),
    .B1(_03236_),
    .X(_03237_));
 sg13g2_nor2_1 _08641_ (.A(_02812_),
    .B(net420),
    .Y(_03238_));
 sg13g2_nor2_1 _08642_ (.A(_02319_),
    .B(_02429_),
    .Y(_03239_));
 sg13g2_nand3_1 _08643_ (.B(_03225_),
    .C(_03239_),
    .A(_03238_),
    .Y(_03240_));
 sg13g2_nand2_1 _08644_ (.Y(_03241_),
    .A(_01925_),
    .B(_02320_));
 sg13g2_nand2_1 _08645_ (.Y(_03242_),
    .A(net391),
    .B(_02441_));
 sg13g2_nor2_1 _08646_ (.A(_01960_),
    .B(net460),
    .Y(_03243_));
 sg13g2_and3_1 _08647_ (.X(_03244_),
    .A(_03241_),
    .B(_03242_),
    .C(_03243_));
 sg13g2_a21oi_1 _08648_ (.A1(_03225_),
    .A2(_03244_),
    .Y(_03245_),
    .B1(net421));
 sg13g2_a22oi_1 _08649_ (.Y(_03246_),
    .B1(_03240_),
    .B2(_03245_),
    .A2(_03237_),
    .A1(net108));
 sg13g2_and2_1 _08650_ (.A(net173),
    .B(_03241_),
    .X(_03247_));
 sg13g2_buf_1 _08651_ (.A(_03247_),
    .X(_03248_));
 sg13g2_nor2_1 _08652_ (.A(net247),
    .B(_03248_),
    .Y(_03249_));
 sg13g2_buf_1 _08653_ (.A(net99),
    .X(_03250_));
 sg13g2_a21oi_1 _08654_ (.A1(net98),
    .A2(_03250_),
    .Y(_03251_),
    .B1(_02967_));
 sg13g2_nor3_1 _08655_ (.A(net424),
    .B(_03249_),
    .C(_03251_),
    .Y(_03252_));
 sg13g2_nor2_2 _08656_ (.A(net296),
    .B(_02359_),
    .Y(_03253_));
 sg13g2_a21oi_1 _08657_ (.A1(net88),
    .A2(net246),
    .Y(_03254_),
    .B1(_03253_));
 sg13g2_a221oi_1 _08658_ (.B2(net245),
    .C1(net198),
    .B1(net204),
    .A1(net76),
    .Y(_03255_),
    .A2(net199));
 sg13g2_o21ai_1 _08659_ (.B1(_03255_),
    .Y(_03256_),
    .A1(_02684_),
    .A2(_03254_));
 sg13g2_o21ai_1 _08660_ (.B1(_03256_),
    .Y(_03257_),
    .A1(net444),
    .A2(_03252_));
 sg13g2_inv_1 _08661_ (.Y(_03258_),
    .A(_03257_));
 sg13g2_a21oi_1 _08662_ (.A1(net60),
    .A2(net80),
    .Y(_03259_),
    .B1(net386));
 sg13g2_nor2_2 _08663_ (.A(_02664_),
    .B(_03259_),
    .Y(_03260_));
 sg13g2_a22oi_1 _08664_ (.Y(_03261_),
    .B1(_03258_),
    .B2(_03260_),
    .A2(_03246_),
    .A1(_03227_));
 sg13g2_nor2_1 _08665_ (.A(_02339_),
    .B(net463),
    .Y(_03262_));
 sg13g2_a221oi_1 _08666_ (.B2(_02383_),
    .C1(net238),
    .B1(_03262_),
    .A1(net240),
    .Y(_03263_),
    .A2(_02710_));
 sg13g2_o21ai_1 _08667_ (.B1(net155),
    .Y(_03264_),
    .A1(_02766_),
    .A2(_03027_));
 sg13g2_o21ai_1 _08668_ (.B1(net287),
    .Y(_03265_),
    .A1(net288),
    .A2(net306));
 sg13g2_nand2_1 _08669_ (.Y(_03266_),
    .A(_02823_),
    .B(_03265_));
 sg13g2_a21oi_1 _08670_ (.A1(_03263_),
    .A2(_03264_),
    .Y(_03267_),
    .B1(_03266_));
 sg13g2_a21oi_1 _08671_ (.A1(net393),
    .A2(_02863_),
    .Y(_03268_),
    .B1(_02355_));
 sg13g2_nor2_1 _08672_ (.A(net300),
    .B(_03268_),
    .Y(_03269_));
 sg13g2_a21oi_1 _08673_ (.A1(net119),
    .A2(net141),
    .Y(_03270_),
    .B1(_03269_));
 sg13g2_nand3_1 _08674_ (.B(net394),
    .C(net379),
    .A(_01766_),
    .Y(_03271_));
 sg13g2_buf_1 _08675_ (.A(_03271_),
    .X(_03272_));
 sg13g2_o21ai_1 _08676_ (.B1(_03272_),
    .Y(_03273_),
    .A1(net282),
    .A2(_03207_));
 sg13g2_a22oi_1 _08677_ (.Y(_03274_),
    .B1(_03273_),
    .B2(_02472_),
    .A2(_02731_),
    .A1(net176));
 sg13g2_o21ai_1 _08678_ (.B1(_03274_),
    .Y(_03275_),
    .A1(net126),
    .A2(_03270_));
 sg13g2_nand3_1 _08679_ (.B(_02684_),
    .C(_02864_),
    .A(net208),
    .Y(_03276_));
 sg13g2_nor2_1 _08680_ (.A(_02733_),
    .B(_02936_),
    .Y(_03277_));
 sg13g2_nor2_1 _08681_ (.A(net120),
    .B(net299),
    .Y(_03278_));
 sg13g2_o21ai_1 _08682_ (.B1(_02612_),
    .Y(_03279_),
    .A1(_02628_),
    .A2(net321));
 sg13g2_nand2b_1 _08683_ (.Y(_03280_),
    .B(_03279_),
    .A_N(_03278_));
 sg13g2_o21ai_1 _08684_ (.B1(net313),
    .Y(_03281_),
    .A1(_02336_),
    .A2(net306));
 sg13g2_nand2_1 _08685_ (.Y(_03282_),
    .A(_01976_),
    .B(_02847_));
 sg13g2_o21ai_1 _08686_ (.B1(_02799_),
    .Y(_03283_),
    .A1(_03281_),
    .A2(_03282_));
 sg13g2_a221oi_1 _08687_ (.B2(net320),
    .C1(_03283_),
    .B1(_03280_),
    .A1(_03276_),
    .Y(_03284_),
    .A2(_03277_));
 sg13g2_nand2_1 _08688_ (.Y(_03285_),
    .A(net317),
    .B(_02355_));
 sg13g2_nor2b_1 _08689_ (.A(_03281_),
    .B_N(_03285_),
    .Y(_03286_));
 sg13g2_nor2_1 _08690_ (.A(net142),
    .B(_03106_),
    .Y(_03287_));
 sg13g2_nor3_1 _08691_ (.A(_02749_),
    .B(_03286_),
    .C(_03287_),
    .Y(_03288_));
 sg13g2_a22oi_1 _08692_ (.Y(_03289_),
    .B1(_03284_),
    .B2(_03288_),
    .A2(_03275_),
    .A1(_03267_));
 sg13g2_o21ai_1 _08693_ (.B1(net140),
    .Y(_03290_),
    .A1(_03267_),
    .A2(_03284_));
 sg13g2_nand2_1 _08694_ (.Y(_03291_),
    .A(_03289_),
    .B(_03290_));
 sg13g2_nand2_1 _08695_ (.Y(_03292_),
    .A(_02489_),
    .B(_02603_));
 sg13g2_and2_1 _08696_ (.A(_01885_),
    .B(net383),
    .X(_03293_));
 sg13g2_buf_1 _08697_ (.A(_03293_),
    .X(_03294_));
 sg13g2_o21ai_1 _08698_ (.B1(_02373_),
    .Y(_03295_),
    .A1(_03294_),
    .A2(net190));
 sg13g2_a21oi_1 _08699_ (.A1(net60),
    .A2(_03295_),
    .Y(_03296_),
    .B1(net386));
 sg13g2_nor2_1 _08700_ (.A(_03292_),
    .B(_03296_),
    .Y(_03297_));
 sg13g2_buf_1 _08701_ (.A(_03161_),
    .X(_03298_));
 sg13g2_buf_1 _08702_ (.A(net168),
    .X(_03299_));
 sg13g2_nand2_1 _08703_ (.Y(_03300_),
    .A(_02298_),
    .B(net427));
 sg13g2_a21oi_1 _08704_ (.A1(net97),
    .A2(_03300_),
    .Y(_03301_),
    .B1(_02570_));
 sg13g2_nor3_1 _08705_ (.A(_02717_),
    .B(net334),
    .C(net283),
    .Y(_03302_));
 sg13g2_o21ai_1 _08706_ (.B1(_02584_),
    .Y(_03303_),
    .A1(net133),
    .A2(_03302_));
 sg13g2_o21ai_1 _08707_ (.B1(_03303_),
    .Y(_03304_),
    .A1(net58),
    .A2(_03301_));
 sg13g2_buf_1 _08708_ (.A(net319),
    .X(_03305_));
 sg13g2_buf_1 _08709_ (.A(net165),
    .X(_03306_));
 sg13g2_a21oi_1 _08710_ (.A1(net207),
    .A2(net136),
    .Y(_03307_),
    .B1(_03306_));
 sg13g2_o21ai_1 _08711_ (.B1(net245),
    .Y(_03308_),
    .A1(net322),
    .A2(_03307_));
 sg13g2_nor2_1 _08712_ (.A(_02468_),
    .B(_02852_),
    .Y(_03309_));
 sg13g2_o21ai_1 _08713_ (.B1(_02637_),
    .Y(_03310_),
    .A1(net219),
    .A2(_03309_));
 sg13g2_nand2_1 _08714_ (.Y(_03311_),
    .A(_03308_),
    .B(_03310_));
 sg13g2_o21ai_1 _08715_ (.B1(_03311_),
    .Y(_03312_),
    .A1(net252),
    .A2(_03304_));
 sg13g2_nor2_1 _08716_ (.A(net331),
    .B(_02684_),
    .Y(_03313_));
 sg13g2_buf_1 _08717_ (.A(_03313_),
    .X(_03314_));
 sg13g2_nor2_1 _08718_ (.A(net219),
    .B(net95),
    .Y(_03315_));
 sg13g2_nor2_1 _08719_ (.A(net318),
    .B(_03012_),
    .Y(_03316_));
 sg13g2_nor3_1 _08720_ (.A(net313),
    .B(net189),
    .C(_03029_),
    .Y(_03317_));
 sg13g2_nor3_1 _08721_ (.A(net177),
    .B(_03316_),
    .C(_03317_),
    .Y(_03318_));
 sg13g2_nand2_1 _08722_ (.Y(_03319_),
    .A(net333),
    .B(_02383_));
 sg13g2_a22oi_1 _08723_ (.Y(_03320_),
    .B1(net167),
    .B2(net168),
    .A2(_03319_),
    .A1(net328));
 sg13g2_o21ai_1 _08724_ (.B1(net314),
    .Y(_03321_),
    .A1(net105),
    .A2(_03320_));
 sg13g2_o21ai_1 _08725_ (.B1(_03239_),
    .Y(_03322_),
    .A1(_03318_),
    .A2(_03321_));
 sg13g2_a21oi_1 _08726_ (.A1(_03026_),
    .A2(_03315_),
    .Y(_03323_),
    .B1(_03322_));
 sg13g2_nand2_1 _08727_ (.Y(_03324_),
    .A(net307),
    .B(_03022_));
 sg13g2_o21ai_1 _08728_ (.B1(_03243_),
    .Y(_03325_),
    .A1(_03015_),
    .A2(_03324_));
 sg13g2_buf_1 _08729_ (.A(net309),
    .X(_03326_));
 sg13g2_a221oi_1 _08730_ (.B2(net164),
    .C1(_03211_),
    .B1(_03319_),
    .A1(net145),
    .Y(_03327_),
    .A2(net239));
 sg13g2_nor2_1 _08731_ (.A(net433),
    .B(_02614_),
    .Y(_03328_));
 sg13g2_nor3_1 _08732_ (.A(net219),
    .B(_02608_),
    .C(_03328_),
    .Y(_03329_));
 sg13g2_nor3_1 _08733_ (.A(_03325_),
    .B(_03327_),
    .C(_03329_),
    .Y(_03330_));
 sg13g2_nor2_1 _08734_ (.A(_03323_),
    .B(_03330_),
    .Y(_03331_));
 sg13g2_a22oi_1 _08735_ (.Y(_03332_),
    .B1(_03331_),
    .B2(_02507_),
    .A2(_03312_),
    .A1(net109));
 sg13g2_inv_1 _08736_ (.Y(_03333_),
    .A(_02919_));
 sg13g2_a221oi_1 _08737_ (.B2(_03332_),
    .C1(_03333_),
    .B1(_03297_),
    .A1(_02883_),
    .Y(_03334_),
    .A2(_03291_));
 sg13g2_nand4_1 _08738_ (.B(_03223_),
    .C(_03261_),
    .A(_03198_),
    .Y(_03335_),
    .D(_03334_));
 sg13g2_a21oi_1 _08739_ (.A1(net99),
    .A2(_03242_),
    .Y(_03336_),
    .B1(net187));
 sg13g2_a21oi_1 _08740_ (.A1(net154),
    .A2(_02968_),
    .Y(_03337_),
    .B1(_03336_));
 sg13g2_nor2_1 _08741_ (.A(net87),
    .B(net210),
    .Y(_03338_));
 sg13g2_a221oi_1 _08742_ (.B2(net80),
    .C1(net122),
    .B1(_03338_),
    .A1(net87),
    .Y(_03339_),
    .A2(_03337_));
 sg13g2_or2_1 _08743_ (.X(_03340_),
    .B(_03245_),
    .A(_03226_));
 sg13g2_o21ai_1 _08744_ (.B1(_03333_),
    .Y(_03341_),
    .A1(_03339_),
    .A2(_03340_));
 sg13g2_o21ai_1 _08745_ (.B1(_03341_),
    .Y(_03342_),
    .A1(_03169_),
    .A2(_03335_));
 sg13g2_a22oi_1 _08746_ (.Y(_03343_),
    .B1(_03201_),
    .B2(net240),
    .A2(net378),
    .A1(net211));
 sg13g2_nor2_1 _08747_ (.A(net164),
    .B(_03343_),
    .Y(_03344_));
 sg13g2_nor3_1 _08748_ (.A(net249),
    .B(_02860_),
    .C(_03344_),
    .Y(_03345_));
 sg13g2_nand2_1 _08749_ (.Y(_03346_),
    .A(net169),
    .B(net125));
 sg13g2_nand2_1 _08750_ (.Y(_03347_),
    .A(_02839_),
    .B(net201));
 sg13g2_nand3_1 _08751_ (.B(_03346_),
    .C(_03347_),
    .A(net249),
    .Y(_03348_));
 sg13g2_nor2b_1 _08752_ (.A(_03345_),
    .B_N(_03348_),
    .Y(_03349_));
 sg13g2_buf_1 _08753_ (.A(net283),
    .X(_03350_));
 sg13g2_o21ai_1 _08754_ (.B1(net135),
    .Y(_03351_),
    .A1(_02562_),
    .A2(net163));
 sg13g2_a221oi_1 _08755_ (.B2(net78),
    .C1(net236),
    .B1(_03351_),
    .A1(_01942_),
    .Y(_03352_),
    .A2(net107));
 sg13g2_nor2_1 _08756_ (.A(net291),
    .B(_02644_),
    .Y(_03353_));
 sg13g2_o21ai_1 _08757_ (.B1(net149),
    .Y(_03354_),
    .A1(_03352_),
    .A2(_03353_));
 sg13g2_o21ai_1 _08758_ (.B1(_03354_),
    .Y(_03355_),
    .A1(net140),
    .A2(_03349_));
 sg13g2_nand2_1 _08759_ (.Y(_03356_),
    .A(_01913_),
    .B(_03355_));
 sg13g2_o21ai_1 _08760_ (.B1(net135),
    .Y(_03357_),
    .A1(net210),
    .A2(net174));
 sg13g2_nand2_1 _08761_ (.Y(_03358_),
    .A(net210),
    .B(net204));
 sg13g2_nor2_1 _08762_ (.A(_03358_),
    .B(net281),
    .Y(_03359_));
 sg13g2_a21oi_1 _08763_ (.A1(net58),
    .A2(_03357_),
    .Y(_03360_),
    .B1(_03359_));
 sg13g2_nor2_2 _08764_ (.A(_01929_),
    .B(_01899_),
    .Y(_03361_));
 sg13g2_a21oi_1 _08765_ (.A1(_02647_),
    .A2(net173),
    .Y(_03362_),
    .B1(_01952_));
 sg13g2_nand2b_1 _08766_ (.Y(_03363_),
    .B(_03362_),
    .A_N(_03361_));
 sg13g2_nor2_1 _08767_ (.A(net140),
    .B(_03363_),
    .Y(_03364_));
 sg13g2_a21oi_1 _08768_ (.A1(net87),
    .A2(_03360_),
    .Y(_03365_),
    .B1(_03364_));
 sg13g2_nor2_1 _08769_ (.A(net134),
    .B(_02687_),
    .Y(_03366_));
 sg13g2_a22oi_1 _08770_ (.Y(_03367_),
    .B1(_03365_),
    .B2(_03366_),
    .A2(_03356_),
    .A1(net400));
 sg13g2_nor2_1 _08771_ (.A(_02949_),
    .B(_03367_),
    .Y(_03368_));
 sg13g2_o21ai_1 _08772_ (.B1(net192),
    .Y(_03369_),
    .A1(net114),
    .A2(_02614_));
 sg13g2_o21ai_1 _08773_ (.B1(_02836_),
    .Y(_03370_),
    .A1(net169),
    .A2(net221));
 sg13g2_nor3_1 _08774_ (.A(net285),
    .B(_02601_),
    .C(_03370_),
    .Y(_03371_));
 sg13g2_a21o_1 _08775_ (.A2(_03369_),
    .A1(net202),
    .B1(_03371_),
    .X(_03372_));
 sg13g2_a21oi_1 _08776_ (.A1(_02610_),
    .A2(_03372_),
    .Y(_03373_),
    .B1(net421));
 sg13g2_nor2_1 _08777_ (.A(_02619_),
    .B(net101),
    .Y(_03374_));
 sg13g2_nor3_1 _08778_ (.A(_00091_),
    .B(_02812_),
    .C(net420),
    .Y(_03375_));
 sg13g2_a21oi_1 _08779_ (.A1(_03374_),
    .A2(_03375_),
    .Y(_03376_),
    .B1(_02704_));
 sg13g2_nor3_1 _08780_ (.A(_02605_),
    .B(_03373_),
    .C(_03376_),
    .Y(_03377_));
 sg13g2_a22oi_1 _08781_ (.Y(_03378_),
    .B1(_03358_),
    .B2(net154),
    .A2(net210),
    .A1(net433));
 sg13g2_a21oi_1 _08782_ (.A1(net372),
    .A2(_02697_),
    .Y(_03379_),
    .B1(_02703_));
 sg13g2_o21ai_1 _08783_ (.B1(_03379_),
    .Y(_03380_),
    .A1(net117),
    .A2(_03378_));
 sg13g2_nor2_2 _08784_ (.A(_01960_),
    .B(net459),
    .Y(_03381_));
 sg13g2_nand2_1 _08785_ (.Y(_03382_),
    .A(_02647_),
    .B(_03381_));
 sg13g2_o21ai_1 _08786_ (.B1(_03382_),
    .Y(_03383_),
    .A1(net238),
    .A2(net187));
 sg13g2_nand3_1 _08787_ (.B(net290),
    .C(_03383_),
    .A(net80),
    .Y(_03384_));
 sg13g2_a21oi_1 _08788_ (.A1(_03380_),
    .A2(_03384_),
    .Y(_03385_),
    .B1(_02664_));
 sg13g2_nand2_1 _08789_ (.Y(_03386_),
    .A(_02503_),
    .B(_02772_));
 sg13g2_nand2_1 _08790_ (.Y(_03387_),
    .A(net328),
    .B(_02720_));
 sg13g2_o21ai_1 _08791_ (.B1(_03387_),
    .Y(_03388_),
    .A1(net302),
    .A2(_02570_));
 sg13g2_and2_1 _08792_ (.A(net293),
    .B(net461),
    .X(_03389_));
 sg13g2_a221oi_1 _08793_ (.B2(net289),
    .C1(_03142_),
    .B1(_03389_),
    .A1(net170),
    .Y(_03390_),
    .A2(_02383_));
 sg13g2_a221oi_1 _08794_ (.B2(_03390_),
    .C1(_03231_),
    .B1(net171),
    .A1(net209),
    .Y(_03391_),
    .A2(_03388_));
 sg13g2_buf_1 _08795_ (.A(_02636_),
    .X(_03392_));
 sg13g2_nand2_1 _08796_ (.Y(_03393_),
    .A(net288),
    .B(_02377_));
 sg13g2_nand2_1 _08797_ (.Y(_03394_),
    .A(net112),
    .B(net227));
 sg13g2_nand4_1 _08798_ (.B(net106),
    .C(_03393_),
    .A(net280),
    .Y(_03395_),
    .D(_03394_));
 sg13g2_o21ai_1 _08799_ (.B1(_03395_),
    .Y(_03396_),
    .A1(_02638_),
    .A2(_03391_));
 sg13g2_buf_1 _08800_ (.A(net288),
    .X(_03397_));
 sg13g2_o21ai_1 _08801_ (.B1(net345),
    .Y(_03398_),
    .A1(_02708_),
    .A2(net162));
 sg13g2_nor2_1 _08802_ (.A(net112),
    .B(net111),
    .Y(_03399_));
 sg13g2_a21oi_1 _08803_ (.A1(net58),
    .A2(_03398_),
    .Y(_03400_),
    .B1(_03399_));
 sg13g2_nand2_1 _08804_ (.Y(_03401_),
    .A(net313),
    .B(_02684_));
 sg13g2_o21ai_1 _08805_ (.B1(_03401_),
    .Y(_03402_),
    .A1(net162),
    .A2(net163));
 sg13g2_a221oi_1 _08806_ (.B2(net78),
    .C1(net98),
    .B1(_03402_),
    .A1(net167),
    .Y(_03403_),
    .A2(_03262_));
 sg13g2_a21oi_1 _08807_ (.A1(net132),
    .A2(_03400_),
    .Y(_03404_),
    .B1(_03403_));
 sg13g2_a22oi_1 _08808_ (.Y(_03405_),
    .B1(_02795_),
    .B2(_03404_),
    .A2(_03396_),
    .A1(net109));
 sg13g2_nor2_1 _08809_ (.A(_03386_),
    .B(_03405_),
    .Y(_03406_));
 sg13g2_nor2_1 _08810_ (.A(net373),
    .B(net321),
    .Y(_03407_));
 sg13g2_a22oi_1 _08811_ (.Y(_03408_),
    .B1(_03407_),
    .B2(net101),
    .A2(net321),
    .A1(net107));
 sg13g2_a21oi_1 _08812_ (.A1(net228),
    .A2(_03408_),
    .Y(_03409_),
    .B1(net229));
 sg13g2_o21ai_1 _08813_ (.B1(net283),
    .Y(_03410_),
    .A1(net230),
    .A2(_02378_));
 sg13g2_nand3_1 _08814_ (.B(net197),
    .C(_03062_),
    .A(net77),
    .Y(_03411_));
 sg13g2_o21ai_1 _08815_ (.B1(_03411_),
    .Y(_03412_),
    .A1(net78),
    .A2(_03410_));
 sg13g2_nand3_1 _08816_ (.B(_02388_),
    .C(_02832_),
    .A(net423),
    .Y(_03413_));
 sg13g2_a21oi_1 _08817_ (.A1(net328),
    .A2(_03413_),
    .Y(_03414_),
    .B1(_02748_));
 sg13g2_o21ai_1 _08818_ (.B1(_03414_),
    .Y(_03415_),
    .A1(net131),
    .A2(_02728_));
 sg13g2_a22oi_1 _08819_ (.Y(_03416_),
    .B1(_03415_),
    .B2(_02901_),
    .A2(_03412_),
    .A1(net188));
 sg13g2_a21oi_1 _08820_ (.A1(_02707_),
    .A2(net227),
    .Y(_03417_),
    .B1(net335));
 sg13g2_a21oi_1 _08821_ (.A1(net283),
    .A2(_02732_),
    .Y(_03418_),
    .B1(net208));
 sg13g2_nor3_1 _08822_ (.A(net325),
    .B(_03417_),
    .C(_03418_),
    .Y(_03419_));
 sg13g2_nor2_1 _08823_ (.A(net319),
    .B(net304),
    .Y(_03420_));
 sg13g2_o21ai_1 _08824_ (.B1(_01916_),
    .Y(_03421_),
    .A1(net196),
    .A2(_03420_));
 sg13g2_a21oi_1 _08825_ (.A1(_01976_),
    .A2(_03421_),
    .Y(_03422_),
    .B1(_02703_));
 sg13g2_nor2b_1 _08826_ (.A(_03419_),
    .B_N(_03422_),
    .Y(_03423_));
 sg13g2_o21ai_1 _08827_ (.B1(net133),
    .Y(_03424_),
    .A1(net96),
    .A2(net210));
 sg13g2_nand2_1 _08828_ (.Y(_03425_),
    .A(net323),
    .B(net168));
 sg13g2_nor2b_1 _08829_ (.A(_03425_),
    .B_N(_02511_),
    .Y(_03426_));
 sg13g2_o21ai_1 _08830_ (.B1(net144),
    .Y(_03427_),
    .A1(net170),
    .A2(_03426_));
 sg13g2_nand3_1 _08831_ (.B(_03424_),
    .C(_03427_),
    .A(net123),
    .Y(_03428_));
 sg13g2_a22oi_1 _08832_ (.Y(_03429_),
    .B1(_03423_),
    .B2(_03428_),
    .A2(_03416_),
    .A1(_03409_));
 sg13g2_o21ai_1 _08833_ (.B1(net59),
    .Y(_03430_),
    .A1(_02887_),
    .A2(_03429_));
 sg13g2_nor4_1 _08834_ (.A(_03377_),
    .B(_03385_),
    .C(_03406_),
    .D(_03430_),
    .Y(_03431_));
 sg13g2_a21oi_1 _08835_ (.A1(net131),
    .A2(net180),
    .Y(_03432_),
    .B1(_02805_));
 sg13g2_nand2_1 _08836_ (.Y(_03433_),
    .A(_03218_),
    .B(net133));
 sg13g2_nand2_2 _08837_ (.Y(_03434_),
    .A(_02450_),
    .B(_02373_));
 sg13g2_o21ai_1 _08838_ (.B1(net240),
    .Y(_03435_),
    .A1(net211),
    .A2(_03434_));
 sg13g2_nor2_1 _08839_ (.A(_02461_),
    .B(_02414_),
    .Y(_03436_));
 sg13g2_a221oi_1 _08840_ (.B2(net150),
    .C1(net205),
    .B1(_03436_),
    .A1(_03433_),
    .Y(_03437_),
    .A2(_03435_));
 sg13g2_a21oi_1 _08841_ (.A1(net118),
    .A2(_03432_),
    .Y(_03438_),
    .B1(_03437_));
 sg13g2_o21ai_1 _08842_ (.B1(_02454_),
    .Y(_03439_),
    .A1(net203),
    .A2(net97));
 sg13g2_a21oi_1 _08843_ (.A1(_03425_),
    .A2(_03439_),
    .Y(_03440_),
    .B1(net180));
 sg13g2_nand2_1 _08844_ (.Y(_03441_),
    .A(net172),
    .B(_03440_));
 sg13g2_o21ai_1 _08845_ (.B1(_03441_),
    .Y(_03442_),
    .A1(net117),
    .A2(_03438_));
 sg13g2_a221oi_1 _08846_ (.B2(net311),
    .C1(net315),
    .B1(_02564_),
    .A1(net193),
    .Y(_03443_),
    .A2(net221));
 sg13g2_or3_1 _08847_ (.A(net300),
    .B(_02560_),
    .C(_03443_),
    .X(_03444_));
 sg13g2_nand2_1 _08848_ (.Y(_03445_),
    .A(_02844_),
    .B(net214));
 sg13g2_nand3_1 _08849_ (.B(_03445_),
    .C(_02456_),
    .A(net186),
    .Y(_03446_));
 sg13g2_nand2_1 _08850_ (.Y(_03447_),
    .A(_03444_),
    .B(_03446_));
 sg13g2_o21ai_1 _08851_ (.B1(_03393_),
    .Y(_03448_),
    .A1(net239),
    .A2(net162));
 sg13g2_o21ai_1 _08852_ (.B1(_02574_),
    .Y(_03449_),
    .A1(net224),
    .A2(_02466_));
 sg13g2_a22oi_1 _08853_ (.Y(_03450_),
    .B1(_03449_),
    .B2(net292),
    .A2(_03448_),
    .A1(net298));
 sg13g2_o21ai_1 _08854_ (.B1(_03450_),
    .Y(_03451_),
    .A1(net206),
    .A2(_03447_));
 sg13g2_nand3_1 _08855_ (.B(net60),
    .C(_02589_),
    .A(net401),
    .Y(_03452_));
 sg13g2_o21ai_1 _08856_ (.B1(_03452_),
    .Y(_03453_),
    .A1(net401),
    .A2(_03451_));
 sg13g2_a22oi_1 _08857_ (.Y(_03454_),
    .B1(_03453_),
    .B2(net444),
    .A2(_03442_),
    .A1(net290));
 sg13g2_and2_1 _08858_ (.A(_02489_),
    .B(_02595_),
    .X(_03455_));
 sg13g2_buf_1 _08859_ (.A(_03455_),
    .X(_03456_));
 sg13g2_nand2b_1 _08860_ (.Y(_03457_),
    .B(_03456_),
    .A_N(_03454_));
 sg13g2_inv_1 _08861_ (.Y(_03458_),
    .A(_02536_));
 sg13g2_a21oi_1 _08862_ (.A1(net128),
    .A2(net419),
    .Y(_03459_),
    .B1(_03105_));
 sg13g2_a221oi_1 _08863_ (.B2(_03459_),
    .C1(net151),
    .B1(_03458_),
    .A1(net82),
    .Y(_03460_),
    .A2(_02645_));
 sg13g2_o21ai_1 _08864_ (.B1(net98),
    .Y(_03461_),
    .A1(net162),
    .A2(_02674_));
 sg13g2_o21ai_1 _08865_ (.B1(_02795_),
    .Y(_03462_),
    .A1(_03399_),
    .A2(_03461_));
 sg13g2_nand2_1 _08866_ (.Y(_03463_),
    .A(_02470_),
    .B(net284));
 sg13g2_nand2_1 _08867_ (.Y(_03464_),
    .A(_01885_),
    .B(net427));
 sg13g2_a21oi_1 _08868_ (.A1(_03463_),
    .A2(_03464_),
    .Y(_03465_),
    .B1(net168));
 sg13g2_nor2_1 _08869_ (.A(net310),
    .B(_03465_),
    .Y(_03466_));
 sg13g2_nand2_1 _08870_ (.Y(_03467_),
    .A(net241),
    .B(_02642_));
 sg13g2_o21ai_1 _08871_ (.B1(_03467_),
    .Y(_03468_),
    .A1(net103),
    .A2(_03466_));
 sg13g2_o21ai_1 _08872_ (.B1(net178),
    .Y(_03469_),
    .A1(net200),
    .A2(net183));
 sg13g2_a221oi_1 _08873_ (.B2(net97),
    .C1(net219),
    .B1(_03469_),
    .A1(net103),
    .Y(_03470_),
    .A2(_03034_));
 sg13g2_a21oi_1 _08874_ (.A1(net118),
    .A2(_03468_),
    .Y(_03471_),
    .B1(_03470_));
 sg13g2_o21ai_1 _08875_ (.B1(_02784_),
    .Y(_03472_),
    .A1(net149),
    .A2(_03471_));
 sg13g2_o21ai_1 _08876_ (.B1(_03472_),
    .Y(_03473_),
    .A1(_03460_),
    .A2(_03462_));
 sg13g2_nand4_1 _08877_ (.B(net467),
    .C(_02812_),
    .A(_02283_),
    .Y(_03474_),
    .D(_02576_));
 sg13g2_nand2_1 _08878_ (.Y(_03475_),
    .A(_01886_),
    .B(net233));
 sg13g2_nand2_1 _08879_ (.Y(_03476_),
    .A(net315),
    .B(net101));
 sg13g2_o21ai_1 _08880_ (.B1(_03476_),
    .Y(_03477_),
    .A1(net241),
    .A2(_03475_));
 sg13g2_a221oi_1 _08881_ (.B2(net374),
    .C1(net192),
    .B1(_03477_),
    .A1(_01786_),
    .Y(_03478_),
    .A2(net112));
 sg13g2_a21oi_1 _08882_ (.A1(net98),
    .A2(_03474_),
    .Y(_03479_),
    .B1(_03478_));
 sg13g2_nand3_1 _08883_ (.B(_02389_),
    .C(_03106_),
    .A(_01917_),
    .Y(_03480_));
 sg13g2_nand2_1 _08884_ (.Y(_03481_),
    .A(net216),
    .B(_03119_));
 sg13g2_a22oi_1 _08885_ (.Y(_03482_),
    .B1(_03481_),
    .B2(net199),
    .A2(_03480_),
    .A1(net192));
 sg13g2_nand2b_1 _08886_ (.Y(_03483_),
    .B(net206),
    .A_N(_03482_));
 sg13g2_o21ai_1 _08887_ (.B1(_03483_),
    .Y(_03484_),
    .A1(net172),
    .A2(_03479_));
 sg13g2_o21ai_1 _08888_ (.B1(net109),
    .Y(_03485_),
    .A1(_01771_),
    .A2(_02879_));
 sg13g2_o21ai_1 _08889_ (.B1(net211),
    .Y(_03486_),
    .A1(net176),
    .A2(_03159_));
 sg13g2_nand3_1 _08890_ (.B(_03463_),
    .C(_03486_),
    .A(net163),
    .Y(_03487_));
 sg13g2_o21ai_1 _08891_ (.B1(_02390_),
    .Y(_03488_),
    .A1(_03294_),
    .A2(_03012_));
 sg13g2_nor2_1 _08892_ (.A(net143),
    .B(_03015_),
    .Y(_03489_));
 sg13g2_a221oi_1 _08893_ (.B2(_03489_),
    .C1(net420),
    .B1(_03488_),
    .A1(net100),
    .Y(_03490_),
    .A2(_03487_));
 sg13g2_nor2_1 _08894_ (.A(net311),
    .B(_01786_),
    .Y(_03491_));
 sg13g2_a21oi_1 _08895_ (.A1(_01887_),
    .A2(_02642_),
    .Y(_03492_),
    .B1(_03491_));
 sg13g2_a21oi_1 _08896_ (.A1(_02583_),
    .A2(net197),
    .Y(_03493_),
    .B1(_02352_));
 sg13g2_a22oi_1 _08897_ (.Y(_03494_),
    .B1(_03174_),
    .B2(_03493_),
    .A2(_03492_),
    .A1(_02994_));
 sg13g2_nand3_1 _08898_ (.B(_03458_),
    .C(_02545_),
    .A(net119),
    .Y(_03495_));
 sg13g2_nand4_1 _08899_ (.B(net127),
    .C(_03150_),
    .A(net200),
    .Y(_03496_),
    .D(net167));
 sg13g2_and2_1 _08900_ (.A(net320),
    .B(_03496_),
    .X(_03497_));
 sg13g2_a221oi_1 _08901_ (.B2(_03497_),
    .C1(_02433_),
    .B1(_03495_),
    .A1(net188),
    .Y(_03498_),
    .A2(_03494_));
 sg13g2_o21ai_1 _08902_ (.B1(_03498_),
    .Y(_03499_),
    .A1(net117),
    .A2(_03490_));
 sg13g2_o21ai_1 _08903_ (.B1(_03499_),
    .Y(_03500_),
    .A1(_03484_),
    .A2(_03485_));
 sg13g2_nand2_1 _08904_ (.Y(_03501_),
    .A(_02284_),
    .B(net345));
 sg13g2_o21ai_1 _08905_ (.B1(net227),
    .Y(_03502_),
    .A1(net297),
    .A2(_03501_));
 sg13g2_nor2_1 _08906_ (.A(net372),
    .B(net180),
    .Y(_03503_));
 sg13g2_a22oi_1 _08907_ (.Y(_03504_),
    .B1(_03503_),
    .B2(_02732_),
    .A2(_03502_),
    .A1(net89));
 sg13g2_nor2_1 _08908_ (.A(_02679_),
    .B(net234),
    .Y(_03505_));
 sg13g2_mux2_1 _08909_ (.A0(_02728_),
    .A1(_03184_),
    .S(_02745_),
    .X(_03506_));
 sg13g2_a221oi_1 _08910_ (.B2(_03506_),
    .C1(net205),
    .B1(_03505_),
    .A1(_02718_),
    .Y(_03507_),
    .A2(_02549_));
 sg13g2_a21oi_1 _08911_ (.A1(net132),
    .A2(_03504_),
    .Y(_03508_),
    .B1(_03507_));
 sg13g2_a21oi_1 _08912_ (.A1(net342),
    .A2(net425),
    .Y(_03509_),
    .B1(_03214_));
 sg13g2_nand2_1 _08913_ (.Y(_03510_),
    .A(net313),
    .B(_03171_));
 sg13g2_o21ai_1 _08914_ (.B1(_03510_),
    .Y(_03511_),
    .A1(_02803_),
    .A2(_03509_));
 sg13g2_nand2_1 _08915_ (.Y(_03512_),
    .A(net96),
    .B(_03511_));
 sg13g2_nand2b_1 _08916_ (.Y(_03513_),
    .B(net381),
    .A_N(net432));
 sg13g2_a21oi_1 _08917_ (.A1(net233),
    .A2(_03513_),
    .Y(_03514_),
    .B1(net326));
 sg13g2_nor2_1 _08918_ (.A(net342),
    .B(net233),
    .Y(_03515_));
 sg13g2_o21ai_1 _08919_ (.B1(net242),
    .Y(_03516_),
    .A1(_03514_),
    .A2(_03515_));
 sg13g2_a21oi_1 _08920_ (.A1(_03512_),
    .A2(_03516_),
    .Y(_03517_),
    .B1(_01912_));
 sg13g2_nand2_1 _08921_ (.Y(_03518_),
    .A(net244),
    .B(net169));
 sg13g2_a21oi_1 _08922_ (.A1(net425),
    .A2(net182),
    .Y(_03519_),
    .B1(net242));
 sg13g2_a221oi_1 _08923_ (.B2(_03519_),
    .C1(net238),
    .B1(_03518_),
    .A1(net110),
    .Y(_03520_),
    .A2(_03063_));
 sg13g2_o21ai_1 _08924_ (.B1(_02799_),
    .Y(_03521_),
    .A1(_01978_),
    .A2(_03184_));
 sg13g2_o21ai_1 _08925_ (.B1(net233),
    .Y(_03522_),
    .A1(net312),
    .A2(net307));
 sg13g2_nor2_1 _08926_ (.A(net241),
    .B(_02447_),
    .Y(_03523_));
 sg13g2_o21ai_1 _08927_ (.B1(_03523_),
    .Y(_03524_),
    .A1(_03306_),
    .A2(_03522_));
 sg13g2_a21oi_1 _08928_ (.A1(net217),
    .A2(net425),
    .Y(_03525_),
    .B1(net459));
 sg13g2_a21oi_1 _08929_ (.A1(_03524_),
    .A2(_03525_),
    .Y(_03526_),
    .B1(net280));
 sg13g2_nor4_1 _08930_ (.A(_03517_),
    .B(_03520_),
    .C(_03521_),
    .D(_03526_),
    .Y(_03527_));
 sg13g2_a21oi_1 _08931_ (.A1(_02916_),
    .A2(_03508_),
    .Y(_03528_),
    .B1(_03527_));
 sg13g2_a221oi_1 _08932_ (.B2(net329),
    .C1(net313),
    .B1(net213),
    .A1(net342),
    .Y(_03529_),
    .A2(net376));
 sg13g2_or2_1 _08933_ (.X(_03530_),
    .B(_02345_),
    .A(net394));
 sg13g2_nand3_1 _08934_ (.B(_02404_),
    .C(_03530_),
    .A(net390),
    .Y(_03531_));
 sg13g2_nand2_1 _08935_ (.Y(_03532_),
    .A(net165),
    .B(_03531_));
 sg13g2_nand3_1 _08936_ (.B(net337),
    .C(net221),
    .A(net220),
    .Y(_03533_));
 sg13g2_o21ai_1 _08937_ (.B1(_03533_),
    .Y(_03534_),
    .A1(_03529_),
    .A2(_03532_));
 sg13g2_nor2_1 _08938_ (.A(_02564_),
    .B(_02991_),
    .Y(_03535_));
 sg13g2_a21oi_1 _08939_ (.A1(net321),
    .A2(_03535_),
    .Y(_03536_),
    .B1(net300));
 sg13g2_a221oi_1 _08940_ (.B2(_02419_),
    .C1(net301),
    .B1(_03536_),
    .A1(net192),
    .Y(_03537_),
    .A2(_03534_));
 sg13g2_nor3_1 _08941_ (.A(net330),
    .B(net312),
    .C(net419),
    .Y(_03538_));
 sg13g2_a21oi_1 _08942_ (.A1(net254),
    .A2(net110),
    .Y(_03539_),
    .B1(_03538_));
 sg13g2_o21ai_1 _08943_ (.B1(net287),
    .Y(_03540_),
    .A1(net207),
    .A2(_03539_));
 sg13g2_a21oi_1 _08944_ (.A1(net419),
    .A2(_03513_),
    .Y(_03541_),
    .B1(net318));
 sg13g2_a21oi_1 _08945_ (.A1(net194),
    .A2(net308),
    .Y(_03542_),
    .B1(_03541_));
 sg13g2_nor2_1 _08946_ (.A(net104),
    .B(_03542_),
    .Y(_03543_));
 sg13g2_nor2_1 _08947_ (.A(_03540_),
    .B(_03543_),
    .Y(_03544_));
 sg13g2_o21ai_1 _08948_ (.B1(net320),
    .Y(_03545_),
    .A1(net180),
    .A2(_02892_));
 sg13g2_nand2_1 _08949_ (.Y(_03546_),
    .A(net290),
    .B(_03545_));
 sg13g2_nor3_1 _08950_ (.A(_03537_),
    .B(_03544_),
    .C(_03546_),
    .Y(_03547_));
 sg13g2_nor2_2 _08951_ (.A(net293),
    .B(net338),
    .Y(_03548_));
 sg13g2_nor2_1 _08952_ (.A(net431),
    .B(_03272_),
    .Y(_03549_));
 sg13g2_o21ai_1 _08953_ (.B1(net105),
    .Y(_03550_),
    .A1(_03548_),
    .A2(_03549_));
 sg13g2_nand2_1 _08954_ (.Y(_03551_),
    .A(net431),
    .B(net230));
 sg13g2_nand3_1 _08955_ (.B(_02707_),
    .C(_02375_),
    .A(net382),
    .Y(_03552_));
 sg13g2_nand3_1 _08956_ (.B(_03551_),
    .C(_03552_),
    .A(net130),
    .Y(_03553_));
 sg13g2_nand3_1 _08957_ (.B(_03550_),
    .C(_03553_),
    .A(net186),
    .Y(_03554_));
 sg13g2_nand2_1 _08958_ (.Y(_03555_),
    .A(net390),
    .B(_02844_));
 sg13g2_nand2_1 _08959_ (.Y(_03556_),
    .A(net393),
    .B(_03159_));
 sg13g2_nand3_1 _08960_ (.B(_03555_),
    .C(_03556_),
    .A(net212),
    .Y(_03557_));
 sg13g2_nand2_1 _08961_ (.Y(_03558_),
    .A(_03445_),
    .B(_02574_));
 sg13g2_a221oi_1 _08962_ (.B2(_02554_),
    .C1(net446),
    .B1(_03558_),
    .A1(net399),
    .Y(_03559_),
    .A2(_03557_));
 sg13g2_a22oi_1 _08963_ (.Y(_03560_),
    .B1(_02593_),
    .B2(net79),
    .A2(_03559_),
    .A1(_03554_));
 sg13g2_nor2_1 _08964_ (.A(_02428_),
    .B(_03560_),
    .Y(_03561_));
 sg13g2_inv_1 _08965_ (.Y(_03562_),
    .A(_02504_));
 sg13g2_o21ai_1 _08966_ (.B1(_03562_),
    .Y(_03563_),
    .A1(_03547_),
    .A2(_03561_));
 sg13g2_o21ai_1 _08967_ (.B1(_03563_),
    .Y(_03564_),
    .A1(_02773_),
    .A2(_03528_));
 sg13g2_a221oi_1 _08968_ (.B2(_03500_),
    .C1(_03564_),
    .B1(_02883_),
    .A1(_02779_),
    .Y(_03565_),
    .A2(_03473_));
 sg13g2_nand3_1 _08969_ (.B(_03457_),
    .C(_03565_),
    .A(_03431_),
    .Y(_03566_));
 sg13g2_nand2_1 _08970_ (.Y(_03567_),
    .A(_02926_),
    .B(_02561_));
 sg13g2_buf_2 _08971_ (.A(_03567_),
    .X(_03568_));
 sg13g2_a21oi_1 _08972_ (.A1(net115),
    .A2(_03568_),
    .Y(_03569_),
    .B1(net286));
 sg13g2_o21ai_1 _08973_ (.B1(_02959_),
    .Y(_03570_),
    .A1(net136),
    .A2(_03569_));
 sg13g2_nor2_2 _08974_ (.A(net467),
    .B(_02812_),
    .Y(_03571_));
 sg13g2_nor2_1 _08975_ (.A(net392),
    .B(_03571_),
    .Y(_03572_));
 sg13g2_o21ai_1 _08976_ (.B1(net297),
    .Y(_03573_),
    .A1(net115),
    .A2(_03572_));
 sg13g2_nor2_1 _08977_ (.A(_01952_),
    .B(_03474_),
    .Y(_03574_));
 sg13g2_nor2_1 _08978_ (.A(net297),
    .B(_03574_),
    .Y(_03575_));
 sg13g2_nand3_1 _08979_ (.B(_02964_),
    .C(_03575_),
    .A(_03568_),
    .Y(_03576_));
 sg13g2_nand2_1 _08980_ (.Y(_03577_),
    .A(_03573_),
    .B(_03576_));
 sg13g2_a221oi_1 _08981_ (.B2(_03577_),
    .C1(_02953_),
    .B1(net108),
    .A1(net316),
    .Y(_03578_),
    .A2(_03570_));
 sg13g2_or2_1 _08982_ (.X(_03579_),
    .B(_03578_),
    .A(net59));
 sg13g2_o21ai_1 _08983_ (.B1(_03579_),
    .Y(_03580_),
    .A1(_03368_),
    .A2(_03566_));
 sg13g2_nand2_1 _08984_ (.Y(_03581_),
    .A(net230),
    .B(_02578_));
 sg13g2_a21oi_1 _08985_ (.A1(net60),
    .A2(_03581_),
    .Y(_03582_),
    .B1(net386));
 sg13g2_and2_1 _08986_ (.A(net132),
    .B(_03571_),
    .X(_03583_));
 sg13g2_a22oi_1 _08987_ (.Y(_03584_),
    .B1(_03581_),
    .B2(_03583_),
    .A2(net76),
    .A1(net139));
 sg13g2_a22oi_1 _08988_ (.Y(_03585_),
    .B1(_03584_),
    .B2(net87),
    .A2(net81),
    .A1(net215));
 sg13g2_nand3_1 _08989_ (.B(_03568_),
    .C(_03474_),
    .A(net246),
    .Y(_03586_));
 sg13g2_a21oi_1 _08990_ (.A1(_03585_),
    .A2(_03586_),
    .Y(_03587_),
    .B1(net122));
 sg13g2_a22oi_1 _08991_ (.Y(_03588_),
    .B1(_02782_),
    .B2(_03225_),
    .A2(_02860_),
    .A1(net205));
 sg13g2_nor2_2 _08992_ (.A(net285),
    .B(net459),
    .Y(_03589_));
 sg13g2_nand3_1 _08993_ (.B(_03571_),
    .C(_03589_),
    .A(net80),
    .Y(_03590_));
 sg13g2_o21ai_1 _08994_ (.B1(_03590_),
    .Y(_03591_),
    .A1(net87),
    .A2(_03588_));
 sg13g2_a21oi_1 _08995_ (.A1(_02430_),
    .A2(_03591_),
    .Y(_03592_),
    .B1(_01763_));
 sg13g2_nor3_1 _08996_ (.A(_03582_),
    .B(_03587_),
    .C(_03592_),
    .Y(_03593_));
 sg13g2_o21ai_1 _08997_ (.B1(net81),
    .Y(_03594_),
    .A1(net154),
    .A2(net199));
 sg13g2_o21ai_1 _08998_ (.B1(_03594_),
    .Y(_03595_),
    .A1(net140),
    .A2(_03248_));
 sg13g2_nor2_1 _08999_ (.A(net226),
    .B(_02960_),
    .Y(_03596_));
 sg13g2_o21ai_1 _09000_ (.B1(net322),
    .Y(_03597_),
    .A1(_03253_),
    .A2(_03596_));
 sg13g2_nor2_1 _09001_ (.A(net401),
    .B(net80),
    .Y(_03598_));
 sg13g2_a21o_1 _09002_ (.A2(_03598_),
    .A1(_03597_),
    .B1(net375),
    .X(_03599_));
 sg13g2_o21ai_1 _09003_ (.B1(_03599_),
    .Y(_03600_),
    .A1(net134),
    .A2(_03595_));
 sg13g2_o21ai_1 _09004_ (.B1(net253),
    .Y(_03601_),
    .A1(net195),
    .A2(net115));
 sg13g2_a21oi_1 _09005_ (.A1(_02402_),
    .A2(_03601_),
    .Y(_03602_),
    .B1(_01983_));
 sg13g2_nor2_1 _09006_ (.A(_02947_),
    .B(_03602_),
    .Y(_03603_));
 sg13g2_a22oi_1 _09007_ (.Y(_03604_),
    .B1(_03228_),
    .B2(net143),
    .A2(_02939_),
    .A1(_01888_));
 sg13g2_inv_1 _09008_ (.Y(_03605_),
    .A(_03604_));
 sg13g2_a22oi_1 _09009_ (.Y(_03606_),
    .B1(_03605_),
    .B2(net132),
    .A2(net79),
    .A1(net166));
 sg13g2_nand2_1 _09010_ (.Y(_03607_),
    .A(_01931_),
    .B(net99));
 sg13g2_a21oi_1 _09011_ (.A1(net81),
    .A2(_03607_),
    .Y(_03608_),
    .B1(_03193_));
 sg13g2_nor3_1 _09012_ (.A(_03010_),
    .B(_03234_),
    .C(_03608_),
    .Y(_03609_));
 sg13g2_a21o_1 _09013_ (.A2(_03606_),
    .A1(net140),
    .B1(_03609_),
    .X(_03610_));
 sg13g2_nand2_1 _09014_ (.Y(_03611_),
    .A(_03569_),
    .B(_03589_));
 sg13g2_o21ai_1 _09015_ (.B1(_03611_),
    .Y(_03612_),
    .A1(net172),
    .A2(_03588_));
 sg13g2_a21oi_1 _09016_ (.A1(_02430_),
    .A2(_03612_),
    .Y(_03613_),
    .B1(net444));
 sg13g2_a21oi_1 _09017_ (.A1(net108),
    .A2(_03610_),
    .Y(_03614_),
    .B1(_03613_));
 sg13g2_a22oi_1 _09018_ (.Y(_03615_),
    .B1(_03603_),
    .B2(_03614_),
    .A2(_03600_),
    .A1(_03260_));
 sg13g2_o21ai_1 _09019_ (.B1(net446),
    .Y(_03616_),
    .A1(_02322_),
    .A2(_02614_));
 sg13g2_and2_1 _09020_ (.A(net474),
    .B(_03616_),
    .X(_03617_));
 sg13g2_a21oi_1 _09021_ (.A1(net104),
    .A2(_01978_),
    .Y(_03618_),
    .B1(net126));
 sg13g2_nor3_1 _09022_ (.A(net334),
    .B(_01978_),
    .C(_03350_),
    .Y(_03619_));
 sg13g2_nor2_1 _09023_ (.A(net446),
    .B(_03619_),
    .Y(_03620_));
 sg13g2_o21ai_1 _09024_ (.B1(_03620_),
    .Y(_03621_),
    .A1(net58),
    .A2(_03618_));
 sg13g2_o21ai_1 _09025_ (.B1(net335),
    .Y(_03622_),
    .A1(net293),
    .A2(_02781_));
 sg13g2_a221oi_1 _09026_ (.B2(net221),
    .C1(_02408_),
    .B1(_03622_),
    .A1(_02647_),
    .Y(_03623_),
    .A2(_02461_));
 sg13g2_nor2_1 _09027_ (.A(net134),
    .B(_03623_),
    .Y(_03624_));
 sg13g2_o21ai_1 _09028_ (.B1(net179),
    .Y(_03625_),
    .A1(net195),
    .A2(net227));
 sg13g2_a221oi_1 _09029_ (.B2(net119),
    .C1(net238),
    .B1(_03625_),
    .A1(net164),
    .Y(_03626_),
    .A2(_02612_));
 sg13g2_o21ai_1 _09030_ (.B1(net145),
    .Y(_03627_),
    .A1(_03305_),
    .A2(net153));
 sg13g2_a221oi_1 _09031_ (.B2(net164),
    .C1(net226),
    .B1(_03627_),
    .A1(net96),
    .Y(_03628_),
    .A2(net209));
 sg13g2_a21oi_1 _09032_ (.A1(net230),
    .A2(_03272_),
    .Y(_03629_),
    .B1(net120));
 sg13g2_nand2b_1 _09033_ (.Y(_03630_),
    .B(_02867_),
    .A_N(_03629_));
 sg13g2_a21oi_1 _09034_ (.A1(net244),
    .A2(_03012_),
    .Y(_03631_),
    .B1(net221));
 sg13g2_nor2_1 _09035_ (.A(net200),
    .B(net299),
    .Y(_03632_));
 sg13g2_a21oi_1 _09036_ (.A1(net103),
    .A2(_03631_),
    .Y(_03633_),
    .B1(_03632_));
 sg13g2_nor2_1 _09037_ (.A(_03630_),
    .B(_03633_),
    .Y(_03634_));
 sg13g2_nor3_1 _09038_ (.A(_03626_),
    .B(_03628_),
    .C(_03634_),
    .Y(_03635_));
 sg13g2_a22oi_1 _09039_ (.Y(_03636_),
    .B1(_03624_),
    .B2(_03635_),
    .A2(_03621_),
    .A1(_03617_));
 sg13g2_nor2_1 _09040_ (.A(_03292_),
    .B(_03636_),
    .Y(_03637_));
 sg13g2_a21oi_1 _09041_ (.A1(net218),
    .A2(net105),
    .Y(_03638_),
    .B1(net242));
 sg13g2_nand2_1 _09042_ (.Y(_03639_),
    .A(net200),
    .B(net239));
 sg13g2_nand2_1 _09043_ (.Y(_03640_),
    .A(net330),
    .B(_02863_));
 sg13g2_nand3_1 _09044_ (.B(_03639_),
    .C(_03640_),
    .A(net207),
    .Y(_03641_));
 sg13g2_o21ai_1 _09045_ (.B1(_03641_),
    .Y(_03642_),
    .A1(net97),
    .A2(_03638_));
 sg13g2_o21ai_1 _09046_ (.B1(net175),
    .Y(_03643_),
    .A1(net420),
    .A2(_03642_));
 sg13g2_o21ai_1 _09047_ (.B1(net251),
    .Y(_03644_),
    .A1(net201),
    .A2(_02727_));
 sg13g2_a21oi_1 _09048_ (.A1(net288),
    .A2(_02644_),
    .Y(_03645_),
    .B1(_02359_));
 sg13g2_nand2_1 _09049_ (.Y(_03646_),
    .A(net162),
    .B(_03066_));
 sg13g2_nand3_1 _09050_ (.B(_03645_),
    .C(_03646_),
    .A(_03644_),
    .Y(_03647_));
 sg13g2_nand3_1 _09051_ (.B(_03062_),
    .C(_03067_),
    .A(net188),
    .Y(_03648_));
 sg13g2_nand4_1 _09052_ (.B(_03643_),
    .C(_03647_),
    .A(net290),
    .Y(_03649_),
    .D(_03648_));
 sg13g2_a22oi_1 _09053_ (.Y(_03650_),
    .B1(_02847_),
    .B2(net327),
    .A2(_02576_),
    .A1(net429));
 sg13g2_o21ai_1 _09054_ (.B1(_02823_),
    .Y(_03651_),
    .A1(_01771_),
    .A2(_03650_));
 sg13g2_nand3_1 _09055_ (.B(net308),
    .C(net178),
    .A(net89),
    .Y(_03652_));
 sg13g2_o21ai_1 _09056_ (.B1(net232),
    .Y(_03653_),
    .A1(net433),
    .A2(net166));
 sg13g2_nand2_1 _09057_ (.Y(_03654_),
    .A(net387),
    .B(_02339_));
 sg13g2_nand2_1 _09058_ (.Y(_03655_),
    .A(_02733_),
    .B(_03654_));
 sg13g2_a221oi_1 _09059_ (.B2(net129),
    .C1(net301),
    .B1(_03655_),
    .A1(_03066_),
    .Y(_03656_),
    .A2(_03653_));
 sg13g2_a221oi_1 _09060_ (.B2(net188),
    .C1(_03656_),
    .B1(_03652_),
    .A1(net152),
    .Y(_03657_),
    .A2(_03101_));
 sg13g2_nand2b_1 _09061_ (.Y(_03658_),
    .B(_03657_),
    .A_N(_03651_));
 sg13g2_a21oi_1 _09062_ (.A1(_03649_),
    .A2(_03658_),
    .Y(_03659_),
    .B1(_02887_));
 sg13g2_a21oi_1 _09063_ (.A1(net217),
    .A2(_03214_),
    .Y(_03660_),
    .B1(_02511_));
 sg13g2_nand2_1 _09064_ (.Y(_03661_),
    .A(net193),
    .B(_02719_));
 sg13g2_a22oi_1 _09065_ (.Y(_03662_),
    .B1(_03661_),
    .B2(_01930_),
    .A2(_03135_),
    .A1(net289));
 sg13g2_or2_1 _09066_ (.X(_03663_),
    .B(_03662_),
    .A(net77));
 sg13g2_o21ai_1 _09067_ (.B1(_03663_),
    .Y(_03664_),
    .A1(_02988_),
    .A2(_03660_));
 sg13g2_a21oi_1 _09068_ (.A1(_02836_),
    .A2(_03664_),
    .Y(_03665_),
    .B1(net172));
 sg13g2_o21ai_1 _09069_ (.B1(_02386_),
    .Y(_03666_),
    .A1(_02689_),
    .A2(_02909_));
 sg13g2_nand3_1 _09070_ (.B(net224),
    .C(net183),
    .A(_02889_),
    .Y(_03667_));
 sg13g2_o21ai_1 _09071_ (.B1(_03667_),
    .Y(_03668_),
    .A1(net207),
    .A2(_03666_));
 sg13g2_nand2_1 _09072_ (.Y(_03669_),
    .A(net178),
    .B(_03668_));
 sg13g2_a221oi_1 _09073_ (.B2(net188),
    .C1(net134),
    .B1(_03669_),
    .A1(_03346_),
    .Y(_03670_),
    .A2(_03101_));
 sg13g2_nand2b_1 _09074_ (.Y(_03671_),
    .B(_03670_),
    .A_N(_03665_));
 sg13g2_o21ai_1 _09075_ (.B1(_03190_),
    .Y(_03672_),
    .A1(net77),
    .A2(_03012_));
 sg13g2_a21oi_1 _09076_ (.A1(net191),
    .A2(net309),
    .Y(_03673_),
    .B1(_03121_));
 sg13g2_a21oi_1 _09077_ (.A1(net114),
    .A2(_03673_),
    .Y(_03674_),
    .B1(net97));
 sg13g2_o21ai_1 _09078_ (.B1(_03674_),
    .Y(_03675_),
    .A1(net142),
    .A2(_03672_));
 sg13g2_o21ai_1 _09079_ (.B1(net248),
    .Y(_03676_),
    .A1(_02356_),
    .A2(net225));
 sg13g2_nand3_1 _09080_ (.B(_03675_),
    .C(_03676_),
    .A(net228),
    .Y(_03677_));
 sg13g2_nand2_1 _09081_ (.Y(_03678_),
    .A(net121),
    .B(net209));
 sg13g2_nand3_1 _09082_ (.B(net174),
    .C(_03678_),
    .A(net175),
    .Y(_03679_));
 sg13g2_nand3_1 _09083_ (.B(_03679_),
    .C(_03117_),
    .A(_03677_),
    .Y(_03680_));
 sg13g2_a21oi_1 _09084_ (.A1(_03671_),
    .A2(_03680_),
    .Y(_03681_),
    .B1(_02773_));
 sg13g2_nor4_1 _09085_ (.A(_03333_),
    .B(_03637_),
    .C(_03659_),
    .D(_03681_),
    .Y(_03682_));
 sg13g2_o21ai_1 _09086_ (.B1(net119),
    .Y(_03683_),
    .A1(_01926_),
    .A2(_02895_));
 sg13g2_nor2_1 _09087_ (.A(_01936_),
    .B(_03052_),
    .Y(_03684_));
 sg13g2_a21oi_1 _09088_ (.A1(_03683_),
    .A2(_03684_),
    .Y(_03685_),
    .B1(_02366_));
 sg13g2_a21oi_1 _09089_ (.A1(_02712_),
    .A2(_02567_),
    .Y(_03686_),
    .B1(_02517_));
 sg13g2_o21ai_1 _09090_ (.B1(_02381_),
    .Y(_03687_),
    .A1(_02989_),
    .A2(_03686_));
 sg13g2_nand2_1 _09091_ (.Y(_03688_),
    .A(net143),
    .B(net179));
 sg13g2_nand3_1 _09092_ (.B(_03687_),
    .C(_03688_),
    .A(net98),
    .Y(_03689_));
 sg13g2_nand2_1 _09093_ (.Y(_03690_),
    .A(_03685_),
    .B(_03689_));
 sg13g2_o21ai_1 _09094_ (.B1(_01976_),
    .Y(_03691_),
    .A1(net427),
    .A2(_02450_));
 sg13g2_a21oi_1 _09095_ (.A1(net326),
    .A2(_02991_),
    .Y(_03692_),
    .B1(_03691_));
 sg13g2_o21ai_1 _09096_ (.B1(net399),
    .Y(_03693_),
    .A1(net338),
    .A2(net179));
 sg13g2_a21oi_1 _09097_ (.A1(net248),
    .A2(_02564_),
    .Y(_03694_),
    .B1(_03693_));
 sg13g2_nor3_1 _09098_ (.A(net460),
    .B(_03692_),
    .C(_03694_),
    .Y(_03695_));
 sg13g2_nand2_1 _09099_ (.Y(_03696_),
    .A(_03690_),
    .B(_03695_));
 sg13g2_nand2_1 _09100_ (.Y(_03697_),
    .A(net80),
    .B(_02521_));
 sg13g2_nor3_1 _09101_ (.A(net323),
    .B(_02674_),
    .C(net286),
    .Y(_03698_));
 sg13g2_nor2_1 _09102_ (.A(_02520_),
    .B(_02989_),
    .Y(_03699_));
 sg13g2_nor2_1 _09103_ (.A(_02408_),
    .B(net190),
    .Y(_03700_));
 sg13g2_o21ai_1 _09104_ (.B1(_03700_),
    .Y(_03701_),
    .A1(net79),
    .A2(_03699_));
 sg13g2_nor2b_1 _09105_ (.A(_03698_),
    .B_N(_03701_),
    .Y(_03702_));
 sg13g2_nor2_1 _09106_ (.A(_01941_),
    .B(net124),
    .Y(_03703_));
 sg13g2_o21ai_1 _09107_ (.B1(net247),
    .Y(_03704_),
    .A1(net205),
    .A2(_03703_));
 sg13g2_a22oi_1 _09108_ (.Y(_03705_),
    .B1(_03702_),
    .B2(_03704_),
    .A2(_02982_),
    .A1(_03697_));
 sg13g2_o21ai_1 _09109_ (.B1(_01762_),
    .Y(_03706_),
    .A1(net346),
    .A2(_03705_));
 sg13g2_o21ai_1 _09110_ (.B1(_03706_),
    .Y(_03707_),
    .A1(net444),
    .A2(_03696_));
 sg13g2_nand2_1 _09111_ (.Y(_03708_),
    .A(net222),
    .B(_02629_));
 sg13g2_o21ai_1 _09112_ (.B1(_02423_),
    .Y(_03709_),
    .A1(net163),
    .A2(_03708_));
 sg13g2_or2_1 _09113_ (.X(_03710_),
    .B(_02410_),
    .A(net390));
 sg13g2_o21ai_1 _09114_ (.B1(_03710_),
    .Y(_03711_),
    .A1(_02468_),
    .A2(net223));
 sg13g2_a22oi_1 _09115_ (.Y(_03712_),
    .B1(_03711_),
    .B2(net339),
    .A2(_02518_),
    .A1(net303));
 sg13g2_inv_1 _09116_ (.Y(_03713_),
    .A(_03712_));
 sg13g2_a22oi_1 _09117_ (.Y(_03714_),
    .B1(_03713_),
    .B2(_02301_),
    .A2(_03709_),
    .A1(net58));
 sg13g2_nor2_1 _09118_ (.A(net89),
    .B(_03350_),
    .Y(_03715_));
 sg13g2_o21ai_1 _09119_ (.B1(_02820_),
    .Y(_03716_),
    .A1(net95),
    .A2(_03715_));
 sg13g2_o21ai_1 _09120_ (.B1(_03716_),
    .Y(_03717_),
    .A1(_03010_),
    .A2(_03714_));
 sg13g2_nor2_1 _09121_ (.A(net325),
    .B(net299),
    .Y(_03718_));
 sg13g2_nand2_1 _09122_ (.Y(_03719_),
    .A(_02556_),
    .B(_03718_));
 sg13g2_a21oi_1 _09123_ (.A1(net89),
    .A2(_03106_),
    .Y(_03720_),
    .B1(_03719_));
 sg13g2_o21ai_1 _09124_ (.B1(net142),
    .Y(_03721_),
    .A1(net128),
    .A2(_02549_));
 sg13g2_a21oi_1 _09125_ (.A1(net293),
    .A2(net335),
    .Y(_03722_),
    .B1(net333));
 sg13g2_nor2_1 _09126_ (.A(net332),
    .B(net288),
    .Y(_03723_));
 sg13g2_o21ai_1 _09127_ (.B1(net78),
    .Y(_03724_),
    .A1(_03722_),
    .A2(_03723_));
 sg13g2_nand3_1 _09128_ (.B(_03640_),
    .C(_03724_),
    .A(net236),
    .Y(_03725_));
 sg13g2_a221oi_1 _09129_ (.B2(net171),
    .C1(_03392_),
    .B1(_03136_),
    .A1(net210),
    .Y(_03726_),
    .A2(_02976_));
 sg13g2_a22oi_1 _09130_ (.Y(_03727_),
    .B1(_03725_),
    .B2(_03726_),
    .A2(_03721_),
    .A1(_03720_));
 sg13g2_inv_1 _09131_ (.Y(_03728_),
    .A(_03727_));
 sg13g2_a22oi_1 _09132_ (.Y(_03729_),
    .B1(_03728_),
    .B2(_02779_),
    .A2(_03717_),
    .A1(_02828_));
 sg13g2_inv_1 _09133_ (.Y(_03730_),
    .A(_03729_));
 sg13g2_a22oi_1 _09134_ (.Y(_03731_),
    .B1(_03730_),
    .B2(net108),
    .A2(_03707_),
    .A1(_02978_));
 sg13g2_nand3_1 _09135_ (.B(net179),
    .C(_02682_),
    .A(net98),
    .Y(_03732_));
 sg13g2_nand2_1 _09136_ (.Y(_03733_),
    .A(_02706_),
    .B(_03092_));
 sg13g2_a221oi_1 _09137_ (.B2(_03733_),
    .C1(net149),
    .B1(_03732_),
    .A1(net88),
    .Y(_03734_),
    .A2(net176));
 sg13g2_nand2_1 _09138_ (.Y(_03735_),
    .A(net332),
    .B(_02297_));
 sg13g2_a22oi_1 _09139_ (.Y(_03736_),
    .B1(_03735_),
    .B2(net228),
    .A2(_02642_),
    .A1(_02760_));
 sg13g2_a22oi_1 _09140_ (.Y(_03737_),
    .B1(net102),
    .B2(_01937_),
    .A2(_03083_),
    .A1(_03230_));
 sg13g2_nand2_1 _09141_ (.Y(_03738_),
    .A(_03505_),
    .B(_03737_));
 sg13g2_o21ai_1 _09142_ (.B1(_03738_),
    .Y(_03739_),
    .A1(_02343_),
    .A2(_03736_));
 sg13g2_o21ai_1 _09143_ (.B1(_02922_),
    .Y(_03740_),
    .A1(_03734_),
    .A2(_03739_));
 sg13g2_nor2_2 _09144_ (.A(net394),
    .B(net383),
    .Y(_03741_));
 sg13g2_nor2_1 _09145_ (.A(net137),
    .B(_03741_),
    .Y(_03742_));
 sg13g2_o21ai_1 _09146_ (.B1(net301),
    .Y(_03743_),
    .A1(_03324_),
    .A2(_03742_));
 sg13g2_nand2_1 _09147_ (.Y(_03744_),
    .A(_02368_),
    .B(_02601_));
 sg13g2_o21ai_1 _09148_ (.B1(_03744_),
    .Y(_03745_),
    .A1(net166),
    .A2(net102));
 sg13g2_a21oi_1 _09149_ (.A1(net222),
    .A2(net307),
    .Y(_03746_),
    .B1(_02601_));
 sg13g2_o21ai_1 _09150_ (.B1(_02900_),
    .Y(_03747_),
    .A1(net166),
    .A2(_03746_));
 sg13g2_nand2b_1 _09151_ (.Y(_03748_),
    .B(_03220_),
    .A_N(_03747_));
 sg13g2_o21ai_1 _09152_ (.B1(_03748_),
    .Y(_03749_),
    .A1(_03743_),
    .A2(_03745_));
 sg13g2_a21oi_1 _09153_ (.A1(_03200_),
    .A2(_03749_),
    .Y(_03750_),
    .B1(_02660_));
 sg13g2_a21oi_1 _09154_ (.A1(net60),
    .A2(net102),
    .Y(_03751_),
    .B1(net386));
 sg13g2_or2_1 _09155_ (.X(_03752_),
    .B(_03751_),
    .A(_02504_));
 sg13g2_nor2_1 _09156_ (.A(_03750_),
    .B(_03752_),
    .Y(_03753_));
 sg13g2_o21ai_1 _09157_ (.B1(net145),
    .Y(_03754_),
    .A1(net203),
    .A2(_03106_));
 sg13g2_o21ai_1 _09158_ (.B1(_02291_),
    .Y(_03755_),
    .A1(net138),
    .A2(_02871_));
 sg13g2_a22oi_1 _09159_ (.Y(_03756_),
    .B1(_03755_),
    .B2(net121),
    .A2(_03754_),
    .A1(_01932_));
 sg13g2_nand2_2 _09160_ (.Y(_03757_),
    .A(_02375_),
    .B(net231));
 sg13g2_nand2_1 _09161_ (.Y(_03758_),
    .A(net311),
    .B(_02613_));
 sg13g2_o21ai_1 _09162_ (.B1(_03758_),
    .Y(_03759_),
    .A1(net254),
    .A2(_03757_));
 sg13g2_and2_1 _09163_ (.A(net250),
    .B(_03759_),
    .X(_03760_));
 sg13g2_nor4_1 _09164_ (.A(net247),
    .B(_02749_),
    .C(_03760_),
    .D(_03286_),
    .Y(_03761_));
 sg13g2_a21oi_1 _09165_ (.A1(net117),
    .A2(_03756_),
    .Y(_03762_),
    .B1(_03761_));
 sg13g2_o21ai_1 _09166_ (.B1(_03393_),
    .Y(_03763_),
    .A1(net162),
    .A2(_02626_));
 sg13g2_nor2_1 _09167_ (.A(net137),
    .B(_02570_),
    .Y(_03764_));
 sg13g2_nor2_1 _09168_ (.A(_02651_),
    .B(_03764_),
    .Y(_03765_));
 sg13g2_a22oi_1 _09169_ (.Y(_03766_),
    .B1(_03765_),
    .B2(_02443_),
    .A2(_03763_),
    .A1(net118));
 sg13g2_nor2_1 _09170_ (.A(_02842_),
    .B(_02625_),
    .Y(_03767_));
 sg13g2_nor2_1 _09171_ (.A(net250),
    .B(_03767_),
    .Y(_03768_));
 sg13g2_nand2_1 _09172_ (.Y(_03769_),
    .A(net222),
    .B(_02377_));
 sg13g2_a21oi_1 _09173_ (.A1(net155),
    .A2(net137),
    .Y(_03770_),
    .B1(_02763_));
 sg13g2_a22oi_1 _09174_ (.Y(_03771_),
    .B1(_03769_),
    .B2(_03770_),
    .A2(_03768_),
    .A1(_03758_));
 sg13g2_a21oi_1 _09175_ (.A1(net228),
    .A2(_03771_),
    .Y(_03772_),
    .B1(_03266_));
 sg13g2_o21ai_1 _09176_ (.B1(_03772_),
    .Y(_03773_),
    .A1(_02737_),
    .A2(_03766_));
 sg13g2_o21ai_1 _09177_ (.B1(_03773_),
    .Y(_03774_),
    .A1(_03283_),
    .A2(_03762_));
 sg13g2_o21ai_1 _09178_ (.B1(_03206_),
    .Y(_03775_),
    .A1(net88),
    .A2(_02535_));
 sg13g2_o21ai_1 _09179_ (.B1(_01931_),
    .Y(_03776_),
    .A1(net77),
    .A2(_03214_));
 sg13g2_o21ai_1 _09180_ (.B1(net97),
    .Y(_03777_),
    .A1(_02568_),
    .A2(_02473_));
 sg13g2_nand4_1 _09181_ (.B(_02924_),
    .C(_03776_),
    .A(net121),
    .Y(_03778_),
    .D(_03777_));
 sg13g2_o21ai_1 _09182_ (.B1(_03778_),
    .Y(_03779_),
    .A1(net139),
    .A2(_03775_));
 sg13g2_nor2_1 _09183_ (.A(net244),
    .B(_03741_),
    .Y(_03780_));
 sg13g2_o21ai_1 _09184_ (.B1(_03160_),
    .Y(_03781_),
    .A1(net250),
    .A2(_03780_));
 sg13g2_a22oi_1 _09185_ (.Y(_03782_),
    .B1(_03781_),
    .B2(net245),
    .A2(_02667_),
    .A1(net100));
 sg13g2_a21oi_1 _09186_ (.A1(_02667_),
    .A2(_03230_),
    .Y(_03783_),
    .B1(_03361_));
 sg13g2_inv_1 _09187_ (.Y(_03784_),
    .A(_03783_));
 sg13g2_o21ai_1 _09188_ (.B1(net113),
    .Y(_03785_),
    .A1(_02379_),
    .A2(net231));
 sg13g2_a22oi_1 _09189_ (.Y(_03786_),
    .B1(_03785_),
    .B2(net118),
    .A2(_03784_),
    .A1(net90));
 sg13g2_o21ai_1 _09190_ (.B1(_03786_),
    .Y(_03787_),
    .A1(_02527_),
    .A2(_03782_));
 sg13g2_a22oi_1 _09191_ (.Y(_03788_),
    .B1(_03787_),
    .B2(_02828_),
    .A2(_03779_),
    .A1(_02779_));
 sg13g2_nor2_1 _09192_ (.A(net185),
    .B(_03788_),
    .Y(_03789_));
 sg13g2_a221oi_1 _09193_ (.B2(_02883_),
    .C1(_03789_),
    .B1(_03774_),
    .A1(_03740_),
    .Y(_03790_),
    .A2(_03753_));
 sg13g2_nand4_1 _09194_ (.B(_03682_),
    .C(_03731_),
    .A(_03615_),
    .Y(_03791_),
    .D(_03790_));
 sg13g2_o21ai_1 _09195_ (.B1(_03791_),
    .Y(_03792_),
    .A1(net59),
    .A2(_03593_));
 sg13g2_mux4_1 _09196_ (.S0(_01892_),
    .A0(_02975_),
    .A1(_03342_),
    .A2(_03580_),
    .A3(_03792_),
    .S1(net469),
    .X(_03793_));
 sg13g2_nand2b_1 _09197_ (.Y(_03794_),
    .B(_03793_),
    .A_N(_01890_));
 sg13g2_nor2b_1 _09198_ (.A(net422),
    .B_N(net380),
    .Y(_03795_));
 sg13g2_o21ai_1 _09199_ (.B1(net243),
    .Y(_03796_),
    .A1(net289),
    .A2(net223));
 sg13g2_o21ai_1 _09200_ (.B1(net212),
    .Y(_03797_),
    .A1(net340),
    .A2(_02297_));
 sg13g2_a21oi_1 _09201_ (.A1(net179),
    .A2(_02439_),
    .Y(_03798_),
    .B1(net218));
 sg13g2_a221oi_1 _09202_ (.B2(net195),
    .C1(_03798_),
    .B1(_03797_),
    .A1(_03795_),
    .Y(_03799_),
    .A2(_03796_));
 sg13g2_o21ai_1 _09203_ (.B1(net175),
    .Y(_03800_),
    .A1(net420),
    .A2(_03799_));
 sg13g2_a221oi_1 _09204_ (.B2(net213),
    .C1(net341),
    .B1(_01786_),
    .A1(net334),
    .Y(_03801_),
    .A2(net244));
 sg13g2_a21o_1 _09205_ (.A2(_02304_),
    .A1(net345),
    .B1(net240),
    .X(_03802_));
 sg13g2_a21oi_1 _09206_ (.A1(net193),
    .A2(net338),
    .Y(_03803_),
    .B1(net333));
 sg13g2_o21ai_1 _09207_ (.B1(net334),
    .Y(_03804_),
    .A1(net177),
    .A2(_03548_));
 sg13g2_o21ai_1 _09208_ (.B1(_03804_),
    .Y(_03805_),
    .A1(net334),
    .A2(_03803_));
 sg13g2_a221oi_1 _09209_ (.B2(net298),
    .C1(net229),
    .B1(_03805_),
    .A1(_03801_),
    .Y(_03806_),
    .A2(_03802_));
 sg13g2_nor2_1 _09210_ (.A(_02445_),
    .B(net176),
    .Y(_03807_));
 sg13g2_a221oi_1 _09211_ (.B2(net324),
    .C1(net192),
    .B1(_03417_),
    .A1(net170),
    .Y(_03808_),
    .A2(_03387_));
 sg13g2_a21oi_1 _09212_ (.A1(_03069_),
    .A2(_03807_),
    .Y(_03809_),
    .B1(_03808_));
 sg13g2_a22oi_1 _09213_ (.Y(_03810_),
    .B1(_03809_),
    .B2(_03422_),
    .A2(_03806_),
    .A1(_03800_));
 sg13g2_o21ai_1 _09214_ (.B1(net59),
    .Y(_03811_),
    .A1(_02887_),
    .A2(_03810_));
 sg13g2_a22oi_1 _09215_ (.Y(_03812_),
    .B1(_03571_),
    .B2(_02526_),
    .A2(_02955_),
    .A1(net76));
 sg13g2_a21oi_1 _09216_ (.A1(net154),
    .A2(net174),
    .Y(_03813_),
    .B1(_03812_));
 sg13g2_o21ai_1 _09217_ (.B1(_03379_),
    .Y(_03814_),
    .A1(net149),
    .A2(_03813_));
 sg13g2_nor2_1 _09218_ (.A(_01901_),
    .B(net112),
    .Y(_03815_));
 sg13g2_nand2_1 _09219_ (.Y(_03816_),
    .A(net236),
    .B(_02812_));
 sg13g2_nor2_1 _09220_ (.A(net433),
    .B(_03037_),
    .Y(_03817_));
 sg13g2_nor3_1 _09221_ (.A(net336),
    .B(net115),
    .C(_03817_),
    .Y(_03818_));
 sg13g2_a22oi_1 _09222_ (.Y(_03819_),
    .B1(_03816_),
    .B2(_03818_),
    .A2(_03815_),
    .A1(_03589_));
 sg13g2_nand2b_1 _09223_ (.Y(_03820_),
    .B(net290),
    .A_N(_03819_));
 sg13g2_a21oi_1 _09224_ (.A1(_03814_),
    .A2(_03820_),
    .Y(_03821_),
    .B1(_02664_));
 sg13g2_nand2_1 _09225_ (.Y(_03822_),
    .A(_02436_),
    .B(_03127_));
 sg13g2_o21ai_1 _09226_ (.B1(net128),
    .Y(_03823_),
    .A1(net216),
    .A2(net107));
 sg13g2_a21oi_1 _09227_ (.A1(_02653_),
    .A2(_03823_),
    .Y(_03824_),
    .B1(net100));
 sg13g2_nand2b_1 _09228_ (.Y(_03825_),
    .B(net305),
    .A_N(_03083_));
 sg13g2_nand2_1 _09229_ (.Y(_03826_),
    .A(_03150_),
    .B(_03464_));
 sg13g2_a22oi_1 _09230_ (.Y(_03827_),
    .B1(_03826_),
    .B2(net303),
    .A2(_03655_),
    .A1(net378));
 sg13g2_nand4_1 _09231_ (.B(net163),
    .C(_03825_),
    .A(_03028_),
    .Y(_03828_),
    .D(_03827_));
 sg13g2_nand3_1 _09232_ (.B(net170),
    .C(net181),
    .A(_01919_),
    .Y(_03829_));
 sg13g2_a22oi_1 _09233_ (.Y(_03830_),
    .B1(_03829_),
    .B2(_03266_),
    .A2(_03828_),
    .A1(net175));
 sg13g2_o21ai_1 _09234_ (.B1(_03830_),
    .Y(_03831_),
    .A1(_03822_),
    .A2(_03824_));
 sg13g2_nor2_1 _09235_ (.A(_02688_),
    .B(_02744_),
    .Y(_03832_));
 sg13g2_nand2_1 _09236_ (.Y(_03833_),
    .A(net326),
    .B(_02864_));
 sg13g2_nand2b_1 _09237_ (.Y(_03834_),
    .B(_03833_),
    .A_N(_03832_));
 sg13g2_a22oi_1 _09238_ (.Y(_03835_),
    .B1(_03834_),
    .B2(_02988_),
    .A2(_03083_),
    .A1(net112));
 sg13g2_and2_1 _09239_ (.A(net292),
    .B(_03496_),
    .X(_03836_));
 sg13g2_o21ai_1 _09240_ (.B1(_03836_),
    .Y(_03837_),
    .A1(net58),
    .A2(_03835_));
 sg13g2_o21ai_1 _09241_ (.B1(net216),
    .Y(_03838_),
    .A1(_03012_),
    .A2(_03699_));
 sg13g2_nor2_1 _09242_ (.A(net374),
    .B(_01918_),
    .Y(_03839_));
 sg13g2_o21ai_1 _09243_ (.B1(net170),
    .Y(_03840_),
    .A1(_03723_),
    .A2(_03839_));
 sg13g2_nand3_1 _09244_ (.B(_03838_),
    .C(_03840_),
    .A(_02436_),
    .Y(_03841_));
 sg13g2_nor2_1 _09245_ (.A(net119),
    .B(net216),
    .Y(_03842_));
 sg13g2_o21ai_1 _09246_ (.B1(net175),
    .Y(_03843_),
    .A1(_03107_),
    .A2(_03842_));
 sg13g2_nand4_1 _09247_ (.B(_03837_),
    .C(_03841_),
    .A(net290),
    .Y(_03844_),
    .D(_03843_));
 sg13g2_a21oi_1 _09248_ (.A1(_03831_),
    .A2(_03844_),
    .Y(_03845_),
    .B1(_02773_));
 sg13g2_nor2_1 _09249_ (.A(net387),
    .B(_02456_),
    .Y(_03846_));
 sg13g2_a21oi_1 _09250_ (.A1(net323),
    .A2(_02453_),
    .Y(_03847_),
    .B1(_03846_));
 sg13g2_nand3_1 _09251_ (.B(net302),
    .C(_02453_),
    .A(net372),
    .Y(_03848_));
 sg13g2_o21ai_1 _09252_ (.B1(_03848_),
    .Y(_03849_),
    .A1(net336),
    .A2(_03847_));
 sg13g2_and2_1 _09253_ (.A(net152),
    .B(_03849_),
    .X(_03850_));
 sg13g2_inv_1 _09254_ (.Y(_03851_),
    .A(_02456_));
 sg13g2_a22oi_1 _09255_ (.Y(_03852_),
    .B1(_02453_),
    .B2(net116),
    .A2(_03851_),
    .A1(net150));
 sg13g2_o21ai_1 _09256_ (.B1(_03043_),
    .Y(_03853_),
    .A1(net136),
    .A2(_03852_));
 sg13g2_o21ai_1 _09257_ (.B1(net109),
    .Y(_03854_),
    .A1(_03850_),
    .A2(_03853_));
 sg13g2_nand2_1 _09258_ (.Y(_03855_),
    .A(net251),
    .B(net304));
 sg13g2_o21ai_1 _09259_ (.B1(_03855_),
    .Y(_03856_),
    .A1(net419),
    .A2(net251));
 sg13g2_a221oi_1 _09260_ (.B2(net165),
    .C1(net282),
    .B1(_03856_),
    .A1(net177),
    .Y(_03857_),
    .A2(net176));
 sg13g2_a21oi_1 _09261_ (.A1(net214),
    .A2(net102),
    .Y(_03858_),
    .B1(_03005_));
 sg13g2_o21ai_1 _09262_ (.B1(net282),
    .Y(_03859_),
    .A1(net286),
    .A2(_03858_));
 sg13g2_nor2b_1 _09263_ (.A(_03857_),
    .B_N(_03859_),
    .Y(_03860_));
 sg13g2_o21ai_1 _09264_ (.B1(net120),
    .Y(_03861_),
    .A1(net168),
    .A2(_03548_));
 sg13g2_o21ai_1 _09265_ (.B1(_03861_),
    .Y(_03862_),
    .A1(net105),
    .A2(_03803_));
 sg13g2_a21oi_1 _09266_ (.A1(_02556_),
    .A2(_03530_),
    .Y(_03863_),
    .B1(net332));
 sg13g2_o21ai_1 _09267_ (.B1(_03204_),
    .Y(_03864_),
    .A1(_03203_),
    .A2(_03863_));
 sg13g2_a221oi_1 _09268_ (.B2(net320),
    .C1(net460),
    .B1(_03864_),
    .A1(net292),
    .Y(_03865_),
    .A2(_03862_));
 sg13g2_o21ai_1 _09269_ (.B1(_03865_),
    .Y(_03866_),
    .A1(net237),
    .A2(_03860_));
 sg13g2_nand2_1 _09270_ (.Y(_03867_),
    .A(net375),
    .B(_03866_));
 sg13g2_and3_1 _09271_ (.X(_03868_),
    .A(_03009_),
    .B(_03854_),
    .C(_03867_));
 sg13g2_or4_1 _09272_ (.A(_03811_),
    .B(_03821_),
    .C(_03845_),
    .D(_03868_),
    .X(_03869_));
 sg13g2_and2_1 _09273_ (.A(_02417_),
    .B(_02896_),
    .X(_03870_));
 sg13g2_a21oi_1 _09274_ (.A1(_02622_),
    .A2(_03870_),
    .Y(_03871_),
    .B1(net185));
 sg13g2_a22oi_1 _09275_ (.Y(_03872_),
    .B1(_03475_),
    .B2(_02301_),
    .A2(_02684_),
    .A1(net245));
 sg13g2_a21oi_1 _09276_ (.A1(net227),
    .A2(_03175_),
    .Y(_03873_),
    .B1(net90));
 sg13g2_a221oi_1 _09277_ (.B2(net82),
    .C1(_03873_),
    .B1(_03872_),
    .A1(net376),
    .Y(_03874_),
    .A2(_03832_));
 sg13g2_a21oi_1 _09278_ (.A1(net90),
    .A2(net295),
    .Y(_03875_),
    .B1(_01786_));
 sg13g2_o21ai_1 _09279_ (.B1(net113),
    .Y(_03876_),
    .A1(net58),
    .A2(_03875_));
 sg13g2_a22oi_1 _09280_ (.Y(_03877_),
    .B1(_03876_),
    .B2(net171),
    .A2(_03874_),
    .A1(net139));
 sg13g2_o21ai_1 _09281_ (.B1(_03022_),
    .Y(_03878_),
    .A1(_03389_),
    .A2(_02757_));
 sg13g2_nand2_1 _09282_ (.Y(_03879_),
    .A(net297),
    .B(_03878_));
 sg13g2_nand2_1 _09283_ (.Y(_03880_),
    .A(_03076_),
    .B(net167));
 sg13g2_nand2_1 _09284_ (.Y(_03881_),
    .A(_03139_),
    .B(_02752_));
 sg13g2_nand3_1 _09285_ (.B(_03880_),
    .C(_03881_),
    .A(_01900_),
    .Y(_03882_));
 sg13g2_nand2_1 _09286_ (.Y(_03883_),
    .A(net131),
    .B(_03390_));
 sg13g2_o21ai_1 _09287_ (.B1(_03883_),
    .Y(_03884_),
    .A1(net100),
    .A2(_03882_));
 sg13g2_nor2_1 _09288_ (.A(net78),
    .B(_02398_),
    .Y(_03885_));
 sg13g2_nand2_1 _09289_ (.Y(_03886_),
    .A(net163),
    .B(_02945_));
 sg13g2_o21ai_1 _09290_ (.B1(net210),
    .Y(_03887_),
    .A1(_03885_),
    .A2(_03886_));
 sg13g2_o21ai_1 _09291_ (.B1(_03887_),
    .Y(_03888_),
    .A1(_01938_),
    .A2(_03884_));
 sg13g2_nor2_1 _09292_ (.A(net325),
    .B(net225),
    .Y(_03889_));
 sg13g2_o21ai_1 _09293_ (.B1(net82),
    .Y(_03890_),
    .A1(_01889_),
    .A2(_02398_));
 sg13g2_nand2_1 _09294_ (.Y(_03891_),
    .A(_03214_),
    .B(_03469_));
 sg13g2_nand2_1 _09295_ (.Y(_03892_),
    .A(net419),
    .B(_03121_));
 sg13g2_nand4_1 _09296_ (.B(_03890_),
    .C(_03891_),
    .A(_03889_),
    .Y(_03893_),
    .D(_03892_));
 sg13g2_o21ai_1 _09297_ (.B1(_03893_),
    .Y(_03894_),
    .A1(_03879_),
    .A2(_03888_));
 sg13g2_a22oi_1 _09298_ (.Y(_03895_),
    .B1(_03894_),
    .B2(_02922_),
    .A2(_03877_),
    .A1(_03871_));
 sg13g2_nor2_1 _09299_ (.A(_03386_),
    .B(_03895_),
    .Y(_03896_));
 sg13g2_nand2_1 _09300_ (.Y(_03897_),
    .A(net135),
    .B(_02682_));
 sg13g2_a221oi_1 _09301_ (.B2(net78),
    .C1(net226),
    .B1(_03897_),
    .A1(_01919_),
    .Y(_03898_),
    .A2(_02452_));
 sg13g2_o21ai_1 _09302_ (.B1(net250),
    .Y(_03899_),
    .A1(_02300_),
    .A2(_03214_));
 sg13g2_nor3_1 _09303_ (.A(net334),
    .B(net189),
    .C(_02892_),
    .Y(_03900_));
 sg13g2_a221oi_1 _09304_ (.B2(_03900_),
    .C1(_01912_),
    .B1(_03899_),
    .A1(net150),
    .Y(_03901_),
    .A2(_02713_));
 sg13g2_nand2_1 _09305_ (.Y(_03902_),
    .A(net120),
    .B(_03014_));
 sg13g2_nor2_1 _09306_ (.A(_01959_),
    .B(net333),
    .Y(_03903_));
 sg13g2_and2_1 _09307_ (.A(_03902_),
    .B(_03903_),
    .X(_03904_));
 sg13g2_nor2_1 _09308_ (.A(net342),
    .B(_03300_),
    .Y(_03905_));
 sg13g2_a21oi_1 _09309_ (.A1(_02842_),
    .A2(net284),
    .Y(_03906_),
    .B1(_03905_));
 sg13g2_a21oi_1 _09310_ (.A1(_02522_),
    .A2(_02989_),
    .Y(_03907_),
    .B1(net127));
 sg13g2_mux2_1 _09311_ (.A0(_03906_),
    .A1(_03907_),
    .S(_02717_),
    .X(_03908_));
 sg13g2_a221oi_1 _09312_ (.B2(_03908_),
    .C1(_01937_),
    .B1(_03904_),
    .A1(net301),
    .Y(_03909_),
    .A2(net201));
 sg13g2_nor4_1 _09313_ (.A(net401),
    .B(_03898_),
    .C(_03901_),
    .D(_03909_),
    .Y(_03910_));
 sg13g2_a21o_1 _09314_ (.A2(_03466_),
    .A1(_02593_),
    .B1(_03910_),
    .X(_03911_));
 sg13g2_a21o_1 _09315_ (.A2(_03518_),
    .A1(net121),
    .B1(_03063_),
    .X(_03912_));
 sg13g2_a22oi_1 _09316_ (.Y(_03913_),
    .B1(_03912_),
    .B2(_02357_),
    .A2(_03817_),
    .A1(_03005_));
 sg13g2_o21ai_1 _09317_ (.B1(_02413_),
    .Y(_03914_),
    .A1(net116),
    .A2(_02375_));
 sg13g2_nand2_1 _09318_ (.Y(_03915_),
    .A(_01932_),
    .B(_03914_));
 sg13g2_o21ai_1 _09319_ (.B1(_02357_),
    .Y(_03916_),
    .A1(net143),
    .A2(_03214_));
 sg13g2_a21oi_1 _09320_ (.A1(_03915_),
    .A2(_03916_),
    .Y(_03917_),
    .B1(net139));
 sg13g2_a21oi_1 _09321_ (.A1(net312),
    .A2(net180),
    .Y(_03918_),
    .B1(_02531_));
 sg13g2_nor2b_1 _09322_ (.A(_03918_),
    .B_N(_03684_),
    .Y(_03919_));
 sg13g2_nor3_1 _09323_ (.A(_02737_),
    .B(_03917_),
    .C(_03919_),
    .Y(_03920_));
 sg13g2_a21oi_1 _09324_ (.A1(_01964_),
    .A2(_03913_),
    .Y(_03921_),
    .B1(_03920_));
 sg13g2_a22oi_1 _09325_ (.Y(_03922_),
    .B1(_03921_),
    .B2(_02830_),
    .A2(_03911_),
    .A1(_01762_));
 sg13g2_nor2_1 _09326_ (.A(_02596_),
    .B(_03922_),
    .Y(_03923_));
 sg13g2_nor2_1 _09327_ (.A(_03305_),
    .B(net153),
    .Y(_03924_));
 sg13g2_nand2_1 _09328_ (.Y(_03925_),
    .A(net373),
    .B(_03924_));
 sg13g2_a221oi_1 _09329_ (.B2(net133),
    .C1(net252),
    .B1(_03925_),
    .A1(net88),
    .Y(_03926_),
    .A2(_03434_));
 sg13g2_a21oi_1 _09330_ (.A1(_01786_),
    .A2(_02322_),
    .Y(_03927_),
    .B1(_03501_));
 sg13g2_nor2_1 _09331_ (.A(net188),
    .B(_03927_),
    .Y(_03928_));
 sg13g2_o21ai_1 _09332_ (.B1(net108),
    .Y(_03929_),
    .A1(_03926_),
    .A2(_03928_));
 sg13g2_a221oi_1 _09333_ (.B2(net164),
    .C1(net126),
    .B1(_03924_),
    .A1(net119),
    .Y(_03930_),
    .A2(net239));
 sg13g2_a21oi_1 _09334_ (.A1(net126),
    .A2(net178),
    .Y(_03931_),
    .B1(_03930_));
 sg13g2_nor2_1 _09335_ (.A(net151),
    .B(_03931_),
    .Y(_03932_));
 sg13g2_a21oi_1 _09336_ (.A1(net180),
    .A2(_03086_),
    .Y(_03933_),
    .B1(net300));
 sg13g2_o21ai_1 _09337_ (.B1(_03137_),
    .Y(_03934_),
    .A1(_02600_),
    .A2(net171));
 sg13g2_nor3_1 _09338_ (.A(_03325_),
    .B(_03933_),
    .C(_03934_),
    .Y(_03935_));
 sg13g2_nor2_1 _09339_ (.A(net421),
    .B(_03935_),
    .Y(_03936_));
 sg13g2_o21ai_1 _09340_ (.B1(_03936_),
    .Y(_03937_),
    .A1(_03322_),
    .A2(_03932_));
 sg13g2_nand3_1 _09341_ (.B(_03929_),
    .C(_03937_),
    .A(_03297_),
    .Y(_03938_));
 sg13g2_nand3_1 _09342_ (.B(_02555_),
    .C(_03225_),
    .A(net138),
    .Y(_03939_));
 sg13g2_o21ai_1 _09343_ (.B1(net253),
    .Y(_03940_),
    .A1(_02923_),
    .A2(net281));
 sg13g2_nand3_1 _09344_ (.B(_03238_),
    .C(_03940_),
    .A(net117),
    .Y(_03941_));
 sg13g2_nand3_1 _09345_ (.B(_03939_),
    .C(_03941_),
    .A(net108),
    .Y(_03942_));
 sg13g2_a22oi_1 _09346_ (.Y(_03943_),
    .B1(_03225_),
    .B2(_02537_),
    .A2(_03142_),
    .A1(_02714_));
 sg13g2_inv_1 _09347_ (.Y(_03944_),
    .A(_03943_));
 sg13g2_nor2_1 _09348_ (.A(net253),
    .B(_03397_),
    .Y(_03945_));
 sg13g2_a22oi_1 _09349_ (.Y(_03946_),
    .B1(_03945_),
    .B2(net205),
    .A2(_03225_),
    .A1(_02782_));
 sg13g2_nor2_1 _09350_ (.A(net237),
    .B(_03946_),
    .Y(_03947_));
 sg13g2_a21oi_1 _09351_ (.A1(_03589_),
    .A2(_03944_),
    .Y(_03948_),
    .B1(_03947_));
 sg13g2_o21ai_1 _09352_ (.B1(net316),
    .Y(_03949_),
    .A1(net424),
    .A2(_03948_));
 sg13g2_nand3_1 _09353_ (.B(_03942_),
    .C(_03949_),
    .A(_03227_),
    .Y(_03950_));
 sg13g2_nor2_1 _09354_ (.A(net300),
    .B(_02853_),
    .Y(_03951_));
 sg13g2_nand2_1 _09355_ (.Y(_03952_),
    .A(net333),
    .B(_01949_));
 sg13g2_nand2_1 _09356_ (.Y(_03953_),
    .A(_02286_),
    .B(_03952_));
 sg13g2_nand3_1 _09357_ (.B(_02835_),
    .C(_03953_),
    .A(net162),
    .Y(_03954_));
 sg13g2_nand3_1 _09358_ (.B(_03568_),
    .C(_02653_),
    .A(net98),
    .Y(_03955_));
 sg13g2_nand3_1 _09359_ (.B(net181),
    .C(_03955_),
    .A(net123),
    .Y(_03956_));
 sg13g2_a21oi_1 _09360_ (.A1(_03951_),
    .A2(_03954_),
    .Y(_03957_),
    .B1(_03956_));
 sg13g2_o21ai_1 _09361_ (.B1(net310),
    .Y(_03958_),
    .A1(_02587_),
    .A2(_01918_));
 sg13g2_nor2_1 _09362_ (.A(net341),
    .B(_03309_),
    .Y(_03959_));
 sg13g2_a221oi_1 _09363_ (.B2(_02786_),
    .C1(_02432_),
    .B1(_03959_),
    .A1(_02435_),
    .Y(_03960_),
    .A2(_03958_));
 sg13g2_o21ai_1 _09364_ (.B1(net340),
    .Y(_03961_),
    .A1(_01967_),
    .A2(_03741_));
 sg13g2_o21ai_1 _09365_ (.B1(_03961_),
    .Y(_03962_),
    .A1(net314),
    .A2(_03294_));
 sg13g2_a21o_1 _09366_ (.A2(net153),
    .A1(net314),
    .B1(_01950_),
    .X(_03963_));
 sg13g2_a22oi_1 _09367_ (.Y(_03964_),
    .B1(_03963_),
    .B2(net176),
    .A2(_03962_),
    .A1(net216));
 sg13g2_nor2_1 _09368_ (.A(net198),
    .B(_03964_),
    .Y(_03965_));
 sg13g2_nor2_1 _09369_ (.A(_03960_),
    .B(_03965_),
    .Y(_03966_));
 sg13g2_nand2_1 _09370_ (.Y(_03967_),
    .A(net319),
    .B(net463));
 sg13g2_o21ai_1 _09371_ (.B1(_03967_),
    .Y(_03968_),
    .A1(_02467_),
    .A2(_03735_));
 sg13g2_a21oi_1 _09372_ (.A1(_02994_),
    .A2(_03968_),
    .Y(_03969_),
    .B1(net459));
 sg13g2_nor2_1 _09373_ (.A(net313),
    .B(_02863_),
    .Y(_03970_));
 sg13g2_nand2_1 _09374_ (.Y(_03971_),
    .A(net141),
    .B(_03513_));
 sg13g2_nand2_1 _09375_ (.Y(_03972_),
    .A(_03970_),
    .B(_03971_));
 sg13g2_nand3_1 _09376_ (.B(_03960_),
    .C(_03972_),
    .A(_03969_),
    .Y(_03973_));
 sg13g2_o21ai_1 _09377_ (.B1(_03973_),
    .Y(_03974_),
    .A1(_02681_),
    .A2(_03966_));
 sg13g2_o21ai_1 _09378_ (.B1(_02883_),
    .Y(_03975_),
    .A1(_03957_),
    .A2(_03974_));
 sg13g2_a21oi_1 _09379_ (.A1(net419),
    .A2(_03121_),
    .Y(_03976_),
    .B1(_03767_));
 sg13g2_a21oi_1 _09380_ (.A1(_02944_),
    .A2(_03976_),
    .Y(_03977_),
    .B1(net232));
 sg13g2_nor2_1 _09381_ (.A(net142),
    .B(net107),
    .Y(_03978_));
 sg13g2_a221oi_1 _09382_ (.B2(_02845_),
    .C1(_02370_),
    .B1(_03978_),
    .A1(net100),
    .Y(_03979_),
    .A2(_02589_));
 sg13g2_inv_1 _09383_ (.Y(_03980_),
    .A(_03654_));
 sg13g2_nand2_1 _09384_ (.Y(_03981_),
    .A(_02584_),
    .B(_02911_));
 sg13g2_and4_1 _09385_ (.A(_02291_),
    .B(_03980_),
    .C(_03902_),
    .D(_03981_),
    .X(_03982_));
 sg13g2_nor4_1 _09386_ (.A(net185),
    .B(_03977_),
    .C(_03979_),
    .D(_03982_),
    .Y(_03983_));
 sg13g2_nand3_1 _09387_ (.B(net191),
    .C(_02373_),
    .A(net218),
    .Y(_03984_));
 sg13g2_o21ai_1 _09388_ (.B1(_03984_),
    .Y(_03985_),
    .A1(net114),
    .A2(_02655_));
 sg13g2_a22oi_1 _09389_ (.Y(_03986_),
    .B1(_03985_),
    .B2(net190),
    .A2(_02580_),
    .A1(_01943_));
 sg13g2_nor3_1 _09390_ (.A(net133),
    .B(_03515_),
    .C(_03654_),
    .Y(_03987_));
 sg13g2_nand2b_1 _09391_ (.Y(_03988_),
    .B(_03881_),
    .A_N(_02757_));
 sg13g2_a221oi_1 _09392_ (.B2(net199),
    .C1(net247),
    .B1(_03988_),
    .A1(net96),
    .Y(_03989_),
    .A2(_03987_));
 sg13g2_o21ai_1 _09393_ (.B1(_03989_),
    .Y(_03990_),
    .A1(_02370_),
    .A2(_03986_));
 sg13g2_o21ai_1 _09394_ (.B1(_02509_),
    .Y(_03991_),
    .A1(net317),
    .A2(_02421_));
 sg13g2_nand3_1 _09395_ (.B(_03153_),
    .C(_03026_),
    .A(_02671_),
    .Y(_03992_));
 sg13g2_a21o_1 _09396_ (.A2(_03991_),
    .A1(_02286_),
    .B1(_03992_),
    .X(_03993_));
 sg13g2_a21oi_1 _09397_ (.A1(_03990_),
    .A2(_03993_),
    .Y(_03994_),
    .B1(_02705_));
 sg13g2_o21ai_1 _09398_ (.B1(_02779_),
    .Y(_03995_),
    .A1(_03983_),
    .A2(_03994_));
 sg13g2_nand4_1 _09399_ (.B(_03950_),
    .C(_03975_),
    .A(_03938_),
    .Y(_03996_),
    .D(_03995_));
 sg13g2_nor4_1 _09400_ (.A(_03869_),
    .B(_03896_),
    .C(_03923_),
    .D(_03996_),
    .Y(_03997_));
 sg13g2_o21ai_1 _09401_ (.B1(_02964_),
    .Y(_03998_),
    .A1(net154),
    .A2(net89));
 sg13g2_a221oi_1 _09402_ (.B2(net87),
    .C1(net122),
    .B1(_03998_),
    .A1(_03241_),
    .Y(_03999_),
    .A2(_03818_));
 sg13g2_nand2_1 _09403_ (.Y(_04000_),
    .A(net297),
    .B(_02430_));
 sg13g2_a21oi_1 _09404_ (.A1(net151),
    .A2(_03607_),
    .Y(_04001_),
    .B1(_04000_));
 sg13g2_a21oi_1 _09405_ (.A1(_03363_),
    .A2(_04001_),
    .Y(_04002_),
    .B1(_01763_));
 sg13g2_nor3_1 _09406_ (.A(_02953_),
    .B(_03999_),
    .C(_04002_),
    .Y(_04003_));
 sg13g2_o21ai_1 _09407_ (.B1(net469),
    .Y(_04004_),
    .A1(net59),
    .A2(_04003_));
 sg13g2_a22oi_1 _09408_ (.Y(_04005_),
    .B1(_03940_),
    .B2(net305),
    .A2(_03242_),
    .A1(net125));
 sg13g2_a21oi_1 _09409_ (.A1(net337),
    .A2(net173),
    .Y(_04006_),
    .B1(net99));
 sg13g2_nor2_1 _09410_ (.A(_02525_),
    .B(_04006_),
    .Y(_04007_));
 sg13g2_nor3_1 _09411_ (.A(net336),
    .B(_03698_),
    .C(_04007_),
    .Y(_04008_));
 sg13g2_a21o_1 _09412_ (.A2(_04005_),
    .A1(net247),
    .B1(_04008_),
    .X(_04009_));
 sg13g2_nor2_1 _09413_ (.A(net325),
    .B(net125),
    .Y(_04010_));
 sg13g2_a221oi_1 _09414_ (.B2(net173),
    .C1(net341),
    .B1(net130),
    .A1(net105),
    .Y(_04011_),
    .A2(net322));
 sg13g2_nor2_1 _09415_ (.A(net328),
    .B(net99),
    .Y(_04012_));
 sg13g2_nand3_1 _09416_ (.B(net423),
    .C(_02624_),
    .A(net432),
    .Y(_04013_));
 sg13g2_buf_1 _09417_ (.A(_04013_),
    .X(_04014_));
 sg13g2_nand3_1 _09418_ (.B(net331),
    .C(_02612_),
    .A(net317),
    .Y(_04015_));
 sg13g2_and3_1 _09419_ (.X(_04016_),
    .A(net296),
    .B(_04014_),
    .C(_04015_));
 sg13g2_o21ai_1 _09420_ (.B1(_02630_),
    .Y(_04017_),
    .A1(_04012_),
    .A2(_04016_));
 sg13g2_a21oi_1 _09421_ (.A1(_03363_),
    .A2(_04017_),
    .Y(_04018_),
    .B1(net336));
 sg13g2_or4_1 _09422_ (.A(_02429_),
    .B(_04010_),
    .C(_04011_),
    .D(_04018_),
    .X(_04019_));
 sg13g2_a22oi_1 _09423_ (.Y(_04020_),
    .B1(_04019_),
    .B2(net375),
    .A2(_04009_),
    .A1(net181));
 sg13g2_nand2_1 _09424_ (.Y(_04021_),
    .A(net235),
    .B(net113));
 sg13g2_o21ai_1 _09425_ (.B1(_04021_),
    .Y(_04022_),
    .A1(net224),
    .A2(_02804_));
 sg13g2_a21oi_1 _09426_ (.A1(net320),
    .A2(_04022_),
    .Y(_04023_),
    .B1(net446));
 sg13g2_a221oi_1 _09427_ (.B2(_02517_),
    .C1(_02340_),
    .B1(_03464_),
    .A1(net389),
    .Y(_04024_),
    .A2(_02991_));
 sg13g2_or3_1 _09428_ (.A(net291),
    .B(_02560_),
    .C(_04024_),
    .X(_04025_));
 sg13g2_nor3_1 _09429_ (.A(net387),
    .B(_02290_),
    .C(_03268_),
    .Y(_04026_));
 sg13g2_nor2_1 _09430_ (.A(net372),
    .B(_04026_),
    .Y(_04027_));
 sg13g2_o21ai_1 _09431_ (.B1(_03285_),
    .Y(_04028_),
    .A1(net222),
    .A2(net101));
 sg13g2_a22oi_1 _09432_ (.Y(_04029_),
    .B1(_03918_),
    .B2(_03769_),
    .A2(_04028_),
    .A1(_02532_));
 sg13g2_a22oi_1 _09433_ (.Y(_04030_),
    .B1(_04029_),
    .B2(net292),
    .A2(_04027_),
    .A1(_04025_));
 sg13g2_o21ai_1 _09434_ (.B1(net190),
    .Y(_04031_),
    .A1(net137),
    .A2(_03121_));
 sg13g2_a22oi_1 _09435_ (.Y(_04032_),
    .B1(_04031_),
    .B2(_02593_),
    .A2(_04030_),
    .A1(_04023_));
 sg13g2_a221oi_1 _09436_ (.B2(net314),
    .C1(net180),
    .B1(_02732_),
    .A1(net244),
    .Y(_04033_),
    .A2(net130));
 sg13g2_mux2_1 _09437_ (.A0(net319),
    .A1(_02576_),
    .S(_01916_),
    .X(_04034_));
 sg13g2_a22oi_1 _09438_ (.Y(_04035_),
    .B1(_04034_),
    .B2(net127),
    .A2(_03757_),
    .A1(net182));
 sg13g2_nand2_1 _09439_ (.Y(_04036_),
    .A(net230),
    .B(net233));
 sg13g2_a221oi_1 _09440_ (.B2(net248),
    .C1(net291),
    .B1(_04036_),
    .A1(net288),
    .Y(_04037_),
    .A2(_03434_));
 sg13g2_a21oi_1 _09441_ (.A1(net339),
    .A2(_04035_),
    .Y(_04038_),
    .B1(_04037_));
 sg13g2_mux2_1 _09442_ (.A0(_04033_),
    .A1(_04038_),
    .S(net285),
    .X(_04039_));
 sg13g2_nand2_1 _09443_ (.Y(_04040_),
    .A(net290),
    .B(_04039_));
 sg13g2_o21ai_1 _09444_ (.B1(_04040_),
    .Y(_04041_),
    .A1(net375),
    .A2(_04032_));
 sg13g2_nand2b_1 _09445_ (.Y(_04042_),
    .B(net462),
    .A_N(net468));
 sg13g2_nand2_1 _09446_ (.Y(_04043_),
    .A(net381),
    .B(_04042_));
 sg13g2_nand2_1 _09447_ (.Y(_04044_),
    .A(net382),
    .B(_01786_));
 sg13g2_nor2_1 _09448_ (.A(net317),
    .B(_02437_),
    .Y(_04045_));
 sg13g2_a221oi_1 _09449_ (.B2(_04045_),
    .C1(net385),
    .B1(_04044_),
    .A1(net294),
    .Y(_04046_),
    .A2(_04043_));
 sg13g2_a22oi_1 _09450_ (.Y(_04047_),
    .B1(_02809_),
    .B2(net389),
    .A2(_02576_),
    .A1(net429));
 sg13g2_o21ai_1 _09451_ (.B1(net296),
    .Y(_04048_),
    .A1(net382),
    .A2(_04047_));
 sg13g2_nand2_1 _09452_ (.Y(_04049_),
    .A(net330),
    .B(net243));
 sg13g2_o21ai_1 _09453_ (.B1(_04049_),
    .Y(_04050_),
    .A1(_04046_),
    .A2(_04048_));
 sg13g2_nand3_1 _09454_ (.B(net182),
    .C(net183),
    .A(net253),
    .Y(_04051_));
 sg13g2_a221oi_1 _09455_ (.B2(net287),
    .C1(_02703_),
    .B1(_04051_),
    .A1(net282),
    .Y(_04052_),
    .A2(_04050_));
 sg13g2_xnor2_1 _09456_ (.Y(_04053_),
    .A(net207),
    .B(_03548_));
 sg13g2_o21ai_1 _09457_ (.B1(net249),
    .Y(_04054_),
    .A1(net164),
    .A2(_04053_));
 sg13g2_mux2_1 _09458_ (.A0(_02296_),
    .A1(_02877_),
    .S(_02470_),
    .X(_04055_));
 sg13g2_a221oi_1 _09459_ (.B2(_02863_),
    .C1(_01953_),
    .B1(_03513_),
    .A1(net378),
    .Y(_04056_),
    .A2(net281));
 sg13g2_a21oi_1 _09460_ (.A1(net313),
    .A2(_04055_),
    .Y(_04057_),
    .B1(_04056_));
 sg13g2_nor2b_1 _09461_ (.A(net381),
    .B_N(net432),
    .Y(_04058_));
 sg13g2_a221oi_1 _09462_ (.B2(net380),
    .C1(net293),
    .B1(_04058_),
    .A1(net461),
    .Y(_04059_),
    .A2(_01948_));
 sg13g2_nor3_1 _09463_ (.A(_02288_),
    .B(net338),
    .C(_02809_),
    .Y(_04060_));
 sg13g2_or3_1 _09464_ (.A(net391),
    .B(_04059_),
    .C(_04060_),
    .X(_04061_));
 sg13g2_o21ai_1 _09465_ (.B1(_04061_),
    .Y(_04062_),
    .A1(net323),
    .A2(_04057_));
 sg13g2_a21oi_1 _09466_ (.A1(net324),
    .A2(_04062_),
    .Y(_04063_),
    .B1(_02432_));
 sg13g2_nand2_1 _09467_ (.Y(_04064_),
    .A(net425),
    .B(net189));
 sg13g2_o21ai_1 _09468_ (.B1(_04064_),
    .Y(_04065_),
    .A1(net310),
    .A2(net189));
 sg13g2_o21ai_1 _09469_ (.B1(net311),
    .Y(_04066_),
    .A1(_01786_),
    .A2(_02447_));
 sg13g2_and2_1 _09470_ (.A(_03970_),
    .B(_04066_),
    .X(_04067_));
 sg13g2_a221oi_1 _09471_ (.B2(_03285_),
    .C1(_02748_),
    .B1(_04067_),
    .A1(net131),
    .Y(_04068_),
    .A2(_04065_));
 sg13g2_a22oi_1 _09472_ (.Y(_04069_),
    .B1(_04063_),
    .B2(_04068_),
    .A2(_04054_),
    .A1(_04052_));
 sg13g2_o21ai_1 _09473_ (.B1(net172),
    .Y(_04070_),
    .A1(_04052_),
    .A2(_04063_));
 sg13g2_a21oi_1 _09474_ (.A1(_04069_),
    .A2(_04070_),
    .Y(_04071_),
    .B1(_02773_));
 sg13g2_a221oi_1 _09475_ (.B2(_03456_),
    .C1(_04071_),
    .B1(_04041_),
    .A1(_03227_),
    .Y(_04072_),
    .A2(_04020_));
 sg13g2_a21oi_1 _09476_ (.A1(_03746_),
    .A2(_03229_),
    .Y(_04073_),
    .B1(_03574_));
 sg13g2_a221oi_1 _09477_ (.B2(_02731_),
    .C1(net336),
    .B1(net176),
    .A1(_02285_),
    .Y(_04074_),
    .A2(net204));
 sg13g2_a21oi_1 _09478_ (.A1(net280),
    .A2(_04073_),
    .Y(_04075_),
    .B1(_04074_));
 sg13g2_o21ai_1 _09479_ (.B1(_01761_),
    .Y(_04076_),
    .A1(_01755_),
    .A2(_04075_));
 sg13g2_nand2_1 _09480_ (.Y(_04077_),
    .A(net223),
    .B(_03208_));
 sg13g2_a21oi_1 _09481_ (.A1(_02383_),
    .A2(_03555_),
    .Y(_04078_),
    .B1(net203));
 sg13g2_nor3_1 _09482_ (.A(_04077_),
    .B(_03933_),
    .C(_04078_),
    .Y(_04079_));
 sg13g2_nand3_1 _09483_ (.B(net243),
    .C(net169),
    .A(net242),
    .Y(_04080_));
 sg13g2_nand2_1 _09484_ (.Y(_04081_),
    .A(net295),
    .B(_02511_));
 sg13g2_a221oi_1 _09485_ (.B2(net298),
    .C1(net229),
    .B1(_04081_),
    .A1(_02840_),
    .Y(_04082_),
    .A2(_04080_));
 sg13g2_o21ai_1 _09486_ (.B1(_04082_),
    .Y(_04083_),
    .A1(net206),
    .A2(_04079_));
 sg13g2_nand2_1 _09487_ (.Y(_04084_),
    .A(_04076_),
    .B(_04083_));
 sg13g2_nor2_1 _09488_ (.A(net193),
    .B(_02517_),
    .Y(_04085_));
 sg13g2_a221oi_1 _09489_ (.B2(_02785_),
    .C1(net314),
    .B1(_04085_),
    .A1(net165),
    .Y(_04086_),
    .A2(net419));
 sg13g2_o21ai_1 _09490_ (.B1(net291),
    .Y(_04087_),
    .A1(net337),
    .A2(net178));
 sg13g2_a21oi_1 _09491_ (.A1(net224),
    .A2(_02453_),
    .Y(_04088_),
    .B1(_04087_));
 sg13g2_or3_1 _09492_ (.A(net324),
    .B(_04086_),
    .C(_04088_),
    .X(_04089_));
 sg13g2_nand2_1 _09493_ (.Y(_04090_),
    .A(net340),
    .B(net284));
 sg13g2_o21ai_1 _09494_ (.B1(_04090_),
    .Y(_04091_),
    .A1(net194),
    .A2(_03757_));
 sg13g2_nand3_1 _09495_ (.B(net137),
    .C(net307),
    .A(net248),
    .Y(_04092_));
 sg13g2_nand2_1 _09496_ (.Y(_04093_),
    .A(net235),
    .B(_03159_));
 sg13g2_nand3_1 _09497_ (.B(_04092_),
    .C(_04093_),
    .A(_03115_),
    .Y(_04094_));
 sg13g2_a221oi_1 _09498_ (.B2(net292),
    .C1(net446),
    .B1(_04094_),
    .A1(net320),
    .Y(_04095_),
    .A2(_04091_));
 sg13g2_a22oi_1 _09499_ (.Y(_04096_),
    .B1(_04089_),
    .B2(_04095_),
    .A2(_02593_),
    .A1(_03005_));
 sg13g2_nand2_1 _09500_ (.Y(_04097_),
    .A(_02561_),
    .B(_03159_));
 sg13g2_o21ai_1 _09501_ (.B1(net101),
    .Y(_04098_),
    .A1(net332),
    .A2(_01971_));
 sg13g2_and2_1 _09502_ (.A(_04097_),
    .B(_04098_),
    .X(_04099_));
 sg13g2_a21oi_1 _09503_ (.A1(net326),
    .A2(net304),
    .Y(_04100_),
    .B1(_03262_));
 sg13g2_o21ai_1 _09504_ (.B1(_03889_),
    .Y(_04101_),
    .A1(_02300_),
    .A2(_04100_));
 sg13g2_o21ai_1 _09505_ (.B1(_04101_),
    .Y(_04102_),
    .A1(net341),
    .A2(_04099_));
 sg13g2_nor2_1 _09506_ (.A(_01940_),
    .B(net286),
    .Y(_04103_));
 sg13g2_a221oi_1 _09507_ (.B2(_04103_),
    .C1(net291),
    .B1(_03005_),
    .A1(net248),
    .Y(_04104_),
    .A2(_02414_));
 sg13g2_a21oi_1 _09508_ (.A1(net300),
    .A2(_02453_),
    .Y(_04105_),
    .B1(_04104_));
 sg13g2_nor2_1 _09509_ (.A(net301),
    .B(_04105_),
    .Y(_04106_));
 sg13g2_or4_1 _09510_ (.A(net474),
    .B(net460),
    .C(_04102_),
    .D(_04106_),
    .X(_04107_));
 sg13g2_o21ai_1 _09511_ (.B1(_04107_),
    .Y(_04108_),
    .A1(net375),
    .A2(_04096_));
 sg13g2_a22oi_1 _09512_ (.Y(_04109_),
    .B1(_04108_),
    .B2(_03562_),
    .A2(_04084_),
    .A1(_02606_));
 sg13g2_o21ai_1 _09513_ (.B1(net302),
    .Y(_04110_),
    .A1(net235),
    .A2(_03175_));
 sg13g2_a221oi_1 _09514_ (.B2(_02454_),
    .C1(_04110_),
    .B1(_03434_),
    .A1(net165),
    .Y(_04111_),
    .A2(_02518_));
 sg13g2_nand2_1 _09515_ (.Y(_04112_),
    .A(net311),
    .B(_03434_));
 sg13g2_a21oi_1 _09516_ (.A1(_02945_),
    .A2(_04112_),
    .Y(_04113_),
    .B1(net194));
 sg13g2_a21oi_1 _09517_ (.A1(net241),
    .A2(net167),
    .Y(_04114_),
    .B1(net419));
 sg13g2_nor3_1 _09518_ (.A(net186),
    .B(_04113_),
    .C(_04114_),
    .Y(_04115_));
 sg13g2_nor3_1 _09519_ (.A(net185),
    .B(_04111_),
    .C(_04115_),
    .Y(_04116_));
 sg13g2_nand2_1 _09520_ (.Y(_04117_),
    .A(_02756_),
    .B(net463));
 sg13g2_nand2_1 _09521_ (.Y(_04118_),
    .A(_02809_),
    .B(_03214_));
 sg13g2_a22oi_1 _09522_ (.Y(_04119_),
    .B1(_04118_),
    .B2(_02334_),
    .A2(_04117_),
    .A1(net321));
 sg13g2_nor3_1 _09523_ (.A(net294),
    .B(net193),
    .C(net376),
    .Y(_04120_));
 sg13g2_or4_1 _09524_ (.A(_02791_),
    .B(_02991_),
    .C(_04119_),
    .D(_04120_),
    .X(_04121_));
 sg13g2_a21oi_1 _09525_ (.A1(net254),
    .A2(net310),
    .Y(_04122_),
    .B1(_02467_));
 sg13g2_a21oi_1 _09526_ (.A1(_03285_),
    .A2(_04117_),
    .Y(_04123_),
    .B1(net326));
 sg13g2_nor2_1 _09527_ (.A(_02757_),
    .B(_04123_),
    .Y(_04124_));
 sg13g2_o21ai_1 _09528_ (.B1(_04124_),
    .Y(_04125_),
    .A1(net250),
    .A2(_04122_));
 sg13g2_nand2_1 _09529_ (.Y(_04126_),
    .A(_01935_),
    .B(_02607_));
 sg13g2_nor2_1 _09530_ (.A(net390),
    .B(_02618_),
    .Y(_04127_));
 sg13g2_a21oi_1 _09531_ (.A1(net326),
    .A2(_02908_),
    .Y(_04128_),
    .B1(_04127_));
 sg13g2_nor2_1 _09532_ (.A(net177),
    .B(_04128_),
    .Y(_04129_));
 sg13g2_o21ai_1 _09533_ (.B1(_02823_),
    .Y(_04130_),
    .A1(_04126_),
    .A2(_04129_));
 sg13g2_a221oi_1 _09534_ (.B2(net215),
    .C1(_04130_),
    .B1(_04125_),
    .A1(net301),
    .Y(_04131_),
    .A2(_04121_));
 sg13g2_o21ai_1 _09535_ (.B1(_02779_),
    .Y(_04132_),
    .A1(_04116_),
    .A2(_04131_));
 sg13g2_nand2_1 _09536_ (.Y(_04133_),
    .A(_02684_),
    .B(_02864_));
 sg13g2_o21ai_1 _09537_ (.B1(net309),
    .Y(_04134_),
    .A1(net184),
    .A2(_04133_));
 sg13g2_nand3_1 _09538_ (.B(net330),
    .C(_03149_),
    .A(_01959_),
    .Y(_04135_));
 sg13g2_o21ai_1 _09539_ (.B1(_04135_),
    .Y(_04136_),
    .A1(net388),
    .A2(_02612_));
 sg13g2_a22oi_1 _09540_ (.Y(_04137_),
    .B1(_04136_),
    .B2(net203),
    .A2(_04134_),
    .A1(net285));
 sg13g2_o21ai_1 _09541_ (.B1(net385),
    .Y(_04138_),
    .A1(net329),
    .A2(_03741_));
 sg13g2_nand4_1 _09542_ (.B(net233),
    .C(_03464_),
    .A(net184),
    .Y(_04139_),
    .D(_04138_));
 sg13g2_a21oi_1 _09543_ (.A1(net101),
    .A2(_03080_),
    .Y(_04140_),
    .B1(net325));
 sg13g2_o21ai_1 _09544_ (.B1(net101),
    .Y(_04141_),
    .A1(_02570_),
    .A2(_03795_));
 sg13g2_a21oi_1 _09545_ (.A1(_02712_),
    .A2(_02511_),
    .Y(_04142_),
    .B1(net341));
 sg13g2_a221oi_1 _09546_ (.B2(_04142_),
    .C1(_02432_),
    .B1(_04141_),
    .A1(_04139_),
    .Y(_04143_),
    .A2(_04140_));
 sg13g2_a22oi_1 _09547_ (.Y(_04144_),
    .B1(_02908_),
    .B2(_02864_),
    .A2(net233),
    .A1(net193));
 sg13g2_o21ai_1 _09548_ (.B1(_03414_),
    .Y(_04145_),
    .A1(net241),
    .A2(_04144_));
 sg13g2_nand2_1 _09549_ (.Y(_04146_),
    .A(net285),
    .B(_04145_));
 sg13g2_a22oi_1 _09550_ (.Y(_04147_),
    .B1(_04143_),
    .B2(_04146_),
    .A2(_04137_),
    .A1(_03423_));
 sg13g2_or2_1 _09551_ (.X(_04148_),
    .B(_04147_),
    .A(_02887_));
 sg13g2_a21oi_1 _09552_ (.A1(_02630_),
    .A2(net299),
    .Y(_04149_),
    .B1(net99));
 sg13g2_o21ai_1 _09553_ (.B1(net285),
    .Y(_04150_),
    .A1(_03336_),
    .A2(_04149_));
 sg13g2_nand2_1 _09554_ (.Y(_04151_),
    .A(_03379_),
    .B(_04150_));
 sg13g2_o21ai_1 _09555_ (.B1(_03575_),
    .Y(_04152_),
    .A1(_02963_),
    .A2(_03568_));
 sg13g2_nand3_1 _09556_ (.B(_02830_),
    .C(_04152_),
    .A(_03573_),
    .Y(_04153_));
 sg13g2_a21o_1 _09557_ (.A2(_04153_),
    .A1(_04151_),
    .B1(_02664_),
    .X(_04154_));
 sg13g2_and4_1 _09558_ (.A(_02919_),
    .B(_04132_),
    .C(_04148_),
    .D(_04154_),
    .X(_04155_));
 sg13g2_o21ai_1 _09559_ (.B1(_02847_),
    .Y(_04156_),
    .A1(net289),
    .A2(net197));
 sg13g2_o21ai_1 _09560_ (.B1(_02791_),
    .Y(_04157_),
    .A1(net200),
    .A2(net373));
 sg13g2_a22oi_1 _09561_ (.Y(_04158_),
    .B1(_04157_),
    .B2(net216),
    .A2(_04156_),
    .A1(net305));
 sg13g2_inv_1 _09562_ (.Y(_04159_),
    .A(_04158_));
 sg13g2_nor2_1 _09563_ (.A(net280),
    .B(_04067_),
    .Y(_04160_));
 sg13g2_a22oi_1 _09564_ (.Y(_04161_),
    .B1(_03969_),
    .B2(_04160_),
    .A2(_04159_),
    .A1(net237));
 sg13g2_nor2_1 _09565_ (.A(net335),
    .B(_02877_),
    .Y(_04162_));
 sg13g2_a21oi_1 _09566_ (.A1(net310),
    .A2(_01949_),
    .Y(_04163_),
    .B1(_04162_));
 sg13g2_mux2_1 _09567_ (.A0(_03480_),
    .A1(_04163_),
    .S(net282),
    .X(_04164_));
 sg13g2_nand2_1 _09568_ (.Y(_04165_),
    .A(_02299_),
    .B(net251));
 sg13g2_o21ai_1 _09569_ (.B1(_04165_),
    .Y(_04166_),
    .A1(_02816_),
    .A2(_03156_));
 sg13g2_a221oi_1 _09570_ (.B2(_03230_),
    .C1(_01961_),
    .B1(_04166_),
    .A1(_02544_),
    .Y(_04167_),
    .A2(_03708_));
 sg13g2_a21oi_1 _09571_ (.A1(_03392_),
    .A2(_04164_),
    .Y(_04168_),
    .B1(_04167_));
 sg13g2_nand2_1 _09572_ (.Y(_04169_),
    .A(net181),
    .B(_04168_));
 sg13g2_o21ai_1 _09573_ (.B1(_04169_),
    .Y(_04170_),
    .A1(net134),
    .A2(_04161_));
 sg13g2_o21ai_1 _09574_ (.B1(_02375_),
    .Y(_04171_),
    .A1(_03115_),
    .A2(_03151_));
 sg13g2_a22oi_1 _09575_ (.Y(_04172_),
    .B1(_03175_),
    .B2(_03276_),
    .A2(_02896_),
    .A1(net222));
 sg13g2_nand2_1 _09576_ (.Y(_04173_),
    .A(_02621_),
    .B(_02896_));
 sg13g2_o21ai_1 _09577_ (.B1(_04173_),
    .Y(_04174_),
    .A1(_02400_),
    .A2(_04172_));
 sg13g2_a221oi_1 _09578_ (.B2(_03980_),
    .C1(_03879_),
    .B1(_03882_),
    .A1(_02903_),
    .Y(_04175_),
    .A2(_04174_));
 sg13g2_a21oi_1 _09579_ (.A1(_02820_),
    .A2(_04171_),
    .Y(_04176_),
    .B1(_04175_));
 sg13g2_nor2_1 _09580_ (.A(_02763_),
    .B(_02472_),
    .Y(_04177_));
 sg13g2_a21oi_1 _09581_ (.A1(_02353_),
    .A2(_02536_),
    .Y(_04178_),
    .B1(_04177_));
 sg13g2_inv_1 _09582_ (.Y(_04179_),
    .A(_02954_));
 sg13g2_a21oi_1 _09583_ (.A1(_04179_),
    .A2(_03870_),
    .Y(_04180_),
    .B1(net185));
 sg13g2_o21ai_1 _09584_ (.B1(_04180_),
    .Y(_04181_),
    .A1(_02527_),
    .A2(_04178_));
 sg13g2_o21ai_1 _09585_ (.B1(_04181_),
    .Y(_04182_),
    .A1(net198),
    .A2(_04176_));
 sg13g2_a22oi_1 _09586_ (.Y(_04183_),
    .B1(_04182_),
    .B2(_02828_),
    .A2(_04170_),
    .A1(_02883_));
 sg13g2_and4_1 _09587_ (.A(_04072_),
    .B(_04109_),
    .C(_04155_),
    .D(_04183_),
    .X(_04184_));
 sg13g2_nor2_1 _09588_ (.A(_02725_),
    .B(_04015_),
    .Y(_04185_));
 sg13g2_o21ai_1 _09589_ (.B1(net152),
    .Y(_04186_),
    .A1(_02675_),
    .A2(_04185_));
 sg13g2_o21ai_1 _09590_ (.B1(_04186_),
    .Y(_04187_),
    .A1(net151),
    .A2(_03346_));
 sg13g2_o21ai_1 _09591_ (.B1(net205),
    .Y(_04188_),
    .A1(net154),
    .A2(_03397_));
 sg13g2_o21ai_1 _09592_ (.B1(_03363_),
    .Y(_04189_),
    .A1(_02819_),
    .A2(_04188_));
 sg13g2_nor2_1 _09593_ (.A(net117),
    .B(_04189_),
    .Y(_04190_));
 sg13g2_a21oi_1 _09594_ (.A1(net140),
    .A2(_04187_),
    .Y(_04191_),
    .B1(_04190_));
 sg13g2_o21ai_1 _09595_ (.B1(net316),
    .Y(_04192_),
    .A1(net424),
    .A2(_04191_));
 sg13g2_o21ai_1 _09596_ (.B1(net87),
    .Y(_04193_),
    .A1(_02965_),
    .A2(_03361_));
 sg13g2_and2_1 _09597_ (.A(net80),
    .B(_03816_),
    .X(_04194_));
 sg13g2_a21oi_1 _09598_ (.A1(net123),
    .A2(_04194_),
    .Y(_04195_),
    .B1(net122));
 sg13g2_a21oi_1 _09599_ (.A1(_04193_),
    .A2(_04195_),
    .Y(_04196_),
    .B1(_02953_));
 sg13g2_a21oi_1 _09600_ (.A1(_04192_),
    .A2(_04196_),
    .Y(_04197_),
    .B1(_02920_));
 sg13g2_or3_1 _09601_ (.A(net469),
    .B(_04184_),
    .C(_04197_),
    .X(_04198_));
 sg13g2_o21ai_1 _09602_ (.B1(_04198_),
    .Y(_04199_),
    .A1(_03997_),
    .A2(_04004_));
 sg13g2_nor3_1 _09603_ (.A(net169),
    .B(net79),
    .C(_04085_),
    .Y(_04200_));
 sg13g2_nor2_1 _09604_ (.A(_02627_),
    .B(net374),
    .Y(_04201_));
 sg13g2_nand2b_1 _09605_ (.Y(_04202_),
    .B(net331),
    .A_N(_02347_));
 sg13g2_o21ai_1 _09606_ (.B1(_03014_),
    .Y(_04203_),
    .A1(_01955_),
    .A2(_04202_));
 sg13g2_nand2b_1 _09607_ (.Y(_04204_),
    .B(_02348_),
    .A_N(net331));
 sg13g2_a21oi_1 _09608_ (.A1(_02460_),
    .A2(_04204_),
    .Y(_04205_),
    .B1(_02688_));
 sg13g2_a221oi_1 _09609_ (.B2(_02351_),
    .C1(_04205_),
    .B1(_04203_),
    .A1(net222),
    .Y(_04206_),
    .A2(_04201_));
 sg13g2_o21ai_1 _09610_ (.B1(_03676_),
    .Y(_04207_),
    .A1(net207),
    .A2(_04206_));
 sg13g2_mux2_1 _09611_ (.A0(_04200_),
    .A1(_04207_),
    .S(net236),
    .X(_04208_));
 sg13g2_nor2_1 _09612_ (.A(_02378_),
    .B(_03233_),
    .Y(_04209_));
 sg13g2_a221oi_1 _09613_ (.B2(_02619_),
    .C1(net104),
    .B1(_04209_),
    .A1(net77),
    .Y(_04210_),
    .A2(net106));
 sg13g2_nor3_1 _09614_ (.A(net247),
    .B(net126),
    .C(_04210_),
    .Y(_04211_));
 sg13g2_a21oi_1 _09615_ (.A1(net172),
    .A2(_04208_),
    .Y(_04212_),
    .B1(_04211_));
 sg13g2_a21oi_1 _09616_ (.A1(net212),
    .A2(_03967_),
    .Y(_04213_),
    .B1(net254));
 sg13g2_o21ai_1 _09617_ (.B1(net312),
    .Y(_04214_),
    .A1(net329),
    .A2(net284));
 sg13g2_nand2_1 _09618_ (.Y(_04215_),
    .A(_02304_),
    .B(_04214_));
 sg13g2_o21ai_1 _09619_ (.B1(net305),
    .Y(_04216_),
    .A1(_04213_),
    .A2(_04215_));
 sg13g2_nand3_1 _09620_ (.B(net171),
    .C(net231),
    .A(net113),
    .Y(_04217_));
 sg13g2_o21ai_1 _09621_ (.B1(_03353_),
    .Y(_04218_),
    .A1(_03086_),
    .A2(_03077_));
 sg13g2_nand4_1 _09622_ (.B(_04216_),
    .C(_04217_),
    .A(net280),
    .Y(_04219_),
    .D(_04218_));
 sg13g2_nor2_1 _09623_ (.A(_02520_),
    .B(_02613_),
    .Y(_04220_));
 sg13g2_o21ai_1 _09624_ (.B1(_02386_),
    .Y(_04221_),
    .A1(net294),
    .A2(_04202_));
 sg13g2_nor2_1 _09625_ (.A(net281),
    .B(_03795_),
    .Y(_04222_));
 sg13g2_a21oi_1 _09626_ (.A1(_02341_),
    .A2(_04221_),
    .Y(_04223_),
    .B1(_04222_));
 sg13g2_nor2_1 _09627_ (.A(net97),
    .B(_04223_),
    .Y(_04224_));
 sg13g2_o21ai_1 _09628_ (.B1(_03381_),
    .Y(_04225_),
    .A1(_04220_),
    .A2(_04224_));
 sg13g2_a21o_1 _09629_ (.A2(_04225_),
    .A1(_04219_),
    .B1(_02434_),
    .X(_04226_));
 sg13g2_o21ai_1 _09630_ (.B1(_04226_),
    .Y(_04227_),
    .A1(_02705_),
    .A2(_04212_));
 sg13g2_nor2_1 _09631_ (.A(net297),
    .B(net173),
    .Y(_04228_));
 sg13g2_nor2_1 _09632_ (.A(_02446_),
    .B(net95),
    .Y(_04229_));
 sg13g2_a221oi_1 _09633_ (.B2(net299),
    .C1(net322),
    .B1(net309),
    .A1(net297),
    .Y(_04230_),
    .A2(_02368_));
 sg13g2_a221oi_1 _09634_ (.B2(net224),
    .C1(_04230_),
    .B1(_04229_),
    .A1(net232),
    .Y(_04231_),
    .A2(_04228_));
 sg13g2_o21ai_1 _09635_ (.B1(_04231_),
    .Y(_04232_),
    .A1(_02409_),
    .A2(_02967_));
 sg13g2_nand3_1 _09636_ (.B(_01957_),
    .C(_03708_),
    .A(_03250_),
    .Y(_04233_));
 sg13g2_a21oi_1 _09637_ (.A1(net81),
    .A2(_04233_),
    .Y(_04234_),
    .B1(net175));
 sg13g2_o21ai_1 _09638_ (.B1(_02430_),
    .Y(_04235_),
    .A1(_03248_),
    .A2(_04234_));
 sg13g2_a22oi_1 _09639_ (.Y(_04236_),
    .B1(_04235_),
    .B2(net316),
    .A2(_04232_),
    .A1(net109));
 sg13g2_o21ai_1 _09640_ (.B1(net183),
    .Y(_04237_),
    .A1(net222),
    .A2(net223));
 sg13g2_a22oi_1 _09641_ (.Y(_04238_),
    .B1(_04237_),
    .B2(net314),
    .A2(net284),
    .A1(net254));
 sg13g2_nor2b_1 _09642_ (.A(net208),
    .B_N(_01909_),
    .Y(_04239_));
 sg13g2_nand2_1 _09643_ (.Y(_04240_),
    .A(net326),
    .B(_04239_));
 sg13g2_a221oi_1 _09644_ (.B2(net177),
    .C1(net297),
    .B1(_04240_),
    .A1(net165),
    .Y(_04241_),
    .A2(_04239_));
 sg13g2_o21ai_1 _09645_ (.B1(_04241_),
    .Y(_04242_),
    .A1(net250),
    .A2(_04238_));
 sg13g2_a22oi_1 _09646_ (.Y(_04243_),
    .B1(_03757_),
    .B2(net194),
    .A2(_02337_),
    .A1(_03463_));
 sg13g2_nand2b_1 _09647_ (.Y(_04244_),
    .B(_03381_),
    .A_N(_04243_));
 sg13g2_a21oi_1 _09648_ (.A1(_04242_),
    .A2(_04244_),
    .Y(_04245_),
    .B1(net229));
 sg13g2_o21ai_1 _09649_ (.B1(net304),
    .Y(_04246_),
    .A1(_02720_),
    .A2(_02849_));
 sg13g2_a21oi_1 _09650_ (.A1(_02443_),
    .A2(_04246_),
    .Y(_04247_),
    .B1(net302));
 sg13g2_a21oi_1 _09651_ (.A1(net339),
    .A2(_02804_),
    .Y(_04248_),
    .B1(_04247_));
 sg13g2_o21ai_1 _09652_ (.B1(_02633_),
    .Y(_04249_),
    .A1(net235),
    .A2(net110));
 sg13g2_nand3b_1 _09653_ (.B(_04249_),
    .C(_04097_),
    .Y(_04250_),
    .A_N(_02333_));
 sg13g2_a221oi_1 _09654_ (.B2(net298),
    .C1(_03266_),
    .B1(_04250_),
    .A1(net202),
    .Y(_04251_),
    .A2(_04248_));
 sg13g2_o21ai_1 _09655_ (.B1(_02883_),
    .Y(_04252_),
    .A1(_04245_),
    .A2(_04251_));
 sg13g2_nand2_1 _09656_ (.Y(_04253_),
    .A(net179),
    .B(_02734_));
 sg13g2_nor2_1 _09657_ (.A(net329),
    .B(_02863_),
    .Y(_04254_));
 sg13g2_o21ai_1 _09658_ (.B1(net251),
    .Y(_04255_),
    .A1(net225),
    .A2(_04254_));
 sg13g2_a221oi_1 _09659_ (.B2(_02867_),
    .C1(_03651_),
    .B1(_04255_),
    .A1(_03253_),
    .Y(_04256_),
    .A2(_04253_));
 sg13g2_mux2_1 _09660_ (.A0(_02642_),
    .A1(_03077_),
    .S(net251),
    .X(_04257_));
 sg13g2_a21oi_1 _09661_ (.A1(net153),
    .A2(net129),
    .Y(_04258_),
    .B1(net282));
 sg13g2_a21oi_1 _09662_ (.A1(net203),
    .A2(_04257_),
    .Y(_04259_),
    .B1(_04258_));
 sg13g2_o21ai_1 _09663_ (.B1(_01976_),
    .Y(_04260_),
    .A1(_01788_),
    .A2(net286));
 sg13g2_nand3_1 _09664_ (.B(net385),
    .C(_03022_),
    .A(net431),
    .Y(_04261_));
 sg13g2_nand3_1 _09665_ (.B(_04260_),
    .C(_04261_),
    .A(_02799_),
    .Y(_04262_));
 sg13g2_a21oi_1 _09666_ (.A1(_03644_),
    .A2(_03645_),
    .Y(_04263_),
    .B1(_04262_));
 sg13g2_a21oi_1 _09667_ (.A1(net345),
    .A2(net231),
    .Y(_04264_),
    .B1(net184));
 sg13g2_nor2_1 _09668_ (.A(_02727_),
    .B(_04264_),
    .Y(_04265_));
 sg13g2_nand2_1 _09669_ (.Y(_04266_),
    .A(net318),
    .B(_03014_));
 sg13g2_nand3_1 _09670_ (.B(_03401_),
    .C(_04266_),
    .A(_02983_),
    .Y(_04267_));
 sg13g2_a21oi_1 _09671_ (.A1(_04265_),
    .A2(_04267_),
    .Y(_04268_),
    .B1(net459));
 sg13g2_a22oi_1 _09672_ (.Y(_04269_),
    .B1(_04263_),
    .B2(_04268_),
    .A2(_04259_),
    .A1(_04256_));
 sg13g2_o21ai_1 _09673_ (.B1(net247),
    .Y(_04270_),
    .A1(_04256_),
    .A2(_04263_));
 sg13g2_a21o_1 _09674_ (.A2(_04270_),
    .A1(_04269_),
    .B1(_02887_),
    .X(_04271_));
 sg13g2_a21oi_1 _09675_ (.A1(net220),
    .A2(_01978_),
    .Y(_04272_),
    .B1(_02397_));
 sg13g2_a21oi_1 _09676_ (.A1(_01972_),
    .A2(net299),
    .Y(_04273_),
    .B1(_01754_));
 sg13g2_o21ai_1 _09677_ (.B1(_04273_),
    .Y(_04274_),
    .A1(net78),
    .A2(_04272_));
 sg13g2_and2_1 _09678_ (.A(_03617_),
    .B(_04274_),
    .X(_04275_));
 sg13g2_a22oi_1 _09679_ (.Y(_04276_),
    .B1(_03070_),
    .B2(net246),
    .A2(_03501_),
    .A1(net399));
 sg13g2_nand3b_1 _09680_ (.B(_04276_),
    .C(_02799_),
    .Y(_04277_),
    .A_N(_03623_));
 sg13g2_a22oi_1 _09681_ (.Y(_04278_),
    .B1(_03035_),
    .B2(net300),
    .A2(_02892_),
    .A1(net399));
 sg13g2_nor2_1 _09682_ (.A(net96),
    .B(_04278_),
    .Y(_04279_));
 sg13g2_a21oi_1 _09683_ (.A1(net138),
    .A2(net204),
    .Y(_04280_),
    .B1(_03630_));
 sg13g2_nor3_1 _09684_ (.A(_04277_),
    .B(_04279_),
    .C(_04280_),
    .Y(_04281_));
 sg13g2_o21ai_1 _09685_ (.B1(_02604_),
    .Y(_04282_),
    .A1(_04275_),
    .A2(_04281_));
 sg13g2_nand4_1 _09686_ (.B(_04252_),
    .C(_04271_),
    .A(net59),
    .Y(_04283_),
    .D(_04282_));
 sg13g2_a221oi_1 _09687_ (.B2(_03260_),
    .C1(_04283_),
    .B1(_04236_),
    .A1(_02774_),
    .Y(_04284_),
    .A2(_04227_));
 sg13g2_nand2_1 _09688_ (.Y(_04285_),
    .A(net103),
    .B(net145));
 sg13g2_xnor2_1 _09689_ (.Y(_04286_),
    .A(_02285_),
    .B(_03029_));
 sg13g2_nand2_1 _09690_ (.Y(_04287_),
    .A(net197),
    .B(_02858_));
 sg13g2_a21oi_1 _09691_ (.A1(net244),
    .A2(_03741_),
    .Y(_04288_),
    .B1(_04287_));
 sg13g2_nor2_1 _09692_ (.A(net339),
    .B(_04288_),
    .Y(_04289_));
 sg13g2_o21ai_1 _09693_ (.B1(_04289_),
    .Y(_04290_),
    .A1(_04285_),
    .A2(_04286_));
 sg13g2_o21ai_1 _09694_ (.B1(net155),
    .Y(_04291_),
    .A1(_02686_),
    .A2(_02452_));
 sg13g2_nand3_1 _09695_ (.B(_02656_),
    .C(_04291_),
    .A(_03023_),
    .Y(_04292_));
 sg13g2_nand2_1 _09696_ (.Y(_04293_),
    .A(_03028_),
    .B(_02510_));
 sg13g2_nand3_1 _09697_ (.B(_02413_),
    .C(_04293_),
    .A(_02622_),
    .Y(_04294_));
 sg13g2_nand4_1 _09698_ (.B(_04290_),
    .C(_04292_),
    .A(_02795_),
    .Y(_04295_),
    .D(_04294_));
 sg13g2_o21ai_1 _09699_ (.B1(_02845_),
    .Y(_04296_),
    .A1(_02849_),
    .A2(net179));
 sg13g2_a21oi_1 _09700_ (.A1(_02633_),
    .A2(_04296_),
    .Y(_04297_),
    .B1(net186));
 sg13g2_nor2_1 _09701_ (.A(net234),
    .B(net212),
    .Y(_04298_));
 sg13g2_nor3_1 _09702_ (.A(_02689_),
    .B(_02876_),
    .C(_02878_),
    .Y(_04299_));
 sg13g2_nor3_1 _09703_ (.A(net203),
    .B(_04298_),
    .C(_04299_),
    .Y(_04300_));
 sg13g2_nor3_1 _09704_ (.A(net280),
    .B(_04297_),
    .C(_04300_),
    .Y(_04301_));
 sg13g2_nand3_1 _09705_ (.B(net106),
    .C(_02647_),
    .A(net372),
    .Y(_04302_));
 sg13g2_a21oi_1 _09706_ (.A1(net174),
    .A2(_02903_),
    .Y(_04303_),
    .B1(_04302_));
 sg13g2_o21ai_1 _09707_ (.B1(net181),
    .Y(_04304_),
    .A1(_04301_),
    .A2(_04303_));
 sg13g2_a21oi_1 _09708_ (.A1(_04295_),
    .A2(_04304_),
    .Y(_04305_),
    .B1(_03386_));
 sg13g2_xnor2_1 _09709_ (.Y(_04306_),
    .A(net309),
    .B(_01941_));
 sg13g2_nor2_1 _09710_ (.A(_01910_),
    .B(net173),
    .Y(_04307_));
 sg13g2_o21ai_1 _09711_ (.B1(_04307_),
    .Y(_04308_),
    .A1(net135),
    .A2(_04306_));
 sg13g2_mux2_1 _09712_ (.A0(_02417_),
    .A1(_02897_),
    .S(net311),
    .X(_04309_));
 sg13g2_nand2b_1 _09713_ (.Y(_04310_),
    .B(_04309_),
    .A_N(_01771_));
 sg13g2_o21ai_1 _09714_ (.B1(net111),
    .Y(_04311_),
    .A1(_03253_),
    .A2(_02861_));
 sg13g2_a22oi_1 _09715_ (.Y(_04312_),
    .B1(_03991_),
    .B2(net184),
    .A2(_02666_),
    .A1(net289));
 sg13g2_a21oi_1 _09716_ (.A1(net340),
    .A2(net99),
    .Y(_04313_),
    .B1(_02408_));
 sg13g2_o21ai_1 _09717_ (.B1(_04313_),
    .Y(_04314_),
    .A1(net105),
    .A2(_04312_));
 sg13g2_nand4_1 _09718_ (.B(_04310_),
    .C(_04311_),
    .A(_04308_),
    .Y(_04315_),
    .D(_04314_));
 sg13g2_o21ai_1 _09719_ (.B1(net283),
    .Y(_04316_),
    .A1(_02534_),
    .A2(_02422_));
 sg13g2_nand2_1 _09720_ (.Y(_04317_),
    .A(net309),
    .B(_04316_));
 sg13g2_o21ai_1 _09721_ (.B1(_03239_),
    .Y(_04318_),
    .A1(net302),
    .A2(net95));
 sg13g2_a221oi_1 _09722_ (.B2(net171),
    .C1(_04318_),
    .B1(_04317_),
    .A1(net305),
    .Y(_04319_),
    .A2(_02929_));
 sg13g2_xor2_1 _09723_ (.B(net208),
    .A(net392),
    .X(_04320_));
 sg13g2_a22oi_1 _09724_ (.Y(_04321_),
    .B1(_02985_),
    .B2(_04320_),
    .A2(net173),
    .A1(net232));
 sg13g2_o21ai_1 _09725_ (.B1(_02428_),
    .Y(_04322_),
    .A1(_04000_),
    .A2(_04321_));
 sg13g2_nor2_1 _09726_ (.A(_04319_),
    .B(_04322_),
    .Y(_04323_));
 sg13g2_a21oi_1 _09727_ (.A1(_02824_),
    .A2(_04315_),
    .Y(_04324_),
    .B1(_04323_));
 sg13g2_a21oi_1 _09728_ (.A1(net293),
    .A2(_02441_),
    .Y(_04325_),
    .B1(net377));
 sg13g2_a21oi_1 _09729_ (.A1(net323),
    .A2(_04325_),
    .Y(_04326_),
    .B1(net388));
 sg13g2_o21ai_1 _09730_ (.B1(net124),
    .Y(_04327_),
    .A1(_03101_),
    .A2(_04326_));
 sg13g2_a21oi_1 _09731_ (.A1(_02388_),
    .A2(_02851_),
    .Y(_04328_),
    .B1(net294));
 sg13g2_o21ai_1 _09732_ (.B1(net315),
    .Y(_04329_),
    .A1(_02991_),
    .A2(_04328_));
 sg13g2_nor3_1 _09733_ (.A(net388),
    .B(net291),
    .C(_04325_),
    .Y(_04330_));
 sg13g2_a221oi_1 _09734_ (.B2(_04329_),
    .C1(_04330_),
    .B1(_04307_),
    .A1(net218),
    .Y(_04331_),
    .A2(_03101_));
 sg13g2_nand2_1 _09735_ (.Y(_04332_),
    .A(_04327_),
    .B(_04331_));
 sg13g2_a21oi_1 _09736_ (.A1(net309),
    .A2(_03722_),
    .Y(_04333_),
    .B1(net304));
 sg13g2_o21ai_1 _09737_ (.B1(net215),
    .Y(_04334_),
    .A1(net286),
    .A2(_04333_));
 sg13g2_nand2_1 _09738_ (.Y(_04335_),
    .A(net308),
    .B(_03723_));
 sg13g2_nand2_1 _09739_ (.Y(_04336_),
    .A(_03807_),
    .B(_04335_));
 sg13g2_nand3_1 _09740_ (.B(_04334_),
    .C(_04336_),
    .A(_03695_),
    .Y(_04337_));
 sg13g2_nand2b_1 _09741_ (.Y(_04338_),
    .B(_03456_),
    .A_N(_02977_));
 sg13g2_a221oi_1 _09742_ (.B2(_02428_),
    .C1(_04338_),
    .B1(_04337_),
    .A1(net181),
    .Y(_04339_),
    .A2(_04332_));
 sg13g2_a21o_1 _09743_ (.A2(_04324_),
    .A1(_03603_),
    .B1(_04339_),
    .X(_04340_));
 sg13g2_nor2_1 _09744_ (.A(_01789_),
    .B(_02816_),
    .Y(_04341_));
 sg13g2_o21ai_1 _09745_ (.B1(_03744_),
    .Y(_04342_),
    .A1(_04126_),
    .A2(_04341_));
 sg13g2_nand3_1 _09746_ (.B(_03687_),
    .C(_03204_),
    .A(_02725_),
    .Y(_04343_));
 sg13g2_a21oi_1 _09747_ (.A1(_02782_),
    .A2(_03003_),
    .Y(_04344_),
    .B1(_02365_));
 sg13g2_a221oi_1 _09748_ (.B2(_04344_),
    .C1(net424),
    .B1(_04343_),
    .A1(net280),
    .Y(_04345_),
    .A2(_04342_));
 sg13g2_nor2_1 _09749_ (.A(_02660_),
    .B(_04345_),
    .Y(_04346_));
 sg13g2_a21o_1 _09750_ (.A2(net102),
    .A1(net289),
    .B1(_02991_),
    .X(_04347_));
 sg13g2_a221oi_1 _09751_ (.B2(net217),
    .C1(net203),
    .B1(_04347_),
    .A1(net374),
    .Y(_04348_),
    .A2(_02519_));
 sg13g2_a21oi_1 _09752_ (.A1(net422),
    .A2(_03075_),
    .Y(_04349_),
    .B1(_02863_));
 sg13g2_o21ai_1 _09753_ (.B1(net385),
    .Y(_04350_),
    .A1(net328),
    .A2(net283));
 sg13g2_a221oi_1 _09754_ (.B2(net191),
    .C1(net314),
    .B1(_04350_),
    .A1(net200),
    .Y(_04351_),
    .A2(_04349_));
 sg13g2_a21oi_1 _09755_ (.A1(_02682_),
    .A2(_04349_),
    .Y(_04352_),
    .B1(net226));
 sg13g2_nand4_1 _09756_ (.B(net303),
    .C(_02642_),
    .A(net195),
    .Y(_04353_),
    .D(_03077_));
 sg13g2_o21ai_1 _09757_ (.B1(_04353_),
    .Y(_04354_),
    .A1(_04351_),
    .A2(_04352_));
 sg13g2_o21ai_1 _09758_ (.B1(_04354_),
    .Y(_04355_),
    .A1(net202),
    .A2(_04348_));
 sg13g2_a21oi_1 _09759_ (.A1(net191),
    .A2(_03135_),
    .Y(_04356_),
    .B1(_02522_));
 sg13g2_o21ai_1 _09760_ (.B1(_03632_),
    .Y(_04357_),
    .A1(net77),
    .A2(_04356_));
 sg13g2_a21o_1 _09761_ (.A2(_04357_),
    .A1(_03467_),
    .B1(net238),
    .X(_04358_));
 sg13g2_a21oi_1 _09762_ (.A1(_04355_),
    .A2(_04358_),
    .Y(_04359_),
    .B1(net198));
 sg13g2_nor3_1 _09763_ (.A(_03752_),
    .B(_04346_),
    .C(_04359_),
    .Y(_04360_));
 sg13g2_a21oi_1 _09764_ (.A1(net128),
    .A2(net141),
    .Y(_04361_),
    .B1(_03078_));
 sg13g2_a21oi_1 _09765_ (.A1(net174),
    .A2(_02858_),
    .Y(_04362_),
    .B1(net205));
 sg13g2_o21ai_1 _09766_ (.B1(_04362_),
    .Y(_04363_),
    .A1(_03833_),
    .A2(_04361_));
 sg13g2_a21oi_1 _09767_ (.A1(net141),
    .A2(_02719_),
    .Y(_04364_),
    .B1(_03211_));
 sg13g2_a21oi_1 _09768_ (.A1(net81),
    .A2(_04364_),
    .Y(_04365_),
    .B1(net185));
 sg13g2_a21oi_1 _09769_ (.A1(net155),
    .A2(_02708_),
    .Y(_04366_),
    .B1(net295));
 sg13g2_o21ai_1 _09770_ (.B1(_03023_),
    .Y(_04367_),
    .A1(net306),
    .A2(_04366_));
 sg13g2_nand3_1 _09771_ (.B(_04365_),
    .C(_04367_),
    .A(_04363_),
    .Y(_04368_));
 sg13g2_a21oi_1 _09772_ (.A1(net213),
    .A2(_03083_),
    .Y(_04369_),
    .B1(_03066_));
 sg13g2_a21oi_1 _09773_ (.A1(net223),
    .A2(net183),
    .Y(_04370_),
    .B1(_02744_));
 sg13g2_nor3_1 _09774_ (.A(net315),
    .B(_02696_),
    .C(_04370_),
    .Y(_04371_));
 sg13g2_a21o_1 _09775_ (.A2(_04369_),
    .A1(net240),
    .B1(_04371_),
    .X(_04372_));
 sg13g2_nand2b_1 _09776_ (.Y(_04373_),
    .B(_03299_),
    .A_N(_03268_));
 sg13g2_a221oi_1 _09777_ (.B2(_03951_),
    .C1(net247),
    .B1(_04373_),
    .A1(_02651_),
    .Y(_04374_),
    .A2(_04372_));
 sg13g2_a21oi_1 _09778_ (.A1(net345),
    .A2(net190),
    .Y(_04375_),
    .B1(_04302_));
 sg13g2_o21ai_1 _09779_ (.B1(_02916_),
    .Y(_04376_),
    .A1(_04374_),
    .A2(_04375_));
 sg13g2_inv_1 _09780_ (.Y(_04377_),
    .A(_02779_));
 sg13g2_a21oi_1 _09781_ (.A1(_04368_),
    .A2(_04376_),
    .Y(_04378_),
    .B1(_04377_));
 sg13g2_nor4_1 _09782_ (.A(_04305_),
    .B(_04340_),
    .C(_04360_),
    .D(_04378_),
    .Y(_04379_));
 sg13g2_a21oi_1 _09783_ (.A1(_03193_),
    .A2(_03361_),
    .Y(_04380_),
    .B1(_03056_));
 sg13g2_a21o_1 _09784_ (.A2(_03581_),
    .A1(_02714_),
    .B1(net79),
    .X(_04381_));
 sg13g2_a221oi_1 _09785_ (.B2(_04381_),
    .C1(net202),
    .B1(_03229_),
    .A1(net76),
    .Y(_04382_),
    .A2(net106));
 sg13g2_a21o_1 _09786_ (.A2(_04380_),
    .A1(_02681_),
    .B1(_04382_),
    .X(_04383_));
 sg13g2_a21oi_1 _09787_ (.A1(_02555_),
    .A2(_03943_),
    .Y(_04384_),
    .B1(net424));
 sg13g2_o21ai_1 _09788_ (.B1(net246),
    .Y(_04385_),
    .A1(net81),
    .A2(net187));
 sg13g2_o21ai_1 _09789_ (.B1(net228),
    .Y(_04386_),
    .A1(net88),
    .A2(net111));
 sg13g2_o21ai_1 _09790_ (.B1(net188),
    .Y(_04387_),
    .A1(net286),
    .A2(net81));
 sg13g2_nand4_1 _09791_ (.B(_04385_),
    .C(_04386_),
    .A(_04384_),
    .Y(_04388_),
    .D(_04387_));
 sg13g2_a221oi_1 _09792_ (.B2(net316),
    .C1(_03582_),
    .B1(_04388_),
    .A1(net108),
    .Y(_04389_),
    .A2(_04383_));
 sg13g2_nor2_1 _09793_ (.A(_02920_),
    .B(_04389_),
    .Y(_04390_));
 sg13g2_a21o_1 _09794_ (.A2(_04379_),
    .A1(_04284_),
    .B1(_04390_),
    .X(_04391_));
 sg13g2_nand2_1 _09795_ (.Y(_04392_),
    .A(net97),
    .B(net306));
 sg13g2_nor2_1 _09796_ (.A(net116),
    .B(net107),
    .Y(_04393_));
 sg13g2_a221oi_1 _09797_ (.B2(_04393_),
    .C1(_01771_),
    .B1(_04392_),
    .A1(net116),
    .Y(_04394_),
    .A2(_03374_));
 sg13g2_a22oi_1 _09798_ (.Y(_04395_),
    .B1(_02871_),
    .B2(net163),
    .A2(_02761_),
    .A1(net166));
 sg13g2_nand2_1 _09799_ (.Y(_04396_),
    .A(_02471_),
    .B(_02666_));
 sg13g2_a21oi_1 _09800_ (.A1(net143),
    .A2(_04396_),
    .Y(_04397_),
    .B1(net219));
 sg13g2_nor3_1 _09801_ (.A(_01962_),
    .B(_04395_),
    .C(_04397_),
    .Y(_04398_));
 sg13g2_nand4_1 _09802_ (.B(_04396_),
    .C(_03101_),
    .A(net119),
    .Y(_04399_),
    .D(_04014_));
 sg13g2_nand2_1 _09803_ (.Y(_04400_),
    .A(_02402_),
    .B(_02979_));
 sg13g2_nand3_1 _09804_ (.B(_04399_),
    .C(_04400_),
    .A(_03117_),
    .Y(_04401_));
 sg13g2_nor3_1 _09805_ (.A(_04394_),
    .B(_04398_),
    .C(_04401_),
    .Y(_04402_));
 sg13g2_nor2_1 _09806_ (.A(_03037_),
    .B(net189),
    .Y(_04403_));
 sg13g2_a21oi_1 _09807_ (.A1(net373),
    .A2(net321),
    .Y(_04404_),
    .B1(net291));
 sg13g2_o21ai_1 _09808_ (.B1(_02626_),
    .Y(_04405_),
    .A1(_04403_),
    .A2(_04404_));
 sg13g2_nor2_1 _09809_ (.A(_02733_),
    .B(_03159_),
    .Y(_04406_));
 sg13g2_o21ai_1 _09810_ (.B1(_04406_),
    .Y(_04407_),
    .A1(_03115_),
    .A2(_03515_));
 sg13g2_nand3_1 _09811_ (.B(net133),
    .C(net189),
    .A(net305),
    .Y(_04408_));
 sg13g2_nand3_1 _09812_ (.B(_04407_),
    .C(_04408_),
    .A(_04405_),
    .Y(_04409_));
 sg13g2_a221oi_1 _09813_ (.B2(net143),
    .C1(_02811_),
    .B1(_03144_),
    .A1(net164),
    .Y(_04410_),
    .A2(_02612_));
 sg13g2_a22oi_1 _09814_ (.Y(_04411_),
    .B1(_04410_),
    .B2(_03381_),
    .A2(_04409_),
    .A1(net206));
 sg13g2_nor2_1 _09815_ (.A(_02434_),
    .B(_04411_),
    .Y(_04412_));
 sg13g2_o21ai_1 _09816_ (.B1(_02774_),
    .Y(_04413_),
    .A1(_04402_),
    .A2(_04412_));
 sg13g2_nor2_1 _09817_ (.A(net163),
    .B(_02788_),
    .Y(_04414_));
 sg13g2_a22oi_1 _09818_ (.Y(_04415_),
    .B1(_04414_),
    .B2(_02726_),
    .A2(net174),
    .A1(_02693_));
 sg13g2_nor3_1 _09819_ (.A(_03298_),
    .B(_02801_),
    .C(_04415_),
    .Y(_04416_));
 sg13g2_nor3_1 _09820_ (.A(net285),
    .B(_04179_),
    .C(_02868_),
    .Y(_04417_));
 sg13g2_nand2_1 _09821_ (.Y(_04418_),
    .A(_01969_),
    .B(_03076_));
 sg13g2_a21oi_1 _09822_ (.A1(_02533_),
    .A2(_03119_),
    .Y(_04419_),
    .B1(_04418_));
 sg13g2_a221oi_1 _09823_ (.B2(_04417_),
    .C1(_04419_),
    .B1(_03278_),
    .A1(_02403_),
    .Y(_04420_),
    .A2(_02565_));
 sg13g2_nor2_1 _09824_ (.A(net198),
    .B(_04420_),
    .Y(_04421_));
 sg13g2_o21ai_1 _09825_ (.B1(_02779_),
    .Y(_04422_),
    .A1(_04416_),
    .A2(_04421_));
 sg13g2_nor2_1 _09826_ (.A(net165),
    .B(net308),
    .Y(_04423_));
 sg13g2_a21oi_1 _09827_ (.A1(net165),
    .A2(net223),
    .Y(_04424_),
    .B1(_04423_));
 sg13g2_a21oi_1 _09828_ (.A1(net112),
    .A2(_04424_),
    .Y(_04425_),
    .B1(net236));
 sg13g2_nand2_1 _09829_ (.Y(_04426_),
    .A(net236),
    .B(_03467_));
 sg13g2_o21ai_1 _09830_ (.B1(_04426_),
    .Y(_04427_),
    .A1(net202),
    .A2(_04425_));
 sg13g2_o21ai_1 _09831_ (.B1(net324),
    .Y(_04428_),
    .A1(net186),
    .A2(net209));
 sg13g2_a221oi_1 _09832_ (.B2(_03903_),
    .C1(net114),
    .B1(net176),
    .A1(net96),
    .Y(_04429_),
    .A2(net209));
 sg13g2_a21oi_1 _09833_ (.A1(_04428_),
    .A2(_04429_),
    .Y(_04430_),
    .B1(_03651_));
 sg13g2_o21ai_1 _09834_ (.B1(_02707_),
    .Y(_04431_),
    .A1(net295),
    .A2(_02441_));
 sg13g2_nand2_1 _09835_ (.Y(_04432_),
    .A(net345),
    .B(net281));
 sg13g2_a221oi_1 _09836_ (.B2(net184),
    .C1(net95),
    .B1(_04432_),
    .A1(net120),
    .Y(_04433_),
    .A2(_04431_));
 sg13g2_a21oi_1 _09837_ (.A1(_02836_),
    .A2(_04433_),
    .Y(_04434_),
    .B1(net324));
 sg13g2_a21oi_1 _09838_ (.A1(net150),
    .A2(net225),
    .Y(_04435_),
    .B1(_04260_));
 sg13g2_nor4_1 _09839_ (.A(net229),
    .B(_04434_),
    .C(_04435_),
    .D(_04010_),
    .Y(_04436_));
 sg13g2_a21oi_1 _09840_ (.A1(_04427_),
    .A2(_04430_),
    .Y(_04437_),
    .B1(_04436_));
 sg13g2_or2_1 _09841_ (.X(_04438_),
    .B(_04437_),
    .A(_02887_));
 sg13g2_nand3_1 _09842_ (.B(_04422_),
    .C(_04438_),
    .A(_04413_),
    .Y(_04439_));
 sg13g2_o21ai_1 _09843_ (.B1(net186),
    .Y(_04440_),
    .A1(_01901_),
    .A2(_02839_));
 sg13g2_o21ai_1 _09844_ (.B1(_04440_),
    .Y(_04441_),
    .A1(_02526_),
    .A2(_02860_));
 sg13g2_a21o_1 _09845_ (.A2(_03581_),
    .A1(_02562_),
    .B1(_02992_),
    .X(_04442_));
 sg13g2_nor2_1 _09846_ (.A(net203),
    .B(_02868_),
    .Y(_04443_));
 sg13g2_a221oi_1 _09847_ (.B2(_04443_),
    .C1(net202),
    .B1(_04442_),
    .A1(net76),
    .Y(_04444_),
    .A2(net106));
 sg13g2_a21o_1 _09848_ (.A2(_04441_),
    .A1(_02901_),
    .B1(_04444_),
    .X(_04445_));
 sg13g2_nand2_1 _09849_ (.Y(_04446_),
    .A(_02533_),
    .B(net95));
 sg13g2_nand2_1 _09850_ (.Y(_04447_),
    .A(_02955_),
    .B(net79));
 sg13g2_a22oi_1 _09851_ (.Y(_04448_),
    .B1(_04447_),
    .B2(_04228_),
    .A2(_04446_),
    .A1(_02861_));
 sg13g2_nand2_1 _09852_ (.Y(_04449_),
    .A(_04384_),
    .B(_04448_));
 sg13g2_a22oi_1 _09853_ (.Y(_04450_),
    .B1(_04449_),
    .B2(net316),
    .A2(_04445_),
    .A1(net109));
 sg13g2_nor2_1 _09854_ (.A(_02919_),
    .B(_03582_),
    .Y(_04451_));
 sg13g2_mux2_1 _09855_ (.A0(net422),
    .A1(_02892_),
    .S(net391),
    .X(_04452_));
 sg13g2_nand2_1 _09856_ (.Y(_04453_),
    .A(net388),
    .B(_04452_));
 sg13g2_o21ai_1 _09857_ (.B1(_04453_),
    .Y(_04454_),
    .A1(net106),
    .A2(_04042_));
 sg13g2_nand2_1 _09858_ (.Y(_04455_),
    .A(net120),
    .B(net337));
 sg13g2_a22oi_1 _09859_ (.Y(_04456_),
    .B1(_04455_),
    .B2(net287),
    .A2(_02333_),
    .A1(_02554_));
 sg13g2_nand2b_1 _09860_ (.Y(_04457_),
    .B(net104),
    .A_N(_04456_));
 sg13g2_a221oi_1 _09861_ (.B2(net190),
    .C1(net446),
    .B1(_04457_),
    .A1(net104),
    .Y(_04458_),
    .A2(_04454_));
 sg13g2_a21oi_1 _09862_ (.A1(net204),
    .A2(net281),
    .Y(_04459_),
    .B1(net79));
 sg13g2_nor2b_1 _09863_ (.A(_04459_),
    .B_N(_02593_),
    .Y(_04460_));
 sg13g2_o21ai_1 _09864_ (.B1(net421),
    .Y(_04461_),
    .A1(_04458_),
    .A2(_04460_));
 sg13g2_a21oi_1 _09865_ (.A1(net312),
    .A2(_02870_),
    .Y(_04462_),
    .B1(_02908_));
 sg13g2_o21ai_1 _09866_ (.B1(_02417_),
    .Y(_04463_),
    .A1(net177),
    .A2(_04462_));
 sg13g2_a21oi_1 _09867_ (.A1(net103),
    .A2(_04463_),
    .Y(_04464_),
    .B1(_03328_));
 sg13g2_o21ai_1 _09868_ (.B1(net242),
    .Y(_04465_),
    .A1(net105),
    .A2(_03063_));
 sg13g2_a21oi_1 _09869_ (.A1(net105),
    .A2(_03952_),
    .Y(_04466_),
    .B1(_02727_));
 sg13g2_nand3_1 _09870_ (.B(_04465_),
    .C(_04466_),
    .A(net219),
    .Y(_04467_));
 sg13g2_o21ai_1 _09871_ (.B1(_04467_),
    .Y(_04468_),
    .A1(net249),
    .A2(_04464_));
 sg13g2_nand2_1 _09872_ (.Y(_04469_),
    .A(net244),
    .B(net167));
 sg13g2_nand3_1 _09873_ (.B(_02523_),
    .C(_04469_),
    .A(_03326_),
    .Y(_04470_));
 sg13g2_nand2_1 _09874_ (.Y(_04471_),
    .A(_03326_),
    .B(_03897_));
 sg13g2_a21oi_1 _09875_ (.A1(_02890_),
    .A2(net110),
    .Y(_04472_),
    .B1(_01911_));
 sg13g2_a221oi_1 _09876_ (.B2(_04472_),
    .C1(net229),
    .B1(_04471_),
    .A1(net298),
    .Y(_04473_),
    .A2(_04470_));
 sg13g2_o21ai_1 _09877_ (.B1(_04473_),
    .Y(_04474_),
    .A1(net172),
    .A2(_04468_));
 sg13g2_a21oi_1 _09878_ (.A1(_04461_),
    .A2(_04474_),
    .Y(_04475_),
    .B1(_03292_));
 sg13g2_a21o_1 _09879_ (.A2(_04451_),
    .A1(_04450_),
    .B1(_04475_),
    .X(_04476_));
 sg13g2_a21oi_1 _09880_ (.A1(net218),
    .A2(net167),
    .Y(_04477_),
    .B1(_03121_));
 sg13g2_nand2_1 _09881_ (.Y(_04478_),
    .A(net145),
    .B(_03387_));
 sg13g2_o21ai_1 _09882_ (.B1(_04478_),
    .Y(_04479_),
    .A1(net145),
    .A2(_04477_));
 sg13g2_a221oi_1 _09883_ (.B2(net245),
    .C1(net121),
    .B1(_04479_),
    .A1(_01943_),
    .Y(_04480_),
    .A2(net209));
 sg13g2_nand2_1 _09884_ (.Y(_04481_),
    .A(net213),
    .B(_04127_));
 sg13g2_o21ai_1 _09885_ (.B1(net334),
    .Y(_04482_),
    .A1(net373),
    .A2(net130));
 sg13g2_a21oi_1 _09886_ (.A1(_04481_),
    .A2(_04482_),
    .Y(_04483_),
    .B1(_02634_));
 sg13g2_o21ai_1 _09887_ (.B1(net206),
    .Y(_04484_),
    .A1(net118),
    .A2(_04483_));
 sg13g2_nand2_1 _09888_ (.Y(_04485_),
    .A(_04058_),
    .B(net110));
 sg13g2_a21oi_1 _09889_ (.A1(net111),
    .A2(_04485_),
    .Y(_04486_),
    .B1(net136));
 sg13g2_o21ai_1 _09890_ (.B1(_03346_),
    .Y(_04487_),
    .A1(net162),
    .A2(_02614_));
 sg13g2_a221oi_1 _09891_ (.B2(net246),
    .C1(net198),
    .B1(_04487_),
    .A1(_02418_),
    .Y(_04488_),
    .A2(_04486_));
 sg13g2_o21ai_1 _09892_ (.B1(_04488_),
    .Y(_04489_),
    .A1(_04480_),
    .A2(_04484_));
 sg13g2_a21oi_1 _09893_ (.A1(net174),
    .A2(_02750_),
    .Y(_04490_),
    .B1(net128));
 sg13g2_o21ai_1 _09894_ (.B1(net137),
    .Y(_04491_),
    .A1(net373),
    .A2(_03020_));
 sg13g2_o21ai_1 _09895_ (.B1(net60),
    .Y(_04492_),
    .A1(_04490_),
    .A2(_04491_));
 sg13g2_nand2b_1 _09896_ (.Y(_04493_),
    .B(_04492_),
    .A_N(_01984_));
 sg13g2_a21oi_1 _09897_ (.A1(net168),
    .A2(net337),
    .Y(_04494_),
    .B1(net220));
 sg13g2_o21ai_1 _09898_ (.B1(net285),
    .Y(_04495_),
    .A1(_03233_),
    .A2(_04494_));
 sg13g2_a21oi_1 _09899_ (.A1(net309),
    .A2(_03272_),
    .Y(_04496_),
    .B1(_02889_));
 sg13g2_o21ai_1 _09900_ (.B1(_02782_),
    .Y(_04497_),
    .A1(_02992_),
    .A2(_04496_));
 sg13g2_nand2b_1 _09901_ (.Y(_04498_),
    .B(_04497_),
    .A_N(_04495_));
 sg13g2_mux2_1 _09902_ (.A0(_02642_),
    .A1(_04349_),
    .S(net235),
    .X(_04499_));
 sg13g2_nand2_1 _09903_ (.Y(_04500_),
    .A(net194),
    .B(net307));
 sg13g2_o21ai_1 _09904_ (.B1(_04500_),
    .Y(_04501_),
    .A1(net194),
    .A2(_03005_));
 sg13g2_a22oi_1 _09905_ (.Y(_04502_),
    .B1(_04501_),
    .B2(net292),
    .A2(_04499_),
    .A1(net298));
 sg13g2_nand3_1 _09906_ (.B(_04498_),
    .C(_04502_),
    .A(_02430_),
    .Y(_04503_));
 sg13g2_a21oi_1 _09907_ (.A1(net375),
    .A2(_04503_),
    .Y(_04504_),
    .B1(_02596_));
 sg13g2_nand3_1 _09908_ (.B(_04493_),
    .C(_04504_),
    .A(_04489_),
    .Y(_04505_));
 sg13g2_nand2_1 _09909_ (.Y(_04506_),
    .A(_02425_),
    .B(_03066_));
 sg13g2_a221oi_1 _09910_ (.B2(_04506_),
    .C1(net185),
    .B1(_04289_),
    .A1(_01938_),
    .Y(_04507_),
    .A2(_03092_));
 sg13g2_nand2_1 _09911_ (.Y(_04508_),
    .A(net114),
    .B(net433));
 sg13g2_o21ai_1 _09912_ (.B1(_03640_),
    .Y(_04509_),
    .A1(net115),
    .A2(_04508_));
 sg13g2_a22oi_1 _09913_ (.Y(_04510_),
    .B1(_04509_),
    .B2(_03381_),
    .A2(_04417_),
    .A1(net95));
 sg13g2_nor2_1 _09914_ (.A(_02704_),
    .B(_04510_),
    .Y(_04511_));
 sg13g2_o21ai_1 _09915_ (.B1(_02828_),
    .Y(_04512_),
    .A1(_04507_),
    .A2(_04511_));
 sg13g2_a21oi_1 _09916_ (.A1(net214),
    .A2(net304),
    .Y(_04513_),
    .B1(net221));
 sg13g2_nor3_1 _09917_ (.A(net242),
    .B(_03101_),
    .C(_04513_),
    .Y(_04514_));
 sg13g2_nand3_1 _09918_ (.B(net332),
    .C(net243),
    .A(net318),
    .Y(_04515_));
 sg13g2_a21oi_1 _09919_ (.A1(_03101_),
    .A2(_04515_),
    .Y(_04516_),
    .B1(net287));
 sg13g2_nand3_1 _09920_ (.B(net305),
    .C(_03294_),
    .A(net243),
    .Y(_04517_));
 sg13g2_o21ai_1 _09921_ (.B1(net170),
    .Y(_04518_),
    .A1(net422),
    .A2(_03037_));
 sg13g2_a21oi_1 _09922_ (.A1(net303),
    .A2(net284),
    .Y(_04519_),
    .B1(net388));
 sg13g2_nand3_1 _09923_ (.B(_04518_),
    .C(_04519_),
    .A(_04517_),
    .Y(_04520_));
 sg13g2_o21ai_1 _09924_ (.B1(_04520_),
    .Y(_04521_),
    .A1(_04514_),
    .A2(_04516_));
 sg13g2_nand3_1 _09925_ (.B(_03522_),
    .C(_02593_),
    .A(net96),
    .Y(_04522_));
 sg13g2_o21ai_1 _09926_ (.B1(_04522_),
    .Y(_04523_),
    .A1(net401),
    .A2(_04521_));
 sg13g2_o21ai_1 _09927_ (.B1(net345),
    .Y(_04524_),
    .A1(net182),
    .A2(net178));
 sg13g2_o21ai_1 _09928_ (.B1(_04524_),
    .Y(_04525_),
    .A1(net224),
    .A2(net284));
 sg13g2_nand3_1 _09929_ (.B(_02647_),
    .C(net308),
    .A(net96),
    .Y(_04526_));
 sg13g2_a221oi_1 _09930_ (.B2(net215),
    .C1(net229),
    .B1(_04526_),
    .A1(_02759_),
    .Y(_04527_),
    .A2(_04525_));
 sg13g2_o21ai_1 _09931_ (.B1(net124),
    .Y(_04528_),
    .A1(net153),
    .A2(_03077_));
 sg13g2_o21ai_1 _09932_ (.B1(_04528_),
    .Y(_04529_),
    .A1(net138),
    .A2(_03066_));
 sg13g2_nand2_1 _09933_ (.Y(_04530_),
    .A(net114),
    .B(net124));
 sg13g2_nand3_1 _09934_ (.B(net111),
    .C(_04485_),
    .A(net250),
    .Y(_04531_));
 sg13g2_a21oi_1 _09935_ (.A1(_04530_),
    .A2(_04531_),
    .Y(_04532_),
    .B1(net226));
 sg13g2_a21oi_1 _09936_ (.A1(net228),
    .A2(_04529_),
    .Y(_04533_),
    .B1(_04532_));
 sg13g2_a22oi_1 _09937_ (.Y(_04534_),
    .B1(_04527_),
    .B2(_04533_),
    .A2(_04523_),
    .A1(net421));
 sg13g2_nand2b_1 _09938_ (.Y(_04535_),
    .B(_03562_),
    .A_N(_04534_));
 sg13g2_nand3_1 _09939_ (.B(_04512_),
    .C(_04535_),
    .A(_04505_),
    .Y(_04536_));
 sg13g2_nand2_1 _09940_ (.Y(_04537_),
    .A(net301),
    .B(net166));
 sg13g2_o21ai_1 _09941_ (.B1(_02430_),
    .Y(_04538_),
    .A1(net95),
    .A2(_04537_));
 sg13g2_a221oi_1 _09942_ (.B2(net100),
    .C1(_02409_),
    .B1(_03940_),
    .A1(_01889_),
    .Y(_04539_),
    .A2(net76));
 sg13g2_a22oi_1 _09943_ (.Y(_04540_),
    .B1(_02929_),
    .B2(_03505_),
    .A2(_02897_),
    .A1(_02680_));
 sg13g2_nor2_1 _09944_ (.A(net139),
    .B(_04540_),
    .Y(_04541_));
 sg13g2_nor4_1 _09945_ (.A(net421),
    .B(_04538_),
    .C(_04539_),
    .D(_04541_),
    .Y(_04542_));
 sg13g2_nor2_1 _09946_ (.A(net135),
    .B(_01957_),
    .Y(_04543_));
 sg13g2_nor2_1 _09947_ (.A(_03314_),
    .B(_04543_),
    .Y(_04544_));
 sg13g2_xnor2_1 _09948_ (.Y(_04545_),
    .A(_02711_),
    .B(_02629_));
 sg13g2_a221oi_1 _09949_ (.B2(net322),
    .C1(_01961_),
    .B1(_04545_),
    .A1(_02939_),
    .Y(_04546_),
    .A2(_03708_));
 sg13g2_a21oi_1 _09950_ (.A1(net280),
    .A2(_04544_),
    .Y(_04547_),
    .B1(_04546_));
 sg13g2_nand2_1 _09951_ (.Y(_04548_),
    .A(_01913_),
    .B(_04547_));
 sg13g2_nand3_1 _09952_ (.B(net76),
    .C(_02403_),
    .A(net401),
    .Y(_04549_));
 sg13g2_a21oi_1 _09953_ (.A1(_04548_),
    .A2(_04549_),
    .Y(_04550_),
    .B1(_02506_));
 sg13g2_o21ai_1 _09954_ (.B1(_02948_),
    .Y(_04551_),
    .A1(_04542_),
    .A2(_04550_));
 sg13g2_a21oi_1 _09955_ (.A1(net76),
    .A2(net166),
    .Y(_04552_),
    .B1(_02936_));
 sg13g2_a21oi_1 _09956_ (.A1(net115),
    .A2(_03568_),
    .Y(_04553_),
    .B1(_03362_));
 sg13g2_nor2_1 _09957_ (.A(net206),
    .B(_04553_),
    .Y(_04554_));
 sg13g2_nor3_1 _09958_ (.A(net134),
    .B(_04552_),
    .C(_04554_),
    .Y(_04555_));
 sg13g2_a21o_1 _09959_ (.A2(_03410_),
    .A1(net164),
    .B1(net136),
    .X(_04556_));
 sg13g2_a21oi_1 _09960_ (.A1(_04231_),
    .A2(_04556_),
    .Y(_04557_),
    .B1(net401));
 sg13g2_nor2_1 _09961_ (.A(_02506_),
    .B(_04557_),
    .Y(_04558_));
 sg13g2_o21ai_1 _09962_ (.B1(_03260_),
    .Y(_04559_),
    .A1(_04555_),
    .A2(_04558_));
 sg13g2_nand3_1 _09963_ (.B(_02304_),
    .C(_02579_),
    .A(net130),
    .Y(_04560_));
 sg13g2_nand3b_1 _09964_ (.B(_04560_),
    .C(_02435_),
    .Y(_04561_),
    .A_N(_03703_));
 sg13g2_nand3_1 _09965_ (.B(net182),
    .C(_02810_),
    .A(_01789_),
    .Y(_04562_));
 sg13g2_a21oi_1 _09966_ (.A1(net292),
    .A2(_04562_),
    .Y(_04563_),
    .B1(_02703_));
 sg13g2_nand2_1 _09967_ (.Y(_04564_),
    .A(_04561_),
    .B(_04563_));
 sg13g2_o21ai_1 _09968_ (.B1(_02656_),
    .Y(_04565_),
    .A1(_02745_),
    .A2(net113));
 sg13g2_nand3_1 _09969_ (.B(_02945_),
    .C(_04014_),
    .A(net300),
    .Y(_04566_));
 sg13g2_o21ai_1 _09970_ (.B1(_04566_),
    .Y(_04567_),
    .A1(_02792_),
    .A2(_04565_));
 sg13g2_and2_1 _09971_ (.A(net100),
    .B(_04567_),
    .X(_04568_));
 sg13g2_nand2_1 _09972_ (.Y(_04569_),
    .A(_01936_),
    .B(_02510_));
 sg13g2_o21ai_1 _09973_ (.B1(_04569_),
    .Y(_04570_),
    .A1(_02792_),
    .A2(_03156_));
 sg13g2_a221oi_1 _09974_ (.B2(_03298_),
    .C1(_02343_),
    .B1(_04570_),
    .A1(_02706_),
    .Y(_04571_),
    .A2(net129));
 sg13g2_nor3_1 _09975_ (.A(_04564_),
    .B(_04568_),
    .C(_04571_),
    .Y(_04572_));
 sg13g2_nor2_1 _09976_ (.A(net234),
    .B(_03691_),
    .Y(_04573_));
 sg13g2_a221oi_1 _09977_ (.B2(_02656_),
    .C1(_02432_),
    .B1(_04573_),
    .A1(_03718_),
    .Y(_04574_),
    .A2(_03089_));
 sg13g2_nand4_1 _09978_ (.B(net171),
    .C(_04396_),
    .A(net324),
    .Y(_04575_),
    .D(_04014_));
 sg13g2_a22oi_1 _09979_ (.Y(_04576_),
    .B1(_04574_),
    .B2(_04575_),
    .A2(_04563_),
    .A1(_04561_));
 sg13g2_nor2_1 _09980_ (.A(net127),
    .B(net373),
    .Y(_04577_));
 sg13g2_a21oi_1 _09981_ (.A1(net321),
    .A2(_04577_),
    .Y(_04578_),
    .B1(_04220_));
 sg13g2_a21oi_1 _09982_ (.A1(_02634_),
    .A2(_04578_),
    .Y(_04579_),
    .B1(net459));
 sg13g2_nor2_1 _09983_ (.A(net191),
    .B(_04204_),
    .Y(_04580_));
 sg13g2_a21oi_1 _09984_ (.A1(net77),
    .A2(net374),
    .Y(_04581_),
    .B1(_04580_));
 sg13g2_a21oi_1 _09985_ (.A1(net110),
    .A2(_03832_),
    .Y(_04582_),
    .B1(_03299_));
 sg13g2_o21ai_1 _09986_ (.B1(_04582_),
    .Y(_04583_),
    .A1(_02718_),
    .A2(_04581_));
 sg13g2_nand4_1 _09987_ (.B(_04575_),
    .C(_04579_),
    .A(_04574_),
    .Y(_04584_),
    .D(_04583_));
 sg13g2_o21ai_1 _09988_ (.B1(_04584_),
    .Y(_04585_),
    .A1(net123),
    .A2(_04576_));
 sg13g2_o21ai_1 _09989_ (.B1(_02883_),
    .Y(_04586_),
    .A1(_04572_),
    .A2(_04585_));
 sg13g2_nand3_1 _09990_ (.B(_04559_),
    .C(_04586_),
    .A(_04551_),
    .Y(_04587_));
 sg13g2_nor4_1 _09991_ (.A(_04439_),
    .B(_04476_),
    .C(_04536_),
    .D(_04587_),
    .Y(_04588_));
 sg13g2_mux2_1 _09992_ (.A0(_04391_),
    .A1(_04588_),
    .S(_01891_),
    .X(_04589_));
 sg13g2_nand2_1 _09993_ (.Y(_04590_),
    .A(_01892_),
    .B(_04589_));
 sg13g2_o21ai_1 _09994_ (.B1(_04590_),
    .Y(_04591_),
    .A1(_01892_),
    .A2(_04199_));
 sg13g2_nand2_1 _09995_ (.Y(_04592_),
    .A(_01890_),
    .B(_04591_));
 sg13g2_a21oi_1 _09996_ (.A1(_02663_),
    .A2(_02603_),
    .Y(_04593_),
    .B1(_02918_));
 sg13g2_nand3_1 _09997_ (.B(_04592_),
    .C(_04593_),
    .A(_03794_),
    .Y(_04594_));
 sg13g2_buf_1 _09998_ (.A(_04594_),
    .X(_04595_));
 sg13g2_nor2_1 _09999_ (.A(_02331_),
    .B(_04595_),
    .Y(_04596_));
 sg13g2_nor3_1 _10000_ (.A(\draw_game_inst.new_tiles_counter[0] ),
    .B(_01795_),
    .C(_01796_),
    .Y(_04597_));
 sg13g2_mux4_1 _10001_ (.S0(net398),
    .A0(\draw_game_inst.new_tiles[9] ),
    .A1(\draw_game_inst.new_tiles[11] ),
    .A2(\draw_game_inst.new_tiles[10] ),
    .A3(\draw_game_inst.new_tiles[8] ),
    .S1(net397),
    .X(_04598_));
 sg13g2_mux4_1 _10002_ (.S0(net398),
    .A0(\draw_game_inst.new_tiles[1] ),
    .A1(\draw_game_inst.new_tiles[3] ),
    .A2(\draw_game_inst.new_tiles[2] ),
    .A3(\draw_game_inst.new_tiles[0] ),
    .S1(net397),
    .X(_04599_));
 sg13g2_mux4_1 _10003_ (.S0(net398),
    .A0(\draw_game_inst.new_tiles[13] ),
    .A1(\draw_game_inst.new_tiles[15] ),
    .A2(\draw_game_inst.new_tiles[14] ),
    .A3(\draw_game_inst.new_tiles[12] ),
    .S1(net397),
    .X(_04600_));
 sg13g2_mux4_1 _10004_ (.S0(net398),
    .A0(\draw_game_inst.new_tiles[5] ),
    .A1(\draw_game_inst.new_tiles[7] ),
    .A2(\draw_game_inst.new_tiles[6] ),
    .A3(\draw_game_inst.new_tiles[4] ),
    .S1(net397),
    .X(_04601_));
 sg13g2_mux4_1 _10005_ (.S0(net445),
    .A0(_04598_),
    .A1(_04599_),
    .A2(_04600_),
    .A3(_04601_),
    .S1(net475),
    .X(_04602_));
 sg13g2_nand2b_1 _10006_ (.Y(_04603_),
    .B(_04602_),
    .A_N(_04597_));
 sg13g2_nor2_1 _10007_ (.A(_00087_),
    .B(_04603_),
    .Y(_04604_));
 sg13g2_a21oi_1 _10008_ (.A1(net5),
    .A2(_04603_),
    .Y(_04605_),
    .B1(_04604_));
 sg13g2_nand4_1 _10009_ (.B(net346),
    .C(_01914_),
    .A(net6),
    .Y(_04606_),
    .D(_02314_));
 sg13g2_nor3_1 _10010_ (.A(_01774_),
    .B(_01752_),
    .C(_04606_),
    .Y(_04607_));
 sg13g2_and2_1 _10011_ (.A(_02331_),
    .B(_04607_),
    .X(_04608_));
 sg13g2_buf_1 _10012_ (.A(_04608_),
    .X(_04609_));
 sg13g2_inv_1 _10013_ (.Y(_04610_),
    .A(net5));
 sg13g2_inv_1 _10014_ (.Y(_04611_),
    .A(_02331_));
 sg13g2_nor4_1 _10015_ (.A(_01890_),
    .B(net469),
    .C(_01892_),
    .D(net144),
    .Y(_04612_));
 sg13g2_and2_1 _10016_ (.A(net170),
    .B(_04612_),
    .X(_04613_));
 sg13g2_or4_1 _10017_ (.A(_01985_),
    .B(_02305_),
    .C(_02323_),
    .D(_04613_),
    .X(_04614_));
 sg13g2_buf_1 _10018_ (.A(_04614_),
    .X(_04615_));
 sg13g2_and4_1 _10019_ (.A(_04610_),
    .B(_04611_),
    .C(_04595_),
    .D(_04615_),
    .X(_04616_));
 sg13g2_buf_1 _10020_ (.A(_04616_),
    .X(_04617_));
 sg13g2_a221oi_1 _10021_ (.B2(net58),
    .C1(_04617_),
    .B1(_04609_),
    .A1(_04596_),
    .Y(_04618_),
    .A2(_04605_));
 sg13g2_nor2_1 _10022_ (.A(_02317_),
    .B(_04618_),
    .Y(_00171_));
 sg13g2_nand2_1 _10023_ (.Y(_04619_),
    .A(_01795_),
    .B(_04602_));
 sg13g2_a221oi_1 _10024_ (.B2(_04596_),
    .C1(_04617_),
    .B1(_04619_),
    .A1(net126),
    .Y(_04620_),
    .A2(_04609_));
 sg13g2_nor2_1 _10025_ (.A(_02317_),
    .B(_04620_),
    .Y(_00172_));
 sg13g2_nand2_1 _10026_ (.Y(_04621_),
    .A(_01796_),
    .B(_04602_));
 sg13g2_or2_1 _10027_ (.X(_04622_),
    .B(_04621_),
    .A(_04595_));
 sg13g2_nand2_1 _10028_ (.Y(_04623_),
    .A(_04610_),
    .B(_04615_));
 sg13g2_inv_1 _10029_ (.Y(_04624_),
    .A(_04615_));
 sg13g2_nand3_1 _10030_ (.B(net5),
    .C(_04624_),
    .A(net469),
    .Y(_04625_));
 sg13g2_nand3_1 _10031_ (.B(_04623_),
    .C(_04625_),
    .A(_04595_),
    .Y(_04626_));
 sg13g2_nand3_1 _10032_ (.B(_04622_),
    .C(_04626_),
    .A(_04611_),
    .Y(_04627_));
 sg13g2_nand3_1 _10033_ (.B(_02331_),
    .C(_04607_),
    .A(net144),
    .Y(_04628_));
 sg13g2_a21oi_1 _10034_ (.A1(_04627_),
    .A2(_04628_),
    .Y(_00173_),
    .B1(_02317_));
 sg13g2_nor2_1 _10035_ (.A(_02331_),
    .B(_04615_),
    .Y(_04629_));
 sg13g2_nand2_1 _10036_ (.Y(_04630_),
    .A(_01780_),
    .B(_04607_));
 sg13g2_a221oi_1 _10037_ (.B2(_02331_),
    .C1(_02317_),
    .B1(_04630_),
    .A1(_04595_),
    .Y(_00174_),
    .A2(_04629_));
 sg13g2_a21oi_1 _10038_ (.A1(_01777_),
    .A2(_04609_),
    .Y(_04631_),
    .B1(_04617_));
 sg13g2_nor2_1 _10039_ (.A(_02317_),
    .B(_04631_),
    .Y(_00175_));
 sg13g2_nand3_1 _10040_ (.B(_04596_),
    .C(_04603_),
    .A(net5),
    .Y(_04632_));
 sg13g2_a21oi_1 _10041_ (.A1(_01772_),
    .A2(_04609_),
    .Y(_04633_),
    .B1(_04617_));
 sg13g2_a21oi_1 _10042_ (.A1(_04632_),
    .A2(_04633_),
    .Y(_00176_),
    .B1(_02317_));
 sg13g2_buf_1 _10043_ (.A(net407),
    .X(_04634_));
 sg13g2_and2_1 _10044_ (.A(net279),
    .B(net2),
    .X(_00177_));
 sg13g2_and2_1 _10045_ (.A(net279),
    .B(\btn_down_debounce.button_sync_0 ),
    .X(_00178_));
 sg13g2_mux2_1 _10046_ (.A0(\btn_down_debounce.button_sync_1 ),
    .A1(_05073_),
    .S(_02066_),
    .X(_04635_));
 sg13g2_and2_1 _10047_ (.A(net279),
    .B(_04635_),
    .X(_00197_));
 sg13g2_and2_1 _10048_ (.A(_04634_),
    .B(net3),
    .X(_00198_));
 sg13g2_buf_1 _10049_ (.A(net403),
    .X(_04636_));
 sg13g2_and2_1 _10050_ (.A(_04636_),
    .B(\btn_left_debounce.button_sync_0 ),
    .X(_00199_));
 sg13g2_nand2_1 _10051_ (.Y(_04637_),
    .A(\btn_left_debounce.button_sync_1 ),
    .B(_02120_));
 sg13g2_nand2b_1 _10052_ (.Y(_04638_),
    .B(_05066_),
    .A_N(_02120_));
 sg13g2_buf_1 _10053_ (.A(net405),
    .X(_04639_));
 sg13g2_a21oi_1 _10054_ (.A1(_04637_),
    .A2(_04638_),
    .Y(_00218_),
    .B1(net277));
 sg13g2_and2_1 _10055_ (.A(net278),
    .B(net4),
    .X(_00219_));
 sg13g2_and2_1 _10056_ (.A(net278),
    .B(\btn_right_debounce.button_sync_0 ),
    .X(_00220_));
 sg13g2_nand2_1 _10057_ (.Y(_04640_),
    .A(\btn_right_debounce.button_sync_1 ),
    .B(_02177_));
 sg13g2_nand2b_1 _10058_ (.Y(_04641_),
    .B(_05065_),
    .A_N(_02177_));
 sg13g2_a21oi_1 _10059_ (.A1(_04640_),
    .A2(_04641_),
    .Y(_00239_),
    .B1(net277));
 sg13g2_and2_1 _10060_ (.A(net278),
    .B(net1),
    .X(_00240_));
 sg13g2_and2_1 _10061_ (.A(_04636_),
    .B(\btn_up_debounce.button_sync_0 ),
    .X(_00241_));
 sg13g2_nand2_1 _10062_ (.Y(_04642_),
    .A(\btn_up_debounce.button_sync_1 ),
    .B(_02234_));
 sg13g2_nand2b_1 _10063_ (.Y(_04643_),
    .B(_05070_),
    .A_N(_02234_));
 sg13g2_a21oi_1 _10064_ (.A1(_04642_),
    .A2(_04643_),
    .Y(_00260_),
    .B1(net277));
 sg13g2_buf_1 _10065_ (.A(\debug_controller_inst.grid_addr[0] ),
    .X(_04644_));
 sg13g2_buf_1 _10066_ (.A(_04644_),
    .X(_04645_));
 sg13g2_buf_1 _10067_ (.A(\debug_controller_inst.grid_addr[1] ),
    .X(_04646_));
 sg13g2_buf_1 _10068_ (.A(_04646_),
    .X(_04647_));
 sg13g2_mux4_1 _10069_ (.S0(net418),
    .A0(_05215_),
    .A1(_05216_),
    .A2(_05161_),
    .A3(_05160_),
    .S1(net417),
    .X(_04648_));
 sg13g2_mux4_1 _10070_ (.S0(net418),
    .A0(_00468_),
    .A1(_00469_),
    .A2(_05198_),
    .A3(_05197_),
    .S1(net417),
    .X(_04649_));
 sg13g2_buf_2 _10071_ (.A(_04644_),
    .X(_04650_));
 sg13g2_mux4_1 _10072_ (.S0(_04650_),
    .A0(_05222_),
    .A1(_05223_),
    .A2(_05142_),
    .A3(_05141_),
    .S1(net458),
    .X(_04651_));
 sg13g2_mux4_1 _10073_ (.S0(_04650_),
    .A0(_00471_),
    .A1(_00472_),
    .A2(_05208_),
    .A3(_05207_),
    .S1(_04646_),
    .X(_04652_));
 sg13g2_buf_4 _10074_ (.X(_04653_),
    .A(\debug_controller_inst.grid_addr[2] ));
 sg13g2_buf_2 _10075_ (.A(\debug_controller_inst.grid_addr[3] ),
    .X(_04654_));
 sg13g2_mux4_1 _10076_ (.S0(_04653_),
    .A0(_04648_),
    .A1(_04649_),
    .A2(_04651_),
    .A3(_04652_),
    .S1(_04654_),
    .X(_04655_));
 sg13g2_buf_1 _10077_ (.A(uio_in[1]),
    .X(_04656_));
 sg13g2_nand2b_1 _10078_ (.Y(_04657_),
    .B(net6),
    .A_N(net9));
 sg13g2_buf_1 _10079_ (.A(_04657_),
    .X(_04658_));
 sg13g2_nor2_1 _10080_ (.A(net8),
    .B(_04658_),
    .Y(_04659_));
 sg13g2_nand2_1 _10081_ (.Y(_04660_),
    .A(net7),
    .B(_04659_));
 sg13g2_buf_2 _10082_ (.A(_04660_),
    .X(_04661_));
 sg13g2_nor2_1 _10083_ (.A(net481),
    .B(_04661_),
    .Y(_04662_));
 sg13g2_nand2_1 _10084_ (.Y(_04663_),
    .A(_04655_),
    .B(_04662_));
 sg13g2_o21ai_1 _10085_ (.B1(net18),
    .Y(_04664_),
    .A1(_04656_),
    .A2(_04661_));
 sg13g2_a21oi_1 _10086_ (.A1(_04663_),
    .A2(_04664_),
    .Y(_00261_),
    .B1(net277));
 sg13g2_mux4_1 _10087_ (.S0(net418),
    .A0(_05218_),
    .A1(_05219_),
    .A2(_05182_),
    .A3(_05181_),
    .S1(net417),
    .X(_04665_));
 sg13g2_mux4_1 _10088_ (.S0(net418),
    .A0(_05122_),
    .A1(_05123_),
    .A2(_05126_),
    .A3(_05125_),
    .S1(net417),
    .X(_04666_));
 sg13g2_mux4_1 _10089_ (.S0(net416),
    .A0(_05225_),
    .A1(_05226_),
    .A2(_05188_),
    .A3(_05187_),
    .S1(net458),
    .X(_04667_));
 sg13g2_mux4_1 _10090_ (.S0(net416),
    .A0(_05128_),
    .A1(_05129_),
    .A2(_05132_),
    .A3(_05131_),
    .S1(net458),
    .X(_04668_));
 sg13g2_mux4_1 _10091_ (.S0(_04653_),
    .A0(_04665_),
    .A1(_04666_),
    .A2(_04667_),
    .A3(_04668_),
    .S1(_04654_),
    .X(_04669_));
 sg13g2_nand2_1 _10092_ (.Y(_04670_),
    .A(_04662_),
    .B(_04669_));
 sg13g2_o21ai_1 _10093_ (.B1(net19),
    .Y(_04671_),
    .A1(net481),
    .A2(_04661_));
 sg13g2_buf_1 _10094_ (.A(net413),
    .X(_04672_));
 sg13g2_a21oi_1 _10095_ (.A1(_04670_),
    .A2(_04671_),
    .Y(_00262_),
    .B1(net276));
 sg13g2_mux4_1 _10096_ (.S0(net416),
    .A0(_05178_),
    .A1(_05179_),
    .A2(_00460_),
    .A3(_00459_),
    .S1(net417),
    .X(_04673_));
 sg13g2_mux4_1 _10097_ (.S0(net418),
    .A0(_05201_),
    .A1(_05202_),
    .A2(_05195_),
    .A3(_05194_),
    .S1(net417),
    .X(_04674_));
 sg13g2_mux4_1 _10098_ (.S0(net416),
    .A0(_05184_),
    .A1(_05185_),
    .A2(_00463_),
    .A3(_00462_),
    .S1(net458),
    .X(_04675_));
 sg13g2_mux4_1 _10099_ (.S0(net416),
    .A0(_05211_),
    .A1(_05212_),
    .A2(_05205_),
    .A3(_05204_),
    .S1(net458),
    .X(_04676_));
 sg13g2_mux4_1 _10100_ (.S0(_04653_),
    .A0(_04673_),
    .A1(_04674_),
    .A2(_04675_),
    .A3(_04676_),
    .S1(_04654_),
    .X(_04677_));
 sg13g2_nand2_1 _10101_ (.Y(_04678_),
    .A(_04662_),
    .B(_04677_));
 sg13g2_o21ai_1 _10102_ (.B1(net20),
    .Y(_04679_),
    .A1(net481),
    .A2(_04661_));
 sg13g2_a21oi_1 _10103_ (.A1(_04678_),
    .A2(_04679_),
    .Y(_00263_),
    .B1(_04672_));
 sg13g2_mux4_1 _10104_ (.S0(net416),
    .A0(_05149_),
    .A1(_05150_),
    .A2(_05158_),
    .A3(_05157_),
    .S1(net458),
    .X(_04680_));
 sg13g2_mux4_1 _10105_ (.S0(net418),
    .A0(_05165_),
    .A1(_05166_),
    .A2(_05169_),
    .A3(_05168_),
    .S1(net417),
    .X(_04681_));
 sg13g2_mux4_1 _10106_ (.S0(net416),
    .A0(_05152_),
    .A1(_05153_),
    .A2(_05145_),
    .A3(_05144_),
    .S1(net458),
    .X(_04682_));
 sg13g2_mux4_1 _10107_ (.S0(net416),
    .A0(_05171_),
    .A1(_05172_),
    .A2(_05175_),
    .A3(_05174_),
    .S1(net458),
    .X(_04683_));
 sg13g2_mux4_1 _10108_ (.S0(_04653_),
    .A0(_04680_),
    .A1(_04681_),
    .A2(_04682_),
    .A3(_04683_),
    .S1(_04654_),
    .X(_04684_));
 sg13g2_nand2_1 _10109_ (.Y(_04685_),
    .A(_04662_),
    .B(_04684_));
 sg13g2_o21ai_1 _10110_ (.B1(net21),
    .Y(_04686_),
    .A1(net481),
    .A2(_04661_));
 sg13g2_a21oi_1 _10111_ (.A1(_04685_),
    .A2(_04686_),
    .Y(_00264_),
    .B1(_04672_));
 sg13g2_nor3_1 _10112_ (.A(net481),
    .B(net344),
    .C(_04661_),
    .Y(_00265_));
 sg13g2_nor2_1 _10113_ (.A(net7),
    .B(net481),
    .Y(_04687_));
 sg13g2_nand3_1 _10114_ (.B(net447),
    .C(_04687_),
    .A(net8),
    .Y(_04688_));
 sg13g2_nor2_1 _10115_ (.A(_04658_),
    .B(_04688_),
    .Y(_04689_));
 sg13g2_and2_1 _10116_ (.A(net10),
    .B(_04689_),
    .X(_00266_));
 sg13g2_and2_1 _10117_ (.A(net11),
    .B(_04689_),
    .X(_00267_));
 sg13g2_and2_1 _10118_ (.A(net12),
    .B(_04689_),
    .X(_00268_));
 sg13g2_and2_1 _10119_ (.A(net13),
    .B(_04689_),
    .X(_00269_));
 sg13g2_nor3_1 _10120_ (.A(net8),
    .B(_04658_),
    .C(_04687_),
    .Y(_04690_));
 sg13g2_buf_2 _10121_ (.A(_04690_),
    .X(_04691_));
 sg13g2_inv_1 _10122_ (.Y(_04692_),
    .A(net481));
 sg13g2_nor2_1 _10123_ (.A(_04692_),
    .B(_04661_),
    .Y(_04693_));
 sg13g2_buf_2 _10124_ (.A(_04693_),
    .X(_04694_));
 sg13g2_nand2_1 _10125_ (.Y(_04695_),
    .A(net10),
    .B(_04694_));
 sg13g2_nand3_1 _10126_ (.B(net481),
    .C(_04659_),
    .A(net7),
    .Y(_04696_));
 sg13g2_nand2_1 _10127_ (.Y(_04697_),
    .A(_00088_),
    .B(_04696_));
 sg13g2_nand3_1 _10128_ (.B(_04695_),
    .C(_04697_),
    .A(_04691_),
    .Y(_04698_));
 sg13g2_o21ai_1 _10129_ (.B1(_04698_),
    .Y(_04699_),
    .A1(net418),
    .A2(_04691_));
 sg13g2_nor2_1 _10130_ (.A(net361),
    .B(_04699_),
    .Y(_00270_));
 sg13g2_nand2b_1 _10131_ (.Y(_04700_),
    .B(net418),
    .A_N(net417));
 sg13g2_nand2_1 _10132_ (.Y(_04701_),
    .A(net11),
    .B(_04694_));
 sg13g2_o21ai_1 _10133_ (.B1(_04701_),
    .Y(_04702_),
    .A1(_04694_),
    .A2(_04700_));
 sg13g2_o21ai_1 _10134_ (.B1(_04691_),
    .Y(_04703_),
    .A1(_04645_),
    .A2(_04694_));
 sg13g2_a22oi_1 _10135_ (.Y(_04704_),
    .B1(_04703_),
    .B2(_04647_),
    .A2(_04702_),
    .A1(_04691_));
 sg13g2_nor2_1 _10136_ (.A(net361),
    .B(_04704_),
    .Y(_00271_));
 sg13g2_and2_1 _10137_ (.A(\debug_controller_inst.grid_addr[1] ),
    .B(_04644_),
    .X(_04705_));
 sg13g2_buf_1 _10138_ (.A(_04705_),
    .X(_04706_));
 sg13g2_nor2b_1 _10139_ (.A(_04653_),
    .B_N(_04706_),
    .Y(_04707_));
 sg13g2_mux2_1 _10140_ (.A0(net12),
    .A1(_04707_),
    .S(_04696_),
    .X(_04708_));
 sg13g2_o21ai_1 _10141_ (.B1(_04691_),
    .Y(_04709_),
    .A1(_04694_),
    .A2(_04706_));
 sg13g2_a22oi_1 _10142_ (.Y(_04710_),
    .B1(_04709_),
    .B2(_04653_),
    .A2(_04708_),
    .A1(_04691_));
 sg13g2_nor2_1 _10143_ (.A(net277),
    .B(_04710_),
    .Y(_00272_));
 sg13g2_nand2_1 _10144_ (.Y(_04711_),
    .A(_04653_),
    .B(_04706_));
 sg13g2_nor3_1 _10145_ (.A(_04654_),
    .B(_04694_),
    .C(_04711_),
    .Y(_04712_));
 sg13g2_a21o_1 _10146_ (.A2(_04694_),
    .A1(net13),
    .B1(_04712_),
    .X(_04713_));
 sg13g2_nand2_1 _10147_ (.Y(_04714_),
    .A(_04696_),
    .B(_04711_));
 sg13g2_nand2_1 _10148_ (.Y(_04715_),
    .A(_04691_),
    .B(_04714_));
 sg13g2_a22oi_1 _10149_ (.Y(_04716_),
    .B1(_04715_),
    .B2(_04654_),
    .A2(_04713_),
    .A1(_04691_));
 sg13g2_nor2_1 _10150_ (.A(net277),
    .B(_04716_),
    .Y(_00273_));
 sg13g2_nor4_1 _10151_ (.A(net7),
    .B(_04692_),
    .C(net8),
    .D(_04658_),
    .Y(_04717_));
 sg13g2_buf_1 _10152_ (.A(_04717_),
    .X(_04718_));
 sg13g2_buf_1 _10153_ (.A(_04718_),
    .X(_04719_));
 sg13g2_nand2_1 _10154_ (.Y(_04720_),
    .A(_04645_),
    .B(net275));
 sg13g2_nand2b_1 _10155_ (.Y(_04721_),
    .B(net450),
    .A_N(net275));
 sg13g2_a21oi_1 _10156_ (.A1(_04720_),
    .A2(_04721_),
    .Y(_00274_),
    .B1(net276));
 sg13g2_nand2_1 _10157_ (.Y(_04722_),
    .A(_04647_),
    .B(net275));
 sg13g2_nand2b_1 _10158_ (.Y(_04723_),
    .B(_05094_),
    .A_N(_04718_));
 sg13g2_a21oi_1 _10159_ (.A1(_04722_),
    .A2(_04723_),
    .Y(_00275_),
    .B1(net276));
 sg13g2_nand2_1 _10160_ (.Y(_04724_),
    .A(_04653_),
    .B(_04719_));
 sg13g2_nand2b_1 _10161_ (.Y(_04725_),
    .B(_05093_),
    .A_N(_04718_));
 sg13g2_a21oi_1 _10162_ (.A1(_04724_),
    .A2(_04725_),
    .Y(_00276_),
    .B1(net276));
 sg13g2_nand2_1 _10163_ (.Y(_04726_),
    .A(_04654_),
    .B(_04719_));
 sg13g2_nand2b_1 _10164_ (.Y(_04727_),
    .B(_05091_),
    .A_N(_04718_));
 sg13g2_a21oi_1 _10165_ (.A1(_04726_),
    .A2(_04727_),
    .Y(_00277_),
    .B1(net276));
 sg13g2_nand2_1 _10166_ (.Y(_04728_),
    .A(net10),
    .B(net275));
 sg13g2_nand2b_1 _10167_ (.Y(_04729_),
    .B(_00895_),
    .A_N(_04718_));
 sg13g2_a21oi_1 _10168_ (.A1(_04728_),
    .A2(_04729_),
    .Y(_00278_),
    .B1(net276));
 sg13g2_nand2_1 _10169_ (.Y(_04730_),
    .A(net11),
    .B(net275));
 sg13g2_nand2b_1 _10170_ (.Y(_04731_),
    .B(_00921_),
    .A_N(_04718_));
 sg13g2_a21oi_1 _10171_ (.A1(_04730_),
    .A2(_04731_),
    .Y(_00279_),
    .B1(net276));
 sg13g2_nand2_1 _10172_ (.Y(_04732_),
    .A(net12),
    .B(net275));
 sg13g2_nand2b_1 _10173_ (.Y(_04733_),
    .B(net477),
    .A_N(_04718_));
 sg13g2_a21oi_1 _10174_ (.A1(_04732_),
    .A2(_04733_),
    .Y(_00280_),
    .B1(net276));
 sg13g2_nand2_1 _10175_ (.Y(_04734_),
    .A(net13),
    .B(net275));
 sg13g2_nand2b_1 _10176_ (.Y(_04735_),
    .B(net476),
    .A_N(_04718_));
 sg13g2_buf_1 _10177_ (.A(net405),
    .X(_04736_));
 sg13g2_a21oi_1 _10178_ (.A1(_04734_),
    .A2(_04735_),
    .Y(_00281_),
    .B1(_04736_));
 sg13g2_and2_1 _10179_ (.A(net278),
    .B(net275),
    .X(_00282_));
 sg13g2_xor2_1 _10180_ (.B(_01175_),
    .A(_00512_),
    .X(_04737_));
 sg13g2_nand3_1 _10181_ (.B(_00512_),
    .C(_01169_),
    .A(net69),
    .Y(_04738_));
 sg13g2_o21ai_1 _10182_ (.B1(_04738_),
    .Y(_04739_),
    .A1(net69),
    .A2(_04737_));
 sg13g2_nor2_1 _10183_ (.A(_01128_),
    .B(_01164_),
    .Y(_04740_));
 sg13g2_a21oi_1 _10184_ (.A1(_01167_),
    .A2(_01128_),
    .Y(_04741_),
    .B1(_04740_));
 sg13g2_nor3_1 _10185_ (.A(_00514_),
    .B(_01058_),
    .C(_04741_),
    .Y(_04742_));
 sg13g2_a21o_1 _10186_ (.A2(_01061_),
    .A1(_01050_),
    .B1(_01167_),
    .X(_04743_));
 sg13g2_nand3_1 _10187_ (.B(_01158_),
    .C(_01159_),
    .A(_01061_),
    .Y(_04744_));
 sg13g2_nand3b_1 _10188_ (.B(_04743_),
    .C(_04744_),
    .Y(_04745_),
    .A_N(_00514_));
 sg13g2_inv_1 _10189_ (.Y(_04746_),
    .A(_02276_));
 sg13g2_o21ai_1 _10190_ (.B1(_00848_),
    .Y(_04747_),
    .A1(_00069_),
    .A2(_01623_));
 sg13g2_o21ai_1 _10191_ (.B1(_04747_),
    .Y(_04748_),
    .A1(_04746_),
    .A2(_00844_));
 sg13g2_nand3_1 _10192_ (.B(_04745_),
    .C(_04748_),
    .A(net360),
    .Y(_04749_));
 sg13g2_o21ai_1 _10193_ (.B1(_00664_),
    .Y(_04750_),
    .A1(_01273_),
    .A2(_01274_));
 sg13g2_o21ai_1 _10194_ (.B1(_04750_),
    .Y(_04751_),
    .A1(_01210_),
    .A2(_01263_));
 sg13g2_nor4_1 _10195_ (.A(_04739_),
    .B(_04742_),
    .C(_04749_),
    .D(_04751_),
    .Y(_04752_));
 sg13g2_nand2_1 _10196_ (.Y(_04753_),
    .A(_05120_),
    .B(_00807_));
 sg13g2_inv_1 _10197_ (.Y(_04754_),
    .A(_00548_));
 sg13g2_or4_1 _10198_ (.A(net160),
    .B(_00511_),
    .C(_04754_),
    .D(_01173_),
    .X(_04755_));
 sg13g2_o21ai_1 _10199_ (.B1(_04755_),
    .Y(_04756_),
    .A1(_01146_),
    .A2(_04753_));
 sg13g2_nand2_1 _10200_ (.Y(_04757_),
    .A(_00555_),
    .B(net32));
 sg13g2_o21ai_1 _10201_ (.B1(_04757_),
    .Y(_04758_),
    .A1(_00548_),
    .A2(_00733_));
 sg13g2_nor2_1 _10202_ (.A(_00958_),
    .B(_04758_),
    .Y(_04759_));
 sg13g2_nand2_1 _10203_ (.Y(_04760_),
    .A(net158),
    .B(_00836_));
 sg13g2_nand2_1 _10204_ (.Y(_04761_),
    .A(_00607_),
    .B(_04760_));
 sg13g2_nand2b_1 _10205_ (.Y(_04762_),
    .B(_00610_),
    .A_N(_01260_));
 sg13g2_nand2_1 _10206_ (.Y(_04763_),
    .A(_00779_),
    .B(_00794_));
 sg13g2_a21oi_1 _10207_ (.A1(_04761_),
    .A2(_04762_),
    .Y(_04764_),
    .B1(_04763_));
 sg13g2_nand2b_1 _10208_ (.Y(_04765_),
    .B(_00953_),
    .A_N(_04758_));
 sg13g2_or4_1 _10209_ (.A(net54),
    .B(_00765_),
    .C(_01134_),
    .D(_01110_),
    .X(_04766_));
 sg13g2_nand2_1 _10210_ (.Y(_04767_),
    .A(net260),
    .B(_00630_));
 sg13g2_inv_1 _10211_ (.Y(_04768_),
    .A(_04767_));
 sg13g2_nor3_2 _10212_ (.A(net158),
    .B(_00548_),
    .C(_00951_),
    .Y(_04769_));
 sg13g2_nand2b_1 _10213_ (.Y(_04770_),
    .B(_04769_),
    .A_N(net33));
 sg13g2_nand2b_1 _10214_ (.Y(_04771_),
    .B(_00683_),
    .A_N(_00938_));
 sg13g2_inv_1 _10215_ (.Y(_04772_),
    .A(_04771_));
 sg13g2_o21ai_1 _10216_ (.B1(_00907_),
    .Y(_04773_),
    .A1(_04769_),
    .A2(_04772_));
 sg13g2_nand2b_1 _10217_ (.Y(_04774_),
    .B(_04772_),
    .A_N(_00934_));
 sg13g2_nand3_1 _10218_ (.B(_04773_),
    .C(_04774_),
    .A(_04770_),
    .Y(_04775_));
 sg13g2_o21ai_1 _10219_ (.B1(net260),
    .Y(_04776_),
    .A1(_00610_),
    .A2(_00733_));
 sg13g2_nor3_1 _10220_ (.A(net260),
    .B(_00511_),
    .C(_01044_),
    .Y(_04777_));
 sg13g2_o21ai_1 _10221_ (.B1(_04777_),
    .Y(_04778_),
    .A1(net71),
    .A2(_01142_));
 sg13g2_o21ai_1 _10222_ (.B1(_04778_),
    .Y(_04779_),
    .A1(net32),
    .A2(_04776_));
 sg13g2_nor4_1 _10223_ (.A(net158),
    .B(_00497_),
    .C(_01061_),
    .D(_01018_),
    .Y(_04780_));
 sg13g2_or3_1 _10224_ (.A(\game_logic_inst.valid_move ),
    .B(_04779_),
    .C(_04780_),
    .X(_04781_));
 sg13g2_a221oi_1 _10225_ (.B2(_00789_),
    .C1(_04781_),
    .B1(_04775_),
    .A1(_04768_),
    .Y(_04782_),
    .A2(_01110_));
 sg13g2_a21oi_1 _10226_ (.A1(_00635_),
    .A2(_00636_),
    .Y(_04783_),
    .B1(_01110_));
 sg13g2_and3_1 _10227_ (.X(_04784_),
    .A(_00498_),
    .B(_00664_),
    .C(_00788_));
 sg13g2_nand3b_1 _10228_ (.B(_00934_),
    .C(_04769_),
    .Y(_04785_),
    .A_N(net33));
 sg13g2_o21ai_1 _10229_ (.B1(_04785_),
    .Y(_04786_),
    .A1(_00926_),
    .A2(_04774_));
 sg13g2_a221oi_1 _10230_ (.B2(_01050_),
    .C1(_04786_),
    .B1(_04784_),
    .A1(_01058_),
    .Y(_04787_),
    .A2(_04783_));
 sg13g2_nand4_1 _10231_ (.B(_04766_),
    .C(_04782_),
    .A(_04765_),
    .Y(_04788_),
    .D(_04787_));
 sg13g2_nor4_1 _10232_ (.A(_04756_),
    .B(_04759_),
    .C(_04764_),
    .D(_04788_),
    .Y(_04789_));
 sg13g2_nand2_1 _10233_ (.Y(_04790_),
    .A(_00548_),
    .B(_04761_));
 sg13g2_o21ai_1 _10234_ (.B1(_00511_),
    .Y(_04791_),
    .A1(_01044_),
    .A2(_01171_));
 sg13g2_a21oi_1 _10235_ (.A1(_04761_),
    .A2(_04791_),
    .Y(_04792_),
    .B1(net160));
 sg13g2_o21ai_1 _10236_ (.B1(_04792_),
    .Y(_04793_),
    .A1(_01173_),
    .A2(_04790_));
 sg13g2_nand4_1 _10237_ (.B(_00907_),
    .C(_00954_),
    .A(net33),
    .Y(_04794_),
    .D(_04769_));
 sg13g2_mux2_1 _10238_ (.A0(_04794_),
    .A1(_04770_),
    .S(_00928_),
    .X(_04795_));
 sg13g2_nand3_1 _10239_ (.B(_00926_),
    .C(_00934_),
    .A(_00907_),
    .Y(_04796_));
 sg13g2_mux2_1 _10240_ (.A0(_04796_),
    .A1(_04774_),
    .S(_01050_),
    .X(_04797_));
 sg13g2_nor2_1 _10241_ (.A(_04767_),
    .B(_01058_),
    .Y(_04798_));
 sg13g2_a22oi_1 _10242_ (.Y(_04799_),
    .B1(_01211_),
    .B2(_04798_),
    .A2(_00795_),
    .A1(_00799_));
 sg13g2_nand4_1 _10243_ (.B(_04795_),
    .C(_04797_),
    .A(_04793_),
    .Y(_04800_),
    .D(_04799_));
 sg13g2_a221oi_1 _10244_ (.B2(_00628_),
    .C1(_04800_),
    .B1(_01368_),
    .A1(_00639_),
    .Y(_04801_),
    .A2(_00800_));
 sg13g2_nand2_1 _10245_ (.Y(_04802_),
    .A(_01125_),
    .B(_01130_));
 sg13g2_nand2_1 _10246_ (.Y(_04803_),
    .A(net160),
    .B(_00497_));
 sg13g2_a221oi_1 _10247_ (.B2(_01050_),
    .C1(_04803_),
    .B1(_01131_),
    .A1(_01098_),
    .Y(_04804_),
    .A2(_01124_));
 sg13g2_and3_1 _10248_ (.X(_04805_),
    .A(_00498_),
    .B(_01125_),
    .C(_01130_));
 sg13g2_a21oi_1 _10249_ (.A1(_04802_),
    .A2(_04804_),
    .Y(_04806_),
    .B1(_04805_));
 sg13g2_a21o_1 _10250_ (.A2(_00937_),
    .A1(_00935_),
    .B1(_00941_),
    .X(_04807_));
 sg13g2_a21oi_1 _10251_ (.A1(net30),
    .A2(_01030_),
    .Y(_04808_),
    .B1(_01210_));
 sg13g2_nand2_1 _10252_ (.Y(_04809_),
    .A(_00630_),
    .B(net31));
 sg13g2_o21ai_1 _10253_ (.B1(_00630_),
    .Y(_04810_),
    .A1(net93),
    .A2(_01110_));
 sg13g2_o21ai_1 _10254_ (.B1(_04810_),
    .Y(_04811_),
    .A1(_04808_),
    .A2(_04809_));
 sg13g2_mux2_1 _10255_ (.A0(_04811_),
    .A1(_00993_),
    .S(_01101_),
    .X(_04812_));
 sg13g2_a221oi_1 _10256_ (.B2(_00663_),
    .C1(_04812_),
    .B1(_04807_),
    .A1(_00608_),
    .Y(_04813_),
    .A2(_00913_));
 sg13g2_nand4_1 _10257_ (.B(_04801_),
    .C(_04806_),
    .A(_04789_),
    .Y(_04814_),
    .D(_04813_));
 sg13g2_nand3b_1 _10258_ (.B(_01064_),
    .C(_01048_),
    .Y(_04815_),
    .A_N(_00570_));
 sg13g2_or3_1 _10259_ (.A(_00571_),
    .B(_01064_),
    .C(_01048_),
    .X(_04816_));
 sg13g2_a21o_1 _10260_ (.A2(_04816_),
    .A1(_04815_),
    .B1(net69),
    .X(_04817_));
 sg13g2_xnor2_1 _10261_ (.Y(_04818_),
    .A(_00481_),
    .B(_01048_));
 sg13g2_or2_1 _10262_ (.X(_04819_),
    .B(_01064_),
    .A(_00479_));
 sg13g2_a21oi_1 _10263_ (.A1(_00570_),
    .A2(_00571_),
    .Y(_04820_),
    .B1(net93));
 sg13g2_a21oi_1 _10264_ (.A1(_00479_),
    .A2(_01064_),
    .Y(_04821_),
    .B1(_04820_));
 sg13g2_nand3_1 _10265_ (.B(_04819_),
    .C(_04821_),
    .A(_04818_),
    .Y(_04822_));
 sg13g2_nand2b_1 _10266_ (.Y(_04823_),
    .B(_00911_),
    .A_N(_00608_));
 sg13g2_nor2_1 _10267_ (.A(_00733_),
    .B(_00953_),
    .Y(_04824_));
 sg13g2_o21ai_1 _10268_ (.B1(net93),
    .Y(_04825_),
    .A1(_04754_),
    .A2(_00837_));
 sg13g2_a221oi_1 _10269_ (.B2(_04824_),
    .C1(_04825_),
    .B1(_00958_),
    .A1(_01210_),
    .Y(_04826_),
    .A2(_00911_));
 sg13g2_xnor2_1 _10270_ (.Y(_04827_),
    .A(_00497_),
    .B(_01146_));
 sg13g2_a22oi_1 _10271_ (.Y(_04828_),
    .B1(_04826_),
    .B2(_04827_),
    .A2(_04823_),
    .A1(net94));
 sg13g2_a21o_1 _10272_ (.A2(_04822_),
    .A1(_04817_),
    .B1(_04828_),
    .X(_04829_));
 sg13g2_nand2b_1 _10273_ (.Y(_04830_),
    .B(_01146_),
    .A_N(_00807_));
 sg13g2_xor2_1 _10274_ (.B(_01169_),
    .A(_00511_),
    .X(_04831_));
 sg13g2_a21oi_1 _10275_ (.A1(_04830_),
    .A2(_04831_),
    .Y(_04832_),
    .B1(_00949_));
 sg13g2_xor2_1 _10276_ (.B(_01133_),
    .A(_00807_),
    .X(_04833_));
 sg13g2_nor2_1 _10277_ (.A(net94),
    .B(_04833_),
    .Y(_04834_));
 sg13g2_nor4_2 _10278_ (.A(_04814_),
    .B(_04829_),
    .C(_04832_),
    .Y(_04835_),
    .D(_04834_));
 sg13g2_nand3_1 _10279_ (.B(_00889_),
    .C(_01074_),
    .A(_01079_),
    .Y(_04836_));
 sg13g2_nand2_1 _10280_ (.Y(_04837_),
    .A(_04748_),
    .B(_04836_));
 sg13g2_inv_1 _10281_ (.Y(_04838_),
    .A(\game_logic_inst.debug_move_reg ));
 sg13g2_nor2_1 _10282_ (.A(_05100_),
    .B(\game_logic_inst.add_new_tiles[0] ),
    .Y(_04839_));
 sg13g2_a21oi_1 _10283_ (.A1(net412),
    .A2(_04838_),
    .Y(_04840_),
    .B1(_04839_));
 sg13g2_nor3_1 _10284_ (.A(_01077_),
    .B(_04837_),
    .C(_04840_),
    .Y(_04841_));
 sg13g2_and2_1 _10285_ (.A(\game_logic_inst.add_new_tiles[0] ),
    .B(_04837_),
    .X(_04842_));
 sg13g2_o21ai_1 _10286_ (.B1(net402),
    .Y(_04843_),
    .A1(_04841_),
    .A2(_04842_));
 sg13g2_a21oi_1 _10287_ (.A1(_04752_),
    .A2(_04835_),
    .Y(_00283_),
    .B1(_04843_));
 sg13g2_and2_1 _10288_ (.A(\game_logic_inst.add_new_tiles[0] ),
    .B(_00069_),
    .X(_04844_));
 sg13g2_o21ai_1 _10289_ (.B1(\game_logic_inst.add_new_tiles[1] ),
    .Y(_04845_),
    .A1(_04837_),
    .A2(_04844_));
 sg13g2_a21oi_1 _10290_ (.A1(_00069_),
    .A2(_00864_),
    .Y(_04846_),
    .B1(_02276_));
 sg13g2_or2_1 _10291_ (.X(_04847_),
    .B(_04846_),
    .A(_04837_));
 sg13g2_a21oi_1 _10292_ (.A1(_04845_),
    .A2(_04847_),
    .Y(_00284_),
    .B1(_04736_));
 sg13g2_nand2b_1 _10293_ (.Y(_04848_),
    .B(net480),
    .A_N(net349));
 sg13g2_o21ai_1 _10294_ (.B1(net360),
    .Y(_04849_),
    .A1(_01614_),
    .A2(_04848_));
 sg13g2_a21oi_1 _10295_ (.A1(_05080_),
    .A2(_04849_),
    .Y(_00289_),
    .B1(net274));
 sg13g2_o21ai_1 _10296_ (.B1(_04746_),
    .Y(_04850_),
    .A1(_05078_),
    .A2(_01424_));
 sg13g2_nand2_1 _10297_ (.Y(_04851_),
    .A(_05107_),
    .B(_04850_));
 sg13g2_nor2_1 _10298_ (.A(_02276_),
    .B(_01228_),
    .Y(_04852_));
 sg13g2_nand3_1 _10299_ (.B(_00844_),
    .C(_04852_),
    .A(_01302_),
    .Y(_04853_));
 sg13g2_a21oi_1 _10300_ (.A1(_04851_),
    .A2(_04853_),
    .Y(_00290_),
    .B1(net274));
 sg13g2_nand2_1 _10301_ (.Y(_04854_),
    .A(_05107_),
    .B(_01089_));
 sg13g2_nor3_1 _10302_ (.A(_02276_),
    .B(_05113_),
    .C(_04854_),
    .Y(_04855_));
 sg13g2_a21oi_1 _10303_ (.A1(_05113_),
    .A2(_04854_),
    .Y(_04856_),
    .B1(_04855_));
 sg13g2_nor2_1 _10304_ (.A(_05078_),
    .B(_04856_),
    .Y(_04857_));
 sg13g2_a21oi_1 _10305_ (.A1(_02276_),
    .A2(net161),
    .Y(_04858_),
    .B1(_04857_));
 sg13g2_nor2_1 _10306_ (.A(net277),
    .B(_04858_),
    .Y(_00291_));
 sg13g2_nor4_1 _10307_ (.A(debug_btn_up),
    .B(debug_btn_right),
    .C(debug_btn_down),
    .D(debug_btn_left),
    .Y(_04859_));
 sg13g2_nor2_1 _10308_ (.A(_02276_),
    .B(_00844_),
    .Y(_04860_));
 sg13g2_mux2_1 _10309_ (.A0(_04838_),
    .A1(_04859_),
    .S(_04860_),
    .X(_04861_));
 sg13g2_nor2_1 _10310_ (.A(net277),
    .B(_04861_),
    .Y(_00292_));
 sg13g2_o21ai_1 _10311_ (.B1(net343),
    .Y(_04862_),
    .A1(net480),
    .A2(_05078_));
 sg13g2_inv_1 _10312_ (.Y(_00293_),
    .A(_04862_));
 sg13g2_and2_1 _10313_ (.A(net278),
    .B(_00170_),
    .X(_00294_));
 sg13g2_xor2_1 _10314_ (.B(_00851_),
    .A(_00850_),
    .X(_04863_));
 sg13g2_nor2_1 _10315_ (.A(_04639_),
    .B(_04863_),
    .Y(_00295_));
 sg13g2_and2_1 _10316_ (.A(net278),
    .B(_05076_),
    .X(_00296_));
 sg13g2_nand2_1 _10317_ (.Y(_04864_),
    .A(_05075_),
    .B(_05078_));
 sg13g2_a21oi_1 _10318_ (.A1(net480),
    .A2(_04864_),
    .Y(_04865_),
    .B1(_01298_));
 sg13g2_o21ai_1 _10319_ (.B1(_01727_),
    .Y(_04866_),
    .A1(_05062_),
    .A2(\game_logic_inst.current_direction[1] ));
 sg13g2_a21oi_1 _10320_ (.A1(net49),
    .A2(_04866_),
    .Y(_04867_),
    .B1(net413));
 sg13g2_nor2b_1 _10321_ (.A(_04865_),
    .B_N(_04867_),
    .Y(_00297_));
 sg13g2_o21ai_1 _10322_ (.B1(net403),
    .Y(_04868_),
    .A1(\game_logic_inst.valid_move ),
    .A2(_04852_));
 sg13g2_nor3_1 _10323_ (.A(_04835_),
    .B(_04860_),
    .C(_04868_),
    .Y(_00298_));
 sg13g2_buf_1 _10324_ (.A(_05071_),
    .X(_04869_));
 sg13g2_buf_1 _10325_ (.A(net415),
    .X(_04870_));
 sg13g2_buf_1 _10326_ (.A(net479),
    .X(_04871_));
 sg13g2_buf_1 _10327_ (.A(net438),
    .X(_04872_));
 sg13g2_a21o_1 _10328_ (.A2(\welcome_screen_grid[0] ),
    .A1(_04871_),
    .B1(_04872_),
    .X(_04873_));
 sg13g2_a21oi_1 _10329_ (.A1(net371),
    .A2(_05215_),
    .Y(_04874_),
    .B1(_04873_));
 sg13g2_buf_1 _10330_ (.A(net396),
    .X(_04875_));
 sg13g2_o21ai_1 _10331_ (.B1(net343),
    .Y(_04876_),
    .A1(\draw_game_inst.grid[0] ),
    .A2(net273));
 sg13g2_nor2_1 _10332_ (.A(_04874_),
    .B(_04876_),
    .Y(_00299_));
 sg13g2_buf_1 _10333_ (.A(net395),
    .X(_04877_));
 sg13g2_nand2_1 _10334_ (.Y(_04878_),
    .A(\draw_game_inst.grid[10] ),
    .B(net272));
 sg13g2_buf_1 _10335_ (.A(net415),
    .X(_04879_));
 sg13g2_buf_1 _10336_ (.A(_01793_),
    .X(_04880_));
 sg13g2_nand3_1 _10337_ (.B(_00460_),
    .C(net368),
    .A(net369),
    .Y(_04881_));
 sg13g2_a21oi_1 _10338_ (.A1(_04878_),
    .A2(_04881_),
    .Y(_00300_),
    .B1(net274));
 sg13g2_a21o_1 _10339_ (.A2(\welcome_screen_grid[11] ),
    .A1(net414),
    .B1(net370),
    .X(_04882_));
 sg13g2_a21oi_1 _10340_ (.A1(_04870_),
    .A2(_05158_),
    .Y(_04883_),
    .B1(_04882_));
 sg13g2_o21ai_1 _10341_ (.B1(net343),
    .Y(_04884_),
    .A1(\draw_game_inst.grid[11] ),
    .A2(_04875_));
 sg13g2_nor2_1 _10342_ (.A(_04883_),
    .B(_04884_),
    .Y(_00301_));
 sg13g2_a21o_1 _10343_ (.A2(\welcome_screen_grid[12] ),
    .A1(net414),
    .B1(net370),
    .X(_04885_));
 sg13g2_a21oi_1 _10344_ (.A1(net371),
    .A2(_05160_),
    .Y(_04886_),
    .B1(_04885_));
 sg13g2_o21ai_1 _10345_ (.B1(net343),
    .Y(_04887_),
    .A1(\draw_game_inst.grid[12] ),
    .A2(net273));
 sg13g2_nor2_1 _10346_ (.A(_04886_),
    .B(_04887_),
    .Y(_00302_));
 sg13g2_a21oi_1 _10347_ (.A1(net371),
    .A2(_05181_),
    .Y(_04888_),
    .B1(_04885_));
 sg13g2_buf_1 _10348_ (.A(net407),
    .X(_04889_));
 sg13g2_o21ai_1 _10349_ (.B1(_04889_),
    .Y(_04890_),
    .A1(\draw_game_inst.grid[13] ),
    .A2(net273));
 sg13g2_nor2_1 _10350_ (.A(_04888_),
    .B(_04890_),
    .Y(_00303_));
 sg13g2_nand2_1 _10351_ (.Y(_04891_),
    .A(\draw_game_inst.grid[14] ),
    .B(net272));
 sg13g2_buf_1 _10352_ (.A(_01793_),
    .X(_04892_));
 sg13g2_nand3_1 _10353_ (.B(_00459_),
    .C(net367),
    .A(net369),
    .Y(_04893_));
 sg13g2_a21oi_1 _10354_ (.A1(_04891_),
    .A2(_04893_),
    .Y(_00304_),
    .B1(net274));
 sg13g2_a21oi_1 _10355_ (.A1(_04870_),
    .A2(_05157_),
    .Y(_04894_),
    .B1(_04885_));
 sg13g2_o21ai_1 _10356_ (.B1(net271),
    .Y(_04895_),
    .A1(\draw_game_inst.grid[15] ),
    .A2(_04875_));
 sg13g2_nor2_1 _10357_ (.A(_04894_),
    .B(_04895_),
    .Y(_00305_));
 sg13g2_a21o_1 _10358_ (.A2(\welcome_screen_grid[16] ),
    .A1(net414),
    .B1(net370),
    .X(_04896_));
 sg13g2_a21oi_1 _10359_ (.A1(net371),
    .A2(_00468_),
    .Y(_04897_),
    .B1(_04896_));
 sg13g2_o21ai_1 _10360_ (.B1(net271),
    .Y(_04898_),
    .A1(\draw_game_inst.grid[16] ),
    .A2(net273));
 sg13g2_nor2_1 _10361_ (.A(_04897_),
    .B(_04898_),
    .Y(_00306_));
 sg13g2_a21oi_1 _10362_ (.A1(net371),
    .A2(_05122_),
    .Y(_04899_),
    .B1(_04896_));
 sg13g2_o21ai_1 _10363_ (.B1(net271),
    .Y(_04900_),
    .A1(\draw_game_inst.grid[17] ),
    .A2(net273));
 sg13g2_nor2_1 _10364_ (.A(_04899_),
    .B(_04900_),
    .Y(_00307_));
 sg13g2_nand2_1 _10365_ (.Y(_04901_),
    .A(\draw_game_inst.grid[18] ),
    .B(net272));
 sg13g2_buf_1 _10366_ (.A(net415),
    .X(_04902_));
 sg13g2_nand3_1 _10367_ (.B(_05201_),
    .C(net367),
    .A(net366),
    .Y(_04903_));
 sg13g2_a21oi_1 _10368_ (.A1(_04901_),
    .A2(_04903_),
    .Y(_00308_),
    .B1(net274));
 sg13g2_a21oi_1 _10369_ (.A1(net371),
    .A2(_05165_),
    .Y(_04904_),
    .B1(_04896_));
 sg13g2_o21ai_1 _10370_ (.B1(net271),
    .Y(_04905_),
    .A1(\draw_game_inst.grid[19] ),
    .A2(net273));
 sg13g2_nor2_1 _10371_ (.A(_04904_),
    .B(_04905_),
    .Y(_00309_));
 sg13g2_a21oi_1 _10372_ (.A1(net371),
    .A2(_05218_),
    .Y(_04906_),
    .B1(_04873_));
 sg13g2_o21ai_1 _10373_ (.B1(_04889_),
    .Y(_04907_),
    .A1(\draw_game_inst.grid[1] ),
    .A2(net273));
 sg13g2_nor2_1 _10374_ (.A(_04906_),
    .B(_04907_),
    .Y(_00310_));
 sg13g2_a21o_1 _10375_ (.A2(\welcome_screen_grid[20] ),
    .A1(net414),
    .B1(net370),
    .X(_04908_));
 sg13g2_a21oi_1 _10376_ (.A1(net371),
    .A2(_00469_),
    .Y(_04909_),
    .B1(_04908_));
 sg13g2_o21ai_1 _10377_ (.B1(net271),
    .Y(_04910_),
    .A1(\draw_game_inst.grid[20] ),
    .A2(net273));
 sg13g2_nor2_1 _10378_ (.A(_04909_),
    .B(_04910_),
    .Y(_00311_));
 sg13g2_buf_1 _10379_ (.A(net415),
    .X(_04911_));
 sg13g2_a21oi_1 _10380_ (.A1(net365),
    .A2(_05123_),
    .Y(_04912_),
    .B1(_04908_));
 sg13g2_buf_1 _10381_ (.A(net396),
    .X(_04913_));
 sg13g2_o21ai_1 _10382_ (.B1(net271),
    .Y(_04914_),
    .A1(\draw_game_inst.grid[21] ),
    .A2(net270));
 sg13g2_nor2_1 _10383_ (.A(_04912_),
    .B(_04914_),
    .Y(_00312_));
 sg13g2_nand2_1 _10384_ (.Y(_04915_),
    .A(\draw_game_inst.grid[22] ),
    .B(_04877_));
 sg13g2_nand3_1 _10385_ (.B(_05202_),
    .C(_04892_),
    .A(net366),
    .Y(_04916_));
 sg13g2_a21oi_1 _10386_ (.A1(_04915_),
    .A2(_04916_),
    .Y(_00313_),
    .B1(net274));
 sg13g2_a21oi_1 _10387_ (.A1(net365),
    .A2(_05166_),
    .Y(_04917_),
    .B1(_04908_));
 sg13g2_o21ai_1 _10388_ (.B1(net271),
    .Y(_04918_),
    .A1(\draw_game_inst.grid[23] ),
    .A2(net270));
 sg13g2_nor2_1 _10389_ (.A(_04917_),
    .B(_04918_),
    .Y(_00314_));
 sg13g2_a21o_1 _10390_ (.A2(\welcome_screen_grid[24] ),
    .A1(net414),
    .B1(net370),
    .X(_04919_));
 sg13g2_a21oi_1 _10391_ (.A1(net365),
    .A2(_05198_),
    .Y(_04920_),
    .B1(_04919_));
 sg13g2_o21ai_1 _10392_ (.B1(net271),
    .Y(_04921_),
    .A1(\draw_game_inst.grid[24] ),
    .A2(net270));
 sg13g2_nor2_1 _10393_ (.A(_04920_),
    .B(_04921_),
    .Y(_00315_));
 sg13g2_a21oi_1 _10394_ (.A1(net365),
    .A2(_05126_),
    .Y(_04922_),
    .B1(_04919_));
 sg13g2_buf_1 _10395_ (.A(net407),
    .X(_04923_));
 sg13g2_o21ai_1 _10396_ (.B1(net269),
    .Y(_04924_),
    .A1(\draw_game_inst.grid[25] ),
    .A2(net270));
 sg13g2_nor2_1 _10397_ (.A(_04922_),
    .B(_04924_),
    .Y(_00316_));
 sg13g2_nand2_1 _10398_ (.Y(_04925_),
    .A(\draw_game_inst.grid[26] ),
    .B(_04877_));
 sg13g2_nand3_1 _10399_ (.B(_05195_),
    .C(_04892_),
    .A(_04902_),
    .Y(_04926_));
 sg13g2_a21oi_1 _10400_ (.A1(_04925_),
    .A2(_04926_),
    .Y(_00317_),
    .B1(net274));
 sg13g2_a21oi_1 _10401_ (.A1(net365),
    .A2(_05169_),
    .Y(_04927_),
    .B1(_04919_));
 sg13g2_o21ai_1 _10402_ (.B1(net269),
    .Y(_04928_),
    .A1(\draw_game_inst.grid[27] ),
    .A2(net270));
 sg13g2_nor2_1 _10403_ (.A(_04927_),
    .B(_04928_),
    .Y(_00318_));
 sg13g2_a21o_1 _10404_ (.A2(\welcome_screen_grid[28] ),
    .A1(net414),
    .B1(net370),
    .X(_04929_));
 sg13g2_a21oi_1 _10405_ (.A1(net365),
    .A2(_05197_),
    .Y(_04930_),
    .B1(_04929_));
 sg13g2_o21ai_1 _10406_ (.B1(net269),
    .Y(_04931_),
    .A1(\draw_game_inst.grid[28] ),
    .A2(net270));
 sg13g2_nor2_1 _10407_ (.A(_04930_),
    .B(_04931_),
    .Y(_00319_));
 sg13g2_a21oi_1 _10408_ (.A1(net365),
    .A2(_05125_),
    .Y(_04932_),
    .B1(_04929_));
 sg13g2_o21ai_1 _10409_ (.B1(net269),
    .Y(_04933_),
    .A1(\draw_game_inst.grid[29] ),
    .A2(net270));
 sg13g2_nor2_1 _10410_ (.A(_04932_),
    .B(_04933_),
    .Y(_00320_));
 sg13g2_nand2_1 _10411_ (.Y(_04934_),
    .A(\draw_game_inst.grid[2] ),
    .B(net272));
 sg13g2_nand3_1 _10412_ (.B(_05178_),
    .C(net367),
    .A(net366),
    .Y(_04935_));
 sg13g2_a21oi_1 _10413_ (.A1(_04934_),
    .A2(_04935_),
    .Y(_00321_),
    .B1(net274));
 sg13g2_nand2_1 _10414_ (.Y(_04936_),
    .A(\draw_game_inst.grid[30] ),
    .B(net272));
 sg13g2_nand3_1 _10415_ (.B(_05194_),
    .C(net367),
    .A(_04902_),
    .Y(_04937_));
 sg13g2_buf_1 _10416_ (.A(_01120_),
    .X(_04938_));
 sg13g2_a21oi_1 _10417_ (.A1(_04936_),
    .A2(_04937_),
    .Y(_00322_),
    .B1(net268));
 sg13g2_a21oi_1 _10418_ (.A1(net365),
    .A2(_05168_),
    .Y(_04939_),
    .B1(_04929_));
 sg13g2_o21ai_1 _10419_ (.B1(net269),
    .Y(_04940_),
    .A1(\draw_game_inst.grid[31] ),
    .A2(net270));
 sg13g2_nor2_1 _10420_ (.A(_04939_),
    .B(_04940_),
    .Y(_00323_));
 sg13g2_a21o_1 _10421_ (.A2(\welcome_screen_grid[32] ),
    .A1(net414),
    .B1(net370),
    .X(_04941_));
 sg13g2_a21oi_1 _10422_ (.A1(_04911_),
    .A2(_05222_),
    .Y(_04942_),
    .B1(_04941_));
 sg13g2_o21ai_1 _10423_ (.B1(net269),
    .Y(_04943_),
    .A1(\draw_game_inst.grid[32] ),
    .A2(_04913_));
 sg13g2_nor2_1 _10424_ (.A(_04942_),
    .B(_04943_),
    .Y(_00324_));
 sg13g2_a21oi_1 _10425_ (.A1(_04911_),
    .A2(_05225_),
    .Y(_04944_),
    .B1(_04941_));
 sg13g2_o21ai_1 _10426_ (.B1(net269),
    .Y(_04945_),
    .A1(\draw_game_inst.grid[33] ),
    .A2(_04913_));
 sg13g2_nor2_1 _10427_ (.A(_04944_),
    .B(_04945_),
    .Y(_00325_));
 sg13g2_nand2_1 _10428_ (.Y(_04946_),
    .A(\draw_game_inst.grid[34] ),
    .B(net272));
 sg13g2_nand3_1 _10429_ (.B(_05184_),
    .C(net367),
    .A(net366),
    .Y(_04947_));
 sg13g2_a21oi_1 _10430_ (.A1(_04946_),
    .A2(_04947_),
    .Y(_00326_),
    .B1(net268));
 sg13g2_buf_1 _10431_ (.A(net415),
    .X(_04948_));
 sg13g2_a21oi_1 _10432_ (.A1(net364),
    .A2(_05152_),
    .Y(_04949_),
    .B1(_04941_));
 sg13g2_buf_1 _10433_ (.A(net396),
    .X(_04950_));
 sg13g2_o21ai_1 _10434_ (.B1(_04923_),
    .Y(_04951_),
    .A1(\draw_game_inst.grid[35] ),
    .A2(net267));
 sg13g2_nor2_1 _10435_ (.A(_04949_),
    .B(_04951_),
    .Y(_00327_));
 sg13g2_a21o_1 _10436_ (.A2(\welcome_screen_grid[36] ),
    .A1(net414),
    .B1(net370),
    .X(_04952_));
 sg13g2_a21oi_1 _10437_ (.A1(net364),
    .A2(_05223_),
    .Y(_04953_),
    .B1(_04952_));
 sg13g2_o21ai_1 _10438_ (.B1(net269),
    .Y(_04954_),
    .A1(\draw_game_inst.grid[36] ),
    .A2(net267));
 sg13g2_nor2_1 _10439_ (.A(_04953_),
    .B(_04954_),
    .Y(_00328_));
 sg13g2_a21oi_1 _10440_ (.A1(net364),
    .A2(_05226_),
    .Y(_04955_),
    .B1(_04952_));
 sg13g2_o21ai_1 _10441_ (.B1(_04923_),
    .Y(_04956_),
    .A1(\draw_game_inst.grid[37] ),
    .A2(net267));
 sg13g2_nor2_1 _10442_ (.A(_04955_),
    .B(_04956_),
    .Y(_00329_));
 sg13g2_nand2_1 _10443_ (.Y(_04957_),
    .A(\draw_game_inst.grid[38] ),
    .B(net272));
 sg13g2_nand3_1 _10444_ (.B(_05185_),
    .C(net367),
    .A(net366),
    .Y(_04958_));
 sg13g2_a21oi_1 _10445_ (.A1(_04957_),
    .A2(_04958_),
    .Y(_00330_),
    .B1(_04938_));
 sg13g2_a21oi_1 _10446_ (.A1(_04948_),
    .A2(_05153_),
    .Y(_04959_),
    .B1(_04952_));
 sg13g2_buf_1 _10447_ (.A(_00919_),
    .X(_04960_));
 sg13g2_o21ai_1 _10448_ (.B1(net266),
    .Y(_04961_),
    .A1(\draw_game_inst.grid[39] ),
    .A2(_04950_));
 sg13g2_nor2_1 _10449_ (.A(_04959_),
    .B(_04961_),
    .Y(_00331_));
 sg13g2_a21oi_1 _10450_ (.A1(net364),
    .A2(_05149_),
    .Y(_04962_),
    .B1(_04873_));
 sg13g2_o21ai_1 _10451_ (.B1(net266),
    .Y(_04963_),
    .A1(\draw_game_inst.grid[3] ),
    .A2(net267));
 sg13g2_nor2_1 _10452_ (.A(_04962_),
    .B(_04963_),
    .Y(_00332_));
 sg13g2_a21o_1 _10453_ (.A2(\welcome_screen_grid[40] ),
    .A1(net479),
    .B1(_04872_),
    .X(_04964_));
 sg13g2_a21oi_1 _10454_ (.A1(net364),
    .A2(_05142_),
    .Y(_04965_),
    .B1(_04964_));
 sg13g2_o21ai_1 _10455_ (.B1(net266),
    .Y(_04966_),
    .A1(\draw_game_inst.grid[40] ),
    .A2(net267));
 sg13g2_nor2_1 _10456_ (.A(_04965_),
    .B(_04966_),
    .Y(_00333_));
 sg13g2_a21oi_1 _10457_ (.A1(net364),
    .A2(_05188_),
    .Y(_04967_),
    .B1(_04964_));
 sg13g2_o21ai_1 _10458_ (.B1(net266),
    .Y(_04968_),
    .A1(\draw_game_inst.grid[41] ),
    .A2(net267));
 sg13g2_nor2_1 _10459_ (.A(_04967_),
    .B(_04968_),
    .Y(_00334_));
 sg13g2_nand2_1 _10460_ (.Y(_04969_),
    .A(\draw_game_inst.grid[42] ),
    .B(net272));
 sg13g2_nand3_1 _10461_ (.B(_00463_),
    .C(net367),
    .A(net366),
    .Y(_04970_));
 sg13g2_a21oi_1 _10462_ (.A1(_04969_),
    .A2(_04970_),
    .Y(_00335_),
    .B1(net268));
 sg13g2_a21oi_1 _10463_ (.A1(_04948_),
    .A2(_05145_),
    .Y(_04971_),
    .B1(_04964_));
 sg13g2_o21ai_1 _10464_ (.B1(_04960_),
    .Y(_04972_),
    .A1(\draw_game_inst.grid[43] ),
    .A2(_04950_));
 sg13g2_nor2_1 _10465_ (.A(_04971_),
    .B(_04972_),
    .Y(_00336_));
 sg13g2_a21o_1 _10466_ (.A2(\welcome_screen_grid[44] ),
    .A1(net479),
    .B1(net438),
    .X(_04973_));
 sg13g2_a21oi_1 _10467_ (.A1(net364),
    .A2(_05141_),
    .Y(_04974_),
    .B1(_04973_));
 sg13g2_o21ai_1 _10468_ (.B1(net266),
    .Y(_04975_),
    .A1(\draw_game_inst.grid[44] ),
    .A2(net267));
 sg13g2_nor2_1 _10469_ (.A(_04974_),
    .B(_04975_),
    .Y(_00337_));
 sg13g2_a21oi_1 _10470_ (.A1(net364),
    .A2(_05187_),
    .Y(_04976_),
    .B1(_04973_));
 sg13g2_o21ai_1 _10471_ (.B1(net266),
    .Y(_04977_),
    .A1(\draw_game_inst.grid[45] ),
    .A2(net267));
 sg13g2_nor2_1 _10472_ (.A(_04976_),
    .B(_04977_),
    .Y(_00338_));
 sg13g2_nand2_1 _10473_ (.Y(_04978_),
    .A(\draw_game_inst.grid[46] ),
    .B(net395));
 sg13g2_nand3_1 _10474_ (.B(_00462_),
    .C(net367),
    .A(net366),
    .Y(_04979_));
 sg13g2_a21oi_1 _10475_ (.A1(_04978_),
    .A2(_04979_),
    .Y(_00339_),
    .B1(net268));
 sg13g2_buf_1 _10476_ (.A(net415),
    .X(_04980_));
 sg13g2_a21oi_1 _10477_ (.A1(net363),
    .A2(_05144_),
    .Y(_04981_),
    .B1(_04973_));
 sg13g2_buf_1 _10478_ (.A(_01793_),
    .X(_04982_));
 sg13g2_o21ai_1 _10479_ (.B1(_04960_),
    .Y(_04983_),
    .A1(\draw_game_inst.grid[47] ),
    .A2(net362));
 sg13g2_nor2_1 _10480_ (.A(_04981_),
    .B(_04983_),
    .Y(_00340_));
 sg13g2_a21o_1 _10481_ (.A2(\welcome_screen_grid[48] ),
    .A1(net479),
    .B1(net438),
    .X(_04984_));
 sg13g2_a21oi_1 _10482_ (.A1(net363),
    .A2(_00471_),
    .Y(_04985_),
    .B1(_04984_));
 sg13g2_o21ai_1 _10483_ (.B1(net266),
    .Y(_04986_),
    .A1(\draw_game_inst.grid[48] ),
    .A2(net362));
 sg13g2_nor2_1 _10484_ (.A(_04985_),
    .B(_04986_),
    .Y(_00341_));
 sg13g2_a21oi_1 _10485_ (.A1(net363),
    .A2(_05128_),
    .Y(_04987_),
    .B1(_04984_));
 sg13g2_o21ai_1 _10486_ (.B1(net266),
    .Y(_04988_),
    .A1(\draw_game_inst.grid[49] ),
    .A2(net362));
 sg13g2_nor2_1 _10487_ (.A(_04987_),
    .B(_04988_),
    .Y(_00342_));
 sg13g2_a21o_1 _10488_ (.A2(\welcome_screen_grid[4] ),
    .A1(net479),
    .B1(net438),
    .X(_04989_));
 sg13g2_a21oi_1 _10489_ (.A1(net363),
    .A2(_05216_),
    .Y(_04990_),
    .B1(_04989_));
 sg13g2_buf_1 _10490_ (.A(net407),
    .X(_04991_));
 sg13g2_o21ai_1 _10491_ (.B1(net265),
    .Y(_04992_),
    .A1(\draw_game_inst.grid[4] ),
    .A2(net362));
 sg13g2_nor2_1 _10492_ (.A(_04990_),
    .B(_04992_),
    .Y(_00343_));
 sg13g2_nand2_1 _10493_ (.Y(_04993_),
    .A(\draw_game_inst.grid[50] ),
    .B(net395));
 sg13g2_nand3_1 _10494_ (.B(_05211_),
    .C(net396),
    .A(net366),
    .Y(_04994_));
 sg13g2_a21oi_1 _10495_ (.A1(_04993_),
    .A2(_04994_),
    .Y(_00344_),
    .B1(net268));
 sg13g2_a21oi_1 _10496_ (.A1(_04980_),
    .A2(_05171_),
    .Y(_04995_),
    .B1(_04984_));
 sg13g2_o21ai_1 _10497_ (.B1(net265),
    .Y(_04996_),
    .A1(\draw_game_inst.grid[51] ),
    .A2(net362));
 sg13g2_nor2_1 _10498_ (.A(_04995_),
    .B(_04996_),
    .Y(_00345_));
 sg13g2_a21o_1 _10499_ (.A2(\welcome_screen_grid[52] ),
    .A1(net479),
    .B1(net438),
    .X(_04997_));
 sg13g2_a21oi_1 _10500_ (.A1(net363),
    .A2(_00472_),
    .Y(_04998_),
    .B1(_04997_));
 sg13g2_o21ai_1 _10501_ (.B1(net265),
    .Y(_04999_),
    .A1(\draw_game_inst.grid[52] ),
    .A2(net362));
 sg13g2_nor2_1 _10502_ (.A(_04998_),
    .B(_04999_),
    .Y(_00346_));
 sg13g2_a21oi_1 _10503_ (.A1(net363),
    .A2(_05129_),
    .Y(_05000_),
    .B1(_04997_));
 sg13g2_o21ai_1 _10504_ (.B1(net265),
    .Y(_05001_),
    .A1(\draw_game_inst.grid[53] ),
    .A2(net362));
 sg13g2_nor2_1 _10505_ (.A(_05000_),
    .B(_05001_),
    .Y(_00347_));
 sg13g2_nand2_1 _10506_ (.Y(_05002_),
    .A(\draw_game_inst.grid[54] ),
    .B(net395));
 sg13g2_nand3_1 _10507_ (.B(_05212_),
    .C(net396),
    .A(net415),
    .Y(_05003_));
 sg13g2_a21oi_1 _10508_ (.A1(_05002_),
    .A2(_05003_),
    .Y(_00348_),
    .B1(net268));
 sg13g2_a21oi_1 _10509_ (.A1(net363),
    .A2(_05172_),
    .Y(_05004_),
    .B1(_04997_));
 sg13g2_o21ai_1 _10510_ (.B1(net265),
    .Y(_05005_),
    .A1(\draw_game_inst.grid[55] ),
    .A2(_04982_));
 sg13g2_nor2_1 _10511_ (.A(_05004_),
    .B(_05005_),
    .Y(_00349_));
 sg13g2_a21o_1 _10512_ (.A2(\welcome_screen_grid[56] ),
    .A1(net479),
    .B1(net438),
    .X(_05006_));
 sg13g2_a21oi_1 _10513_ (.A1(_04980_),
    .A2(_05208_),
    .Y(_05007_),
    .B1(_05006_));
 sg13g2_o21ai_1 _10514_ (.B1(net265),
    .Y(_05008_),
    .A1(\draw_game_inst.grid[56] ),
    .A2(net362));
 sg13g2_nor2_1 _10515_ (.A(_05007_),
    .B(_05008_),
    .Y(_00350_));
 sg13g2_a21oi_1 _10516_ (.A1(net363),
    .A2(_05132_),
    .Y(_05009_),
    .B1(_05006_));
 sg13g2_o21ai_1 _10517_ (.B1(net265),
    .Y(_05010_),
    .A1(\draw_game_inst.grid[57] ),
    .A2(_04982_));
 sg13g2_nor2_1 _10518_ (.A(_05009_),
    .B(_05010_),
    .Y(_00351_));
 sg13g2_nand2_1 _10519_ (.Y(_05011_),
    .A(\draw_game_inst.grid[58] ),
    .B(net395));
 sg13g2_nand3_1 _10520_ (.B(_05205_),
    .C(net396),
    .A(net415),
    .Y(_05012_));
 sg13g2_a21oi_1 _10521_ (.A1(_05011_),
    .A2(_05012_),
    .Y(_00352_),
    .B1(net268));
 sg13g2_a21oi_1 _10522_ (.A1(net369),
    .A2(_05175_),
    .Y(_05013_),
    .B1(_05006_));
 sg13g2_o21ai_1 _10523_ (.B1(_04991_),
    .Y(_05014_),
    .A1(\draw_game_inst.grid[59] ),
    .A2(net368));
 sg13g2_nor2_1 _10524_ (.A(_05013_),
    .B(_05014_),
    .Y(_00353_));
 sg13g2_a21oi_1 _10525_ (.A1(net369),
    .A2(_05219_),
    .Y(_05015_),
    .B1(_04989_));
 sg13g2_o21ai_1 _10526_ (.B1(net265),
    .Y(_05016_),
    .A1(\draw_game_inst.grid[5] ),
    .A2(net368));
 sg13g2_nor2_1 _10527_ (.A(_05015_),
    .B(_05016_),
    .Y(_00354_));
 sg13g2_a21o_1 _10528_ (.A2(\welcome_screen_grid[60] ),
    .A1(net479),
    .B1(net438),
    .X(_05017_));
 sg13g2_a21oi_1 _10529_ (.A1(net369),
    .A2(_05207_),
    .Y(_05018_),
    .B1(_05017_));
 sg13g2_o21ai_1 _10530_ (.B1(_04991_),
    .Y(_05019_),
    .A1(\draw_game_inst.grid[60] ),
    .A2(net368));
 sg13g2_nor2_1 _10531_ (.A(_05018_),
    .B(_05019_),
    .Y(_00355_));
 sg13g2_a21oi_1 _10532_ (.A1(_04879_),
    .A2(_05131_),
    .Y(_05020_),
    .B1(_05017_));
 sg13g2_o21ai_1 _10533_ (.B1(net402),
    .Y(_05021_),
    .A1(\draw_game_inst.grid[61] ),
    .A2(net368));
 sg13g2_nor2_1 _10534_ (.A(_05020_),
    .B(_05021_),
    .Y(_00356_));
 sg13g2_nand2_1 _10535_ (.Y(_05022_),
    .A(\draw_game_inst.grid[62] ),
    .B(net395));
 sg13g2_nand3_1 _10536_ (.B(_05204_),
    .C(_01794_),
    .A(_04869_),
    .Y(_05023_));
 sg13g2_a21oi_1 _10537_ (.A1(_05022_),
    .A2(_05023_),
    .Y(_00357_),
    .B1(net268));
 sg13g2_a21oi_1 _10538_ (.A1(_04879_),
    .A2(_05174_),
    .Y(_05024_),
    .B1(_05017_));
 sg13g2_o21ai_1 _10539_ (.B1(net402),
    .Y(_05025_),
    .A1(\draw_game_inst.grid[63] ),
    .A2(_04880_));
 sg13g2_nor2_1 _10540_ (.A(_05024_),
    .B(_05025_),
    .Y(_00358_));
 sg13g2_nand2_1 _10541_ (.Y(_05026_),
    .A(\draw_game_inst.grid[6] ),
    .B(net395));
 sg13g2_nand3_1 _10542_ (.B(_05179_),
    .C(_01794_),
    .A(_04869_),
    .Y(_05027_));
 sg13g2_a21oi_1 _10543_ (.A1(_05026_),
    .A2(_05027_),
    .Y(_00359_),
    .B1(_04938_));
 sg13g2_a21oi_1 _10544_ (.A1(net369),
    .A2(_05150_),
    .Y(_05028_),
    .B1(_04989_));
 sg13g2_o21ai_1 _10545_ (.B1(net402),
    .Y(_05029_),
    .A1(\draw_game_inst.grid[7] ),
    .A2(net368));
 sg13g2_nor2_1 _10546_ (.A(_05028_),
    .B(_05029_),
    .Y(_00360_));
 sg13g2_a21oi_1 _10547_ (.A1(net369),
    .A2(_05161_),
    .Y(_05030_),
    .B1(_04882_));
 sg13g2_o21ai_1 _10548_ (.B1(net402),
    .Y(_05031_),
    .A1(\draw_game_inst.grid[8] ),
    .A2(net368));
 sg13g2_nor2_1 _10549_ (.A(_05030_),
    .B(_05031_),
    .Y(_00361_));
 sg13g2_a21oi_1 _10550_ (.A1(net369),
    .A2(_05182_),
    .Y(_05032_),
    .B1(_04882_));
 sg13g2_o21ai_1 _10551_ (.B1(net402),
    .Y(_05033_),
    .A1(\draw_game_inst.grid[9] ),
    .A2(net368));
 sg13g2_nor2_1 _10552_ (.A(_05032_),
    .B(_05033_),
    .Y(_00362_));
 sg13g2_xnor2_1 _10553_ (.Y(_05034_),
    .A(\game_logic_inst.lfsr_value[0] ),
    .B(\game_logic_inst.lfsr_value[1] ));
 sg13g2_xnor2_1 _10554_ (.Y(_05035_),
    .A(_02010_),
    .B(\lfsr_inst.lfsr[21] ));
 sg13g2_xnor2_1 _10555_ (.Y(_05036_),
    .A(_05034_),
    .B(_05035_));
 sg13g2_nor2_1 _10556_ (.A(_04639_),
    .B(_05036_),
    .Y(_00363_));
 sg13g2_and2_1 _10557_ (.A(net278),
    .B(\game_logic_inst.lfsr_value[9] ),
    .X(_00364_));
 sg13g2_buf_1 _10558_ (.A(net403),
    .X(_05037_));
 sg13g2_nand2b_1 _10559_ (.Y(_00365_),
    .B(net264),
    .A_N(\game_logic_inst.lfsr_value[10] ));
 sg13g2_nand2b_1 _10560_ (.Y(_00366_),
    .B(net264),
    .A_N(\game_logic_inst.lfsr_value[11] ));
 sg13g2_nand2b_1 _10561_ (.Y(_00367_),
    .B(net264),
    .A_N(\game_logic_inst.lfsr_value[12] ));
 sg13g2_nand2b_1 _10562_ (.Y(_00368_),
    .B(net264),
    .A_N(\game_logic_inst.lfsr_value[13] ));
 sg13g2_nand2b_1 _10563_ (.Y(_00369_),
    .B(_05037_),
    .A_N(\game_logic_inst.lfsr_value[14] ));
 sg13g2_and2_1 _10564_ (.A(net278),
    .B(\game_logic_inst.lfsr_value[15] ),
    .X(_00370_));
 sg13g2_buf_1 _10565_ (.A(net403),
    .X(_05038_));
 sg13g2_and2_1 _10566_ (.A(net263),
    .B(\lfsr_inst.lfsr[16] ),
    .X(_00371_));
 sg13g2_and2_1 _10567_ (.A(net263),
    .B(\lfsr_inst.lfsr[17] ),
    .X(_00372_));
 sg13g2_nand2b_1 _10568_ (.Y(_00373_),
    .B(net264),
    .A_N(\lfsr_inst.lfsr[18] ));
 sg13g2_nand2b_1 _10569_ (.Y(_00374_),
    .B(_05037_),
    .A_N(\game_logic_inst.lfsr_value[0] ));
 sg13g2_and2_1 _10570_ (.A(_05038_),
    .B(\lfsr_inst.lfsr[19] ),
    .X(_00375_));
 sg13g2_and2_1 _10571_ (.A(net263),
    .B(\lfsr_inst.lfsr[20] ),
    .X(_00376_));
 sg13g2_nand2b_1 _10572_ (.Y(_00377_),
    .B(net264),
    .A_N(\lfsr_inst.lfsr[21] ));
 sg13g2_and2_1 _10573_ (.A(_05038_),
    .B(\lfsr_inst.lfsr[22] ),
    .X(_00378_));
 sg13g2_and2_1 _10574_ (.A(net263),
    .B(\lfsr_inst.lfsr[23] ),
    .X(_00379_));
 sg13g2_and2_1 _10575_ (.A(net263),
    .B(\lfsr_inst.lfsr[24] ),
    .X(_00380_));
 sg13g2_and2_1 _10576_ (.A(net263),
    .B(\lfsr_inst.lfsr[25] ),
    .X(_00381_));
 sg13g2_and2_1 _10577_ (.A(net263),
    .B(\lfsr_inst.lfsr[26] ),
    .X(_00382_));
 sg13g2_and2_1 _10578_ (.A(net263),
    .B(\lfsr_inst.lfsr[27] ),
    .X(_00383_));
 sg13g2_nand2b_1 _10579_ (.Y(_00384_),
    .B(net264),
    .A_N(_02003_));
 sg13g2_and2_1 _10580_ (.A(net343),
    .B(\game_logic_inst.lfsr_value[1] ),
    .X(_00385_));
 sg13g2_and2_1 _10581_ (.A(net343),
    .B(net466),
    .X(_00386_));
 sg13g2_and2_1 _10582_ (.A(net343),
    .B(net465),
    .X(_00387_));
 sg13g2_nand2b_1 _10583_ (.Y(_00388_),
    .B(net279),
    .A_N(\game_logic_inst.lfsr_value[2] ));
 sg13g2_nand2b_1 _10584_ (.Y(_00389_),
    .B(net279),
    .A_N(\game_logic_inst.lfsr_value[3] ));
 sg13g2_nand2b_1 _10585_ (.Y(_00390_),
    .B(net279),
    .A_N(\game_logic_inst.lfsr_value[4] ));
 sg13g2_nand2b_1 _10586_ (.Y(_00391_),
    .B(net279),
    .A_N(\game_logic_inst.lfsr_value[5] ));
 sg13g2_nand2b_1 _10587_ (.Y(_00392_),
    .B(net279),
    .A_N(\game_logic_inst.lfsr_value[6] ));
 sg13g2_and2_1 _10588_ (.A(_01864_),
    .B(\game_logic_inst.lfsr_value[7] ),
    .X(_00393_));
 sg13g2_nand2b_1 _10589_ (.Y(_00394_),
    .B(_04634_),
    .A_N(\game_logic_inst.lfsr_value[8] ));
 sg13g2_nor4_1 _10590_ (.A(_05070_),
    .B(_05065_),
    .C(_05073_),
    .D(_05066_),
    .Y(_05039_));
 sg13g2_o21ai_1 _10591_ (.B1(_04871_),
    .Y(_05040_),
    .A1(net395),
    .A2(_05039_));
 sg13g2_nand2_1 _10592_ (.Y(_00416_),
    .A(net264),
    .B(_05040_));
 sg13g2_and2_1 _10593_ (.A(_01864_),
    .B(\vga_sync_gen.vsync ),
    .X(_00437_));
 sg13g2_nand3b_1 _10594_ (.B(_04880_),
    .C(_02015_),
    .Y(_05041_),
    .A_N(_02001_));
 sg13g2_nand2_1 _10595_ (.Y(_05042_),
    .A(_02001_),
    .B(_01878_));
 sg13g2_a21oi_1 _10596_ (.A1(_05041_),
    .A2(_05042_),
    .Y(_00454_),
    .B1(net344));
 sg13g2_nand2_1 _10597_ (.Y(_05043_),
    .A(_02001_),
    .B(_01793_));
 sg13g2_o21ai_1 _10598_ (.B1(_01565_),
    .Y(_05044_),
    .A1(_02012_),
    .A2(_05043_));
 sg13g2_nand3b_1 _10599_ (.B(_05043_),
    .C(_02012_),
    .Y(_05045_),
    .A_N(_02016_));
 sg13g2_nand2b_1 _10600_ (.Y(_00455_),
    .B(_05045_),
    .A_N(_05044_));
 sg13g2_nand3_1 _10601_ (.B(_02001_),
    .C(_01793_),
    .A(_02012_),
    .Y(_05046_));
 sg13g2_o21ai_1 _10602_ (.B1(_01565_),
    .Y(_05047_),
    .A1(_02014_),
    .A2(_05046_));
 sg13g2_nand3b_1 _10603_ (.B(_05046_),
    .C(_02014_),
    .Y(_05048_),
    .A_N(_02016_));
 sg13g2_nand2b_1 _10604_ (.Y(_00456_),
    .B(_05048_),
    .A_N(_05047_));
 sg13g2_nand4_1 _10605_ (.B(_02001_),
    .C(_02014_),
    .A(_02012_),
    .Y(_05049_),
    .D(_01793_));
 sg13g2_buf_1 _10606_ (.A(_05049_),
    .X(_05050_));
 sg13g2_o21ai_1 _10607_ (.B1(_01367_),
    .Y(_05051_),
    .A1(_02013_),
    .A2(_05050_));
 sg13g2_nand3b_1 _10608_ (.B(_05050_),
    .C(_02013_),
    .Y(_05052_),
    .A_N(_02016_));
 sg13g2_nand2b_1 _10609_ (.Y(_00457_),
    .B(_05052_),
    .A_N(_05051_));
 sg13g2_inv_1 _10610_ (.Y(_05053_),
    .A(_05050_));
 sg13g2_o21ai_1 _10611_ (.B1(_02013_),
    .Y(_05054_),
    .A1(_02016_),
    .A2(_05053_));
 sg13g2_nand2b_1 _10612_ (.Y(_05055_),
    .B(_02013_),
    .A_N(\welcome_screen_inst.welcome_counter[4] ));
 sg13g2_o21ai_1 _10613_ (.B1(_01367_),
    .Y(_05056_),
    .A1(_05050_),
    .A2(_05055_));
 sg13g2_a21o_1 _10614_ (.A2(_05054_),
    .A1(\welcome_screen_inst.welcome_counter[4] ),
    .B1(_05056_),
    .X(_00458_));
 sg13g2_buf_4 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_tiehi \B[0]$_SDFF_PN0__490  (.L_HI(net490));
 sg13g2_buf_1 _10617_ (.A(net482),
    .X(uio_oe[0]));
 sg13g2_buf_1 _10618_ (.A(net483),
    .X(uio_oe[1]));
 sg13g2_buf_1 _10619_ (.A(net484),
    .X(uio_oe[2]));
 sg13g2_buf_1 _10620_ (.A(net485),
    .X(uio_oe[3]));
 sg13g2_buf_1 _10621_ (.A(\debug_controller_inst.data_out_en ),
    .X(net14));
 sg13g2_buf_1 _10622_ (.A(\debug_controller_inst.data_out_en ),
    .X(net15));
 sg13g2_buf_1 _10623_ (.A(\debug_controller_inst.data_out_en ),
    .X(net16));
 sg13g2_buf_1 _10624_ (.A(\debug_controller_inst.data_out_en ),
    .X(net17));
 sg13g2_buf_1 _10625_ (.A(net486),
    .X(uio_out[0]));
 sg13g2_buf_1 _10626_ (.A(net487),
    .X(uio_out[1]));
 sg13g2_buf_1 _10627_ (.A(net488),
    .X(uio_out[2]));
 sg13g2_buf_1 _10628_ (.A(net489),
    .X(uio_out[3]));
 sg13g2_buf_1 _10629_ (.A(\vga_sync_gen.vsync ),
    .X(net25));
 sg13g2_buf_1 _10630_ (.A(hsync),
    .X(net29));
 sg13g2_dfrbp_1 \btn_down_debounce.button_sync_0$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net496),
    .D(_00177_),
    .Q_N(_05474_),
    .Q(\btn_down_debounce.button_sync_0 ));
 sg13g2_dfrbp_1 \btn_down_debounce.button_sync_1$_SDFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net497),
    .D(_00178_),
    .Q_N(_05473_),
    .Q(\btn_down_debounce.button_sync_1 ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[0]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net498),
    .D(_00179_),
    .Q_N(_00166_),
    .Q(\btn_down_debounce.debounce_counter[0] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[10]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net499),
    .D(_00180_),
    .Q_N(_05472_),
    .Q(\btn_down_debounce.debounce_counter[10] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[11]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net500),
    .D(_00181_),
    .Q_N(_05471_),
    .Q(\btn_down_debounce.debounce_counter[11] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[12]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net501),
    .D(_00182_),
    .Q_N(_05470_),
    .Q(\btn_down_debounce.debounce_counter[12] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[13]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net502),
    .D(_00183_),
    .Q_N(_05469_),
    .Q(\btn_down_debounce.debounce_counter[13] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[14]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net503),
    .D(_00184_),
    .Q_N(_05468_),
    .Q(\btn_down_debounce.debounce_counter[14] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[15]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net504),
    .D(_00185_),
    .Q_N(_05467_),
    .Q(\btn_down_debounce.debounce_counter[15] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[16]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net505),
    .D(_00186_),
    .Q_N(_05466_),
    .Q(\btn_down_debounce.debounce_counter[16] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[17]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net506),
    .D(_00187_),
    .Q_N(_05465_),
    .Q(\btn_down_debounce.debounce_counter[17] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[1]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net507),
    .D(_00188_),
    .Q_N(_05464_),
    .Q(\btn_down_debounce.debounce_counter[1] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[2]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net508),
    .D(_00189_),
    .Q_N(_05463_),
    .Q(\btn_down_debounce.debounce_counter[2] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[3]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net509),
    .D(_00190_),
    .Q_N(_05462_),
    .Q(\btn_down_debounce.debounce_counter[3] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[4]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net510),
    .D(_00191_),
    .Q_N(_05461_),
    .Q(\btn_down_debounce.debounce_counter[4] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[5]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net511),
    .D(_00192_),
    .Q_N(_05460_),
    .Q(\btn_down_debounce.debounce_counter[5] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[6]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net512),
    .D(_00193_),
    .Q_N(_05459_),
    .Q(\btn_down_debounce.debounce_counter[6] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[7]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net513),
    .D(_00194_),
    .Q_N(_05458_),
    .Q(\btn_down_debounce.debounce_counter[7] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[8]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net514),
    .D(_00195_),
    .Q_N(_05457_),
    .Q(\btn_down_debounce.debounce_counter[8] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounce_counter[9]$_SDFF_PP0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net515),
    .D(_00196_),
    .Q_N(_05456_),
    .Q(\btn_down_debounce.debounce_counter[9] ));
 sg13g2_dfrbp_1 \btn_down_debounce.debounced$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net516),
    .D(_00197_),
    .Q_N(_05455_),
    .Q(btn_down));
 sg13g2_dfrbp_1 \btn_left_debounce.button_sync_0$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net517),
    .D(_00198_),
    .Q_N(_05454_),
    .Q(\btn_left_debounce.button_sync_0 ));
 sg13g2_dfrbp_1 \btn_left_debounce.button_sync_1$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net518),
    .D(_00199_),
    .Q_N(_05453_),
    .Q(\btn_left_debounce.button_sync_1 ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[0]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net519),
    .D(_00200_),
    .Q_N(_00167_),
    .Q(\btn_left_debounce.debounce_counter[0] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[10]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net520),
    .D(_00201_),
    .Q_N(_05452_),
    .Q(\btn_left_debounce.debounce_counter[10] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[11]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net521),
    .D(_00202_),
    .Q_N(_05451_),
    .Q(\btn_left_debounce.debounce_counter[11] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[12]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net522),
    .D(_00203_),
    .Q_N(_05450_),
    .Q(\btn_left_debounce.debounce_counter[12] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[13]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net523),
    .D(_00204_),
    .Q_N(_05449_),
    .Q(\btn_left_debounce.debounce_counter[13] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[14]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net524),
    .D(_00205_),
    .Q_N(_05448_),
    .Q(\btn_left_debounce.debounce_counter[14] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[15]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net525),
    .D(_00206_),
    .Q_N(_05447_),
    .Q(\btn_left_debounce.debounce_counter[15] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[16]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net526),
    .D(_00207_),
    .Q_N(_05446_),
    .Q(\btn_left_debounce.debounce_counter[16] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[17]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net527),
    .D(_00208_),
    .Q_N(_05445_),
    .Q(\btn_left_debounce.debounce_counter[17] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[1]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net528),
    .D(_00209_),
    .Q_N(_05444_),
    .Q(\btn_left_debounce.debounce_counter[1] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[2]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net529),
    .D(_00210_),
    .Q_N(_05443_),
    .Q(\btn_left_debounce.debounce_counter[2] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[3]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net530),
    .D(_00211_),
    .Q_N(_05442_),
    .Q(\btn_left_debounce.debounce_counter[3] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[4]$_SDFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net531),
    .D(_00212_),
    .Q_N(_05441_),
    .Q(\btn_left_debounce.debounce_counter[4] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[5]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net532),
    .D(_00213_),
    .Q_N(_05440_),
    .Q(\btn_left_debounce.debounce_counter[5] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[6]$_SDFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net533),
    .D(_00214_),
    .Q_N(_05439_),
    .Q(\btn_left_debounce.debounce_counter[6] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[7]$_SDFF_PP0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net534),
    .D(_00215_),
    .Q_N(_05438_),
    .Q(\btn_left_debounce.debounce_counter[7] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[8]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net535),
    .D(_00216_),
    .Q_N(_05437_),
    .Q(\btn_left_debounce.debounce_counter[8] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounce_counter[9]$_SDFF_PP0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net536),
    .D(_00217_),
    .Q_N(_05436_),
    .Q(\btn_left_debounce.debounce_counter[9] ));
 sg13g2_dfrbp_1 \btn_left_debounce.debounced$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net537),
    .D(_00218_),
    .Q_N(_05435_),
    .Q(btn_left));
 sg13g2_dfrbp_1 \btn_right_debounce.button_sync_0$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net538),
    .D(_00219_),
    .Q_N(_05434_),
    .Q(\btn_right_debounce.button_sync_0 ));
 sg13g2_dfrbp_1 \btn_right_debounce.button_sync_1$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net539),
    .D(_00220_),
    .Q_N(_05433_),
    .Q(\btn_right_debounce.button_sync_1 ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[0]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net540),
    .D(_00221_),
    .Q_N(_00168_),
    .Q(\btn_right_debounce.debounce_counter[0] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[10]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net541),
    .D(_00222_),
    .Q_N(_05432_),
    .Q(\btn_right_debounce.debounce_counter[10] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[11]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net542),
    .D(_00223_),
    .Q_N(_05431_),
    .Q(\btn_right_debounce.debounce_counter[11] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[12]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net543),
    .D(_00224_),
    .Q_N(_05430_),
    .Q(\btn_right_debounce.debounce_counter[12] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[13]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net544),
    .D(_00225_),
    .Q_N(_05429_),
    .Q(\btn_right_debounce.debounce_counter[13] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[14]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net545),
    .D(_00226_),
    .Q_N(_05428_),
    .Q(\btn_right_debounce.debounce_counter[14] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[15]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net546),
    .D(_00227_),
    .Q_N(_05427_),
    .Q(\btn_right_debounce.debounce_counter[15] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[16]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net547),
    .D(_00228_),
    .Q_N(_05426_),
    .Q(\btn_right_debounce.debounce_counter[16] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[17]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net548),
    .D(_00229_),
    .Q_N(_05425_),
    .Q(\btn_right_debounce.debounce_counter[17] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[1]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net549),
    .D(_00230_),
    .Q_N(_05424_),
    .Q(\btn_right_debounce.debounce_counter[1] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[2]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net550),
    .D(_00231_),
    .Q_N(_05423_),
    .Q(\btn_right_debounce.debounce_counter[2] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[3]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net551),
    .D(_00232_),
    .Q_N(_05422_),
    .Q(\btn_right_debounce.debounce_counter[3] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[4]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net552),
    .D(_00233_),
    .Q_N(_05421_),
    .Q(\btn_right_debounce.debounce_counter[4] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[5]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net553),
    .D(_00234_),
    .Q_N(_05420_),
    .Q(\btn_right_debounce.debounce_counter[5] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[6]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net554),
    .D(_00235_),
    .Q_N(_05419_),
    .Q(\btn_right_debounce.debounce_counter[6] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[7]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net555),
    .D(_00236_),
    .Q_N(_05418_),
    .Q(\btn_right_debounce.debounce_counter[7] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[8]$_SDFF_PP0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net556),
    .D(_00237_),
    .Q_N(_05417_),
    .Q(\btn_right_debounce.debounce_counter[8] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounce_counter[9]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net557),
    .D(_00238_),
    .Q_N(_05416_),
    .Q(\btn_right_debounce.debounce_counter[9] ));
 sg13g2_dfrbp_1 \btn_right_debounce.debounced$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net558),
    .D(_00239_),
    .Q_N(_05415_),
    .Q(btn_right));
 sg13g2_dfrbp_1 \btn_up_debounce.button_sync_0$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net559),
    .D(_00240_),
    .Q_N(_05414_),
    .Q(\btn_up_debounce.button_sync_0 ));
 sg13g2_dfrbp_1 \btn_up_debounce.button_sync_1$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net560),
    .D(_00241_),
    .Q_N(_05413_),
    .Q(\btn_up_debounce.button_sync_1 ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[0]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net561),
    .D(_00242_),
    .Q_N(_00169_),
    .Q(\btn_up_debounce.debounce_counter[0] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[10]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net562),
    .D(_00243_),
    .Q_N(_05412_),
    .Q(\btn_up_debounce.debounce_counter[10] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[11]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net563),
    .D(_00244_),
    .Q_N(_05411_),
    .Q(\btn_up_debounce.debounce_counter[11] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[12]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net564),
    .D(_00245_),
    .Q_N(_05410_),
    .Q(\btn_up_debounce.debounce_counter[12] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[13]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net565),
    .D(_00246_),
    .Q_N(_05409_),
    .Q(\btn_up_debounce.debounce_counter[13] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[14]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net566),
    .D(_00247_),
    .Q_N(_05408_),
    .Q(\btn_up_debounce.debounce_counter[14] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[15]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net567),
    .D(_00248_),
    .Q_N(_05407_),
    .Q(\btn_up_debounce.debounce_counter[15] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[16]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net568),
    .D(_00249_),
    .Q_N(_05406_),
    .Q(\btn_up_debounce.debounce_counter[16] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[17]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net569),
    .D(_00250_),
    .Q_N(_05405_),
    .Q(\btn_up_debounce.debounce_counter[17] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[1]$_SDFF_PP0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net570),
    .D(_00251_),
    .Q_N(_05404_),
    .Q(\btn_up_debounce.debounce_counter[1] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[2]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net571),
    .D(_00252_),
    .Q_N(_05403_),
    .Q(\btn_up_debounce.debounce_counter[2] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[3]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net572),
    .D(_00253_),
    .Q_N(_05402_),
    .Q(\btn_up_debounce.debounce_counter[3] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[4]$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net573),
    .D(_00254_),
    .Q_N(_05401_),
    .Q(\btn_up_debounce.debounce_counter[4] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[5]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net574),
    .D(_00255_),
    .Q_N(_05400_),
    .Q(\btn_up_debounce.debounce_counter[5] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[6]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net575),
    .D(_00256_),
    .Q_N(_05399_),
    .Q(\btn_up_debounce.debounce_counter[6] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[7]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net576),
    .D(_00257_),
    .Q_N(_05398_),
    .Q(\btn_up_debounce.debounce_counter[7] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[8]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net577),
    .D(_00258_),
    .Q_N(_05397_),
    .Q(\btn_up_debounce.debounce_counter[8] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounce_counter[9]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net578),
    .D(_00259_),
    .Q_N(_05396_),
    .Q(\btn_up_debounce.debounce_counter[9] ));
 sg13g2_dfrbp_1 \btn_up_debounce.debounced$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net579),
    .D(_00260_),
    .Q_N(_05395_),
    .Q(btn_up));
 sg13g2_dfrbp_1 \debug_controller_inst.data_out[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net580),
    .D(_00261_),
    .Q_N(_05394_),
    .Q(net18));
 sg13g2_dfrbp_1 \debug_controller_inst.data_out[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net581),
    .D(_00262_),
    .Q_N(_05393_),
    .Q(net19));
 sg13g2_dfrbp_1 \debug_controller_inst.data_out[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net582),
    .D(_00263_),
    .Q_N(_05392_),
    .Q(net20));
 sg13g2_dfrbp_1 \debug_controller_inst.data_out[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net583),
    .D(_00264_),
    .Q_N(_05391_),
    .Q(net21));
 sg13g2_dfrbp_1 \debug_controller_inst.data_out_en$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net584),
    .D(_00265_),
    .Q_N(_05390_),
    .Q(\debug_controller_inst.data_out_en ));
 sg13g2_dfrbp_1 \debug_controller_inst.force_move[0]$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net585),
    .D(_00266_),
    .Q_N(_05389_),
    .Q(debug_btn_up));
 sg13g2_dfrbp_1 \debug_controller_inst.force_move[1]$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net586),
    .D(_00267_),
    .Q_N(_05388_),
    .Q(debug_btn_down));
 sg13g2_dfrbp_1 \debug_controller_inst.force_move[2]$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net587),
    .D(_00268_),
    .Q_N(_05387_),
    .Q(debug_btn_left));
 sg13g2_dfrbp_1 \debug_controller_inst.force_move[3]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net588),
    .D(_00269_),
    .Q_N(_05386_),
    .Q(debug_btn_right));
 sg13g2_dfrbp_1 \debug_controller_inst.grid_addr[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net589),
    .D(_00270_),
    .Q_N(_00088_),
    .Q(\debug_controller_inst.grid_addr[0] ));
 sg13g2_dfrbp_1 \debug_controller_inst.grid_addr[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net590),
    .D(_00271_),
    .Q_N(_05385_),
    .Q(\debug_controller_inst.grid_addr[1] ));
 sg13g2_dfrbp_1 \debug_controller_inst.grid_addr[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net591),
    .D(_00272_),
    .Q_N(_05384_),
    .Q(\debug_controller_inst.grid_addr[2] ));
 sg13g2_dfrbp_1 \debug_controller_inst.grid_addr[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net592),
    .D(_00273_),
    .Q_N(_05383_),
    .Q(\debug_controller_inst.grid_addr[3] ));
 sg13g2_dfrbp_1 \debug_controller_inst.grid_out_addr[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net593),
    .D(_00274_),
    .Q_N(_00099_),
    .Q(\debug_controller_inst.grid_out_addr[0] ));
 sg13g2_dfrbp_1 \debug_controller_inst.grid_out_addr[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net594),
    .D(_00275_),
    .Q_N(_05382_),
    .Q(\debug_controller_inst.grid_out_addr[1] ));
 sg13g2_dfrbp_1 \debug_controller_inst.grid_out_addr[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net595),
    .D(_00276_),
    .Q_N(_05381_),
    .Q(\debug_controller_inst.grid_out_addr[2] ));
 sg13g2_dfrbp_1 \debug_controller_inst.grid_out_addr[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net596),
    .D(_00277_),
    .Q_N(_05380_),
    .Q(\debug_controller_inst.grid_out_addr[3] ));
 sg13g2_dfrbp_1 \debug_controller_inst.grid_out_data[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net597),
    .D(_00278_),
    .Q_N(_05379_),
    .Q(\debug_controller_inst.grid_out_data[0] ));
 sg13g2_dfrbp_1 \debug_controller_inst.grid_out_data[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net598),
    .D(_00279_),
    .Q_N(_05378_),
    .Q(\debug_controller_inst.grid_out_data[1] ));
 sg13g2_dfrbp_1 \debug_controller_inst.grid_out_data[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net599),
    .D(_00280_),
    .Q_N(_05377_),
    .Q(\debug_controller_inst.grid_out_data[2] ));
 sg13g2_dfrbp_1 \debug_controller_inst.grid_out_data[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net600),
    .D(_00281_),
    .Q_N(_05376_),
    .Q(\debug_controller_inst.grid_out_data[3] ));
 sg13g2_dfrbp_1 \debug_controller_inst.grid_out_valid$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net601),
    .D(_00282_),
    .Q_N(_05375_),
    .Q(\debug_controller_inst.grid_out_valid ));
 sg13g2_dfrbp_1 \game_logic_inst.add_new_tiles[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net602),
    .D(_00283_),
    .Q_N(_05374_),
    .Q(\game_logic_inst.add_new_tiles[0] ));
 sg13g2_dfrbp_1 \game_logic_inst.add_new_tiles[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net603),
    .D(_00284_),
    .Q_N(_05373_),
    .Q(\game_logic_inst.add_new_tiles[1] ));
 sg13g2_dfrbp_1 \game_logic_inst.added_tile_index[0]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net604),
    .D(_00285_),
    .Q_N(_05372_),
    .Q(\game_logic_inst.added_tile_index[0] ));
 sg13g2_dfrbp_1 \game_logic_inst.added_tile_index[1]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net605),
    .D(_00286_),
    .Q_N(_05371_),
    .Q(\game_logic_inst.added_tile_index[1] ));
 sg13g2_dfrbp_1 \game_logic_inst.added_tile_index[2]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net606),
    .D(_00287_),
    .Q_N(_05370_),
    .Q(\game_logic_inst.added_tile_index[2] ));
 sg13g2_dfrbp_1 \game_logic_inst.added_tile_index[3]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net607),
    .D(_00288_),
    .Q_N(_05369_),
    .Q(\game_logic_inst.added_tile_index[3] ));
 sg13g2_dfrbp_1 \game_logic_inst.calculate_move$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net608),
    .D(_00289_),
    .Q_N(_00069_),
    .Q(\game_logic_inst.calculate_move ));
 sg13g2_dfrbp_1 \game_logic_inst.current_direction[1]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net609),
    .D(_00000_),
    .Q_N(_05481_),
    .Q(\game_logic_inst.current_direction[1] ));
 sg13g2_dfrbp_1 \game_logic_inst.current_direction[2]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net610),
    .D(_00001_),
    .Q_N(_05482_),
    .Q(\game_logic_inst.current_direction[2] ));
 sg13g2_dfrbp_1 \game_logic_inst.current_direction[3]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net611),
    .D(_00002_),
    .Q_N(_05368_),
    .Q(\game_logic_inst.current_direction[3] ));
 sg13g2_dfrbp_1 \game_logic_inst.current_row_index[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net612),
    .D(_00290_),
    .Q_N(_00097_),
    .Q(\game_logic_inst.current_row_index[0] ));
 sg13g2_dfrbp_1 \game_logic_inst.current_row_index[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net613),
    .D(_00291_),
    .Q_N(_05367_),
    .Q(\game_logic_inst.current_row_index[1] ));
 sg13g2_dfrbp_1 \game_logic_inst.debug_move_reg$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net614),
    .D(_00292_),
    .Q_N(_05366_),
    .Q(\game_logic_inst.debug_move_reg ));
 sg13g2_dfrbp_1 \game_logic_inst.game_started$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net615),
    .D(_00293_),
    .Q_N(_00163_),
    .Q(\game_logic_inst.game_started ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[0]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net616),
    .D(_00003_),
    .Q_N(_00098_),
    .Q(\debug_controller_inst.grid_in[0] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[10]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net617),
    .D(_00004_),
    .Q_N(_00115_),
    .Q(\debug_controller_inst.grid_in[10] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[11]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net618),
    .D(_00005_),
    .Q_N(_00117_),
    .Q(\debug_controller_inst.grid_in[11] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[12]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net619),
    .D(_00006_),
    .Q_N(_00119_),
    .Q(\debug_controller_inst.grid_in[12] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[13]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net620),
    .D(_00007_),
    .Q_N(_00121_),
    .Q(\debug_controller_inst.grid_in[13] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[14]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net621),
    .D(_00008_),
    .Q_N(_00123_),
    .Q(\debug_controller_inst.grid_in[14] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[15]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net622),
    .D(_00009_),
    .Q_N(_00125_),
    .Q(\debug_controller_inst.grid_in[15] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[16]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net623),
    .D(_00010_),
    .Q_N(_00104_),
    .Q(\debug_controller_inst.grid_in[16] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[17]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net624),
    .D(_00011_),
    .Q_N(_00106_),
    .Q(\debug_controller_inst.grid_in[17] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[18]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net625),
    .D(_00012_),
    .Q_N(_00108_),
    .Q(\debug_controller_inst.grid_in[18] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[19]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net626),
    .D(_00013_),
    .Q_N(_00110_),
    .Q(\debug_controller_inst.grid_in[19] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[1]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net627),
    .D(_00014_),
    .Q_N(_00100_),
    .Q(\debug_controller_inst.grid_in[1] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[20]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net628),
    .D(_00015_),
    .Q_N(_00127_),
    .Q(\debug_controller_inst.grid_in[20] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[21]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net629),
    .D(_00016_),
    .Q_N(_00128_),
    .Q(\debug_controller_inst.grid_in[21] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[22]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net630),
    .D(_00017_),
    .Q_N(_00129_),
    .Q(\debug_controller_inst.grid_in[22] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[23]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net631),
    .D(_00018_),
    .Q_N(_00130_),
    .Q(\debug_controller_inst.grid_in[23] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[24]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net632),
    .D(_00019_),
    .Q_N(_00131_),
    .Q(\debug_controller_inst.grid_in[24] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[25]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net633),
    .D(_00020_),
    .Q_N(_00133_),
    .Q(\debug_controller_inst.grid_in[25] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[26]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net634),
    .D(_00021_),
    .Q_N(_00135_),
    .Q(\debug_controller_inst.grid_in[26] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[27]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net635),
    .D(_00022_),
    .Q_N(_00137_),
    .Q(\debug_controller_inst.grid_in[27] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[28]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net636),
    .D(_00023_),
    .Q_N(_00139_),
    .Q(\debug_controller_inst.grid_in[28] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[29]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net637),
    .D(_00024_),
    .Q_N(_00141_),
    .Q(\debug_controller_inst.grid_in[29] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[2]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net638),
    .D(_00025_),
    .Q_N(_00101_),
    .Q(\debug_controller_inst.grid_in[2] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[30]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net639),
    .D(_00026_),
    .Q_N(_00143_),
    .Q(\debug_controller_inst.grid_in[30] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[31]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net640),
    .D(_00027_),
    .Q_N(_00145_),
    .Q(\debug_controller_inst.grid_in[31] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[32]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net641),
    .D(_00028_),
    .Q_N(_00112_),
    .Q(\debug_controller_inst.grid_in[32] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[33]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net642),
    .D(_00029_),
    .Q_N(_00114_),
    .Q(\debug_controller_inst.grid_in[33] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[34]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net643),
    .D(_00030_),
    .Q_N(_00116_),
    .Q(\debug_controller_inst.grid_in[34] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[35]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net644),
    .D(_00031_),
    .Q_N(_00118_),
    .Q(\debug_controller_inst.grid_in[35] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[36]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net645),
    .D(_00032_),
    .Q_N(_00132_),
    .Q(\debug_controller_inst.grid_in[36] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[37]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net646),
    .D(_00033_),
    .Q_N(_00134_),
    .Q(\debug_controller_inst.grid_in[37] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[38]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net647),
    .D(_00034_),
    .Q_N(_00136_),
    .Q(\debug_controller_inst.grid_in[38] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[39]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net648),
    .D(_00035_),
    .Q_N(_00138_),
    .Q(\debug_controller_inst.grid_in[39] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[3]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net649),
    .D(_00036_),
    .Q_N(_00102_),
    .Q(\debug_controller_inst.grid_in[3] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[40]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net650),
    .D(_00037_),
    .Q_N(_00147_),
    .Q(\debug_controller_inst.grid_in[40] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[41]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net651),
    .D(_00038_),
    .Q_N(_00148_),
    .Q(\debug_controller_inst.grid_in[41] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[42]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net652),
    .D(_00039_),
    .Q_N(_00149_),
    .Q(\debug_controller_inst.grid_in[42] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[43]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net653),
    .D(_00040_),
    .Q_N(_00150_),
    .Q(\debug_controller_inst.grid_in[43] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[44]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net654),
    .D(_00041_),
    .Q_N(_00151_),
    .Q(\debug_controller_inst.grid_in[44] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[45]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net655),
    .D(_00042_),
    .Q_N(_00153_),
    .Q(\debug_controller_inst.grid_in[45] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[46]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net656),
    .D(_00043_),
    .Q_N(_00155_),
    .Q(\debug_controller_inst.grid_in[46] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[47]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net657),
    .D(_00044_),
    .Q_N(_00157_),
    .Q(\debug_controller_inst.grid_in[47] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[48]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net658),
    .D(_00045_),
    .Q_N(_00120_),
    .Q(\debug_controller_inst.grid_in[48] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[49]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net659),
    .D(_00046_),
    .Q_N(_00122_),
    .Q(\debug_controller_inst.grid_in[49] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[4]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net660),
    .D(_00047_),
    .Q_N(_00103_),
    .Q(\debug_controller_inst.grid_in[4] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[50]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net661),
    .D(_00048_),
    .Q_N(_00124_),
    .Q(\debug_controller_inst.grid_in[50] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[51]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net662),
    .D(_00049_),
    .Q_N(_00126_),
    .Q(\debug_controller_inst.grid_in[51] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[52]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net663),
    .D(_00050_),
    .Q_N(_00140_),
    .Q(\debug_controller_inst.grid_in[52] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[53]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net664),
    .D(_00051_),
    .Q_N(_00142_),
    .Q(\debug_controller_inst.grid_in[53] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[54]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net665),
    .D(_00052_),
    .Q_N(_00144_),
    .Q(\debug_controller_inst.grid_in[54] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[55]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net666),
    .D(_00053_),
    .Q_N(_00146_),
    .Q(\debug_controller_inst.grid_in[55] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[56]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net667),
    .D(_00054_),
    .Q_N(_00152_),
    .Q(\debug_controller_inst.grid_in[56] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[57]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net668),
    .D(_00055_),
    .Q_N(_00154_),
    .Q(\debug_controller_inst.grid_in[57] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[58]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net669),
    .D(_00056_),
    .Q_N(_00156_),
    .Q(\debug_controller_inst.grid_in[58] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[59]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net670),
    .D(_00057_),
    .Q_N(_00158_),
    .Q(\debug_controller_inst.grid_in[59] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[5]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net671),
    .D(_00058_),
    .Q_N(_00105_),
    .Q(\debug_controller_inst.grid_in[5] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[60]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net672),
    .D(_00059_),
    .Q_N(_00159_),
    .Q(\debug_controller_inst.grid_in[60] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[61]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net673),
    .D(_00060_),
    .Q_N(_00160_),
    .Q(\debug_controller_inst.grid_in[61] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[62]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net674),
    .D(_00061_),
    .Q_N(_00161_),
    .Q(\debug_controller_inst.grid_in[62] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[63]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net675),
    .D(_00062_),
    .Q_N(_00162_),
    .Q(\debug_controller_inst.grid_in[63] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[6]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net676),
    .D(_00063_),
    .Q_N(_00107_),
    .Q(\debug_controller_inst.grid_in[6] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[7]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net677),
    .D(_00064_),
    .Q_N(_00109_),
    .Q(\debug_controller_inst.grid_in[7] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[8]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net678),
    .D(_00065_),
    .Q_N(_00111_),
    .Q(\debug_controller_inst.grid_in[8] ));
 sg13g2_dfrbp_1 \game_logic_inst.grid[9]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net679),
    .D(_00066_),
    .Q_N(_00113_),
    .Q(\debug_controller_inst.grid_in[9] ));
 sg13g2_dfrbp_1 \game_logic_inst.lfsr_shift[0]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net680),
    .D(_00294_),
    .Q_N(_00170_),
    .Q(\game_logic_inst.lfsr_shift[0] ));
 sg13g2_dfrbp_1 \game_logic_inst.lfsr_shift[1]$_SDFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net681),
    .D(_00295_),
    .Q_N(_05365_),
    .Q(\game_logic_inst.lfsr_shift[1] ));
 sg13g2_dfrbp_1 \game_logic_inst.prev_any_button_pressed$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net682),
    .D(_00296_),
    .Q_N(_05364_),
    .Q(\game_logic_inst.prev_any_button_pressed ));
 sg13g2_dfrbp_1 \game_logic_inst.should_transpose$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net683),
    .D(_00297_),
    .Q_N(_05363_),
    .Q(\game_logic_inst.should_transpose ));
 sg13g2_dfrbp_1 \game_logic_inst.valid_move$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net684),
    .D(_00298_),
    .Q_N(_05362_),
    .Q(\game_logic_inst.valid_move ));
 sg13g2_dfrbp_1 \grid[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net685),
    .D(_00299_),
    .Q_N(_05361_),
    .Q(\draw_game_inst.grid[0] ));
 sg13g2_dfrbp_1 \grid[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net686),
    .D(_00300_),
    .Q_N(_05360_),
    .Q(\draw_game_inst.grid[10] ));
 sg13g2_dfrbp_1 \grid[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net687),
    .D(_00301_),
    .Q_N(_05359_),
    .Q(\draw_game_inst.grid[11] ));
 sg13g2_dfrbp_1 \grid[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net688),
    .D(_00302_),
    .Q_N(_05358_),
    .Q(\draw_game_inst.grid[12] ));
 sg13g2_dfrbp_1 \grid[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net689),
    .D(_00303_),
    .Q_N(_05357_),
    .Q(\draw_game_inst.grid[13] ));
 sg13g2_dfrbp_1 \grid[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net690),
    .D(_00304_),
    .Q_N(_05356_),
    .Q(\draw_game_inst.grid[14] ));
 sg13g2_dfrbp_1 \grid[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net691),
    .D(_00305_),
    .Q_N(_05355_),
    .Q(\draw_game_inst.grid[15] ));
 sg13g2_dfrbp_1 \grid[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net692),
    .D(_00306_),
    .Q_N(_05354_),
    .Q(\draw_game_inst.grid[16] ));
 sg13g2_dfrbp_1 \grid[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net693),
    .D(_00307_),
    .Q_N(_05353_),
    .Q(\draw_game_inst.grid[17] ));
 sg13g2_dfrbp_1 \grid[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net694),
    .D(_00308_),
    .Q_N(_05352_),
    .Q(\draw_game_inst.grid[18] ));
 sg13g2_dfrbp_1 \grid[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net695),
    .D(_00309_),
    .Q_N(_05351_),
    .Q(\draw_game_inst.grid[19] ));
 sg13g2_dfrbp_1 \grid[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net696),
    .D(_00310_),
    .Q_N(_05350_),
    .Q(\draw_game_inst.grid[1] ));
 sg13g2_dfrbp_1 \grid[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net697),
    .D(_00311_),
    .Q_N(_05349_),
    .Q(\draw_game_inst.grid[20] ));
 sg13g2_dfrbp_1 \grid[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net698),
    .D(_00312_),
    .Q_N(_05348_),
    .Q(\draw_game_inst.grid[21] ));
 sg13g2_dfrbp_1 \grid[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net699),
    .D(_00313_),
    .Q_N(_05347_),
    .Q(\draw_game_inst.grid[22] ));
 sg13g2_dfrbp_1 \grid[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net700),
    .D(_00314_),
    .Q_N(_05346_),
    .Q(\draw_game_inst.grid[23] ));
 sg13g2_dfrbp_1 \grid[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net701),
    .D(_00315_),
    .Q_N(_05345_),
    .Q(\draw_game_inst.grid[24] ));
 sg13g2_dfrbp_1 \grid[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net702),
    .D(_00316_),
    .Q_N(_05344_),
    .Q(\draw_game_inst.grid[25] ));
 sg13g2_dfrbp_1 \grid[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net703),
    .D(_00317_),
    .Q_N(_05343_),
    .Q(\draw_game_inst.grid[26] ));
 sg13g2_dfrbp_1 \grid[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net704),
    .D(_00318_),
    .Q_N(_05342_),
    .Q(\draw_game_inst.grid[27] ));
 sg13g2_dfrbp_1 \grid[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net705),
    .D(_00319_),
    .Q_N(_05341_),
    .Q(\draw_game_inst.grid[28] ));
 sg13g2_dfrbp_1 \grid[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net706),
    .D(_00320_),
    .Q_N(_05340_),
    .Q(\draw_game_inst.grid[29] ));
 sg13g2_dfrbp_1 \grid[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net707),
    .D(_00321_),
    .Q_N(_05339_),
    .Q(\draw_game_inst.grid[2] ));
 sg13g2_dfrbp_1 \grid[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net708),
    .D(_00322_),
    .Q_N(_05338_),
    .Q(\draw_game_inst.grid[30] ));
 sg13g2_dfrbp_1 \grid[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net709),
    .D(_00323_),
    .Q_N(_05337_),
    .Q(\draw_game_inst.grid[31] ));
 sg13g2_dfrbp_1 \grid[32]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net710),
    .D(_00324_),
    .Q_N(_05336_),
    .Q(\draw_game_inst.grid[32] ));
 sg13g2_dfrbp_1 \grid[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net711),
    .D(_00325_),
    .Q_N(_05335_),
    .Q(\draw_game_inst.grid[33] ));
 sg13g2_dfrbp_1 \grid[34]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net712),
    .D(_00326_),
    .Q_N(_05334_),
    .Q(\draw_game_inst.grid[34] ));
 sg13g2_dfrbp_1 \grid[35]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net713),
    .D(_00327_),
    .Q_N(_05333_),
    .Q(\draw_game_inst.grid[35] ));
 sg13g2_dfrbp_1 \grid[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net714),
    .D(_00328_),
    .Q_N(_05332_),
    .Q(\draw_game_inst.grid[36] ));
 sg13g2_dfrbp_1 \grid[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net715),
    .D(_00329_),
    .Q_N(_05331_),
    .Q(\draw_game_inst.grid[37] ));
 sg13g2_dfrbp_1 \grid[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net716),
    .D(_00330_),
    .Q_N(_05330_),
    .Q(\draw_game_inst.grid[38] ));
 sg13g2_dfrbp_1 \grid[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net717),
    .D(_00331_),
    .Q_N(_05329_),
    .Q(\draw_game_inst.grid[39] ));
 sg13g2_dfrbp_1 \grid[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net718),
    .D(_00332_),
    .Q_N(_05328_),
    .Q(\draw_game_inst.grid[3] ));
 sg13g2_dfrbp_1 \grid[40]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net719),
    .D(_00333_),
    .Q_N(_05327_),
    .Q(\draw_game_inst.grid[40] ));
 sg13g2_dfrbp_1 \grid[41]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net720),
    .D(_00334_),
    .Q_N(_05326_),
    .Q(\draw_game_inst.grid[41] ));
 sg13g2_dfrbp_1 \grid[42]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net721),
    .D(_00335_),
    .Q_N(_05325_),
    .Q(\draw_game_inst.grid[42] ));
 sg13g2_dfrbp_1 \grid[43]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net722),
    .D(_00336_),
    .Q_N(_05324_),
    .Q(\draw_game_inst.grid[43] ));
 sg13g2_dfrbp_1 \grid[44]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net723),
    .D(_00337_),
    .Q_N(_05323_),
    .Q(\draw_game_inst.grid[44] ));
 sg13g2_dfrbp_1 \grid[45]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net724),
    .D(_00338_),
    .Q_N(_05322_),
    .Q(\draw_game_inst.grid[45] ));
 sg13g2_dfrbp_1 \grid[46]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net725),
    .D(_00339_),
    .Q_N(_05321_),
    .Q(\draw_game_inst.grid[46] ));
 sg13g2_dfrbp_1 \grid[47]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net726),
    .D(_00340_),
    .Q_N(_05320_),
    .Q(\draw_game_inst.grid[47] ));
 sg13g2_dfrbp_1 \grid[48]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net727),
    .D(_00341_),
    .Q_N(_05319_),
    .Q(\draw_game_inst.grid[48] ));
 sg13g2_dfrbp_1 \grid[49]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net728),
    .D(_00342_),
    .Q_N(_05318_),
    .Q(\draw_game_inst.grid[49] ));
 sg13g2_dfrbp_1 \grid[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net729),
    .D(_00343_),
    .Q_N(_05317_),
    .Q(\draw_game_inst.grid[4] ));
 sg13g2_dfrbp_1 \grid[50]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net730),
    .D(_00344_),
    .Q_N(_05316_),
    .Q(\draw_game_inst.grid[50] ));
 sg13g2_dfrbp_1 \grid[51]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net731),
    .D(_00345_),
    .Q_N(_05315_),
    .Q(\draw_game_inst.grid[51] ));
 sg13g2_dfrbp_1 \grid[52]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net732),
    .D(_00346_),
    .Q_N(_05314_),
    .Q(\draw_game_inst.grid[52] ));
 sg13g2_dfrbp_1 \grid[53]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net733),
    .D(_00347_),
    .Q_N(_05313_),
    .Q(\draw_game_inst.grid[53] ));
 sg13g2_dfrbp_1 \grid[54]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net734),
    .D(_00348_),
    .Q_N(_05312_),
    .Q(\draw_game_inst.grid[54] ));
 sg13g2_dfrbp_1 \grid[55]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net735),
    .D(_00349_),
    .Q_N(_05311_),
    .Q(\draw_game_inst.grid[55] ));
 sg13g2_dfrbp_1 \grid[56]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net736),
    .D(_00350_),
    .Q_N(_05310_),
    .Q(\draw_game_inst.grid[56] ));
 sg13g2_dfrbp_1 \grid[57]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net737),
    .D(_00351_),
    .Q_N(_05309_),
    .Q(\draw_game_inst.grid[57] ));
 sg13g2_dfrbp_1 \grid[58]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net738),
    .D(_00352_),
    .Q_N(_05308_),
    .Q(\draw_game_inst.grid[58] ));
 sg13g2_dfrbp_1 \grid[59]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net739),
    .D(_00353_),
    .Q_N(_05307_),
    .Q(\draw_game_inst.grid[59] ));
 sg13g2_dfrbp_1 \grid[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net740),
    .D(_00354_),
    .Q_N(_05306_),
    .Q(\draw_game_inst.grid[5] ));
 sg13g2_dfrbp_1 \grid[60]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net741),
    .D(_00355_),
    .Q_N(_05305_),
    .Q(\draw_game_inst.grid[60] ));
 sg13g2_dfrbp_1 \grid[61]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net742),
    .D(_00356_),
    .Q_N(_05304_),
    .Q(\draw_game_inst.grid[61] ));
 sg13g2_dfrbp_1 \grid[62]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net743),
    .D(_00357_),
    .Q_N(_05303_),
    .Q(\draw_game_inst.grid[62] ));
 sg13g2_dfrbp_1 \grid[63]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net744),
    .D(_00358_),
    .Q_N(_05302_),
    .Q(\draw_game_inst.grid[63] ));
 sg13g2_dfrbp_1 \grid[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net745),
    .D(_00359_),
    .Q_N(_05301_),
    .Q(\draw_game_inst.grid[6] ));
 sg13g2_dfrbp_1 \grid[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net746),
    .D(_00360_),
    .Q_N(_05300_),
    .Q(\draw_game_inst.grid[7] ));
 sg13g2_dfrbp_1 \grid[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net747),
    .D(_00361_),
    .Q_N(_05299_),
    .Q(\draw_game_inst.grid[8] ));
 sg13g2_dfrbp_1 \grid[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net748),
    .D(_00362_),
    .Q_N(_05298_),
    .Q(\draw_game_inst.grid[9] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[0]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net749),
    .D(_00363_),
    .Q_N(_05297_),
    .Q(\game_logic_inst.lfsr_value[0] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[10]$_SDFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net750),
    .D(_00364_),
    .Q_N(_05296_),
    .Q(\game_logic_inst.lfsr_value[10] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[11]$_SDFF_PN1_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net751),
    .D(_00365_),
    .Q_N(_05295_),
    .Q(\game_logic_inst.lfsr_value[11] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[12]$_SDFF_PN1_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net752),
    .D(_00366_),
    .Q_N(_05294_),
    .Q(\game_logic_inst.lfsr_value[12] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[13]$_SDFF_PN1_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net753),
    .D(_00367_),
    .Q_N(_05293_),
    .Q(\game_logic_inst.lfsr_value[13] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[14]$_SDFF_PN1_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net754),
    .D(_00368_),
    .Q_N(_05292_),
    .Q(\game_logic_inst.lfsr_value[14] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[15]$_SDFF_PN1_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net755),
    .D(_00369_),
    .Q_N(_05291_),
    .Q(\game_logic_inst.lfsr_value[15] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[16]$_SDFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net756),
    .D(_00370_),
    .Q_N(_05290_),
    .Q(\lfsr_inst.lfsr[16] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[17]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net757),
    .D(_00371_),
    .Q_N(_05289_),
    .Q(\lfsr_inst.lfsr[17] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[18]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net758),
    .D(_00372_),
    .Q_N(_05288_),
    .Q(\lfsr_inst.lfsr[18] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[19]$_SDFF_PN1_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net759),
    .D(_00373_),
    .Q_N(_05287_),
    .Q(\lfsr_inst.lfsr[19] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[1]$_SDFF_PN1_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net760),
    .D(_00374_),
    .Q_N(_05286_),
    .Q(\game_logic_inst.lfsr_value[1] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[20]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net761),
    .D(_00375_),
    .Q_N(_05285_),
    .Q(\lfsr_inst.lfsr[20] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[21]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net762),
    .D(_00376_),
    .Q_N(_05284_),
    .Q(\lfsr_inst.lfsr[21] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[22]$_SDFF_PN1_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net763),
    .D(_00377_),
    .Q_N(_05283_),
    .Q(\lfsr_inst.lfsr[22] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[23]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net764),
    .D(_00378_),
    .Q_N(_05282_),
    .Q(\lfsr_inst.lfsr[23] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[24]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net765),
    .D(_00379_),
    .Q_N(_05281_),
    .Q(\lfsr_inst.lfsr[24] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[25]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net766),
    .D(_00380_),
    .Q_N(_05280_),
    .Q(\lfsr_inst.lfsr[25] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[26]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net767),
    .D(_00381_),
    .Q_N(_05279_),
    .Q(\lfsr_inst.lfsr[26] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[27]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net768),
    .D(_00382_),
    .Q_N(_05278_),
    .Q(\lfsr_inst.lfsr[27] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[28]$_SDFF_PN0_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net769),
    .D(_00383_),
    .Q_N(_00070_),
    .Q(\lfsr_inst.lfsr[28] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[29]$_SDFF_PN1_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net770),
    .D(_00384_),
    .Q_N(_05277_),
    .Q(\lfsr_inst.lfsr[29] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[2]$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net771),
    .D(_00385_),
    .Q_N(_05276_),
    .Q(\game_logic_inst.lfsr_value[2] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[30]$_SDFF_PN0_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net772),
    .D(_00386_),
    .Q_N(_05275_),
    .Q(\lfsr_inst.lfsr[30] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[31]$_SDFF_PN0_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net773),
    .D(_00387_),
    .Q_N(_05274_),
    .Q(\lfsr_inst.lfsr[31] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[3]$_SDFF_PN1_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net774),
    .D(_00388_),
    .Q_N(_05273_),
    .Q(\game_logic_inst.lfsr_value[3] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[4]$_SDFF_PN1_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net775),
    .D(_00389_),
    .Q_N(_05272_),
    .Q(\game_logic_inst.lfsr_value[4] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[5]$_SDFF_PN1_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net776),
    .D(_00390_),
    .Q_N(_05271_),
    .Q(\game_logic_inst.lfsr_value[5] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[6]$_SDFF_PN1_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net777),
    .D(_00391_),
    .Q_N(_05270_),
    .Q(\game_logic_inst.lfsr_value[6] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[7]$_SDFF_PN1_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net778),
    .D(_00392_),
    .Q_N(_05269_),
    .Q(\game_logic_inst.lfsr_value[7] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[8]$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net779),
    .D(_00393_),
    .Q_N(_05268_),
    .Q(\game_logic_inst.lfsr_value[8] ));
 sg13g2_dfrbp_1 \lfsr_inst.lfsr[9]$_SDFF_PN1_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net780),
    .D(_00394_),
    .Q_N(_05267_),
    .Q(\game_logic_inst.lfsr_value[9] ));
 sg13g2_dfrbp_1 \new_tiles[0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net781),
    .D(_00395_),
    .Q_N(_05266_),
    .Q(\draw_game_inst.new_tiles[0] ));
 sg13g2_dfrbp_1 \new_tiles[10]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net782),
    .D(_00396_),
    .Q_N(_00080_),
    .Q(\draw_game_inst.new_tiles[10] ));
 sg13g2_dfrbp_1 \new_tiles[11]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net783),
    .D(_00397_),
    .Q_N(_00081_),
    .Q(\draw_game_inst.new_tiles[11] ));
 sg13g2_dfrbp_1 \new_tiles[12]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net784),
    .D(_00398_),
    .Q_N(_00082_),
    .Q(\draw_game_inst.new_tiles[12] ));
 sg13g2_dfrbp_1 \new_tiles[13]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net785),
    .D(_00399_),
    .Q_N(_00083_),
    .Q(\draw_game_inst.new_tiles[13] ));
 sg13g2_dfrbp_1 \new_tiles[14]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net786),
    .D(_00400_),
    .Q_N(_00084_),
    .Q(\draw_game_inst.new_tiles[14] ));
 sg13g2_dfrbp_1 \new_tiles[15]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net787),
    .D(_00401_),
    .Q_N(_00085_),
    .Q(\draw_game_inst.new_tiles[15] ));
 sg13g2_dfrbp_1 \new_tiles[1]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net788),
    .D(_00402_),
    .Q_N(_00071_),
    .Q(\draw_game_inst.new_tiles[1] ));
 sg13g2_dfrbp_1 \new_tiles[2]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net789),
    .D(_00403_),
    .Q_N(_00072_),
    .Q(\draw_game_inst.new_tiles[2] ));
 sg13g2_dfrbp_1 \new_tiles[3]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net790),
    .D(_00404_),
    .Q_N(_00073_),
    .Q(\draw_game_inst.new_tiles[3] ));
 sg13g2_dfrbp_1 \new_tiles[4]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net791),
    .D(_00405_),
    .Q_N(_00074_),
    .Q(\draw_game_inst.new_tiles[4] ));
 sg13g2_dfrbp_1 \new_tiles[5]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net792),
    .D(_00406_),
    .Q_N(_00075_),
    .Q(\draw_game_inst.new_tiles[5] ));
 sg13g2_dfrbp_1 \new_tiles[6]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net793),
    .D(_00407_),
    .Q_N(_00076_),
    .Q(\draw_game_inst.new_tiles[6] ));
 sg13g2_dfrbp_1 \new_tiles[7]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net794),
    .D(_00408_),
    .Q_N(_00077_),
    .Q(\draw_game_inst.new_tiles[7] ));
 sg13g2_dfrbp_1 \new_tiles[8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net795),
    .D(_00409_),
    .Q_N(_00078_),
    .Q(\draw_game_inst.new_tiles[8] ));
 sg13g2_dfrbp_1 \new_tiles[9]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net796),
    .D(_00410_),
    .Q_N(_00079_),
    .Q(\draw_game_inst.new_tiles[9] ));
 sg13g2_dfrbp_1 \new_tiles_counter[0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net797),
    .D(_00411_),
    .Q_N(_00086_),
    .Q(\new_tiles_counter[0] ));
 sg13g2_dfrbp_1 \new_tiles_counter[1]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net798),
    .D(_00412_),
    .Q_N(_00087_),
    .Q(\draw_game_inst.new_tiles_counter[0] ));
 sg13g2_dfrbp_1 \new_tiles_counter[2]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net799),
    .D(_00413_),
    .Q_N(_05265_),
    .Q(\draw_game_inst.new_tiles_counter[1] ));
 sg13g2_dfrbp_1 \new_tiles_counter[3]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net800),
    .D(_00414_),
    .Q_N(_05264_),
    .Q(\draw_game_inst.new_tiles_counter[2] ));
 sg13g2_dfrbp_1 \new_tiles_counter[4]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net801),
    .D(_00415_),
    .Q_N(_05263_),
    .Q(\new_tiles_counter[4] ));
 sg13g2_dfrbp_1 \show_welcome_screen$_SDFFE_PN1P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net802),
    .D(_00416_),
    .Q_N(_05262_),
    .Q(show_welcome_screen));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[0]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net803),
    .D(_00417_),
    .Q_N(_00165_),
    .Q(\draw_game_inst.board_x[0] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[1]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net804),
    .D(_00418_),
    .Q_N(_05261_),
    .Q(\draw_game_inst.board_x[1] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[2]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net805),
    .D(_00419_),
    .Q_N(_05260_),
    .Q(\draw_game_inst.board_x[2] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[3]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net806),
    .D(_00420_),
    .Q_N(_00095_),
    .Q(\draw_game_inst.board_x[3] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[4]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net807),
    .D(_00421_),
    .Q_N(_00096_),
    .Q(\draw_game_inst.board_x[4] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[5]$_SDFF_PP0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net808),
    .D(_00422_),
    .Q_N(_00094_),
    .Q(\draw_game_inst.board_x[5] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[6]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net809),
    .D(_00423_),
    .Q_N(_05259_),
    .Q(\draw_game_inst.x[6] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[7]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net810),
    .D(_00424_),
    .Q_N(_05258_),
    .Q(\draw_game_inst.x[7] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[8]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net811),
    .D(_00425_),
    .Q_N(_05257_),
    .Q(\draw_game_inst.x[8] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[9]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net812),
    .D(_00426_),
    .Q_N(_05483_),
    .Q(\draw_game_inst.x[9] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hsync$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net813),
    .D(_00067_),
    .Q_N(_05256_),
    .Q(hsync));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net814),
    .D(_00427_),
    .Q_N(_00164_),
    .Q(\draw_game_inst.board_y[0] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net815),
    .D(_00428_),
    .Q_N(_00093_),
    .Q(\draw_game_inst.board_y[1] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net816),
    .D(_00429_),
    .Q_N(_00092_),
    .Q(\draw_game_inst.board_y[2] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net817),
    .D(_00430_),
    .Q_N(_00091_),
    .Q(\draw_game_inst.board_y[3] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[4]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net818),
    .D(_00431_),
    .Q_N(_00090_),
    .Q(\draw_game_inst.board_y[4] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[5]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net819),
    .D(_00432_),
    .Q_N(_05255_),
    .Q(\draw_game_inst.board_y[5] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[6]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net820),
    .D(_00433_),
    .Q_N(_05254_),
    .Q(\draw_game_inst.board_y[6] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[7]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net821),
    .D(_00434_),
    .Q_N(_00089_),
    .Q(\draw_game_inst.y[7] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[8]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net822),
    .D(_00435_),
    .Q_N(_05253_),
    .Q(\draw_game_inst.y[8] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[9]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net823),
    .D(_00436_),
    .Q_N(_05484_),
    .Q(\draw_game_inst.y[9] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vsync$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net824),
    .D(_00068_),
    .Q_N(_05252_),
    .Q(\vga_sync_gen.vsync ));
 sg13g2_dfrbp_1 \vsync_prev$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net825),
    .D(_00437_),
    .Q_N(_05251_),
    .Q(vsync_prev));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[11]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net826),
    .D(_00438_),
    .Q_N(_05250_),
    .Q(\welcome_screen_grid[11] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[15]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net827),
    .D(_00439_),
    .Q_N(_05249_),
    .Q(\welcome_screen_grid[12] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[19]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net828),
    .D(_00440_),
    .Q_N(_05248_),
    .Q(\welcome_screen_grid[16] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[23]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net829),
    .D(_00441_),
    .Q_N(_05247_),
    .Q(\welcome_screen_grid[20] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[27]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net830),
    .D(_00442_),
    .Q_N(_05246_),
    .Q(\welcome_screen_grid[24] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[31]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net831),
    .D(_00443_),
    .Q_N(_05245_),
    .Q(\welcome_screen_grid[28] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[35]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net832),
    .D(_00444_),
    .Q_N(_05244_),
    .Q(\welcome_screen_grid[32] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[39]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net833),
    .D(_00445_),
    .Q_N(_05243_),
    .Q(\welcome_screen_grid[36] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net834),
    .D(_00446_),
    .Q_N(_05242_),
    .Q(\welcome_screen_grid[0] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[43]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net835),
    .D(_00447_),
    .Q_N(_05241_),
    .Q(\welcome_screen_grid[40] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[47]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net836),
    .D(_00448_),
    .Q_N(_05240_),
    .Q(\welcome_screen_grid[44] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[51]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net837),
    .D(_00449_),
    .Q_N(_05239_),
    .Q(\welcome_screen_grid[48] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[55]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net838),
    .D(_00450_),
    .Q_N(_05238_),
    .Q(\welcome_screen_grid[52] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[59]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net839),
    .D(_00451_),
    .Q_N(_05237_),
    .Q(\welcome_screen_grid[56] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[61]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net840),
    .D(_00452_),
    .Q_N(_05236_),
    .Q(\welcome_screen_grid[60] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.grid[7]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net841),
    .D(_00453_),
    .Q_N(_05235_),
    .Q(\welcome_screen_grid[4] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.welcome_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net842),
    .D(_00454_),
    .Q_N(_05234_),
    .Q(\welcome_screen_inst.welcome_counter[0] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.welcome_counter[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net843),
    .D(_00455_),
    .Q_N(_05233_),
    .Q(\welcome_screen_inst.welcome_counter[1] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.welcome_counter[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net844),
    .D(_00456_),
    .Q_N(_05232_),
    .Q(\welcome_screen_inst.welcome_counter[2] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.welcome_counter[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net845),
    .D(_00457_),
    .Q_N(_05231_),
    .Q(\welcome_screen_inst.welcome_counter[3] ));
 sg13g2_dfrbp_1 \welcome_screen_inst.welcome_counter[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net846),
    .D(_00458_),
    .Q_N(_05230_),
    .Q(\welcome_screen_inst.welcome_counter[4] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[0]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[5]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[6]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_oe[4]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[5]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_oe[6]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_oe[7]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[4]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[5]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[6]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[7]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[0]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[1]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[2]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[3]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[4]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[5]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[6]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout30 (.A(_01013_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_01036_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_00837_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_00747_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_00771_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_00661_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_00785_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_00654_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_01924_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_01240_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_00982_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_00813_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_00685_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_00682_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_00671_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_01233_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_00981_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_01304_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_01186_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_01119_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_00980_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_00765_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_00649_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_01118_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_00675_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_00667_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_00621_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_00563_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_03298_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_02920_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_02403_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_02069_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_02027_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_02020_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_02019_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_01624_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_01614_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_01471_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_01306_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_00949_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_00900_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_00602_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_00484_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_00477_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_05193_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_05115_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_03250_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_03161_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_03028_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_02992_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_02967_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_02944_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_02343_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_02238_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_02181_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_02124_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_02068_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_01964_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_01943_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_01919_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_01889_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_01812_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_00978_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_00936_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_05121_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_03314_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_03306_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_03299_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_03193_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_03142_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_03105_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_03052_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_03003_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_02994_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_02988_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_02983_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_02955_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_02939_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_02922_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_02916_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_02909_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_02903_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_02839_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_02818_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_02763_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_02761_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_02741_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_02737_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_02726_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_02718_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_02711_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_02706_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_02705_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_02681_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_02674_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_02645_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_02634_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_02628_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_02584_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_02565_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_02562_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_02533_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_02527_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_02519_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_02434_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_02423_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_02409_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_02390_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_02379_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_02370_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_02367_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_02357_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_02353_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_02342_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_02301_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_02291_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_02237_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_02180_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_02123_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_01963_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_01942_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_01938_),
    .X(net151));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(_01932_));
 sg13g2_buf_2 fanout153 (.A(_01918_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_01901_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_01888_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_01424_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_01287_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_00662_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_00568_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_05120_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_05113_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_03397_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_03350_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_03326_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_03305_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_03211_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_03190_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_03150_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_03086_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_03076_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_03023_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_03010_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_02928_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_02924_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_02901_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_02895_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_02889_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_02871_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_02852_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_02845_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_02824_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_02816_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_02810_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_02803_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_02801_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_02792_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_02788_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_02760_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_02752_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_02750_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_02745_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_02725_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_02720_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_02717_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_02714_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_02710_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_02708_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_02704_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_02693_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_02689_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_02686_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_02680_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_02672_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_02667_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_02651_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_02638_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_02633_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_02627_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_02626_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_02622_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_02583_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_02578_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_02568_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_02561_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_02555_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_02549_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_02537_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_02532_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_02526_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_02522_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_02518_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_02471_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_02466_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_02454_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_02452_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_02446_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_02439_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_02436_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_02433_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_02422_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_02413_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_02400_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_02389_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_02381_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_02378_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_02369_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_02366_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_02361_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_02356_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_02352_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_02341_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_02300_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_02297_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_02290_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_02286_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_01969_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_01962_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_01941_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_01937_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_01931_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_01917_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_01912_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_01900_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_01887_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_01504_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_01324_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_01247_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_01228_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_00482_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_05119_),
    .X(net260));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(_05112_));
 sg13g2_buf_2 fanout262 (.A(_05107_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_05038_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_05037_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_04991_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_04960_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_04950_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_04938_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_04923_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_04913_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_04889_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_04877_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_04875_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_04736_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_04719_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_04672_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_04639_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_04636_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_04634_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_03392_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_03020_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_02963_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_02923_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_02911_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_02900_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_02868_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_02867_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_02849_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_02842_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_02830_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_02791_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_02759_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_02756_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_02744_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_02712_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_02688_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_02679_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_02671_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_02666_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_02650_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_02637_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_02630_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_02629_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_02625_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_02621_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_02613_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_02607_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_02600_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_02585_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_02548_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_02538_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_02534_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_02531_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_02525_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_02520_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_02507_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_02470_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_02468_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_02460_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_02435_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_02425_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_02398_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_02368_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_02365_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_02360_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_02351_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_02344_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_02340_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_02336_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_02334_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_02332_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_02299_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_02289_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_02285_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_01971_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_01961_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_01949_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_01940_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_01936_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_01930_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_01911_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_01886_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_01864_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_01802_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_01789_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_01756_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_01398_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_01298_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_01286_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_01153_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_01089_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_01074_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_00987_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_05140_),
    .X(net354));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(_05139_));
 sg13g2_buf_4 fanout356 (.X(net356),
    .A(_05136_));
 sg13g2_buf_2 fanout357 (.A(_05118_),
    .X(net357));
 sg13g2_buf_4 fanout358 (.X(net358),
    .A(_05111_));
 sg13g2_buf_4 fanout359 (.X(net359),
    .A(_05106_));
 sg13g2_buf_2 fanout360 (.A(_05102_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_05061_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_04982_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_04980_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_04948_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_04911_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_04902_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_04892_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_04880_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_04879_),
    .X(net369));
 sg13g2_buf_1 fanout370 (.A(_04872_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_04870_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_02636_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_02619_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_02587_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_02506_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_02472_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_02450_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_02397_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_02382_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_02339_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_02335_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_02319_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_02298_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_02295_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_02284_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_01984_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_01967_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_01960_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_01955_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_01953_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_01952_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_01935_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_01929_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_01885_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_01878_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_01794_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_01780_),
    .X(net397));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(_01777_));
 sg13g2_buf_2 fanout399 (.A(_01769_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_01763_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_01755_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_01565_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_01367_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_01181_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_01120_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_00984_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_00919_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_05155_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_05117_),
    .X(net409));
 sg13g2_buf_4 fanout410 (.X(net410),
    .A(_05110_));
 sg13g2_buf_4 fanout411 (.X(net411),
    .A(_05105_));
 sg13g2_buf_2 fanout412 (.A(_05101_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_05060_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_04871_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_04869_),
    .X(net415));
 sg13g2_buf_4 fanout416 (.X(net416),
    .A(_04650_));
 sg13g2_buf_2 fanout417 (.A(_04647_),
    .X(net417));
 sg13g2_buf_4 fanout418 (.X(net418),
    .A(_04645_));
 sg13g2_buf_2 fanout419 (.A(_03139_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_02749_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_02660_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_02618_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_02586_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_02530_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_02513_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_02371_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_02348_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_02294_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_02283_),
    .X(net429));
 sg13g2_buf_4 fanout430 (.X(net430),
    .A(_02003_));
 sg13g2_buf_2 fanout431 (.A(_01959_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_01954_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_01926_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_01909_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_01897_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_01895_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_01884_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_01861_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_01784_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_01782_),
    .X(net440));
 sg13g2_buf_4 fanout441 (.X(net441),
    .A(_01779_));
 sg13g2_buf_8 fanout442 (.A(_01776_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_01766_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_01762_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_01759_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_01754_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_01253_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_01180_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_00983_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_00968_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_00922_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_00918_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_00896_),
    .X(net453));
 sg13g2_buf_4 fanout454 (.X(net454),
    .A(_05109_));
 sg13g2_buf_4 fanout455 (.X(net455),
    .A(_05104_));
 sg13g2_buf_2 fanout456 (.A(_05100_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_05059_),
    .X(net457));
 sg13g2_buf_4 fanout458 (.X(net458),
    .A(_04646_));
 sg13g2_buf_2 fanout459 (.A(_02748_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_02429_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_02410_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_02347_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_02345_),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_02010_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_02009_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_02004_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_01925_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_01908_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_01891_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_01783_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_01781_),
    .X(net471));
 sg13g2_buf_4 fanout472 (.X(net472),
    .A(_01778_));
 sg13g2_buf_4 fanout473 (.X(net473),
    .A(_01775_));
 sg13g2_buf_2 fanout474 (.A(_01761_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_01760_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_00948_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_00946_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_00917_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_05064_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_05063_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_04656_),
    .X(net481));
 sg13g2_tielo _10617__482 (.L_LO(net482));
 sg13g2_tielo _10618__483 (.L_LO(net483));
 sg13g2_tielo _10619__484 (.L_LO(net484));
 sg13g2_tielo _10620__485 (.L_LO(net485));
 sg13g2_tielo _10625__486 (.L_LO(net486));
 sg13g2_tielo _10626__487 (.L_LO(net487));
 sg13g2_tielo _10627__488 (.L_LO(net488));
 sg13g2_tielo _10628__489 (.L_LO(net489));
 sg13g2_tiehi \B[1]$_SDFF_PN0__491  (.L_HI(net491));
 sg13g2_tiehi \G[0]$_SDFF_PN0__492  (.L_HI(net492));
 sg13g2_tiehi \G[1]$_SDFF_PN0__493  (.L_HI(net493));
 sg13g2_tiehi \R[0]$_SDFF_PN0__494  (.L_HI(net494));
 sg13g2_tiehi \R[1]$_SDFF_PN0__495  (.L_HI(net495));
 sg13g2_tiehi \btn_down_debounce.button_sync_0$_SDFF_PN0__496  (.L_HI(net496));
 sg13g2_tiehi \btn_down_debounce.button_sync_1$_SDFF_PN0__497  (.L_HI(net497));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[0]$_SDFF_PP0__498  (.L_HI(net498));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[10]$_SDFF_PP0__499  (.L_HI(net499));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[11]$_SDFF_PP0__500  (.L_HI(net500));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[12]$_SDFF_PP0__501  (.L_HI(net501));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[13]$_SDFF_PP0__502  (.L_HI(net502));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[14]$_SDFF_PP0__503  (.L_HI(net503));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[15]$_SDFF_PP0__504  (.L_HI(net504));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[16]$_SDFF_PP0__505  (.L_HI(net505));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[17]$_SDFF_PP0__506  (.L_HI(net506));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[1]$_SDFF_PP0__507  (.L_HI(net507));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[2]$_SDFF_PP0__508  (.L_HI(net508));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[3]$_SDFF_PP0__509  (.L_HI(net509));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[4]$_SDFF_PP0__510  (.L_HI(net510));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[5]$_SDFF_PP0__511  (.L_HI(net511));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[6]$_SDFF_PP0__512  (.L_HI(net512));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[7]$_SDFF_PP0__513  (.L_HI(net513));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[8]$_SDFF_PP0__514  (.L_HI(net514));
 sg13g2_tiehi \btn_down_debounce.debounce_counter[9]$_SDFF_PP0__515  (.L_HI(net515));
 sg13g2_tiehi \btn_down_debounce.debounced$_SDFFE_PN0P__516  (.L_HI(net516));
 sg13g2_tiehi \btn_left_debounce.button_sync_0$_SDFF_PN0__517  (.L_HI(net517));
 sg13g2_tiehi \btn_left_debounce.button_sync_1$_SDFF_PN0__518  (.L_HI(net518));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[0]$_SDFF_PP0__519  (.L_HI(net519));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[10]$_SDFF_PP0__520  (.L_HI(net520));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[11]$_SDFF_PP0__521  (.L_HI(net521));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[12]$_SDFF_PP0__522  (.L_HI(net522));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[13]$_SDFF_PP0__523  (.L_HI(net523));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[14]$_SDFF_PP0__524  (.L_HI(net524));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[15]$_SDFF_PP0__525  (.L_HI(net525));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[16]$_SDFF_PP0__526  (.L_HI(net526));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[17]$_SDFF_PP0__527  (.L_HI(net527));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[1]$_SDFF_PP0__528  (.L_HI(net528));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[2]$_SDFF_PP0__529  (.L_HI(net529));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[3]$_SDFF_PP0__530  (.L_HI(net530));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[4]$_SDFF_PP0__531  (.L_HI(net531));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[5]$_SDFF_PP0__532  (.L_HI(net532));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[6]$_SDFF_PP0__533  (.L_HI(net533));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[7]$_SDFF_PP0__534  (.L_HI(net534));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[8]$_SDFF_PP0__535  (.L_HI(net535));
 sg13g2_tiehi \btn_left_debounce.debounce_counter[9]$_SDFF_PP0__536  (.L_HI(net536));
 sg13g2_tiehi \btn_left_debounce.debounced$_SDFFE_PN0P__537  (.L_HI(net537));
 sg13g2_tiehi \btn_right_debounce.button_sync_0$_SDFF_PN0__538  (.L_HI(net538));
 sg13g2_tiehi \btn_right_debounce.button_sync_1$_SDFF_PN0__539  (.L_HI(net539));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[0]$_SDFF_PP0__540  (.L_HI(net540));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[10]$_SDFF_PP0__541  (.L_HI(net541));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[11]$_SDFF_PP0__542  (.L_HI(net542));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[12]$_SDFF_PP0__543  (.L_HI(net543));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[13]$_SDFF_PP0__544  (.L_HI(net544));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[14]$_SDFF_PP0__545  (.L_HI(net545));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[15]$_SDFF_PP0__546  (.L_HI(net546));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[16]$_SDFF_PP0__547  (.L_HI(net547));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[17]$_SDFF_PP0__548  (.L_HI(net548));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[1]$_SDFF_PP0__549  (.L_HI(net549));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[2]$_SDFF_PP0__550  (.L_HI(net550));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[3]$_SDFF_PP0__551  (.L_HI(net551));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[4]$_SDFF_PP0__552  (.L_HI(net552));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[5]$_SDFF_PP0__553  (.L_HI(net553));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[6]$_SDFF_PP0__554  (.L_HI(net554));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[7]$_SDFF_PP0__555  (.L_HI(net555));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[8]$_SDFF_PP0__556  (.L_HI(net556));
 sg13g2_tiehi \btn_right_debounce.debounce_counter[9]$_SDFF_PP0__557  (.L_HI(net557));
 sg13g2_tiehi \btn_right_debounce.debounced$_SDFFE_PN0P__558  (.L_HI(net558));
 sg13g2_tiehi \btn_up_debounce.button_sync_0$_SDFF_PN0__559  (.L_HI(net559));
 sg13g2_tiehi \btn_up_debounce.button_sync_1$_SDFF_PN0__560  (.L_HI(net560));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[0]$_SDFF_PP0__561  (.L_HI(net561));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[10]$_SDFF_PP0__562  (.L_HI(net562));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[11]$_SDFF_PP0__563  (.L_HI(net563));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[12]$_SDFF_PP0__564  (.L_HI(net564));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[13]$_SDFF_PP0__565  (.L_HI(net565));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[14]$_SDFF_PP0__566  (.L_HI(net566));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[15]$_SDFF_PP0__567  (.L_HI(net567));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[16]$_SDFF_PP0__568  (.L_HI(net568));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[17]$_SDFF_PP0__569  (.L_HI(net569));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[1]$_SDFF_PP0__570  (.L_HI(net570));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[2]$_SDFF_PP0__571  (.L_HI(net571));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[3]$_SDFF_PP0__572  (.L_HI(net572));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[4]$_SDFF_PP0__573  (.L_HI(net573));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[5]$_SDFF_PP0__574  (.L_HI(net574));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[6]$_SDFF_PP0__575  (.L_HI(net575));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[7]$_SDFF_PP0__576  (.L_HI(net576));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[8]$_SDFF_PP0__577  (.L_HI(net577));
 sg13g2_tiehi \btn_up_debounce.debounce_counter[9]$_SDFF_PP0__578  (.L_HI(net578));
 sg13g2_tiehi \btn_up_debounce.debounced$_SDFFE_PN0P__579  (.L_HI(net579));
 sg13g2_tiehi \debug_controller_inst.data_out[0]$_SDFFE_PN0P__580  (.L_HI(net580));
 sg13g2_tiehi \debug_controller_inst.data_out[1]$_SDFFE_PN0P__581  (.L_HI(net581));
 sg13g2_tiehi \debug_controller_inst.data_out[2]$_SDFFE_PN0P__582  (.L_HI(net582));
 sg13g2_tiehi \debug_controller_inst.data_out[3]$_SDFFE_PN0P__583  (.L_HI(net583));
 sg13g2_tiehi \debug_controller_inst.data_out_en$_SDFF_PN0__584  (.L_HI(net584));
 sg13g2_tiehi \debug_controller_inst.force_move[0]$_SDFF_PN0__585  (.L_HI(net585));
 sg13g2_tiehi \debug_controller_inst.force_move[1]$_SDFF_PN0__586  (.L_HI(net586));
 sg13g2_tiehi \debug_controller_inst.force_move[2]$_SDFF_PN0__587  (.L_HI(net587));
 sg13g2_tiehi \debug_controller_inst.force_move[3]$_SDFF_PN0__588  (.L_HI(net588));
 sg13g2_tiehi \debug_controller_inst.grid_addr[0]$_SDFFE_PN0P__589  (.L_HI(net589));
 sg13g2_tiehi \debug_controller_inst.grid_addr[1]$_SDFFE_PN0P__590  (.L_HI(net590));
 sg13g2_tiehi \debug_controller_inst.grid_addr[2]$_SDFFE_PN0P__591  (.L_HI(net591));
 sg13g2_tiehi \debug_controller_inst.grid_addr[3]$_SDFFE_PN0P__592  (.L_HI(net592));
 sg13g2_tiehi \debug_controller_inst.grid_out_addr[0]$_SDFFE_PN0P__593  (.L_HI(net593));
 sg13g2_tiehi \debug_controller_inst.grid_out_addr[1]$_SDFFE_PN0P__594  (.L_HI(net594));
 sg13g2_tiehi \debug_controller_inst.grid_out_addr[2]$_SDFFE_PN0P__595  (.L_HI(net595));
 sg13g2_tiehi \debug_controller_inst.grid_out_addr[3]$_SDFFE_PN0P__596  (.L_HI(net596));
 sg13g2_tiehi \debug_controller_inst.grid_out_data[0]$_SDFFE_PN0P__597  (.L_HI(net597));
 sg13g2_tiehi \debug_controller_inst.grid_out_data[1]$_SDFFE_PN0P__598  (.L_HI(net598));
 sg13g2_tiehi \debug_controller_inst.grid_out_data[2]$_SDFFE_PN0P__599  (.L_HI(net599));
 sg13g2_tiehi \debug_controller_inst.grid_out_data[3]$_SDFFE_PN0P__600  (.L_HI(net600));
 sg13g2_tiehi \debug_controller_inst.grid_out_valid$_SDFF_PN0__601  (.L_HI(net601));
 sg13g2_tiehi \game_logic_inst.add_new_tiles[0]$_SDFFE_PN0P__602  (.L_HI(net602));
 sg13g2_tiehi \game_logic_inst.add_new_tiles[1]$_SDFFE_PN0P__603  (.L_HI(net603));
 sg13g2_tiehi \game_logic_inst.added_tile_index[0]$_SDFF_PP0__604  (.L_HI(net604));
 sg13g2_tiehi \game_logic_inst.added_tile_index[1]$_SDFF_PP0__605  (.L_HI(net605));
 sg13g2_tiehi \game_logic_inst.added_tile_index[2]$_SDFF_PP0__606  (.L_HI(net606));
 sg13g2_tiehi \game_logic_inst.added_tile_index[3]$_SDFF_PP0__607  (.L_HI(net607));
 sg13g2_tiehi \game_logic_inst.calculate_move$_SDFFE_PN0P__608  (.L_HI(net608));
 sg13g2_tiehi \game_logic_inst.current_direction[1]$_DFF_P__609  (.L_HI(net609));
 sg13g2_tiehi \game_logic_inst.current_direction[2]$_DFF_P__610  (.L_HI(net610));
 sg13g2_tiehi \game_logic_inst.current_direction[3]$_DFF_P__611  (.L_HI(net611));
 sg13g2_tiehi \game_logic_inst.current_row_index[0]$_SDFFE_PN0P__612  (.L_HI(net612));
 sg13g2_tiehi \game_logic_inst.current_row_index[1]$_SDFFE_PN0P__613  (.L_HI(net613));
 sg13g2_tiehi \game_logic_inst.debug_move_reg$_SDFFE_PN0P__614  (.L_HI(net614));
 sg13g2_tiehi \game_logic_inst.game_started$_SDFF_PN0__615  (.L_HI(net615));
 sg13g2_tiehi \game_logic_inst.grid[0]$_DFF_P__616  (.L_HI(net616));
 sg13g2_tiehi \game_logic_inst.grid[10]$_DFF_P__617  (.L_HI(net617));
 sg13g2_tiehi \game_logic_inst.grid[11]$_DFF_P__618  (.L_HI(net618));
 sg13g2_tiehi \game_logic_inst.grid[12]$_DFF_P__619  (.L_HI(net619));
 sg13g2_tiehi \game_logic_inst.grid[13]$_DFF_P__620  (.L_HI(net620));
 sg13g2_tiehi \game_logic_inst.grid[14]$_DFF_P__621  (.L_HI(net621));
 sg13g2_tiehi \game_logic_inst.grid[15]$_DFF_P__622  (.L_HI(net622));
 sg13g2_tiehi \game_logic_inst.grid[16]$_DFF_P__623  (.L_HI(net623));
 sg13g2_tiehi \game_logic_inst.grid[17]$_DFF_P__624  (.L_HI(net624));
 sg13g2_tiehi \game_logic_inst.grid[18]$_DFF_P__625  (.L_HI(net625));
 sg13g2_tiehi \game_logic_inst.grid[19]$_DFF_P__626  (.L_HI(net626));
 sg13g2_tiehi \game_logic_inst.grid[1]$_DFF_P__627  (.L_HI(net627));
 sg13g2_tiehi \game_logic_inst.grid[20]$_DFF_P__628  (.L_HI(net628));
 sg13g2_tiehi \game_logic_inst.grid[21]$_DFF_P__629  (.L_HI(net629));
 sg13g2_tiehi \game_logic_inst.grid[22]$_DFF_P__630  (.L_HI(net630));
 sg13g2_tiehi \game_logic_inst.grid[23]$_DFF_P__631  (.L_HI(net631));
 sg13g2_tiehi \game_logic_inst.grid[24]$_DFF_P__632  (.L_HI(net632));
 sg13g2_tiehi \game_logic_inst.grid[25]$_DFF_P__633  (.L_HI(net633));
 sg13g2_tiehi \game_logic_inst.grid[26]$_DFF_P__634  (.L_HI(net634));
 sg13g2_tiehi \game_logic_inst.grid[27]$_DFF_P__635  (.L_HI(net635));
 sg13g2_tiehi \game_logic_inst.grid[28]$_DFF_P__636  (.L_HI(net636));
 sg13g2_tiehi \game_logic_inst.grid[29]$_DFF_P__637  (.L_HI(net637));
 sg13g2_tiehi \game_logic_inst.grid[2]$_DFF_P__638  (.L_HI(net638));
 sg13g2_tiehi \game_logic_inst.grid[30]$_DFF_P__639  (.L_HI(net639));
 sg13g2_tiehi \game_logic_inst.grid[31]$_DFF_P__640  (.L_HI(net640));
 sg13g2_tiehi \game_logic_inst.grid[32]$_DFF_P__641  (.L_HI(net641));
 sg13g2_tiehi \game_logic_inst.grid[33]$_DFF_P__642  (.L_HI(net642));
 sg13g2_tiehi \game_logic_inst.grid[34]$_DFF_P__643  (.L_HI(net643));
 sg13g2_tiehi \game_logic_inst.grid[35]$_DFF_P__644  (.L_HI(net644));
 sg13g2_tiehi \game_logic_inst.grid[36]$_DFF_P__645  (.L_HI(net645));
 sg13g2_tiehi \game_logic_inst.grid[37]$_DFF_P__646  (.L_HI(net646));
 sg13g2_tiehi \game_logic_inst.grid[38]$_DFF_P__647  (.L_HI(net647));
 sg13g2_tiehi \game_logic_inst.grid[39]$_DFF_P__648  (.L_HI(net648));
 sg13g2_tiehi \game_logic_inst.grid[3]$_DFF_P__649  (.L_HI(net649));
 sg13g2_tiehi \game_logic_inst.grid[40]$_DFF_P__650  (.L_HI(net650));
 sg13g2_tiehi \game_logic_inst.grid[41]$_DFF_P__651  (.L_HI(net651));
 sg13g2_tiehi \game_logic_inst.grid[42]$_DFF_P__652  (.L_HI(net652));
 sg13g2_tiehi \game_logic_inst.grid[43]$_DFF_P__653  (.L_HI(net653));
 sg13g2_tiehi \game_logic_inst.grid[44]$_DFF_P__654  (.L_HI(net654));
 sg13g2_tiehi \game_logic_inst.grid[45]$_DFF_P__655  (.L_HI(net655));
 sg13g2_tiehi \game_logic_inst.grid[46]$_DFF_P__656  (.L_HI(net656));
 sg13g2_tiehi \game_logic_inst.grid[47]$_DFF_P__657  (.L_HI(net657));
 sg13g2_tiehi \game_logic_inst.grid[48]$_DFF_P__658  (.L_HI(net658));
 sg13g2_tiehi \game_logic_inst.grid[49]$_DFF_P__659  (.L_HI(net659));
 sg13g2_tiehi \game_logic_inst.grid[4]$_DFF_P__660  (.L_HI(net660));
 sg13g2_tiehi \game_logic_inst.grid[50]$_DFF_P__661  (.L_HI(net661));
 sg13g2_tiehi \game_logic_inst.grid[51]$_DFF_P__662  (.L_HI(net662));
 sg13g2_tiehi \game_logic_inst.grid[52]$_DFF_P__663  (.L_HI(net663));
 sg13g2_tiehi \game_logic_inst.grid[53]$_DFF_P__664  (.L_HI(net664));
 sg13g2_tiehi \game_logic_inst.grid[54]$_DFF_P__665  (.L_HI(net665));
 sg13g2_tiehi \game_logic_inst.grid[55]$_DFF_P__666  (.L_HI(net666));
 sg13g2_tiehi \game_logic_inst.grid[56]$_DFF_P__667  (.L_HI(net667));
 sg13g2_tiehi \game_logic_inst.grid[57]$_DFF_P__668  (.L_HI(net668));
 sg13g2_tiehi \game_logic_inst.grid[58]$_DFF_P__669  (.L_HI(net669));
 sg13g2_tiehi \game_logic_inst.grid[59]$_DFF_P__670  (.L_HI(net670));
 sg13g2_tiehi \game_logic_inst.grid[5]$_DFF_P__671  (.L_HI(net671));
 sg13g2_tiehi \game_logic_inst.grid[60]$_DFF_P__672  (.L_HI(net672));
 sg13g2_tiehi \game_logic_inst.grid[61]$_DFF_P__673  (.L_HI(net673));
 sg13g2_tiehi \game_logic_inst.grid[62]$_DFF_P__674  (.L_HI(net674));
 sg13g2_tiehi \game_logic_inst.grid[63]$_DFF_P__675  (.L_HI(net675));
 sg13g2_tiehi \game_logic_inst.grid[6]$_DFF_P__676  (.L_HI(net676));
 sg13g2_tiehi \game_logic_inst.grid[7]$_DFF_P__677  (.L_HI(net677));
 sg13g2_tiehi \game_logic_inst.grid[8]$_DFF_P__678  (.L_HI(net678));
 sg13g2_tiehi \game_logic_inst.grid[9]$_DFF_P__679  (.L_HI(net679));
 sg13g2_tiehi \game_logic_inst.lfsr_shift[0]$_SDFF_PN0__680  (.L_HI(net680));
 sg13g2_tiehi \game_logic_inst.lfsr_shift[1]$_SDFF_PN0__681  (.L_HI(net681));
 sg13g2_tiehi \game_logic_inst.prev_any_button_pressed$_SDFF_PN0__682  (.L_HI(net682));
 sg13g2_tiehi \game_logic_inst.should_transpose$_SDFFE_PN0P__683  (.L_HI(net683));
 sg13g2_tiehi \game_logic_inst.valid_move$_SDFFE_PN0P__684  (.L_HI(net684));
 sg13g2_tiehi \grid[0]$_SDFFE_PN0P__685  (.L_HI(net685));
 sg13g2_tiehi \grid[10]$_SDFFE_PN0P__686  (.L_HI(net686));
 sg13g2_tiehi \grid[11]$_SDFFE_PN0P__687  (.L_HI(net687));
 sg13g2_tiehi \grid[12]$_SDFFE_PN0P__688  (.L_HI(net688));
 sg13g2_tiehi \grid[13]$_SDFFE_PN0P__689  (.L_HI(net689));
 sg13g2_tiehi \grid[14]$_SDFFE_PN0P__690  (.L_HI(net690));
 sg13g2_tiehi \grid[15]$_SDFFE_PN0P__691  (.L_HI(net691));
 sg13g2_tiehi \grid[16]$_SDFFE_PN0P__692  (.L_HI(net692));
 sg13g2_tiehi \grid[17]$_SDFFE_PN0P__693  (.L_HI(net693));
 sg13g2_tiehi \grid[18]$_SDFFE_PN0P__694  (.L_HI(net694));
 sg13g2_tiehi \grid[19]$_SDFFE_PN0P__695  (.L_HI(net695));
 sg13g2_tiehi \grid[1]$_SDFFE_PN0P__696  (.L_HI(net696));
 sg13g2_tiehi \grid[20]$_SDFFE_PN0P__697  (.L_HI(net697));
 sg13g2_tiehi \grid[21]$_SDFFE_PN0P__698  (.L_HI(net698));
 sg13g2_tiehi \grid[22]$_SDFFE_PN0P__699  (.L_HI(net699));
 sg13g2_tiehi \grid[23]$_SDFFE_PN0P__700  (.L_HI(net700));
 sg13g2_tiehi \grid[24]$_SDFFE_PN0P__701  (.L_HI(net701));
 sg13g2_tiehi \grid[25]$_SDFFE_PN0P__702  (.L_HI(net702));
 sg13g2_tiehi \grid[26]$_SDFFE_PN0P__703  (.L_HI(net703));
 sg13g2_tiehi \grid[27]$_SDFFE_PN0P__704  (.L_HI(net704));
 sg13g2_tiehi \grid[28]$_SDFFE_PN0P__705  (.L_HI(net705));
 sg13g2_tiehi \grid[29]$_SDFFE_PN0P__706  (.L_HI(net706));
 sg13g2_tiehi \grid[2]$_SDFFE_PN0P__707  (.L_HI(net707));
 sg13g2_tiehi \grid[30]$_SDFFE_PN0P__708  (.L_HI(net708));
 sg13g2_tiehi \grid[31]$_SDFFE_PN0P__709  (.L_HI(net709));
 sg13g2_tiehi \grid[32]$_SDFFE_PN0P__710  (.L_HI(net710));
 sg13g2_tiehi \grid[33]$_SDFFE_PN0P__711  (.L_HI(net711));
 sg13g2_tiehi \grid[34]$_SDFFE_PN0P__712  (.L_HI(net712));
 sg13g2_tiehi \grid[35]$_SDFFE_PN0P__713  (.L_HI(net713));
 sg13g2_tiehi \grid[36]$_SDFFE_PN0P__714  (.L_HI(net714));
 sg13g2_tiehi \grid[37]$_SDFFE_PN0P__715  (.L_HI(net715));
 sg13g2_tiehi \grid[38]$_SDFFE_PN0P__716  (.L_HI(net716));
 sg13g2_tiehi \grid[39]$_SDFFE_PN0P__717  (.L_HI(net717));
 sg13g2_tiehi \grid[3]$_SDFFE_PN0P__718  (.L_HI(net718));
 sg13g2_tiehi \grid[40]$_SDFFE_PN0P__719  (.L_HI(net719));
 sg13g2_tiehi \grid[41]$_SDFFE_PN0P__720  (.L_HI(net720));
 sg13g2_tiehi \grid[42]$_SDFFE_PN0P__721  (.L_HI(net721));
 sg13g2_tiehi \grid[43]$_SDFFE_PN0P__722  (.L_HI(net722));
 sg13g2_tiehi \grid[44]$_SDFFE_PN0P__723  (.L_HI(net723));
 sg13g2_tiehi \grid[45]$_SDFFE_PN0P__724  (.L_HI(net724));
 sg13g2_tiehi \grid[46]$_SDFFE_PN0P__725  (.L_HI(net725));
 sg13g2_tiehi \grid[47]$_SDFFE_PN0P__726  (.L_HI(net726));
 sg13g2_tiehi \grid[48]$_SDFFE_PN0P__727  (.L_HI(net727));
 sg13g2_tiehi \grid[49]$_SDFFE_PN0P__728  (.L_HI(net728));
 sg13g2_tiehi \grid[4]$_SDFFE_PN0P__729  (.L_HI(net729));
 sg13g2_tiehi \grid[50]$_SDFFE_PN0P__730  (.L_HI(net730));
 sg13g2_tiehi \grid[51]$_SDFFE_PN0P__731  (.L_HI(net731));
 sg13g2_tiehi \grid[52]$_SDFFE_PN0P__732  (.L_HI(net732));
 sg13g2_tiehi \grid[53]$_SDFFE_PN0P__733  (.L_HI(net733));
 sg13g2_tiehi \grid[54]$_SDFFE_PN0P__734  (.L_HI(net734));
 sg13g2_tiehi \grid[55]$_SDFFE_PN0P__735  (.L_HI(net735));
 sg13g2_tiehi \grid[56]$_SDFFE_PN0P__736  (.L_HI(net736));
 sg13g2_tiehi \grid[57]$_SDFFE_PN0P__737  (.L_HI(net737));
 sg13g2_tiehi \grid[58]$_SDFFE_PN0P__738  (.L_HI(net738));
 sg13g2_tiehi \grid[59]$_SDFFE_PN0P__739  (.L_HI(net739));
 sg13g2_tiehi \grid[5]$_SDFFE_PN0P__740  (.L_HI(net740));
 sg13g2_tiehi \grid[60]$_SDFFE_PN0P__741  (.L_HI(net741));
 sg13g2_tiehi \grid[61]$_SDFFE_PN0P__742  (.L_HI(net742));
 sg13g2_tiehi \grid[62]$_SDFFE_PN0P__743  (.L_HI(net743));
 sg13g2_tiehi \grid[63]$_SDFFE_PN0P__744  (.L_HI(net744));
 sg13g2_tiehi \grid[6]$_SDFFE_PN0P__745  (.L_HI(net745));
 sg13g2_tiehi \grid[7]$_SDFFE_PN0P__746  (.L_HI(net746));
 sg13g2_tiehi \grid[8]$_SDFFE_PN0P__747  (.L_HI(net747));
 sg13g2_tiehi \grid[9]$_SDFFE_PN0P__748  (.L_HI(net748));
 sg13g2_tiehi \lfsr_inst.lfsr[0]$_SDFF_PN0__749  (.L_HI(net749));
 sg13g2_tiehi \lfsr_inst.lfsr[10]$_SDFF_PN0__750  (.L_HI(net750));
 sg13g2_tiehi \lfsr_inst.lfsr[11]$_SDFF_PN1__751  (.L_HI(net751));
 sg13g2_tiehi \lfsr_inst.lfsr[12]$_SDFF_PN1__752  (.L_HI(net752));
 sg13g2_tiehi \lfsr_inst.lfsr[13]$_SDFF_PN1__753  (.L_HI(net753));
 sg13g2_tiehi \lfsr_inst.lfsr[14]$_SDFF_PN1__754  (.L_HI(net754));
 sg13g2_tiehi \lfsr_inst.lfsr[15]$_SDFF_PN1__755  (.L_HI(net755));
 sg13g2_tiehi \lfsr_inst.lfsr[16]$_SDFF_PN0__756  (.L_HI(net756));
 sg13g2_tiehi \lfsr_inst.lfsr[17]$_SDFF_PN0__757  (.L_HI(net757));
 sg13g2_tiehi \lfsr_inst.lfsr[18]$_SDFF_PN0__758  (.L_HI(net758));
 sg13g2_tiehi \lfsr_inst.lfsr[19]$_SDFF_PN1__759  (.L_HI(net759));
 sg13g2_tiehi \lfsr_inst.lfsr[1]$_SDFF_PN1__760  (.L_HI(net760));
 sg13g2_tiehi \lfsr_inst.lfsr[20]$_SDFF_PN0__761  (.L_HI(net761));
 sg13g2_tiehi \lfsr_inst.lfsr[21]$_SDFF_PN0__762  (.L_HI(net762));
 sg13g2_tiehi \lfsr_inst.lfsr[22]$_SDFF_PN1__763  (.L_HI(net763));
 sg13g2_tiehi \lfsr_inst.lfsr[23]$_SDFF_PN0__764  (.L_HI(net764));
 sg13g2_tiehi \lfsr_inst.lfsr[24]$_SDFF_PN0__765  (.L_HI(net765));
 sg13g2_tiehi \lfsr_inst.lfsr[25]$_SDFF_PN0__766  (.L_HI(net766));
 sg13g2_tiehi \lfsr_inst.lfsr[26]$_SDFF_PN0__767  (.L_HI(net767));
 sg13g2_tiehi \lfsr_inst.lfsr[27]$_SDFF_PN0__768  (.L_HI(net768));
 sg13g2_tiehi \lfsr_inst.lfsr[28]$_SDFF_PN0__769  (.L_HI(net769));
 sg13g2_tiehi \lfsr_inst.lfsr[29]$_SDFF_PN1__770  (.L_HI(net770));
 sg13g2_tiehi \lfsr_inst.lfsr[2]$_SDFF_PN0__771  (.L_HI(net771));
 sg13g2_tiehi \lfsr_inst.lfsr[30]$_SDFF_PN0__772  (.L_HI(net772));
 sg13g2_tiehi \lfsr_inst.lfsr[31]$_SDFF_PN0__773  (.L_HI(net773));
 sg13g2_tiehi \lfsr_inst.lfsr[3]$_SDFF_PN1__774  (.L_HI(net774));
 sg13g2_tiehi \lfsr_inst.lfsr[4]$_SDFF_PN1__775  (.L_HI(net775));
 sg13g2_tiehi \lfsr_inst.lfsr[5]$_SDFF_PN1__776  (.L_HI(net776));
 sg13g2_tiehi \lfsr_inst.lfsr[6]$_SDFF_PN1__777  (.L_HI(net777));
 sg13g2_tiehi \lfsr_inst.lfsr[7]$_SDFF_PN1__778  (.L_HI(net778));
 sg13g2_tiehi \lfsr_inst.lfsr[8]$_SDFF_PN0__779  (.L_HI(net779));
 sg13g2_tiehi \lfsr_inst.lfsr[9]$_SDFF_PN1__780  (.L_HI(net780));
 sg13g2_tiehi \new_tiles[0]$_DFFE_PP__781  (.L_HI(net781));
 sg13g2_tiehi \new_tiles[10]$_DFFE_PP__782  (.L_HI(net782));
 sg13g2_tiehi \new_tiles[11]$_DFFE_PP__783  (.L_HI(net783));
 sg13g2_tiehi \new_tiles[12]$_DFFE_PP__784  (.L_HI(net784));
 sg13g2_tiehi \new_tiles[13]$_DFFE_PP__785  (.L_HI(net785));
 sg13g2_tiehi \new_tiles[14]$_DFFE_PP__786  (.L_HI(net786));
 sg13g2_tiehi \new_tiles[15]$_DFFE_PP__787  (.L_HI(net787));
 sg13g2_tiehi \new_tiles[1]$_DFFE_PP__788  (.L_HI(net788));
 sg13g2_tiehi \new_tiles[2]$_DFFE_PP__789  (.L_HI(net789));
 sg13g2_tiehi \new_tiles[3]$_DFFE_PP__790  (.L_HI(net790));
 sg13g2_tiehi \new_tiles[4]$_DFFE_PP__791  (.L_HI(net791));
 sg13g2_tiehi \new_tiles[5]$_DFFE_PP__792  (.L_HI(net792));
 sg13g2_tiehi \new_tiles[6]$_DFFE_PP__793  (.L_HI(net793));
 sg13g2_tiehi \new_tiles[7]$_DFFE_PP__794  (.L_HI(net794));
 sg13g2_tiehi \new_tiles[8]$_DFFE_PP__795  (.L_HI(net795));
 sg13g2_tiehi \new_tiles[9]$_DFFE_PP__796  (.L_HI(net796));
 sg13g2_tiehi \new_tiles_counter[0]$_DFFE_PP__797  (.L_HI(net797));
 sg13g2_tiehi \new_tiles_counter[1]$_DFFE_PP__798  (.L_HI(net798));
 sg13g2_tiehi \new_tiles_counter[2]$_DFFE_PP__799  (.L_HI(net799));
 sg13g2_tiehi \new_tiles_counter[3]$_DFFE_PP__800  (.L_HI(net800));
 sg13g2_tiehi \new_tiles_counter[4]$_DFFE_PP__801  (.L_HI(net801));
 sg13g2_tiehi \show_welcome_screen$_SDFFE_PN1P__802  (.L_HI(net802));
 sg13g2_tiehi \vga_sync_gen.hpos[0]$_SDFF_PP0__803  (.L_HI(net803));
 sg13g2_tiehi \vga_sync_gen.hpos[1]$_SDFF_PP0__804  (.L_HI(net804));
 sg13g2_tiehi \vga_sync_gen.hpos[2]$_SDFF_PP0__805  (.L_HI(net805));
 sg13g2_tiehi \vga_sync_gen.hpos[3]$_SDFF_PP0__806  (.L_HI(net806));
 sg13g2_tiehi \vga_sync_gen.hpos[4]$_SDFF_PP0__807  (.L_HI(net807));
 sg13g2_tiehi \vga_sync_gen.hpos[5]$_SDFF_PP0__808  (.L_HI(net808));
 sg13g2_tiehi \vga_sync_gen.hpos[6]$_SDFF_PP0__809  (.L_HI(net809));
 sg13g2_tiehi \vga_sync_gen.hpos[7]$_SDFF_PP0__810  (.L_HI(net810));
 sg13g2_tiehi \vga_sync_gen.hpos[8]$_SDFF_PP0__811  (.L_HI(net811));
 sg13g2_tiehi \vga_sync_gen.hpos[9]$_SDFF_PP0__812  (.L_HI(net812));
 sg13g2_tiehi \vga_sync_gen.hsync$_DFF_P__813  (.L_HI(net813));
 sg13g2_tiehi \vga_sync_gen.vpos[0]$_SDFFCE_PP0P__814  (.L_HI(net814));
 sg13g2_tiehi \vga_sync_gen.vpos[1]$_SDFFCE_PP0P__815  (.L_HI(net815));
 sg13g2_tiehi \vga_sync_gen.vpos[2]$_SDFFCE_PP0P__816  (.L_HI(net816));
 sg13g2_tiehi \vga_sync_gen.vpos[3]$_SDFFCE_PP0P__817  (.L_HI(net817));
 sg13g2_tiehi \vga_sync_gen.vpos[4]$_SDFFCE_PP0P__818  (.L_HI(net818));
 sg13g2_tiehi \vga_sync_gen.vpos[5]$_SDFFCE_PP0P__819  (.L_HI(net819));
 sg13g2_tiehi \vga_sync_gen.vpos[6]$_SDFFCE_PP0P__820  (.L_HI(net820));
 sg13g2_tiehi \vga_sync_gen.vpos[7]$_SDFFCE_PP0P__821  (.L_HI(net821));
 sg13g2_tiehi \vga_sync_gen.vpos[8]$_SDFFCE_PP0P__822  (.L_HI(net822));
 sg13g2_tiehi \vga_sync_gen.vpos[9]$_SDFFCE_PP0P__823  (.L_HI(net823));
 sg13g2_tiehi \vga_sync_gen.vsync$_DFF_P__824  (.L_HI(net824));
 sg13g2_tiehi \vsync_prev$_SDFF_PN0__825  (.L_HI(net825));
 sg13g2_tiehi \welcome_screen_inst.grid[11]$_SDFFCE_PP0P__826  (.L_HI(net826));
 sg13g2_tiehi \welcome_screen_inst.grid[15]$_SDFFCE_PP0P__827  (.L_HI(net827));
 sg13g2_tiehi \welcome_screen_inst.grid[19]$_SDFFCE_PP0P__828  (.L_HI(net828));
 sg13g2_tiehi \welcome_screen_inst.grid[23]$_SDFFCE_PP0P__829  (.L_HI(net829));
 sg13g2_tiehi \welcome_screen_inst.grid[27]$_SDFFCE_PP0P__830  (.L_HI(net830));
 sg13g2_tiehi \welcome_screen_inst.grid[31]$_SDFFCE_PP0P__831  (.L_HI(net831));
 sg13g2_tiehi \welcome_screen_inst.grid[35]$_SDFFCE_PP0P__832  (.L_HI(net832));
 sg13g2_tiehi \welcome_screen_inst.grid[39]$_SDFFCE_PP0P__833  (.L_HI(net833));
 sg13g2_tiehi \welcome_screen_inst.grid[3]$_SDFFCE_PP0P__834  (.L_HI(net834));
 sg13g2_tiehi \welcome_screen_inst.grid[43]$_SDFFCE_PP0P__835  (.L_HI(net835));
 sg13g2_tiehi \welcome_screen_inst.grid[47]$_SDFFCE_PP0P__836  (.L_HI(net836));
 sg13g2_tiehi \welcome_screen_inst.grid[51]$_SDFFCE_PP0P__837  (.L_HI(net837));
 sg13g2_tiehi \welcome_screen_inst.grid[55]$_SDFFCE_PP0P__838  (.L_HI(net838));
 sg13g2_tiehi \welcome_screen_inst.grid[59]$_SDFFCE_PP0P__839  (.L_HI(net839));
 sg13g2_tiehi \welcome_screen_inst.grid[61]$_SDFFCE_PP0P__840  (.L_HI(net840));
 sg13g2_tiehi \welcome_screen_inst.grid[7]$_SDFFCE_PP0P__841  (.L_HI(net841));
 sg13g2_tiehi \welcome_screen_inst.welcome_counter[0]$_SDFFE_PN0P__842  (.L_HI(net842));
 sg13g2_tiehi \welcome_screen_inst.welcome_counter[1]$_SDFFE_PN1P__843  (.L_HI(net843));
 sg13g2_tiehi \welcome_screen_inst.welcome_counter[2]$_SDFFE_PN1P__844  (.L_HI(net844));
 sg13g2_tiehi \welcome_screen_inst.welcome_counter[3]$_SDFFE_PN1P__845  (.L_HI(net845));
 sg13g2_tiehi \welcome_screen_inst.welcome_counter[4]$_SDFFE_PN1P__846  (.L_HI(net846));
 sg13g2_buf_4 clkbuf_leaf_1_clk (.X(clknet_leaf_1_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_3_clk (.X(clknet_leaf_3_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkbuf_leaf_5_clk (.X(clknet_leaf_5_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_9_clk (.X(clknet_leaf_9_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_10_clk (.X(clknet_leaf_10_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_11_clk (.X(clknet_leaf_11_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_15_clk (.X(clknet_leaf_15_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_19_clk (.X(clknet_leaf_19_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_22_clk (.X(clknet_leaf_22_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_24_clk (.X(clknet_leaf_24_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_25_clk (.X(clknet_leaf_25_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_26_clk (.X(clknet_leaf_26_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_27_clk (.X(clknet_leaf_27_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_28_clk (.X(clknet_leaf_28_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_29_clk (.X(clknet_leaf_29_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_30_clk (.X(clknet_leaf_30_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_31_clk (.X(clknet_leaf_31_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_32_clk (.X(clknet_leaf_32_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_33_clk (.X(clknet_leaf_33_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_34_clk (.X(clknet_leaf_34_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_35_clk (.X(clknet_leaf_35_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_36_clk (.X(clknet_leaf_36_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_37_clk (.X(clknet_leaf_37_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_38_clk (.X(clknet_leaf_38_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_39_clk (.X(clknet_leaf_39_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_40_clk (.X(clknet_leaf_40_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_41_clk (.X(clknet_leaf_41_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_42_clk (.X(clknet_leaf_42_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_43_clk (.X(clknet_leaf_43_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_44_clk (.X(clknet_leaf_44_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_45_clk (.X(clknet_leaf_45_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_46_clk (.X(clknet_leaf_46_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_47_clk (.X(clknet_leaf_47_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_48_clk (.X(clknet_leaf_48_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_49_clk (.X(clknet_leaf_49_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_50_clk (.X(clknet_leaf_50_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_51_clk (.X(clknet_leaf_51_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_52_clk (.X(clknet_leaf_52_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_53_clk (.X(clknet_leaf_53_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_54_clk (.X(clknet_leaf_54_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_55_clk (.X(clknet_leaf_55_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_56_clk (.X(clknet_leaf_56_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_57_clk (.X(clknet_leaf_57_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_0_0_clk (.X(clknet_4_0_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_1_0_clk (.X(clknet_4_1_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_2_0_clk (.X(clknet_4_2_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_3_0_clk (.X(clknet_4_3_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_4_0_clk (.X(clknet_4_4_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_5_0_clk (.X(clknet_4_5_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_6_0_clk (.X(clknet_4_6_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_7_0_clk (.X(clknet_4_7_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_8_0_clk (.X(clknet_4_8_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_9_0_clk (.X(clknet_4_9_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_10_0_clk (.X(clknet_4_10_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_11_0_clk (.X(clknet_4_11_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_12_0_clk (.X(clknet_4_12_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_13_0_clk (.X(clknet_4_13_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_14_0_clk (.X(clknet_4_14_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_15_0_clk (.X(clknet_4_15_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkload3 (.A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkload4 (.A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkload5 (.A(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_4_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_57_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_leaf_6_clk));
 sg13g2_buf_16 clkload10 (.A(clknet_leaf_7_clk));
 sg13g2_buf_16 clkload11 (.A(clknet_leaf_8_clk));
 sg13g2_buf_16 clkload12 (.A(clknet_leaf_1_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_2_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_56_clk));
 sg13g2_buf_8 clkload15 (.A(clknet_leaf_3_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_21_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_12_clk));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_13_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_20_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_11_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_15_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_18_clk));
 sg13g2_inv_2 clkload23 (.A(clknet_leaf_27_clk));
 sg13g2_inv_4 clkload24 (.A(clknet_leaf_41_clk));
 sg13g2_inv_2 clkload25 (.A(clknet_leaf_43_clk));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_45_clk));
 sg13g2_inv_1 clkload27 (.A(clknet_leaf_51_clk));
 sg13g2_inv_1 clkload28 (.A(clknet_leaf_52_clk));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_39_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_42_clk));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_46_clk));
 sg13g2_inv_1 clkload32 (.A(clknet_leaf_34_clk));
 sg13g2_buf_16 clkload33 (.A(clknet_leaf_35_clk));
 sg13g2_inv_2 clkload34 (.A(clknet_leaf_48_clk));
 sg13g2_inv_2 clkload35 (.A(clknet_leaf_49_clk));
 sg13g2_inv_1 clkload36 (.A(clknet_leaf_24_clk));
 sg13g2_buf_8 clkload37 (.A(clknet_leaf_25_clk));
 sg13g2_buf_8 clkload38 (.A(clknet_leaf_26_clk));
 sg13g2_inv_2 clkload39 (.A(clknet_leaf_30_clk));
 sg13g2_buf_16 clkload40 (.A(clknet_leaf_31_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00383_));
 sg13g2_antennanp ANTENNA_2 (.A(_00420_));
 sg13g2_antennanp ANTENNA_3 (.A(_00422_));
 sg13g2_antennanp ANTENNA_4 (.A(_02067_));
 sg13g2_antennanp ANTENNA_5 (.A(_02067_));
 sg13g2_antennanp ANTENNA_6 (.A(_02400_));
 sg13g2_antennanp ANTENNA_7 (.A(_02400_));
 sg13g2_antennanp ANTENNA_8 (.A(_02400_));
 sg13g2_antennanp ANTENNA_9 (.A(_02672_));
 sg13g2_antennanp ANTENNA_10 (.A(_02672_));
 sg13g2_antennanp ANTENNA_11 (.A(_02672_));
 sg13g2_antennanp ANTENNA_12 (.A(_05057_));
 sg13g2_antennanp ANTENNA_13 (.A(_05057_));
 sg13g2_antennanp ANTENNA_14 (.A(_05057_));
 sg13g2_antennanp ANTENNA_15 (.A(_05057_));
 sg13g2_antennanp ANTENNA_16 (.A(_05057_));
 sg13g2_antennanp ANTENNA_17 (.A(_05057_));
 sg13g2_antennanp ANTENNA_18 (.A(clk));
 sg13g2_antennanp ANTENNA_19 (.A(net22));
 sg13g2_antennanp ANTENNA_20 (.A(net22));
 sg13g2_antennanp ANTENNA_21 (.A(net23));
 sg13g2_antennanp ANTENNA_22 (.A(net23));
 sg13g2_antennanp ANTENNA_23 (.A(net24));
 sg13g2_antennanp ANTENNA_24 (.A(net24));
 sg13g2_antennanp ANTENNA_25 (.A(net403));
 sg13g2_antennanp ANTENNA_26 (.A(net403));
 sg13g2_antennanp ANTENNA_27 (.A(net403));
 sg13g2_antennanp ANTENNA_28 (.A(net403));
 sg13g2_antennanp ANTENNA_29 (.A(net403));
 sg13g2_antennanp ANTENNA_30 (.A(net403));
 sg13g2_antennanp ANTENNA_31 (.A(net403));
 sg13g2_antennanp ANTENNA_32 (.A(net403));
 sg13g2_antennanp ANTENNA_33 (.A(net447));
 sg13g2_antennanp ANTENNA_34 (.A(net447));
 sg13g2_antennanp ANTENNA_35 (.A(net447));
 sg13g2_antennanp ANTENNA_36 (.A(net447));
 sg13g2_antennanp ANTENNA_37 (.A(net447));
 sg13g2_antennanp ANTENNA_38 (.A(net447));
 sg13g2_antennanp ANTENNA_39 (.A(net447));
 sg13g2_antennanp ANTENNA_40 (.A(net447));
 sg13g2_antennanp ANTENNA_41 (.A(net447));
 sg13g2_antennanp ANTENNA_42 (.A(net447));
 sg13g2_antennanp ANTENNA_43 (.A(net447));
 sg13g2_antennanp ANTENNA_44 (.A(net447));
 sg13g2_antennanp ANTENNA_45 (.A(net447));
 sg13g2_antennanp ANTENNA_46 (.A(net447));
 sg13g2_antennanp ANTENNA_47 (.A(net447));
 sg13g2_antennanp ANTENNA_48 (.A(net447));
 sg13g2_antennanp ANTENNA_49 (.A(net447));
 sg13g2_antennanp ANTENNA_50 (.A(net447));
 sg13g2_antennanp ANTENNA_51 (.A(net447));
 sg13g2_antennanp ANTENNA_52 (.A(net447));
 sg13g2_antennanp ANTENNA_53 (.A(net447));
 sg13g2_antennanp ANTENNA_54 (.A(net447));
 sg13g2_antennanp ANTENNA_55 (.A(net447));
 sg13g2_antennanp ANTENNA_56 (.A(_00383_));
 sg13g2_antennanp ANTENNA_57 (.A(_00422_));
 sg13g2_antennanp ANTENNA_58 (.A(_02067_));
 sg13g2_antennanp ANTENNA_59 (.A(_02067_));
 sg13g2_antennanp ANTENNA_60 (.A(_02400_));
 sg13g2_antennanp ANTENNA_61 (.A(_02400_));
 sg13g2_antennanp ANTENNA_62 (.A(_05057_));
 sg13g2_antennanp ANTENNA_63 (.A(_05057_));
 sg13g2_antennanp ANTENNA_64 (.A(_05057_));
 sg13g2_antennanp ANTENNA_65 (.A(_05057_));
 sg13g2_antennanp ANTENNA_66 (.A(_05057_));
 sg13g2_antennanp ANTENNA_67 (.A(_05057_));
 sg13g2_antennanp ANTENNA_68 (.A(clk));
 sg13g2_antennanp ANTENNA_69 (.A(clk));
 sg13g2_antennanp ANTENNA_70 (.A(net22));
 sg13g2_antennanp ANTENNA_71 (.A(net22));
 sg13g2_antennanp ANTENNA_72 (.A(net23));
 sg13g2_antennanp ANTENNA_73 (.A(net23));
 sg13g2_antennanp ANTENNA_74 (.A(net24));
 sg13g2_antennanp ANTENNA_75 (.A(net24));
 sg13g2_antennanp ANTENNA_76 (.A(net447));
 sg13g2_antennanp ANTENNA_77 (.A(net447));
 sg13g2_antennanp ANTENNA_78 (.A(net447));
 sg13g2_antennanp ANTENNA_79 (.A(net447));
 sg13g2_antennanp ANTENNA_80 (.A(net447));
 sg13g2_antennanp ANTENNA_81 (.A(net447));
 sg13g2_antennanp ANTENNA_82 (.A(net447));
 sg13g2_antennanp ANTENNA_83 (.A(net447));
 sg13g2_antennanp ANTENNA_84 (.A(net447));
 sg13g2_antennanp ANTENNA_85 (.A(_00383_));
 sg13g2_antennanp ANTENNA_86 (.A(_00422_));
 sg13g2_antennanp ANTENNA_87 (.A(_02067_));
 sg13g2_antennanp ANTENNA_88 (.A(_02067_));
 sg13g2_antennanp ANTENNA_89 (.A(_02400_));
 sg13g2_antennanp ANTENNA_90 (.A(_02400_));
 sg13g2_antennanp ANTENNA_91 (.A(_05057_));
 sg13g2_antennanp ANTENNA_92 (.A(_05057_));
 sg13g2_antennanp ANTENNA_93 (.A(_05057_));
 sg13g2_antennanp ANTENNA_94 (.A(_05057_));
 sg13g2_antennanp ANTENNA_95 (.A(_05057_));
 sg13g2_antennanp ANTENNA_96 (.A(_05057_));
 sg13g2_antennanp ANTENNA_97 (.A(clk));
 sg13g2_antennanp ANTENNA_98 (.A(clk));
 sg13g2_antennanp ANTENNA_99 (.A(net22));
 sg13g2_antennanp ANTENNA_100 (.A(net22));
 sg13g2_antennanp ANTENNA_101 (.A(net23));
 sg13g2_antennanp ANTENNA_102 (.A(net23));
 sg13g2_antennanp ANTENNA_103 (.A(net24));
 sg13g2_antennanp ANTENNA_104 (.A(net24));
 sg13g2_antennanp ANTENNA_105 (.A(_00383_));
 sg13g2_antennanp ANTENNA_106 (.A(_00422_));
 sg13g2_antennanp ANTENNA_107 (.A(_02067_));
 sg13g2_antennanp ANTENNA_108 (.A(_02067_));
 sg13g2_antennanp ANTENNA_109 (.A(_02400_));
 sg13g2_antennanp ANTENNA_110 (.A(_02400_));
 sg13g2_antennanp ANTENNA_111 (.A(_05057_));
 sg13g2_antennanp ANTENNA_112 (.A(_05057_));
 sg13g2_antennanp ANTENNA_113 (.A(_05057_));
 sg13g2_antennanp ANTENNA_114 (.A(_05057_));
 sg13g2_antennanp ANTENNA_115 (.A(_05057_));
 sg13g2_antennanp ANTENNA_116 (.A(_05057_));
 sg13g2_antennanp ANTENNA_117 (.A(clk));
 sg13g2_antennanp ANTENNA_118 (.A(clk));
 sg13g2_antennanp ANTENNA_119 (.A(net22));
 sg13g2_antennanp ANTENNA_120 (.A(net22));
 sg13g2_antennanp ANTENNA_121 (.A(net23));
 sg13g2_antennanp ANTENNA_122 (.A(net23));
 sg13g2_antennanp ANTENNA_123 (.A(net24));
 sg13g2_antennanp ANTENNA_124 (.A(net24));
 sg13g2_antennanp ANTENNA_125 (.A(_00383_));
 sg13g2_antennanp ANTENNA_126 (.A(_00422_));
 sg13g2_antennanp ANTENNA_127 (.A(_02067_));
 sg13g2_antennanp ANTENNA_128 (.A(_02067_));
 sg13g2_antennanp ANTENNA_129 (.A(_02400_));
 sg13g2_antennanp ANTENNA_130 (.A(_02400_));
 sg13g2_antennanp ANTENNA_131 (.A(_05057_));
 sg13g2_antennanp ANTENNA_132 (.A(_05057_));
 sg13g2_antennanp ANTENNA_133 (.A(_05057_));
 sg13g2_antennanp ANTENNA_134 (.A(_05057_));
 sg13g2_antennanp ANTENNA_135 (.A(_05057_));
 sg13g2_antennanp ANTENNA_136 (.A(_05057_));
 sg13g2_antennanp ANTENNA_137 (.A(clk));
 sg13g2_antennanp ANTENNA_138 (.A(clk));
 sg13g2_antennanp ANTENNA_139 (.A(net22));
 sg13g2_antennanp ANTENNA_140 (.A(net22));
 sg13g2_antennanp ANTENNA_141 (.A(net23));
 sg13g2_antennanp ANTENNA_142 (.A(net23));
 sg13g2_antennanp ANTENNA_143 (.A(net24));
 sg13g2_antennanp ANTENNA_144 (.A(net24));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_945 ();
 sg13g2_decap_8 FILLER_0_952 ();
 sg13g2_decap_8 FILLER_0_959 ();
 sg13g2_decap_8 FILLER_0_966 ();
 sg13g2_decap_8 FILLER_0_973 ();
 sg13g2_decap_8 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_987 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_decap_8 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1008 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1022 ();
 sg13g2_decap_8 FILLER_0_1029 ();
 sg13g2_decap_8 FILLER_0_1036 ();
 sg13g2_decap_8 FILLER_0_1043 ();
 sg13g2_decap_8 FILLER_0_1050 ();
 sg13g2_fill_2 FILLER_0_1057 ();
 sg13g2_fill_2 FILLER_0_1063 ();
 sg13g2_decap_8 FILLER_0_1068 ();
 sg13g2_decap_8 FILLER_0_1075 ();
 sg13g2_decap_8 FILLER_0_1082 ();
 sg13g2_decap_8 FILLER_0_1089 ();
 sg13g2_decap_8 FILLER_0_1096 ();
 sg13g2_decap_8 FILLER_0_1103 ();
 sg13g2_decap_8 FILLER_0_1110 ();
 sg13g2_decap_8 FILLER_0_1117 ();
 sg13g2_decap_8 FILLER_0_1124 ();
 sg13g2_decap_8 FILLER_0_1131 ();
 sg13g2_decap_8 FILLER_0_1138 ();
 sg13g2_decap_8 FILLER_0_1145 ();
 sg13g2_decap_8 FILLER_0_1152 ();
 sg13g2_decap_8 FILLER_0_1159 ();
 sg13g2_decap_8 FILLER_0_1166 ();
 sg13g2_decap_8 FILLER_0_1173 ();
 sg13g2_decap_8 FILLER_0_1180 ();
 sg13g2_decap_8 FILLER_0_1187 ();
 sg13g2_decap_8 FILLER_0_1194 ();
 sg13g2_decap_8 FILLER_0_1201 ();
 sg13g2_decap_8 FILLER_0_1208 ();
 sg13g2_decap_8 FILLER_0_1215 ();
 sg13g2_decap_8 FILLER_0_1222 ();
 sg13g2_decap_8 FILLER_0_1229 ();
 sg13g2_decap_8 FILLER_0_1236 ();
 sg13g2_decap_8 FILLER_0_1243 ();
 sg13g2_decap_8 FILLER_0_1250 ();
 sg13g2_decap_8 FILLER_0_1257 ();
 sg13g2_decap_8 FILLER_0_1264 ();
 sg13g2_decap_8 FILLER_0_1271 ();
 sg13g2_decap_8 FILLER_0_1278 ();
 sg13g2_decap_8 FILLER_0_1285 ();
 sg13g2_decap_8 FILLER_0_1292 ();
 sg13g2_decap_8 FILLER_0_1299 ();
 sg13g2_decap_8 FILLER_0_1306 ();
 sg13g2_decap_8 FILLER_0_1313 ();
 sg13g2_decap_4 FILLER_0_1320 ();
 sg13g2_fill_2 FILLER_0_1324 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_94 ();
 sg13g2_decap_8 FILLER_1_101 ();
 sg13g2_decap_8 FILLER_1_108 ();
 sg13g2_decap_8 FILLER_1_115 ();
 sg13g2_decap_8 FILLER_1_122 ();
 sg13g2_decap_8 FILLER_1_129 ();
 sg13g2_decap_8 FILLER_1_136 ();
 sg13g2_decap_8 FILLER_1_143 ();
 sg13g2_decap_8 FILLER_1_150 ();
 sg13g2_decap_8 FILLER_1_157 ();
 sg13g2_decap_8 FILLER_1_164 ();
 sg13g2_decap_8 FILLER_1_171 ();
 sg13g2_decap_4 FILLER_1_178 ();
 sg13g2_fill_1 FILLER_1_182 ();
 sg13g2_fill_1 FILLER_1_195 ();
 sg13g2_fill_1 FILLER_1_208 ();
 sg13g2_decap_8 FILLER_1_212 ();
 sg13g2_decap_8 FILLER_1_219 ();
 sg13g2_decap_8 FILLER_1_226 ();
 sg13g2_decap_4 FILLER_1_233 ();
 sg13g2_decap_8 FILLER_1_249 ();
 sg13g2_decap_8 FILLER_1_256 ();
 sg13g2_decap_8 FILLER_1_263 ();
 sg13g2_decap_8 FILLER_1_270 ();
 sg13g2_decap_8 FILLER_1_277 ();
 sg13g2_decap_8 FILLER_1_284 ();
 sg13g2_decap_8 FILLER_1_291 ();
 sg13g2_decap_8 FILLER_1_298 ();
 sg13g2_decap_8 FILLER_1_305 ();
 sg13g2_decap_8 FILLER_1_312 ();
 sg13g2_decap_8 FILLER_1_319 ();
 sg13g2_decap_8 FILLER_1_326 ();
 sg13g2_decap_8 FILLER_1_333 ();
 sg13g2_decap_8 FILLER_1_340 ();
 sg13g2_decap_8 FILLER_1_347 ();
 sg13g2_decap_8 FILLER_1_354 ();
 sg13g2_decap_8 FILLER_1_361 ();
 sg13g2_decap_8 FILLER_1_368 ();
 sg13g2_decap_4 FILLER_1_375 ();
 sg13g2_fill_2 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_fill_1 FILLER_1_430 ();
 sg13g2_decap_8 FILLER_1_435 ();
 sg13g2_decap_4 FILLER_1_442 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_509 ();
 sg13g2_fill_1 FILLER_1_516 ();
 sg13g2_fill_1 FILLER_1_522 ();
 sg13g2_decap_8 FILLER_1_535 ();
 sg13g2_decap_8 FILLER_1_542 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_4 FILLER_1_574 ();
 sg13g2_fill_2 FILLER_1_578 ();
 sg13g2_decap_8 FILLER_1_606 ();
 sg13g2_decap_8 FILLER_1_613 ();
 sg13g2_decap_8 FILLER_1_620 ();
 sg13g2_decap_8 FILLER_1_627 ();
 sg13g2_fill_1 FILLER_1_634 ();
 sg13g2_decap_8 FILLER_1_643 ();
 sg13g2_decap_8 FILLER_1_650 ();
 sg13g2_decap_8 FILLER_1_657 ();
 sg13g2_decap_8 FILLER_1_664 ();
 sg13g2_decap_8 FILLER_1_671 ();
 sg13g2_fill_2 FILLER_1_678 ();
 sg13g2_decap_8 FILLER_1_706 ();
 sg13g2_decap_8 FILLER_1_713 ();
 sg13g2_decap_8 FILLER_1_720 ();
 sg13g2_decap_8 FILLER_1_727 ();
 sg13g2_decap_8 FILLER_1_734 ();
 sg13g2_decap_8 FILLER_1_741 ();
 sg13g2_decap_4 FILLER_1_748 ();
 sg13g2_fill_2 FILLER_1_752 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_4 FILLER_1_826 ();
 sg13g2_fill_2 FILLER_1_830 ();
 sg13g2_decap_8 FILLER_1_858 ();
 sg13g2_decap_8 FILLER_1_865 ();
 sg13g2_decap_8 FILLER_1_905 ();
 sg13g2_fill_2 FILLER_1_912 ();
 sg13g2_fill_1 FILLER_1_914 ();
 sg13g2_decap_4 FILLER_1_949 ();
 sg13g2_fill_2 FILLER_1_953 ();
 sg13g2_decap_8 FILLER_1_959 ();
 sg13g2_decap_8 FILLER_1_966 ();
 sg13g2_decap_8 FILLER_1_973 ();
 sg13g2_decap_8 FILLER_1_980 ();
 sg13g2_decap_4 FILLER_1_987 ();
 sg13g2_fill_2 FILLER_1_991 ();
 sg13g2_decap_8 FILLER_1_997 ();
 sg13g2_decap_4 FILLER_1_1004 ();
 sg13g2_decap_8 FILLER_1_1034 ();
 sg13g2_decap_8 FILLER_1_1041 ();
 sg13g2_decap_4 FILLER_1_1048 ();
 sg13g2_fill_2 FILLER_1_1052 ();
 sg13g2_decap_8 FILLER_1_1080 ();
 sg13g2_decap_8 FILLER_1_1087 ();
 sg13g2_fill_1 FILLER_1_1094 ();
 sg13g2_decap_8 FILLER_1_1099 ();
 sg13g2_decap_8 FILLER_1_1106 ();
 sg13g2_fill_2 FILLER_1_1113 ();
 sg13g2_fill_1 FILLER_1_1115 ();
 sg13g2_decap_8 FILLER_1_1120 ();
 sg13g2_decap_8 FILLER_1_1131 ();
 sg13g2_decap_4 FILLER_1_1138 ();
 sg13g2_fill_1 FILLER_1_1142 ();
 sg13g2_decap_8 FILLER_1_1147 ();
 sg13g2_decap_8 FILLER_1_1158 ();
 sg13g2_decap_4 FILLER_1_1165 ();
 sg13g2_decap_8 FILLER_1_1173 ();
 sg13g2_decap_8 FILLER_1_1184 ();
 sg13g2_decap_8 FILLER_1_1191 ();
 sg13g2_decap_8 FILLER_1_1198 ();
 sg13g2_decap_8 FILLER_1_1205 ();
 sg13g2_decap_8 FILLER_1_1212 ();
 sg13g2_decap_8 FILLER_1_1219 ();
 sg13g2_decap_8 FILLER_1_1226 ();
 sg13g2_decap_8 FILLER_1_1233 ();
 sg13g2_decap_8 FILLER_1_1240 ();
 sg13g2_decap_8 FILLER_1_1247 ();
 sg13g2_decap_8 FILLER_1_1254 ();
 sg13g2_decap_8 FILLER_1_1261 ();
 sg13g2_decap_8 FILLER_1_1268 ();
 sg13g2_decap_8 FILLER_1_1275 ();
 sg13g2_decap_8 FILLER_1_1282 ();
 sg13g2_decap_8 FILLER_1_1289 ();
 sg13g2_decap_8 FILLER_1_1296 ();
 sg13g2_decap_8 FILLER_1_1303 ();
 sg13g2_decap_8 FILLER_1_1310 ();
 sg13g2_decap_8 FILLER_1_1317 ();
 sg13g2_fill_2 FILLER_1_1324 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_4 FILLER_2_56 ();
 sg13g2_fill_1 FILLER_2_60 ();
 sg13g2_decap_4 FILLER_2_69 ();
 sg13g2_fill_2 FILLER_2_73 ();
 sg13g2_decap_4 FILLER_2_90 ();
 sg13g2_fill_1 FILLER_2_103 ();
 sg13g2_fill_1 FILLER_2_108 ();
 sg13g2_decap_8 FILLER_2_117 ();
 sg13g2_fill_1 FILLER_2_124 ();
 sg13g2_decap_8 FILLER_2_134 ();
 sg13g2_decap_4 FILLER_2_141 ();
 sg13g2_fill_1 FILLER_2_145 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_fill_2 FILLER_2_178 ();
 sg13g2_fill_1 FILLER_2_180 ();
 sg13g2_fill_1 FILLER_2_194 ();
 sg13g2_fill_1 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_fill_2 FILLER_2_221 ();
 sg13g2_fill_1 FILLER_2_223 ();
 sg13g2_fill_2 FILLER_2_228 ();
 sg13g2_fill_1 FILLER_2_230 ();
 sg13g2_decap_8 FILLER_2_244 ();
 sg13g2_fill_1 FILLER_2_260 ();
 sg13g2_decap_4 FILLER_2_266 ();
 sg13g2_decap_4 FILLER_2_282 ();
 sg13g2_fill_1 FILLER_2_286 ();
 sg13g2_decap_4 FILLER_2_291 ();
 sg13g2_fill_1 FILLER_2_295 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_4 FILLER_2_378 ();
 sg13g2_decap_4 FILLER_2_421 ();
 sg13g2_decap_8 FILLER_2_460 ();
 sg13g2_decap_8 FILLER_2_467 ();
 sg13g2_decap_8 FILLER_2_474 ();
 sg13g2_decap_8 FILLER_2_481 ();
 sg13g2_fill_2 FILLER_2_492 ();
 sg13g2_decap_4 FILLER_2_576 ();
 sg13g2_fill_2 FILLER_2_580 ();
 sg13g2_fill_1 FILLER_2_631 ();
 sg13g2_fill_1 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_649 ();
 sg13g2_decap_8 FILLER_2_656 ();
 sg13g2_decap_8 FILLER_2_663 ();
 sg13g2_decap_8 FILLER_2_670 ();
 sg13g2_fill_1 FILLER_2_677 ();
 sg13g2_decap_8 FILLER_2_682 ();
 sg13g2_fill_1 FILLER_2_689 ();
 sg13g2_decap_8 FILLER_2_694 ();
 sg13g2_fill_2 FILLER_2_701 ();
 sg13g2_fill_1 FILLER_2_707 ();
 sg13g2_decap_4 FILLER_2_723 ();
 sg13g2_fill_2 FILLER_2_757 ();
 sg13g2_decap_8 FILLER_2_789 ();
 sg13g2_decap_8 FILLER_2_796 ();
 sg13g2_decap_8 FILLER_2_829 ();
 sg13g2_fill_1 FILLER_2_836 ();
 sg13g2_decap_8 FILLER_2_841 ();
 sg13g2_fill_2 FILLER_2_848 ();
 sg13g2_decap_8 FILLER_2_853 ();
 sg13g2_decap_8 FILLER_2_860 ();
 sg13g2_decap_8 FILLER_2_867 ();
 sg13g2_decap_4 FILLER_2_874 ();
 sg13g2_decap_8 FILLER_2_886 ();
 sg13g2_decap_8 FILLER_2_893 ();
 sg13g2_decap_8 FILLER_2_900 ();
 sg13g2_decap_8 FILLER_2_907 ();
 sg13g2_fill_2 FILLER_2_914 ();
 sg13g2_fill_2 FILLER_2_928 ();
 sg13g2_fill_2 FILLER_2_934 ();
 sg13g2_fill_1 FILLER_2_936 ();
 sg13g2_fill_1 FILLER_2_945 ();
 sg13g2_fill_2 FILLER_2_972 ();
 sg13g2_fill_1 FILLER_2_974 ();
 sg13g2_fill_2 FILLER_2_1005 ();
 sg13g2_fill_1 FILLER_2_1007 ();
 sg13g2_decap_4 FILLER_2_1012 ();
 sg13g2_fill_2 FILLER_2_1016 ();
 sg13g2_decap_8 FILLER_2_1026 ();
 sg13g2_decap_4 FILLER_2_1033 ();
 sg13g2_fill_1 FILLER_2_1037 ();
 sg13g2_decap_8 FILLER_2_1042 ();
 sg13g2_decap_8 FILLER_2_1049 ();
 sg13g2_decap_8 FILLER_2_1056 ();
 sg13g2_decap_8 FILLER_2_1067 ();
 sg13g2_decap_8 FILLER_2_1074 ();
 sg13g2_decap_4 FILLER_2_1081 ();
 sg13g2_fill_1 FILLER_2_1085 ();
 sg13g2_decap_8 FILLER_2_1202 ();
 sg13g2_decap_8 FILLER_2_1209 ();
 sg13g2_decap_8 FILLER_2_1216 ();
 sg13g2_decap_8 FILLER_2_1223 ();
 sg13g2_decap_8 FILLER_2_1230 ();
 sg13g2_decap_8 FILLER_2_1237 ();
 sg13g2_decap_8 FILLER_2_1244 ();
 sg13g2_decap_8 FILLER_2_1251 ();
 sg13g2_decap_8 FILLER_2_1258 ();
 sg13g2_decap_8 FILLER_2_1265 ();
 sg13g2_decap_8 FILLER_2_1272 ();
 sg13g2_decap_8 FILLER_2_1279 ();
 sg13g2_decap_8 FILLER_2_1286 ();
 sg13g2_decap_8 FILLER_2_1293 ();
 sg13g2_decap_8 FILLER_2_1300 ();
 sg13g2_decap_8 FILLER_2_1307 ();
 sg13g2_decap_8 FILLER_2_1314 ();
 sg13g2_decap_4 FILLER_2_1321 ();
 sg13g2_fill_1 FILLER_2_1325 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_4 FILLER_3_49 ();
 sg13g2_fill_2 FILLER_3_53 ();
 sg13g2_fill_1 FILLER_3_66 ();
 sg13g2_decap_4 FILLER_3_87 ();
 sg13g2_decap_8 FILLER_3_96 ();
 sg13g2_decap_4 FILLER_3_103 ();
 sg13g2_fill_2 FILLER_3_112 ();
 sg13g2_fill_1 FILLER_3_114 ();
 sg13g2_fill_2 FILLER_3_119 ();
 sg13g2_fill_1 FILLER_3_121 ();
 sg13g2_decap_4 FILLER_3_142 ();
 sg13g2_fill_1 FILLER_3_154 ();
 sg13g2_decap_4 FILLER_3_159 ();
 sg13g2_decap_8 FILLER_3_173 ();
 sg13g2_decap_4 FILLER_3_180 ();
 sg13g2_fill_2 FILLER_3_184 ();
 sg13g2_fill_1 FILLER_3_214 ();
 sg13g2_decap_4 FILLER_3_225 ();
 sg13g2_fill_2 FILLER_3_229 ();
 sg13g2_decap_8 FILLER_3_265 ();
 sg13g2_decap_4 FILLER_3_272 ();
 sg13g2_fill_1 FILLER_3_276 ();
 sg13g2_decap_8 FILLER_3_281 ();
 sg13g2_fill_2 FILLER_3_288 ();
 sg13g2_fill_1 FILLER_3_290 ();
 sg13g2_decap_4 FILLER_3_305 ();
 sg13g2_fill_2 FILLER_3_314 ();
 sg13g2_decap_8 FILLER_3_330 ();
 sg13g2_decap_8 FILLER_3_337 ();
 sg13g2_decap_8 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_351 ();
 sg13g2_decap_8 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_fill_2 FILLER_3_393 ();
 sg13g2_fill_1 FILLER_3_395 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_3_414 ();
 sg13g2_fill_2 FILLER_3_421 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_4 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_443 ();
 sg13g2_decap_8 FILLER_3_450 ();
 sg13g2_decap_8 FILLER_3_457 ();
 sg13g2_decap_8 FILLER_3_464 ();
 sg13g2_decap_8 FILLER_3_471 ();
 sg13g2_decap_8 FILLER_3_487 ();
 sg13g2_decap_8 FILLER_3_494 ();
 sg13g2_fill_2 FILLER_3_501 ();
 sg13g2_fill_1 FILLER_3_503 ();
 sg13g2_decap_8 FILLER_3_508 ();
 sg13g2_decap_8 FILLER_3_515 ();
 sg13g2_decap_8 FILLER_3_526 ();
 sg13g2_decap_4 FILLER_3_533 ();
 sg13g2_fill_1 FILLER_3_563 ();
 sg13g2_decap_8 FILLER_3_568 ();
 sg13g2_decap_8 FILLER_3_575 ();
 sg13g2_decap_8 FILLER_3_582 ();
 sg13g2_decap_4 FILLER_3_589 ();
 sg13g2_decap_4 FILLER_3_597 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_4 FILLER_3_616 ();
 sg13g2_fill_1 FILLER_3_620 ();
 sg13g2_fill_2 FILLER_3_647 ();
 sg13g2_fill_1 FILLER_3_649 ();
 sg13g2_decap_4 FILLER_3_654 ();
 sg13g2_decap_4 FILLER_3_662 ();
 sg13g2_fill_2 FILLER_3_674 ();
 sg13g2_decap_8 FILLER_3_684 ();
 sg13g2_decap_8 FILLER_3_691 ();
 sg13g2_fill_2 FILLER_3_698 ();
 sg13g2_fill_1 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_743 ();
 sg13g2_fill_1 FILLER_3_750 ();
 sg13g2_fill_1 FILLER_3_755 ();
 sg13g2_decap_8 FILLER_3_760 ();
 sg13g2_fill_2 FILLER_3_767 ();
 sg13g2_fill_1 FILLER_3_769 ();
 sg13g2_decap_8 FILLER_3_800 ();
 sg13g2_fill_2 FILLER_3_807 ();
 sg13g2_decap_8 FILLER_3_813 ();
 sg13g2_decap_4 FILLER_3_820 ();
 sg13g2_fill_1 FILLER_3_824 ();
 sg13g2_fill_1 FILLER_3_829 ();
 sg13g2_fill_2 FILLER_3_834 ();
 sg13g2_fill_1 FILLER_3_844 ();
 sg13g2_fill_2 FILLER_3_871 ();
 sg13g2_decap_8 FILLER_3_879 ();
 sg13g2_decap_8 FILLER_3_886 ();
 sg13g2_decap_8 FILLER_3_898 ();
 sg13g2_fill_2 FILLER_3_905 ();
 sg13g2_decap_8 FILLER_3_919 ();
 sg13g2_fill_1 FILLER_3_926 ();
 sg13g2_fill_1 FILLER_3_935 ();
 sg13g2_decap_8 FILLER_3_941 ();
 sg13g2_decap_8 FILLER_3_948 ();
 sg13g2_decap_8 FILLER_3_955 ();
 sg13g2_decap_8 FILLER_3_962 ();
 sg13g2_decap_8 FILLER_3_969 ();
 sg13g2_decap_4 FILLER_3_976 ();
 sg13g2_fill_2 FILLER_3_980 ();
 sg13g2_decap_8 FILLER_3_986 ();
 sg13g2_fill_2 FILLER_3_993 ();
 sg13g2_decap_4 FILLER_3_1003 ();
 sg13g2_decap_8 FILLER_3_1019 ();
 sg13g2_decap_4 FILLER_3_1026 ();
 sg13g2_fill_1 FILLER_3_1030 ();
 sg13g2_decap_8 FILLER_3_1061 ();
 sg13g2_decap_8 FILLER_3_1068 ();
 sg13g2_decap_8 FILLER_3_1075 ();
 sg13g2_decap_8 FILLER_3_1082 ();
 sg13g2_fill_1 FILLER_3_1089 ();
 sg13g2_decap_8 FILLER_3_1094 ();
 sg13g2_fill_2 FILLER_3_1101 ();
 sg13g2_fill_1 FILLER_3_1115 ();
 sg13g2_decap_8 FILLER_3_1120 ();
 sg13g2_decap_8 FILLER_3_1127 ();
 sg13g2_decap_4 FILLER_3_1134 ();
 sg13g2_fill_2 FILLER_3_1138 ();
 sg13g2_decap_8 FILLER_3_1151 ();
 sg13g2_decap_8 FILLER_3_1158 ();
 sg13g2_decap_8 FILLER_3_1165 ();
 sg13g2_decap_8 FILLER_3_1180 ();
 sg13g2_decap_8 FILLER_3_1187 ();
 sg13g2_decap_8 FILLER_3_1194 ();
 sg13g2_decap_8 FILLER_3_1201 ();
 sg13g2_decap_8 FILLER_3_1208 ();
 sg13g2_decap_8 FILLER_3_1215 ();
 sg13g2_decap_8 FILLER_3_1222 ();
 sg13g2_decap_8 FILLER_3_1229 ();
 sg13g2_decap_8 FILLER_3_1236 ();
 sg13g2_decap_8 FILLER_3_1243 ();
 sg13g2_decap_8 FILLER_3_1250 ();
 sg13g2_decap_8 FILLER_3_1257 ();
 sg13g2_decap_8 FILLER_3_1264 ();
 sg13g2_decap_8 FILLER_3_1271 ();
 sg13g2_decap_8 FILLER_3_1278 ();
 sg13g2_decap_8 FILLER_3_1285 ();
 sg13g2_decap_8 FILLER_3_1292 ();
 sg13g2_decap_8 FILLER_3_1299 ();
 sg13g2_decap_8 FILLER_3_1306 ();
 sg13g2_decap_8 FILLER_3_1313 ();
 sg13g2_decap_4 FILLER_3_1320 ();
 sg13g2_fill_2 FILLER_3_1324 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_4 FILLER_4_49 ();
 sg13g2_decap_4 FILLER_4_58 ();
 sg13g2_fill_2 FILLER_4_62 ();
 sg13g2_fill_1 FILLER_4_71 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_fill_2 FILLER_4_112 ();
 sg13g2_fill_1 FILLER_4_114 ();
 sg13g2_fill_1 FILLER_4_130 ();
 sg13g2_fill_2 FILLER_4_159 ();
 sg13g2_fill_1 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_170 ();
 sg13g2_fill_1 FILLER_4_177 ();
 sg13g2_decap_8 FILLER_4_186 ();
 sg13g2_decap_8 FILLER_4_193 ();
 sg13g2_decap_8 FILLER_4_200 ();
 sg13g2_decap_8 FILLER_4_207 ();
 sg13g2_decap_8 FILLER_4_214 ();
 sg13g2_decap_8 FILLER_4_221 ();
 sg13g2_decap_8 FILLER_4_228 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_4 FILLER_4_273 ();
 sg13g2_fill_1 FILLER_4_277 ();
 sg13g2_decap_4 FILLER_4_288 ();
 sg13g2_decap_4 FILLER_4_313 ();
 sg13g2_fill_1 FILLER_4_317 ();
 sg13g2_fill_2 FILLER_4_333 ();
 sg13g2_fill_1 FILLER_4_335 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_fill_1 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_355 ();
 sg13g2_decap_8 FILLER_4_362 ();
 sg13g2_decap_4 FILLER_4_369 ();
 sg13g2_fill_2 FILLER_4_373 ();
 sg13g2_fill_1 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_411 ();
 sg13g2_decap_8 FILLER_4_418 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_4_443 ();
 sg13g2_decap_8 FILLER_4_450 ();
 sg13g2_decap_8 FILLER_4_457 ();
 sg13g2_decap_8 FILLER_4_485 ();
 sg13g2_decap_8 FILLER_4_492 ();
 sg13g2_decap_8 FILLER_4_499 ();
 sg13g2_decap_8 FILLER_4_506 ();
 sg13g2_decap_8 FILLER_4_513 ();
 sg13g2_decap_8 FILLER_4_520 ();
 sg13g2_decap_8 FILLER_4_527 ();
 sg13g2_decap_8 FILLER_4_534 ();
 sg13g2_decap_8 FILLER_4_541 ();
 sg13g2_fill_2 FILLER_4_548 ();
 sg13g2_fill_1 FILLER_4_550 ();
 sg13g2_decap_8 FILLER_4_556 ();
 sg13g2_decap_8 FILLER_4_563 ();
 sg13g2_decap_8 FILLER_4_570 ();
 sg13g2_decap_8 FILLER_4_577 ();
 sg13g2_decap_8 FILLER_4_584 ();
 sg13g2_decap_8 FILLER_4_591 ();
 sg13g2_fill_2 FILLER_4_598 ();
 sg13g2_fill_1 FILLER_4_600 ();
 sg13g2_decap_4 FILLER_4_609 ();
 sg13g2_fill_2 FILLER_4_613 ();
 sg13g2_fill_2 FILLER_4_620 ();
 sg13g2_fill_1 FILLER_4_622 ();
 sg13g2_decap_8 FILLER_4_628 ();
 sg13g2_decap_4 FILLER_4_635 ();
 sg13g2_fill_2 FILLER_4_639 ();
 sg13g2_fill_2 FILLER_4_647 ();
 sg13g2_decap_8 FILLER_4_684 ();
 sg13g2_decap_8 FILLER_4_691 ();
 sg13g2_decap_8 FILLER_4_698 ();
 sg13g2_decap_4 FILLER_4_705 ();
 sg13g2_fill_1 FILLER_4_709 ();
 sg13g2_fill_1 FILLER_4_716 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_4 FILLER_4_761 ();
 sg13g2_fill_2 FILLER_4_765 ();
 sg13g2_decap_8 FILLER_4_775 ();
 sg13g2_decap_8 FILLER_4_782 ();
 sg13g2_fill_1 FILLER_4_789 ();
 sg13g2_decap_8 FILLER_4_793 ();
 sg13g2_fill_1 FILLER_4_800 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_fill_1 FILLER_4_819 ();
 sg13g2_decap_4 FILLER_4_832 ();
 sg13g2_fill_1 FILLER_4_836 ();
 sg13g2_decap_4 FILLER_4_841 ();
 sg13g2_decap_4 FILLER_4_853 ();
 sg13g2_fill_1 FILLER_4_857 ();
 sg13g2_fill_2 FILLER_4_871 ();
 sg13g2_decap_4 FILLER_4_877 ();
 sg13g2_fill_2 FILLER_4_885 ();
 sg13g2_fill_1 FILLER_4_887 ();
 sg13g2_decap_8 FILLER_4_892 ();
 sg13g2_fill_2 FILLER_4_899 ();
 sg13g2_fill_1 FILLER_4_906 ();
 sg13g2_decap_8 FILLER_4_941 ();
 sg13g2_decap_8 FILLER_4_948 ();
 sg13g2_decap_8 FILLER_4_955 ();
 sg13g2_decap_8 FILLER_4_962 ();
 sg13g2_decap_8 FILLER_4_969 ();
 sg13g2_decap_8 FILLER_4_976 ();
 sg13g2_decap_8 FILLER_4_983 ();
 sg13g2_fill_2 FILLER_4_990 ();
 sg13g2_fill_1 FILLER_4_996 ();
 sg13g2_fill_2 FILLER_4_1010 ();
 sg13g2_fill_1 FILLER_4_1012 ();
 sg13g2_fill_2 FILLER_4_1019 ();
 sg13g2_decap_4 FILLER_4_1024 ();
 sg13g2_decap_4 FILLER_4_1032 ();
 sg13g2_decap_4 FILLER_4_1044 ();
 sg13g2_decap_8 FILLER_4_1067 ();
 sg13g2_decap_4 FILLER_4_1074 ();
 sg13g2_fill_1 FILLER_4_1078 ();
 sg13g2_decap_8 FILLER_4_1083 ();
 sg13g2_decap_8 FILLER_4_1090 ();
 sg13g2_decap_8 FILLER_4_1097 ();
 sg13g2_decap_8 FILLER_4_1104 ();
 sg13g2_decap_4 FILLER_4_1111 ();
 sg13g2_fill_1 FILLER_4_1115 ();
 sg13g2_decap_8 FILLER_4_1121 ();
 sg13g2_decap_8 FILLER_4_1128 ();
 sg13g2_decap_4 FILLER_4_1135 ();
 sg13g2_fill_2 FILLER_4_1139 ();
 sg13g2_decap_8 FILLER_4_1147 ();
 sg13g2_decap_8 FILLER_4_1154 ();
 sg13g2_decap_8 FILLER_4_1161 ();
 sg13g2_decap_4 FILLER_4_1168 ();
 sg13g2_fill_2 FILLER_4_1172 ();
 sg13g2_decap_8 FILLER_4_1178 ();
 sg13g2_decap_8 FILLER_4_1185 ();
 sg13g2_decap_8 FILLER_4_1192 ();
 sg13g2_decap_8 FILLER_4_1199 ();
 sg13g2_decap_8 FILLER_4_1206 ();
 sg13g2_decap_8 FILLER_4_1213 ();
 sg13g2_decap_8 FILLER_4_1220 ();
 sg13g2_decap_8 FILLER_4_1227 ();
 sg13g2_decap_8 FILLER_4_1234 ();
 sg13g2_decap_8 FILLER_4_1241 ();
 sg13g2_decap_8 FILLER_4_1248 ();
 sg13g2_decap_8 FILLER_4_1255 ();
 sg13g2_decap_8 FILLER_4_1262 ();
 sg13g2_decap_8 FILLER_4_1269 ();
 sg13g2_decap_8 FILLER_4_1276 ();
 sg13g2_decap_8 FILLER_4_1283 ();
 sg13g2_decap_8 FILLER_4_1290 ();
 sg13g2_decap_8 FILLER_4_1297 ();
 sg13g2_decap_8 FILLER_4_1304 ();
 sg13g2_decap_8 FILLER_4_1311 ();
 sg13g2_decap_8 FILLER_4_1318 ();
 sg13g2_fill_1 FILLER_4_1325 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_fill_1 FILLER_5_56 ();
 sg13g2_fill_1 FILLER_5_65 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_fill_2 FILLER_5_84 ();
 sg13g2_fill_1 FILLER_5_86 ();
 sg13g2_decap_8 FILLER_5_93 ();
 sg13g2_decap_8 FILLER_5_100 ();
 sg13g2_decap_8 FILLER_5_107 ();
 sg13g2_decap_8 FILLER_5_114 ();
 sg13g2_decap_8 FILLER_5_121 ();
 sg13g2_decap_8 FILLER_5_128 ();
 sg13g2_decap_8 FILLER_5_135 ();
 sg13g2_decap_8 FILLER_5_142 ();
 sg13g2_decap_4 FILLER_5_149 ();
 sg13g2_fill_1 FILLER_5_153 ();
 sg13g2_decap_8 FILLER_5_158 ();
 sg13g2_decap_4 FILLER_5_165 ();
 sg13g2_fill_2 FILLER_5_169 ();
 sg13g2_decap_8 FILLER_5_183 ();
 sg13g2_decap_8 FILLER_5_190 ();
 sg13g2_decap_8 FILLER_5_197 ();
 sg13g2_decap_8 FILLER_5_204 ();
 sg13g2_fill_2 FILLER_5_211 ();
 sg13g2_fill_1 FILLER_5_213 ();
 sg13g2_decap_8 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_229 ();
 sg13g2_fill_1 FILLER_5_236 ();
 sg13g2_decap_4 FILLER_5_242 ();
 sg13g2_fill_1 FILLER_5_246 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_fill_2 FILLER_5_266 ();
 sg13g2_fill_2 FILLER_5_286 ();
 sg13g2_fill_1 FILLER_5_288 ();
 sg13g2_fill_2 FILLER_5_294 ();
 sg13g2_fill_1 FILLER_5_296 ();
 sg13g2_decap_8 FILLER_5_302 ();
 sg13g2_decap_4 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_317 ();
 sg13g2_decap_8 FILLER_5_324 ();
 sg13g2_decap_8 FILLER_5_331 ();
 sg13g2_decap_8 FILLER_5_338 ();
 sg13g2_decap_4 FILLER_5_371 ();
 sg13g2_fill_2 FILLER_5_379 ();
 sg13g2_fill_1 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_4 FILLER_5_398 ();
 sg13g2_fill_1 FILLER_5_402 ();
 sg13g2_fill_2 FILLER_5_424 ();
 sg13g2_fill_1 FILLER_5_426 ();
 sg13g2_fill_1 FILLER_5_453 ();
 sg13g2_decap_8 FILLER_5_480 ();
 sg13g2_decap_8 FILLER_5_487 ();
 sg13g2_decap_8 FILLER_5_494 ();
 sg13g2_decap_8 FILLER_5_501 ();
 sg13g2_decap_4 FILLER_5_508 ();
 sg13g2_decap_8 FILLER_5_517 ();
 sg13g2_decap_8 FILLER_5_524 ();
 sg13g2_decap_8 FILLER_5_531 ();
 sg13g2_decap_8 FILLER_5_538 ();
 sg13g2_decap_8 FILLER_5_545 ();
 sg13g2_decap_8 FILLER_5_552 ();
 sg13g2_decap_8 FILLER_5_559 ();
 sg13g2_decap_8 FILLER_5_566 ();
 sg13g2_decap_8 FILLER_5_573 ();
 sg13g2_decap_8 FILLER_5_580 ();
 sg13g2_decap_8 FILLER_5_587 ();
 sg13g2_decap_8 FILLER_5_594 ();
 sg13g2_decap_8 FILLER_5_601 ();
 sg13g2_fill_2 FILLER_5_608 ();
 sg13g2_decap_4 FILLER_5_614 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_fill_2 FILLER_5_700 ();
 sg13g2_fill_1 FILLER_5_702 ();
 sg13g2_decap_8 FILLER_5_715 ();
 sg13g2_decap_8 FILLER_5_722 ();
 sg13g2_decap_8 FILLER_5_729 ();
 sg13g2_decap_8 FILLER_5_736 ();
 sg13g2_decap_8 FILLER_5_743 ();
 sg13g2_decap_8 FILLER_5_750 ();
 sg13g2_decap_4 FILLER_5_757 ();
 sg13g2_fill_2 FILLER_5_761 ();
 sg13g2_decap_8 FILLER_5_767 ();
 sg13g2_decap_8 FILLER_5_774 ();
 sg13g2_decap_8 FILLER_5_781 ();
 sg13g2_decap_8 FILLER_5_788 ();
 sg13g2_decap_8 FILLER_5_795 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_decap_8 FILLER_5_809 ();
 sg13g2_decap_8 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_823 ();
 sg13g2_decap_8 FILLER_5_830 ();
 sg13g2_decap_8 FILLER_5_837 ();
 sg13g2_decap_8 FILLER_5_844 ();
 sg13g2_decap_8 FILLER_5_851 ();
 sg13g2_decap_8 FILLER_5_858 ();
 sg13g2_decap_4 FILLER_5_865 ();
 sg13g2_decap_8 FILLER_5_907 ();
 sg13g2_fill_2 FILLER_5_914 ();
 sg13g2_fill_1 FILLER_5_916 ();
 sg13g2_decap_8 FILLER_5_921 ();
 sg13g2_decap_8 FILLER_5_928 ();
 sg13g2_decap_8 FILLER_5_935 ();
 sg13g2_decap_4 FILLER_5_942 ();
 sg13g2_fill_2 FILLER_5_946 ();
 sg13g2_decap_4 FILLER_5_952 ();
 sg13g2_fill_1 FILLER_5_956 ();
 sg13g2_decap_8 FILLER_5_961 ();
 sg13g2_decap_8 FILLER_5_968 ();
 sg13g2_decap_4 FILLER_5_975 ();
 sg13g2_fill_1 FILLER_5_979 ();
 sg13g2_decap_8 FILLER_5_1006 ();
 sg13g2_decap_8 FILLER_5_1013 ();
 sg13g2_fill_2 FILLER_5_1020 ();
 sg13g2_fill_1 FILLER_5_1022 ();
 sg13g2_decap_8 FILLER_5_1029 ();
 sg13g2_decap_8 FILLER_5_1036 ();
 sg13g2_fill_1 FILLER_5_1055 ();
 sg13g2_fill_2 FILLER_5_1082 ();
 sg13g2_fill_1 FILLER_5_1084 ();
 sg13g2_decap_8 FILLER_5_1090 ();
 sg13g2_decap_4 FILLER_5_1097 ();
 sg13g2_fill_1 FILLER_5_1101 ();
 sg13g2_decap_8 FILLER_5_1117 ();
 sg13g2_decap_8 FILLER_5_1124 ();
 sg13g2_decap_4 FILLER_5_1131 ();
 sg13g2_fill_2 FILLER_5_1135 ();
 sg13g2_decap_8 FILLER_5_1143 ();
 sg13g2_decap_8 FILLER_5_1150 ();
 sg13g2_decap_8 FILLER_5_1157 ();
 sg13g2_decap_4 FILLER_5_1164 ();
 sg13g2_decap_4 FILLER_5_1180 ();
 sg13g2_fill_1 FILLER_5_1184 ();
 sg13g2_decap_8 FILLER_5_1195 ();
 sg13g2_decap_8 FILLER_5_1202 ();
 sg13g2_decap_8 FILLER_5_1209 ();
 sg13g2_decap_8 FILLER_5_1216 ();
 sg13g2_decap_8 FILLER_5_1223 ();
 sg13g2_decap_8 FILLER_5_1230 ();
 sg13g2_decap_8 FILLER_5_1237 ();
 sg13g2_decap_8 FILLER_5_1244 ();
 sg13g2_decap_8 FILLER_5_1251 ();
 sg13g2_decap_8 FILLER_5_1258 ();
 sg13g2_decap_8 FILLER_5_1265 ();
 sg13g2_decap_8 FILLER_5_1272 ();
 sg13g2_decap_8 FILLER_5_1279 ();
 sg13g2_decap_8 FILLER_5_1286 ();
 sg13g2_decap_8 FILLER_5_1293 ();
 sg13g2_decap_8 FILLER_5_1300 ();
 sg13g2_decap_8 FILLER_5_1307 ();
 sg13g2_decap_8 FILLER_5_1314 ();
 sg13g2_decap_4 FILLER_5_1321 ();
 sg13g2_fill_1 FILLER_5_1325 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_4 FILLER_6_54 ();
 sg13g2_fill_2 FILLER_6_62 ();
 sg13g2_decap_4 FILLER_6_68 ();
 sg13g2_decap_4 FILLER_6_91 ();
 sg13g2_fill_2 FILLER_6_95 ();
 sg13g2_decap_4 FILLER_6_101 ();
 sg13g2_fill_2 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_114 ();
 sg13g2_decap_8 FILLER_6_121 ();
 sg13g2_fill_2 FILLER_6_128 ();
 sg13g2_decap_8 FILLER_6_135 ();
 sg13g2_decap_8 FILLER_6_142 ();
 sg13g2_decap_4 FILLER_6_149 ();
 sg13g2_fill_1 FILLER_6_153 ();
 sg13g2_decap_8 FILLER_6_159 ();
 sg13g2_decap_8 FILLER_6_166 ();
 sg13g2_fill_1 FILLER_6_173 ();
 sg13g2_fill_1 FILLER_6_183 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_228 ();
 sg13g2_fill_2 FILLER_6_235 ();
 sg13g2_fill_2 FILLER_6_249 ();
 sg13g2_fill_1 FILLER_6_251 ();
 sg13g2_decap_8 FILLER_6_257 ();
 sg13g2_decap_4 FILLER_6_264 ();
 sg13g2_fill_2 FILLER_6_268 ();
 sg13g2_fill_1 FILLER_6_284 ();
 sg13g2_decap_8 FILLER_6_299 ();
 sg13g2_decap_8 FILLER_6_306 ();
 sg13g2_decap_8 FILLER_6_313 ();
 sg13g2_decap_4 FILLER_6_320 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_4 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_431 ();
 sg13g2_decap_8 FILLER_6_436 ();
 sg13g2_decap_8 FILLER_6_443 ();
 sg13g2_fill_1 FILLER_6_450 ();
 sg13g2_decap_8 FILLER_6_464 ();
 sg13g2_decap_8 FILLER_6_471 ();
 sg13g2_fill_2 FILLER_6_478 ();
 sg13g2_decap_8 FILLER_6_489 ();
 sg13g2_fill_2 FILLER_6_496 ();
 sg13g2_fill_1 FILLER_6_498 ();
 sg13g2_decap_4 FILLER_6_529 ();
 sg13g2_fill_1 FILLER_6_533 ();
 sg13g2_fill_1 FILLER_6_539 ();
 sg13g2_decap_4 FILLER_6_561 ();
 sg13g2_fill_2 FILLER_6_565 ();
 sg13g2_decap_8 FILLER_6_571 ();
 sg13g2_decap_8 FILLER_6_578 ();
 sg13g2_decap_8 FILLER_6_585 ();
 sg13g2_decap_8 FILLER_6_592 ();
 sg13g2_fill_2 FILLER_6_599 ();
 sg13g2_fill_1 FILLER_6_601 ();
 sg13g2_decap_8 FILLER_6_614 ();
 sg13g2_decap_8 FILLER_6_621 ();
 sg13g2_fill_2 FILLER_6_628 ();
 sg13g2_fill_1 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_647 ();
 sg13g2_decap_4 FILLER_6_657 ();
 sg13g2_fill_2 FILLER_6_673 ();
 sg13g2_decap_8 FILLER_6_685 ();
 sg13g2_decap_4 FILLER_6_692 ();
 sg13g2_decap_4 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_712 ();
 sg13g2_decap_4 FILLER_6_719 ();
 sg13g2_decap_8 FILLER_6_727 ();
 sg13g2_decap_8 FILLER_6_734 ();
 sg13g2_decap_8 FILLER_6_741 ();
 sg13g2_decap_8 FILLER_6_748 ();
 sg13g2_fill_1 FILLER_6_755 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_4 FILLER_6_805 ();
 sg13g2_fill_1 FILLER_6_809 ();
 sg13g2_fill_2 FILLER_6_814 ();
 sg13g2_fill_1 FILLER_6_816 ();
 sg13g2_decap_8 FILLER_6_834 ();
 sg13g2_decap_8 FILLER_6_841 ();
 sg13g2_decap_8 FILLER_6_848 ();
 sg13g2_decap_8 FILLER_6_855 ();
 sg13g2_decap_8 FILLER_6_862 ();
 sg13g2_decap_8 FILLER_6_869 ();
 sg13g2_decap_8 FILLER_6_876 ();
 sg13g2_decap_8 FILLER_6_883 ();
 sg13g2_decap_8 FILLER_6_890 ();
 sg13g2_fill_2 FILLER_6_897 ();
 sg13g2_fill_1 FILLER_6_899 ();
 sg13g2_decap_8 FILLER_6_904 ();
 sg13g2_decap_8 FILLER_6_911 ();
 sg13g2_decap_8 FILLER_6_918 ();
 sg13g2_decap_8 FILLER_6_925 ();
 sg13g2_decap_4 FILLER_6_932 ();
 sg13g2_fill_1 FILLER_6_936 ();
 sg13g2_decap_8 FILLER_6_976 ();
 sg13g2_fill_1 FILLER_6_983 ();
 sg13g2_decap_8 FILLER_6_988 ();
 sg13g2_decap_8 FILLER_6_995 ();
 sg13g2_decap_8 FILLER_6_1002 ();
 sg13g2_decap_8 FILLER_6_1009 ();
 sg13g2_decap_8 FILLER_6_1016 ();
 sg13g2_decap_8 FILLER_6_1023 ();
 sg13g2_decap_8 FILLER_6_1030 ();
 sg13g2_decap_8 FILLER_6_1037 ();
 sg13g2_decap_8 FILLER_6_1044 ();
 sg13g2_fill_1 FILLER_6_1051 ();
 sg13g2_decap_8 FILLER_6_1056 ();
 sg13g2_decap_8 FILLER_6_1063 ();
 sg13g2_decap_8 FILLER_6_1070 ();
 sg13g2_decap_8 FILLER_6_1077 ();
 sg13g2_decap_8 FILLER_6_1084 ();
 sg13g2_decap_4 FILLER_6_1091 ();
 sg13g2_decap_4 FILLER_6_1100 ();
 sg13g2_fill_1 FILLER_6_1104 ();
 sg13g2_decap_8 FILLER_6_1115 ();
 sg13g2_decap_8 FILLER_6_1122 ();
 sg13g2_decap_8 FILLER_6_1129 ();
 sg13g2_fill_2 FILLER_6_1136 ();
 sg13g2_decap_8 FILLER_6_1155 ();
 sg13g2_decap_8 FILLER_6_1162 ();
 sg13g2_decap_8 FILLER_6_1199 ();
 sg13g2_decap_8 FILLER_6_1206 ();
 sg13g2_decap_8 FILLER_6_1213 ();
 sg13g2_decap_8 FILLER_6_1220 ();
 sg13g2_decap_8 FILLER_6_1227 ();
 sg13g2_decap_8 FILLER_6_1234 ();
 sg13g2_decap_8 FILLER_6_1241 ();
 sg13g2_decap_8 FILLER_6_1248 ();
 sg13g2_decap_8 FILLER_6_1255 ();
 sg13g2_decap_8 FILLER_6_1262 ();
 sg13g2_decap_8 FILLER_6_1269 ();
 sg13g2_decap_8 FILLER_6_1276 ();
 sg13g2_decap_8 FILLER_6_1283 ();
 sg13g2_decap_8 FILLER_6_1290 ();
 sg13g2_decap_8 FILLER_6_1297 ();
 sg13g2_decap_8 FILLER_6_1304 ();
 sg13g2_decap_8 FILLER_6_1311 ();
 sg13g2_decap_8 FILLER_6_1318 ();
 sg13g2_fill_1 FILLER_6_1325 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_fill_2 FILLER_7_72 ();
 sg13g2_fill_1 FILLER_7_107 ();
 sg13g2_decap_4 FILLER_7_113 ();
 sg13g2_fill_2 FILLER_7_117 ();
 sg13g2_decap_8 FILLER_7_122 ();
 sg13g2_fill_2 FILLER_7_129 ();
 sg13g2_fill_2 FILLER_7_137 ();
 sg13g2_decap_8 FILLER_7_162 ();
 sg13g2_fill_1 FILLER_7_169 ();
 sg13g2_decap_8 FILLER_7_185 ();
 sg13g2_decap_8 FILLER_7_192 ();
 sg13g2_decap_8 FILLER_7_199 ();
 sg13g2_decap_4 FILLER_7_206 ();
 sg13g2_fill_1 FILLER_7_210 ();
 sg13g2_fill_1 FILLER_7_237 ();
 sg13g2_fill_2 FILLER_7_243 ();
 sg13g2_fill_1 FILLER_7_245 ();
 sg13g2_decap_4 FILLER_7_262 ();
 sg13g2_fill_2 FILLER_7_270 ();
 sg13g2_decap_8 FILLER_7_277 ();
 sg13g2_fill_1 FILLER_7_284 ();
 sg13g2_decap_8 FILLER_7_289 ();
 sg13g2_decap_8 FILLER_7_296 ();
 sg13g2_decap_8 FILLER_7_303 ();
 sg13g2_decap_8 FILLER_7_310 ();
 sg13g2_decap_8 FILLER_7_317 ();
 sg13g2_decap_8 FILLER_7_324 ();
 sg13g2_decap_8 FILLER_7_331 ();
 sg13g2_decap_8 FILLER_7_338 ();
 sg13g2_decap_8 FILLER_7_345 ();
 sg13g2_decap_8 FILLER_7_352 ();
 sg13g2_decap_8 FILLER_7_359 ();
 sg13g2_decap_8 FILLER_7_366 ();
 sg13g2_decap_8 FILLER_7_373 ();
 sg13g2_decap_8 FILLER_7_380 ();
 sg13g2_decap_8 FILLER_7_387 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_decap_8 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_7_415 ();
 sg13g2_decap_8 FILLER_7_422 ();
 sg13g2_decap_8 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_7_436 ();
 sg13g2_decap_8 FILLER_7_443 ();
 sg13g2_decap_8 FILLER_7_450 ();
 sg13g2_decap_8 FILLER_7_457 ();
 sg13g2_decap_8 FILLER_7_464 ();
 sg13g2_fill_2 FILLER_7_471 ();
 sg13g2_fill_1 FILLER_7_473 ();
 sg13g2_decap_4 FILLER_7_504 ();
 sg13g2_fill_2 FILLER_7_508 ();
 sg13g2_decap_8 FILLER_7_514 ();
 sg13g2_fill_1 FILLER_7_521 ();
 sg13g2_fill_2 FILLER_7_557 ();
 sg13g2_fill_1 FILLER_7_559 ();
 sg13g2_decap_8 FILLER_7_586 ();
 sg13g2_decap_4 FILLER_7_593 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_fill_2 FILLER_7_630 ();
 sg13g2_decap_4 FILLER_7_689 ();
 sg13g2_decap_8 FILLER_7_727 ();
 sg13g2_decap_8 FILLER_7_739 ();
 sg13g2_decap_8 FILLER_7_746 ();
 sg13g2_decap_4 FILLER_7_753 ();
 sg13g2_decap_8 FILLER_7_792 ();
 sg13g2_decap_4 FILLER_7_799 ();
 sg13g2_decap_8 FILLER_7_834 ();
 sg13g2_decap_8 FILLER_7_841 ();
 sg13g2_decap_8 FILLER_7_848 ();
 sg13g2_decap_8 FILLER_7_855 ();
 sg13g2_decap_8 FILLER_7_862 ();
 sg13g2_decap_8 FILLER_7_869 ();
 sg13g2_decap_8 FILLER_7_876 ();
 sg13g2_decap_8 FILLER_7_883 ();
 sg13g2_decap_8 FILLER_7_890 ();
 sg13g2_decap_8 FILLER_7_897 ();
 sg13g2_decap_8 FILLER_7_904 ();
 sg13g2_decap_8 FILLER_7_911 ();
 sg13g2_decap_8 FILLER_7_918 ();
 sg13g2_decap_8 FILLER_7_925 ();
 sg13g2_decap_8 FILLER_7_932 ();
 sg13g2_fill_2 FILLER_7_939 ();
 sg13g2_fill_1 FILLER_7_941 ();
 sg13g2_decap_8 FILLER_7_948 ();
 sg13g2_decap_8 FILLER_7_955 ();
 sg13g2_decap_8 FILLER_7_962 ();
 sg13g2_decap_8 FILLER_7_969 ();
 sg13g2_decap_8 FILLER_7_976 ();
 sg13g2_decap_8 FILLER_7_983 ();
 sg13g2_decap_8 FILLER_7_990 ();
 sg13g2_fill_1 FILLER_7_997 ();
 sg13g2_decap_8 FILLER_7_1003 ();
 sg13g2_fill_2 FILLER_7_1010 ();
 sg13g2_fill_1 FILLER_7_1012 ();
 sg13g2_decap_8 FILLER_7_1042 ();
 sg13g2_decap_8 FILLER_7_1049 ();
 sg13g2_decap_4 FILLER_7_1056 ();
 sg13g2_fill_2 FILLER_7_1060 ();
 sg13g2_decap_4 FILLER_7_1066 ();
 sg13g2_decap_8 FILLER_7_1078 ();
 sg13g2_fill_1 FILLER_7_1089 ();
 sg13g2_decap_8 FILLER_7_1094 ();
 sg13g2_decap_4 FILLER_7_1101 ();
 sg13g2_fill_1 FILLER_7_1105 ();
 sg13g2_fill_1 FILLER_7_1132 ();
 sg13g2_decap_4 FILLER_7_1137 ();
 sg13g2_decap_8 FILLER_7_1149 ();
 sg13g2_decap_8 FILLER_7_1156 ();
 sg13g2_decap_8 FILLER_7_1201 ();
 sg13g2_decap_8 FILLER_7_1208 ();
 sg13g2_decap_8 FILLER_7_1215 ();
 sg13g2_decap_8 FILLER_7_1222 ();
 sg13g2_decap_8 FILLER_7_1229 ();
 sg13g2_decap_8 FILLER_7_1236 ();
 sg13g2_decap_8 FILLER_7_1243 ();
 sg13g2_decap_8 FILLER_7_1250 ();
 sg13g2_decap_8 FILLER_7_1257 ();
 sg13g2_decap_8 FILLER_7_1264 ();
 sg13g2_decap_8 FILLER_7_1271 ();
 sg13g2_decap_8 FILLER_7_1278 ();
 sg13g2_decap_8 FILLER_7_1285 ();
 sg13g2_decap_8 FILLER_7_1292 ();
 sg13g2_decap_8 FILLER_7_1299 ();
 sg13g2_decap_8 FILLER_7_1306 ();
 sg13g2_decap_8 FILLER_7_1313 ();
 sg13g2_decap_4 FILLER_7_1320 ();
 sg13g2_fill_2 FILLER_7_1324 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_4 FILLER_8_49 ();
 sg13g2_fill_2 FILLER_8_53 ();
 sg13g2_decap_8 FILLER_8_71 ();
 sg13g2_decap_4 FILLER_8_78 ();
 sg13g2_fill_2 FILLER_8_82 ();
 sg13g2_fill_1 FILLER_8_97 ();
 sg13g2_fill_2 FILLER_8_111 ();
 sg13g2_decap_8 FILLER_8_117 ();
 sg13g2_fill_1 FILLER_8_124 ();
 sg13g2_fill_2 FILLER_8_137 ();
 sg13g2_fill_1 FILLER_8_139 ();
 sg13g2_fill_2 FILLER_8_145 ();
 sg13g2_fill_2 FILLER_8_151 ();
 sg13g2_fill_1 FILLER_8_153 ();
 sg13g2_decap_4 FILLER_8_176 ();
 sg13g2_fill_1 FILLER_8_180 ();
 sg13g2_decap_8 FILLER_8_185 ();
 sg13g2_decap_8 FILLER_8_192 ();
 sg13g2_fill_2 FILLER_8_199 ();
 sg13g2_fill_1 FILLER_8_201 ();
 sg13g2_decap_4 FILLER_8_206 ();
 sg13g2_fill_2 FILLER_8_210 ();
 sg13g2_fill_2 FILLER_8_234 ();
 sg13g2_fill_1 FILLER_8_240 ();
 sg13g2_decap_8 FILLER_8_246 ();
 sg13g2_decap_8 FILLER_8_253 ();
 sg13g2_decap_4 FILLER_8_260 ();
 sg13g2_decap_8 FILLER_8_278 ();
 sg13g2_decap_4 FILLER_8_285 ();
 sg13g2_fill_2 FILLER_8_289 ();
 sg13g2_decap_4 FILLER_8_299 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_fill_2 FILLER_8_314 ();
 sg13g2_fill_1 FILLER_8_316 ();
 sg13g2_fill_1 FILLER_8_320 ();
 sg13g2_decap_8 FILLER_8_331 ();
 sg13g2_decap_8 FILLER_8_338 ();
 sg13g2_decap_8 FILLER_8_345 ();
 sg13g2_decap_8 FILLER_8_352 ();
 sg13g2_decap_8 FILLER_8_359 ();
 sg13g2_decap_4 FILLER_8_366 ();
 sg13g2_fill_2 FILLER_8_370 ();
 sg13g2_fill_2 FILLER_8_378 ();
 sg13g2_fill_1 FILLER_8_380 ();
 sg13g2_fill_2 FILLER_8_390 ();
 sg13g2_fill_1 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_fill_1 FILLER_8_404 ();
 sg13g2_fill_2 FILLER_8_410 ();
 sg13g2_decap_8 FILLER_8_433 ();
 sg13g2_decap_8 FILLER_8_440 ();
 sg13g2_decap_8 FILLER_8_447 ();
 sg13g2_decap_8 FILLER_8_454 ();
 sg13g2_decap_8 FILLER_8_461 ();
 sg13g2_decap_8 FILLER_8_468 ();
 sg13g2_decap_8 FILLER_8_475 ();
 sg13g2_decap_8 FILLER_8_482 ();
 sg13g2_decap_8 FILLER_8_489 ();
 sg13g2_decap_8 FILLER_8_496 ();
 sg13g2_decap_8 FILLER_8_503 ();
 sg13g2_fill_2 FILLER_8_510 ();
 sg13g2_decap_8 FILLER_8_517 ();
 sg13g2_decap_8 FILLER_8_524 ();
 sg13g2_fill_2 FILLER_8_531 ();
 sg13g2_decap_8 FILLER_8_537 ();
 sg13g2_decap_8 FILLER_8_544 ();
 sg13g2_fill_2 FILLER_8_551 ();
 sg13g2_decap_8 FILLER_8_557 ();
 sg13g2_decap_8 FILLER_8_564 ();
 sg13g2_decap_8 FILLER_8_571 ();
 sg13g2_decap_8 FILLER_8_578 ();
 sg13g2_decap_8 FILLER_8_585 ();
 sg13g2_decap_8 FILLER_8_592 ();
 sg13g2_decap_4 FILLER_8_599 ();
 sg13g2_fill_2 FILLER_8_603 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_fill_1 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_642 ();
 sg13g2_decap_8 FILLER_8_649 ();
 sg13g2_decap_8 FILLER_8_656 ();
 sg13g2_fill_1 FILLER_8_663 ();
 sg13g2_decap_8 FILLER_8_668 ();
 sg13g2_decap_8 FILLER_8_675 ();
 sg13g2_decap_8 FILLER_8_682 ();
 sg13g2_decap_4 FILLER_8_689 ();
 sg13g2_fill_2 FILLER_8_693 ();
 sg13g2_fill_2 FILLER_8_703 ();
 sg13g2_fill_1 FILLER_8_705 ();
 sg13g2_decap_4 FILLER_8_709 ();
 sg13g2_fill_2 FILLER_8_713 ();
 sg13g2_fill_1 FILLER_8_724 ();
 sg13g2_decap_8 FILLER_8_730 ();
 sg13g2_decap_4 FILLER_8_737 ();
 sg13g2_decap_8 FILLER_8_745 ();
 sg13g2_decap_8 FILLER_8_752 ();
 sg13g2_fill_2 FILLER_8_759 ();
 sg13g2_decap_8 FILLER_8_765 ();
 sg13g2_fill_1 FILLER_8_772 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_4 FILLER_8_805 ();
 sg13g2_fill_2 FILLER_8_809 ();
 sg13g2_decap_8 FILLER_8_815 ();
 sg13g2_decap_8 FILLER_8_822 ();
 sg13g2_decap_8 FILLER_8_829 ();
 sg13g2_decap_8 FILLER_8_836 ();
 sg13g2_decap_4 FILLER_8_843 ();
 sg13g2_decap_8 FILLER_8_873 ();
 sg13g2_fill_2 FILLER_8_880 ();
 sg13g2_fill_1 FILLER_8_882 ();
 sg13g2_decap_8 FILLER_8_892 ();
 sg13g2_decap_4 FILLER_8_899 ();
 sg13g2_fill_1 FILLER_8_903 ();
 sg13g2_decap_8 FILLER_8_916 ();
 sg13g2_decap_8 FILLER_8_923 ();
 sg13g2_fill_2 FILLER_8_943 ();
 sg13g2_decap_4 FILLER_8_957 ();
 sg13g2_fill_2 FILLER_8_961 ();
 sg13g2_decap_8 FILLER_8_974 ();
 sg13g2_decap_8 FILLER_8_981 ();
 sg13g2_decap_4 FILLER_8_988 ();
 sg13g2_fill_1 FILLER_8_992 ();
 sg13g2_decap_8 FILLER_8_1002 ();
 sg13g2_fill_2 FILLER_8_1009 ();
 sg13g2_fill_1 FILLER_8_1011 ();
 sg13g2_decap_8 FILLER_8_1020 ();
 sg13g2_decap_8 FILLER_8_1027 ();
 sg13g2_decap_8 FILLER_8_1042 ();
 sg13g2_decap_8 FILLER_8_1049 ();
 sg13g2_decap_4 FILLER_8_1056 ();
 sg13g2_fill_1 FILLER_8_1060 ();
 sg13g2_fill_2 FILLER_8_1087 ();
 sg13g2_decap_8 FILLER_8_1097 ();
 sg13g2_decap_8 FILLER_8_1104 ();
 sg13g2_fill_1 FILLER_8_1111 ();
 sg13g2_decap_8 FILLER_8_1116 ();
 sg13g2_decap_8 FILLER_8_1123 ();
 sg13g2_fill_2 FILLER_8_1130 ();
 sg13g2_decap_8 FILLER_8_1158 ();
 sg13g2_decap_8 FILLER_8_1165 ();
 sg13g2_fill_1 FILLER_8_1172 ();
 sg13g2_decap_8 FILLER_8_1177 ();
 sg13g2_decap_8 FILLER_8_1184 ();
 sg13g2_decap_8 FILLER_8_1191 ();
 sg13g2_decap_8 FILLER_8_1198 ();
 sg13g2_decap_8 FILLER_8_1205 ();
 sg13g2_decap_8 FILLER_8_1212 ();
 sg13g2_decap_8 FILLER_8_1219 ();
 sg13g2_decap_8 FILLER_8_1226 ();
 sg13g2_decap_8 FILLER_8_1233 ();
 sg13g2_decap_8 FILLER_8_1240 ();
 sg13g2_decap_8 FILLER_8_1247 ();
 sg13g2_decap_8 FILLER_8_1254 ();
 sg13g2_decap_8 FILLER_8_1261 ();
 sg13g2_decap_8 FILLER_8_1268 ();
 sg13g2_decap_8 FILLER_8_1275 ();
 sg13g2_decap_8 FILLER_8_1282 ();
 sg13g2_decap_8 FILLER_8_1289 ();
 sg13g2_decap_8 FILLER_8_1296 ();
 sg13g2_decap_8 FILLER_8_1303 ();
 sg13g2_decap_8 FILLER_8_1310 ();
 sg13g2_decap_8 FILLER_8_1317 ();
 sg13g2_fill_2 FILLER_8_1324 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_fill_1 FILLER_9_42 ();
 sg13g2_decap_4 FILLER_9_56 ();
 sg13g2_fill_2 FILLER_9_60 ();
 sg13g2_decap_4 FILLER_9_79 ();
 sg13g2_fill_1 FILLER_9_83 ();
 sg13g2_decap_8 FILLER_9_113 ();
 sg13g2_decap_8 FILLER_9_120 ();
 sg13g2_decap_8 FILLER_9_127 ();
 sg13g2_decap_8 FILLER_9_138 ();
 sg13g2_decap_8 FILLER_9_145 ();
 sg13g2_decap_8 FILLER_9_152 ();
 sg13g2_fill_2 FILLER_9_159 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_fill_2 FILLER_9_167 ();
 sg13g2_decap_8 FILLER_9_173 ();
 sg13g2_decap_8 FILLER_9_180 ();
 sg13g2_decap_8 FILLER_9_187 ();
 sg13g2_decap_8 FILLER_9_194 ();
 sg13g2_decap_8 FILLER_9_201 ();
 sg13g2_decap_8 FILLER_9_208 ();
 sg13g2_decap_8 FILLER_9_215 ();
 sg13g2_decap_8 FILLER_9_222 ();
 sg13g2_decap_8 FILLER_9_229 ();
 sg13g2_decap_8 FILLER_9_236 ();
 sg13g2_decap_8 FILLER_9_243 ();
 sg13g2_decap_8 FILLER_9_264 ();
 sg13g2_fill_1 FILLER_9_271 ();
 sg13g2_decap_4 FILLER_9_282 ();
 sg13g2_fill_2 FILLER_9_300 ();
 sg13g2_fill_1 FILLER_9_307 ();
 sg13g2_fill_1 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_327 ();
 sg13g2_decap_8 FILLER_9_334 ();
 sg13g2_fill_1 FILLER_9_341 ();
 sg13g2_fill_2 FILLER_9_419 ();
 sg13g2_decap_8 FILLER_9_447 ();
 sg13g2_decap_4 FILLER_9_454 ();
 sg13g2_fill_1 FILLER_9_458 ();
 sg13g2_decap_8 FILLER_9_468 ();
 sg13g2_decap_8 FILLER_9_475 ();
 sg13g2_decap_8 FILLER_9_482 ();
 sg13g2_decap_8 FILLER_9_489 ();
 sg13g2_decap_8 FILLER_9_496 ();
 sg13g2_decap_8 FILLER_9_503 ();
 sg13g2_decap_8 FILLER_9_510 ();
 sg13g2_decap_8 FILLER_9_517 ();
 sg13g2_decap_8 FILLER_9_524 ();
 sg13g2_decap_8 FILLER_9_531 ();
 sg13g2_decap_8 FILLER_9_538 ();
 sg13g2_decap_8 FILLER_9_545 ();
 sg13g2_decap_8 FILLER_9_552 ();
 sg13g2_decap_8 FILLER_9_559 ();
 sg13g2_fill_2 FILLER_9_566 ();
 sg13g2_decap_8 FILLER_9_572 ();
 sg13g2_decap_8 FILLER_9_579 ();
 sg13g2_decap_8 FILLER_9_586 ();
 sg13g2_decap_8 FILLER_9_593 ();
 sg13g2_decap_8 FILLER_9_600 ();
 sg13g2_decap_8 FILLER_9_607 ();
 sg13g2_fill_2 FILLER_9_614 ();
 sg13g2_fill_1 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_621 ();
 sg13g2_decap_8 FILLER_9_628 ();
 sg13g2_decap_8 FILLER_9_635 ();
 sg13g2_decap_4 FILLER_9_642 ();
 sg13g2_fill_1 FILLER_9_646 ();
 sg13g2_decap_8 FILLER_9_655 ();
 sg13g2_decap_8 FILLER_9_662 ();
 sg13g2_decap_8 FILLER_9_669 ();
 sg13g2_decap_8 FILLER_9_676 ();
 sg13g2_fill_2 FILLER_9_683 ();
 sg13g2_fill_1 FILLER_9_685 ();
 sg13g2_decap_8 FILLER_9_712 ();
 sg13g2_decap_4 FILLER_9_719 ();
 sg13g2_fill_2 FILLER_9_723 ();
 sg13g2_decap_8 FILLER_9_729 ();
 sg13g2_fill_1 FILLER_9_769 ();
 sg13g2_fill_2 FILLER_9_796 ();
 sg13g2_fill_1 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_813 ();
 sg13g2_decap_8 FILLER_9_820 ();
 sg13g2_decap_8 FILLER_9_827 ();
 sg13g2_decap_4 FILLER_9_834 ();
 sg13g2_fill_1 FILLER_9_853 ();
 sg13g2_fill_2 FILLER_9_858 ();
 sg13g2_fill_1 FILLER_9_860 ();
 sg13g2_decap_8 FILLER_9_869 ();
 sg13g2_decap_8 FILLER_9_876 ();
 sg13g2_fill_2 FILLER_9_883 ();
 sg13g2_decap_8 FILLER_9_894 ();
 sg13g2_decap_4 FILLER_9_901 ();
 sg13g2_decap_8 FILLER_9_943 ();
 sg13g2_fill_2 FILLER_9_950 ();
 sg13g2_fill_2 FILLER_9_956 ();
 sg13g2_fill_2 FILLER_9_984 ();
 sg13g2_fill_1 FILLER_9_1022 ();
 sg13g2_decap_8 FILLER_9_1053 ();
 sg13g2_decap_8 FILLER_9_1060 ();
 sg13g2_fill_2 FILLER_9_1067 ();
 sg13g2_fill_1 FILLER_9_1069 ();
 sg13g2_decap_4 FILLER_9_1074 ();
 sg13g2_fill_1 FILLER_9_1082 ();
 sg13g2_decap_8 FILLER_9_1109 ();
 sg13g2_decap_8 FILLER_9_1116 ();
 sg13g2_decap_8 FILLER_9_1123 ();
 sg13g2_decap_8 FILLER_9_1130 ();
 sg13g2_decap_8 FILLER_9_1141 ();
 sg13g2_decap_8 FILLER_9_1148 ();
 sg13g2_decap_8 FILLER_9_1155 ();
 sg13g2_decap_8 FILLER_9_1162 ();
 sg13g2_decap_8 FILLER_9_1169 ();
 sg13g2_decap_8 FILLER_9_1176 ();
 sg13g2_decap_8 FILLER_9_1183 ();
 sg13g2_decap_8 FILLER_9_1190 ();
 sg13g2_decap_8 FILLER_9_1197 ();
 sg13g2_decap_8 FILLER_9_1204 ();
 sg13g2_decap_8 FILLER_9_1211 ();
 sg13g2_decap_8 FILLER_9_1218 ();
 sg13g2_decap_8 FILLER_9_1225 ();
 sg13g2_decap_8 FILLER_9_1232 ();
 sg13g2_decap_8 FILLER_9_1239 ();
 sg13g2_decap_8 FILLER_9_1246 ();
 sg13g2_decap_8 FILLER_9_1253 ();
 sg13g2_decap_8 FILLER_9_1260 ();
 sg13g2_decap_8 FILLER_9_1267 ();
 sg13g2_decap_8 FILLER_9_1274 ();
 sg13g2_decap_8 FILLER_9_1281 ();
 sg13g2_decap_8 FILLER_9_1288 ();
 sg13g2_decap_8 FILLER_9_1295 ();
 sg13g2_decap_8 FILLER_9_1302 ();
 sg13g2_decap_8 FILLER_9_1309 ();
 sg13g2_decap_8 FILLER_9_1316 ();
 sg13g2_fill_2 FILLER_9_1323 ();
 sg13g2_fill_1 FILLER_9_1325 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_4 FILLER_10_21 ();
 sg13g2_fill_1 FILLER_10_25 ();
 sg13g2_decap_8 FILLER_10_31 ();
 sg13g2_decap_8 FILLER_10_38 ();
 sg13g2_decap_8 FILLER_10_45 ();
 sg13g2_fill_1 FILLER_10_52 ();
 sg13g2_fill_2 FILLER_10_58 ();
 sg13g2_fill_2 FILLER_10_71 ();
 sg13g2_fill_1 FILLER_10_73 ();
 sg13g2_decap_4 FILLER_10_79 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_107 ();
 sg13g2_decap_8 FILLER_10_118 ();
 sg13g2_decap_4 FILLER_10_125 ();
 sg13g2_decap_8 FILLER_10_138 ();
 sg13g2_fill_2 FILLER_10_145 ();
 sg13g2_fill_1 FILLER_10_147 ();
 sg13g2_decap_4 FILLER_10_153 ();
 sg13g2_fill_2 FILLER_10_157 ();
 sg13g2_decap_4 FILLER_10_163 ();
 sg13g2_fill_2 FILLER_10_167 ();
 sg13g2_decap_8 FILLER_10_173 ();
 sg13g2_decap_8 FILLER_10_180 ();
 sg13g2_decap_8 FILLER_10_187 ();
 sg13g2_decap_8 FILLER_10_194 ();
 sg13g2_decap_8 FILLER_10_201 ();
 sg13g2_decap_4 FILLER_10_208 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_4 FILLER_10_235 ();
 sg13g2_fill_1 FILLER_10_239 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_fill_1 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_279 ();
 sg13g2_fill_1 FILLER_10_286 ();
 sg13g2_decap_8 FILLER_10_292 ();
 sg13g2_decap_8 FILLER_10_299 ();
 sg13g2_fill_2 FILLER_10_306 ();
 sg13g2_decap_8 FILLER_10_327 ();
 sg13g2_decap_8 FILLER_10_334 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_decap_8 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_408 ();
 sg13g2_decap_4 FILLER_10_415 ();
 sg13g2_fill_2 FILLER_10_423 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_fill_1 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_484 ();
 sg13g2_decap_8 FILLER_10_491 ();
 sg13g2_fill_2 FILLER_10_498 ();
 sg13g2_fill_1 FILLER_10_500 ();
 sg13g2_decap_8 FILLER_10_505 ();
 sg13g2_fill_1 FILLER_10_512 ();
 sg13g2_decap_4 FILLER_10_522 ();
 sg13g2_decap_8 FILLER_10_534 ();
 sg13g2_fill_2 FILLER_10_541 ();
 sg13g2_fill_1 FILLER_10_543 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_fill_1 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_587 ();
 sg13g2_decap_8 FILLER_10_594 ();
 sg13g2_decap_8 FILLER_10_601 ();
 sg13g2_fill_2 FILLER_10_608 ();
 sg13g2_fill_1 FILLER_10_610 ();
 sg13g2_decap_8 FILLER_10_615 ();
 sg13g2_decap_8 FILLER_10_622 ();
 sg13g2_decap_8 FILLER_10_629 ();
 sg13g2_decap_8 FILLER_10_636 ();
 sg13g2_decap_8 FILLER_10_643 ();
 sg13g2_decap_8 FILLER_10_650 ();
 sg13g2_decap_8 FILLER_10_657 ();
 sg13g2_decap_4 FILLER_10_664 ();
 sg13g2_fill_2 FILLER_10_668 ();
 sg13g2_decap_8 FILLER_10_678 ();
 sg13g2_decap_8 FILLER_10_685 ();
 sg13g2_fill_2 FILLER_10_692 ();
 sg13g2_fill_1 FILLER_10_694 ();
 sg13g2_decap_8 FILLER_10_699 ();
 sg13g2_decap_8 FILLER_10_706 ();
 sg13g2_decap_8 FILLER_10_713 ();
 sg13g2_decap_4 FILLER_10_720 ();
 sg13g2_fill_1 FILLER_10_724 ();
 sg13g2_decap_8 FILLER_10_755 ();
 sg13g2_fill_1 FILLER_10_766 ();
 sg13g2_decap_4 FILLER_10_771 ();
 sg13g2_fill_2 FILLER_10_775 ();
 sg13g2_decap_8 FILLER_10_781 ();
 sg13g2_decap_8 FILLER_10_788 ();
 sg13g2_decap_8 FILLER_10_795 ();
 sg13g2_decap_8 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_809 ();
 sg13g2_decap_4 FILLER_10_816 ();
 sg13g2_fill_1 FILLER_10_820 ();
 sg13g2_decap_8 FILLER_10_846 ();
 sg13g2_decap_8 FILLER_10_853 ();
 sg13g2_decap_4 FILLER_10_860 ();
 sg13g2_fill_1 FILLER_10_864 ();
 sg13g2_fill_1 FILLER_10_869 ();
 sg13g2_decap_8 FILLER_10_879 ();
 sg13g2_fill_1 FILLER_10_886 ();
 sg13g2_fill_2 FILLER_10_899 ();
 sg13g2_decap_8 FILLER_10_905 ();
 sg13g2_fill_2 FILLER_10_912 ();
 sg13g2_decap_8 FILLER_10_918 ();
 sg13g2_fill_2 FILLER_10_925 ();
 sg13g2_fill_1 FILLER_10_927 ();
 sg13g2_decap_8 FILLER_10_954 ();
 sg13g2_fill_2 FILLER_10_961 ();
 sg13g2_fill_1 FILLER_10_963 ();
 sg13g2_decap_8 FILLER_10_968 ();
 sg13g2_decap_8 FILLER_10_975 ();
 sg13g2_decap_4 FILLER_10_982 ();
 sg13g2_fill_1 FILLER_10_986 ();
 sg13g2_fill_2 FILLER_10_1000 ();
 sg13g2_decap_8 FILLER_10_1012 ();
 sg13g2_decap_8 FILLER_10_1019 ();
 sg13g2_decap_8 FILLER_10_1026 ();
 sg13g2_fill_2 FILLER_10_1033 ();
 sg13g2_fill_1 FILLER_10_1035 ();
 sg13g2_decap_8 FILLER_10_1040 ();
 sg13g2_decap_8 FILLER_10_1047 ();
 sg13g2_decap_8 FILLER_10_1054 ();
 sg13g2_decap_8 FILLER_10_1061 ();
 sg13g2_decap_8 FILLER_10_1068 ();
 sg13g2_decap_8 FILLER_10_1075 ();
 sg13g2_decap_8 FILLER_10_1082 ();
 sg13g2_decap_8 FILLER_10_1093 ();
 sg13g2_decap_8 FILLER_10_1100 ();
 sg13g2_decap_8 FILLER_10_1107 ();
 sg13g2_decap_8 FILLER_10_1114 ();
 sg13g2_decap_8 FILLER_10_1121 ();
 sg13g2_decap_8 FILLER_10_1128 ();
 sg13g2_decap_8 FILLER_10_1135 ();
 sg13g2_decap_8 FILLER_10_1142 ();
 sg13g2_decap_8 FILLER_10_1149 ();
 sg13g2_decap_8 FILLER_10_1156 ();
 sg13g2_decap_8 FILLER_10_1163 ();
 sg13g2_decap_8 FILLER_10_1170 ();
 sg13g2_decap_8 FILLER_10_1177 ();
 sg13g2_decap_8 FILLER_10_1184 ();
 sg13g2_decap_8 FILLER_10_1191 ();
 sg13g2_decap_8 FILLER_10_1198 ();
 sg13g2_decap_8 FILLER_10_1205 ();
 sg13g2_decap_8 FILLER_10_1212 ();
 sg13g2_decap_8 FILLER_10_1219 ();
 sg13g2_decap_8 FILLER_10_1226 ();
 sg13g2_decap_8 FILLER_10_1233 ();
 sg13g2_decap_8 FILLER_10_1240 ();
 sg13g2_decap_8 FILLER_10_1247 ();
 sg13g2_decap_8 FILLER_10_1254 ();
 sg13g2_decap_8 FILLER_10_1261 ();
 sg13g2_decap_8 FILLER_10_1268 ();
 sg13g2_decap_8 FILLER_10_1275 ();
 sg13g2_decap_8 FILLER_10_1282 ();
 sg13g2_decap_8 FILLER_10_1289 ();
 sg13g2_decap_8 FILLER_10_1296 ();
 sg13g2_decap_8 FILLER_10_1303 ();
 sg13g2_decap_8 FILLER_10_1310 ();
 sg13g2_decap_8 FILLER_10_1317 ();
 sg13g2_fill_2 FILLER_10_1324 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_14 ();
 sg13g2_decap_4 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_43 ();
 sg13g2_decap_8 FILLER_11_50 ();
 sg13g2_decap_8 FILLER_11_57 ();
 sg13g2_decap_8 FILLER_11_64 ();
 sg13g2_decap_8 FILLER_11_71 ();
 sg13g2_decap_4 FILLER_11_78 ();
 sg13g2_fill_2 FILLER_11_82 ();
 sg13g2_decap_4 FILLER_11_90 ();
 sg13g2_fill_1 FILLER_11_94 ();
 sg13g2_decap_8 FILLER_11_100 ();
 sg13g2_decap_4 FILLER_11_107 ();
 sg13g2_fill_1 FILLER_11_111 ();
 sg13g2_decap_8 FILLER_11_116 ();
 sg13g2_decap_8 FILLER_11_123 ();
 sg13g2_decap_4 FILLER_11_130 ();
 sg13g2_fill_2 FILLER_11_134 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_fill_2 FILLER_11_161 ();
 sg13g2_fill_1 FILLER_11_163 ();
 sg13g2_decap_8 FILLER_11_177 ();
 sg13g2_decap_8 FILLER_11_184 ();
 sg13g2_decap_8 FILLER_11_197 ();
 sg13g2_decap_8 FILLER_11_204 ();
 sg13g2_decap_8 FILLER_11_211 ();
 sg13g2_decap_8 FILLER_11_218 ();
 sg13g2_decap_8 FILLER_11_225 ();
 sg13g2_decap_8 FILLER_11_232 ();
 sg13g2_decap_8 FILLER_11_239 ();
 sg13g2_decap_8 FILLER_11_246 ();
 sg13g2_decap_8 FILLER_11_253 ();
 sg13g2_decap_8 FILLER_11_260 ();
 sg13g2_decap_8 FILLER_11_267 ();
 sg13g2_decap_8 FILLER_11_274 ();
 sg13g2_decap_8 FILLER_11_281 ();
 sg13g2_decap_8 FILLER_11_288 ();
 sg13g2_decap_8 FILLER_11_295 ();
 sg13g2_decap_4 FILLER_11_302 ();
 sg13g2_fill_1 FILLER_11_306 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_fill_2 FILLER_11_375 ();
 sg13g2_fill_2 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_decap_8 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_11_415 ();
 sg13g2_decap_8 FILLER_11_422 ();
 sg13g2_decap_8 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_11_436 ();
 sg13g2_decap_8 FILLER_11_443 ();
 sg13g2_fill_2 FILLER_11_450 ();
 sg13g2_decap_8 FILLER_11_456 ();
 sg13g2_decap_4 FILLER_11_463 ();
 sg13g2_decap_4 FILLER_11_472 ();
 sg13g2_fill_2 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_482 ();
 sg13g2_decap_4 FILLER_11_559 ();
 sg13g2_fill_1 FILLER_11_563 ();
 sg13g2_decap_8 FILLER_11_585 ();
 sg13g2_decap_8 FILLER_11_592 ();
 sg13g2_decap_4 FILLER_11_599 ();
 sg13g2_fill_1 FILLER_11_603 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_fill_2 FILLER_11_637 ();
 sg13g2_fill_1 FILLER_11_639 ();
 sg13g2_decap_8 FILLER_11_666 ();
 sg13g2_decap_8 FILLER_11_677 ();
 sg13g2_decap_8 FILLER_11_684 ();
 sg13g2_decap_8 FILLER_11_691 ();
 sg13g2_decap_8 FILLER_11_698 ();
 sg13g2_decap_8 FILLER_11_705 ();
 sg13g2_decap_8 FILLER_11_712 ();
 sg13g2_decap_8 FILLER_11_719 ();
 sg13g2_decap_4 FILLER_11_726 ();
 sg13g2_fill_1 FILLER_11_730 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_782 ();
 sg13g2_decap_8 FILLER_11_789 ();
 sg13g2_fill_1 FILLER_11_796 ();
 sg13g2_fill_2 FILLER_11_830 ();
 sg13g2_fill_1 FILLER_11_832 ();
 sg13g2_fill_2 FILLER_11_856 ();
 sg13g2_fill_1 FILLER_11_858 ();
 sg13g2_fill_1 FILLER_11_867 ();
 sg13g2_decap_8 FILLER_11_894 ();
 sg13g2_decap_8 FILLER_11_901 ();
 sg13g2_decap_8 FILLER_11_908 ();
 sg13g2_decap_8 FILLER_11_915 ();
 sg13g2_decap_8 FILLER_11_922 ();
 sg13g2_decap_4 FILLER_11_929 ();
 sg13g2_decap_8 FILLER_11_937 ();
 sg13g2_decap_8 FILLER_11_944 ();
 sg13g2_decap_4 FILLER_11_951 ();
 sg13g2_fill_2 FILLER_11_955 ();
 sg13g2_decap_8 FILLER_11_971 ();
 sg13g2_decap_8 FILLER_11_978 ();
 sg13g2_decap_8 FILLER_11_985 ();
 sg13g2_decap_8 FILLER_11_992 ();
 sg13g2_decap_8 FILLER_11_999 ();
 sg13g2_decap_8 FILLER_11_1006 ();
 sg13g2_decap_8 FILLER_11_1013 ();
 sg13g2_decap_8 FILLER_11_1020 ();
 sg13g2_decap_8 FILLER_11_1027 ();
 sg13g2_decap_8 FILLER_11_1034 ();
 sg13g2_decap_8 FILLER_11_1041 ();
 sg13g2_decap_8 FILLER_11_1048 ();
 sg13g2_decap_8 FILLER_11_1055 ();
 sg13g2_decap_8 FILLER_11_1062 ();
 sg13g2_decap_8 FILLER_11_1069 ();
 sg13g2_decap_8 FILLER_11_1076 ();
 sg13g2_decap_8 FILLER_11_1083 ();
 sg13g2_decap_8 FILLER_11_1090 ();
 sg13g2_decap_8 FILLER_11_1097 ();
 sg13g2_decap_8 FILLER_11_1104 ();
 sg13g2_decap_8 FILLER_11_1111 ();
 sg13g2_decap_8 FILLER_11_1118 ();
 sg13g2_decap_8 FILLER_11_1125 ();
 sg13g2_decap_8 FILLER_11_1132 ();
 sg13g2_decap_8 FILLER_11_1139 ();
 sg13g2_decap_8 FILLER_11_1146 ();
 sg13g2_decap_4 FILLER_11_1153 ();
 sg13g2_fill_2 FILLER_11_1157 ();
 sg13g2_decap_8 FILLER_11_1163 ();
 sg13g2_decap_8 FILLER_11_1170 ();
 sg13g2_decap_8 FILLER_11_1177 ();
 sg13g2_decap_8 FILLER_11_1184 ();
 sg13g2_decap_8 FILLER_11_1191 ();
 sg13g2_decap_8 FILLER_11_1198 ();
 sg13g2_decap_8 FILLER_11_1205 ();
 sg13g2_decap_8 FILLER_11_1212 ();
 sg13g2_decap_8 FILLER_11_1219 ();
 sg13g2_decap_8 FILLER_11_1226 ();
 sg13g2_decap_8 FILLER_11_1233 ();
 sg13g2_decap_8 FILLER_11_1240 ();
 sg13g2_decap_8 FILLER_11_1247 ();
 sg13g2_decap_8 FILLER_11_1254 ();
 sg13g2_decap_8 FILLER_11_1261 ();
 sg13g2_decap_8 FILLER_11_1268 ();
 sg13g2_decap_8 FILLER_11_1275 ();
 sg13g2_decap_8 FILLER_11_1282 ();
 sg13g2_decap_8 FILLER_11_1289 ();
 sg13g2_decap_8 FILLER_11_1296 ();
 sg13g2_decap_8 FILLER_11_1303 ();
 sg13g2_decap_8 FILLER_11_1310 ();
 sg13g2_decap_8 FILLER_11_1317 ();
 sg13g2_fill_2 FILLER_11_1324 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_14 ();
 sg13g2_decap_4 FILLER_12_31 ();
 sg13g2_fill_1 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_48 ();
 sg13g2_decap_8 FILLER_12_55 ();
 sg13g2_decap_8 FILLER_12_62 ();
 sg13g2_decap_4 FILLER_12_81 ();
 sg13g2_fill_2 FILLER_12_97 ();
 sg13g2_fill_1 FILLER_12_99 ();
 sg13g2_fill_2 FILLER_12_121 ();
 sg13g2_fill_1 FILLER_12_123 ();
 sg13g2_decap_4 FILLER_12_128 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_4 FILLER_12_158 ();
 sg13g2_fill_1 FILLER_12_162 ();
 sg13g2_fill_1 FILLER_12_185 ();
 sg13g2_fill_1 FILLER_12_190 ();
 sg13g2_fill_1 FILLER_12_195 ();
 sg13g2_decap_4 FILLER_12_205 ();
 sg13g2_fill_1 FILLER_12_213 ();
 sg13g2_fill_2 FILLER_12_222 ();
 sg13g2_fill_2 FILLER_12_236 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_4 FILLER_12_263 ();
 sg13g2_fill_1 FILLER_12_267 ();
 sg13g2_decap_8 FILLER_12_271 ();
 sg13g2_decap_8 FILLER_12_278 ();
 sg13g2_decap_8 FILLER_12_285 ();
 sg13g2_fill_2 FILLER_12_292 ();
 sg13g2_fill_1 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_decap_8 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_338 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_decap_8 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_12_415 ();
 sg13g2_decap_8 FILLER_12_431 ();
 sg13g2_decap_8 FILLER_12_438 ();
 sg13g2_decap_4 FILLER_12_445 ();
 sg13g2_fill_1 FILLER_12_449 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_fill_1 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_509 ();
 sg13g2_decap_8 FILLER_12_516 ();
 sg13g2_decap_8 FILLER_12_523 ();
 sg13g2_decap_8 FILLER_12_534 ();
 sg13g2_decap_4 FILLER_12_541 ();
 sg13g2_fill_1 FILLER_12_545 ();
 sg13g2_decap_4 FILLER_12_551 ();
 sg13g2_fill_1 FILLER_12_555 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_4 FILLER_12_581 ();
 sg13g2_fill_2 FILLER_12_585 ();
 sg13g2_fill_2 FILLER_12_594 ();
 sg13g2_decap_4 FILLER_12_603 ();
 sg13g2_decap_4 FILLER_12_614 ();
 sg13g2_decap_4 FILLER_12_644 ();
 sg13g2_fill_2 FILLER_12_652 ();
 sg13g2_decap_4 FILLER_12_661 ();
 sg13g2_fill_1 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_692 ();
 sg13g2_decap_8 FILLER_12_699 ();
 sg13g2_decap_8 FILLER_12_706 ();
 sg13g2_decap_8 FILLER_12_713 ();
 sg13g2_decap_8 FILLER_12_720 ();
 sg13g2_decap_8 FILLER_12_727 ();
 sg13g2_decap_8 FILLER_12_734 ();
 sg13g2_decap_8 FILLER_12_741 ();
 sg13g2_decap_8 FILLER_12_748 ();
 sg13g2_decap_8 FILLER_12_755 ();
 sg13g2_decap_8 FILLER_12_762 ();
 sg13g2_decap_8 FILLER_12_769 ();
 sg13g2_decap_8 FILLER_12_776 ();
 sg13g2_decap_8 FILLER_12_783 ();
 sg13g2_decap_8 FILLER_12_790 ();
 sg13g2_decap_4 FILLER_12_797 ();
 sg13g2_fill_2 FILLER_12_801 ();
 sg13g2_decap_8 FILLER_12_807 ();
 sg13g2_decap_8 FILLER_12_814 ();
 sg13g2_decap_4 FILLER_12_821 ();
 sg13g2_fill_2 FILLER_12_825 ();
 sg13g2_decap_8 FILLER_12_853 ();
 sg13g2_fill_2 FILLER_12_860 ();
 sg13g2_decap_8 FILLER_12_866 ();
 sg13g2_decap_8 FILLER_12_873 ();
 sg13g2_decap_4 FILLER_12_880 ();
 sg13g2_decap_8 FILLER_12_888 ();
 sg13g2_decap_8 FILLER_12_895 ();
 sg13g2_decap_8 FILLER_12_902 ();
 sg13g2_decap_8 FILLER_12_909 ();
 sg13g2_decap_8 FILLER_12_916 ();
 sg13g2_decap_8 FILLER_12_923 ();
 sg13g2_decap_8 FILLER_12_930 ();
 sg13g2_decap_8 FILLER_12_937 ();
 sg13g2_decap_4 FILLER_12_944 ();
 sg13g2_fill_1 FILLER_12_948 ();
 sg13g2_decap_8 FILLER_12_953 ();
 sg13g2_decap_8 FILLER_12_960 ();
 sg13g2_decap_8 FILLER_12_967 ();
 sg13g2_decap_8 FILLER_12_974 ();
 sg13g2_decap_4 FILLER_12_981 ();
 sg13g2_decap_8 FILLER_12_993 ();
 sg13g2_decap_8 FILLER_12_1000 ();
 sg13g2_decap_8 FILLER_12_1007 ();
 sg13g2_decap_8 FILLER_12_1014 ();
 sg13g2_decap_8 FILLER_12_1021 ();
 sg13g2_decap_8 FILLER_12_1028 ();
 sg13g2_decap_8 FILLER_12_1035 ();
 sg13g2_decap_8 FILLER_12_1042 ();
 sg13g2_decap_8 FILLER_12_1049 ();
 sg13g2_decap_8 FILLER_12_1056 ();
 sg13g2_decap_8 FILLER_12_1063 ();
 sg13g2_decap_8 FILLER_12_1070 ();
 sg13g2_decap_8 FILLER_12_1077 ();
 sg13g2_decap_8 FILLER_12_1084 ();
 sg13g2_decap_8 FILLER_12_1091 ();
 sg13g2_fill_2 FILLER_12_1098 ();
 sg13g2_decap_8 FILLER_12_1114 ();
 sg13g2_decap_8 FILLER_12_1121 ();
 sg13g2_decap_8 FILLER_12_1133 ();
 sg13g2_decap_8 FILLER_12_1140 ();
 sg13g2_decap_8 FILLER_12_1147 ();
 sg13g2_decap_4 FILLER_12_1164 ();
 sg13g2_decap_4 FILLER_12_1189 ();
 sg13g2_decap_8 FILLER_12_1198 ();
 sg13g2_decap_8 FILLER_12_1205 ();
 sg13g2_decap_8 FILLER_12_1212 ();
 sg13g2_decap_8 FILLER_12_1219 ();
 sg13g2_decap_8 FILLER_12_1226 ();
 sg13g2_decap_8 FILLER_12_1233 ();
 sg13g2_decap_8 FILLER_12_1240 ();
 sg13g2_decap_8 FILLER_12_1247 ();
 sg13g2_decap_8 FILLER_12_1254 ();
 sg13g2_decap_8 FILLER_12_1261 ();
 sg13g2_decap_8 FILLER_12_1268 ();
 sg13g2_decap_8 FILLER_12_1275 ();
 sg13g2_decap_8 FILLER_12_1282 ();
 sg13g2_decap_8 FILLER_12_1289 ();
 sg13g2_decap_8 FILLER_12_1296 ();
 sg13g2_decap_8 FILLER_12_1303 ();
 sg13g2_decap_8 FILLER_12_1310 ();
 sg13g2_decap_8 FILLER_12_1317 ();
 sg13g2_fill_2 FILLER_12_1324 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_43 ();
 sg13g2_decap_8 FILLER_13_50 ();
 sg13g2_decap_8 FILLER_13_57 ();
 sg13g2_decap_8 FILLER_13_64 ();
 sg13g2_decap_4 FILLER_13_76 ();
 sg13g2_decap_8 FILLER_13_93 ();
 sg13g2_decap_4 FILLER_13_100 ();
 sg13g2_decap_4 FILLER_13_119 ();
 sg13g2_fill_1 FILLER_13_123 ();
 sg13g2_decap_4 FILLER_13_129 ();
 sg13g2_fill_1 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_142 ();
 sg13g2_decap_8 FILLER_13_149 ();
 sg13g2_fill_2 FILLER_13_156 ();
 sg13g2_fill_2 FILLER_13_172 ();
 sg13g2_fill_1 FILLER_13_174 ();
 sg13g2_fill_1 FILLER_13_190 ();
 sg13g2_fill_1 FILLER_13_207 ();
 sg13g2_decap_4 FILLER_13_216 ();
 sg13g2_fill_2 FILLER_13_231 ();
 sg13g2_fill_1 FILLER_13_236 ();
 sg13g2_decap_4 FILLER_13_241 ();
 sg13g2_fill_2 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_251 ();
 sg13g2_decap_8 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_265 ();
 sg13g2_decap_8 FILLER_13_272 ();
 sg13g2_fill_2 FILLER_13_279 ();
 sg13g2_fill_1 FILLER_13_281 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_4 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_330 ();
 sg13g2_fill_2 FILLER_13_337 ();
 sg13g2_fill_1 FILLER_13_339 ();
 sg13g2_fill_2 FILLER_13_343 ();
 sg13g2_fill_1 FILLER_13_345 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_4 FILLER_13_371 ();
 sg13g2_fill_1 FILLER_13_375 ();
 sg13g2_fill_2 FILLER_13_386 ();
 sg13g2_fill_1 FILLER_13_398 ();
 sg13g2_fill_2 FILLER_13_414 ();
 sg13g2_fill_1 FILLER_13_416 ();
 sg13g2_decap_8 FILLER_13_422 ();
 sg13g2_decap_8 FILLER_13_429 ();
 sg13g2_decap_4 FILLER_13_436 ();
 sg13g2_fill_1 FILLER_13_440 ();
 sg13g2_fill_2 FILLER_13_446 ();
 sg13g2_decap_4 FILLER_13_452 ();
 sg13g2_fill_1 FILLER_13_456 ();
 sg13g2_decap_4 FILLER_13_461 ();
 sg13g2_decap_8 FILLER_13_470 ();
 sg13g2_decap_8 FILLER_13_477 ();
 sg13g2_decap_8 FILLER_13_484 ();
 sg13g2_fill_2 FILLER_13_491 ();
 sg13g2_fill_2 FILLER_13_497 ();
 sg13g2_fill_1 FILLER_13_499 ();
 sg13g2_fill_2 FILLER_13_531 ();
 sg13g2_fill_1 FILLER_13_533 ();
 sg13g2_decap_4 FILLER_13_542 ();
 sg13g2_decap_8 FILLER_13_576 ();
 sg13g2_decap_4 FILLER_13_583 ();
 sg13g2_fill_2 FILLER_13_587 ();
 sg13g2_decap_8 FILLER_13_603 ();
 sg13g2_decap_4 FILLER_13_610 ();
 sg13g2_fill_2 FILLER_13_614 ();
 sg13g2_fill_2 FILLER_13_627 ();
 sg13g2_fill_1 FILLER_13_629 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_fill_2 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_674 ();
 sg13g2_decap_8 FILLER_13_681 ();
 sg13g2_decap_8 FILLER_13_688 ();
 sg13g2_decap_8 FILLER_13_695 ();
 sg13g2_decap_8 FILLER_13_702 ();
 sg13g2_decap_8 FILLER_13_709 ();
 sg13g2_decap_8 FILLER_13_716 ();
 sg13g2_decap_8 FILLER_13_723 ();
 sg13g2_decap_8 FILLER_13_730 ();
 sg13g2_decap_8 FILLER_13_737 ();
 sg13g2_decap_8 FILLER_13_744 ();
 sg13g2_decap_8 FILLER_13_751 ();
 sg13g2_decap_8 FILLER_13_758 ();
 sg13g2_decap_8 FILLER_13_765 ();
 sg13g2_decap_8 FILLER_13_772 ();
 sg13g2_decap_8 FILLER_13_779 ();
 sg13g2_decap_8 FILLER_13_786 ();
 sg13g2_fill_2 FILLER_13_793 ();
 sg13g2_fill_1 FILLER_13_795 ();
 sg13g2_decap_8 FILLER_13_800 ();
 sg13g2_decap_8 FILLER_13_807 ();
 sg13g2_decap_8 FILLER_13_814 ();
 sg13g2_decap_8 FILLER_13_821 ();
 sg13g2_decap_8 FILLER_13_828 ();
 sg13g2_decap_8 FILLER_13_839 ();
 sg13g2_decap_8 FILLER_13_846 ();
 sg13g2_decap_8 FILLER_13_853 ();
 sg13g2_fill_1 FILLER_13_860 ();
 sg13g2_decap_8 FILLER_13_887 ();
 sg13g2_decap_8 FILLER_13_894 ();
 sg13g2_decap_8 FILLER_13_901 ();
 sg13g2_decap_8 FILLER_13_908 ();
 sg13g2_decap_8 FILLER_13_915 ();
 sg13g2_fill_2 FILLER_13_922 ();
 sg13g2_fill_1 FILLER_13_924 ();
 sg13g2_decap_4 FILLER_13_928 ();
 sg13g2_fill_1 FILLER_13_932 ();
 sg13g2_decap_8 FILLER_13_937 ();
 sg13g2_decap_8 FILLER_13_944 ();
 sg13g2_decap_4 FILLER_13_951 ();
 sg13g2_fill_2 FILLER_13_955 ();
 sg13g2_decap_8 FILLER_13_967 ();
 sg13g2_decap_8 FILLER_13_974 ();
 sg13g2_decap_8 FILLER_13_981 ();
 sg13g2_fill_2 FILLER_13_988 ();
 sg13g2_decap_8 FILLER_13_995 ();
 sg13g2_decap_8 FILLER_13_1002 ();
 sg13g2_decap_8 FILLER_13_1009 ();
 sg13g2_decap_8 FILLER_13_1016 ();
 sg13g2_decap_8 FILLER_13_1023 ();
 sg13g2_decap_8 FILLER_13_1030 ();
 sg13g2_decap_8 FILLER_13_1037 ();
 sg13g2_fill_2 FILLER_13_1044 ();
 sg13g2_fill_1 FILLER_13_1046 ();
 sg13g2_decap_4 FILLER_13_1052 ();
 sg13g2_decap_8 FILLER_13_1060 ();
 sg13g2_decap_4 FILLER_13_1067 ();
 sg13g2_fill_2 FILLER_13_1071 ();
 sg13g2_fill_2 FILLER_13_1084 ();
 sg13g2_fill_1 FILLER_13_1086 ();
 sg13g2_decap_8 FILLER_13_1091 ();
 sg13g2_decap_4 FILLER_13_1098 ();
 sg13g2_fill_1 FILLER_13_1117 ();
 sg13g2_fill_2 FILLER_13_1122 ();
 sg13g2_decap_8 FILLER_13_1133 ();
 sg13g2_decap_8 FILLER_13_1140 ();
 sg13g2_decap_4 FILLER_13_1152 ();
 sg13g2_fill_1 FILLER_13_1156 ();
 sg13g2_decap_4 FILLER_13_1175 ();
 sg13g2_fill_2 FILLER_13_1195 ();
 sg13g2_fill_1 FILLER_13_1197 ();
 sg13g2_fill_2 FILLER_13_1205 ();
 sg13g2_decap_4 FILLER_13_1212 ();
 sg13g2_fill_1 FILLER_13_1216 ();
 sg13g2_decap_8 FILLER_13_1224 ();
 sg13g2_decap_8 FILLER_13_1231 ();
 sg13g2_decap_8 FILLER_13_1238 ();
 sg13g2_decap_8 FILLER_13_1245 ();
 sg13g2_decap_8 FILLER_13_1252 ();
 sg13g2_decap_8 FILLER_13_1259 ();
 sg13g2_decap_8 FILLER_13_1266 ();
 sg13g2_decap_8 FILLER_13_1273 ();
 sg13g2_decap_8 FILLER_13_1280 ();
 sg13g2_decap_8 FILLER_13_1287 ();
 sg13g2_decap_8 FILLER_13_1294 ();
 sg13g2_decap_8 FILLER_13_1301 ();
 sg13g2_decap_8 FILLER_13_1308 ();
 sg13g2_decap_8 FILLER_13_1315 ();
 sg13g2_decap_4 FILLER_13_1322 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_4 FILLER_14_105 ();
 sg13g2_fill_2 FILLER_14_109 ();
 sg13g2_decap_8 FILLER_14_125 ();
 sg13g2_decap_8 FILLER_14_132 ();
 sg13g2_decap_8 FILLER_14_139 ();
 sg13g2_decap_8 FILLER_14_146 ();
 sg13g2_decap_8 FILLER_14_153 ();
 sg13g2_decap_8 FILLER_14_160 ();
 sg13g2_decap_8 FILLER_14_171 ();
 sg13g2_decap_8 FILLER_14_178 ();
 sg13g2_decap_8 FILLER_14_185 ();
 sg13g2_decap_8 FILLER_14_192 ();
 sg13g2_decap_8 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_decap_4 FILLER_14_213 ();
 sg13g2_fill_1 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_226 ();
 sg13g2_decap_8 FILLER_14_233 ();
 sg13g2_decap_4 FILLER_14_240 ();
 sg13g2_fill_2 FILLER_14_244 ();
 sg13g2_decap_8 FILLER_14_251 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_decap_8 FILLER_14_267 ();
 sg13g2_decap_8 FILLER_14_274 ();
 sg13g2_decap_8 FILLER_14_281 ();
 sg13g2_decap_8 FILLER_14_288 ();
 sg13g2_decap_8 FILLER_14_295 ();
 sg13g2_decap_4 FILLER_14_302 ();
 sg13g2_fill_2 FILLER_14_306 ();
 sg13g2_decap_8 FILLER_14_321 ();
 sg13g2_decap_8 FILLER_14_328 ();
 sg13g2_decap_8 FILLER_14_335 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_356 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_4 FILLER_14_377 ();
 sg13g2_fill_2 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_400 ();
 sg13g2_decap_8 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_14_414 ();
 sg13g2_fill_2 FILLER_14_421 ();
 sg13g2_fill_1 FILLER_14_423 ();
 sg13g2_decap_8 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_14_436 ();
 sg13g2_fill_1 FILLER_14_443 ();
 sg13g2_decap_8 FILLER_14_449 ();
 sg13g2_decap_8 FILLER_14_456 ();
 sg13g2_decap_8 FILLER_14_463 ();
 sg13g2_decap_8 FILLER_14_470 ();
 sg13g2_decap_8 FILLER_14_477 ();
 sg13g2_decap_8 FILLER_14_484 ();
 sg13g2_decap_8 FILLER_14_491 ();
 sg13g2_decap_8 FILLER_14_498 ();
 sg13g2_decap_8 FILLER_14_505 ();
 sg13g2_decap_8 FILLER_14_512 ();
 sg13g2_decap_8 FILLER_14_519 ();
 sg13g2_decap_8 FILLER_14_526 ();
 sg13g2_decap_8 FILLER_14_533 ();
 sg13g2_decap_8 FILLER_14_540 ();
 sg13g2_fill_1 FILLER_14_547 ();
 sg13g2_fill_1 FILLER_14_552 ();
 sg13g2_decap_8 FILLER_14_562 ();
 sg13g2_decap_8 FILLER_14_569 ();
 sg13g2_decap_8 FILLER_14_576 ();
 sg13g2_decap_8 FILLER_14_583 ();
 sg13g2_decap_8 FILLER_14_590 ();
 sg13g2_decap_8 FILLER_14_597 ();
 sg13g2_decap_8 FILLER_14_604 ();
 sg13g2_decap_8 FILLER_14_611 ();
 sg13g2_decap_8 FILLER_14_618 ();
 sg13g2_decap_8 FILLER_14_625 ();
 sg13g2_decap_8 FILLER_14_632 ();
 sg13g2_decap_8 FILLER_14_639 ();
 sg13g2_decap_8 FILLER_14_646 ();
 sg13g2_fill_2 FILLER_14_653 ();
 sg13g2_decap_4 FILLER_14_675 ();
 sg13g2_fill_2 FILLER_14_679 ();
 sg13g2_decap_4 FILLER_14_711 ();
 sg13g2_fill_1 FILLER_14_715 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_4 FILLER_14_798 ();
 sg13g2_fill_2 FILLER_14_802 ();
 sg13g2_decap_8 FILLER_14_830 ();
 sg13g2_fill_2 FILLER_14_837 ();
 sg13g2_fill_1 FILLER_14_839 ();
 sg13g2_decap_8 FILLER_14_848 ();
 sg13g2_decap_8 FILLER_14_855 ();
 sg13g2_decap_4 FILLER_14_862 ();
 sg13g2_fill_2 FILLER_14_866 ();
 sg13g2_decap_8 FILLER_14_872 ();
 sg13g2_decap_8 FILLER_14_879 ();
 sg13g2_decap_8 FILLER_14_886 ();
 sg13g2_decap_8 FILLER_14_893 ();
 sg13g2_decap_8 FILLER_14_900 ();
 sg13g2_decap_8 FILLER_14_907 ();
 sg13g2_fill_1 FILLER_14_914 ();
 sg13g2_decap_4 FILLER_14_920 ();
 sg13g2_fill_1 FILLER_14_924 ();
 sg13g2_decap_8 FILLER_14_951 ();
 sg13g2_decap_8 FILLER_14_970 ();
 sg13g2_decap_8 FILLER_14_977 ();
 sg13g2_decap_8 FILLER_14_984 ();
 sg13g2_decap_8 FILLER_14_999 ();
 sg13g2_decap_8 FILLER_14_1006 ();
 sg13g2_decap_4 FILLER_14_1013 ();
 sg13g2_fill_2 FILLER_14_1017 ();
 sg13g2_decap_8 FILLER_14_1024 ();
 sg13g2_decap_8 FILLER_14_1031 ();
 sg13g2_decap_8 FILLER_14_1043 ();
 sg13g2_decap_8 FILLER_14_1053 ();
 sg13g2_fill_1 FILLER_14_1060 ();
 sg13g2_decap_8 FILLER_14_1069 ();
 sg13g2_decap_4 FILLER_14_1076 ();
 sg13g2_decap_8 FILLER_14_1093 ();
 sg13g2_fill_1 FILLER_14_1104 ();
 sg13g2_fill_2 FILLER_14_1109 ();
 sg13g2_decap_4 FILLER_14_1116 ();
 sg13g2_decap_8 FILLER_14_1130 ();
 sg13g2_fill_1 FILLER_14_1141 ();
 sg13g2_fill_2 FILLER_14_1147 ();
 sg13g2_fill_1 FILLER_14_1149 ();
 sg13g2_fill_1 FILLER_14_1166 ();
 sg13g2_fill_2 FILLER_14_1172 ();
 sg13g2_fill_1 FILLER_14_1178 ();
 sg13g2_decap_4 FILLER_14_1184 ();
 sg13g2_fill_2 FILLER_14_1193 ();
 sg13g2_fill_1 FILLER_14_1200 ();
 sg13g2_decap_4 FILLER_14_1206 ();
 sg13g2_fill_1 FILLER_14_1210 ();
 sg13g2_fill_1 FILLER_14_1216 ();
 sg13g2_decap_8 FILLER_14_1232 ();
 sg13g2_decap_8 FILLER_14_1239 ();
 sg13g2_decap_8 FILLER_14_1246 ();
 sg13g2_decap_8 FILLER_14_1253 ();
 sg13g2_decap_8 FILLER_14_1260 ();
 sg13g2_decap_8 FILLER_14_1267 ();
 sg13g2_decap_8 FILLER_14_1274 ();
 sg13g2_decap_8 FILLER_14_1281 ();
 sg13g2_decap_8 FILLER_14_1288 ();
 sg13g2_decap_8 FILLER_14_1295 ();
 sg13g2_decap_8 FILLER_14_1302 ();
 sg13g2_decap_8 FILLER_14_1309 ();
 sg13g2_decap_8 FILLER_14_1316 ();
 sg13g2_fill_2 FILLER_14_1323 ();
 sg13g2_fill_1 FILLER_14_1325 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_64 ();
 sg13g2_decap_8 FILLER_15_71 ();
 sg13g2_decap_8 FILLER_15_78 ();
 sg13g2_decap_8 FILLER_15_85 ();
 sg13g2_decap_8 FILLER_15_92 ();
 sg13g2_decap_8 FILLER_15_99 ();
 sg13g2_decap_4 FILLER_15_106 ();
 sg13g2_fill_2 FILLER_15_110 ();
 sg13g2_decap_4 FILLER_15_117 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_fill_2 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_173 ();
 sg13g2_decap_8 FILLER_15_180 ();
 sg13g2_decap_8 FILLER_15_187 ();
 sg13g2_decap_8 FILLER_15_194 ();
 sg13g2_decap_8 FILLER_15_201 ();
 sg13g2_decap_8 FILLER_15_208 ();
 sg13g2_decap_4 FILLER_15_215 ();
 sg13g2_decap_8 FILLER_15_223 ();
 sg13g2_decap_8 FILLER_15_230 ();
 sg13g2_decap_4 FILLER_15_247 ();
 sg13g2_fill_2 FILLER_15_251 ();
 sg13g2_decap_8 FILLER_15_268 ();
 sg13g2_decap_8 FILLER_15_275 ();
 sg13g2_fill_2 FILLER_15_282 ();
 sg13g2_fill_1 FILLER_15_284 ();
 sg13g2_decap_4 FILLER_15_290 ();
 sg13g2_fill_1 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_305 ();
 sg13g2_fill_2 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_fill_2 FILLER_15_357 ();
 sg13g2_fill_1 FILLER_15_359 ();
 sg13g2_fill_1 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_decap_8 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_15_414 ();
 sg13g2_decap_8 FILLER_15_421 ();
 sg13g2_decap_8 FILLER_15_428 ();
 sg13g2_fill_1 FILLER_15_435 ();
 sg13g2_fill_1 FILLER_15_444 ();
 sg13g2_decap_8 FILLER_15_450 ();
 sg13g2_decap_8 FILLER_15_457 ();
 sg13g2_decap_4 FILLER_15_464 ();
 sg13g2_fill_2 FILLER_15_468 ();
 sg13g2_decap_4 FILLER_15_484 ();
 sg13g2_fill_2 FILLER_15_488 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_4 FILLER_15_651 ();
 sg13g2_fill_2 FILLER_15_655 ();
 sg13g2_fill_1 FILLER_15_662 ();
 sg13g2_decap_4 FILLER_15_676 ();
 sg13g2_fill_1 FILLER_15_680 ();
 sg13g2_fill_1 FILLER_15_686 ();
 sg13g2_fill_2 FILLER_15_692 ();
 sg13g2_decap_8 FILLER_15_708 ();
 sg13g2_decap_8 FILLER_15_715 ();
 sg13g2_decap_8 FILLER_15_726 ();
 sg13g2_decap_8 FILLER_15_733 ();
 sg13g2_decap_8 FILLER_15_740 ();
 sg13g2_decap_8 FILLER_15_747 ();
 sg13g2_fill_2 FILLER_15_754 ();
 sg13g2_fill_1 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_fill_1 FILLER_15_805 ();
 sg13g2_fill_2 FILLER_15_810 ();
 sg13g2_fill_1 FILLER_15_816 ();
 sg13g2_decap_8 FILLER_15_820 ();
 sg13g2_decap_8 FILLER_15_827 ();
 sg13g2_decap_8 FILLER_15_834 ();
 sg13g2_decap_8 FILLER_15_841 ();
 sg13g2_decap_8 FILLER_15_848 ();
 sg13g2_decap_8 FILLER_15_855 ();
 sg13g2_decap_8 FILLER_15_862 ();
 sg13g2_decap_8 FILLER_15_869 ();
 sg13g2_decap_8 FILLER_15_876 ();
 sg13g2_decap_8 FILLER_15_883 ();
 sg13g2_decap_8 FILLER_15_890 ();
 sg13g2_decap_8 FILLER_15_897 ();
 sg13g2_fill_2 FILLER_15_904 ();
 sg13g2_fill_1 FILLER_15_906 ();
 sg13g2_fill_1 FILLER_15_912 ();
 sg13g2_decap_4 FILLER_15_937 ();
 sg13g2_fill_1 FILLER_15_941 ();
 sg13g2_decap_8 FILLER_15_946 ();
 sg13g2_decap_4 FILLER_15_953 ();
 sg13g2_fill_2 FILLER_15_957 ();
 sg13g2_decap_8 FILLER_15_969 ();
 sg13g2_decap_8 FILLER_15_976 ();
 sg13g2_decap_8 FILLER_15_983 ();
 sg13g2_decap_8 FILLER_15_990 ();
 sg13g2_fill_2 FILLER_15_997 ();
 sg13g2_fill_1 FILLER_15_999 ();
 sg13g2_decap_8 FILLER_15_1014 ();
 sg13g2_fill_2 FILLER_15_1021 ();
 sg13g2_fill_2 FILLER_15_1027 ();
 sg13g2_fill_1 FILLER_15_1033 ();
 sg13g2_fill_2 FILLER_15_1051 ();
 sg13g2_fill_2 FILLER_15_1065 ();
 sg13g2_fill_2 FILLER_15_1076 ();
 sg13g2_decap_8 FILLER_15_1082 ();
 sg13g2_fill_1 FILLER_15_1089 ();
 sg13g2_decap_8 FILLER_15_1098 ();
 sg13g2_fill_1 FILLER_15_1105 ();
 sg13g2_fill_2 FILLER_15_1116 ();
 sg13g2_decap_8 FILLER_15_1122 ();
 sg13g2_decap_8 FILLER_15_1129 ();
 sg13g2_decap_8 FILLER_15_1136 ();
 sg13g2_decap_8 FILLER_15_1143 ();
 sg13g2_decap_8 FILLER_15_1150 ();
 sg13g2_decap_8 FILLER_15_1157 ();
 sg13g2_decap_8 FILLER_15_1164 ();
 sg13g2_decap_8 FILLER_15_1171 ();
 sg13g2_fill_2 FILLER_15_1178 ();
 sg13g2_decap_8 FILLER_15_1184 ();
 sg13g2_decap_8 FILLER_15_1191 ();
 sg13g2_decap_8 FILLER_15_1198 ();
 sg13g2_decap_8 FILLER_15_1205 ();
 sg13g2_decap_8 FILLER_15_1212 ();
 sg13g2_decap_4 FILLER_15_1219 ();
 sg13g2_decap_4 FILLER_15_1232 ();
 sg13g2_fill_1 FILLER_15_1236 ();
 sg13g2_decap_8 FILLER_15_1242 ();
 sg13g2_decap_8 FILLER_15_1249 ();
 sg13g2_decap_8 FILLER_15_1256 ();
 sg13g2_decap_8 FILLER_15_1263 ();
 sg13g2_decap_8 FILLER_15_1270 ();
 sg13g2_decap_8 FILLER_15_1277 ();
 sg13g2_decap_8 FILLER_15_1284 ();
 sg13g2_decap_8 FILLER_15_1291 ();
 sg13g2_decap_8 FILLER_15_1298 ();
 sg13g2_decap_8 FILLER_15_1305 ();
 sg13g2_decap_8 FILLER_15_1312 ();
 sg13g2_decap_8 FILLER_15_1319 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_4 FILLER_16_31 ();
 sg13g2_decap_8 FILLER_16_60 ();
 sg13g2_decap_8 FILLER_16_67 ();
 sg13g2_decap_8 FILLER_16_74 ();
 sg13g2_decap_8 FILLER_16_81 ();
 sg13g2_decap_4 FILLER_16_88 ();
 sg13g2_fill_1 FILLER_16_92 ();
 sg13g2_fill_1 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_116 ();
 sg13g2_fill_2 FILLER_16_121 ();
 sg13g2_fill_1 FILLER_16_123 ();
 sg13g2_decap_8 FILLER_16_128 ();
 sg13g2_decap_8 FILLER_16_144 ();
 sg13g2_decap_8 FILLER_16_151 ();
 sg13g2_fill_1 FILLER_16_163 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_fill_1 FILLER_16_220 ();
 sg13g2_fill_2 FILLER_16_226 ();
 sg13g2_fill_2 FILLER_16_235 ();
 sg13g2_fill_1 FILLER_16_237 ();
 sg13g2_decap_8 FILLER_16_253 ();
 sg13g2_decap_8 FILLER_16_260 ();
 sg13g2_decap_8 FILLER_16_267 ();
 sg13g2_decap_4 FILLER_16_274 ();
 sg13g2_decap_8 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_316 ();
 sg13g2_decap_4 FILLER_16_323 ();
 sg13g2_decap_8 FILLER_16_337 ();
 sg13g2_fill_1 FILLER_16_344 ();
 sg13g2_fill_1 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_decap_8 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_16_415 ();
 sg13g2_decap_8 FILLER_16_422 ();
 sg13g2_fill_2 FILLER_16_429 ();
 sg13g2_decap_4 FILLER_16_462 ();
 sg13g2_fill_1 FILLER_16_466 ();
 sg13g2_decap_4 FILLER_16_471 ();
 sg13g2_fill_2 FILLER_16_492 ();
 sg13g2_decap_8 FILLER_16_499 ();
 sg13g2_decap_4 FILLER_16_506 ();
 sg13g2_decap_8 FILLER_16_514 ();
 sg13g2_decap_8 FILLER_16_526 ();
 sg13g2_decap_8 FILLER_16_533 ();
 sg13g2_decap_4 FILLER_16_540 ();
 sg13g2_decap_8 FILLER_16_570 ();
 sg13g2_decap_8 FILLER_16_577 ();
 sg13g2_decap_8 FILLER_16_584 ();
 sg13g2_fill_2 FILLER_16_591 ();
 sg13g2_decap_8 FILLER_16_619 ();
 sg13g2_decap_8 FILLER_16_633 ();
 sg13g2_decap_8 FILLER_16_640 ();
 sg13g2_fill_2 FILLER_16_647 ();
 sg13g2_fill_1 FILLER_16_649 ();
 sg13g2_decap_4 FILLER_16_663 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_fill_1 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_699 ();
 sg13g2_decap_4 FILLER_16_706 ();
 sg13g2_fill_1 FILLER_16_710 ();
 sg13g2_decap_8 FILLER_16_715 ();
 sg13g2_decap_8 FILLER_16_722 ();
 sg13g2_decap_8 FILLER_16_729 ();
 sg13g2_decap_8 FILLER_16_736 ();
 sg13g2_decap_8 FILLER_16_743 ();
 sg13g2_decap_8 FILLER_16_750 ();
 sg13g2_decap_4 FILLER_16_757 ();
 sg13g2_fill_2 FILLER_16_761 ();
 sg13g2_decap_8 FILLER_16_767 ();
 sg13g2_fill_2 FILLER_16_774 ();
 sg13g2_fill_1 FILLER_16_806 ();
 sg13g2_decap_8 FILLER_16_815 ();
 sg13g2_fill_1 FILLER_16_822 ();
 sg13g2_decap_8 FILLER_16_853 ();
 sg13g2_decap_8 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_16_867 ();
 sg13g2_decap_8 FILLER_16_878 ();
 sg13g2_decap_8 FILLER_16_885 ();
 sg13g2_decap_8 FILLER_16_892 ();
 sg13g2_decap_8 FILLER_16_899 ();
 sg13g2_decap_8 FILLER_16_906 ();
 sg13g2_decap_8 FILLER_16_913 ();
 sg13g2_fill_2 FILLER_16_920 ();
 sg13g2_fill_1 FILLER_16_922 ();
 sg13g2_decap_8 FILLER_16_931 ();
 sg13g2_decap_8 FILLER_16_938 ();
 sg13g2_decap_8 FILLER_16_945 ();
 sg13g2_decap_8 FILLER_16_952 ();
 sg13g2_decap_8 FILLER_16_959 ();
 sg13g2_decap_8 FILLER_16_966 ();
 sg13g2_decap_4 FILLER_16_973 ();
 sg13g2_decap_8 FILLER_16_985 ();
 sg13g2_decap_8 FILLER_16_992 ();
 sg13g2_decap_8 FILLER_16_999 ();
 sg13g2_decap_8 FILLER_16_1014 ();
 sg13g2_decap_4 FILLER_16_1021 ();
 sg13g2_decap_8 FILLER_16_1029 ();
 sg13g2_decap_8 FILLER_16_1036 ();
 sg13g2_fill_2 FILLER_16_1043 ();
 sg13g2_fill_1 FILLER_16_1050 ();
 sg13g2_decap_4 FILLER_16_1056 ();
 sg13g2_fill_1 FILLER_16_1060 ();
 sg13g2_decap_8 FILLER_16_1070 ();
 sg13g2_fill_1 FILLER_16_1077 ();
 sg13g2_decap_8 FILLER_16_1100 ();
 sg13g2_decap_8 FILLER_16_1107 ();
 sg13g2_decap_4 FILLER_16_1114 ();
 sg13g2_fill_1 FILLER_16_1118 ();
 sg13g2_decap_8 FILLER_16_1123 ();
 sg13g2_decap_8 FILLER_16_1130 ();
 sg13g2_decap_8 FILLER_16_1137 ();
 sg13g2_decap_8 FILLER_16_1144 ();
 sg13g2_fill_2 FILLER_16_1151 ();
 sg13g2_fill_1 FILLER_16_1153 ();
 sg13g2_decap_8 FILLER_16_1158 ();
 sg13g2_fill_2 FILLER_16_1169 ();
 sg13g2_decap_8 FILLER_16_1175 ();
 sg13g2_fill_2 FILLER_16_1182 ();
 sg13g2_fill_1 FILLER_16_1184 ();
 sg13g2_decap_8 FILLER_16_1193 ();
 sg13g2_decap_8 FILLER_16_1200 ();
 sg13g2_decap_8 FILLER_16_1207 ();
 sg13g2_decap_8 FILLER_16_1214 ();
 sg13g2_decap_4 FILLER_16_1221 ();
 sg13g2_fill_1 FILLER_16_1229 ();
 sg13g2_fill_2 FILLER_16_1244 ();
 sg13g2_decap_8 FILLER_16_1249 ();
 sg13g2_decap_8 FILLER_16_1256 ();
 sg13g2_decap_8 FILLER_16_1263 ();
 sg13g2_decap_8 FILLER_16_1270 ();
 sg13g2_decap_8 FILLER_16_1277 ();
 sg13g2_decap_8 FILLER_16_1284 ();
 sg13g2_decap_8 FILLER_16_1291 ();
 sg13g2_decap_8 FILLER_16_1298 ();
 sg13g2_decap_8 FILLER_16_1305 ();
 sg13g2_decap_8 FILLER_16_1312 ();
 sg13g2_decap_8 FILLER_16_1319 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_27 ();
 sg13g2_decap_4 FILLER_17_33 ();
 sg13g2_fill_2 FILLER_17_37 ();
 sg13g2_fill_2 FILLER_17_47 ();
 sg13g2_fill_1 FILLER_17_49 ();
 sg13g2_fill_1 FILLER_17_59 ();
 sg13g2_fill_2 FILLER_17_66 ();
 sg13g2_fill_1 FILLER_17_82 ();
 sg13g2_fill_2 FILLER_17_88 ();
 sg13g2_fill_1 FILLER_17_90 ();
 sg13g2_fill_2 FILLER_17_104 ();
 sg13g2_decap_8 FILLER_17_123 ();
 sg13g2_fill_2 FILLER_17_130 ();
 sg13g2_fill_1 FILLER_17_132 ();
 sg13g2_fill_1 FILLER_17_141 ();
 sg13g2_decap_8 FILLER_17_174 ();
 sg13g2_decap_8 FILLER_17_181 ();
 sg13g2_decap_8 FILLER_17_188 ();
 sg13g2_decap_8 FILLER_17_195 ();
 sg13g2_decap_8 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_216 ();
 sg13g2_fill_1 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_234 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_4 FILLER_17_273 ();
 sg13g2_fill_1 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_313 ();
 sg13g2_decap_4 FILLER_17_348 ();
 sg13g2_fill_1 FILLER_17_352 ();
 sg13g2_fill_1 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_8 FILLER_17_404 ();
 sg13g2_decap_8 FILLER_17_411 ();
 sg13g2_decap_8 FILLER_17_418 ();
 sg13g2_decap_8 FILLER_17_425 ();
 sg13g2_decap_4 FILLER_17_432 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_453 ();
 sg13g2_decap_8 FILLER_17_460 ();
 sg13g2_fill_2 FILLER_17_467 ();
 sg13g2_fill_1 FILLER_17_469 ();
 sg13g2_decap_4 FILLER_17_506 ();
 sg13g2_fill_2 FILLER_17_520 ();
 sg13g2_fill_1 FILLER_17_537 ();
 sg13g2_decap_8 FILLER_17_543 ();
 sg13g2_fill_1 FILLER_17_550 ();
 sg13g2_fill_1 FILLER_17_555 ();
 sg13g2_decap_8 FILLER_17_582 ();
 sg13g2_fill_2 FILLER_17_603 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_fill_2 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_4 FILLER_17_679 ();
 sg13g2_fill_2 FILLER_17_683 ();
 sg13g2_decap_8 FILLER_17_697 ();
 sg13g2_fill_1 FILLER_17_704 ();
 sg13g2_decap_8 FILLER_17_731 ();
 sg13g2_decap_4 FILLER_17_738 ();
 sg13g2_fill_2 FILLER_17_742 ();
 sg13g2_fill_2 FILLER_17_752 ();
 sg13g2_fill_1 FILLER_17_754 ();
 sg13g2_decap_8 FILLER_17_758 ();
 sg13g2_decap_4 FILLER_17_765 ();
 sg13g2_fill_2 FILLER_17_769 ();
 sg13g2_fill_1 FILLER_17_783 ();
 sg13g2_decap_8 FILLER_17_797 ();
 sg13g2_decap_4 FILLER_17_804 ();
 sg13g2_fill_2 FILLER_17_818 ();
 sg13g2_decap_4 FILLER_17_828 ();
 sg13g2_fill_1 FILLER_17_832 ();
 sg13g2_decap_8 FILLER_17_837 ();
 sg13g2_decap_8 FILLER_17_844 ();
 sg13g2_decap_8 FILLER_17_851 ();
 sg13g2_fill_2 FILLER_17_858 ();
 sg13g2_fill_1 FILLER_17_864 ();
 sg13g2_decap_8 FILLER_17_895 ();
 sg13g2_decap_8 FILLER_17_902 ();
 sg13g2_fill_2 FILLER_17_909 ();
 sg13g2_decap_8 FILLER_17_915 ();
 sg13g2_fill_2 FILLER_17_922 ();
 sg13g2_fill_1 FILLER_17_924 ();
 sg13g2_fill_1 FILLER_17_929 ();
 sg13g2_decap_8 FILLER_17_934 ();
 sg13g2_fill_1 FILLER_17_956 ();
 sg13g2_fill_2 FILLER_17_978 ();
 sg13g2_fill_1 FILLER_17_980 ();
 sg13g2_fill_2 FILLER_17_986 ();
 sg13g2_fill_1 FILLER_17_988 ();
 sg13g2_decap_8 FILLER_17_994 ();
 sg13g2_decap_8 FILLER_17_1001 ();
 sg13g2_decap_8 FILLER_17_1008 ();
 sg13g2_decap_8 FILLER_17_1015 ();
 sg13g2_fill_2 FILLER_17_1022 ();
 sg13g2_fill_1 FILLER_17_1024 ();
 sg13g2_decap_4 FILLER_17_1030 ();
 sg13g2_decap_8 FILLER_17_1038 ();
 sg13g2_decap_8 FILLER_17_1045 ();
 sg13g2_decap_8 FILLER_17_1052 ();
 sg13g2_decap_4 FILLER_17_1059 ();
 sg13g2_fill_2 FILLER_17_1073 ();
 sg13g2_fill_1 FILLER_17_1075 ();
 sg13g2_decap_8 FILLER_17_1080 ();
 sg13g2_fill_1 FILLER_17_1092 ();
 sg13g2_decap_8 FILLER_17_1097 ();
 sg13g2_decap_8 FILLER_17_1104 ();
 sg13g2_decap_4 FILLER_17_1111 ();
 sg13g2_decap_8 FILLER_17_1124 ();
 sg13g2_decap_8 FILLER_17_1131 ();
 sg13g2_decap_4 FILLER_17_1138 ();
 sg13g2_fill_2 FILLER_17_1142 ();
 sg13g2_decap_4 FILLER_17_1148 ();
 sg13g2_fill_2 FILLER_17_1166 ();
 sg13g2_fill_1 FILLER_17_1168 ();
 sg13g2_fill_2 FILLER_17_1179 ();
 sg13g2_decap_8 FILLER_17_1185 ();
 sg13g2_fill_2 FILLER_17_1192 ();
 sg13g2_decap_8 FILLER_17_1199 ();
 sg13g2_decap_8 FILLER_17_1206 ();
 sg13g2_decap_8 FILLER_17_1213 ();
 sg13g2_decap_4 FILLER_17_1220 ();
 sg13g2_fill_1 FILLER_17_1224 ();
 sg13g2_fill_1 FILLER_17_1230 ();
 sg13g2_fill_2 FILLER_17_1235 ();
 sg13g2_fill_2 FILLER_17_1247 ();
 sg13g2_fill_1 FILLER_17_1249 ();
 sg13g2_fill_2 FILLER_17_1254 ();
 sg13g2_decap_4 FILLER_17_1264 ();
 sg13g2_fill_2 FILLER_17_1268 ();
 sg13g2_decap_8 FILLER_17_1275 ();
 sg13g2_decap_8 FILLER_17_1282 ();
 sg13g2_decap_8 FILLER_17_1289 ();
 sg13g2_decap_8 FILLER_17_1296 ();
 sg13g2_decap_8 FILLER_17_1303 ();
 sg13g2_decap_8 FILLER_17_1310 ();
 sg13g2_decap_8 FILLER_17_1317 ();
 sg13g2_fill_2 FILLER_17_1324 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_4 FILLER_18_35 ();
 sg13g2_fill_2 FILLER_18_39 ();
 sg13g2_fill_2 FILLER_18_44 ();
 sg13g2_fill_1 FILLER_18_46 ();
 sg13g2_decap_8 FILLER_18_52 ();
 sg13g2_decap_8 FILLER_18_59 ();
 sg13g2_decap_8 FILLER_18_66 ();
 sg13g2_decap_8 FILLER_18_73 ();
 sg13g2_decap_8 FILLER_18_80 ();
 sg13g2_decap_4 FILLER_18_87 ();
 sg13g2_fill_2 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_115 ();
 sg13g2_decap_8 FILLER_18_122 ();
 sg13g2_decap_8 FILLER_18_129 ();
 sg13g2_decap_8 FILLER_18_136 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_decap_8 FILLER_18_150 ();
 sg13g2_decap_4 FILLER_18_157 ();
 sg13g2_decap_8 FILLER_18_177 ();
 sg13g2_decap_8 FILLER_18_184 ();
 sg13g2_decap_8 FILLER_18_191 ();
 sg13g2_decap_8 FILLER_18_198 ();
 sg13g2_decap_8 FILLER_18_205 ();
 sg13g2_decap_8 FILLER_18_212 ();
 sg13g2_decap_8 FILLER_18_219 ();
 sg13g2_decap_8 FILLER_18_226 ();
 sg13g2_decap_8 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_240 ();
 sg13g2_decap_4 FILLER_18_247 ();
 sg13g2_fill_2 FILLER_18_251 ();
 sg13g2_decap_8 FILLER_18_257 ();
 sg13g2_decap_8 FILLER_18_264 ();
 sg13g2_decap_8 FILLER_18_271 ();
 sg13g2_decap_8 FILLER_18_278 ();
 sg13g2_decap_4 FILLER_18_285 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_decap_8 FILLER_18_300 ();
 sg13g2_decap_8 FILLER_18_307 ();
 sg13g2_decap_4 FILLER_18_314 ();
 sg13g2_fill_2 FILLER_18_318 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_fill_2 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_8 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_18_412 ();
 sg13g2_decap_8 FILLER_18_419 ();
 sg13g2_decap_8 FILLER_18_426 ();
 sg13g2_decap_4 FILLER_18_433 ();
 sg13g2_fill_1 FILLER_18_437 ();
 sg13g2_decap_4 FILLER_18_443 ();
 sg13g2_fill_1 FILLER_18_447 ();
 sg13g2_fill_2 FILLER_18_453 ();
 sg13g2_decap_8 FILLER_18_460 ();
 sg13g2_fill_2 FILLER_18_467 ();
 sg13g2_decap_4 FILLER_18_473 ();
 sg13g2_fill_2 FILLER_18_482 ();
 sg13g2_decap_8 FILLER_18_487 ();
 sg13g2_decap_8 FILLER_18_494 ();
 sg13g2_decap_8 FILLER_18_501 ();
 sg13g2_decap_8 FILLER_18_508 ();
 sg13g2_decap_8 FILLER_18_515 ();
 sg13g2_decap_8 FILLER_18_522 ();
 sg13g2_decap_8 FILLER_18_529 ();
 sg13g2_decap_8 FILLER_18_536 ();
 sg13g2_fill_2 FILLER_18_547 ();
 sg13g2_fill_1 FILLER_18_554 ();
 sg13g2_fill_2 FILLER_18_564 ();
 sg13g2_fill_1 FILLER_18_566 ();
 sg13g2_decap_8 FILLER_18_571 ();
 sg13g2_decap_8 FILLER_18_578 ();
 sg13g2_decap_8 FILLER_18_585 ();
 sg13g2_fill_1 FILLER_18_592 ();
 sg13g2_fill_1 FILLER_18_607 ();
 sg13g2_decap_8 FILLER_18_612 ();
 sg13g2_decap_8 FILLER_18_619 ();
 sg13g2_decap_8 FILLER_18_626 ();
 sg13g2_decap_8 FILLER_18_633 ();
 sg13g2_decap_4 FILLER_18_640 ();
 sg13g2_fill_2 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_671 ();
 sg13g2_decap_8 FILLER_18_678 ();
 sg13g2_decap_8 FILLER_18_685 ();
 sg13g2_decap_8 FILLER_18_718 ();
 sg13g2_decap_8 FILLER_18_725 ();
 sg13g2_decap_4 FILLER_18_732 ();
 sg13g2_fill_1 FILLER_18_736 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_fill_1 FILLER_18_784 ();
 sg13g2_decap_4 FILLER_18_789 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_4 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_821 ();
 sg13g2_decap_8 FILLER_18_828 ();
 sg13g2_decap_8 FILLER_18_835 ();
 sg13g2_decap_8 FILLER_18_842 ();
 sg13g2_fill_2 FILLER_18_849 ();
 sg13g2_decap_8 FILLER_18_866 ();
 sg13g2_decap_8 FILLER_18_873 ();
 sg13g2_decap_8 FILLER_18_880 ();
 sg13g2_decap_8 FILLER_18_887 ();
 sg13g2_decap_8 FILLER_18_894 ();
 sg13g2_decap_8 FILLER_18_901 ();
 sg13g2_decap_8 FILLER_18_908 ();
 sg13g2_decap_8 FILLER_18_915 ();
 sg13g2_decap_8 FILLER_18_922 ();
 sg13g2_fill_2 FILLER_18_929 ();
 sg13g2_fill_1 FILLER_18_936 ();
 sg13g2_fill_2 FILLER_18_941 ();
 sg13g2_fill_1 FILLER_18_943 ();
 sg13g2_fill_1 FILLER_18_949 ();
 sg13g2_fill_1 FILLER_18_966 ();
 sg13g2_fill_2 FILLER_18_983 ();
 sg13g2_fill_1 FILLER_18_985 ();
 sg13g2_decap_8 FILLER_18_990 ();
 sg13g2_decap_4 FILLER_18_997 ();
 sg13g2_fill_1 FILLER_18_1001 ();
 sg13g2_fill_1 FILLER_18_1011 ();
 sg13g2_decap_4 FILLER_18_1017 ();
 sg13g2_fill_2 FILLER_18_1021 ();
 sg13g2_decap_4 FILLER_18_1028 ();
 sg13g2_fill_2 FILLER_18_1032 ();
 sg13g2_decap_4 FILLER_18_1039 ();
 sg13g2_decap_8 FILLER_18_1058 ();
 sg13g2_decap_8 FILLER_18_1065 ();
 sg13g2_decap_8 FILLER_18_1072 ();
 sg13g2_fill_2 FILLER_18_1079 ();
 sg13g2_decap_8 FILLER_18_1086 ();
 sg13g2_fill_1 FILLER_18_1093 ();
 sg13g2_decap_4 FILLER_18_1100 ();
 sg13g2_fill_2 FILLER_18_1104 ();
 sg13g2_fill_1 FILLER_18_1115 ();
 sg13g2_fill_2 FILLER_18_1121 ();
 sg13g2_decap_4 FILLER_18_1132 ();
 sg13g2_decap_8 FILLER_18_1141 ();
 sg13g2_fill_2 FILLER_18_1148 ();
 sg13g2_decap_8 FILLER_18_1159 ();
 sg13g2_decap_4 FILLER_18_1174 ();
 sg13g2_fill_1 FILLER_18_1178 ();
 sg13g2_decap_4 FILLER_18_1183 ();
 sg13g2_decap_8 FILLER_18_1212 ();
 sg13g2_decap_4 FILLER_18_1219 ();
 sg13g2_fill_1 FILLER_18_1223 ();
 sg13g2_decap_4 FILLER_18_1229 ();
 sg13g2_fill_1 FILLER_18_1233 ();
 sg13g2_decap_8 FILLER_18_1244 ();
 sg13g2_decap_8 FILLER_18_1251 ();
 sg13g2_fill_1 FILLER_18_1258 ();
 sg13g2_fill_2 FILLER_18_1262 ();
 sg13g2_decap_8 FILLER_18_1281 ();
 sg13g2_decap_8 FILLER_18_1288 ();
 sg13g2_decap_8 FILLER_18_1295 ();
 sg13g2_decap_8 FILLER_18_1302 ();
 sg13g2_decap_8 FILLER_18_1309 ();
 sg13g2_decap_8 FILLER_18_1316 ();
 sg13g2_fill_2 FILLER_18_1323 ();
 sg13g2_fill_1 FILLER_18_1325 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_20 ();
 sg13g2_decap_8 FILLER_19_27 ();
 sg13g2_fill_2 FILLER_19_34 ();
 sg13g2_decap_4 FILLER_19_41 ();
 sg13g2_fill_2 FILLER_19_45 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_4 FILLER_19_77 ();
 sg13g2_fill_1 FILLER_19_81 ();
 sg13g2_decap_8 FILLER_19_87 ();
 sg13g2_decap_8 FILLER_19_94 ();
 sg13g2_decap_8 FILLER_19_101 ();
 sg13g2_decap_8 FILLER_19_108 ();
 sg13g2_decap_8 FILLER_19_115 ();
 sg13g2_decap_8 FILLER_19_122 ();
 sg13g2_decap_8 FILLER_19_129 ();
 sg13g2_decap_8 FILLER_19_136 ();
 sg13g2_decap_8 FILLER_19_143 ();
 sg13g2_fill_2 FILLER_19_150 ();
 sg13g2_decap_4 FILLER_19_170 ();
 sg13g2_decap_8 FILLER_19_184 ();
 sg13g2_decap_8 FILLER_19_191 ();
 sg13g2_decap_4 FILLER_19_198 ();
 sg13g2_fill_2 FILLER_19_202 ();
 sg13g2_decap_8 FILLER_19_209 ();
 sg13g2_decap_8 FILLER_19_216 ();
 sg13g2_fill_2 FILLER_19_223 ();
 sg13g2_fill_1 FILLER_19_225 ();
 sg13g2_decap_4 FILLER_19_252 ();
 sg13g2_fill_2 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_299 ();
 sg13g2_decap_8 FILLER_19_306 ();
 sg13g2_decap_8 FILLER_19_313 ();
 sg13g2_decap_8 FILLER_19_320 ();
 sg13g2_fill_1 FILLER_19_327 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_decap_8 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_fill_2 FILLER_19_354 ();
 sg13g2_decap_4 FILLER_19_360 ();
 sg13g2_fill_1 FILLER_19_364 ();
 sg13g2_fill_1 FILLER_19_369 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_fill_2 FILLER_19_392 ();
 sg13g2_fill_1 FILLER_19_394 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_decap_8 FILLER_19_415 ();
 sg13g2_decap_8 FILLER_19_422 ();
 sg13g2_decap_8 FILLER_19_429 ();
 sg13g2_fill_2 FILLER_19_436 ();
 sg13g2_fill_1 FILLER_19_442 ();
 sg13g2_decap_8 FILLER_19_452 ();
 sg13g2_fill_2 FILLER_19_459 ();
 sg13g2_fill_2 FILLER_19_465 ();
 sg13g2_decap_8 FILLER_19_477 ();
 sg13g2_decap_8 FILLER_19_484 ();
 sg13g2_decap_8 FILLER_19_491 ();
 sg13g2_decap_8 FILLER_19_498 ();
 sg13g2_decap_8 FILLER_19_505 ();
 sg13g2_decap_4 FILLER_19_512 ();
 sg13g2_fill_1 FILLER_19_516 ();
 sg13g2_decap_8 FILLER_19_527 ();
 sg13g2_fill_2 FILLER_19_534 ();
 sg13g2_fill_1 FILLER_19_536 ();
 sg13g2_decap_8 FILLER_19_547 ();
 sg13g2_decap_8 FILLER_19_554 ();
 sg13g2_decap_8 FILLER_19_561 ();
 sg13g2_decap_8 FILLER_19_568 ();
 sg13g2_decap_8 FILLER_19_575 ();
 sg13g2_decap_8 FILLER_19_582 ();
 sg13g2_fill_1 FILLER_19_589 ();
 sg13g2_decap_8 FILLER_19_606 ();
 sg13g2_decap_8 FILLER_19_613 ();
 sg13g2_decap_8 FILLER_19_620 ();
 sg13g2_decap_4 FILLER_19_627 ();
 sg13g2_decap_8 FILLER_19_652 ();
 sg13g2_decap_8 FILLER_19_680 ();
 sg13g2_decap_4 FILLER_19_687 ();
 sg13g2_fill_1 FILLER_19_691 ();
 sg13g2_decap_8 FILLER_19_703 ();
 sg13g2_decap_8 FILLER_19_710 ();
 sg13g2_decap_8 FILLER_19_717 ();
 sg13g2_decap_8 FILLER_19_724 ();
 sg13g2_decap_8 FILLER_19_731 ();
 sg13g2_decap_8 FILLER_19_738 ();
 sg13g2_decap_8 FILLER_19_745 ();
 sg13g2_decap_4 FILLER_19_752 ();
 sg13g2_fill_2 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_762 ();
 sg13g2_decap_8 FILLER_19_769 ();
 sg13g2_decap_8 FILLER_19_776 ();
 sg13g2_decap_8 FILLER_19_783 ();
 sg13g2_decap_8 FILLER_19_790 ();
 sg13g2_decap_8 FILLER_19_797 ();
 sg13g2_decap_8 FILLER_19_804 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_4 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_877 ();
 sg13g2_decap_8 FILLER_19_884 ();
 sg13g2_decap_8 FILLER_19_891 ();
 sg13g2_decap_8 FILLER_19_898 ();
 sg13g2_decap_8 FILLER_19_905 ();
 sg13g2_decap_8 FILLER_19_912 ();
 sg13g2_decap_8 FILLER_19_919 ();
 sg13g2_decap_8 FILLER_19_926 ();
 sg13g2_fill_2 FILLER_19_933 ();
 sg13g2_fill_1 FILLER_19_935 ();
 sg13g2_decap_8 FILLER_19_940 ();
 sg13g2_fill_2 FILLER_19_947 ();
 sg13g2_decap_4 FILLER_19_958 ();
 sg13g2_fill_2 FILLER_19_962 ();
 sg13g2_decap_8 FILLER_19_983 ();
 sg13g2_decap_8 FILLER_19_990 ();
 sg13g2_fill_2 FILLER_19_997 ();
 sg13g2_fill_2 FILLER_19_1003 ();
 sg13g2_fill_1 FILLER_19_1005 ();
 sg13g2_fill_1 FILLER_19_1010 ();
 sg13g2_fill_1 FILLER_19_1015 ();
 sg13g2_fill_1 FILLER_19_1021 ();
 sg13g2_decap_8 FILLER_19_1030 ();
 sg13g2_fill_2 FILLER_19_1037 ();
 sg13g2_decap_8 FILLER_19_1048 ();
 sg13g2_decap_8 FILLER_19_1055 ();
 sg13g2_fill_2 FILLER_19_1062 ();
 sg13g2_decap_4 FILLER_19_1068 ();
 sg13g2_fill_1 FILLER_19_1077 ();
 sg13g2_fill_2 FILLER_19_1083 ();
 sg13g2_fill_1 FILLER_19_1085 ();
 sg13g2_decap_4 FILLER_19_1099 ();
 sg13g2_fill_2 FILLER_19_1113 ();
 sg13g2_fill_1 FILLER_19_1119 ();
 sg13g2_fill_2 FILLER_19_1128 ();
 sg13g2_fill_1 FILLER_19_1130 ();
 sg13g2_fill_2 FILLER_19_1137 ();
 sg13g2_decap_8 FILLER_19_1143 ();
 sg13g2_decap_4 FILLER_19_1159 ();
 sg13g2_fill_1 FILLER_19_1167 ();
 sg13g2_decap_8 FILLER_19_1172 ();
 sg13g2_decap_4 FILLER_19_1184 ();
 sg13g2_fill_1 FILLER_19_1188 ();
 sg13g2_fill_1 FILLER_19_1198 ();
 sg13g2_decap_4 FILLER_19_1203 ();
 sg13g2_fill_2 FILLER_19_1207 ();
 sg13g2_decap_8 FILLER_19_1213 ();
 sg13g2_fill_1 FILLER_19_1220 ();
 sg13g2_fill_2 FILLER_19_1234 ();
 sg13g2_decap_4 FILLER_19_1241 ();
 sg13g2_fill_1 FILLER_19_1245 ();
 sg13g2_decap_4 FILLER_19_1252 ();
 sg13g2_decap_8 FILLER_19_1265 ();
 sg13g2_decap_8 FILLER_19_1272 ();
 sg13g2_fill_2 FILLER_19_1279 ();
 sg13g2_decap_8 FILLER_19_1285 ();
 sg13g2_decap_8 FILLER_19_1292 ();
 sg13g2_decap_8 FILLER_19_1299 ();
 sg13g2_decap_8 FILLER_19_1306 ();
 sg13g2_decap_8 FILLER_19_1313 ();
 sg13g2_decap_4 FILLER_19_1320 ();
 sg13g2_fill_2 FILLER_19_1324 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_21 ();
 sg13g2_fill_1 FILLER_20_25 ();
 sg13g2_decap_8 FILLER_20_41 ();
 sg13g2_fill_2 FILLER_20_48 ();
 sg13g2_fill_2 FILLER_20_71 ();
 sg13g2_fill_2 FILLER_20_77 ();
 sg13g2_fill_1 FILLER_20_79 ();
 sg13g2_decap_8 FILLER_20_95 ();
 sg13g2_decap_8 FILLER_20_102 ();
 sg13g2_decap_4 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_120 ();
 sg13g2_decap_8 FILLER_20_145 ();
 sg13g2_decap_8 FILLER_20_159 ();
 sg13g2_fill_2 FILLER_20_172 ();
 sg13g2_fill_1 FILLER_20_174 ();
 sg13g2_fill_2 FILLER_20_180 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_fill_2 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_decap_4 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_265 ();
 sg13g2_decap_8 FILLER_20_272 ();
 sg13g2_decap_4 FILLER_20_279 ();
 sg13g2_decap_8 FILLER_20_295 ();
 sg13g2_decap_8 FILLER_20_302 ();
 sg13g2_decap_8 FILLER_20_309 ();
 sg13g2_decap_4 FILLER_20_316 ();
 sg13g2_fill_1 FILLER_20_320 ();
 sg13g2_decap_4 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_decap_4 FILLER_20_379 ();
 sg13g2_fill_2 FILLER_20_383 ();
 sg13g2_decap_4 FILLER_20_393 ();
 sg13g2_fill_2 FILLER_20_434 ();
 sg13g2_fill_1 FILLER_20_436 ();
 sg13g2_fill_2 FILLER_20_463 ();
 sg13g2_decap_8 FILLER_20_491 ();
 sg13g2_decap_8 FILLER_20_498 ();
 sg13g2_decap_8 FILLER_20_505 ();
 sg13g2_decap_8 FILLER_20_516 ();
 sg13g2_decap_8 FILLER_20_523 ();
 sg13g2_decap_8 FILLER_20_530 ();
 sg13g2_decap_8 FILLER_20_537 ();
 sg13g2_decap_8 FILLER_20_544 ();
 sg13g2_decap_8 FILLER_20_551 ();
 sg13g2_decap_8 FILLER_20_558 ();
 sg13g2_decap_8 FILLER_20_565 ();
 sg13g2_decap_8 FILLER_20_572 ();
 sg13g2_decap_8 FILLER_20_579 ();
 sg13g2_decap_8 FILLER_20_586 ();
 sg13g2_decap_8 FILLER_20_593 ();
 sg13g2_decap_8 FILLER_20_600 ();
 sg13g2_decap_8 FILLER_20_607 ();
 sg13g2_decap_8 FILLER_20_614 ();
 sg13g2_decap_8 FILLER_20_621 ();
 sg13g2_decap_8 FILLER_20_628 ();
 sg13g2_decap_8 FILLER_20_635 ();
 sg13g2_decap_8 FILLER_20_642 ();
 sg13g2_decap_8 FILLER_20_649 ();
 sg13g2_decap_8 FILLER_20_656 ();
 sg13g2_decap_8 FILLER_20_663 ();
 sg13g2_decap_8 FILLER_20_670 ();
 sg13g2_decap_8 FILLER_20_677 ();
 sg13g2_decap_8 FILLER_20_684 ();
 sg13g2_decap_8 FILLER_20_691 ();
 sg13g2_decap_8 FILLER_20_698 ();
 sg13g2_decap_8 FILLER_20_705 ();
 sg13g2_decap_8 FILLER_20_712 ();
 sg13g2_decap_8 FILLER_20_719 ();
 sg13g2_decap_8 FILLER_20_726 ();
 sg13g2_decap_8 FILLER_20_733 ();
 sg13g2_decap_4 FILLER_20_740 ();
 sg13g2_fill_1 FILLER_20_744 ();
 sg13g2_decap_8 FILLER_20_757 ();
 sg13g2_decap_8 FILLER_20_764 ();
 sg13g2_decap_4 FILLER_20_771 ();
 sg13g2_fill_2 FILLER_20_775 ();
 sg13g2_decap_8 FILLER_20_793 ();
 sg13g2_decap_8 FILLER_20_800 ();
 sg13g2_decap_4 FILLER_20_807 ();
 sg13g2_fill_1 FILLER_20_811 ();
 sg13g2_decap_8 FILLER_20_842 ();
 sg13g2_decap_8 FILLER_20_849 ();
 sg13g2_fill_2 FILLER_20_856 ();
 sg13g2_decap_8 FILLER_20_862 ();
 sg13g2_decap_8 FILLER_20_869 ();
 sg13g2_decap_8 FILLER_20_876 ();
 sg13g2_decap_8 FILLER_20_883 ();
 sg13g2_fill_2 FILLER_20_890 ();
 sg13g2_decap_4 FILLER_20_896 ();
 sg13g2_decap_8 FILLER_20_904 ();
 sg13g2_fill_2 FILLER_20_911 ();
 sg13g2_fill_1 FILLER_20_913 ();
 sg13g2_decap_4 FILLER_20_923 ();
 sg13g2_fill_1 FILLER_20_927 ();
 sg13g2_decap_4 FILLER_20_933 ();
 sg13g2_decap_8 FILLER_20_945 ();
 sg13g2_decap_8 FILLER_20_952 ();
 sg13g2_fill_2 FILLER_20_959 ();
 sg13g2_fill_1 FILLER_20_961 ();
 sg13g2_fill_2 FILLER_20_971 ();
 sg13g2_decap_4 FILLER_20_977 ();
 sg13g2_fill_2 FILLER_20_981 ();
 sg13g2_decap_8 FILLER_20_989 ();
 sg13g2_decap_8 FILLER_20_996 ();
 sg13g2_fill_2 FILLER_20_1007 ();
 sg13g2_fill_1 FILLER_20_1009 ();
 sg13g2_decap_4 FILLER_20_1015 ();
 sg13g2_fill_1 FILLER_20_1019 ();
 sg13g2_decap_4 FILLER_20_1038 ();
 sg13g2_decap_8 FILLER_20_1046 ();
 sg13g2_decap_4 FILLER_20_1053 ();
 sg13g2_decap_8 FILLER_20_1062 ();
 sg13g2_fill_1 FILLER_20_1076 ();
 sg13g2_decap_4 FILLER_20_1091 ();
 sg13g2_fill_1 FILLER_20_1095 ();
 sg13g2_fill_2 FILLER_20_1101 ();
 sg13g2_fill_1 FILLER_20_1103 ();
 sg13g2_decap_4 FILLER_20_1113 ();
 sg13g2_fill_1 FILLER_20_1117 ();
 sg13g2_decap_4 FILLER_20_1123 ();
 sg13g2_fill_1 FILLER_20_1127 ();
 sg13g2_fill_2 FILLER_20_1133 ();
 sg13g2_decap_8 FILLER_20_1140 ();
 sg13g2_decap_8 FILLER_20_1147 ();
 sg13g2_fill_1 FILLER_20_1162 ();
 sg13g2_fill_2 FILLER_20_1171 ();
 sg13g2_fill_1 FILLER_20_1178 ();
 sg13g2_fill_2 FILLER_20_1183 ();
 sg13g2_decap_4 FILLER_20_1190 ();
 sg13g2_fill_1 FILLER_20_1194 ();
 sg13g2_decap_8 FILLER_20_1200 ();
 sg13g2_decap_8 FILLER_20_1207 ();
 sg13g2_fill_2 FILLER_20_1214 ();
 sg13g2_fill_1 FILLER_20_1228 ();
 sg13g2_decap_8 FILLER_20_1238 ();
 sg13g2_decap_8 FILLER_20_1245 ();
 sg13g2_decap_4 FILLER_20_1252 ();
 sg13g2_fill_2 FILLER_20_1256 ();
 sg13g2_fill_1 FILLER_20_1262 ();
 sg13g2_fill_2 FILLER_20_1267 ();
 sg13g2_decap_8 FILLER_20_1273 ();
 sg13g2_decap_8 FILLER_20_1280 ();
 sg13g2_decap_8 FILLER_20_1287 ();
 sg13g2_decap_8 FILLER_20_1294 ();
 sg13g2_decap_8 FILLER_20_1301 ();
 sg13g2_decap_8 FILLER_20_1308 ();
 sg13g2_decap_8 FILLER_20_1315 ();
 sg13g2_decap_4 FILLER_20_1322 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_14 ();
 sg13g2_decap_4 FILLER_21_27 ();
 sg13g2_decap_8 FILLER_21_46 ();
 sg13g2_decap_4 FILLER_21_53 ();
 sg13g2_fill_2 FILLER_21_57 ();
 sg13g2_decap_8 FILLER_21_68 ();
 sg13g2_decap_8 FILLER_21_75 ();
 sg13g2_decap_8 FILLER_21_82 ();
 sg13g2_fill_1 FILLER_21_89 ();
 sg13g2_decap_8 FILLER_21_94 ();
 sg13g2_fill_1 FILLER_21_101 ();
 sg13g2_decap_8 FILLER_21_109 ();
 sg13g2_decap_4 FILLER_21_116 ();
 sg13g2_fill_2 FILLER_21_120 ();
 sg13g2_decap_4 FILLER_21_145 ();
 sg13g2_decap_8 FILLER_21_158 ();
 sg13g2_decap_8 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_172 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_fill_2 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_214 ();
 sg13g2_decap_8 FILLER_21_221 ();
 sg13g2_decap_8 FILLER_21_228 ();
 sg13g2_decap_8 FILLER_21_235 ();
 sg13g2_decap_8 FILLER_21_242 ();
 sg13g2_decap_4 FILLER_21_249 ();
 sg13g2_fill_2 FILLER_21_253 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_fill_1 FILLER_21_266 ();
 sg13g2_decap_4 FILLER_21_292 ();
 sg13g2_decap_4 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_327 ();
 sg13g2_decap_8 FILLER_21_334 ();
 sg13g2_decap_8 FILLER_21_341 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_fill_1 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_21_409 ();
 sg13g2_decap_8 FILLER_21_416 ();
 sg13g2_decap_8 FILLER_21_423 ();
 sg13g2_decap_8 FILLER_21_430 ();
 sg13g2_decap_8 FILLER_21_437 ();
 sg13g2_decap_8 FILLER_21_444 ();
 sg13g2_decap_8 FILLER_21_451 ();
 sg13g2_decap_8 FILLER_21_458 ();
 sg13g2_decap_4 FILLER_21_465 ();
 sg13g2_fill_2 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_475 ();
 sg13g2_decap_4 FILLER_21_482 ();
 sg13g2_fill_2 FILLER_21_507 ();
 sg13g2_decap_8 FILLER_21_535 ();
 sg13g2_decap_8 FILLER_21_542 ();
 sg13g2_decap_8 FILLER_21_549 ();
 sg13g2_decap_4 FILLER_21_577 ();
 sg13g2_decap_4 FILLER_21_602 ();
 sg13g2_fill_2 FILLER_21_606 ();
 sg13g2_decap_8 FILLER_21_645 ();
 sg13g2_decap_4 FILLER_21_652 ();
 sg13g2_fill_1 FILLER_21_656 ();
 sg13g2_fill_1 FILLER_21_663 ();
 sg13g2_decap_8 FILLER_21_668 ();
 sg13g2_decap_8 FILLER_21_675 ();
 sg13g2_decap_8 FILLER_21_682 ();
 sg13g2_decap_4 FILLER_21_689 ();
 sg13g2_fill_2 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_699 ();
 sg13g2_decap_8 FILLER_21_706 ();
 sg13g2_decap_8 FILLER_21_713 ();
 sg13g2_decap_8 FILLER_21_720 ();
 sg13g2_decap_8 FILLER_21_727 ();
 sg13g2_fill_2 FILLER_21_734 ();
 sg13g2_fill_1 FILLER_21_736 ();
 sg13g2_fill_1 FILLER_21_771 ();
 sg13g2_decap_8 FILLER_21_802 ();
 sg13g2_decap_8 FILLER_21_809 ();
 sg13g2_fill_2 FILLER_21_816 ();
 sg13g2_fill_1 FILLER_21_818 ();
 sg13g2_decap_8 FILLER_21_827 ();
 sg13g2_decap_8 FILLER_21_834 ();
 sg13g2_decap_8 FILLER_21_841 ();
 sg13g2_decap_8 FILLER_21_848 ();
 sg13g2_decap_8 FILLER_21_855 ();
 sg13g2_decap_8 FILLER_21_862 ();
 sg13g2_decap_8 FILLER_21_869 ();
 sg13g2_decap_8 FILLER_21_876 ();
 sg13g2_decap_8 FILLER_21_883 ();
 sg13g2_decap_8 FILLER_21_890 ();
 sg13g2_decap_8 FILLER_21_897 ();
 sg13g2_decap_8 FILLER_21_904 ();
 sg13g2_decap_4 FILLER_21_911 ();
 sg13g2_decap_4 FILLER_21_924 ();
 sg13g2_fill_2 FILLER_21_933 ();
 sg13g2_fill_2 FILLER_21_940 ();
 sg13g2_fill_1 FILLER_21_942 ();
 sg13g2_decap_8 FILLER_21_958 ();
 sg13g2_fill_2 FILLER_21_965 ();
 sg13g2_fill_1 FILLER_21_967 ();
 sg13g2_decap_8 FILLER_21_973 ();
 sg13g2_fill_2 FILLER_21_980 ();
 sg13g2_decap_4 FILLER_21_991 ();
 sg13g2_decap_4 FILLER_21_1000 ();
 sg13g2_decap_8 FILLER_21_1008 ();
 sg13g2_decap_8 FILLER_21_1015 ();
 sg13g2_decap_8 FILLER_21_1027 ();
 sg13g2_decap_8 FILLER_21_1034 ();
 sg13g2_decap_8 FILLER_21_1041 ();
 sg13g2_decap_8 FILLER_21_1048 ();
 sg13g2_decap_4 FILLER_21_1055 ();
 sg13g2_fill_2 FILLER_21_1064 ();
 sg13g2_decap_8 FILLER_21_1071 ();
 sg13g2_decap_4 FILLER_21_1078 ();
 sg13g2_decap_8 FILLER_21_1086 ();
 sg13g2_decap_8 FILLER_21_1101 ();
 sg13g2_decap_8 FILLER_21_1108 ();
 sg13g2_decap_8 FILLER_21_1115 ();
 sg13g2_fill_1 FILLER_21_1122 ();
 sg13g2_decap_8 FILLER_21_1127 ();
 sg13g2_fill_2 FILLER_21_1134 ();
 sg13g2_decap_8 FILLER_21_1140 ();
 sg13g2_decap_4 FILLER_21_1147 ();
 sg13g2_fill_1 FILLER_21_1151 ();
 sg13g2_fill_2 FILLER_21_1163 ();
 sg13g2_fill_1 FILLER_21_1165 ();
 sg13g2_fill_2 FILLER_21_1171 ();
 sg13g2_fill_1 FILLER_21_1186 ();
 sg13g2_decap_4 FILLER_21_1191 ();
 sg13g2_decap_4 FILLER_21_1204 ();
 sg13g2_fill_2 FILLER_21_1208 ();
 sg13g2_fill_2 FILLER_21_1233 ();
 sg13g2_decap_8 FILLER_21_1239 ();
 sg13g2_decap_8 FILLER_21_1246 ();
 sg13g2_fill_1 FILLER_21_1253 ();
 sg13g2_fill_2 FILLER_21_1261 ();
 sg13g2_fill_1 FILLER_21_1263 ();
 sg13g2_decap_8 FILLER_21_1268 ();
 sg13g2_decap_8 FILLER_21_1275 ();
 sg13g2_decap_8 FILLER_21_1282 ();
 sg13g2_decap_8 FILLER_21_1289 ();
 sg13g2_decap_8 FILLER_21_1296 ();
 sg13g2_decap_8 FILLER_21_1303 ();
 sg13g2_decap_8 FILLER_21_1310 ();
 sg13g2_decap_8 FILLER_21_1317 ();
 sg13g2_fill_2 FILLER_21_1324 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_4 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_4 FILLER_22_49 ();
 sg13g2_fill_1 FILLER_22_53 ();
 sg13g2_fill_2 FILLER_22_69 ();
 sg13g2_decap_4 FILLER_22_77 ();
 sg13g2_fill_1 FILLER_22_81 ();
 sg13g2_fill_2 FILLER_22_86 ();
 sg13g2_fill_1 FILLER_22_88 ();
 sg13g2_decap_8 FILLER_22_92 ();
 sg13g2_decap_8 FILLER_22_99 ();
 sg13g2_fill_1 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_114 ();
 sg13g2_decap_8 FILLER_22_121 ();
 sg13g2_decap_8 FILLER_22_128 ();
 sg13g2_fill_1 FILLER_22_135 ();
 sg13g2_decap_8 FILLER_22_141 ();
 sg13g2_decap_8 FILLER_22_148 ();
 sg13g2_decap_8 FILLER_22_155 ();
 sg13g2_decap_8 FILLER_22_162 ();
 sg13g2_decap_8 FILLER_22_169 ();
 sg13g2_decap_4 FILLER_22_176 ();
 sg13g2_decap_8 FILLER_22_185 ();
 sg13g2_decap_8 FILLER_22_192 ();
 sg13g2_decap_8 FILLER_22_199 ();
 sg13g2_decap_8 FILLER_22_206 ();
 sg13g2_decap_8 FILLER_22_213 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_fill_2 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_251 ();
 sg13g2_decap_8 FILLER_22_262 ();
 sg13g2_decap_8 FILLER_22_269 ();
 sg13g2_fill_2 FILLER_22_276 ();
 sg13g2_decap_8 FILLER_22_283 ();
 sg13g2_fill_2 FILLER_22_290 ();
 sg13g2_decap_8 FILLER_22_313 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_decap_8 FILLER_22_341 ();
 sg13g2_fill_2 FILLER_22_348 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_fill_2 FILLER_22_391 ();
 sg13g2_fill_1 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_22_414 ();
 sg13g2_decap_8 FILLER_22_421 ();
 sg13g2_decap_8 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_22_435 ();
 sg13g2_decap_8 FILLER_22_442 ();
 sg13g2_decap_8 FILLER_22_449 ();
 sg13g2_decap_8 FILLER_22_456 ();
 sg13g2_decap_8 FILLER_22_463 ();
 sg13g2_decap_8 FILLER_22_470 ();
 sg13g2_decap_8 FILLER_22_477 ();
 sg13g2_decap_8 FILLER_22_484 ();
 sg13g2_decap_8 FILLER_22_491 ();
 sg13g2_decap_8 FILLER_22_498 ();
 sg13g2_decap_8 FILLER_22_505 ();
 sg13g2_fill_1 FILLER_22_512 ();
 sg13g2_decap_4 FILLER_22_521 ();
 sg13g2_fill_1 FILLER_22_530 ();
 sg13g2_decap_8 FILLER_22_536 ();
 sg13g2_decap_8 FILLER_22_543 ();
 sg13g2_fill_2 FILLER_22_550 ();
 sg13g2_decap_8 FILLER_22_573 ();
 sg13g2_decap_8 FILLER_22_580 ();
 sg13g2_decap_8 FILLER_22_587 ();
 sg13g2_decap_8 FILLER_22_594 ();
 sg13g2_decap_8 FILLER_22_601 ();
 sg13g2_decap_8 FILLER_22_608 ();
 sg13g2_decap_8 FILLER_22_615 ();
 sg13g2_decap_8 FILLER_22_622 ();
 sg13g2_decap_8 FILLER_22_629 ();
 sg13g2_decap_8 FILLER_22_636 ();
 sg13g2_decap_8 FILLER_22_643 ();
 sg13g2_decap_8 FILLER_22_650 ();
 sg13g2_fill_2 FILLER_22_657 ();
 sg13g2_decap_8 FILLER_22_669 ();
 sg13g2_fill_1 FILLER_22_680 ();
 sg13g2_fill_1 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_694 ();
 sg13g2_fill_1 FILLER_22_701 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_fill_1 FILLER_22_777 ();
 sg13g2_decap_4 FILLER_22_783 ();
 sg13g2_fill_1 FILLER_22_787 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_fill_1 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_830 ();
 sg13g2_decap_8 FILLER_22_837 ();
 sg13g2_decap_8 FILLER_22_844 ();
 sg13g2_decap_8 FILLER_22_851 ();
 sg13g2_decap_8 FILLER_22_858 ();
 sg13g2_decap_8 FILLER_22_865 ();
 sg13g2_decap_8 FILLER_22_872 ();
 sg13g2_decap_8 FILLER_22_879 ();
 sg13g2_decap_8 FILLER_22_886 ();
 sg13g2_fill_2 FILLER_22_893 ();
 sg13g2_fill_1 FILLER_22_895 ();
 sg13g2_decap_4 FILLER_22_901 ();
 sg13g2_fill_1 FILLER_22_905 ();
 sg13g2_decap_8 FILLER_22_929 ();
 sg13g2_fill_1 FILLER_22_936 ();
 sg13g2_fill_2 FILLER_22_942 ();
 sg13g2_fill_1 FILLER_22_961 ();
 sg13g2_fill_2 FILLER_22_967 ();
 sg13g2_fill_1 FILLER_22_969 ();
 sg13g2_fill_2 FILLER_22_982 ();
 sg13g2_fill_1 FILLER_22_984 ();
 sg13g2_fill_2 FILLER_22_1005 ();
 sg13g2_decap_4 FILLER_22_1012 ();
 sg13g2_fill_2 FILLER_22_1016 ();
 sg13g2_decap_8 FILLER_22_1023 ();
 sg13g2_decap_8 FILLER_22_1030 ();
 sg13g2_decap_8 FILLER_22_1037 ();
 sg13g2_decap_8 FILLER_22_1044 ();
 sg13g2_decap_4 FILLER_22_1072 ();
 sg13g2_fill_1 FILLER_22_1076 ();
 sg13g2_decap_4 FILLER_22_1097 ();
 sg13g2_fill_2 FILLER_22_1111 ();
 sg13g2_fill_1 FILLER_22_1121 ();
 sg13g2_decap_8 FILLER_22_1129 ();
 sg13g2_decap_4 FILLER_22_1136 ();
 sg13g2_decap_8 FILLER_22_1150 ();
 sg13g2_decap_8 FILLER_22_1157 ();
 sg13g2_decap_8 FILLER_22_1164 ();
 sg13g2_decap_8 FILLER_22_1171 ();
 sg13g2_fill_2 FILLER_22_1178 ();
 sg13g2_fill_1 FILLER_22_1180 ();
 sg13g2_decap_8 FILLER_22_1186 ();
 sg13g2_decap_4 FILLER_22_1193 ();
 sg13g2_fill_2 FILLER_22_1197 ();
 sg13g2_decap_8 FILLER_22_1204 ();
 sg13g2_decap_8 FILLER_22_1211 ();
 sg13g2_decap_8 FILLER_22_1222 ();
 sg13g2_decap_4 FILLER_22_1229 ();
 sg13g2_fill_1 FILLER_22_1233 ();
 sg13g2_decap_4 FILLER_22_1244 ();
 sg13g2_fill_1 FILLER_22_1248 ();
 sg13g2_decap_4 FILLER_22_1259 ();
 sg13g2_decap_4 FILLER_22_1267 ();
 sg13g2_fill_2 FILLER_22_1276 ();
 sg13g2_fill_1 FILLER_22_1278 ();
 sg13g2_decap_8 FILLER_22_1284 ();
 sg13g2_decap_8 FILLER_22_1291 ();
 sg13g2_decap_8 FILLER_22_1298 ();
 sg13g2_decap_8 FILLER_22_1305 ();
 sg13g2_decap_8 FILLER_22_1312 ();
 sg13g2_decap_8 FILLER_22_1319 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_4 FILLER_23_56 ();
 sg13g2_fill_1 FILLER_23_60 ();
 sg13g2_fill_2 FILLER_23_65 ();
 sg13g2_decap_8 FILLER_23_71 ();
 sg13g2_decap_8 FILLER_23_78 ();
 sg13g2_fill_2 FILLER_23_85 ();
 sg13g2_fill_1 FILLER_23_95 ();
 sg13g2_decap_8 FILLER_23_102 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_decap_4 FILLER_23_116 ();
 sg13g2_fill_2 FILLER_23_120 ();
 sg13g2_decap_8 FILLER_23_129 ();
 sg13g2_fill_1 FILLER_23_136 ();
 sg13g2_decap_8 FILLER_23_142 ();
 sg13g2_decap_8 FILLER_23_149 ();
 sg13g2_decap_8 FILLER_23_156 ();
 sg13g2_decap_4 FILLER_23_163 ();
 sg13g2_fill_2 FILLER_23_167 ();
 sg13g2_decap_8 FILLER_23_174 ();
 sg13g2_decap_8 FILLER_23_181 ();
 sg13g2_decap_8 FILLER_23_188 ();
 sg13g2_decap_8 FILLER_23_195 ();
 sg13g2_decap_8 FILLER_23_202 ();
 sg13g2_decap_8 FILLER_23_209 ();
 sg13g2_decap_8 FILLER_23_216 ();
 sg13g2_decap_8 FILLER_23_223 ();
 sg13g2_decap_8 FILLER_23_230 ();
 sg13g2_decap_8 FILLER_23_237 ();
 sg13g2_decap_8 FILLER_23_244 ();
 sg13g2_decap_8 FILLER_23_255 ();
 sg13g2_decap_8 FILLER_23_262 ();
 sg13g2_fill_1 FILLER_23_269 ();
 sg13g2_decap_8 FILLER_23_296 ();
 sg13g2_decap_8 FILLER_23_303 ();
 sg13g2_decap_8 FILLER_23_310 ();
 sg13g2_decap_8 FILLER_23_317 ();
 sg13g2_decap_8 FILLER_23_324 ();
 sg13g2_fill_2 FILLER_23_331 ();
 sg13g2_decap_8 FILLER_23_346 ();
 sg13g2_fill_2 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_decap_4 FILLER_23_390 ();
 sg13g2_fill_1 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_411 ();
 sg13g2_fill_2 FILLER_23_418 ();
 sg13g2_decap_8 FILLER_23_428 ();
 sg13g2_decap_8 FILLER_23_435 ();
 sg13g2_decap_8 FILLER_23_442 ();
 sg13g2_decap_8 FILLER_23_449 ();
 sg13g2_decap_8 FILLER_23_456 ();
 sg13g2_decap_8 FILLER_23_463 ();
 sg13g2_fill_2 FILLER_23_470 ();
 sg13g2_fill_1 FILLER_23_472 ();
 sg13g2_decap_4 FILLER_23_477 ();
 sg13g2_fill_2 FILLER_23_481 ();
 sg13g2_decap_8 FILLER_23_487 ();
 sg13g2_decap_8 FILLER_23_494 ();
 sg13g2_decap_8 FILLER_23_501 ();
 sg13g2_decap_4 FILLER_23_508 ();
 sg13g2_fill_2 FILLER_23_512 ();
 sg13g2_decap_8 FILLER_23_519 ();
 sg13g2_fill_1 FILLER_23_556 ();
 sg13g2_decap_8 FILLER_23_583 ();
 sg13g2_decap_8 FILLER_23_590 ();
 sg13g2_decap_8 FILLER_23_597 ();
 sg13g2_fill_1 FILLER_23_604 ();
 sg13g2_decap_8 FILLER_23_612 ();
 sg13g2_decap_8 FILLER_23_619 ();
 sg13g2_decap_8 FILLER_23_626 ();
 sg13g2_decap_8 FILLER_23_633 ();
 sg13g2_decap_4 FILLER_23_640 ();
 sg13g2_decap_8 FILLER_23_670 ();
 sg13g2_fill_2 FILLER_23_677 ();
 sg13g2_fill_1 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_fill_1 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_698 ();
 sg13g2_decap_4 FILLER_23_705 ();
 sg13g2_decap_8 FILLER_23_713 ();
 sg13g2_decap_8 FILLER_23_720 ();
 sg13g2_decap_8 FILLER_23_727 ();
 sg13g2_decap_8 FILLER_23_734 ();
 sg13g2_decap_8 FILLER_23_741 ();
 sg13g2_decap_8 FILLER_23_748 ();
 sg13g2_decap_8 FILLER_23_755 ();
 sg13g2_decap_8 FILLER_23_762 ();
 sg13g2_decap_4 FILLER_23_777 ();
 sg13g2_fill_1 FILLER_23_781 ();
 sg13g2_fill_1 FILLER_23_787 ();
 sg13g2_decap_8 FILLER_23_794 ();
 sg13g2_decap_8 FILLER_23_801 ();
 sg13g2_decap_8 FILLER_23_816 ();
 sg13g2_fill_1 FILLER_23_823 ();
 sg13g2_decap_8 FILLER_23_828 ();
 sg13g2_decap_8 FILLER_23_835 ();
 sg13g2_decap_8 FILLER_23_842 ();
 sg13g2_decap_8 FILLER_23_849 ();
 sg13g2_decap_8 FILLER_23_856 ();
 sg13g2_decap_8 FILLER_23_863 ();
 sg13g2_decap_8 FILLER_23_870 ();
 sg13g2_decap_8 FILLER_23_877 ();
 sg13g2_decap_8 FILLER_23_884 ();
 sg13g2_decap_4 FILLER_23_891 ();
 sg13g2_fill_2 FILLER_23_895 ();
 sg13g2_fill_1 FILLER_23_910 ();
 sg13g2_fill_2 FILLER_23_916 ();
 sg13g2_fill_1 FILLER_23_918 ();
 sg13g2_decap_8 FILLER_23_927 ();
 sg13g2_fill_1 FILLER_23_934 ();
 sg13g2_decap_4 FILLER_23_941 ();
 sg13g2_decap_8 FILLER_23_949 ();
 sg13g2_decap_8 FILLER_23_956 ();
 sg13g2_decap_8 FILLER_23_963 ();
 sg13g2_fill_2 FILLER_23_970 ();
 sg13g2_decap_8 FILLER_23_981 ();
 sg13g2_fill_2 FILLER_23_998 ();
 sg13g2_fill_2 FILLER_23_1005 ();
 sg13g2_fill_1 FILLER_23_1007 ();
 sg13g2_decap_8 FILLER_23_1013 ();
 sg13g2_decap_8 FILLER_23_1020 ();
 sg13g2_decap_8 FILLER_23_1027 ();
 sg13g2_fill_2 FILLER_23_1034 ();
 sg13g2_decap_4 FILLER_23_1040 ();
 sg13g2_fill_1 FILLER_23_1044 ();
 sg13g2_decap_4 FILLER_23_1049 ();
 sg13g2_fill_1 FILLER_23_1053 ();
 sg13g2_decap_8 FILLER_23_1070 ();
 sg13g2_decap_4 FILLER_23_1077 ();
 sg13g2_fill_1 FILLER_23_1081 ();
 sg13g2_decap_8 FILLER_23_1087 ();
 sg13g2_decap_4 FILLER_23_1094 ();
 sg13g2_fill_1 FILLER_23_1098 ();
 sg13g2_fill_1 FILLER_23_1118 ();
 sg13g2_fill_2 FILLER_23_1143 ();
 sg13g2_fill_1 FILLER_23_1145 ();
 sg13g2_decap_8 FILLER_23_1172 ();
 sg13g2_decap_8 FILLER_23_1179 ();
 sg13g2_decap_8 FILLER_23_1186 ();
 sg13g2_decap_8 FILLER_23_1193 ();
 sg13g2_decap_4 FILLER_23_1200 ();
 sg13g2_fill_2 FILLER_23_1204 ();
 sg13g2_decap_8 FILLER_23_1215 ();
 sg13g2_decap_4 FILLER_23_1231 ();
 sg13g2_fill_2 FILLER_23_1235 ();
 sg13g2_decap_4 FILLER_23_1245 ();
 sg13g2_fill_1 FILLER_23_1249 ();
 sg13g2_decap_4 FILLER_23_1255 ();
 sg13g2_decap_4 FILLER_23_1272 ();
 sg13g2_decap_8 FILLER_23_1280 ();
 sg13g2_fill_2 FILLER_23_1287 ();
 sg13g2_fill_1 FILLER_23_1289 ();
 sg13g2_decap_8 FILLER_23_1294 ();
 sg13g2_decap_8 FILLER_23_1301 ();
 sg13g2_decap_8 FILLER_23_1308 ();
 sg13g2_decap_8 FILLER_23_1315 ();
 sg13g2_decap_4 FILLER_23_1322 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_37 ();
 sg13g2_fill_1 FILLER_24_44 ();
 sg13g2_decap_8 FILLER_24_62 ();
 sg13g2_decap_8 FILLER_24_73 ();
 sg13g2_fill_2 FILLER_24_80 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_decap_4 FILLER_24_88 ();
 sg13g2_fill_1 FILLER_24_92 ();
 sg13g2_decap_4 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_114 ();
 sg13g2_fill_2 FILLER_24_128 ();
 sg13g2_fill_2 FILLER_24_134 ();
 sg13g2_decap_8 FILLER_24_145 ();
 sg13g2_fill_2 FILLER_24_152 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_4 FILLER_24_175 ();
 sg13g2_fill_2 FILLER_24_184 ();
 sg13g2_decap_8 FILLER_24_194 ();
 sg13g2_decap_8 FILLER_24_201 ();
 sg13g2_fill_2 FILLER_24_208 ();
 sg13g2_fill_1 FILLER_24_210 ();
 sg13g2_fill_2 FILLER_24_221 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_decap_4 FILLER_24_239 ();
 sg13g2_fill_1 FILLER_24_243 ();
 sg13g2_decap_8 FILLER_24_253 ();
 sg13g2_decap_8 FILLER_24_260 ();
 sg13g2_decap_4 FILLER_24_267 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_decap_8 FILLER_24_299 ();
 sg13g2_decap_8 FILLER_24_306 ();
 sg13g2_decap_8 FILLER_24_313 ();
 sg13g2_decap_8 FILLER_24_320 ();
 sg13g2_decap_8 FILLER_24_327 ();
 sg13g2_decap_8 FILLER_24_334 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_fill_2 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_372 ();
 sg13g2_decap_8 FILLER_24_379 ();
 sg13g2_decap_4 FILLER_24_386 ();
 sg13g2_fill_1 FILLER_24_390 ();
 sg13g2_fill_1 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_24_411 ();
 sg13g2_fill_2 FILLER_24_418 ();
 sg13g2_decap_8 FILLER_24_435 ();
 sg13g2_decap_8 FILLER_24_442 ();
 sg13g2_decap_8 FILLER_24_449 ();
 sg13g2_decap_8 FILLER_24_456 ();
 sg13g2_fill_1 FILLER_24_463 ();
 sg13g2_fill_2 FILLER_24_473 ();
 sg13g2_fill_1 FILLER_24_475 ();
 sg13g2_decap_4 FILLER_24_507 ();
 sg13g2_fill_1 FILLER_24_511 ();
 sg13g2_decap_8 FILLER_24_517 ();
 sg13g2_decap_8 FILLER_24_524 ();
 sg13g2_decap_4 FILLER_24_531 ();
 sg13g2_fill_1 FILLER_24_535 ();
 sg13g2_decap_8 FILLER_24_545 ();
 sg13g2_fill_2 FILLER_24_552 ();
 sg13g2_fill_2 FILLER_24_558 ();
 sg13g2_fill_1 FILLER_24_560 ();
 sg13g2_fill_2 FILLER_24_566 ();
 sg13g2_decap_8 FILLER_24_572 ();
 sg13g2_decap_8 FILLER_24_579 ();
 sg13g2_decap_8 FILLER_24_586 ();
 sg13g2_decap_4 FILLER_24_593 ();
 sg13g2_fill_2 FILLER_24_597 ();
 sg13g2_decap_8 FILLER_24_613 ();
 sg13g2_decap_4 FILLER_24_620 ();
 sg13g2_fill_2 FILLER_24_624 ();
 sg13g2_decap_8 FILLER_24_652 ();
 sg13g2_decap_4 FILLER_24_659 ();
 sg13g2_decap_4 FILLER_24_670 ();
 sg13g2_fill_1 FILLER_24_674 ();
 sg13g2_decap_8 FILLER_24_713 ();
 sg13g2_decap_8 FILLER_24_720 ();
 sg13g2_decap_8 FILLER_24_727 ();
 sg13g2_decap_8 FILLER_24_734 ();
 sg13g2_fill_1 FILLER_24_741 ();
 sg13g2_fill_2 FILLER_24_758 ();
 sg13g2_fill_2 FILLER_24_771 ();
 sg13g2_decap_8 FILLER_24_785 ();
 sg13g2_decap_8 FILLER_24_792 ();
 sg13g2_decap_8 FILLER_24_799 ();
 sg13g2_fill_2 FILLER_24_806 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_fill_2 FILLER_24_819 ();
 sg13g2_fill_1 FILLER_24_821 ();
 sg13g2_decap_8 FILLER_24_852 ();
 sg13g2_decap_8 FILLER_24_859 ();
 sg13g2_decap_8 FILLER_24_866 ();
 sg13g2_decap_8 FILLER_24_873 ();
 sg13g2_decap_8 FILLER_24_880 ();
 sg13g2_decap_8 FILLER_24_887 ();
 sg13g2_fill_2 FILLER_24_894 ();
 sg13g2_fill_1 FILLER_24_896 ();
 sg13g2_decap_4 FILLER_24_906 ();
 sg13g2_fill_1 FILLER_24_910 ();
 sg13g2_fill_2 FILLER_24_924 ();
 sg13g2_fill_1 FILLER_24_941 ();
 sg13g2_fill_2 FILLER_24_946 ();
 sg13g2_fill_1 FILLER_24_948 ();
 sg13g2_decap_8 FILLER_24_954 ();
 sg13g2_fill_2 FILLER_24_961 ();
 sg13g2_decap_8 FILLER_24_967 ();
 sg13g2_decap_8 FILLER_24_974 ();
 sg13g2_decap_4 FILLER_24_985 ();
 sg13g2_fill_1 FILLER_24_989 ();
 sg13g2_fill_2 FILLER_24_1005 ();
 sg13g2_fill_1 FILLER_24_1007 ();
 sg13g2_fill_2 FILLER_24_1013 ();
 sg13g2_fill_2 FILLER_24_1026 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_decap_8 FILLER_24_1037 ();
 sg13g2_decap_4 FILLER_24_1044 ();
 sg13g2_fill_2 FILLER_24_1048 ();
 sg13g2_decap_8 FILLER_24_1066 ();
 sg13g2_decap_4 FILLER_24_1073 ();
 sg13g2_fill_1 FILLER_24_1077 ();
 sg13g2_decap_4 FILLER_24_1095 ();
 sg13g2_fill_1 FILLER_24_1099 ();
 sg13g2_fill_1 FILLER_24_1110 ();
 sg13g2_decap_8 FILLER_24_1125 ();
 sg13g2_decap_8 FILLER_24_1142 ();
 sg13g2_fill_1 FILLER_24_1170 ();
 sg13g2_fill_1 FILLER_24_1176 ();
 sg13g2_fill_2 FILLER_24_1187 ();
 sg13g2_decap_8 FILLER_24_1200 ();
 sg13g2_decap_4 FILLER_24_1207 ();
 sg13g2_fill_2 FILLER_24_1211 ();
 sg13g2_fill_2 FILLER_24_1218 ();
 sg13g2_fill_2 FILLER_24_1229 ();
 sg13g2_fill_2 FILLER_24_1240 ();
 sg13g2_fill_2 FILLER_24_1247 ();
 sg13g2_fill_1 FILLER_24_1249 ();
 sg13g2_decap_4 FILLER_24_1256 ();
 sg13g2_fill_1 FILLER_24_1260 ();
 sg13g2_fill_1 FILLER_24_1271 ();
 sg13g2_decap_8 FILLER_24_1282 ();
 sg13g2_decap_8 FILLER_24_1289 ();
 sg13g2_decap_8 FILLER_24_1296 ();
 sg13g2_decap_8 FILLER_24_1303 ();
 sg13g2_decap_8 FILLER_24_1310 ();
 sg13g2_decap_8 FILLER_24_1317 ();
 sg13g2_fill_2 FILLER_24_1324 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_fill_2 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_23 ();
 sg13g2_decap_8 FILLER_25_34 ();
 sg13g2_decap_4 FILLER_25_41 ();
 sg13g2_fill_1 FILLER_25_49 ();
 sg13g2_fill_2 FILLER_25_55 ();
 sg13g2_fill_1 FILLER_25_62 ();
 sg13g2_decap_8 FILLER_25_68 ();
 sg13g2_decap_4 FILLER_25_75 ();
 sg13g2_fill_2 FILLER_25_79 ();
 sg13g2_decap_4 FILLER_25_86 ();
 sg13g2_fill_1 FILLER_25_90 ();
 sg13g2_decap_8 FILLER_25_96 ();
 sg13g2_fill_2 FILLER_25_103 ();
 sg13g2_fill_1 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_115 ();
 sg13g2_decap_4 FILLER_25_126 ();
 sg13g2_fill_2 FILLER_25_130 ();
 sg13g2_decap_8 FILLER_25_142 ();
 sg13g2_decap_4 FILLER_25_149 ();
 sg13g2_fill_2 FILLER_25_153 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_decap_8 FILLER_25_194 ();
 sg13g2_decap_8 FILLER_25_201 ();
 sg13g2_decap_8 FILLER_25_208 ();
 sg13g2_decap_8 FILLER_25_215 ();
 sg13g2_decap_4 FILLER_25_222 ();
 sg13g2_fill_1 FILLER_25_226 ();
 sg13g2_decap_8 FILLER_25_237 ();
 sg13g2_decap_4 FILLER_25_244 ();
 sg13g2_decap_8 FILLER_25_253 ();
 sg13g2_decap_8 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_267 ();
 sg13g2_fill_1 FILLER_25_269 ();
 sg13g2_fill_2 FILLER_25_280 ();
 sg13g2_fill_1 FILLER_25_282 ();
 sg13g2_decap_8 FILLER_25_288 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_324 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_8 FILLER_25_338 ();
 sg13g2_fill_2 FILLER_25_345 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_decap_4 FILLER_25_352 ();
 sg13g2_fill_1 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_fill_2 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_2 FILLER_25_408 ();
 sg13g2_fill_1 FILLER_25_410 ();
 sg13g2_fill_1 FILLER_25_424 ();
 sg13g2_decap_4 FILLER_25_430 ();
 sg13g2_fill_1 FILLER_25_434 ();
 sg13g2_fill_2 FILLER_25_443 ();
 sg13g2_fill_1 FILLER_25_492 ();
 sg13g2_decap_8 FILLER_25_498 ();
 sg13g2_decap_8 FILLER_25_505 ();
 sg13g2_decap_4 FILLER_25_512 ();
 sg13g2_fill_2 FILLER_25_516 ();
 sg13g2_decap_8 FILLER_25_529 ();
 sg13g2_decap_8 FILLER_25_536 ();
 sg13g2_decap_8 FILLER_25_543 ();
 sg13g2_decap_8 FILLER_25_550 ();
 sg13g2_decap_8 FILLER_25_557 ();
 sg13g2_fill_2 FILLER_25_564 ();
 sg13g2_decap_8 FILLER_25_587 ();
 sg13g2_decap_8 FILLER_25_594 ();
 sg13g2_decap_8 FILLER_25_601 ();
 sg13g2_decap_8 FILLER_25_608 ();
 sg13g2_decap_8 FILLER_25_615 ();
 sg13g2_decap_8 FILLER_25_622 ();
 sg13g2_fill_2 FILLER_25_629 ();
 sg13g2_fill_1 FILLER_25_631 ();
 sg13g2_decap_8 FILLER_25_636 ();
 sg13g2_decap_8 FILLER_25_643 ();
 sg13g2_fill_2 FILLER_25_650 ();
 sg13g2_decap_8 FILLER_25_663 ();
 sg13g2_decap_4 FILLER_25_670 ();
 sg13g2_decap_8 FILLER_25_683 ();
 sg13g2_decap_8 FILLER_25_690 ();
 sg13g2_decap_8 FILLER_25_697 ();
 sg13g2_decap_8 FILLER_25_704 ();
 sg13g2_decap_8 FILLER_25_711 ();
 sg13g2_decap_8 FILLER_25_718 ();
 sg13g2_decap_8 FILLER_25_725 ();
 sg13g2_decap_4 FILLER_25_766 ();
 sg13g2_decap_4 FILLER_25_796 ();
 sg13g2_decap_4 FILLER_25_805 ();
 sg13g2_fill_1 FILLER_25_835 ();
 sg13g2_decap_8 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_decap_8 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_25_868 ();
 sg13g2_decap_8 FILLER_25_875 ();
 sg13g2_decap_8 FILLER_25_882 ();
 sg13g2_decap_8 FILLER_25_889 ();
 sg13g2_fill_1 FILLER_25_896 ();
 sg13g2_fill_2 FILLER_25_902 ();
 sg13g2_fill_1 FILLER_25_904 ();
 sg13g2_decap_8 FILLER_25_910 ();
 sg13g2_fill_2 FILLER_25_921 ();
 sg13g2_fill_2 FILLER_25_931 ();
 sg13g2_fill_1 FILLER_25_933 ();
 sg13g2_decap_4 FILLER_25_943 ();
 sg13g2_fill_1 FILLER_25_947 ();
 sg13g2_decap_8 FILLER_25_961 ();
 sg13g2_decap_8 FILLER_25_973 ();
 sg13g2_fill_1 FILLER_25_980 ();
 sg13g2_fill_2 FILLER_25_991 ();
 sg13g2_fill_1 FILLER_25_993 ();
 sg13g2_fill_1 FILLER_25_998 ();
 sg13g2_decap_4 FILLER_25_1012 ();
 sg13g2_fill_2 FILLER_25_1016 ();
 sg13g2_fill_2 FILLER_25_1036 ();
 sg13g2_fill_1 FILLER_25_1042 ();
 sg13g2_decap_4 FILLER_25_1049 ();
 sg13g2_fill_1 FILLER_25_1053 ();
 sg13g2_fill_1 FILLER_25_1059 ();
 sg13g2_decap_8 FILLER_25_1072 ();
 sg13g2_decap_4 FILLER_25_1079 ();
 sg13g2_decap_4 FILLER_25_1091 ();
 sg13g2_decap_8 FILLER_25_1100 ();
 sg13g2_fill_2 FILLER_25_1107 ();
 sg13g2_fill_1 FILLER_25_1109 ();
 sg13g2_decap_8 FILLER_25_1115 ();
 sg13g2_decap_8 FILLER_25_1122 ();
 sg13g2_decap_4 FILLER_25_1129 ();
 sg13g2_decap_4 FILLER_25_1143 ();
 sg13g2_fill_1 FILLER_25_1147 ();
 sg13g2_decap_8 FILLER_25_1169 ();
 sg13g2_fill_1 FILLER_25_1176 ();
 sg13g2_fill_2 FILLER_25_1192 ();
 sg13g2_fill_1 FILLER_25_1194 ();
 sg13g2_decap_8 FILLER_25_1205 ();
 sg13g2_fill_2 FILLER_25_1212 ();
 sg13g2_decap_8 FILLER_25_1218 ();
 sg13g2_fill_1 FILLER_25_1225 ();
 sg13g2_decap_4 FILLER_25_1230 ();
 sg13g2_fill_1 FILLER_25_1234 ();
 sg13g2_fill_2 FILLER_25_1239 ();
 sg13g2_fill_1 FILLER_25_1241 ();
 sg13g2_fill_2 FILLER_25_1247 ();
 sg13g2_fill_2 FILLER_25_1259 ();
 sg13g2_decap_8 FILLER_25_1283 ();
 sg13g2_decap_8 FILLER_25_1290 ();
 sg13g2_decap_8 FILLER_25_1297 ();
 sg13g2_decap_8 FILLER_25_1304 ();
 sg13g2_decap_8 FILLER_25_1311 ();
 sg13g2_decap_8 FILLER_25_1318 ();
 sg13g2_fill_1 FILLER_25_1325 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_24 ();
 sg13g2_decap_8 FILLER_26_31 ();
 sg13g2_fill_2 FILLER_26_38 ();
 sg13g2_fill_1 FILLER_26_40 ();
 sg13g2_decap_4 FILLER_26_46 ();
 sg13g2_fill_1 FILLER_26_50 ();
 sg13g2_fill_2 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_58 ();
 sg13g2_fill_2 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_65 ();
 sg13g2_decap_4 FILLER_26_75 ();
 sg13g2_decap_4 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_100 ();
 sg13g2_decap_8 FILLER_26_107 ();
 sg13g2_decap_8 FILLER_26_114 ();
 sg13g2_fill_2 FILLER_26_127 ();
 sg13g2_fill_2 FILLER_26_134 ();
 sg13g2_fill_1 FILLER_26_136 ();
 sg13g2_decap_8 FILLER_26_143 ();
 sg13g2_decap_8 FILLER_26_150 ();
 sg13g2_decap_8 FILLER_26_157 ();
 sg13g2_decap_8 FILLER_26_164 ();
 sg13g2_fill_2 FILLER_26_171 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_decap_8 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_195 ();
 sg13g2_decap_8 FILLER_26_202 ();
 sg13g2_decap_8 FILLER_26_209 ();
 sg13g2_decap_4 FILLER_26_216 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_decap_8 FILLER_26_229 ();
 sg13g2_decap_8 FILLER_26_236 ();
 sg13g2_decap_8 FILLER_26_243 ();
 sg13g2_decap_8 FILLER_26_250 ();
 sg13g2_decap_8 FILLER_26_257 ();
 sg13g2_decap_8 FILLER_26_264 ();
 sg13g2_decap_8 FILLER_26_271 ();
 sg13g2_decap_8 FILLER_26_278 ();
 sg13g2_decap_8 FILLER_26_285 ();
 sg13g2_fill_2 FILLER_26_292 ();
 sg13g2_fill_1 FILLER_26_299 ();
 sg13g2_decap_4 FILLER_26_321 ();
 sg13g2_fill_2 FILLER_26_354 ();
 sg13g2_decap_4 FILLER_26_360 ();
 sg13g2_fill_2 FILLER_26_364 ();
 sg13g2_fill_2 FILLER_26_375 ();
 sg13g2_fill_1 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_fill_1 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_26_414 ();
 sg13g2_decap_8 FILLER_26_421 ();
 sg13g2_decap_8 FILLER_26_428 ();
 sg13g2_decap_8 FILLER_26_435 ();
 sg13g2_decap_8 FILLER_26_442 ();
 sg13g2_fill_2 FILLER_26_449 ();
 sg13g2_decap_8 FILLER_26_455 ();
 sg13g2_fill_2 FILLER_26_462 ();
 sg13g2_fill_1 FILLER_26_464 ();
 sg13g2_fill_1 FILLER_26_470 ();
 sg13g2_fill_1 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_482 ();
 sg13g2_fill_2 FILLER_26_489 ();
 sg13g2_fill_1 FILLER_26_491 ();
 sg13g2_fill_2 FILLER_26_496 ();
 sg13g2_fill_1 FILLER_26_498 ();
 sg13g2_decap_8 FILLER_26_525 ();
 sg13g2_decap_4 FILLER_26_532 ();
 sg13g2_fill_2 FILLER_26_536 ();
 sg13g2_decap_8 FILLER_26_543 ();
 sg13g2_decap_8 FILLER_26_550 ();
 sg13g2_decap_8 FILLER_26_557 ();
 sg13g2_decap_4 FILLER_26_564 ();
 sg13g2_fill_1 FILLER_26_568 ();
 sg13g2_fill_2 FILLER_26_573 ();
 sg13g2_fill_1 FILLER_26_575 ();
 sg13g2_fill_1 FILLER_26_602 ();
 sg13g2_decap_8 FILLER_26_610 ();
 sg13g2_decap_8 FILLER_26_617 ();
 sg13g2_decap_8 FILLER_26_624 ();
 sg13g2_decap_8 FILLER_26_631 ();
 sg13g2_decap_8 FILLER_26_638 ();
 sg13g2_decap_8 FILLER_26_645 ();
 sg13g2_fill_1 FILLER_26_652 ();
 sg13g2_fill_2 FILLER_26_669 ();
 sg13g2_fill_2 FILLER_26_680 ();
 sg13g2_decap_4 FILLER_26_686 ();
 sg13g2_fill_1 FILLER_26_690 ();
 sg13g2_decap_8 FILLER_26_697 ();
 sg13g2_decap_8 FILLER_26_704 ();
 sg13g2_decap_8 FILLER_26_711 ();
 sg13g2_decap_8 FILLER_26_718 ();
 sg13g2_decap_8 FILLER_26_725 ();
 sg13g2_decap_4 FILLER_26_732 ();
 sg13g2_fill_2 FILLER_26_736 ();
 sg13g2_decap_8 FILLER_26_742 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_756 ();
 sg13g2_decap_8 FILLER_26_763 ();
 sg13g2_decap_4 FILLER_26_770 ();
 sg13g2_fill_1 FILLER_26_774 ();
 sg13g2_fill_2 FILLER_26_779 ();
 sg13g2_fill_2 FILLER_26_789 ();
 sg13g2_decap_4 FILLER_26_795 ();
 sg13g2_fill_2 FILLER_26_799 ();
 sg13g2_decap_8 FILLER_26_805 ();
 sg13g2_fill_2 FILLER_26_812 ();
 sg13g2_decap_8 FILLER_26_843 ();
 sg13g2_decap_8 FILLER_26_850 ();
 sg13g2_decap_8 FILLER_26_857 ();
 sg13g2_decap_8 FILLER_26_864 ();
 sg13g2_decap_8 FILLER_26_871 ();
 sg13g2_decap_8 FILLER_26_878 ();
 sg13g2_decap_8 FILLER_26_885 ();
 sg13g2_decap_8 FILLER_26_892 ();
 sg13g2_fill_2 FILLER_26_899 ();
 sg13g2_fill_1 FILLER_26_901 ();
 sg13g2_fill_2 FILLER_26_921 ();
 sg13g2_decap_8 FILLER_26_927 ();
 sg13g2_decap_4 FILLER_26_934 ();
 sg13g2_fill_2 FILLER_26_955 ();
 sg13g2_fill_1 FILLER_26_957 ();
 sg13g2_decap_8 FILLER_26_977 ();
 sg13g2_decap_8 FILLER_26_984 ();
 sg13g2_fill_2 FILLER_26_991 ();
 sg13g2_decap_4 FILLER_26_997 ();
 sg13g2_fill_2 FILLER_26_1001 ();
 sg13g2_fill_1 FILLER_26_1008 ();
 sg13g2_fill_1 FILLER_26_1019 ();
 sg13g2_decap_8 FILLER_26_1025 ();
 sg13g2_decap_8 FILLER_26_1032 ();
 sg13g2_fill_1 FILLER_26_1039 ();
 sg13g2_decap_4 FILLER_26_1046 ();
 sg13g2_fill_2 FILLER_26_1050 ();
 sg13g2_decap_4 FILLER_26_1066 ();
 sg13g2_fill_1 FILLER_26_1070 ();
 sg13g2_decap_8 FILLER_26_1087 ();
 sg13g2_decap_8 FILLER_26_1094 ();
 sg13g2_decap_8 FILLER_26_1101 ();
 sg13g2_decap_8 FILLER_26_1108 ();
 sg13g2_decap_8 FILLER_26_1115 ();
 sg13g2_decap_8 FILLER_26_1122 ();
 sg13g2_decap_4 FILLER_26_1129 ();
 sg13g2_fill_1 FILLER_26_1133 ();
 sg13g2_decap_4 FILLER_26_1139 ();
 sg13g2_fill_1 FILLER_26_1143 ();
 sg13g2_fill_1 FILLER_26_1150 ();
 sg13g2_fill_2 FILLER_26_1156 ();
 sg13g2_decap_8 FILLER_26_1163 ();
 sg13g2_decap_8 FILLER_26_1170 ();
 sg13g2_decap_8 FILLER_26_1177 ();
 sg13g2_decap_8 FILLER_26_1184 ();
 sg13g2_decap_8 FILLER_26_1203 ();
 sg13g2_decap_8 FILLER_26_1210 ();
 sg13g2_fill_1 FILLER_26_1217 ();
 sg13g2_decap_8 FILLER_26_1223 ();
 sg13g2_fill_2 FILLER_26_1230 ();
 sg13g2_fill_1 FILLER_26_1241 ();
 sg13g2_fill_2 FILLER_26_1254 ();
 sg13g2_fill_1 FILLER_26_1256 ();
 sg13g2_decap_8 FILLER_26_1262 ();
 sg13g2_fill_1 FILLER_26_1269 ();
 sg13g2_decap_8 FILLER_26_1280 ();
 sg13g2_decap_8 FILLER_26_1287 ();
 sg13g2_decap_8 FILLER_26_1294 ();
 sg13g2_decap_8 FILLER_26_1301 ();
 sg13g2_decap_8 FILLER_26_1308 ();
 sg13g2_decap_8 FILLER_26_1315 ();
 sg13g2_decap_4 FILLER_26_1322 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_23 ();
 sg13g2_decap_8 FILLER_27_33 ();
 sg13g2_decap_8 FILLER_27_40 ();
 sg13g2_decap_8 FILLER_27_47 ();
 sg13g2_decap_4 FILLER_27_54 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_4 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_88 ();
 sg13g2_fill_1 FILLER_27_99 ();
 sg13g2_decap_4 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_109 ();
 sg13g2_decap_8 FILLER_27_114 ();
 sg13g2_decap_8 FILLER_27_121 ();
 sg13g2_decap_8 FILLER_27_128 ();
 sg13g2_fill_2 FILLER_27_135 ();
 sg13g2_decap_8 FILLER_27_145 ();
 sg13g2_decap_8 FILLER_27_152 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_decap_4 FILLER_27_171 ();
 sg13g2_fill_2 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_27_191 ();
 sg13g2_decap_8 FILLER_27_198 ();
 sg13g2_decap_8 FILLER_27_205 ();
 sg13g2_fill_2 FILLER_27_212 ();
 sg13g2_fill_1 FILLER_27_214 ();
 sg13g2_decap_4 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_249 ();
 sg13g2_decap_8 FILLER_27_256 ();
 sg13g2_decap_8 FILLER_27_263 ();
 sg13g2_decap_8 FILLER_27_270 ();
 sg13g2_decap_8 FILLER_27_277 ();
 sg13g2_decap_8 FILLER_27_284 ();
 sg13g2_decap_8 FILLER_27_291 ();
 sg13g2_decap_8 FILLER_27_298 ();
 sg13g2_decap_8 FILLER_27_305 ();
 sg13g2_decap_8 FILLER_27_312 ();
 sg13g2_decap_8 FILLER_27_319 ();
 sg13g2_decap_8 FILLER_27_326 ();
 sg13g2_decap_8 FILLER_27_333 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_fill_2 FILLER_27_347 ();
 sg13g2_decap_8 FILLER_27_355 ();
 sg13g2_decap_8 FILLER_27_362 ();
 sg13g2_decap_8 FILLER_27_369 ();
 sg13g2_decap_8 FILLER_27_376 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_decap_4 FILLER_27_390 ();
 sg13g2_fill_1 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_decap_8 FILLER_27_407 ();
 sg13g2_fill_2 FILLER_27_414 ();
 sg13g2_fill_1 FILLER_27_416 ();
 sg13g2_decap_8 FILLER_27_425 ();
 sg13g2_decap_8 FILLER_27_432 ();
 sg13g2_decap_8 FILLER_27_439 ();
 sg13g2_decap_8 FILLER_27_446 ();
 sg13g2_decap_8 FILLER_27_453 ();
 sg13g2_decap_8 FILLER_27_460 ();
 sg13g2_decap_4 FILLER_27_467 ();
 sg13g2_fill_1 FILLER_27_471 ();
 sg13g2_decap_8 FILLER_27_477 ();
 sg13g2_decap_8 FILLER_27_484 ();
 sg13g2_decap_8 FILLER_27_491 ();
 sg13g2_decap_8 FILLER_27_498 ();
 sg13g2_decap_8 FILLER_27_509 ();
 sg13g2_fill_1 FILLER_27_516 ();
 sg13g2_decap_8 FILLER_27_522 ();
 sg13g2_decap_8 FILLER_27_529 ();
 sg13g2_decap_4 FILLER_27_536 ();
 sg13g2_fill_1 FILLER_27_545 ();
 sg13g2_decap_4 FILLER_27_550 ();
 sg13g2_fill_2 FILLER_27_554 ();
 sg13g2_decap_4 FILLER_27_577 ();
 sg13g2_fill_1 FILLER_27_581 ();
 sg13g2_decap_8 FILLER_27_586 ();
 sg13g2_decap_4 FILLER_27_593 ();
 sg13g2_decap_8 FILLER_27_601 ();
 sg13g2_decap_8 FILLER_27_608 ();
 sg13g2_decap_8 FILLER_27_615 ();
 sg13g2_decap_8 FILLER_27_622 ();
 sg13g2_fill_2 FILLER_27_629 ();
 sg13g2_decap_8 FILLER_27_657 ();
 sg13g2_decap_4 FILLER_27_664 ();
 sg13g2_fill_2 FILLER_27_668 ();
 sg13g2_fill_2 FILLER_27_674 ();
 sg13g2_fill_1 FILLER_27_676 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_4 FILLER_27_707 ();
 sg13g2_fill_2 FILLER_27_711 ();
 sg13g2_decap_8 FILLER_27_717 ();
 sg13g2_decap_8 FILLER_27_724 ();
 sg13g2_decap_8 FILLER_27_731 ();
 sg13g2_decap_8 FILLER_27_738 ();
 sg13g2_fill_2 FILLER_27_745 ();
 sg13g2_fill_1 FILLER_27_747 ();
 sg13g2_decap_8 FILLER_27_752 ();
 sg13g2_decap_8 FILLER_27_759 ();
 sg13g2_decap_8 FILLER_27_766 ();
 sg13g2_decap_8 FILLER_27_773 ();
 sg13g2_decap_8 FILLER_27_810 ();
 sg13g2_fill_1 FILLER_27_817 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_decap_8 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_27_868 ();
 sg13g2_fill_2 FILLER_27_875 ();
 sg13g2_decap_8 FILLER_27_884 ();
 sg13g2_decap_8 FILLER_27_891 ();
 sg13g2_decap_8 FILLER_27_898 ();
 sg13g2_decap_8 FILLER_27_905 ();
 sg13g2_decap_8 FILLER_27_926 ();
 sg13g2_decap_8 FILLER_27_933 ();
 sg13g2_decap_8 FILLER_27_940 ();
 sg13g2_decap_8 FILLER_27_947 ();
 sg13g2_fill_2 FILLER_27_954 ();
 sg13g2_fill_1 FILLER_27_956 ();
 sg13g2_decap_8 FILLER_27_961 ();
 sg13g2_decap_8 FILLER_27_968 ();
 sg13g2_decap_8 FILLER_27_975 ();
 sg13g2_fill_1 FILLER_27_982 ();
 sg13g2_decap_4 FILLER_27_993 ();
 sg13g2_fill_1 FILLER_27_1001 ();
 sg13g2_fill_2 FILLER_27_1016 ();
 sg13g2_decap_8 FILLER_27_1024 ();
 sg13g2_decap_4 FILLER_27_1036 ();
 sg13g2_fill_1 FILLER_27_1040 ();
 sg13g2_decap_8 FILLER_27_1050 ();
 sg13g2_decap_4 FILLER_27_1057 ();
 sg13g2_fill_2 FILLER_27_1076 ();
 sg13g2_decap_8 FILLER_27_1083 ();
 sg13g2_fill_2 FILLER_27_1090 ();
 sg13g2_decap_8 FILLER_27_1096 ();
 sg13g2_decap_8 FILLER_27_1107 ();
 sg13g2_fill_2 FILLER_27_1114 ();
 sg13g2_decap_4 FILLER_27_1124 ();
 sg13g2_decap_4 FILLER_27_1133 ();
 sg13g2_fill_1 FILLER_27_1137 ();
 sg13g2_decap_8 FILLER_27_1156 ();
 sg13g2_decap_4 FILLER_27_1163 ();
 sg13g2_decap_4 FILLER_27_1189 ();
 sg13g2_fill_1 FILLER_27_1193 ();
 sg13g2_fill_1 FILLER_27_1199 ();
 sg13g2_fill_2 FILLER_27_1211 ();
 sg13g2_fill_1 FILLER_27_1213 ();
 sg13g2_decap_8 FILLER_27_1223 ();
 sg13g2_fill_1 FILLER_27_1230 ();
 sg13g2_fill_2 FILLER_27_1247 ();
 sg13g2_fill_1 FILLER_27_1249 ();
 sg13g2_fill_1 FILLER_27_1255 ();
 sg13g2_fill_1 FILLER_27_1265 ();
 sg13g2_fill_2 FILLER_27_1271 ();
 sg13g2_fill_1 FILLER_27_1273 ();
 sg13g2_decap_8 FILLER_27_1279 ();
 sg13g2_decap_8 FILLER_27_1286 ();
 sg13g2_decap_8 FILLER_27_1293 ();
 sg13g2_decap_8 FILLER_27_1300 ();
 sg13g2_decap_8 FILLER_27_1307 ();
 sg13g2_decap_8 FILLER_27_1314 ();
 sg13g2_decap_4 FILLER_27_1321 ();
 sg13g2_fill_1 FILLER_27_1325 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_31 ();
 sg13g2_decap_8 FILLER_28_38 ();
 sg13g2_decap_8 FILLER_28_45 ();
 sg13g2_fill_2 FILLER_28_52 ();
 sg13g2_decap_8 FILLER_28_64 ();
 sg13g2_decap_8 FILLER_28_71 ();
 sg13g2_fill_1 FILLER_28_78 ();
 sg13g2_decap_8 FILLER_28_99 ();
 sg13g2_fill_1 FILLER_28_111 ();
 sg13g2_decap_8 FILLER_28_124 ();
 sg13g2_decap_8 FILLER_28_131 ();
 sg13g2_decap_8 FILLER_28_138 ();
 sg13g2_decap_8 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_162 ();
 sg13g2_fill_1 FILLER_28_169 ();
 sg13g2_decap_8 FILLER_28_174 ();
 sg13g2_decap_8 FILLER_28_181 ();
 sg13g2_decap_8 FILLER_28_188 ();
 sg13g2_decap_8 FILLER_28_195 ();
 sg13g2_decap_8 FILLER_28_202 ();
 sg13g2_decap_8 FILLER_28_209 ();
 sg13g2_fill_2 FILLER_28_224 ();
 sg13g2_fill_1 FILLER_28_226 ();
 sg13g2_decap_8 FILLER_28_256 ();
 sg13g2_decap_8 FILLER_28_263 ();
 sg13g2_decap_8 FILLER_28_270 ();
 sg13g2_decap_4 FILLER_28_277 ();
 sg13g2_fill_2 FILLER_28_281 ();
 sg13g2_decap_8 FILLER_28_295 ();
 sg13g2_decap_8 FILLER_28_302 ();
 sg13g2_decap_4 FILLER_28_309 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_decap_8 FILLER_28_335 ();
 sg13g2_decap_8 FILLER_28_342 ();
 sg13g2_fill_2 FILLER_28_349 ();
 sg13g2_fill_1 FILLER_28_351 ();
 sg13g2_fill_2 FILLER_28_362 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_375 ();
 sg13g2_fill_2 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_4 FILLER_28_420 ();
 sg13g2_fill_1 FILLER_28_424 ();
 sg13g2_decap_8 FILLER_28_441 ();
 sg13g2_decap_8 FILLER_28_448 ();
 sg13g2_decap_8 FILLER_28_455 ();
 sg13g2_decap_8 FILLER_28_462 ();
 sg13g2_decap_4 FILLER_28_469 ();
 sg13g2_fill_2 FILLER_28_477 ();
 sg13g2_fill_1 FILLER_28_479 ();
 sg13g2_decap_4 FILLER_28_485 ();
 sg13g2_fill_1 FILLER_28_489 ();
 sg13g2_decap_8 FILLER_28_495 ();
 sg13g2_decap_8 FILLER_28_502 ();
 sg13g2_decap_4 FILLER_28_509 ();
 sg13g2_fill_1 FILLER_28_513 ();
 sg13g2_decap_8 FILLER_28_575 ();
 sg13g2_decap_8 FILLER_28_582 ();
 sg13g2_decap_8 FILLER_28_589 ();
 sg13g2_decap_4 FILLER_28_596 ();
 sg13g2_decap_8 FILLER_28_607 ();
 sg13g2_decap_8 FILLER_28_614 ();
 sg13g2_decap_8 FILLER_28_621 ();
 sg13g2_decap_8 FILLER_28_628 ();
 sg13g2_decap_4 FILLER_28_635 ();
 sg13g2_decap_4 FILLER_28_643 ();
 sg13g2_fill_2 FILLER_28_647 ();
 sg13g2_fill_1 FILLER_28_654 ();
 sg13g2_fill_2 FILLER_28_686 ();
 sg13g2_fill_1 FILLER_28_688 ();
 sg13g2_fill_1 FILLER_28_697 ();
 sg13g2_decap_8 FILLER_28_731 ();
 sg13g2_decap_8 FILLER_28_738 ();
 sg13g2_fill_2 FILLER_28_745 ();
 sg13g2_fill_2 FILLER_28_751 ();
 sg13g2_fill_1 FILLER_28_753 ();
 sg13g2_decap_8 FILLER_28_773 ();
 sg13g2_decap_8 FILLER_28_780 ();
 sg13g2_decap_8 FILLER_28_787 ();
 sg13g2_fill_1 FILLER_28_794 ();
 sg13g2_decap_8 FILLER_28_804 ();
 sg13g2_fill_1 FILLER_28_811 ();
 sg13g2_decap_8 FILLER_28_816 ();
 sg13g2_decap_8 FILLER_28_823 ();
 sg13g2_decap_8 FILLER_28_830 ();
 sg13g2_decap_8 FILLER_28_837 ();
 sg13g2_decap_8 FILLER_28_844 ();
 sg13g2_decap_8 FILLER_28_851 ();
 sg13g2_decap_8 FILLER_28_858 ();
 sg13g2_decap_8 FILLER_28_865 ();
 sg13g2_decap_8 FILLER_28_872 ();
 sg13g2_decap_8 FILLER_28_879 ();
 sg13g2_decap_8 FILLER_28_886 ();
 sg13g2_decap_8 FILLER_28_893 ();
 sg13g2_fill_2 FILLER_28_900 ();
 sg13g2_decap_4 FILLER_28_907 ();
 sg13g2_fill_2 FILLER_28_926 ();
 sg13g2_fill_2 FILLER_28_937 ();
 sg13g2_decap_8 FILLER_28_943 ();
 sg13g2_fill_1 FILLER_28_950 ();
 sg13g2_decap_4 FILLER_28_961 ();
 sg13g2_fill_1 FILLER_28_965 ();
 sg13g2_decap_8 FILLER_28_971 ();
 sg13g2_fill_1 FILLER_28_978 ();
 sg13g2_fill_1 FILLER_28_993 ();
 sg13g2_fill_2 FILLER_28_998 ();
 sg13g2_decap_8 FILLER_28_1006 ();
 sg13g2_fill_1 FILLER_28_1019 ();
 sg13g2_decap_8 FILLER_28_1024 ();
 sg13g2_decap_8 FILLER_28_1031 ();
 sg13g2_decap_8 FILLER_28_1038 ();
 sg13g2_decap_8 FILLER_28_1045 ();
 sg13g2_decap_8 FILLER_28_1052 ();
 sg13g2_decap_8 FILLER_28_1059 ();
 sg13g2_decap_8 FILLER_28_1066 ();
 sg13g2_decap_8 FILLER_28_1073 ();
 sg13g2_decap_4 FILLER_28_1085 ();
 sg13g2_fill_2 FILLER_28_1089 ();
 sg13g2_decap_8 FILLER_28_1096 ();
 sg13g2_decap_8 FILLER_28_1103 ();
 sg13g2_decap_4 FILLER_28_1110 ();
 sg13g2_fill_2 FILLER_28_1124 ();
 sg13g2_fill_1 FILLER_28_1126 ();
 sg13g2_decap_4 FILLER_28_1135 ();
 sg13g2_decap_8 FILLER_28_1143 ();
 sg13g2_fill_1 FILLER_28_1161 ();
 sg13g2_fill_2 FILLER_28_1167 ();
 sg13g2_fill_1 FILLER_28_1169 ();
 sg13g2_fill_1 FILLER_28_1174 ();
 sg13g2_fill_2 FILLER_28_1185 ();
 sg13g2_decap_8 FILLER_28_1200 ();
 sg13g2_decap_8 FILLER_28_1207 ();
 sg13g2_decap_8 FILLER_28_1214 ();
 sg13g2_decap_8 FILLER_28_1221 ();
 sg13g2_decap_8 FILLER_28_1228 ();
 sg13g2_decap_8 FILLER_28_1235 ();
 sg13g2_decap_4 FILLER_28_1242 ();
 sg13g2_fill_1 FILLER_28_1246 ();
 sg13g2_fill_2 FILLER_28_1252 ();
 sg13g2_fill_2 FILLER_28_1259 ();
 sg13g2_fill_1 FILLER_28_1261 ();
 sg13g2_decap_4 FILLER_28_1267 ();
 sg13g2_fill_1 FILLER_28_1279 ();
 sg13g2_decap_8 FILLER_28_1284 ();
 sg13g2_decap_8 FILLER_28_1291 ();
 sg13g2_decap_8 FILLER_28_1298 ();
 sg13g2_decap_8 FILLER_28_1305 ();
 sg13g2_decap_8 FILLER_28_1312 ();
 sg13g2_decap_8 FILLER_28_1319 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_14 ();
 sg13g2_fill_1 FILLER_29_16 ();
 sg13g2_fill_2 FILLER_29_30 ();
 sg13g2_fill_1 FILLER_29_32 ();
 sg13g2_decap_8 FILLER_29_44 ();
 sg13g2_decap_8 FILLER_29_61 ();
 sg13g2_decap_8 FILLER_29_68 ();
 sg13g2_decap_8 FILLER_29_75 ();
 sg13g2_decap_4 FILLER_29_82 ();
 sg13g2_fill_1 FILLER_29_86 ();
 sg13g2_fill_1 FILLER_29_96 ();
 sg13g2_decap_4 FILLER_29_105 ();
 sg13g2_decap_4 FILLER_29_115 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_129 ();
 sg13g2_decap_8 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_151 ();
 sg13g2_decap_8 FILLER_29_158 ();
 sg13g2_decap_4 FILLER_29_165 ();
 sg13g2_fill_2 FILLER_29_169 ();
 sg13g2_decap_8 FILLER_29_176 ();
 sg13g2_decap_8 FILLER_29_183 ();
 sg13g2_decap_8 FILLER_29_190 ();
 sg13g2_decap_8 FILLER_29_197 ();
 sg13g2_fill_2 FILLER_29_204 ();
 sg13g2_decap_8 FILLER_29_214 ();
 sg13g2_decap_8 FILLER_29_221 ();
 sg13g2_decap_4 FILLER_29_228 ();
 sg13g2_fill_2 FILLER_29_232 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_fill_1 FILLER_29_273 ();
 sg13g2_fill_2 FILLER_29_284 ();
 sg13g2_decap_8 FILLER_29_297 ();
 sg13g2_decap_8 FILLER_29_304 ();
 sg13g2_fill_2 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_313 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_decap_8 FILLER_29_338 ();
 sg13g2_fill_2 FILLER_29_345 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_decap_4 FILLER_29_371 ();
 sg13g2_fill_1 FILLER_29_375 ();
 sg13g2_decap_8 FILLER_29_415 ();
 sg13g2_fill_2 FILLER_29_422 ();
 sg13g2_fill_1 FILLER_29_424 ();
 sg13g2_decap_8 FILLER_29_446 ();
 sg13g2_decap_8 FILLER_29_453 ();
 sg13g2_decap_4 FILLER_29_460 ();
 sg13g2_fill_2 FILLER_29_464 ();
 sg13g2_decap_8 FILLER_29_492 ();
 sg13g2_decap_4 FILLER_29_499 ();
 sg13g2_fill_2 FILLER_29_503 ();
 sg13g2_decap_8 FILLER_29_510 ();
 sg13g2_decap_8 FILLER_29_517 ();
 sg13g2_fill_1 FILLER_29_524 ();
 sg13g2_decap_8 FILLER_29_534 ();
 sg13g2_fill_2 FILLER_29_541 ();
 sg13g2_decap_8 FILLER_29_548 ();
 sg13g2_decap_8 FILLER_29_559 ();
 sg13g2_fill_2 FILLER_29_566 ();
 sg13g2_fill_1 FILLER_29_568 ();
 sg13g2_decap_8 FILLER_29_574 ();
 sg13g2_decap_8 FILLER_29_581 ();
 sg13g2_decap_8 FILLER_29_588 ();
 sg13g2_fill_1 FILLER_29_595 ();
 sg13g2_decap_8 FILLER_29_601 ();
 sg13g2_decap_4 FILLER_29_608 ();
 sg13g2_fill_1 FILLER_29_612 ();
 sg13g2_decap_8 FILLER_29_626 ();
 sg13g2_decap_8 FILLER_29_633 ();
 sg13g2_decap_8 FILLER_29_640 ();
 sg13g2_decap_8 FILLER_29_652 ();
 sg13g2_fill_2 FILLER_29_659 ();
 sg13g2_fill_2 FILLER_29_670 ();
 sg13g2_fill_1 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_677 ();
 sg13g2_decap_8 FILLER_29_684 ();
 sg13g2_decap_8 FILLER_29_691 ();
 sg13g2_decap_8 FILLER_29_698 ();
 sg13g2_decap_8 FILLER_29_705 ();
 sg13g2_decap_8 FILLER_29_712 ();
 sg13g2_decap_8 FILLER_29_719 ();
 sg13g2_decap_8 FILLER_29_726 ();
 sg13g2_fill_2 FILLER_29_733 ();
 sg13g2_fill_1 FILLER_29_735 ();
 sg13g2_decap_8 FILLER_29_766 ();
 sg13g2_decap_4 FILLER_29_773 ();
 sg13g2_fill_2 FILLER_29_777 ();
 sg13g2_decap_8 FILLER_29_800 ();
 sg13g2_decap_8 FILLER_29_807 ();
 sg13g2_decap_8 FILLER_29_814 ();
 sg13g2_decap_8 FILLER_29_821 ();
 sg13g2_decap_8 FILLER_29_828 ();
 sg13g2_decap_8 FILLER_29_835 ();
 sg13g2_decap_8 FILLER_29_842 ();
 sg13g2_decap_4 FILLER_29_849 ();
 sg13g2_decap_4 FILLER_29_858 ();
 sg13g2_fill_2 FILLER_29_862 ();
 sg13g2_decap_4 FILLER_29_869 ();
 sg13g2_decap_8 FILLER_29_878 ();
 sg13g2_fill_2 FILLER_29_889 ();
 sg13g2_fill_1 FILLER_29_899 ();
 sg13g2_decap_4 FILLER_29_904 ();
 sg13g2_decap_4 FILLER_29_942 ();
 sg13g2_fill_1 FILLER_29_957 ();
 sg13g2_decap_4 FILLER_29_963 ();
 sg13g2_fill_1 FILLER_29_967 ();
 sg13g2_fill_2 FILLER_29_987 ();
 sg13g2_fill_2 FILLER_29_997 ();
 sg13g2_decap_8 FILLER_29_1004 ();
 sg13g2_fill_1 FILLER_29_1011 ();
 sg13g2_fill_2 FILLER_29_1017 ();
 sg13g2_decap_8 FILLER_29_1027 ();
 sg13g2_decap_8 FILLER_29_1034 ();
 sg13g2_decap_8 FILLER_29_1041 ();
 sg13g2_decap_8 FILLER_29_1048 ();
 sg13g2_decap_4 FILLER_29_1060 ();
 sg13g2_fill_1 FILLER_29_1064 ();
 sg13g2_decap_8 FILLER_29_1070 ();
 sg13g2_decap_4 FILLER_29_1077 ();
 sg13g2_fill_1 FILLER_29_1081 ();
 sg13g2_decap_8 FILLER_29_1093 ();
 sg13g2_fill_2 FILLER_29_1100 ();
 sg13g2_decap_4 FILLER_29_1107 ();
 sg13g2_fill_1 FILLER_29_1111 ();
 sg13g2_fill_2 FILLER_29_1140 ();
 sg13g2_decap_4 FILLER_29_1147 ();
 sg13g2_fill_1 FILLER_29_1151 ();
 sg13g2_decap_4 FILLER_29_1162 ();
 sg13g2_fill_1 FILLER_29_1166 ();
 sg13g2_decap_4 FILLER_29_1182 ();
 sg13g2_fill_2 FILLER_29_1186 ();
 sg13g2_fill_2 FILLER_29_1203 ();
 sg13g2_decap_4 FILLER_29_1214 ();
 sg13g2_fill_2 FILLER_29_1218 ();
 sg13g2_fill_1 FILLER_29_1228 ();
 sg13g2_fill_2 FILLER_29_1235 ();
 sg13g2_decap_8 FILLER_29_1250 ();
 sg13g2_fill_2 FILLER_29_1257 ();
 sg13g2_fill_1 FILLER_29_1259 ();
 sg13g2_fill_2 FILLER_29_1266 ();
 sg13g2_decap_8 FILLER_29_1282 ();
 sg13g2_decap_8 FILLER_29_1289 ();
 sg13g2_decap_8 FILLER_29_1296 ();
 sg13g2_decap_8 FILLER_29_1303 ();
 sg13g2_decap_8 FILLER_29_1310 ();
 sg13g2_decap_8 FILLER_29_1317 ();
 sg13g2_fill_2 FILLER_29_1324 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_1 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_51 ();
 sg13g2_decap_4 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_73 ();
 sg13g2_decap_4 FILLER_30_78 ();
 sg13g2_decap_8 FILLER_30_87 ();
 sg13g2_fill_2 FILLER_30_94 ();
 sg13g2_decap_8 FILLER_30_100 ();
 sg13g2_decap_8 FILLER_30_107 ();
 sg13g2_decap_8 FILLER_30_114 ();
 sg13g2_decap_4 FILLER_30_128 ();
 sg13g2_fill_1 FILLER_30_132 ();
 sg13g2_decap_8 FILLER_30_155 ();
 sg13g2_decap_8 FILLER_30_162 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_4 FILLER_30_210 ();
 sg13g2_fill_1 FILLER_30_214 ();
 sg13g2_decap_8 FILLER_30_236 ();
 sg13g2_decap_4 FILLER_30_243 ();
 sg13g2_fill_2 FILLER_30_247 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_fill_2 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_268 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_fill_2 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_303 ();
 sg13g2_decap_4 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_334 ();
 sg13g2_fill_2 FILLER_30_341 ();
 sg13g2_fill_1 FILLER_30_343 ();
 sg13g2_fill_2 FILLER_30_349 ();
 sg13g2_decap_8 FILLER_30_355 ();
 sg13g2_decap_8 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_30_369 ();
 sg13g2_decap_8 FILLER_30_376 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_fill_1 FILLER_30_420 ();
 sg13g2_decap_8 FILLER_30_437 ();
 sg13g2_fill_1 FILLER_30_444 ();
 sg13g2_decap_8 FILLER_30_458 ();
 sg13g2_decap_8 FILLER_30_465 ();
 sg13g2_decap_4 FILLER_30_476 ();
 sg13g2_decap_8 FILLER_30_490 ();
 sg13g2_decap_8 FILLER_30_497 ();
 sg13g2_decap_8 FILLER_30_504 ();
 sg13g2_decap_8 FILLER_30_511 ();
 sg13g2_decap_8 FILLER_30_518 ();
 sg13g2_decap_8 FILLER_30_525 ();
 sg13g2_decap_8 FILLER_30_532 ();
 sg13g2_decap_8 FILLER_30_539 ();
 sg13g2_decap_8 FILLER_30_546 ();
 sg13g2_decap_8 FILLER_30_553 ();
 sg13g2_fill_2 FILLER_30_560 ();
 sg13g2_decap_8 FILLER_30_567 ();
 sg13g2_decap_8 FILLER_30_574 ();
 sg13g2_decap_8 FILLER_30_581 ();
 sg13g2_decap_8 FILLER_30_588 ();
 sg13g2_decap_8 FILLER_30_595 ();
 sg13g2_decap_8 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_4 FILLER_30_616 ();
 sg13g2_fill_2 FILLER_30_620 ();
 sg13g2_decap_4 FILLER_30_627 ();
 sg13g2_decap_8 FILLER_30_635 ();
 sg13g2_decap_8 FILLER_30_642 ();
 sg13g2_decap_4 FILLER_30_675 ();
 sg13g2_fill_1 FILLER_30_679 ();
 sg13g2_decap_4 FILLER_30_695 ();
 sg13g2_fill_2 FILLER_30_699 ();
 sg13g2_decap_8 FILLER_30_705 ();
 sg13g2_decap_8 FILLER_30_712 ();
 sg13g2_decap_8 FILLER_30_719 ();
 sg13g2_decap_8 FILLER_30_726 ();
 sg13g2_decap_8 FILLER_30_733 ();
 sg13g2_fill_2 FILLER_30_740 ();
 sg13g2_decap_8 FILLER_30_746 ();
 sg13g2_decap_8 FILLER_30_753 ();
 sg13g2_decap_8 FILLER_30_760 ();
 sg13g2_decap_8 FILLER_30_767 ();
 sg13g2_decap_4 FILLER_30_774 ();
 sg13g2_fill_1 FILLER_30_778 ();
 sg13g2_decap_8 FILLER_30_809 ();
 sg13g2_decap_8 FILLER_30_816 ();
 sg13g2_decap_8 FILLER_30_823 ();
 sg13g2_decap_8 FILLER_30_830 ();
 sg13g2_decap_8 FILLER_30_837 ();
 sg13g2_decap_8 FILLER_30_844 ();
 sg13g2_decap_8 FILLER_30_851 ();
 sg13g2_decap_8 FILLER_30_858 ();
 sg13g2_decap_8 FILLER_30_865 ();
 sg13g2_decap_8 FILLER_30_872 ();
 sg13g2_fill_2 FILLER_30_879 ();
 sg13g2_decap_4 FILLER_30_885 ();
 sg13g2_fill_2 FILLER_30_889 ();
 sg13g2_decap_8 FILLER_30_896 ();
 sg13g2_fill_2 FILLER_30_903 ();
 sg13g2_fill_1 FILLER_30_905 ();
 sg13g2_decap_4 FILLER_30_910 ();
 sg13g2_fill_1 FILLER_30_914 ();
 sg13g2_decap_8 FILLER_30_919 ();
 sg13g2_fill_2 FILLER_30_926 ();
 sg13g2_fill_1 FILLER_30_928 ();
 sg13g2_decap_4 FILLER_30_949 ();
 sg13g2_decap_8 FILLER_30_961 ();
 sg13g2_decap_8 FILLER_30_968 ();
 sg13g2_decap_4 FILLER_30_975 ();
 sg13g2_fill_2 FILLER_30_979 ();
 sg13g2_fill_2 FILLER_30_986 ();
 sg13g2_fill_1 FILLER_30_988 ();
 sg13g2_decap_8 FILLER_30_999 ();
 sg13g2_decap_4 FILLER_30_1006 ();
 sg13g2_fill_2 FILLER_30_1010 ();
 sg13g2_fill_2 FILLER_30_1017 ();
 sg13g2_fill_1 FILLER_30_1019 ();
 sg13g2_decap_8 FILLER_30_1024 ();
 sg13g2_decap_8 FILLER_30_1031 ();
 sg13g2_decap_8 FILLER_30_1038 ();
 sg13g2_fill_2 FILLER_30_1045 ();
 sg13g2_fill_1 FILLER_30_1047 ();
 sg13g2_fill_1 FILLER_30_1065 ();
 sg13g2_decap_8 FILLER_30_1077 ();
 sg13g2_decap_8 FILLER_30_1084 ();
 sg13g2_fill_2 FILLER_30_1091 ();
 sg13g2_fill_1 FILLER_30_1093 ();
 sg13g2_decap_8 FILLER_30_1107 ();
 sg13g2_decap_8 FILLER_30_1114 ();
 sg13g2_decap_8 FILLER_30_1121 ();
 sg13g2_decap_8 FILLER_30_1128 ();
 sg13g2_decap_8 FILLER_30_1140 ();
 sg13g2_fill_2 FILLER_30_1147 ();
 sg13g2_fill_1 FILLER_30_1149 ();
 sg13g2_fill_2 FILLER_30_1154 ();
 sg13g2_fill_1 FILLER_30_1156 ();
 sg13g2_decap_4 FILLER_30_1163 ();
 sg13g2_fill_2 FILLER_30_1167 ();
 sg13g2_fill_1 FILLER_30_1175 ();
 sg13g2_decap_8 FILLER_30_1189 ();
 sg13g2_decap_8 FILLER_30_1196 ();
 sg13g2_decap_8 FILLER_30_1203 ();
 sg13g2_decap_4 FILLER_30_1210 ();
 sg13g2_fill_2 FILLER_30_1214 ();
 sg13g2_decap_4 FILLER_30_1220 ();
 sg13g2_fill_2 FILLER_30_1224 ();
 sg13g2_fill_1 FILLER_30_1231 ();
 sg13g2_fill_2 FILLER_30_1245 ();
 sg13g2_fill_2 FILLER_30_1252 ();
 sg13g2_decap_8 FILLER_30_1259 ();
 sg13g2_decap_8 FILLER_30_1270 ();
 sg13g2_fill_2 FILLER_30_1277 ();
 sg13g2_fill_1 FILLER_30_1279 ();
 sg13g2_decap_8 FILLER_30_1284 ();
 sg13g2_decap_8 FILLER_30_1291 ();
 sg13g2_decap_8 FILLER_30_1298 ();
 sg13g2_decap_8 FILLER_30_1305 ();
 sg13g2_decap_8 FILLER_30_1312 ();
 sg13g2_decap_8 FILLER_30_1319 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_4 FILLER_31_35 ();
 sg13g2_fill_1 FILLER_31_39 ();
 sg13g2_decap_8 FILLER_31_50 ();
 sg13g2_fill_1 FILLER_31_57 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_84 ();
 sg13g2_decap_4 FILLER_31_92 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_decap_8 FILLER_31_102 ();
 sg13g2_decap_8 FILLER_31_109 ();
 sg13g2_decap_8 FILLER_31_116 ();
 sg13g2_decap_4 FILLER_31_123 ();
 sg13g2_decap_8 FILLER_31_132 ();
 sg13g2_fill_1 FILLER_31_139 ();
 sg13g2_decap_4 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_156 ();
 sg13g2_decap_8 FILLER_31_162 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_decap_8 FILLER_31_183 ();
 sg13g2_decap_8 FILLER_31_190 ();
 sg13g2_decap_8 FILLER_31_197 ();
 sg13g2_decap_8 FILLER_31_204 ();
 sg13g2_decap_8 FILLER_31_211 ();
 sg13g2_decap_8 FILLER_31_218 ();
 sg13g2_decap_8 FILLER_31_225 ();
 sg13g2_decap_8 FILLER_31_232 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_decap_8 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_decap_8 FILLER_31_260 ();
 sg13g2_decap_8 FILLER_31_267 ();
 sg13g2_decap_8 FILLER_31_274 ();
 sg13g2_decap_8 FILLER_31_281 ();
 sg13g2_fill_1 FILLER_31_288 ();
 sg13g2_fill_2 FILLER_31_293 ();
 sg13g2_fill_1 FILLER_31_295 ();
 sg13g2_decap_8 FILLER_31_305 ();
 sg13g2_decap_4 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_fill_1 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_363 ();
 sg13g2_decap_8 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_31_384 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_8 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_31_412 ();
 sg13g2_decap_8 FILLER_31_419 ();
 sg13g2_decap_8 FILLER_31_426 ();
 sg13g2_decap_8 FILLER_31_433 ();
 sg13g2_fill_2 FILLER_31_440 ();
 sg13g2_fill_1 FILLER_31_442 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_decap_8 FILLER_31_462 ();
 sg13g2_decap_8 FILLER_31_469 ();
 sg13g2_fill_1 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_516 ();
 sg13g2_fill_2 FILLER_31_528 ();
 sg13g2_fill_1 FILLER_31_530 ();
 sg13g2_decap_4 FILLER_31_539 ();
 sg13g2_fill_2 FILLER_31_543 ();
 sg13g2_decap_8 FILLER_31_549 ();
 sg13g2_decap_8 FILLER_31_556 ();
 sg13g2_fill_1 FILLER_31_563 ();
 sg13g2_fill_2 FILLER_31_573 ();
 sg13g2_fill_2 FILLER_31_596 ();
 sg13g2_fill_1 FILLER_31_598 ();
 sg13g2_decap_8 FILLER_31_634 ();
 sg13g2_decap_8 FILLER_31_641 ();
 sg13g2_decap_8 FILLER_31_648 ();
 sg13g2_decap_8 FILLER_31_659 ();
 sg13g2_decap_4 FILLER_31_666 ();
 sg13g2_fill_2 FILLER_31_670 ();
 sg13g2_decap_8 FILLER_31_706 ();
 sg13g2_decap_8 FILLER_31_713 ();
 sg13g2_decap_8 FILLER_31_720 ();
 sg13g2_decap_8 FILLER_31_727 ();
 sg13g2_decap_8 FILLER_31_734 ();
 sg13g2_decap_8 FILLER_31_741 ();
 sg13g2_decap_8 FILLER_31_748 ();
 sg13g2_decap_8 FILLER_31_755 ();
 sg13g2_decap_8 FILLER_31_762 ();
 sg13g2_decap_8 FILLER_31_769 ();
 sg13g2_decap_8 FILLER_31_776 ();
 sg13g2_decap_8 FILLER_31_783 ();
 sg13g2_decap_8 FILLER_31_794 ();
 sg13g2_decap_8 FILLER_31_801 ();
 sg13g2_decap_8 FILLER_31_808 ();
 sg13g2_decap_8 FILLER_31_815 ();
 sg13g2_decap_8 FILLER_31_822 ();
 sg13g2_decap_8 FILLER_31_829 ();
 sg13g2_decap_8 FILLER_31_836 ();
 sg13g2_decap_8 FILLER_31_843 ();
 sg13g2_decap_8 FILLER_31_850 ();
 sg13g2_decap_8 FILLER_31_857 ();
 sg13g2_fill_2 FILLER_31_864 ();
 sg13g2_fill_1 FILLER_31_866 ();
 sg13g2_decap_8 FILLER_31_874 ();
 sg13g2_fill_2 FILLER_31_881 ();
 sg13g2_fill_1 FILLER_31_887 ();
 sg13g2_decap_8 FILLER_31_898 ();
 sg13g2_decap_8 FILLER_31_905 ();
 sg13g2_decap_8 FILLER_31_912 ();
 sg13g2_fill_1 FILLER_31_919 ();
 sg13g2_decap_8 FILLER_31_928 ();
 sg13g2_decap_8 FILLER_31_935 ();
 sg13g2_decap_8 FILLER_31_942 ();
 sg13g2_fill_2 FILLER_31_949 ();
 sg13g2_fill_1 FILLER_31_951 ();
 sg13g2_fill_2 FILLER_31_963 ();
 sg13g2_decap_8 FILLER_31_974 ();
 sg13g2_decap_8 FILLER_31_981 ();
 sg13g2_decap_4 FILLER_31_988 ();
 sg13g2_fill_2 FILLER_31_992 ();
 sg13g2_decap_4 FILLER_31_1003 ();
 sg13g2_decap_8 FILLER_31_1017 ();
 sg13g2_fill_2 FILLER_31_1024 ();
 sg13g2_fill_1 FILLER_31_1026 ();
 sg13g2_decap_8 FILLER_31_1032 ();
 sg13g2_decap_4 FILLER_31_1039 ();
 sg13g2_decap_8 FILLER_31_1047 ();
 sg13g2_decap_8 FILLER_31_1054 ();
 sg13g2_decap_4 FILLER_31_1061 ();
 sg13g2_decap_4 FILLER_31_1075 ();
 sg13g2_fill_2 FILLER_31_1079 ();
 sg13g2_decap_4 FILLER_31_1086 ();
 sg13g2_fill_1 FILLER_31_1090 ();
 sg13g2_fill_1 FILLER_31_1096 ();
 sg13g2_fill_1 FILLER_31_1106 ();
 sg13g2_decap_4 FILLER_31_1112 ();
 sg13g2_fill_2 FILLER_31_1116 ();
 sg13g2_fill_2 FILLER_31_1140 ();
 sg13g2_decap_8 FILLER_31_1147 ();
 sg13g2_fill_2 FILLER_31_1154 ();
 sg13g2_fill_1 FILLER_31_1156 ();
 sg13g2_fill_2 FILLER_31_1162 ();
 sg13g2_decap_4 FILLER_31_1168 ();
 sg13g2_fill_2 FILLER_31_1172 ();
 sg13g2_decap_8 FILLER_31_1180 ();
 sg13g2_decap_4 FILLER_31_1187 ();
 sg13g2_fill_2 FILLER_31_1191 ();
 sg13g2_decap_8 FILLER_31_1200 ();
 sg13g2_fill_2 FILLER_31_1207 ();
 sg13g2_decap_4 FILLER_31_1213 ();
 sg13g2_decap_8 FILLER_31_1222 ();
 sg13g2_fill_1 FILLER_31_1229 ();
 sg13g2_decap_8 FILLER_31_1242 ();
 sg13g2_decap_4 FILLER_31_1249 ();
 sg13g2_decap_4 FILLER_31_1258 ();
 sg13g2_decap_8 FILLER_31_1267 ();
 sg13g2_decap_8 FILLER_31_1283 ();
 sg13g2_decap_8 FILLER_31_1290 ();
 sg13g2_decap_8 FILLER_31_1297 ();
 sg13g2_decap_8 FILLER_31_1304 ();
 sg13g2_decap_8 FILLER_31_1311 ();
 sg13g2_decap_8 FILLER_31_1318 ();
 sg13g2_fill_1 FILLER_31_1325 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_4 FILLER_32_35 ();
 sg13g2_fill_1 FILLER_32_39 ();
 sg13g2_fill_2 FILLER_32_44 ();
 sg13g2_fill_1 FILLER_32_46 ();
 sg13g2_decap_4 FILLER_32_53 ();
 sg13g2_fill_2 FILLER_32_57 ();
 sg13g2_decap_8 FILLER_32_69 ();
 sg13g2_decap_8 FILLER_32_76 ();
 sg13g2_fill_2 FILLER_32_83 ();
 sg13g2_decap_8 FILLER_32_89 ();
 sg13g2_decap_8 FILLER_32_96 ();
 sg13g2_decap_8 FILLER_32_103 ();
 sg13g2_fill_2 FILLER_32_110 ();
 sg13g2_fill_2 FILLER_32_116 ();
 sg13g2_fill_1 FILLER_32_118 ();
 sg13g2_decap_8 FILLER_32_134 ();
 sg13g2_decap_8 FILLER_32_141 ();
 sg13g2_fill_2 FILLER_32_148 ();
 sg13g2_decap_8 FILLER_32_159 ();
 sg13g2_fill_1 FILLER_32_166 ();
 sg13g2_fill_1 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_4 FILLER_32_203 ();
 sg13g2_fill_1 FILLER_32_207 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_fill_1 FILLER_32_241 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_decap_4 FILLER_32_270 ();
 sg13g2_fill_1 FILLER_32_274 ();
 sg13g2_decap_8 FILLER_32_289 ();
 sg13g2_decap_8 FILLER_32_296 ();
 sg13g2_decap_8 FILLER_32_303 ();
 sg13g2_decap_8 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_decap_8 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_decap_4 FILLER_32_351 ();
 sg13g2_fill_2 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_4 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_decap_4 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_426 ();
 sg13g2_fill_2 FILLER_32_433 ();
 sg13g2_fill_1 FILLER_32_435 ();
 sg13g2_decap_8 FILLER_32_444 ();
 sg13g2_decap_8 FILLER_32_451 ();
 sg13g2_decap_8 FILLER_32_458 ();
 sg13g2_decap_8 FILLER_32_465 ();
 sg13g2_decap_8 FILLER_32_472 ();
 sg13g2_fill_2 FILLER_32_479 ();
 sg13g2_decap_4 FILLER_32_485 ();
 sg13g2_fill_1 FILLER_32_489 ();
 sg13g2_decap_8 FILLER_32_494 ();
 sg13g2_decap_4 FILLER_32_501 ();
 sg13g2_fill_1 FILLER_32_505 ();
 sg13g2_fill_1 FILLER_32_510 ();
 sg13g2_fill_1 FILLER_32_547 ();
 sg13g2_decap_8 FILLER_32_600 ();
 sg13g2_decap_8 FILLER_32_607 ();
 sg13g2_fill_2 FILLER_32_614 ();
 sg13g2_fill_1 FILLER_32_616 ();
 sg13g2_decap_8 FILLER_32_621 ();
 sg13g2_decap_8 FILLER_32_628 ();
 sg13g2_decap_8 FILLER_32_635 ();
 sg13g2_decap_8 FILLER_32_642 ();
 sg13g2_decap_8 FILLER_32_649 ();
 sg13g2_decap_8 FILLER_32_656 ();
 sg13g2_decap_8 FILLER_32_663 ();
 sg13g2_decap_8 FILLER_32_670 ();
 sg13g2_decap_8 FILLER_32_677 ();
 sg13g2_decap_8 FILLER_32_684 ();
 sg13g2_fill_2 FILLER_32_691 ();
 sg13g2_decap_8 FILLER_32_697 ();
 sg13g2_fill_2 FILLER_32_704 ();
 sg13g2_decap_8 FILLER_32_732 ();
 sg13g2_decap_8 FILLER_32_739 ();
 sg13g2_fill_1 FILLER_32_746 ();
 sg13g2_decap_8 FILLER_32_751 ();
 sg13g2_fill_2 FILLER_32_758 ();
 sg13g2_fill_1 FILLER_32_760 ();
 sg13g2_fill_2 FILLER_32_769 ();
 sg13g2_fill_1 FILLER_32_781 ();
 sg13g2_decap_8 FILLER_32_787 ();
 sg13g2_decap_8 FILLER_32_794 ();
 sg13g2_decap_8 FILLER_32_801 ();
 sg13g2_decap_8 FILLER_32_808 ();
 sg13g2_decap_8 FILLER_32_815 ();
 sg13g2_decap_8 FILLER_32_822 ();
 sg13g2_decap_8 FILLER_32_829 ();
 sg13g2_decap_8 FILLER_32_836 ();
 sg13g2_decap_8 FILLER_32_843 ();
 sg13g2_decap_8 FILLER_32_850 ();
 sg13g2_decap_8 FILLER_32_857 ();
 sg13g2_decap_8 FILLER_32_864 ();
 sg13g2_decap_8 FILLER_32_871 ();
 sg13g2_decap_4 FILLER_32_878 ();
 sg13g2_decap_8 FILLER_32_891 ();
 sg13g2_decap_8 FILLER_32_898 ();
 sg13g2_decap_8 FILLER_32_905 ();
 sg13g2_decap_8 FILLER_32_912 ();
 sg13g2_fill_2 FILLER_32_919 ();
 sg13g2_fill_2 FILLER_32_929 ();
 sg13g2_decap_8 FILLER_32_936 ();
 sg13g2_decap_4 FILLER_32_943 ();
 sg13g2_decap_8 FILLER_32_951 ();
 sg13g2_fill_2 FILLER_32_968 ();
 sg13g2_fill_2 FILLER_32_989 ();
 sg13g2_fill_1 FILLER_32_1004 ();
 sg13g2_fill_1 FILLER_32_1013 ();
 sg13g2_decap_8 FILLER_32_1019 ();
 sg13g2_decap_8 FILLER_32_1026 ();
 sg13g2_decap_8 FILLER_32_1033 ();
 sg13g2_decap_4 FILLER_32_1040 ();
 sg13g2_decap_8 FILLER_32_1049 ();
 sg13g2_decap_4 FILLER_32_1056 ();
 sg13g2_decap_8 FILLER_32_1073 ();
 sg13g2_decap_8 FILLER_32_1080 ();
 sg13g2_decap_8 FILLER_32_1087 ();
 sg13g2_fill_2 FILLER_32_1098 ();
 sg13g2_decap_8 FILLER_32_1111 ();
 sg13g2_fill_2 FILLER_32_1118 ();
 sg13g2_fill_1 FILLER_32_1135 ();
 sg13g2_fill_2 FILLER_32_1155 ();
 sg13g2_decap_8 FILLER_32_1162 ();
 sg13g2_decap_4 FILLER_32_1169 ();
 sg13g2_fill_1 FILLER_32_1173 ();
 sg13g2_fill_1 FILLER_32_1192 ();
 sg13g2_decap_8 FILLER_32_1197 ();
 sg13g2_decap_4 FILLER_32_1204 ();
 sg13g2_fill_2 FILLER_32_1218 ();
 sg13g2_fill_1 FILLER_32_1225 ();
 sg13g2_fill_2 FILLER_32_1230 ();
 sg13g2_decap_4 FILLER_32_1241 ();
 sg13g2_decap_8 FILLER_32_1250 ();
 sg13g2_decap_4 FILLER_32_1257 ();
 sg13g2_decap_4 FILLER_32_1265 ();
 sg13g2_fill_1 FILLER_32_1283 ();
 sg13g2_decap_8 FILLER_32_1289 ();
 sg13g2_decap_8 FILLER_32_1296 ();
 sg13g2_decap_8 FILLER_32_1303 ();
 sg13g2_decap_8 FILLER_32_1310 ();
 sg13g2_decap_8 FILLER_32_1317 ();
 sg13g2_fill_2 FILLER_32_1324 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_4 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_60 ();
 sg13g2_decap_4 FILLER_33_65 ();
 sg13g2_decap_8 FILLER_33_73 ();
 sg13g2_decap_8 FILLER_33_80 ();
 sg13g2_decap_8 FILLER_33_87 ();
 sg13g2_decap_8 FILLER_33_94 ();
 sg13g2_decap_8 FILLER_33_101 ();
 sg13g2_decap_8 FILLER_33_108 ();
 sg13g2_decap_8 FILLER_33_115 ();
 sg13g2_decap_8 FILLER_33_132 ();
 sg13g2_decap_8 FILLER_33_139 ();
 sg13g2_decap_4 FILLER_33_146 ();
 sg13g2_fill_1 FILLER_33_150 ();
 sg13g2_decap_8 FILLER_33_159 ();
 sg13g2_decap_8 FILLER_33_166 ();
 sg13g2_decap_8 FILLER_33_173 ();
 sg13g2_decap_8 FILLER_33_180 ();
 sg13g2_decap_8 FILLER_33_187 ();
 sg13g2_decap_8 FILLER_33_194 ();
 sg13g2_decap_8 FILLER_33_201 ();
 sg13g2_decap_8 FILLER_33_208 ();
 sg13g2_decap_8 FILLER_33_215 ();
 sg13g2_decap_8 FILLER_33_222 ();
 sg13g2_decap_8 FILLER_33_229 ();
 sg13g2_decap_8 FILLER_33_236 ();
 sg13g2_decap_8 FILLER_33_243 ();
 sg13g2_decap_8 FILLER_33_250 ();
 sg13g2_decap_8 FILLER_33_257 ();
 sg13g2_decap_4 FILLER_33_264 ();
 sg13g2_fill_1 FILLER_33_282 ();
 sg13g2_decap_8 FILLER_33_304 ();
 sg13g2_decap_8 FILLER_33_311 ();
 sg13g2_decap_8 FILLER_33_318 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_345 ();
 sg13g2_decap_8 FILLER_33_352 ();
 sg13g2_decap_8 FILLER_33_359 ();
 sg13g2_decap_8 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_380 ();
 sg13g2_fill_1 FILLER_33_395 ();
 sg13g2_fill_1 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_409 ();
 sg13g2_decap_8 FILLER_33_431 ();
 sg13g2_fill_2 FILLER_33_438 ();
 sg13g2_fill_1 FILLER_33_440 ();
 sg13g2_decap_8 FILLER_33_453 ();
 sg13g2_decap_8 FILLER_33_460 ();
 sg13g2_decap_8 FILLER_33_467 ();
 sg13g2_decap_8 FILLER_33_474 ();
 sg13g2_decap_8 FILLER_33_481 ();
 sg13g2_decap_8 FILLER_33_488 ();
 sg13g2_decap_8 FILLER_33_495 ();
 sg13g2_decap_8 FILLER_33_502 ();
 sg13g2_decap_8 FILLER_33_509 ();
 sg13g2_decap_8 FILLER_33_516 ();
 sg13g2_fill_2 FILLER_33_523 ();
 sg13g2_decap_8 FILLER_33_529 ();
 sg13g2_decap_8 FILLER_33_536 ();
 sg13g2_decap_8 FILLER_33_543 ();
 sg13g2_decap_4 FILLER_33_550 ();
 sg13g2_fill_2 FILLER_33_554 ();
 sg13g2_decap_8 FILLER_33_560 ();
 sg13g2_fill_1 FILLER_33_567 ();
 sg13g2_decap_8 FILLER_33_573 ();
 sg13g2_decap_8 FILLER_33_584 ();
 sg13g2_decap_8 FILLER_33_591 ();
 sg13g2_decap_8 FILLER_33_598 ();
 sg13g2_decap_8 FILLER_33_605 ();
 sg13g2_decap_8 FILLER_33_612 ();
 sg13g2_decap_8 FILLER_33_619 ();
 sg13g2_decap_8 FILLER_33_626 ();
 sg13g2_decap_8 FILLER_33_633 ();
 sg13g2_decap_8 FILLER_33_679 ();
 sg13g2_fill_2 FILLER_33_686 ();
 sg13g2_fill_1 FILLER_33_688 ();
 sg13g2_decap_4 FILLER_33_710 ();
 sg13g2_fill_1 FILLER_33_714 ();
 sg13g2_decap_8 FILLER_33_719 ();
 sg13g2_decap_8 FILLER_33_726 ();
 sg13g2_decap_8 FILLER_33_733 ();
 sg13g2_decap_8 FILLER_33_770 ();
 sg13g2_fill_2 FILLER_33_777 ();
 sg13g2_fill_1 FILLER_33_779 ();
 sg13g2_decap_8 FILLER_33_788 ();
 sg13g2_fill_2 FILLER_33_795 ();
 sg13g2_decap_8 FILLER_33_800 ();
 sg13g2_decap_8 FILLER_33_807 ();
 sg13g2_decap_8 FILLER_33_814 ();
 sg13g2_fill_2 FILLER_33_821 ();
 sg13g2_decap_8 FILLER_33_827 ();
 sg13g2_decap_8 FILLER_33_834 ();
 sg13g2_decap_8 FILLER_33_841 ();
 sg13g2_decap_8 FILLER_33_848 ();
 sg13g2_decap_8 FILLER_33_855 ();
 sg13g2_decap_8 FILLER_33_862 ();
 sg13g2_decap_4 FILLER_33_869 ();
 sg13g2_fill_2 FILLER_33_873 ();
 sg13g2_decap_4 FILLER_33_884 ();
 sg13g2_fill_1 FILLER_33_888 ();
 sg13g2_decap_8 FILLER_33_894 ();
 sg13g2_fill_2 FILLER_33_901 ();
 sg13g2_fill_1 FILLER_33_903 ();
 sg13g2_fill_2 FILLER_33_912 ();
 sg13g2_decap_4 FILLER_33_920 ();
 sg13g2_fill_1 FILLER_33_929 ();
 sg13g2_decap_4 FILLER_33_935 ();
 sg13g2_fill_2 FILLER_33_947 ();
 sg13g2_fill_1 FILLER_33_949 ();
 sg13g2_fill_1 FILLER_33_955 ();
 sg13g2_decap_4 FILLER_33_985 ();
 sg13g2_fill_1 FILLER_33_989 ();
 sg13g2_fill_2 FILLER_33_995 ();
 sg13g2_fill_2 FILLER_33_1026 ();
 sg13g2_decap_8 FILLER_33_1051 ();
 sg13g2_fill_2 FILLER_33_1058 ();
 sg13g2_decap_4 FILLER_33_1065 ();
 sg13g2_fill_2 FILLER_33_1069 ();
 sg13g2_decap_4 FILLER_33_1079 ();
 sg13g2_fill_1 FILLER_33_1083 ();
 sg13g2_decap_8 FILLER_33_1089 ();
 sg13g2_decap_8 FILLER_33_1096 ();
 sg13g2_decap_8 FILLER_33_1103 ();
 sg13g2_fill_2 FILLER_33_1110 ();
 sg13g2_decap_8 FILLER_33_1116 ();
 sg13g2_fill_2 FILLER_33_1123 ();
 sg13g2_fill_1 FILLER_33_1136 ();
 sg13g2_decap_4 FILLER_33_1141 ();
 sg13g2_fill_1 FILLER_33_1145 ();
 sg13g2_decap_8 FILLER_33_1150 ();
 sg13g2_fill_2 FILLER_33_1157 ();
 sg13g2_fill_1 FILLER_33_1159 ();
 sg13g2_fill_2 FILLER_33_1165 ();
 sg13g2_fill_2 FILLER_33_1172 ();
 sg13g2_fill_1 FILLER_33_1174 ();
 sg13g2_decap_8 FILLER_33_1180 ();
 sg13g2_fill_1 FILLER_33_1187 ();
 sg13g2_decap_8 FILLER_33_1192 ();
 sg13g2_decap_8 FILLER_33_1199 ();
 sg13g2_fill_1 FILLER_33_1206 ();
 sg13g2_fill_1 FILLER_33_1214 ();
 sg13g2_decap_4 FILLER_33_1220 ();
 sg13g2_fill_1 FILLER_33_1224 ();
 sg13g2_fill_2 FILLER_33_1234 ();
 sg13g2_decap_8 FILLER_33_1240 ();
 sg13g2_fill_1 FILLER_33_1247 ();
 sg13g2_fill_2 FILLER_33_1261 ();
 sg13g2_fill_1 FILLER_33_1263 ();
 sg13g2_fill_2 FILLER_33_1278 ();
 sg13g2_decap_8 FILLER_33_1284 ();
 sg13g2_decap_8 FILLER_33_1291 ();
 sg13g2_decap_8 FILLER_33_1298 ();
 sg13g2_decap_8 FILLER_33_1305 ();
 sg13g2_decap_8 FILLER_33_1312 ();
 sg13g2_decap_8 FILLER_33_1319 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_64 ();
 sg13g2_decap_8 FILLER_34_71 ();
 sg13g2_decap_8 FILLER_34_78 ();
 sg13g2_decap_8 FILLER_34_85 ();
 sg13g2_decap_8 FILLER_34_92 ();
 sg13g2_decap_8 FILLER_34_99 ();
 sg13g2_decap_8 FILLER_34_106 ();
 sg13g2_decap_8 FILLER_34_113 ();
 sg13g2_decap_8 FILLER_34_120 ();
 sg13g2_fill_1 FILLER_34_127 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_fill_1 FILLER_34_266 ();
 sg13g2_decap_4 FILLER_34_277 ();
 sg13g2_decap_8 FILLER_34_291 ();
 sg13g2_decap_8 FILLER_34_298 ();
 sg13g2_decap_8 FILLER_34_305 ();
 sg13g2_decap_8 FILLER_34_312 ();
 sg13g2_decap_8 FILLER_34_319 ();
 sg13g2_fill_2 FILLER_34_326 ();
 sg13g2_fill_1 FILLER_34_328 ();
 sg13g2_decap_8 FILLER_34_355 ();
 sg13g2_decap_8 FILLER_34_362 ();
 sg13g2_decap_8 FILLER_34_369 ();
 sg13g2_decap_8 FILLER_34_376 ();
 sg13g2_decap_4 FILLER_34_383 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_410 ();
 sg13g2_decap_8 FILLER_34_417 ();
 sg13g2_decap_8 FILLER_34_424 ();
 sg13g2_decap_8 FILLER_34_431 ();
 sg13g2_decap_8 FILLER_34_438 ();
 sg13g2_decap_8 FILLER_34_445 ();
 sg13g2_decap_8 FILLER_34_452 ();
 sg13g2_decap_8 FILLER_34_459 ();
 sg13g2_decap_8 FILLER_34_466 ();
 sg13g2_decap_4 FILLER_34_473 ();
 sg13g2_fill_2 FILLER_34_477 ();
 sg13g2_decap_8 FILLER_34_484 ();
 sg13g2_decap_8 FILLER_34_491 ();
 sg13g2_fill_2 FILLER_34_498 ();
 sg13g2_decap_8 FILLER_34_505 ();
 sg13g2_decap_8 FILLER_34_512 ();
 sg13g2_decap_8 FILLER_34_519 ();
 sg13g2_decap_8 FILLER_34_526 ();
 sg13g2_decap_8 FILLER_34_533 ();
 sg13g2_decap_8 FILLER_34_540 ();
 sg13g2_decap_8 FILLER_34_547 ();
 sg13g2_decap_8 FILLER_34_554 ();
 sg13g2_decap_4 FILLER_34_561 ();
 sg13g2_decap_8 FILLER_34_569 ();
 sg13g2_decap_8 FILLER_34_576 ();
 sg13g2_decap_8 FILLER_34_583 ();
 sg13g2_decap_8 FILLER_34_590 ();
 sg13g2_decap_8 FILLER_34_597 ();
 sg13g2_decap_8 FILLER_34_604 ();
 sg13g2_decap_8 FILLER_34_611 ();
 sg13g2_decap_8 FILLER_34_618 ();
 sg13g2_decap_4 FILLER_34_625 ();
 sg13g2_fill_1 FILLER_34_629 ();
 sg13g2_fill_2 FILLER_34_654 ();
 sg13g2_fill_1 FILLER_34_656 ();
 sg13g2_decap_8 FILLER_34_661 ();
 sg13g2_decap_8 FILLER_34_668 ();
 sg13g2_decap_8 FILLER_34_675 ();
 sg13g2_decap_8 FILLER_34_682 ();
 sg13g2_fill_2 FILLER_34_689 ();
 sg13g2_fill_1 FILLER_34_691 ();
 sg13g2_decap_8 FILLER_34_696 ();
 sg13g2_decap_8 FILLER_34_703 ();
 sg13g2_decap_8 FILLER_34_710 ();
 sg13g2_decap_8 FILLER_34_717 ();
 sg13g2_decap_8 FILLER_34_724 ();
 sg13g2_decap_4 FILLER_34_731 ();
 sg13g2_decap_4 FILLER_34_742 ();
 sg13g2_decap_4 FILLER_34_754 ();
 sg13g2_fill_2 FILLER_34_758 ();
 sg13g2_decap_4 FILLER_34_768 ();
 sg13g2_fill_1 FILLER_34_772 ();
 sg13g2_decap_8 FILLER_34_808 ();
 sg13g2_fill_2 FILLER_34_815 ();
 sg13g2_fill_1 FILLER_34_817 ();
 sg13g2_decap_8 FILLER_34_847 ();
 sg13g2_decap_8 FILLER_34_854 ();
 sg13g2_decap_8 FILLER_34_861 ();
 sg13g2_fill_1 FILLER_34_868 ();
 sg13g2_fill_2 FILLER_34_874 ();
 sg13g2_fill_1 FILLER_34_876 ();
 sg13g2_fill_2 FILLER_34_883 ();
 sg13g2_fill_1 FILLER_34_885 ();
 sg13g2_fill_1 FILLER_34_890 ();
 sg13g2_fill_2 FILLER_34_900 ();
 sg13g2_fill_1 FILLER_34_902 ();
 sg13g2_fill_2 FILLER_34_908 ();
 sg13g2_fill_1 FILLER_34_925 ();
 sg13g2_decap_8 FILLER_34_929 ();
 sg13g2_decap_8 FILLER_34_952 ();
 sg13g2_fill_1 FILLER_34_959 ();
 sg13g2_decap_8 FILLER_34_965 ();
 sg13g2_decap_8 FILLER_34_976 ();
 sg13g2_fill_2 FILLER_34_983 ();
 sg13g2_fill_1 FILLER_34_985 ();
 sg13g2_decap_4 FILLER_34_990 ();
 sg13g2_fill_2 FILLER_34_994 ();
 sg13g2_decap_8 FILLER_34_1001 ();
 sg13g2_fill_2 FILLER_34_1008 ();
 sg13g2_decap_8 FILLER_34_1014 ();
 sg13g2_decap_8 FILLER_34_1021 ();
 sg13g2_decap_8 FILLER_34_1028 ();
 sg13g2_decap_8 FILLER_34_1040 ();
 sg13g2_decap_8 FILLER_34_1056 ();
 sg13g2_fill_2 FILLER_34_1063 ();
 sg13g2_fill_2 FILLER_34_1070 ();
 sg13g2_fill_1 FILLER_34_1072 ();
 sg13g2_fill_2 FILLER_34_1078 ();
 sg13g2_decap_8 FILLER_34_1086 ();
 sg13g2_decap_8 FILLER_34_1093 ();
 sg13g2_decap_4 FILLER_34_1100 ();
 sg13g2_fill_1 FILLER_34_1104 ();
 sg13g2_decap_8 FILLER_34_1114 ();
 sg13g2_decap_8 FILLER_34_1121 ();
 sg13g2_decap_8 FILLER_34_1128 ();
 sg13g2_decap_8 FILLER_34_1135 ();
 sg13g2_fill_1 FILLER_34_1142 ();
 sg13g2_decap_8 FILLER_34_1149 ();
 sg13g2_decap_8 FILLER_34_1156 ();
 sg13g2_decap_4 FILLER_34_1168 ();
 sg13g2_decap_8 FILLER_34_1177 ();
 sg13g2_fill_2 FILLER_34_1184 ();
 sg13g2_fill_1 FILLER_34_1186 ();
 sg13g2_decap_8 FILLER_34_1195 ();
 sg13g2_decap_8 FILLER_34_1202 ();
 sg13g2_fill_2 FILLER_34_1209 ();
 sg13g2_fill_1 FILLER_34_1225 ();
 sg13g2_fill_1 FILLER_34_1232 ();
 sg13g2_decap_8 FILLER_34_1238 ();
 sg13g2_decap_4 FILLER_34_1245 ();
 sg13g2_fill_2 FILLER_34_1249 ();
 sg13g2_fill_2 FILLER_34_1265 ();
 sg13g2_fill_1 FILLER_34_1267 ();
 sg13g2_fill_1 FILLER_34_1273 ();
 sg13g2_fill_2 FILLER_34_1279 ();
 sg13g2_fill_1 FILLER_34_1281 ();
 sg13g2_decap_8 FILLER_34_1286 ();
 sg13g2_decap_8 FILLER_34_1293 ();
 sg13g2_decap_8 FILLER_34_1300 ();
 sg13g2_decap_8 FILLER_34_1307 ();
 sg13g2_decap_8 FILLER_34_1314 ();
 sg13g2_decap_4 FILLER_34_1321 ();
 sg13g2_fill_1 FILLER_34_1325 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_fill_2 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_76 ();
 sg13g2_decap_8 FILLER_35_83 ();
 sg13g2_decap_8 FILLER_35_90 ();
 sg13g2_decap_8 FILLER_35_97 ();
 sg13g2_decap_8 FILLER_35_104 ();
 sg13g2_decap_8 FILLER_35_111 ();
 sg13g2_decap_8 FILLER_35_118 ();
 sg13g2_decap_4 FILLER_35_125 ();
 sg13g2_decap_8 FILLER_35_134 ();
 sg13g2_decap_8 FILLER_35_141 ();
 sg13g2_decap_8 FILLER_35_148 ();
 sg13g2_decap_8 FILLER_35_155 ();
 sg13g2_decap_8 FILLER_35_162 ();
 sg13g2_decap_8 FILLER_35_169 ();
 sg13g2_decap_8 FILLER_35_176 ();
 sg13g2_decap_8 FILLER_35_183 ();
 sg13g2_decap_8 FILLER_35_190 ();
 sg13g2_fill_2 FILLER_35_197 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_decap_8 FILLER_35_205 ();
 sg13g2_decap_8 FILLER_35_212 ();
 sg13g2_decap_8 FILLER_35_219 ();
 sg13g2_decap_8 FILLER_35_226 ();
 sg13g2_decap_8 FILLER_35_233 ();
 sg13g2_decap_8 FILLER_35_240 ();
 sg13g2_decap_8 FILLER_35_247 ();
 sg13g2_decap_8 FILLER_35_254 ();
 sg13g2_decap_8 FILLER_35_261 ();
 sg13g2_decap_8 FILLER_35_268 ();
 sg13g2_decap_8 FILLER_35_275 ();
 sg13g2_decap_8 FILLER_35_282 ();
 sg13g2_decap_8 FILLER_35_289 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_fill_2 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_345 ();
 sg13g2_decap_8 FILLER_35_352 ();
 sg13g2_decap_8 FILLER_35_359 ();
 sg13g2_decap_8 FILLER_35_366 ();
 sg13g2_decap_8 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_380 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_decap_8 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_35_415 ();
 sg13g2_decap_8 FILLER_35_422 ();
 sg13g2_decap_8 FILLER_35_429 ();
 sg13g2_decap_8 FILLER_35_436 ();
 sg13g2_decap_8 FILLER_35_443 ();
 sg13g2_decap_8 FILLER_35_450 ();
 sg13g2_decap_8 FILLER_35_457 ();
 sg13g2_decap_8 FILLER_35_464 ();
 sg13g2_decap_8 FILLER_35_471 ();
 sg13g2_decap_8 FILLER_35_478 ();
 sg13g2_decap_8 FILLER_35_485 ();
 sg13g2_fill_1 FILLER_35_492 ();
 sg13g2_decap_4 FILLER_35_498 ();
 sg13g2_fill_1 FILLER_35_502 ();
 sg13g2_decap_8 FILLER_35_507 ();
 sg13g2_decap_8 FILLER_35_514 ();
 sg13g2_fill_2 FILLER_35_521 ();
 sg13g2_fill_1 FILLER_35_523 ();
 sg13g2_decap_8 FILLER_35_529 ();
 sg13g2_decap_8 FILLER_35_536 ();
 sg13g2_decap_8 FILLER_35_543 ();
 sg13g2_decap_8 FILLER_35_550 ();
 sg13g2_decap_8 FILLER_35_557 ();
 sg13g2_decap_8 FILLER_35_564 ();
 sg13g2_decap_8 FILLER_35_571 ();
 sg13g2_decap_8 FILLER_35_578 ();
 sg13g2_fill_2 FILLER_35_585 ();
 sg13g2_fill_1 FILLER_35_587 ();
 sg13g2_fill_2 FILLER_35_618 ();
 sg13g2_fill_1 FILLER_35_620 ();
 sg13g2_decap_8 FILLER_35_626 ();
 sg13g2_decap_8 FILLER_35_633 ();
 sg13g2_fill_2 FILLER_35_640 ();
 sg13g2_fill_1 FILLER_35_642 ();
 sg13g2_decap_8 FILLER_35_647 ();
 sg13g2_fill_2 FILLER_35_654 ();
 sg13g2_fill_1 FILLER_35_656 ();
 sg13g2_decap_8 FILLER_35_664 ();
 sg13g2_decap_4 FILLER_35_671 ();
 sg13g2_fill_1 FILLER_35_675 ();
 sg13g2_decap_4 FILLER_35_685 ();
 sg13g2_fill_2 FILLER_35_689 ();
 sg13g2_decap_8 FILLER_35_696 ();
 sg13g2_decap_8 FILLER_35_703 ();
 sg13g2_decap_8 FILLER_35_710 ();
 sg13g2_decap_8 FILLER_35_717 ();
 sg13g2_decap_8 FILLER_35_724 ();
 sg13g2_decap_8 FILLER_35_731 ();
 sg13g2_decap_8 FILLER_35_738 ();
 sg13g2_decap_8 FILLER_35_745 ();
 sg13g2_decap_8 FILLER_35_752 ();
 sg13g2_decap_4 FILLER_35_759 ();
 sg13g2_decap_8 FILLER_35_767 ();
 sg13g2_decap_4 FILLER_35_774 ();
 sg13g2_decap_8 FILLER_35_797 ();
 sg13g2_decap_8 FILLER_35_804 ();
 sg13g2_decap_8 FILLER_35_811 ();
 sg13g2_decap_8 FILLER_35_818 ();
 sg13g2_decap_8 FILLER_35_825 ();
 sg13g2_decap_8 FILLER_35_832 ();
 sg13g2_decap_8 FILLER_35_839 ();
 sg13g2_decap_8 FILLER_35_846 ();
 sg13g2_decap_8 FILLER_35_853 ();
 sg13g2_fill_1 FILLER_35_860 ();
 sg13g2_decap_8 FILLER_35_865 ();
 sg13g2_decap_8 FILLER_35_872 ();
 sg13g2_decap_4 FILLER_35_879 ();
 sg13g2_fill_1 FILLER_35_883 ();
 sg13g2_decap_8 FILLER_35_892 ();
 sg13g2_fill_1 FILLER_35_917 ();
 sg13g2_fill_2 FILLER_35_923 ();
 sg13g2_fill_1 FILLER_35_925 ();
 sg13g2_decap_4 FILLER_35_943 ();
 sg13g2_decap_8 FILLER_35_952 ();
 sg13g2_decap_8 FILLER_35_959 ();
 sg13g2_fill_2 FILLER_35_966 ();
 sg13g2_fill_1 FILLER_35_968 ();
 sg13g2_decap_4 FILLER_35_977 ();
 sg13g2_decap_8 FILLER_35_989 ();
 sg13g2_decap_8 FILLER_35_996 ();
 sg13g2_decap_8 FILLER_35_1008 ();
 sg13g2_decap_8 FILLER_35_1015 ();
 sg13g2_decap_8 FILLER_35_1022 ();
 sg13g2_decap_8 FILLER_35_1029 ();
 sg13g2_decap_8 FILLER_35_1036 ();
 sg13g2_fill_2 FILLER_35_1043 ();
 sg13g2_decap_4 FILLER_35_1049 ();
 sg13g2_fill_1 FILLER_35_1053 ();
 sg13g2_decap_4 FILLER_35_1062 ();
 sg13g2_fill_1 FILLER_35_1066 ();
 sg13g2_decap_8 FILLER_35_1072 ();
 sg13g2_decap_4 FILLER_35_1079 ();
 sg13g2_fill_1 FILLER_35_1092 ();
 sg13g2_fill_1 FILLER_35_1103 ();
 sg13g2_decap_8 FILLER_35_1108 ();
 sg13g2_decap_8 FILLER_35_1115 ();
 sg13g2_decap_8 FILLER_35_1122 ();
 sg13g2_decap_8 FILLER_35_1129 ();
 sg13g2_decap_8 FILLER_35_1136 ();
 sg13g2_fill_2 FILLER_35_1143 ();
 sg13g2_fill_1 FILLER_35_1145 ();
 sg13g2_fill_1 FILLER_35_1153 ();
 sg13g2_decap_8 FILLER_35_1159 ();
 sg13g2_decap_4 FILLER_35_1166 ();
 sg13g2_decap_8 FILLER_35_1180 ();
 sg13g2_decap_8 FILLER_35_1187 ();
 sg13g2_decap_4 FILLER_35_1194 ();
 sg13g2_fill_2 FILLER_35_1198 ();
 sg13g2_decap_4 FILLER_35_1209 ();
 sg13g2_decap_4 FILLER_35_1218 ();
 sg13g2_fill_2 FILLER_35_1226 ();
 sg13g2_fill_2 FILLER_35_1238 ();
 sg13g2_fill_1 FILLER_35_1240 ();
 sg13g2_fill_2 FILLER_35_1246 ();
 sg13g2_decap_8 FILLER_35_1253 ();
 sg13g2_decap_8 FILLER_35_1260 ();
 sg13g2_fill_1 FILLER_35_1267 ();
 sg13g2_fill_1 FILLER_35_1273 ();
 sg13g2_decap_8 FILLER_35_1279 ();
 sg13g2_decap_8 FILLER_35_1286 ();
 sg13g2_decap_8 FILLER_35_1293 ();
 sg13g2_decap_8 FILLER_35_1300 ();
 sg13g2_decap_8 FILLER_35_1307 ();
 sg13g2_decap_8 FILLER_35_1314 ();
 sg13g2_decap_4 FILLER_35_1321 ();
 sg13g2_fill_1 FILLER_35_1325 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_44 ();
 sg13g2_decap_8 FILLER_36_50 ();
 sg13g2_decap_8 FILLER_36_57 ();
 sg13g2_fill_1 FILLER_36_64 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_109 ();
 sg13g2_decap_8 FILLER_36_116 ();
 sg13g2_fill_1 FILLER_36_123 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_154 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_fill_2 FILLER_36_191 ();
 sg13g2_decap_4 FILLER_36_198 ();
 sg13g2_decap_8 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_235 ();
 sg13g2_decap_8 FILLER_36_241 ();
 sg13g2_decap_8 FILLER_36_248 ();
 sg13g2_decap_8 FILLER_36_255 ();
 sg13g2_decap_8 FILLER_36_262 ();
 sg13g2_decap_8 FILLER_36_269 ();
 sg13g2_decap_8 FILLER_36_276 ();
 sg13g2_decap_8 FILLER_36_283 ();
 sg13g2_decap_8 FILLER_36_290 ();
 sg13g2_decap_8 FILLER_36_297 ();
 sg13g2_decap_8 FILLER_36_304 ();
 sg13g2_decap_8 FILLER_36_311 ();
 sg13g2_decap_8 FILLER_36_318 ();
 sg13g2_decap_8 FILLER_36_325 ();
 sg13g2_decap_8 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_339 ();
 sg13g2_decap_8 FILLER_36_346 ();
 sg13g2_decap_8 FILLER_36_353 ();
 sg13g2_decap_8 FILLER_36_360 ();
 sg13g2_decap_8 FILLER_36_367 ();
 sg13g2_decap_8 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_36_409 ();
 sg13g2_decap_4 FILLER_36_416 ();
 sg13g2_fill_1 FILLER_36_420 ();
 sg13g2_decap_8 FILLER_36_442 ();
 sg13g2_fill_2 FILLER_36_467 ();
 sg13g2_decap_8 FILLER_36_475 ();
 sg13g2_decap_4 FILLER_36_487 ();
 sg13g2_fill_1 FILLER_36_491 ();
 sg13g2_fill_1 FILLER_36_523 ();
 sg13g2_fill_2 FILLER_36_554 ();
 sg13g2_decap_8 FILLER_36_582 ();
 sg13g2_fill_2 FILLER_36_589 ();
 sg13g2_fill_1 FILLER_36_591 ();
 sg13g2_decap_8 FILLER_36_596 ();
 sg13g2_decap_4 FILLER_36_603 ();
 sg13g2_decap_8 FILLER_36_616 ();
 sg13g2_decap_8 FILLER_36_623 ();
 sg13g2_decap_8 FILLER_36_630 ();
 sg13g2_decap_8 FILLER_36_637 ();
 sg13g2_decap_8 FILLER_36_644 ();
 sg13g2_decap_8 FILLER_36_651 ();
 sg13g2_decap_8 FILLER_36_658 ();
 sg13g2_decap_8 FILLER_36_665 ();
 sg13g2_fill_1 FILLER_36_672 ();
 sg13g2_decap_4 FILLER_36_685 ();
 sg13g2_fill_2 FILLER_36_699 ();
 sg13g2_fill_1 FILLER_36_701 ();
 sg13g2_decap_8 FILLER_36_708 ();
 sg13g2_decap_8 FILLER_36_715 ();
 sg13g2_decap_8 FILLER_36_722 ();
 sg13g2_decap_8 FILLER_36_729 ();
 sg13g2_decap_8 FILLER_36_736 ();
 sg13g2_fill_2 FILLER_36_743 ();
 sg13g2_fill_1 FILLER_36_745 ();
 sg13g2_decap_8 FILLER_36_753 ();
 sg13g2_decap_8 FILLER_36_760 ();
 sg13g2_fill_1 FILLER_36_767 ();
 sg13g2_decap_8 FILLER_36_772 ();
 sg13g2_decap_8 FILLER_36_779 ();
 sg13g2_decap_8 FILLER_36_786 ();
 sg13g2_decap_8 FILLER_36_793 ();
 sg13g2_decap_8 FILLER_36_800 ();
 sg13g2_decap_8 FILLER_36_807 ();
 sg13g2_decap_8 FILLER_36_814 ();
 sg13g2_decap_8 FILLER_36_821 ();
 sg13g2_decap_8 FILLER_36_844 ();
 sg13g2_decap_8 FILLER_36_851 ();
 sg13g2_decap_8 FILLER_36_858 ();
 sg13g2_decap_8 FILLER_36_865 ();
 sg13g2_decap_8 FILLER_36_872 ();
 sg13g2_decap_8 FILLER_36_879 ();
 sg13g2_decap_8 FILLER_36_886 ();
 sg13g2_fill_2 FILLER_36_893 ();
 sg13g2_decap_4 FILLER_36_904 ();
 sg13g2_fill_1 FILLER_36_908 ();
 sg13g2_fill_1 FILLER_36_920 ();
 sg13g2_decap_8 FILLER_36_936 ();
 sg13g2_decap_4 FILLER_36_943 ();
 sg13g2_fill_1 FILLER_36_947 ();
 sg13g2_decap_8 FILLER_36_952 ();
 sg13g2_decap_8 FILLER_36_959 ();
 sg13g2_fill_2 FILLER_36_966 ();
 sg13g2_decap_8 FILLER_36_973 ();
 sg13g2_fill_2 FILLER_36_980 ();
 sg13g2_fill_1 FILLER_36_982 ();
 sg13g2_decap_8 FILLER_36_995 ();
 sg13g2_fill_1 FILLER_36_1002 ();
 sg13g2_decap_8 FILLER_36_1013 ();
 sg13g2_decap_4 FILLER_36_1020 ();
 sg13g2_decap_8 FILLER_36_1033 ();
 sg13g2_decap_8 FILLER_36_1040 ();
 sg13g2_fill_2 FILLER_36_1047 ();
 sg13g2_fill_1 FILLER_36_1049 ();
 sg13g2_decap_8 FILLER_36_1059 ();
 sg13g2_decap_8 FILLER_36_1066 ();
 sg13g2_decap_8 FILLER_36_1073 ();
 sg13g2_decap_8 FILLER_36_1080 ();
 sg13g2_decap_8 FILLER_36_1087 ();
 sg13g2_decap_8 FILLER_36_1094 ();
 sg13g2_fill_1 FILLER_36_1101 ();
 sg13g2_decap_8 FILLER_36_1106 ();
 sg13g2_fill_2 FILLER_36_1113 ();
 sg13g2_fill_1 FILLER_36_1115 ();
 sg13g2_decap_8 FILLER_36_1120 ();
 sg13g2_fill_1 FILLER_36_1127 ();
 sg13g2_fill_2 FILLER_36_1133 ();
 sg13g2_decap_4 FILLER_36_1140 ();
 sg13g2_fill_1 FILLER_36_1144 ();
 sg13g2_fill_2 FILLER_36_1150 ();
 sg13g2_decap_4 FILLER_36_1157 ();
 sg13g2_fill_1 FILLER_36_1161 ();
 sg13g2_decap_8 FILLER_36_1167 ();
 sg13g2_decap_8 FILLER_36_1174 ();
 sg13g2_fill_2 FILLER_36_1181 ();
 sg13g2_fill_1 FILLER_36_1183 ();
 sg13g2_decap_4 FILLER_36_1188 ();
 sg13g2_fill_1 FILLER_36_1192 ();
 sg13g2_decap_4 FILLER_36_1198 ();
 sg13g2_fill_1 FILLER_36_1202 ();
 sg13g2_decap_4 FILLER_36_1208 ();
 sg13g2_decap_4 FILLER_36_1217 ();
 sg13g2_fill_1 FILLER_36_1221 ();
 sg13g2_decap_8 FILLER_36_1231 ();
 sg13g2_decap_8 FILLER_36_1238 ();
 sg13g2_decap_8 FILLER_36_1245 ();
 sg13g2_decap_8 FILLER_36_1256 ();
 sg13g2_fill_2 FILLER_36_1267 ();
 sg13g2_fill_1 FILLER_36_1269 ();
 sg13g2_decap_8 FILLER_36_1280 ();
 sg13g2_decap_8 FILLER_36_1287 ();
 sg13g2_decap_8 FILLER_36_1294 ();
 sg13g2_decap_8 FILLER_36_1301 ();
 sg13g2_decap_8 FILLER_36_1308 ();
 sg13g2_decap_8 FILLER_36_1315 ();
 sg13g2_decap_4 FILLER_36_1322 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_18 ();
 sg13g2_decap_4 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_4 FILLER_37_91 ();
 sg13g2_fill_2 FILLER_37_95 ();
 sg13g2_fill_2 FILLER_37_149 ();
 sg13g2_fill_1 FILLER_37_151 ();
 sg13g2_decap_4 FILLER_37_204 ();
 sg13g2_fill_2 FILLER_37_208 ();
 sg13g2_fill_2 FILLER_37_214 ();
 sg13g2_decap_4 FILLER_37_221 ();
 sg13g2_decap_4 FILLER_37_229 ();
 sg13g2_fill_2 FILLER_37_233 ();
 sg13g2_decap_8 FILLER_37_240 ();
 sg13g2_decap_8 FILLER_37_247 ();
 sg13g2_decap_4 FILLER_37_254 ();
 sg13g2_decap_8 FILLER_37_263 ();
 sg13g2_decap_8 FILLER_37_270 ();
 sg13g2_decap_8 FILLER_37_277 ();
 sg13g2_fill_2 FILLER_37_284 ();
 sg13g2_decap_8 FILLER_37_291 ();
 sg13g2_decap_8 FILLER_37_303 ();
 sg13g2_decap_8 FILLER_37_310 ();
 sg13g2_decap_8 FILLER_37_317 ();
 sg13g2_decap_8 FILLER_37_324 ();
 sg13g2_decap_8 FILLER_37_331 ();
 sg13g2_fill_2 FILLER_37_338 ();
 sg13g2_fill_1 FILLER_37_340 ();
 sg13g2_decap_4 FILLER_37_351 ();
 sg13g2_fill_2 FILLER_37_355 ();
 sg13g2_decap_8 FILLER_37_361 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_4 FILLER_37_396 ();
 sg13g2_decap_8 FILLER_37_421 ();
 sg13g2_decap_8 FILLER_37_428 ();
 sg13g2_fill_1 FILLER_37_435 ();
 sg13g2_decap_8 FILLER_37_478 ();
 sg13g2_decap_4 FILLER_37_485 ();
 sg13g2_fill_1 FILLER_37_489 ();
 sg13g2_fill_1 FILLER_37_495 ();
 sg13g2_decap_8 FILLER_37_506 ();
 sg13g2_fill_1 FILLER_37_513 ();
 sg13g2_decap_8 FILLER_37_518 ();
 sg13g2_decap_8 FILLER_37_525 ();
 sg13g2_fill_1 FILLER_37_536 ();
 sg13g2_decap_8 FILLER_37_571 ();
 sg13g2_decap_8 FILLER_37_578 ();
 sg13g2_decap_8 FILLER_37_637 ();
 sg13g2_decap_8 FILLER_37_644 ();
 sg13g2_decap_4 FILLER_37_651 ();
 sg13g2_fill_2 FILLER_37_655 ();
 sg13g2_decap_4 FILLER_37_666 ();
 sg13g2_fill_1 FILLER_37_670 ();
 sg13g2_decap_4 FILLER_37_710 ();
 sg13g2_decap_8 FILLER_37_719 ();
 sg13g2_fill_1 FILLER_37_726 ();
 sg13g2_decap_8 FILLER_37_731 ();
 sg13g2_decap_8 FILLER_37_738 ();
 sg13g2_decap_8 FILLER_37_745 ();
 sg13g2_decap_8 FILLER_37_752 ();
 sg13g2_fill_2 FILLER_37_759 ();
 sg13g2_fill_1 FILLER_37_761 ();
 sg13g2_decap_8 FILLER_37_788 ();
 sg13g2_decap_8 FILLER_37_795 ();
 sg13g2_decap_8 FILLER_37_802 ();
 sg13g2_fill_1 FILLER_37_809 ();
 sg13g2_decap_8 FILLER_37_815 ();
 sg13g2_decap_8 FILLER_37_822 ();
 sg13g2_fill_2 FILLER_37_829 ();
 sg13g2_fill_1 FILLER_37_831 ();
 sg13g2_decap_8 FILLER_37_845 ();
 sg13g2_decap_8 FILLER_37_852 ();
 sg13g2_decap_8 FILLER_37_859 ();
 sg13g2_fill_2 FILLER_37_866 ();
 sg13g2_fill_1 FILLER_37_868 ();
 sg13g2_decap_8 FILLER_37_874 ();
 sg13g2_decap_8 FILLER_37_881 ();
 sg13g2_fill_2 FILLER_37_893 ();
 sg13g2_fill_1 FILLER_37_895 ();
 sg13g2_fill_2 FILLER_37_900 ();
 sg13g2_fill_1 FILLER_37_902 ();
 sg13g2_fill_2 FILLER_37_908 ();
 sg13g2_fill_2 FILLER_37_924 ();
 sg13g2_fill_1 FILLER_37_930 ();
 sg13g2_decap_8 FILLER_37_947 ();
 sg13g2_decap_8 FILLER_37_965 ();
 sg13g2_decap_4 FILLER_37_972 ();
 sg13g2_decap_8 FILLER_37_981 ();
 sg13g2_fill_2 FILLER_37_988 ();
 sg13g2_fill_1 FILLER_37_990 ();
 sg13g2_fill_1 FILLER_37_1011 ();
 sg13g2_fill_2 FILLER_37_1041 ();
 sg13g2_fill_1 FILLER_37_1048 ();
 sg13g2_decap_8 FILLER_37_1077 ();
 sg13g2_decap_4 FILLER_37_1084 ();
 sg13g2_fill_1 FILLER_37_1088 ();
 sg13g2_decap_4 FILLER_37_1094 ();
 sg13g2_decap_4 FILLER_37_1106 ();
 sg13g2_decap_4 FILLER_37_1114 ();
 sg13g2_fill_2 FILLER_37_1142 ();
 sg13g2_fill_1 FILLER_37_1144 ();
 sg13g2_fill_2 FILLER_37_1150 ();
 sg13g2_fill_1 FILLER_37_1152 ();
 sg13g2_decap_4 FILLER_37_1157 ();
 sg13g2_fill_1 FILLER_37_1161 ();
 sg13g2_decap_4 FILLER_37_1172 ();
 sg13g2_fill_2 FILLER_37_1176 ();
 sg13g2_fill_2 FILLER_37_1182 ();
 sg13g2_fill_1 FILLER_37_1184 ();
 sg13g2_decap_8 FILLER_37_1189 ();
 sg13g2_decap_4 FILLER_37_1196 ();
 sg13g2_decap_4 FILLER_37_1204 ();
 sg13g2_fill_2 FILLER_37_1218 ();
 sg13g2_fill_2 FILLER_37_1225 ();
 sg13g2_fill_2 FILLER_37_1237 ();
 sg13g2_decap_4 FILLER_37_1243 ();
 sg13g2_fill_1 FILLER_37_1247 ();
 sg13g2_decap_8 FILLER_37_1254 ();
 sg13g2_decap_4 FILLER_37_1261 ();
 sg13g2_fill_2 FILLER_37_1265 ();
 sg13g2_decap_8 FILLER_37_1281 ();
 sg13g2_decap_8 FILLER_37_1288 ();
 sg13g2_decap_8 FILLER_37_1295 ();
 sg13g2_decap_8 FILLER_37_1302 ();
 sg13g2_decap_8 FILLER_37_1309 ();
 sg13g2_decap_8 FILLER_37_1316 ();
 sg13g2_fill_2 FILLER_37_1323 ();
 sg13g2_fill_1 FILLER_37_1325 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_28 ();
 sg13g2_fill_1 FILLER_38_30 ();
 sg13g2_decap_4 FILLER_38_57 ();
 sg13g2_fill_1 FILLER_38_61 ();
 sg13g2_decap_8 FILLER_38_85 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_8 FILLER_38_99 ();
 sg13g2_decap_8 FILLER_38_106 ();
 sg13g2_decap_8 FILLER_38_113 ();
 sg13g2_decap_8 FILLER_38_120 ();
 sg13g2_decap_8 FILLER_38_127 ();
 sg13g2_decap_8 FILLER_38_134 ();
 sg13g2_fill_2 FILLER_38_141 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_fill_2 FILLER_38_152 ();
 sg13g2_decap_8 FILLER_38_159 ();
 sg13g2_decap_8 FILLER_38_166 ();
 sg13g2_decap_8 FILLER_38_173 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_191 ();
 sg13g2_decap_8 FILLER_38_198 ();
 sg13g2_fill_2 FILLER_38_205 ();
 sg13g2_fill_1 FILLER_38_207 ();
 sg13g2_decap_8 FILLER_38_242 ();
 sg13g2_fill_2 FILLER_38_249 ();
 sg13g2_fill_1 FILLER_38_251 ();
 sg13g2_decap_8 FILLER_38_261 ();
 sg13g2_decap_4 FILLER_38_268 ();
 sg13g2_fill_2 FILLER_38_272 ();
 sg13g2_decap_4 FILLER_38_279 ();
 sg13g2_fill_1 FILLER_38_283 ();
 sg13g2_decap_8 FILLER_38_288 ();
 sg13g2_decap_8 FILLER_38_295 ();
 sg13g2_decap_8 FILLER_38_302 ();
 sg13g2_decap_8 FILLER_38_309 ();
 sg13g2_decap_8 FILLER_38_316 ();
 sg13g2_decap_8 FILLER_38_323 ();
 sg13g2_decap_8 FILLER_38_330 ();
 sg13g2_decap_8 FILLER_38_337 ();
 sg13g2_decap_4 FILLER_38_344 ();
 sg13g2_fill_2 FILLER_38_348 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_fill_2 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_8 FILLER_38_404 ();
 sg13g2_decap_4 FILLER_38_411 ();
 sg13g2_decap_8 FILLER_38_436 ();
 sg13g2_decap_8 FILLER_38_443 ();
 sg13g2_decap_8 FILLER_38_450 ();
 sg13g2_decap_8 FILLER_38_457 ();
 sg13g2_decap_8 FILLER_38_464 ();
 sg13g2_decap_8 FILLER_38_471 ();
 sg13g2_fill_2 FILLER_38_478 ();
 sg13g2_decap_8 FILLER_38_492 ();
 sg13g2_decap_8 FILLER_38_499 ();
 sg13g2_decap_8 FILLER_38_506 ();
 sg13g2_decap_8 FILLER_38_513 ();
 sg13g2_decap_8 FILLER_38_520 ();
 sg13g2_decap_8 FILLER_38_527 ();
 sg13g2_decap_8 FILLER_38_534 ();
 sg13g2_decap_8 FILLER_38_541 ();
 sg13g2_decap_8 FILLER_38_548 ();
 sg13g2_decap_8 FILLER_38_555 ();
 sg13g2_decap_8 FILLER_38_562 ();
 sg13g2_decap_8 FILLER_38_569 ();
 sg13g2_decap_8 FILLER_38_576 ();
 sg13g2_fill_2 FILLER_38_583 ();
 sg13g2_fill_1 FILLER_38_585 ();
 sg13g2_fill_1 FILLER_38_591 ();
 sg13g2_decap_8 FILLER_38_596 ();
 sg13g2_decap_8 FILLER_38_603 ();
 sg13g2_decap_4 FILLER_38_610 ();
 sg13g2_fill_1 FILLER_38_614 ();
 sg13g2_fill_2 FILLER_38_623 ();
 sg13g2_fill_1 FILLER_38_651 ();
 sg13g2_decap_8 FILLER_38_682 ();
 sg13g2_decap_4 FILLER_38_693 ();
 sg13g2_fill_2 FILLER_38_697 ();
 sg13g2_fill_2 FILLER_38_719 ();
 sg13g2_decap_8 FILLER_38_747 ();
 sg13g2_decap_8 FILLER_38_754 ();
 sg13g2_decap_8 FILLER_38_761 ();
 sg13g2_decap_8 FILLER_38_768 ();
 sg13g2_decap_8 FILLER_38_775 ();
 sg13g2_decap_8 FILLER_38_782 ();
 sg13g2_decap_8 FILLER_38_789 ();
 sg13g2_decap_8 FILLER_38_796 ();
 sg13g2_decap_8 FILLER_38_803 ();
 sg13g2_decap_8 FILLER_38_810 ();
 sg13g2_fill_2 FILLER_38_817 ();
 sg13g2_fill_1 FILLER_38_819 ();
 sg13g2_decap_8 FILLER_38_824 ();
 sg13g2_decap_8 FILLER_38_831 ();
 sg13g2_decap_8 FILLER_38_838 ();
 sg13g2_decap_4 FILLER_38_849 ();
 sg13g2_fill_2 FILLER_38_853 ();
 sg13g2_decap_8 FILLER_38_859 ();
 sg13g2_fill_2 FILLER_38_866 ();
 sg13g2_fill_1 FILLER_38_868 ();
 sg13g2_decap_8 FILLER_38_872 ();
 sg13g2_fill_2 FILLER_38_884 ();
 sg13g2_fill_1 FILLER_38_902 ();
 sg13g2_decap_4 FILLER_38_910 ();
 sg13g2_fill_1 FILLER_38_914 ();
 sg13g2_fill_1 FILLER_38_927 ();
 sg13g2_decap_8 FILLER_38_934 ();
 sg13g2_decap_8 FILLER_38_945 ();
 sg13g2_decap_8 FILLER_38_952 ();
 sg13g2_fill_1 FILLER_38_959 ();
 sg13g2_decap_4 FILLER_38_978 ();
 sg13g2_decap_4 FILLER_38_986 ();
 sg13g2_fill_1 FILLER_38_990 ();
 sg13g2_fill_2 FILLER_38_1000 ();
 sg13g2_decap_8 FILLER_38_1019 ();
 sg13g2_fill_1 FILLER_38_1026 ();
 sg13g2_decap_8 FILLER_38_1031 ();
 sg13g2_decap_8 FILLER_38_1038 ();
 sg13g2_fill_1 FILLER_38_1045 ();
 sg13g2_decap_4 FILLER_38_1051 ();
 sg13g2_decap_8 FILLER_38_1060 ();
 sg13g2_decap_4 FILLER_38_1067 ();
 sg13g2_fill_2 FILLER_38_1071 ();
 sg13g2_decap_8 FILLER_38_1094 ();
 sg13g2_decap_8 FILLER_38_1101 ();
 sg13g2_decap_8 FILLER_38_1108 ();
 sg13g2_decap_8 FILLER_38_1115 ();
 sg13g2_decap_4 FILLER_38_1122 ();
 sg13g2_fill_1 FILLER_38_1126 ();
 sg13g2_fill_1 FILLER_38_1137 ();
 sg13g2_decap_4 FILLER_38_1143 ();
 sg13g2_fill_1 FILLER_38_1147 ();
 sg13g2_fill_1 FILLER_38_1175 ();
 sg13g2_decap_8 FILLER_38_1189 ();
 sg13g2_fill_2 FILLER_38_1196 ();
 sg13g2_fill_1 FILLER_38_1198 ();
 sg13g2_fill_2 FILLER_38_1204 ();
 sg13g2_decap_8 FILLER_38_1214 ();
 sg13g2_decap_8 FILLER_38_1221 ();
 sg13g2_fill_2 FILLER_38_1228 ();
 sg13g2_fill_1 FILLER_38_1230 ();
 sg13g2_decap_4 FILLER_38_1245 ();
 sg13g2_decap_4 FILLER_38_1254 ();
 sg13g2_fill_2 FILLER_38_1271 ();
 sg13g2_fill_2 FILLER_38_1283 ();
 sg13g2_fill_1 FILLER_38_1285 ();
 sg13g2_decap_8 FILLER_38_1291 ();
 sg13g2_decap_8 FILLER_38_1298 ();
 sg13g2_decap_8 FILLER_38_1305 ();
 sg13g2_decap_8 FILLER_38_1312 ();
 sg13g2_decap_8 FILLER_38_1319 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_fill_2 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_41 ();
 sg13g2_decap_8 FILLER_39_48 ();
 sg13g2_fill_1 FILLER_39_69 ();
 sg13g2_fill_1 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_104 ();
 sg13g2_decap_8 FILLER_39_111 ();
 sg13g2_decap_4 FILLER_39_118 ();
 sg13g2_fill_2 FILLER_39_122 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_4 FILLER_39_147 ();
 sg13g2_fill_2 FILLER_39_151 ();
 sg13g2_decap_8 FILLER_39_157 ();
 sg13g2_decap_8 FILLER_39_164 ();
 sg13g2_decap_8 FILLER_39_171 ();
 sg13g2_fill_2 FILLER_39_178 ();
 sg13g2_fill_1 FILLER_39_180 ();
 sg13g2_decap_8 FILLER_39_185 ();
 sg13g2_decap_4 FILLER_39_192 ();
 sg13g2_fill_2 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_202 ();
 sg13g2_decap_8 FILLER_39_209 ();
 sg13g2_decap_8 FILLER_39_216 ();
 sg13g2_decap_8 FILLER_39_223 ();
 sg13g2_decap_8 FILLER_39_230 ();
 sg13g2_decap_8 FILLER_39_237 ();
 sg13g2_decap_8 FILLER_39_244 ();
 sg13g2_decap_8 FILLER_39_303 ();
 sg13g2_fill_2 FILLER_39_310 ();
 sg13g2_fill_1 FILLER_39_312 ();
 sg13g2_decap_4 FILLER_39_317 ();
 sg13g2_fill_2 FILLER_39_321 ();
 sg13g2_fill_2 FILLER_39_336 ();
 sg13g2_decap_8 FILLER_39_373 ();
 sg13g2_decap_8 FILLER_39_380 ();
 sg13g2_decap_8 FILLER_39_387 ();
 sg13g2_decap_4 FILLER_39_394 ();
 sg13g2_fill_2 FILLER_39_398 ();
 sg13g2_decap_8 FILLER_39_421 ();
 sg13g2_decap_8 FILLER_39_428 ();
 sg13g2_decap_8 FILLER_39_435 ();
 sg13g2_decap_8 FILLER_39_442 ();
 sg13g2_decap_8 FILLER_39_449 ();
 sg13g2_decap_8 FILLER_39_456 ();
 sg13g2_decap_8 FILLER_39_463 ();
 sg13g2_decap_8 FILLER_39_470 ();
 sg13g2_decap_8 FILLER_39_483 ();
 sg13g2_decap_8 FILLER_39_490 ();
 sg13g2_fill_2 FILLER_39_497 ();
 sg13g2_fill_1 FILLER_39_499 ();
 sg13g2_decap_8 FILLER_39_505 ();
 sg13g2_fill_2 FILLER_39_512 ();
 sg13g2_fill_1 FILLER_39_514 ();
 sg13g2_fill_2 FILLER_39_520 ();
 sg13g2_decap_4 FILLER_39_526 ();
 sg13g2_decap_8 FILLER_39_542 ();
 sg13g2_decap_8 FILLER_39_549 ();
 sg13g2_decap_8 FILLER_39_556 ();
 sg13g2_decap_8 FILLER_39_563 ();
 sg13g2_decap_8 FILLER_39_570 ();
 sg13g2_decap_8 FILLER_39_577 ();
 sg13g2_decap_8 FILLER_39_584 ();
 sg13g2_fill_1 FILLER_39_591 ();
 sg13g2_decap_8 FILLER_39_595 ();
 sg13g2_decap_8 FILLER_39_602 ();
 sg13g2_fill_1 FILLER_39_609 ();
 sg13g2_decap_8 FILLER_39_640 ();
 sg13g2_decap_4 FILLER_39_647 ();
 sg13g2_fill_2 FILLER_39_651 ();
 sg13g2_fill_1 FILLER_39_658 ();
 sg13g2_decap_8 FILLER_39_663 ();
 sg13g2_decap_8 FILLER_39_670 ();
 sg13g2_decap_8 FILLER_39_677 ();
 sg13g2_decap_8 FILLER_39_684 ();
 sg13g2_decap_8 FILLER_39_691 ();
 sg13g2_decap_8 FILLER_39_698 ();
 sg13g2_fill_2 FILLER_39_722 ();
 sg13g2_decap_8 FILLER_39_754 ();
 sg13g2_decap_8 FILLER_39_761 ();
 sg13g2_decap_8 FILLER_39_768 ();
 sg13g2_decap_8 FILLER_39_775 ();
 sg13g2_decap_8 FILLER_39_782 ();
 sg13g2_decap_8 FILLER_39_789 ();
 sg13g2_decap_8 FILLER_39_796 ();
 sg13g2_decap_8 FILLER_39_803 ();
 sg13g2_decap_8 FILLER_39_810 ();
 sg13g2_decap_4 FILLER_39_817 ();
 sg13g2_decap_8 FILLER_39_852 ();
 sg13g2_fill_2 FILLER_39_871 ();
 sg13g2_decap_4 FILLER_39_883 ();
 sg13g2_decap_8 FILLER_39_894 ();
 sg13g2_decap_8 FILLER_39_901 ();
 sg13g2_decap_4 FILLER_39_908 ();
 sg13g2_fill_2 FILLER_39_912 ();
 sg13g2_fill_2 FILLER_39_925 ();
 sg13g2_fill_1 FILLER_39_927 ();
 sg13g2_decap_8 FILLER_39_933 ();
 sg13g2_fill_2 FILLER_39_940 ();
 sg13g2_fill_1 FILLER_39_942 ();
 sg13g2_decap_4 FILLER_39_948 ();
 sg13g2_fill_1 FILLER_39_961 ();
 sg13g2_decap_8 FILLER_39_972 ();
 sg13g2_fill_2 FILLER_39_979 ();
 sg13g2_decap_8 FILLER_39_986 ();
 sg13g2_decap_8 FILLER_39_1005 ();
 sg13g2_fill_2 FILLER_39_1012 ();
 sg13g2_fill_1 FILLER_39_1014 ();
 sg13g2_decap_8 FILLER_39_1029 ();
 sg13g2_decap_4 FILLER_39_1036 ();
 sg13g2_decap_8 FILLER_39_1044 ();
 sg13g2_decap_8 FILLER_39_1061 ();
 sg13g2_fill_2 FILLER_39_1068 ();
 sg13g2_fill_1 FILLER_39_1070 ();
 sg13g2_decap_4 FILLER_39_1075 ();
 sg13g2_decap_8 FILLER_39_1084 ();
 sg13g2_fill_2 FILLER_39_1091 ();
 sg13g2_decap_8 FILLER_39_1098 ();
 sg13g2_decap_8 FILLER_39_1105 ();
 sg13g2_decap_8 FILLER_39_1112 ();
 sg13g2_decap_8 FILLER_39_1119 ();
 sg13g2_decap_8 FILLER_39_1126 ();
 sg13g2_decap_8 FILLER_39_1133 ();
 sg13g2_decap_8 FILLER_39_1140 ();
 sg13g2_decap_8 FILLER_39_1147 ();
 sg13g2_fill_1 FILLER_39_1154 ();
 sg13g2_decap_8 FILLER_39_1160 ();
 sg13g2_decap_4 FILLER_39_1167 ();
 sg13g2_decap_4 FILLER_39_1176 ();
 sg13g2_fill_2 FILLER_39_1180 ();
 sg13g2_decap_8 FILLER_39_1187 ();
 sg13g2_decap_4 FILLER_39_1194 ();
 sg13g2_decap_8 FILLER_39_1202 ();
 sg13g2_fill_2 FILLER_39_1209 ();
 sg13g2_decap_4 FILLER_39_1215 ();
 sg13g2_decap_8 FILLER_39_1223 ();
 sg13g2_fill_2 FILLER_39_1230 ();
 sg13g2_decap_8 FILLER_39_1242 ();
 sg13g2_fill_2 FILLER_39_1249 ();
 sg13g2_fill_2 FILLER_39_1256 ();
 sg13g2_decap_4 FILLER_39_1273 ();
 sg13g2_decap_8 FILLER_39_1282 ();
 sg13g2_decap_8 FILLER_39_1289 ();
 sg13g2_decap_8 FILLER_39_1296 ();
 sg13g2_decap_8 FILLER_39_1303 ();
 sg13g2_decap_8 FILLER_39_1310 ();
 sg13g2_decap_8 FILLER_39_1317 ();
 sg13g2_fill_2 FILLER_39_1324 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_fill_2 FILLER_40_21 ();
 sg13g2_fill_1 FILLER_40_28 ();
 sg13g2_fill_1 FILLER_40_34 ();
 sg13g2_fill_1 FILLER_40_46 ();
 sg13g2_fill_2 FILLER_40_61 ();
 sg13g2_fill_1 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_82 ();
 sg13g2_fill_1 FILLER_40_89 ();
 sg13g2_decap_8 FILLER_40_100 ();
 sg13g2_fill_2 FILLER_40_107 ();
 sg13g2_decap_8 FILLER_40_113 ();
 sg13g2_decap_8 FILLER_40_120 ();
 sg13g2_decap_4 FILLER_40_127 ();
 sg13g2_decap_4 FILLER_40_146 ();
 sg13g2_fill_1 FILLER_40_150 ();
 sg13g2_decap_4 FILLER_40_156 ();
 sg13g2_fill_2 FILLER_40_165 ();
 sg13g2_fill_2 FILLER_40_172 ();
 sg13g2_decap_8 FILLER_40_187 ();
 sg13g2_decap_4 FILLER_40_194 ();
 sg13g2_fill_2 FILLER_40_198 ();
 sg13g2_fill_2 FILLER_40_218 ();
 sg13g2_fill_1 FILLER_40_220 ();
 sg13g2_decap_8 FILLER_40_225 ();
 sg13g2_decap_8 FILLER_40_232 ();
 sg13g2_decap_8 FILLER_40_239 ();
 sg13g2_decap_8 FILLER_40_246 ();
 sg13g2_decap_8 FILLER_40_253 ();
 sg13g2_fill_1 FILLER_40_265 ();
 sg13g2_decap_8 FILLER_40_275 ();
 sg13g2_decap_8 FILLER_40_282 ();
 sg13g2_decap_8 FILLER_40_289 ();
 sg13g2_fill_1 FILLER_40_296 ();
 sg13g2_decap_4 FILLER_40_300 ();
 sg13g2_fill_2 FILLER_40_304 ();
 sg13g2_fill_1 FILLER_40_332 ();
 sg13g2_decap_8 FILLER_40_389 ();
 sg13g2_decap_8 FILLER_40_396 ();
 sg13g2_decap_8 FILLER_40_403 ();
 sg13g2_decap_8 FILLER_40_410 ();
 sg13g2_decap_8 FILLER_40_417 ();
 sg13g2_decap_8 FILLER_40_424 ();
 sg13g2_decap_8 FILLER_40_431 ();
 sg13g2_decap_8 FILLER_40_438 ();
 sg13g2_decap_8 FILLER_40_445 ();
 sg13g2_decap_8 FILLER_40_452 ();
 sg13g2_decap_8 FILLER_40_459 ();
 sg13g2_decap_4 FILLER_40_466 ();
 sg13g2_decap_8 FILLER_40_507 ();
 sg13g2_fill_2 FILLER_40_514 ();
 sg13g2_decap_8 FILLER_40_542 ();
 sg13g2_decap_8 FILLER_40_549 ();
 sg13g2_fill_1 FILLER_40_556 ();
 sg13g2_fill_1 FILLER_40_604 ();
 sg13g2_decap_8 FILLER_40_610 ();
 sg13g2_decap_8 FILLER_40_617 ();
 sg13g2_decap_4 FILLER_40_624 ();
 sg13g2_decap_8 FILLER_40_631 ();
 sg13g2_decap_8 FILLER_40_638 ();
 sg13g2_decap_8 FILLER_40_645 ();
 sg13g2_decap_8 FILLER_40_652 ();
 sg13g2_decap_8 FILLER_40_659 ();
 sg13g2_decap_8 FILLER_40_666 ();
 sg13g2_decap_8 FILLER_40_673 ();
 sg13g2_decap_8 FILLER_40_680 ();
 sg13g2_decap_8 FILLER_40_687 ();
 sg13g2_decap_8 FILLER_40_694 ();
 sg13g2_decap_8 FILLER_40_701 ();
 sg13g2_decap_8 FILLER_40_708 ();
 sg13g2_decap_8 FILLER_40_715 ();
 sg13g2_decap_8 FILLER_40_722 ();
 sg13g2_fill_2 FILLER_40_729 ();
 sg13g2_fill_1 FILLER_40_731 ();
 sg13g2_fill_2 FILLER_40_736 ();
 sg13g2_decap_8 FILLER_40_742 ();
 sg13g2_decap_8 FILLER_40_749 ();
 sg13g2_decap_8 FILLER_40_756 ();
 sg13g2_decap_8 FILLER_40_763 ();
 sg13g2_decap_8 FILLER_40_770 ();
 sg13g2_decap_8 FILLER_40_777 ();
 sg13g2_decap_8 FILLER_40_784 ();
 sg13g2_decap_8 FILLER_40_791 ();
 sg13g2_decap_8 FILLER_40_798 ();
 sg13g2_decap_8 FILLER_40_805 ();
 sg13g2_fill_2 FILLER_40_812 ();
 sg13g2_decap_8 FILLER_40_817 ();
 sg13g2_decap_8 FILLER_40_824 ();
 sg13g2_decap_8 FILLER_40_831 ();
 sg13g2_decap_8 FILLER_40_838 ();
 sg13g2_decap_8 FILLER_40_845 ();
 sg13g2_decap_8 FILLER_40_852 ();
 sg13g2_decap_8 FILLER_40_859 ();
 sg13g2_decap_8 FILLER_40_866 ();
 sg13g2_decap_8 FILLER_40_873 ();
 sg13g2_decap_8 FILLER_40_880 ();
 sg13g2_decap_8 FILLER_40_887 ();
 sg13g2_decap_8 FILLER_40_894 ();
 sg13g2_decap_8 FILLER_40_901 ();
 sg13g2_decap_4 FILLER_40_908 ();
 sg13g2_fill_2 FILLER_40_912 ();
 sg13g2_decap_8 FILLER_40_932 ();
 sg13g2_decap_8 FILLER_40_939 ();
 sg13g2_decap_8 FILLER_40_946 ();
 sg13g2_decap_8 FILLER_40_953 ();
 sg13g2_decap_8 FILLER_40_960 ();
 sg13g2_decap_8 FILLER_40_967 ();
 sg13g2_fill_1 FILLER_40_992 ();
 sg13g2_decap_8 FILLER_40_997 ();
 sg13g2_decap_8 FILLER_40_1004 ();
 sg13g2_decap_8 FILLER_40_1011 ();
 sg13g2_fill_1 FILLER_40_1018 ();
 sg13g2_decap_8 FILLER_40_1023 ();
 sg13g2_decap_8 FILLER_40_1030 ();
 sg13g2_decap_8 FILLER_40_1037 ();
 sg13g2_decap_8 FILLER_40_1044 ();
 sg13g2_decap_8 FILLER_40_1051 ();
 sg13g2_decap_8 FILLER_40_1058 ();
 sg13g2_fill_1 FILLER_40_1065 ();
 sg13g2_decap_8 FILLER_40_1073 ();
 sg13g2_decap_8 FILLER_40_1080 ();
 sg13g2_decap_8 FILLER_40_1087 ();
 sg13g2_decap_8 FILLER_40_1099 ();
 sg13g2_decap_8 FILLER_40_1106 ();
 sg13g2_decap_8 FILLER_40_1113 ();
 sg13g2_decap_8 FILLER_40_1120 ();
 sg13g2_decap_8 FILLER_40_1132 ();
 sg13g2_decap_8 FILLER_40_1139 ();
 sg13g2_decap_8 FILLER_40_1146 ();
 sg13g2_decap_8 FILLER_40_1153 ();
 sg13g2_decap_4 FILLER_40_1160 ();
 sg13g2_fill_1 FILLER_40_1164 ();
 sg13g2_fill_2 FILLER_40_1171 ();
 sg13g2_fill_1 FILLER_40_1173 ();
 sg13g2_decap_8 FILLER_40_1178 ();
 sg13g2_fill_1 FILLER_40_1185 ();
 sg13g2_fill_1 FILLER_40_1190 ();
 sg13g2_decap_4 FILLER_40_1196 ();
 sg13g2_fill_2 FILLER_40_1200 ();
 sg13g2_decap_8 FILLER_40_1213 ();
 sg13g2_decap_4 FILLER_40_1220 ();
 sg13g2_fill_2 FILLER_40_1229 ();
 sg13g2_fill_1 FILLER_40_1231 ();
 sg13g2_fill_1 FILLER_40_1242 ();
 sg13g2_fill_2 FILLER_40_1247 ();
 sg13g2_fill_1 FILLER_40_1249 ();
 sg13g2_decap_4 FILLER_40_1254 ();
 sg13g2_fill_2 FILLER_40_1258 ();
 sg13g2_fill_1 FILLER_40_1265 ();
 sg13g2_fill_2 FILLER_40_1271 ();
 sg13g2_fill_1 FILLER_40_1273 ();
 sg13g2_decap_8 FILLER_40_1283 ();
 sg13g2_decap_8 FILLER_40_1290 ();
 sg13g2_decap_8 FILLER_40_1297 ();
 sg13g2_decap_8 FILLER_40_1304 ();
 sg13g2_decap_8 FILLER_40_1311 ();
 sg13g2_decap_8 FILLER_40_1318 ();
 sg13g2_fill_1 FILLER_40_1325 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_fill_1 FILLER_41_21 ();
 sg13g2_fill_1 FILLER_41_26 ();
 sg13g2_fill_2 FILLER_41_37 ();
 sg13g2_decap_4 FILLER_41_44 ();
 sg13g2_fill_1 FILLER_41_56 ();
 sg13g2_fill_2 FILLER_41_62 ();
 sg13g2_fill_1 FILLER_41_69 ();
 sg13g2_decap_4 FILLER_41_75 ();
 sg13g2_fill_1 FILLER_41_79 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_fill_1 FILLER_41_91 ();
 sg13g2_decap_4 FILLER_41_96 ();
 sg13g2_fill_2 FILLER_41_100 ();
 sg13g2_decap_8 FILLER_41_128 ();
 sg13g2_decap_8 FILLER_41_135 ();
 sg13g2_fill_1 FILLER_41_142 ();
 sg13g2_decap_8 FILLER_41_188 ();
 sg13g2_decap_4 FILLER_41_195 ();
 sg13g2_fill_1 FILLER_41_199 ();
 sg13g2_decap_4 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_239 ();
 sg13g2_decap_4 FILLER_41_246 ();
 sg13g2_fill_1 FILLER_41_269 ();
 sg13g2_decap_8 FILLER_41_281 ();
 sg13g2_decap_8 FILLER_41_288 ();
 sg13g2_decap_4 FILLER_41_295 ();
 sg13g2_fill_1 FILLER_41_311 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_4 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_331 ();
 sg13g2_decap_4 FILLER_41_338 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_fill_2 FILLER_41_399 ();
 sg13g2_fill_1 FILLER_41_401 ();
 sg13g2_fill_2 FILLER_41_423 ();
 sg13g2_decap_8 FILLER_41_452 ();
 sg13g2_decap_8 FILLER_41_459 ();
 sg13g2_decap_8 FILLER_41_466 ();
 sg13g2_decap_8 FILLER_41_473 ();
 sg13g2_decap_8 FILLER_41_480 ();
 sg13g2_decap_4 FILLER_41_487 ();
 sg13g2_fill_2 FILLER_41_496 ();
 sg13g2_fill_1 FILLER_41_498 ();
 sg13g2_decap_8 FILLER_41_503 ();
 sg13g2_decap_8 FILLER_41_510 ();
 sg13g2_decap_8 FILLER_41_517 ();
 sg13g2_decap_4 FILLER_41_524 ();
 sg13g2_fill_2 FILLER_41_528 ();
 sg13g2_decap_8 FILLER_41_534 ();
 sg13g2_decap_8 FILLER_41_541 ();
 sg13g2_decap_8 FILLER_41_548 ();
 sg13g2_decap_8 FILLER_41_555 ();
 sg13g2_decap_8 FILLER_41_562 ();
 sg13g2_decap_8 FILLER_41_573 ();
 sg13g2_fill_2 FILLER_41_580 ();
 sg13g2_fill_1 FILLER_41_582 ();
 sg13g2_decap_8 FILLER_41_600 ();
 sg13g2_decap_8 FILLER_41_607 ();
 sg13g2_fill_2 FILLER_41_614 ();
 sg13g2_decap_8 FILLER_41_620 ();
 sg13g2_fill_1 FILLER_41_627 ();
 sg13g2_decap_8 FILLER_41_632 ();
 sg13g2_decap_8 FILLER_41_639 ();
 sg13g2_decap_8 FILLER_41_646 ();
 sg13g2_decap_8 FILLER_41_653 ();
 sg13g2_decap_8 FILLER_41_660 ();
 sg13g2_decap_4 FILLER_41_667 ();
 sg13g2_fill_1 FILLER_41_671 ();
 sg13g2_decap_8 FILLER_41_680 ();
 sg13g2_decap_8 FILLER_41_687 ();
 sg13g2_decap_8 FILLER_41_694 ();
 sg13g2_decap_8 FILLER_41_701 ();
 sg13g2_decap_8 FILLER_41_708 ();
 sg13g2_decap_8 FILLER_41_715 ();
 sg13g2_decap_4 FILLER_41_722 ();
 sg13g2_fill_2 FILLER_41_726 ();
 sg13g2_decap_8 FILLER_41_736 ();
 sg13g2_decap_8 FILLER_41_743 ();
 sg13g2_decap_8 FILLER_41_750 ();
 sg13g2_decap_8 FILLER_41_757 ();
 sg13g2_decap_8 FILLER_41_764 ();
 sg13g2_fill_2 FILLER_41_771 ();
 sg13g2_decap_8 FILLER_41_781 ();
 sg13g2_decap_8 FILLER_41_788 ();
 sg13g2_decap_8 FILLER_41_795 ();
 sg13g2_decap_4 FILLER_41_802 ();
 sg13g2_fill_2 FILLER_41_806 ();
 sg13g2_decap_4 FILLER_41_834 ();
 sg13g2_fill_2 FILLER_41_838 ();
 sg13g2_decap_8 FILLER_41_845 ();
 sg13g2_decap_8 FILLER_41_852 ();
 sg13g2_decap_8 FILLER_41_859 ();
 sg13g2_decap_4 FILLER_41_866 ();
 sg13g2_fill_1 FILLER_41_870 ();
 sg13g2_decap_8 FILLER_41_875 ();
 sg13g2_fill_2 FILLER_41_882 ();
 sg13g2_decap_8 FILLER_41_888 ();
 sg13g2_decap_4 FILLER_41_895 ();
 sg13g2_fill_2 FILLER_41_899 ();
 sg13g2_decap_4 FILLER_41_905 ();
 sg13g2_decap_8 FILLER_41_913 ();
 sg13g2_decap_8 FILLER_41_920 ();
 sg13g2_decap_4 FILLER_41_927 ();
 sg13g2_fill_1 FILLER_41_931 ();
 sg13g2_decap_4 FILLER_41_948 ();
 sg13g2_fill_2 FILLER_41_956 ();
 sg13g2_fill_2 FILLER_41_963 ();
 sg13g2_decap_4 FILLER_41_969 ();
 sg13g2_fill_1 FILLER_41_973 ();
 sg13g2_decap_8 FILLER_41_979 ();
 sg13g2_decap_8 FILLER_41_986 ();
 sg13g2_decap_8 FILLER_41_993 ();
 sg13g2_decap_4 FILLER_41_1000 ();
 sg13g2_fill_2 FILLER_41_1009 ();
 sg13g2_fill_1 FILLER_41_1011 ();
 sg13g2_decap_4 FILLER_41_1024 ();
 sg13g2_fill_1 FILLER_41_1028 ();
 sg13g2_decap_8 FILLER_41_1034 ();
 sg13g2_decap_8 FILLER_41_1041 ();
 sg13g2_fill_2 FILLER_41_1048 ();
 sg13g2_fill_1 FILLER_41_1060 ();
 sg13g2_decap_8 FILLER_41_1065 ();
 sg13g2_decap_8 FILLER_41_1072 ();
 sg13g2_fill_1 FILLER_41_1079 ();
 sg13g2_fill_1 FILLER_41_1085 ();
 sg13g2_decap_4 FILLER_41_1091 ();
 sg13g2_fill_2 FILLER_41_1095 ();
 sg13g2_decap_8 FILLER_41_1104 ();
 sg13g2_decap_8 FILLER_41_1111 ();
 sg13g2_decap_4 FILLER_41_1118 ();
 sg13g2_fill_2 FILLER_41_1122 ();
 sg13g2_decap_8 FILLER_41_1137 ();
 sg13g2_decap_8 FILLER_41_1144 ();
 sg13g2_fill_1 FILLER_41_1151 ();
 sg13g2_fill_2 FILLER_41_1178 ();
 sg13g2_decap_8 FILLER_41_1184 ();
 sg13g2_decap_8 FILLER_41_1191 ();
 sg13g2_decap_8 FILLER_41_1198 ();
 sg13g2_decap_4 FILLER_41_1205 ();
 sg13g2_decap_8 FILLER_41_1217 ();
 sg13g2_decap_4 FILLER_41_1224 ();
 sg13g2_fill_2 FILLER_41_1228 ();
 sg13g2_fill_1 FILLER_41_1240 ();
 sg13g2_decap_4 FILLER_41_1255 ();
 sg13g2_decap_4 FILLER_41_1264 ();
 sg13g2_fill_1 FILLER_41_1268 ();
 sg13g2_decap_8 FILLER_41_1278 ();
 sg13g2_decap_8 FILLER_41_1285 ();
 sg13g2_decap_8 FILLER_41_1292 ();
 sg13g2_decap_8 FILLER_41_1299 ();
 sg13g2_decap_8 FILLER_41_1306 ();
 sg13g2_decap_8 FILLER_41_1313 ();
 sg13g2_decap_4 FILLER_41_1320 ();
 sg13g2_fill_2 FILLER_41_1324 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_fill_2 FILLER_42_21 ();
 sg13g2_decap_4 FILLER_42_33 ();
 sg13g2_decap_4 FILLER_42_44 ();
 sg13g2_fill_1 FILLER_42_48 ();
 sg13g2_decap_4 FILLER_42_57 ();
 sg13g2_fill_2 FILLER_42_61 ();
 sg13g2_decap_8 FILLER_42_68 ();
 sg13g2_decap_8 FILLER_42_75 ();
 sg13g2_decap_8 FILLER_42_82 ();
 sg13g2_decap_8 FILLER_42_89 ();
 sg13g2_decap_8 FILLER_42_96 ();
 sg13g2_decap_8 FILLER_42_103 ();
 sg13g2_decap_8 FILLER_42_118 ();
 sg13g2_decap_8 FILLER_42_125 ();
 sg13g2_decap_4 FILLER_42_132 ();
 sg13g2_decap_8 FILLER_42_141 ();
 sg13g2_decap_8 FILLER_42_148 ();
 sg13g2_fill_1 FILLER_42_155 ();
 sg13g2_decap_8 FILLER_42_166 ();
 sg13g2_decap_4 FILLER_42_173 ();
 sg13g2_fill_1 FILLER_42_177 ();
 sg13g2_fill_2 FILLER_42_188 ();
 sg13g2_fill_2 FILLER_42_193 ();
 sg13g2_fill_1 FILLER_42_195 ();
 sg13g2_fill_2 FILLER_42_203 ();
 sg13g2_fill_1 FILLER_42_210 ();
 sg13g2_fill_2 FILLER_42_220 ();
 sg13g2_fill_1 FILLER_42_222 ();
 sg13g2_decap_8 FILLER_42_228 ();
 sg13g2_decap_8 FILLER_42_235 ();
 sg13g2_decap_8 FILLER_42_242 ();
 sg13g2_decap_8 FILLER_42_249 ();
 sg13g2_decap_4 FILLER_42_256 ();
 sg13g2_decap_8 FILLER_42_270 ();
 sg13g2_decap_8 FILLER_42_277 ();
 sg13g2_decap_8 FILLER_42_284 ();
 sg13g2_decap_8 FILLER_42_291 ();
 sg13g2_decap_8 FILLER_42_298 ();
 sg13g2_decap_4 FILLER_42_305 ();
 sg13g2_fill_2 FILLER_42_309 ();
 sg13g2_fill_2 FILLER_42_317 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_fill_2 FILLER_42_329 ();
 sg13g2_fill_1 FILLER_42_331 ();
 sg13g2_fill_2 FILLER_42_358 ();
 sg13g2_fill_1 FILLER_42_360 ();
 sg13g2_decap_8 FILLER_42_366 ();
 sg13g2_decap_8 FILLER_42_373 ();
 sg13g2_decap_8 FILLER_42_380 ();
 sg13g2_decap_8 FILLER_42_387 ();
 sg13g2_decap_8 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_fill_2 FILLER_42_408 ();
 sg13g2_fill_1 FILLER_42_410 ();
 sg13g2_decap_8 FILLER_42_440 ();
 sg13g2_decap_8 FILLER_42_447 ();
 sg13g2_decap_8 FILLER_42_454 ();
 sg13g2_decap_8 FILLER_42_467 ();
 sg13g2_decap_8 FILLER_42_474 ();
 sg13g2_decap_8 FILLER_42_481 ();
 sg13g2_decap_4 FILLER_42_488 ();
 sg13g2_fill_1 FILLER_42_492 ();
 sg13g2_fill_1 FILLER_42_497 ();
 sg13g2_decap_8 FILLER_42_508 ();
 sg13g2_decap_8 FILLER_42_515 ();
 sg13g2_decap_8 FILLER_42_522 ();
 sg13g2_fill_2 FILLER_42_564 ();
 sg13g2_fill_1 FILLER_42_566 ();
 sg13g2_decap_8 FILLER_42_571 ();
 sg13g2_decap_4 FILLER_42_578 ();
 sg13g2_fill_1 FILLER_42_582 ();
 sg13g2_decap_8 FILLER_42_604 ();
 sg13g2_decap_8 FILLER_42_611 ();
 sg13g2_decap_4 FILLER_42_618 ();
 sg13g2_fill_1 FILLER_42_622 ();
 sg13g2_decap_8 FILLER_42_644 ();
 sg13g2_decap_8 FILLER_42_655 ();
 sg13g2_decap_8 FILLER_42_662 ();
 sg13g2_decap_8 FILLER_42_669 ();
 sg13g2_decap_4 FILLER_42_676 ();
 sg13g2_fill_1 FILLER_42_680 ();
 sg13g2_decap_8 FILLER_42_685 ();
 sg13g2_decap_4 FILLER_42_692 ();
 sg13g2_decap_8 FILLER_42_700 ();
 sg13g2_decap_4 FILLER_42_707 ();
 sg13g2_fill_1 FILLER_42_711 ();
 sg13g2_decap_8 FILLER_42_725 ();
 sg13g2_decap_8 FILLER_42_732 ();
 sg13g2_decap_8 FILLER_42_739 ();
 sg13g2_fill_2 FILLER_42_750 ();
 sg13g2_decap_8 FILLER_42_757 ();
 sg13g2_decap_8 FILLER_42_764 ();
 sg13g2_decap_8 FILLER_42_797 ();
 sg13g2_decap_8 FILLER_42_804 ();
 sg13g2_fill_1 FILLER_42_811 ();
 sg13g2_decap_8 FILLER_42_816 ();
 sg13g2_decap_8 FILLER_42_823 ();
 sg13g2_decap_8 FILLER_42_830 ();
 sg13g2_decap_4 FILLER_42_837 ();
 sg13g2_decap_8 FILLER_42_850 ();
 sg13g2_fill_1 FILLER_42_857 ();
 sg13g2_decap_8 FILLER_42_891 ();
 sg13g2_decap_8 FILLER_42_898 ();
 sg13g2_decap_4 FILLER_42_921 ();
 sg13g2_fill_2 FILLER_42_925 ();
 sg13g2_fill_1 FILLER_42_935 ();
 sg13g2_decap_8 FILLER_42_941 ();
 sg13g2_decap_8 FILLER_42_953 ();
 sg13g2_decap_4 FILLER_42_960 ();
 sg13g2_fill_1 FILLER_42_964 ();
 sg13g2_fill_2 FILLER_42_975 ();
 sg13g2_fill_2 FILLER_42_982 ();
 sg13g2_fill_1 FILLER_42_984 ();
 sg13g2_fill_2 FILLER_42_990 ();
 sg13g2_decap_8 FILLER_42_997 ();
 sg13g2_decap_8 FILLER_42_1004 ();
 sg13g2_decap_8 FILLER_42_1011 ();
 sg13g2_decap_8 FILLER_42_1018 ();
 sg13g2_fill_2 FILLER_42_1025 ();
 sg13g2_fill_1 FILLER_42_1027 ();
 sg13g2_decap_8 FILLER_42_1033 ();
 sg13g2_decap_8 FILLER_42_1040 ();
 sg13g2_decap_4 FILLER_42_1051 ();
 sg13g2_fill_1 FILLER_42_1055 ();
 sg13g2_decap_8 FILLER_42_1067 ();
 sg13g2_decap_4 FILLER_42_1074 ();
 sg13g2_decap_8 FILLER_42_1086 ();
 sg13g2_decap_4 FILLER_42_1093 ();
 sg13g2_fill_1 FILLER_42_1097 ();
 sg13g2_decap_4 FILLER_42_1115 ();
 sg13g2_fill_1 FILLER_42_1119 ();
 sg13g2_decap_8 FILLER_42_1132 ();
 sg13g2_decap_8 FILLER_42_1139 ();
 sg13g2_fill_1 FILLER_42_1146 ();
 sg13g2_fill_2 FILLER_42_1160 ();
 sg13g2_decap_4 FILLER_42_1166 ();
 sg13g2_fill_2 FILLER_42_1170 ();
 sg13g2_decap_8 FILLER_42_1177 ();
 sg13g2_decap_8 FILLER_42_1184 ();
 sg13g2_decap_8 FILLER_42_1191 ();
 sg13g2_decap_4 FILLER_42_1198 ();
 sg13g2_fill_1 FILLER_42_1202 ();
 sg13g2_decap_8 FILLER_42_1211 ();
 sg13g2_decap_8 FILLER_42_1218 ();
 sg13g2_fill_2 FILLER_42_1249 ();
 sg13g2_fill_1 FILLER_42_1266 ();
 sg13g2_fill_2 FILLER_42_1271 ();
 sg13g2_fill_1 FILLER_42_1283 ();
 sg13g2_decap_8 FILLER_42_1287 ();
 sg13g2_decap_8 FILLER_42_1294 ();
 sg13g2_decap_8 FILLER_42_1301 ();
 sg13g2_decap_8 FILLER_42_1308 ();
 sg13g2_decap_8 FILLER_42_1315 ();
 sg13g2_decap_4 FILLER_42_1322 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_4 FILLER_43_46 ();
 sg13g2_fill_1 FILLER_43_50 ();
 sg13g2_decap_8 FILLER_43_55 ();
 sg13g2_decap_8 FILLER_43_62 ();
 sg13g2_decap_8 FILLER_43_69 ();
 sg13g2_decap_8 FILLER_43_76 ();
 sg13g2_decap_8 FILLER_43_83 ();
 sg13g2_decap_8 FILLER_43_90 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_fill_1 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_166 ();
 sg13g2_decap_8 FILLER_43_173 ();
 sg13g2_fill_2 FILLER_43_180 ();
 sg13g2_decap_8 FILLER_43_186 ();
 sg13g2_decap_8 FILLER_43_193 ();
 sg13g2_decap_8 FILLER_43_200 ();
 sg13g2_decap_8 FILLER_43_207 ();
 sg13g2_decap_8 FILLER_43_214 ();
 sg13g2_decap_8 FILLER_43_221 ();
 sg13g2_decap_8 FILLER_43_228 ();
 sg13g2_decap_8 FILLER_43_235 ();
 sg13g2_decap_8 FILLER_43_242 ();
 sg13g2_decap_8 FILLER_43_249 ();
 sg13g2_decap_8 FILLER_43_256 ();
 sg13g2_decap_8 FILLER_43_263 ();
 sg13g2_decap_8 FILLER_43_270 ();
 sg13g2_decap_8 FILLER_43_277 ();
 sg13g2_decap_8 FILLER_43_284 ();
 sg13g2_decap_4 FILLER_43_291 ();
 sg13g2_fill_1 FILLER_43_295 ();
 sg13g2_decap_8 FILLER_43_330 ();
 sg13g2_fill_2 FILLER_43_337 ();
 sg13g2_fill_1 FILLER_43_339 ();
 sg13g2_decap_8 FILLER_43_344 ();
 sg13g2_decap_8 FILLER_43_351 ();
 sg13g2_decap_8 FILLER_43_358 ();
 sg13g2_decap_8 FILLER_43_365 ();
 sg13g2_decap_8 FILLER_43_372 ();
 sg13g2_decap_8 FILLER_43_379 ();
 sg13g2_decap_8 FILLER_43_407 ();
 sg13g2_decap_4 FILLER_43_414 ();
 sg13g2_fill_2 FILLER_43_418 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_8 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_455 ();
 sg13g2_decap_4 FILLER_43_462 ();
 sg13g2_decap_8 FILLER_43_472 ();
 sg13g2_decap_8 FILLER_43_479 ();
 sg13g2_decap_8 FILLER_43_486 ();
 sg13g2_decap_8 FILLER_43_493 ();
 sg13g2_decap_8 FILLER_43_500 ();
 sg13g2_decap_8 FILLER_43_507 ();
 sg13g2_decap_8 FILLER_43_514 ();
 sg13g2_decap_8 FILLER_43_521 ();
 sg13g2_decap_8 FILLER_43_528 ();
 sg13g2_decap_4 FILLER_43_535 ();
 sg13g2_decap_4 FILLER_43_544 ();
 sg13g2_fill_1 FILLER_43_548 ();
 sg13g2_fill_1 FILLER_43_553 ();
 sg13g2_decap_8 FILLER_43_584 ();
 sg13g2_fill_2 FILLER_43_591 ();
 sg13g2_fill_1 FILLER_43_593 ();
 sg13g2_decap_8 FILLER_43_599 ();
 sg13g2_decap_8 FILLER_43_606 ();
 sg13g2_decap_8 FILLER_43_613 ();
 sg13g2_decap_8 FILLER_43_620 ();
 sg13g2_decap_8 FILLER_43_627 ();
 sg13g2_decap_4 FILLER_43_639 ();
 sg13g2_fill_1 FILLER_43_643 ();
 sg13g2_fill_1 FILLER_43_680 ();
 sg13g2_decap_8 FILLER_43_741 ();
 sg13g2_decap_8 FILLER_43_748 ();
 sg13g2_fill_2 FILLER_43_755 ();
 sg13g2_fill_1 FILLER_43_757 ();
 sg13g2_decap_8 FILLER_43_762 ();
 sg13g2_decap_8 FILLER_43_769 ();
 sg13g2_decap_8 FILLER_43_776 ();
 sg13g2_decap_8 FILLER_43_783 ();
 sg13g2_decap_8 FILLER_43_790 ();
 sg13g2_decap_8 FILLER_43_797 ();
 sg13g2_fill_2 FILLER_43_804 ();
 sg13g2_fill_1 FILLER_43_806 ();
 sg13g2_decap_8 FILLER_43_811 ();
 sg13g2_decap_8 FILLER_43_818 ();
 sg13g2_decap_8 FILLER_43_825 ();
 sg13g2_decap_8 FILLER_43_832 ();
 sg13g2_decap_8 FILLER_43_839 ();
 sg13g2_decap_8 FILLER_43_846 ();
 sg13g2_decap_4 FILLER_43_853 ();
 sg13g2_fill_2 FILLER_43_861 ();
 sg13g2_fill_1 FILLER_43_867 ();
 sg13g2_fill_2 FILLER_43_888 ();
 sg13g2_fill_1 FILLER_43_890 ();
 sg13g2_decap_4 FILLER_43_897 ();
 sg13g2_fill_2 FILLER_43_910 ();
 sg13g2_fill_1 FILLER_43_920 ();
 sg13g2_decap_8 FILLER_43_930 ();
 sg13g2_fill_1 FILLER_43_937 ();
 sg13g2_decap_8 FILLER_43_943 ();
 sg13g2_decap_4 FILLER_43_950 ();
 sg13g2_fill_2 FILLER_43_954 ();
 sg13g2_fill_2 FILLER_43_971 ();
 sg13g2_decap_8 FILLER_43_978 ();
 sg13g2_decap_4 FILLER_43_990 ();
 sg13g2_fill_2 FILLER_43_999 ();
 sg13g2_decap_8 FILLER_43_1006 ();
 sg13g2_decap_8 FILLER_43_1013 ();
 sg13g2_decap_8 FILLER_43_1020 ();
 sg13g2_decap_8 FILLER_43_1036 ();
 sg13g2_decap_8 FILLER_43_1043 ();
 sg13g2_fill_1 FILLER_43_1050 ();
 sg13g2_decap_8 FILLER_43_1056 ();
 sg13g2_decap_8 FILLER_43_1063 ();
 sg13g2_fill_2 FILLER_43_1070 ();
 sg13g2_fill_1 FILLER_43_1072 ();
 sg13g2_decap_4 FILLER_43_1083 ();
 sg13g2_fill_1 FILLER_43_1087 ();
 sg13g2_decap_8 FILLER_43_1099 ();
 sg13g2_decap_8 FILLER_43_1106 ();
 sg13g2_decap_8 FILLER_43_1118 ();
 sg13g2_decap_8 FILLER_43_1125 ();
 sg13g2_decap_8 FILLER_43_1132 ();
 sg13g2_decap_4 FILLER_43_1139 ();
 sg13g2_fill_2 FILLER_43_1143 ();
 sg13g2_fill_1 FILLER_43_1164 ();
 sg13g2_decap_4 FILLER_43_1170 ();
 sg13g2_decap_8 FILLER_43_1179 ();
 sg13g2_fill_2 FILLER_43_1186 ();
 sg13g2_decap_4 FILLER_43_1198 ();
 sg13g2_fill_2 FILLER_43_1202 ();
 sg13g2_decap_4 FILLER_43_1208 ();
 sg13g2_fill_2 FILLER_43_1212 ();
 sg13g2_decap_8 FILLER_43_1219 ();
 sg13g2_fill_2 FILLER_43_1226 ();
 sg13g2_fill_2 FILLER_43_1240 ();
 sg13g2_fill_2 FILLER_43_1246 ();
 sg13g2_fill_1 FILLER_43_1248 ();
 sg13g2_decap_4 FILLER_43_1254 ();
 sg13g2_decap_8 FILLER_43_1263 ();
 sg13g2_decap_8 FILLER_43_1282 ();
 sg13g2_decap_8 FILLER_43_1289 ();
 sg13g2_decap_8 FILLER_43_1296 ();
 sg13g2_decap_8 FILLER_43_1303 ();
 sg13g2_decap_8 FILLER_43_1310 ();
 sg13g2_decap_8 FILLER_43_1317 ();
 sg13g2_fill_2 FILLER_43_1324 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_74 ();
 sg13g2_decap_8 FILLER_44_81 ();
 sg13g2_decap_8 FILLER_44_88 ();
 sg13g2_decap_8 FILLER_44_95 ();
 sg13g2_decap_4 FILLER_44_102 ();
 sg13g2_fill_1 FILLER_44_106 ();
 sg13g2_fill_1 FILLER_44_115 ();
 sg13g2_decap_8 FILLER_44_130 ();
 sg13g2_decap_8 FILLER_44_137 ();
 sg13g2_decap_8 FILLER_44_144 ();
 sg13g2_fill_2 FILLER_44_164 ();
 sg13g2_decap_8 FILLER_44_171 ();
 sg13g2_decap_8 FILLER_44_178 ();
 sg13g2_decap_8 FILLER_44_185 ();
 sg13g2_decap_8 FILLER_44_192 ();
 sg13g2_decap_8 FILLER_44_199 ();
 sg13g2_decap_8 FILLER_44_206 ();
 sg13g2_decap_8 FILLER_44_213 ();
 sg13g2_decap_8 FILLER_44_220 ();
 sg13g2_fill_1 FILLER_44_227 ();
 sg13g2_decap_8 FILLER_44_258 ();
 sg13g2_decap_8 FILLER_44_265 ();
 sg13g2_decap_8 FILLER_44_272 ();
 sg13g2_decap_8 FILLER_44_279 ();
 sg13g2_decap_8 FILLER_44_286 ();
 sg13g2_decap_8 FILLER_44_293 ();
 sg13g2_decap_8 FILLER_44_300 ();
 sg13g2_decap_8 FILLER_44_307 ();
 sg13g2_decap_8 FILLER_44_314 ();
 sg13g2_decap_4 FILLER_44_321 ();
 sg13g2_fill_1 FILLER_44_325 ();
 sg13g2_decap_8 FILLER_44_331 ();
 sg13g2_decap_8 FILLER_44_338 ();
 sg13g2_decap_8 FILLER_44_345 ();
 sg13g2_decap_8 FILLER_44_352 ();
 sg13g2_fill_2 FILLER_44_359 ();
 sg13g2_fill_1 FILLER_44_361 ();
 sg13g2_decap_8 FILLER_44_366 ();
 sg13g2_fill_2 FILLER_44_373 ();
 sg13g2_fill_1 FILLER_44_375 ();
 sg13g2_decap_8 FILLER_44_397 ();
 sg13g2_decap_4 FILLER_44_425 ();
 sg13g2_fill_1 FILLER_44_429 ();
 sg13g2_decap_8 FILLER_44_486 ();
 sg13g2_decap_4 FILLER_44_493 ();
 sg13g2_fill_1 FILLER_44_497 ();
 sg13g2_decap_8 FILLER_44_503 ();
 sg13g2_fill_2 FILLER_44_510 ();
 sg13g2_decap_8 FILLER_44_542 ();
 sg13g2_decap_4 FILLER_44_549 ();
 sg13g2_fill_1 FILLER_44_553 ();
 sg13g2_decap_8 FILLER_44_559 ();
 sg13g2_fill_1 FILLER_44_566 ();
 sg13g2_decap_8 FILLER_44_571 ();
 sg13g2_decap_8 FILLER_44_578 ();
 sg13g2_decap_8 FILLER_44_585 ();
 sg13g2_decap_8 FILLER_44_592 ();
 sg13g2_fill_1 FILLER_44_599 ();
 sg13g2_decap_8 FILLER_44_604 ();
 sg13g2_decap_8 FILLER_44_611 ();
 sg13g2_decap_8 FILLER_44_618 ();
 sg13g2_decap_8 FILLER_44_625 ();
 sg13g2_decap_8 FILLER_44_632 ();
 sg13g2_decap_8 FILLER_44_639 ();
 sg13g2_decap_8 FILLER_44_646 ();
 sg13g2_decap_8 FILLER_44_653 ();
 sg13g2_decap_8 FILLER_44_660 ();
 sg13g2_fill_1 FILLER_44_667 ();
 sg13g2_fill_1 FILLER_44_678 ();
 sg13g2_fill_2 FILLER_44_682 ();
 sg13g2_decap_4 FILLER_44_698 ();
 sg13g2_fill_1 FILLER_44_702 ();
 sg13g2_decap_4 FILLER_44_717 ();
 sg13g2_decap_8 FILLER_44_725 ();
 sg13g2_decap_8 FILLER_44_732 ();
 sg13g2_decap_8 FILLER_44_743 ();
 sg13g2_fill_1 FILLER_44_750 ();
 sg13g2_decap_8 FILLER_44_777 ();
 sg13g2_decap_8 FILLER_44_784 ();
 sg13g2_decap_8 FILLER_44_791 ();
 sg13g2_fill_2 FILLER_44_798 ();
 sg13g2_fill_1 FILLER_44_800 ();
 sg13g2_decap_8 FILLER_44_809 ();
 sg13g2_decap_8 FILLER_44_816 ();
 sg13g2_decap_8 FILLER_44_823 ();
 sg13g2_decap_8 FILLER_44_830 ();
 sg13g2_decap_8 FILLER_44_837 ();
 sg13g2_decap_8 FILLER_44_844 ();
 sg13g2_decap_4 FILLER_44_851 ();
 sg13g2_fill_2 FILLER_44_855 ();
 sg13g2_decap_8 FILLER_44_861 ();
 sg13g2_decap_4 FILLER_44_868 ();
 sg13g2_decap_8 FILLER_44_886 ();
 sg13g2_decap_8 FILLER_44_893 ();
 sg13g2_fill_1 FILLER_44_900 ();
 sg13g2_decap_4 FILLER_44_914 ();
 sg13g2_fill_1 FILLER_44_918 ();
 sg13g2_fill_2 FILLER_44_932 ();
 sg13g2_fill_2 FILLER_44_939 ();
 sg13g2_fill_1 FILLER_44_941 ();
 sg13g2_decap_8 FILLER_44_954 ();
 sg13g2_decap_8 FILLER_44_961 ();
 sg13g2_decap_4 FILLER_44_968 ();
 sg13g2_fill_1 FILLER_44_972 ();
 sg13g2_decap_4 FILLER_44_977 ();
 sg13g2_fill_2 FILLER_44_981 ();
 sg13g2_decap_4 FILLER_44_996 ();
 sg13g2_fill_2 FILLER_44_1010 ();
 sg13g2_fill_1 FILLER_44_1012 ();
 sg13g2_decap_4 FILLER_44_1023 ();
 sg13g2_decap_8 FILLER_44_1037 ();
 sg13g2_decap_8 FILLER_44_1044 ();
 sg13g2_fill_2 FILLER_44_1051 ();
 sg13g2_fill_1 FILLER_44_1053 ();
 sg13g2_decap_8 FILLER_44_1059 ();
 sg13g2_fill_2 FILLER_44_1078 ();
 sg13g2_decap_8 FILLER_44_1088 ();
 sg13g2_decap_8 FILLER_44_1095 ();
 sg13g2_decap_8 FILLER_44_1102 ();
 sg13g2_fill_2 FILLER_44_1109 ();
 sg13g2_decap_8 FILLER_44_1117 ();
 sg13g2_decap_4 FILLER_44_1124 ();
 sg13g2_fill_2 FILLER_44_1128 ();
 sg13g2_decap_8 FILLER_44_1135 ();
 sg13g2_decap_8 FILLER_44_1142 ();
 sg13g2_decap_4 FILLER_44_1149 ();
 sg13g2_fill_2 FILLER_44_1159 ();
 sg13g2_fill_1 FILLER_44_1161 ();
 sg13g2_fill_1 FILLER_44_1167 ();
 sg13g2_fill_2 FILLER_44_1172 ();
 sg13g2_fill_1 FILLER_44_1188 ();
 sg13g2_decap_4 FILLER_44_1194 ();
 sg13g2_decap_8 FILLER_44_1215 ();
 sg13g2_decap_4 FILLER_44_1222 ();
 sg13g2_fill_1 FILLER_44_1226 ();
 sg13g2_decap_8 FILLER_44_1232 ();
 sg13g2_decap_4 FILLER_44_1239 ();
 sg13g2_decap_4 FILLER_44_1252 ();
 sg13g2_fill_2 FILLER_44_1256 ();
 sg13g2_decap_8 FILLER_44_1273 ();
 sg13g2_decap_8 FILLER_44_1280 ();
 sg13g2_decap_8 FILLER_44_1287 ();
 sg13g2_decap_8 FILLER_44_1294 ();
 sg13g2_decap_8 FILLER_44_1301 ();
 sg13g2_decap_8 FILLER_44_1308 ();
 sg13g2_decap_8 FILLER_44_1315 ();
 sg13g2_decap_4 FILLER_44_1322 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_fill_2 FILLER_45_63 ();
 sg13g2_fill_2 FILLER_45_77 ();
 sg13g2_fill_2 FILLER_45_83 ();
 sg13g2_fill_1 FILLER_45_85 ();
 sg13g2_decap_8 FILLER_45_90 ();
 sg13g2_decap_8 FILLER_45_97 ();
 sg13g2_fill_2 FILLER_45_104 ();
 sg13g2_fill_1 FILLER_45_106 ();
 sg13g2_decap_8 FILLER_45_114 ();
 sg13g2_fill_2 FILLER_45_121 ();
 sg13g2_fill_1 FILLER_45_123 ();
 sg13g2_decap_8 FILLER_45_134 ();
 sg13g2_decap_8 FILLER_45_176 ();
 sg13g2_decap_8 FILLER_45_183 ();
 sg13g2_decap_8 FILLER_45_190 ();
 sg13g2_decap_8 FILLER_45_197 ();
 sg13g2_decap_8 FILLER_45_204 ();
 sg13g2_decap_8 FILLER_45_211 ();
 sg13g2_decap_8 FILLER_45_218 ();
 sg13g2_decap_8 FILLER_45_225 ();
 sg13g2_decap_8 FILLER_45_232 ();
 sg13g2_decap_8 FILLER_45_243 ();
 sg13g2_decap_8 FILLER_45_250 ();
 sg13g2_decap_8 FILLER_45_257 ();
 sg13g2_decap_8 FILLER_45_264 ();
 sg13g2_fill_2 FILLER_45_271 ();
 sg13g2_fill_1 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_278 ();
 sg13g2_fill_2 FILLER_45_285 ();
 sg13g2_fill_1 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_299 ();
 sg13g2_decap_8 FILLER_45_306 ();
 sg13g2_decap_8 FILLER_45_313 ();
 sg13g2_decap_4 FILLER_45_332 ();
 sg13g2_fill_2 FILLER_45_336 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_fill_1 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_414 ();
 sg13g2_fill_1 FILLER_45_421 ();
 sg13g2_decap_8 FILLER_45_443 ();
 sg13g2_decap_8 FILLER_45_450 ();
 sg13g2_decap_8 FILLER_45_457 ();
 sg13g2_decap_8 FILLER_45_464 ();
 sg13g2_decap_8 FILLER_45_471 ();
 sg13g2_decap_8 FILLER_45_478 ();
 sg13g2_decap_8 FILLER_45_485 ();
 sg13g2_decap_8 FILLER_45_492 ();
 sg13g2_fill_2 FILLER_45_499 ();
 sg13g2_decap_8 FILLER_45_506 ();
 sg13g2_fill_1 FILLER_45_513 ();
 sg13g2_decap_8 FILLER_45_523 ();
 sg13g2_fill_2 FILLER_45_530 ();
 sg13g2_decap_4 FILLER_45_553 ();
 sg13g2_fill_2 FILLER_45_557 ();
 sg13g2_decap_8 FILLER_45_563 ();
 sg13g2_decap_8 FILLER_45_570 ();
 sg13g2_decap_8 FILLER_45_577 ();
 sg13g2_decap_4 FILLER_45_587 ();
 sg13g2_fill_2 FILLER_45_591 ();
 sg13g2_decap_4 FILLER_45_597 ();
 sg13g2_decap_8 FILLER_45_627 ();
 sg13g2_decap_8 FILLER_45_634 ();
 sg13g2_decap_8 FILLER_45_641 ();
 sg13g2_decap_8 FILLER_45_648 ();
 sg13g2_decap_8 FILLER_45_655 ();
 sg13g2_decap_8 FILLER_45_662 ();
 sg13g2_fill_1 FILLER_45_669 ();
 sg13g2_fill_1 FILLER_45_686 ();
 sg13g2_decap_8 FILLER_45_697 ();
 sg13g2_decap_8 FILLER_45_704 ();
 sg13g2_fill_2 FILLER_45_711 ();
 sg13g2_fill_1 FILLER_45_713 ();
 sg13g2_decap_8 FILLER_45_718 ();
 sg13g2_decap_8 FILLER_45_725 ();
 sg13g2_decap_8 FILLER_45_732 ();
 sg13g2_decap_8 FILLER_45_739 ();
 sg13g2_fill_2 FILLER_45_746 ();
 sg13g2_fill_1 FILLER_45_748 ();
 sg13g2_decap_8 FILLER_45_753 ();
 sg13g2_decap_8 FILLER_45_760 ();
 sg13g2_decap_8 FILLER_45_767 ();
 sg13g2_decap_8 FILLER_45_774 ();
 sg13g2_decap_8 FILLER_45_781 ();
 sg13g2_decap_8 FILLER_45_788 ();
 sg13g2_decap_8 FILLER_45_795 ();
 sg13g2_decap_8 FILLER_45_802 ();
 sg13g2_decap_8 FILLER_45_809 ();
 sg13g2_decap_4 FILLER_45_816 ();
 sg13g2_decap_8 FILLER_45_846 ();
 sg13g2_decap_8 FILLER_45_853 ();
 sg13g2_decap_8 FILLER_45_860 ();
 sg13g2_decap_8 FILLER_45_867 ();
 sg13g2_decap_8 FILLER_45_874 ();
 sg13g2_decap_8 FILLER_45_881 ();
 sg13g2_decap_8 FILLER_45_888 ();
 sg13g2_decap_4 FILLER_45_895 ();
 sg13g2_decap_8 FILLER_45_908 ();
 sg13g2_fill_2 FILLER_45_915 ();
 sg13g2_fill_1 FILLER_45_917 ();
 sg13g2_decap_4 FILLER_45_928 ();
 sg13g2_decap_4 FILLER_45_937 ();
 sg13g2_decap_8 FILLER_45_946 ();
 sg13g2_decap_4 FILLER_45_953 ();
 sg13g2_fill_2 FILLER_45_970 ();
 sg13g2_fill_2 FILLER_45_987 ();
 sg13g2_decap_8 FILLER_45_995 ();
 sg13g2_fill_2 FILLER_45_1002 ();
 sg13g2_fill_1 FILLER_45_1004 ();
 sg13g2_decap_8 FILLER_45_1013 ();
 sg13g2_decap_8 FILLER_45_1020 ();
 sg13g2_decap_8 FILLER_45_1027 ();
 sg13g2_decap_8 FILLER_45_1034 ();
 sg13g2_decap_8 FILLER_45_1041 ();
 sg13g2_decap_8 FILLER_45_1048 ();
 sg13g2_fill_1 FILLER_45_1060 ();
 sg13g2_fill_1 FILLER_45_1069 ();
 sg13g2_fill_1 FILLER_45_1074 ();
 sg13g2_fill_1 FILLER_45_1080 ();
 sg13g2_decap_8 FILLER_45_1085 ();
 sg13g2_decap_8 FILLER_45_1092 ();
 sg13g2_fill_2 FILLER_45_1099 ();
 sg13g2_fill_2 FILLER_45_1111 ();
 sg13g2_fill_2 FILLER_45_1118 ();
 sg13g2_fill_1 FILLER_45_1120 ();
 sg13g2_fill_1 FILLER_45_1126 ();
 sg13g2_fill_2 FILLER_45_1133 ();
 sg13g2_fill_1 FILLER_45_1135 ();
 sg13g2_fill_2 FILLER_45_1141 ();
 sg13g2_decap_4 FILLER_45_1148 ();
 sg13g2_decap_4 FILLER_45_1157 ();
 sg13g2_fill_1 FILLER_45_1161 ();
 sg13g2_decap_8 FILLER_45_1167 ();
 sg13g2_fill_2 FILLER_45_1174 ();
 sg13g2_fill_1 FILLER_45_1176 ();
 sg13g2_decap_4 FILLER_45_1181 ();
 sg13g2_fill_2 FILLER_45_1185 ();
 sg13g2_decap_8 FILLER_45_1192 ();
 sg13g2_fill_1 FILLER_45_1199 ();
 sg13g2_fill_2 FILLER_45_1211 ();
 sg13g2_fill_1 FILLER_45_1218 ();
 sg13g2_decap_8 FILLER_45_1224 ();
 sg13g2_decap_8 FILLER_45_1231 ();
 sg13g2_decap_8 FILLER_45_1238 ();
 sg13g2_decap_4 FILLER_45_1245 ();
 sg13g2_fill_2 FILLER_45_1249 ();
 sg13g2_decap_4 FILLER_45_1256 ();
 sg13g2_fill_1 FILLER_45_1260 ();
 sg13g2_decap_4 FILLER_45_1265 ();
 sg13g2_decap_8 FILLER_45_1274 ();
 sg13g2_decap_8 FILLER_45_1281 ();
 sg13g2_decap_8 FILLER_45_1288 ();
 sg13g2_decap_8 FILLER_45_1295 ();
 sg13g2_decap_8 FILLER_45_1302 ();
 sg13g2_decap_8 FILLER_45_1309 ();
 sg13g2_decap_8 FILLER_45_1316 ();
 sg13g2_fill_2 FILLER_45_1323 ();
 sg13g2_fill_1 FILLER_45_1325 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_fill_2 FILLER_46_28 ();
 sg13g2_decap_4 FILLER_46_37 ();
 sg13g2_fill_1 FILLER_46_41 ();
 sg13g2_fill_2 FILLER_46_56 ();
 sg13g2_fill_2 FILLER_46_94 ();
 sg13g2_decap_8 FILLER_46_101 ();
 sg13g2_fill_2 FILLER_46_108 ();
 sg13g2_decap_8 FILLER_46_116 ();
 sg13g2_decap_8 FILLER_46_123 ();
 sg13g2_decap_8 FILLER_46_130 ();
 sg13g2_decap_8 FILLER_46_137 ();
 sg13g2_decap_8 FILLER_46_144 ();
 sg13g2_decap_4 FILLER_46_151 ();
 sg13g2_fill_1 FILLER_46_160 ();
 sg13g2_decap_8 FILLER_46_166 ();
 sg13g2_decap_8 FILLER_46_173 ();
 sg13g2_decap_4 FILLER_46_180 ();
 sg13g2_fill_2 FILLER_46_184 ();
 sg13g2_decap_8 FILLER_46_216 ();
 sg13g2_decap_8 FILLER_46_223 ();
 sg13g2_decap_8 FILLER_46_230 ();
 sg13g2_fill_2 FILLER_46_237 ();
 sg13g2_fill_1 FILLER_46_239 ();
 sg13g2_fill_2 FILLER_46_250 ();
 sg13g2_decap_8 FILLER_46_302 ();
 sg13g2_decap_8 FILLER_46_309 ();
 sg13g2_decap_8 FILLER_46_316 ();
 sg13g2_decap_4 FILLER_46_323 ();
 sg13g2_fill_2 FILLER_46_327 ();
 sg13g2_decap_8 FILLER_46_355 ();
 sg13g2_decap_8 FILLER_46_362 ();
 sg13g2_decap_8 FILLER_46_369 ();
 sg13g2_decap_8 FILLER_46_376 ();
 sg13g2_decap_8 FILLER_46_383 ();
 sg13g2_decap_8 FILLER_46_390 ();
 sg13g2_decap_8 FILLER_46_397 ();
 sg13g2_decap_8 FILLER_46_404 ();
 sg13g2_decap_8 FILLER_46_411 ();
 sg13g2_decap_8 FILLER_46_418 ();
 sg13g2_decap_4 FILLER_46_425 ();
 sg13g2_fill_2 FILLER_46_429 ();
 sg13g2_decap_8 FILLER_46_439 ();
 sg13g2_decap_8 FILLER_46_446 ();
 sg13g2_decap_8 FILLER_46_453 ();
 sg13g2_decap_8 FILLER_46_460 ();
 sg13g2_decap_8 FILLER_46_467 ();
 sg13g2_decap_8 FILLER_46_474 ();
 sg13g2_decap_8 FILLER_46_481 ();
 sg13g2_fill_1 FILLER_46_488 ();
 sg13g2_fill_1 FILLER_46_499 ();
 sg13g2_decap_4 FILLER_46_510 ();
 sg13g2_decap_8 FILLER_46_518 ();
 sg13g2_decap_4 FILLER_46_525 ();
 sg13g2_decap_4 FILLER_46_533 ();
 sg13g2_decap_8 FILLER_46_541 ();
 sg13g2_decap_8 FILLER_46_548 ();
 sg13g2_decap_8 FILLER_46_586 ();
 sg13g2_fill_2 FILLER_46_593 ();
 sg13g2_decap_8 FILLER_46_600 ();
 sg13g2_decap_8 FILLER_46_611 ();
 sg13g2_decap_8 FILLER_46_618 ();
 sg13g2_decap_8 FILLER_46_625 ();
 sg13g2_decap_8 FILLER_46_632 ();
 sg13g2_decap_8 FILLER_46_639 ();
 sg13g2_decap_4 FILLER_46_646 ();
 sg13g2_fill_1 FILLER_46_660 ();
 sg13g2_decap_4 FILLER_46_665 ();
 sg13g2_fill_2 FILLER_46_682 ();
 sg13g2_fill_2 FILLER_46_693 ();
 sg13g2_fill_1 FILLER_46_695 ();
 sg13g2_fill_2 FILLER_46_699 ();
 sg13g2_fill_1 FILLER_46_701 ();
 sg13g2_decap_8 FILLER_46_716 ();
 sg13g2_decap_8 FILLER_46_723 ();
 sg13g2_fill_1 FILLER_46_730 ();
 sg13g2_decap_8 FILLER_46_735 ();
 sg13g2_decap_8 FILLER_46_768 ();
 sg13g2_decap_8 FILLER_46_775 ();
 sg13g2_decap_4 FILLER_46_782 ();
 sg13g2_fill_1 FILLER_46_786 ();
 sg13g2_decap_8 FILLER_46_795 ();
 sg13g2_decap_8 FILLER_46_802 ();
 sg13g2_decap_8 FILLER_46_809 ();
 sg13g2_fill_2 FILLER_46_816 ();
 sg13g2_decap_4 FILLER_46_822 ();
 sg13g2_fill_1 FILLER_46_826 ();
 sg13g2_decap_8 FILLER_46_831 ();
 sg13g2_decap_8 FILLER_46_838 ();
 sg13g2_decap_8 FILLER_46_845 ();
 sg13g2_decap_8 FILLER_46_852 ();
 sg13g2_decap_8 FILLER_46_859 ();
 sg13g2_decap_8 FILLER_46_866 ();
 sg13g2_decap_8 FILLER_46_873 ();
 sg13g2_decap_4 FILLER_46_880 ();
 sg13g2_fill_1 FILLER_46_884 ();
 sg13g2_decap_8 FILLER_46_905 ();
 sg13g2_decap_8 FILLER_46_912 ();
 sg13g2_decap_8 FILLER_46_919 ();
 sg13g2_decap_4 FILLER_46_926 ();
 sg13g2_fill_2 FILLER_46_930 ();
 sg13g2_fill_2 FILLER_46_947 ();
 sg13g2_fill_1 FILLER_46_949 ();
 sg13g2_decap_8 FILLER_46_988 ();
 sg13g2_decap_8 FILLER_46_995 ();
 sg13g2_decap_8 FILLER_46_1002 ();
 sg13g2_decap_8 FILLER_46_1009 ();
 sg13g2_decap_8 FILLER_46_1016 ();
 sg13g2_fill_2 FILLER_46_1023 ();
 sg13g2_decap_8 FILLER_46_1030 ();
 sg13g2_decap_8 FILLER_46_1037 ();
 sg13g2_decap_8 FILLER_46_1044 ();
 sg13g2_decap_4 FILLER_46_1051 ();
 sg13g2_fill_2 FILLER_46_1055 ();
 sg13g2_decap_8 FILLER_46_1061 ();
 sg13g2_decap_8 FILLER_46_1068 ();
 sg13g2_fill_1 FILLER_46_1075 ();
 sg13g2_decap_4 FILLER_46_1080 ();
 sg13g2_decap_4 FILLER_46_1089 ();
 sg13g2_fill_2 FILLER_46_1093 ();
 sg13g2_fill_1 FILLER_46_1139 ();
 sg13g2_decap_4 FILLER_46_1144 ();
 sg13g2_fill_1 FILLER_46_1148 ();
 sg13g2_decap_8 FILLER_46_1153 ();
 sg13g2_fill_2 FILLER_46_1160 ();
 sg13g2_fill_1 FILLER_46_1162 ();
 sg13g2_decap_8 FILLER_46_1167 ();
 sg13g2_decap_4 FILLER_46_1174 ();
 sg13g2_decap_8 FILLER_46_1186 ();
 sg13g2_decap_8 FILLER_46_1193 ();
 sg13g2_decap_4 FILLER_46_1200 ();
 sg13g2_decap_8 FILLER_46_1209 ();
 sg13g2_decap_8 FILLER_46_1216 ();
 sg13g2_decap_8 FILLER_46_1223 ();
 sg13g2_decap_8 FILLER_46_1230 ();
 sg13g2_decap_8 FILLER_46_1237 ();
 sg13g2_decap_8 FILLER_46_1244 ();
 sg13g2_fill_1 FILLER_46_1251 ();
 sg13g2_decap_8 FILLER_46_1262 ();
 sg13g2_fill_1 FILLER_46_1269 ();
 sg13g2_decap_8 FILLER_46_1276 ();
 sg13g2_decap_8 FILLER_46_1283 ();
 sg13g2_decap_8 FILLER_46_1290 ();
 sg13g2_decap_8 FILLER_46_1297 ();
 sg13g2_decap_8 FILLER_46_1304 ();
 sg13g2_decap_8 FILLER_46_1311 ();
 sg13g2_decap_8 FILLER_46_1318 ();
 sg13g2_fill_1 FILLER_46_1325 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_fill_2 FILLER_47_35 ();
 sg13g2_decap_4 FILLER_47_49 ();
 sg13g2_fill_2 FILLER_47_53 ();
 sg13g2_fill_1 FILLER_47_70 ();
 sg13g2_fill_1 FILLER_47_79 ();
 sg13g2_decap_8 FILLER_47_87 ();
 sg13g2_decap_8 FILLER_47_94 ();
 sg13g2_decap_8 FILLER_47_101 ();
 sg13g2_fill_2 FILLER_47_108 ();
 sg13g2_decap_8 FILLER_47_123 ();
 sg13g2_decap_8 FILLER_47_130 ();
 sg13g2_decap_8 FILLER_47_137 ();
 sg13g2_decap_8 FILLER_47_144 ();
 sg13g2_fill_2 FILLER_47_151 ();
 sg13g2_decap_8 FILLER_47_166 ();
 sg13g2_decap_8 FILLER_47_173 ();
 sg13g2_fill_2 FILLER_47_180 ();
 sg13g2_fill_1 FILLER_47_182 ();
 sg13g2_decap_4 FILLER_47_187 ();
 sg13g2_fill_2 FILLER_47_191 ();
 sg13g2_decap_4 FILLER_47_203 ();
 sg13g2_fill_1 FILLER_47_207 ();
 sg13g2_decap_8 FILLER_47_211 ();
 sg13g2_decap_8 FILLER_47_218 ();
 sg13g2_decap_4 FILLER_47_225 ();
 sg13g2_decap_4 FILLER_47_260 ();
 sg13g2_fill_1 FILLER_47_264 ();
 sg13g2_fill_2 FILLER_47_291 ();
 sg13g2_fill_1 FILLER_47_293 ();
 sg13g2_decap_8 FILLER_47_299 ();
 sg13g2_fill_1 FILLER_47_306 ();
 sg13g2_fill_1 FILLER_47_316 ();
 sg13g2_decap_8 FILLER_47_356 ();
 sg13g2_fill_1 FILLER_47_363 ();
 sg13g2_decap_8 FILLER_47_368 ();
 sg13g2_decap_8 FILLER_47_375 ();
 sg13g2_decap_4 FILLER_47_382 ();
 sg13g2_fill_2 FILLER_47_386 ();
 sg13g2_fill_1 FILLER_47_394 ();
 sg13g2_decap_8 FILLER_47_401 ();
 sg13g2_decap_8 FILLER_47_408 ();
 sg13g2_decap_4 FILLER_47_415 ();
 sg13g2_fill_2 FILLER_47_419 ();
 sg13g2_decap_8 FILLER_47_442 ();
 sg13g2_decap_8 FILLER_47_449 ();
 sg13g2_decap_8 FILLER_47_456 ();
 sg13g2_decap_8 FILLER_47_463 ();
 sg13g2_decap_8 FILLER_47_470 ();
 sg13g2_decap_8 FILLER_47_477 ();
 sg13g2_decap_4 FILLER_47_484 ();
 sg13g2_fill_1 FILLER_47_488 ();
 sg13g2_decap_4 FILLER_47_515 ();
 sg13g2_decap_4 FILLER_47_529 ();
 sg13g2_fill_2 FILLER_47_533 ();
 sg13g2_decap_4 FILLER_47_539 ();
 sg13g2_fill_2 FILLER_47_543 ();
 sg13g2_decap_8 FILLER_47_549 ();
 sg13g2_decap_8 FILLER_47_556 ();
 sg13g2_fill_2 FILLER_47_563 ();
 sg13g2_decap_8 FILLER_47_577 ();
 sg13g2_decap_8 FILLER_47_584 ();
 sg13g2_fill_1 FILLER_47_591 ();
 sg13g2_decap_4 FILLER_47_597 ();
 sg13g2_fill_1 FILLER_47_601 ();
 sg13g2_decap_8 FILLER_47_609 ();
 sg13g2_decap_8 FILLER_47_616 ();
 sg13g2_decap_8 FILLER_47_623 ();
 sg13g2_decap_8 FILLER_47_630 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_decap_8 FILLER_47_644 ();
 sg13g2_decap_4 FILLER_47_677 ();
 sg13g2_fill_1 FILLER_47_681 ();
 sg13g2_decap_8 FILLER_47_686 ();
 sg13g2_decap_4 FILLER_47_693 ();
 sg13g2_fill_2 FILLER_47_697 ();
 sg13g2_fill_2 FILLER_47_717 ();
 sg13g2_fill_1 FILLER_47_722 ();
 sg13g2_decap_8 FILLER_47_749 ();
 sg13g2_decap_8 FILLER_47_756 ();
 sg13g2_decap_8 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_decap_8 FILLER_47_777 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_823 ();
 sg13g2_decap_8 FILLER_47_830 ();
 sg13g2_decap_8 FILLER_47_837 ();
 sg13g2_decap_8 FILLER_47_844 ();
 sg13g2_decap_8 FILLER_47_851 ();
 sg13g2_fill_2 FILLER_47_858 ();
 sg13g2_fill_1 FILLER_47_860 ();
 sg13g2_decap_8 FILLER_47_866 ();
 sg13g2_decap_8 FILLER_47_873 ();
 sg13g2_fill_1 FILLER_47_880 ();
 sg13g2_decap_8 FILLER_47_894 ();
 sg13g2_fill_1 FILLER_47_901 ();
 sg13g2_decap_8 FILLER_47_906 ();
 sg13g2_decap_4 FILLER_47_919 ();
 sg13g2_fill_2 FILLER_47_923 ();
 sg13g2_decap_8 FILLER_47_929 ();
 sg13g2_decap_8 FILLER_47_936 ();
 sg13g2_fill_2 FILLER_47_943 ();
 sg13g2_decap_8 FILLER_47_951 ();
 sg13g2_fill_1 FILLER_47_958 ();
 sg13g2_decap_8 FILLER_47_972 ();
 sg13g2_fill_1 FILLER_47_979 ();
 sg13g2_decap_4 FILLER_47_985 ();
 sg13g2_fill_2 FILLER_47_989 ();
 sg13g2_decap_8 FILLER_47_996 ();
 sg13g2_decap_8 FILLER_47_1003 ();
 sg13g2_fill_2 FILLER_47_1010 ();
 sg13g2_fill_1 FILLER_47_1012 ();
 sg13g2_fill_1 FILLER_47_1018 ();
 sg13g2_decap_8 FILLER_47_1036 ();
 sg13g2_decap_8 FILLER_47_1043 ();
 sg13g2_decap_4 FILLER_47_1050 ();
 sg13g2_fill_2 FILLER_47_1054 ();
 sg13g2_decap_8 FILLER_47_1061 ();
 sg13g2_decap_4 FILLER_47_1068 ();
 sg13g2_fill_1 FILLER_47_1072 ();
 sg13g2_decap_8 FILLER_47_1078 ();
 sg13g2_fill_2 FILLER_47_1085 ();
 sg13g2_decap_4 FILLER_47_1092 ();
 sg13g2_decap_4 FILLER_47_1102 ();
 sg13g2_fill_2 FILLER_47_1106 ();
 sg13g2_decap_8 FILLER_47_1118 ();
 sg13g2_decap_8 FILLER_47_1125 ();
 sg13g2_decap_8 FILLER_47_1132 ();
 sg13g2_decap_8 FILLER_47_1139 ();
 sg13g2_decap_8 FILLER_47_1156 ();
 sg13g2_decap_8 FILLER_47_1163 ();
 sg13g2_decap_8 FILLER_47_1170 ();
 sg13g2_decap_8 FILLER_47_1177 ();
 sg13g2_fill_1 FILLER_47_1188 ();
 sg13g2_decap_8 FILLER_47_1193 ();
 sg13g2_decap_4 FILLER_47_1200 ();
 sg13g2_fill_1 FILLER_47_1214 ();
 sg13g2_decap_8 FILLER_47_1224 ();
 sg13g2_decap_8 FILLER_47_1231 ();
 sg13g2_decap_8 FILLER_47_1238 ();
 sg13g2_decap_4 FILLER_47_1245 ();
 sg13g2_fill_2 FILLER_47_1249 ();
 sg13g2_decap_4 FILLER_47_1256 ();
 sg13g2_decap_8 FILLER_47_1270 ();
 sg13g2_decap_8 FILLER_47_1277 ();
 sg13g2_decap_8 FILLER_47_1284 ();
 sg13g2_decap_8 FILLER_47_1291 ();
 sg13g2_decap_8 FILLER_47_1298 ();
 sg13g2_decap_8 FILLER_47_1305 ();
 sg13g2_decap_8 FILLER_47_1312 ();
 sg13g2_decap_8 FILLER_47_1319 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_4 FILLER_48_28 ();
 sg13g2_fill_2 FILLER_48_32 ();
 sg13g2_decap_8 FILLER_48_38 ();
 sg13g2_fill_2 FILLER_48_45 ();
 sg13g2_decap_8 FILLER_48_55 ();
 sg13g2_decap_8 FILLER_48_62 ();
 sg13g2_fill_1 FILLER_48_69 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_fill_2 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_4 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_135 ();
 sg13g2_decap_8 FILLER_48_142 ();
 sg13g2_decap_8 FILLER_48_149 ();
 sg13g2_decap_4 FILLER_48_160 ();
 sg13g2_decap_8 FILLER_48_169 ();
 sg13g2_decap_4 FILLER_48_176 ();
 sg13g2_decap_8 FILLER_48_192 ();
 sg13g2_decap_8 FILLER_48_213 ();
 sg13g2_fill_2 FILLER_48_220 ();
 sg13g2_fill_2 FILLER_48_244 ();
 sg13g2_fill_1 FILLER_48_246 ();
 sg13g2_fill_2 FILLER_48_270 ();
 sg13g2_fill_1 FILLER_48_272 ();
 sg13g2_decap_8 FILLER_48_277 ();
 sg13g2_decap_8 FILLER_48_284 ();
 sg13g2_fill_2 FILLER_48_291 ();
 sg13g2_decap_8 FILLER_48_298 ();
 sg13g2_fill_1 FILLER_48_305 ();
 sg13g2_decap_8 FILLER_48_311 ();
 sg13g2_decap_4 FILLER_48_318 ();
 sg13g2_fill_1 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_327 ();
 sg13g2_decap_8 FILLER_48_334 ();
 sg13g2_fill_2 FILLER_48_341 ();
 sg13g2_decap_8 FILLER_48_348 ();
 sg13g2_fill_2 FILLER_48_355 ();
 sg13g2_fill_1 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_411 ();
 sg13g2_fill_1 FILLER_48_418 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_fill_1 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_456 ();
 sg13g2_decap_8 FILLER_48_463 ();
 sg13g2_fill_2 FILLER_48_470 ();
 sg13g2_fill_2 FILLER_48_497 ();
 sg13g2_fill_1 FILLER_48_499 ();
 sg13g2_fill_2 FILLER_48_545 ();
 sg13g2_fill_1 FILLER_48_547 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_decap_8 FILLER_48_560 ();
 sg13g2_decap_8 FILLER_48_567 ();
 sg13g2_decap_8 FILLER_48_574 ();
 sg13g2_decap_8 FILLER_48_581 ();
 sg13g2_decap_8 FILLER_48_588 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_decap_8 FILLER_48_602 ();
 sg13g2_decap_4 FILLER_48_609 ();
 sg13g2_fill_1 FILLER_48_618 ();
 sg13g2_fill_2 FILLER_48_624 ();
 sg13g2_decap_4 FILLER_48_630 ();
 sg13g2_decap_4 FILLER_48_642 ();
 sg13g2_decap_8 FILLER_48_651 ();
 sg13g2_decap_8 FILLER_48_658 ();
 sg13g2_decap_4 FILLER_48_665 ();
 sg13g2_decap_4 FILLER_48_676 ();
 sg13g2_fill_2 FILLER_48_680 ();
 sg13g2_decap_8 FILLER_48_685 ();
 sg13g2_decap_4 FILLER_48_692 ();
 sg13g2_fill_2 FILLER_48_696 ();
 sg13g2_fill_1 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_715 ();
 sg13g2_decap_8 FILLER_48_722 ();
 sg13g2_decap_8 FILLER_48_733 ();
 sg13g2_decap_4 FILLER_48_740 ();
 sg13g2_fill_2 FILLER_48_744 ();
 sg13g2_decap_4 FILLER_48_750 ();
 sg13g2_fill_2 FILLER_48_754 ();
 sg13g2_decap_4 FILLER_48_760 ();
 sg13g2_fill_1 FILLER_48_764 ();
 sg13g2_fill_1 FILLER_48_768 ();
 sg13g2_decap_8 FILLER_48_773 ();
 sg13g2_decap_8 FILLER_48_780 ();
 sg13g2_decap_8 FILLER_48_787 ();
 sg13g2_decap_4 FILLER_48_798 ();
 sg13g2_fill_2 FILLER_48_802 ();
 sg13g2_decap_8 FILLER_48_808 ();
 sg13g2_decap_8 FILLER_48_820 ();
 sg13g2_decap_8 FILLER_48_827 ();
 sg13g2_decap_8 FILLER_48_834 ();
 sg13g2_decap_8 FILLER_48_846 ();
 sg13g2_fill_2 FILLER_48_853 ();
 sg13g2_fill_1 FILLER_48_855 ();
 sg13g2_fill_2 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_48_867 ();
 sg13g2_decap_4 FILLER_48_874 ();
 sg13g2_fill_2 FILLER_48_878 ();
 sg13g2_fill_1 FILLER_48_885 ();
 sg13g2_decap_4 FILLER_48_891 ();
 sg13g2_fill_2 FILLER_48_895 ();
 sg13g2_decap_8 FILLER_48_901 ();
 sg13g2_decap_8 FILLER_48_908 ();
 sg13g2_decap_8 FILLER_48_915 ();
 sg13g2_decap_8 FILLER_48_934 ();
 sg13g2_decap_4 FILLER_48_941 ();
 sg13g2_decap_4 FILLER_48_948 ();
 sg13g2_decap_4 FILLER_48_957 ();
 sg13g2_decap_8 FILLER_48_966 ();
 sg13g2_decap_8 FILLER_48_973 ();
 sg13g2_decap_8 FILLER_48_980 ();
 sg13g2_decap_4 FILLER_48_987 ();
 sg13g2_fill_1 FILLER_48_995 ();
 sg13g2_decap_4 FILLER_48_1001 ();
 sg13g2_fill_1 FILLER_48_1005 ();
 sg13g2_decap_8 FILLER_48_1026 ();
 sg13g2_decap_4 FILLER_48_1033 ();
 sg13g2_fill_2 FILLER_48_1037 ();
 sg13g2_decap_8 FILLER_48_1044 ();
 sg13g2_decap_8 FILLER_48_1051 ();
 sg13g2_fill_1 FILLER_48_1058 ();
 sg13g2_decap_4 FILLER_48_1070 ();
 sg13g2_fill_2 FILLER_48_1079 ();
 sg13g2_decap_8 FILLER_48_1085 ();
 sg13g2_decap_8 FILLER_48_1092 ();
 sg13g2_decap_8 FILLER_48_1099 ();
 sg13g2_decap_8 FILLER_48_1106 ();
 sg13g2_decap_4 FILLER_48_1113 ();
 sg13g2_fill_1 FILLER_48_1117 ();
 sg13g2_fill_1 FILLER_48_1142 ();
 sg13g2_decap_4 FILLER_48_1155 ();
 sg13g2_fill_1 FILLER_48_1159 ();
 sg13g2_fill_2 FILLER_48_1176 ();
 sg13g2_fill_1 FILLER_48_1178 ();
 sg13g2_decap_8 FILLER_48_1183 ();
 sg13g2_decap_4 FILLER_48_1199 ();
 sg13g2_fill_2 FILLER_48_1203 ();
 sg13g2_decap_4 FILLER_48_1229 ();
 sg13g2_fill_2 FILLER_48_1233 ();
 sg13g2_fill_2 FILLER_48_1249 ();
 sg13g2_fill_1 FILLER_48_1251 ();
 sg13g2_decap_4 FILLER_48_1278 ();
 sg13g2_decap_8 FILLER_48_1287 ();
 sg13g2_decap_8 FILLER_48_1294 ();
 sg13g2_decap_8 FILLER_48_1301 ();
 sg13g2_decap_8 FILLER_48_1308 ();
 sg13g2_decap_8 FILLER_48_1315 ();
 sg13g2_decap_4 FILLER_48_1322 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_4 FILLER_49_21 ();
 sg13g2_fill_2 FILLER_49_25 ();
 sg13g2_decap_8 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_60 ();
 sg13g2_decap_8 FILLER_49_67 ();
 sg13g2_decap_8 FILLER_49_74 ();
 sg13g2_decap_8 FILLER_49_81 ();
 sg13g2_decap_8 FILLER_49_88 ();
 sg13g2_decap_8 FILLER_49_99 ();
 sg13g2_decap_8 FILLER_49_106 ();
 sg13g2_fill_2 FILLER_49_113 ();
 sg13g2_fill_1 FILLER_49_115 ();
 sg13g2_fill_1 FILLER_49_120 ();
 sg13g2_decap_8 FILLER_49_124 ();
 sg13g2_decap_8 FILLER_49_131 ();
 sg13g2_decap_8 FILLER_49_138 ();
 sg13g2_decap_4 FILLER_49_145 ();
 sg13g2_fill_1 FILLER_49_149 ();
 sg13g2_decap_8 FILLER_49_160 ();
 sg13g2_decap_8 FILLER_49_167 ();
 sg13g2_decap_8 FILLER_49_174 ();
 sg13g2_decap_8 FILLER_49_185 ();
 sg13g2_fill_2 FILLER_49_192 ();
 sg13g2_decap_8 FILLER_49_199 ();
 sg13g2_decap_8 FILLER_49_206 ();
 sg13g2_fill_2 FILLER_49_213 ();
 sg13g2_fill_2 FILLER_49_222 ();
 sg13g2_fill_1 FILLER_49_224 ();
 sg13g2_fill_1 FILLER_49_241 ();
 sg13g2_decap_4 FILLER_49_256 ();
 sg13g2_fill_1 FILLER_49_263 ();
 sg13g2_decap_8 FILLER_49_274 ();
 sg13g2_decap_8 FILLER_49_281 ();
 sg13g2_decap_8 FILLER_49_288 ();
 sg13g2_fill_2 FILLER_49_295 ();
 sg13g2_fill_1 FILLER_49_297 ();
 sg13g2_fill_1 FILLER_49_303 ();
 sg13g2_decap_8 FILLER_49_318 ();
 sg13g2_decap_8 FILLER_49_325 ();
 sg13g2_decap_8 FILLER_49_332 ();
 sg13g2_decap_8 FILLER_49_339 ();
 sg13g2_decap_8 FILLER_49_346 ();
 sg13g2_decap_4 FILLER_49_353 ();
 sg13g2_fill_1 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_362 ();
 sg13g2_decap_8 FILLER_49_369 ();
 sg13g2_decap_8 FILLER_49_376 ();
 sg13g2_decap_8 FILLER_49_383 ();
 sg13g2_decap_4 FILLER_49_390 ();
 sg13g2_decap_8 FILLER_49_400 ();
 sg13g2_decap_8 FILLER_49_407 ();
 sg13g2_fill_1 FILLER_49_414 ();
 sg13g2_decap_8 FILLER_49_436 ();
 sg13g2_decap_8 FILLER_49_443 ();
 sg13g2_decap_8 FILLER_49_450 ();
 sg13g2_decap_8 FILLER_49_457 ();
 sg13g2_decap_8 FILLER_49_464 ();
 sg13g2_decap_8 FILLER_49_471 ();
 sg13g2_decap_8 FILLER_49_478 ();
 sg13g2_decap_8 FILLER_49_485 ();
 sg13g2_decap_8 FILLER_49_492 ();
 sg13g2_decap_8 FILLER_49_499 ();
 sg13g2_decap_8 FILLER_49_506 ();
 sg13g2_decap_8 FILLER_49_513 ();
 sg13g2_fill_2 FILLER_49_520 ();
 sg13g2_fill_1 FILLER_49_522 ();
 sg13g2_fill_2 FILLER_49_527 ();
 sg13g2_decap_8 FILLER_49_555 ();
 sg13g2_decap_8 FILLER_49_562 ();
 sg13g2_decap_8 FILLER_49_569 ();
 sg13g2_decap_8 FILLER_49_576 ();
 sg13g2_decap_8 FILLER_49_583 ();
 sg13g2_decap_8 FILLER_49_590 ();
 sg13g2_decap_8 FILLER_49_597 ();
 sg13g2_decap_8 FILLER_49_604 ();
 sg13g2_fill_1 FILLER_49_611 ();
 sg13g2_decap_8 FILLER_49_642 ();
 sg13g2_decap_8 FILLER_49_649 ();
 sg13g2_decap_8 FILLER_49_656 ();
 sg13g2_decap_8 FILLER_49_663 ();
 sg13g2_decap_4 FILLER_49_670 ();
 sg13g2_fill_1 FILLER_49_674 ();
 sg13g2_fill_2 FILLER_49_687 ();
 sg13g2_decap_8 FILLER_49_705 ();
 sg13g2_decap_8 FILLER_49_717 ();
 sg13g2_decap_8 FILLER_49_724 ();
 sg13g2_decap_4 FILLER_49_731 ();
 sg13g2_fill_1 FILLER_49_735 ();
 sg13g2_fill_2 FILLER_49_751 ();
 sg13g2_fill_1 FILLER_49_753 ();
 sg13g2_decap_4 FILLER_49_759 ();
 sg13g2_fill_1 FILLER_49_763 ();
 sg13g2_fill_2 FILLER_49_768 ();
 sg13g2_decap_8 FILLER_49_779 ();
 sg13g2_decap_4 FILLER_49_812 ();
 sg13g2_fill_2 FILLER_49_816 ();
 sg13g2_decap_8 FILLER_49_824 ();
 sg13g2_decap_8 FILLER_49_831 ();
 sg13g2_fill_2 FILLER_49_838 ();
 sg13g2_fill_1 FILLER_49_840 ();
 sg13g2_decap_8 FILLER_49_846 ();
 sg13g2_decap_8 FILLER_49_853 ();
 sg13g2_decap_8 FILLER_49_860 ();
 sg13g2_decap_8 FILLER_49_867 ();
 sg13g2_decap_8 FILLER_49_874 ();
 sg13g2_decap_4 FILLER_49_881 ();
 sg13g2_fill_1 FILLER_49_885 ();
 sg13g2_decap_4 FILLER_49_915 ();
 sg13g2_fill_2 FILLER_49_924 ();
 sg13g2_decap_8 FILLER_49_936 ();
 sg13g2_decap_8 FILLER_49_952 ();
 sg13g2_decap_8 FILLER_49_959 ();
 sg13g2_fill_1 FILLER_49_966 ();
 sg13g2_decap_8 FILLER_49_972 ();
 sg13g2_decap_4 FILLER_49_979 ();
 sg13g2_fill_2 FILLER_49_988 ();
 sg13g2_decap_8 FILLER_49_1004 ();
 sg13g2_fill_2 FILLER_49_1011 ();
 sg13g2_decap_8 FILLER_49_1032 ();
 sg13g2_decap_8 FILLER_49_1039 ();
 sg13g2_decap_8 FILLER_49_1046 ();
 sg13g2_fill_1 FILLER_49_1053 ();
 sg13g2_fill_1 FILLER_49_1059 ();
 sg13g2_decap_4 FILLER_49_1068 ();
 sg13g2_fill_2 FILLER_49_1072 ();
 sg13g2_decap_8 FILLER_49_1080 ();
 sg13g2_decap_8 FILLER_49_1087 ();
 sg13g2_decap_8 FILLER_49_1094 ();
 sg13g2_fill_2 FILLER_49_1101 ();
 sg13g2_fill_1 FILLER_49_1103 ();
 sg13g2_decap_4 FILLER_49_1108 ();
 sg13g2_fill_2 FILLER_49_1112 ();
 sg13g2_decap_8 FILLER_49_1128 ();
 sg13g2_fill_1 FILLER_49_1135 ();
 sg13g2_fill_2 FILLER_49_1145 ();
 sg13g2_decap_8 FILLER_49_1153 ();
 sg13g2_fill_2 FILLER_49_1160 ();
 sg13g2_decap_8 FILLER_49_1166 ();
 sg13g2_fill_2 FILLER_49_1173 ();
 sg13g2_decap_8 FILLER_49_1180 ();
 sg13g2_fill_2 FILLER_49_1187 ();
 sg13g2_fill_1 FILLER_49_1189 ();
 sg13g2_fill_1 FILLER_49_1208 ();
 sg13g2_decap_8 FILLER_49_1213 ();
 sg13g2_fill_2 FILLER_49_1220 ();
 sg13g2_fill_1 FILLER_49_1222 ();
 sg13g2_decap_8 FILLER_49_1227 ();
 sg13g2_fill_2 FILLER_49_1234 ();
 sg13g2_fill_2 FILLER_49_1241 ();
 sg13g2_fill_1 FILLER_49_1249 ();
 sg13g2_decap_4 FILLER_49_1254 ();
 sg13g2_decap_8 FILLER_49_1276 ();
 sg13g2_decap_8 FILLER_49_1283 ();
 sg13g2_decap_8 FILLER_49_1290 ();
 sg13g2_decap_8 FILLER_49_1297 ();
 sg13g2_decap_8 FILLER_49_1304 ();
 sg13g2_decap_8 FILLER_49_1311 ();
 sg13g2_decap_8 FILLER_49_1318 ();
 sg13g2_fill_1 FILLER_49_1325 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_13 ();
 sg13g2_decap_8 FILLER_50_20 ();
 sg13g2_decap_4 FILLER_50_27 ();
 sg13g2_fill_1 FILLER_50_31 ();
 sg13g2_fill_1 FILLER_50_37 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_fill_2 FILLER_50_49 ();
 sg13g2_fill_2 FILLER_50_56 ();
 sg13g2_fill_1 FILLER_50_58 ();
 sg13g2_decap_8 FILLER_50_62 ();
 sg13g2_decap_8 FILLER_50_99 ();
 sg13g2_decap_4 FILLER_50_106 ();
 sg13g2_fill_2 FILLER_50_119 ();
 sg13g2_decap_4 FILLER_50_126 ();
 sg13g2_fill_2 FILLER_50_130 ();
 sg13g2_decap_8 FILLER_50_171 ();
 sg13g2_decap_8 FILLER_50_178 ();
 sg13g2_fill_2 FILLER_50_185 ();
 sg13g2_fill_1 FILLER_50_187 ();
 sg13g2_decap_4 FILLER_50_191 ();
 sg13g2_fill_1 FILLER_50_195 ();
 sg13g2_decap_4 FILLER_50_216 ();
 sg13g2_decap_4 FILLER_50_224 ();
 sg13g2_decap_4 FILLER_50_233 ();
 sg13g2_fill_1 FILLER_50_237 ();
 sg13g2_decap_4 FILLER_50_242 ();
 sg13g2_decap_8 FILLER_50_275 ();
 sg13g2_decap_8 FILLER_50_282 ();
 sg13g2_decap_8 FILLER_50_289 ();
 sg13g2_decap_4 FILLER_50_296 ();
 sg13g2_decap_8 FILLER_50_304 ();
 sg13g2_fill_1 FILLER_50_311 ();
 sg13g2_decap_8 FILLER_50_317 ();
 sg13g2_decap_8 FILLER_50_324 ();
 sg13g2_decap_8 FILLER_50_331 ();
 sg13g2_decap_8 FILLER_50_338 ();
 sg13g2_decap_8 FILLER_50_345 ();
 sg13g2_decap_4 FILLER_50_352 ();
 sg13g2_decap_8 FILLER_50_361 ();
 sg13g2_decap_4 FILLER_50_368 ();
 sg13g2_fill_2 FILLER_50_372 ();
 sg13g2_decap_8 FILLER_50_379 ();
 sg13g2_fill_2 FILLER_50_386 ();
 sg13g2_fill_1 FILLER_50_388 ();
 sg13g2_decap_8 FILLER_50_410 ();
 sg13g2_fill_2 FILLER_50_417 ();
 sg13g2_decap_8 FILLER_50_424 ();
 sg13g2_decap_8 FILLER_50_431 ();
 sg13g2_fill_1 FILLER_50_438 ();
 sg13g2_decap_8 FILLER_50_460 ();
 sg13g2_decap_8 FILLER_50_467 ();
 sg13g2_decap_8 FILLER_50_474 ();
 sg13g2_decap_8 FILLER_50_481 ();
 sg13g2_decap_8 FILLER_50_488 ();
 sg13g2_decap_8 FILLER_50_495 ();
 sg13g2_decap_8 FILLER_50_502 ();
 sg13g2_decap_8 FILLER_50_509 ();
 sg13g2_decap_8 FILLER_50_516 ();
 sg13g2_decap_8 FILLER_50_523 ();
 sg13g2_decap_4 FILLER_50_530 ();
 sg13g2_fill_1 FILLER_50_534 ();
 sg13g2_decap_8 FILLER_50_539 ();
 sg13g2_decap_8 FILLER_50_546 ();
 sg13g2_decap_8 FILLER_50_553 ();
 sg13g2_decap_4 FILLER_50_560 ();
 sg13g2_fill_1 FILLER_50_564 ();
 sg13g2_decap_8 FILLER_50_599 ();
 sg13g2_decap_4 FILLER_50_606 ();
 sg13g2_decap_4 FILLER_50_615 ();
 sg13g2_fill_1 FILLER_50_619 ();
 sg13g2_decap_8 FILLER_50_624 ();
 sg13g2_decap_8 FILLER_50_631 ();
 sg13g2_decap_8 FILLER_50_638 ();
 sg13g2_decap_8 FILLER_50_645 ();
 sg13g2_decap_8 FILLER_50_652 ();
 sg13g2_decap_8 FILLER_50_659 ();
 sg13g2_decap_8 FILLER_50_666 ();
 sg13g2_decap_8 FILLER_50_677 ();
 sg13g2_decap_8 FILLER_50_684 ();
 sg13g2_decap_8 FILLER_50_691 ();
 sg13g2_decap_4 FILLER_50_701 ();
 sg13g2_fill_2 FILLER_50_705 ();
 sg13g2_fill_2 FILLER_50_733 ();
 sg13g2_fill_1 FILLER_50_735 ();
 sg13g2_decap_8 FILLER_50_739 ();
 sg13g2_decap_8 FILLER_50_746 ();
 sg13g2_fill_2 FILLER_50_753 ();
 sg13g2_fill_2 FILLER_50_759 ();
 sg13g2_fill_2 FILLER_50_765 ();
 sg13g2_fill_1 FILLER_50_767 ();
 sg13g2_decap_4 FILLER_50_786 ();
 sg13g2_fill_1 FILLER_50_790 ();
 sg13g2_decap_8 FILLER_50_801 ();
 sg13g2_decap_4 FILLER_50_808 ();
 sg13g2_fill_1 FILLER_50_812 ();
 sg13g2_decap_8 FILLER_50_823 ();
 sg13g2_decap_8 FILLER_50_830 ();
 sg13g2_decap_8 FILLER_50_837 ();
 sg13g2_decap_4 FILLER_50_844 ();
 sg13g2_fill_1 FILLER_50_848 ();
 sg13g2_decap_8 FILLER_50_853 ();
 sg13g2_decap_8 FILLER_50_860 ();
 sg13g2_decap_4 FILLER_50_867 ();
 sg13g2_fill_2 FILLER_50_871 ();
 sg13g2_decap_8 FILLER_50_891 ();
 sg13g2_decap_8 FILLER_50_898 ();
 sg13g2_decap_8 FILLER_50_905 ();
 sg13g2_fill_2 FILLER_50_912 ();
 sg13g2_fill_1 FILLER_50_914 ();
 sg13g2_decap_4 FILLER_50_920 ();
 sg13g2_fill_1 FILLER_50_924 ();
 sg13g2_decap_8 FILLER_50_930 ();
 sg13g2_decap_8 FILLER_50_937 ();
 sg13g2_decap_8 FILLER_50_944 ();
 sg13g2_decap_8 FILLER_50_951 ();
 sg13g2_fill_2 FILLER_50_958 ();
 sg13g2_fill_1 FILLER_50_960 ();
 sg13g2_decap_8 FILLER_50_966 ();
 sg13g2_fill_1 FILLER_50_973 ();
 sg13g2_decap_8 FILLER_50_979 ();
 sg13g2_decap_4 FILLER_50_986 ();
 sg13g2_fill_1 FILLER_50_999 ();
 sg13g2_decap_8 FILLER_50_1005 ();
 sg13g2_decap_8 FILLER_50_1012 ();
 sg13g2_decap_4 FILLER_50_1019 ();
 sg13g2_fill_1 FILLER_50_1023 ();
 sg13g2_decap_8 FILLER_50_1034 ();
 sg13g2_decap_8 FILLER_50_1041 ();
 sg13g2_decap_4 FILLER_50_1048 ();
 sg13g2_fill_1 FILLER_50_1052 ();
 sg13g2_fill_2 FILLER_50_1062 ();
 sg13g2_fill_1 FILLER_50_1064 ();
 sg13g2_decap_8 FILLER_50_1069 ();
 sg13g2_decap_8 FILLER_50_1076 ();
 sg13g2_decap_8 FILLER_50_1083 ();
 sg13g2_decap_4 FILLER_50_1090 ();
 sg13g2_fill_1 FILLER_50_1094 ();
 sg13g2_decap_4 FILLER_50_1100 ();
 sg13g2_fill_1 FILLER_50_1104 ();
 sg13g2_decap_8 FILLER_50_1118 ();
 sg13g2_decap_8 FILLER_50_1125 ();
 sg13g2_fill_2 FILLER_50_1132 ();
 sg13g2_fill_1 FILLER_50_1134 ();
 sg13g2_decap_8 FILLER_50_1140 ();
 sg13g2_decap_8 FILLER_50_1147 ();
 sg13g2_decap_4 FILLER_50_1154 ();
 sg13g2_fill_1 FILLER_50_1162 ();
 sg13g2_decap_8 FILLER_50_1168 ();
 sg13g2_decap_8 FILLER_50_1175 ();
 sg13g2_decap_8 FILLER_50_1182 ();
 sg13g2_decap_8 FILLER_50_1189 ();
 sg13g2_decap_4 FILLER_50_1196 ();
 sg13g2_decap_8 FILLER_50_1205 ();
 sg13g2_fill_1 FILLER_50_1223 ();
 sg13g2_decap_4 FILLER_50_1228 ();
 sg13g2_fill_2 FILLER_50_1232 ();
 sg13g2_decap_8 FILLER_50_1239 ();
 sg13g2_decap_8 FILLER_50_1254 ();
 sg13g2_decap_4 FILLER_50_1261 ();
 sg13g2_fill_2 FILLER_50_1273 ();
 sg13g2_fill_1 FILLER_50_1275 ();
 sg13g2_decap_8 FILLER_50_1285 ();
 sg13g2_decap_8 FILLER_50_1292 ();
 sg13g2_decap_8 FILLER_50_1299 ();
 sg13g2_decap_8 FILLER_50_1306 ();
 sg13g2_decap_8 FILLER_50_1313 ();
 sg13g2_decap_4 FILLER_50_1320 ();
 sg13g2_fill_2 FILLER_50_1324 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_53 ();
 sg13g2_decap_8 FILLER_51_65 ();
 sg13g2_decap_4 FILLER_51_72 ();
 sg13g2_fill_2 FILLER_51_76 ();
 sg13g2_fill_1 FILLER_51_97 ();
 sg13g2_decap_8 FILLER_51_103 ();
 sg13g2_decap_8 FILLER_51_110 ();
 sg13g2_decap_8 FILLER_51_117 ();
 sg13g2_decap_8 FILLER_51_124 ();
 sg13g2_decap_8 FILLER_51_131 ();
 sg13g2_decap_8 FILLER_51_138 ();
 sg13g2_fill_2 FILLER_51_145 ();
 sg13g2_decap_8 FILLER_51_166 ();
 sg13g2_decap_8 FILLER_51_173 ();
 sg13g2_decap_8 FILLER_51_180 ();
 sg13g2_decap_8 FILLER_51_239 ();
 sg13g2_fill_2 FILLER_51_246 ();
 sg13g2_fill_1 FILLER_51_248 ();
 sg13g2_decap_8 FILLER_51_253 ();
 sg13g2_decap_8 FILLER_51_274 ();
 sg13g2_decap_8 FILLER_51_281 ();
 sg13g2_decap_8 FILLER_51_288 ();
 sg13g2_decap_8 FILLER_51_295 ();
 sg13g2_decap_8 FILLER_51_302 ();
 sg13g2_decap_8 FILLER_51_309 ();
 sg13g2_decap_8 FILLER_51_316 ();
 sg13g2_decap_8 FILLER_51_323 ();
 sg13g2_decap_4 FILLER_51_330 ();
 sg13g2_decap_8 FILLER_51_343 ();
 sg13g2_decap_8 FILLER_51_350 ();
 sg13g2_decap_8 FILLER_51_357 ();
 sg13g2_decap_8 FILLER_51_364 ();
 sg13g2_fill_1 FILLER_51_371 ();
 sg13g2_decap_8 FILLER_51_377 ();
 sg13g2_decap_8 FILLER_51_384 ();
 sg13g2_decap_8 FILLER_51_391 ();
 sg13g2_decap_8 FILLER_51_398 ();
 sg13g2_decap_8 FILLER_51_405 ();
 sg13g2_decap_8 FILLER_51_412 ();
 sg13g2_decap_8 FILLER_51_419 ();
 sg13g2_decap_8 FILLER_51_426 ();
 sg13g2_decap_8 FILLER_51_433 ();
 sg13g2_decap_8 FILLER_51_440 ();
 sg13g2_decap_8 FILLER_51_447 ();
 sg13g2_decap_8 FILLER_51_454 ();
 sg13g2_decap_8 FILLER_51_461 ();
 sg13g2_decap_8 FILLER_51_468 ();
 sg13g2_decap_8 FILLER_51_475 ();
 sg13g2_decap_8 FILLER_51_482 ();
 sg13g2_decap_8 FILLER_51_489 ();
 sg13g2_decap_8 FILLER_51_496 ();
 sg13g2_decap_8 FILLER_51_503 ();
 sg13g2_decap_8 FILLER_51_510 ();
 sg13g2_decap_8 FILLER_51_517 ();
 sg13g2_decap_8 FILLER_51_524 ();
 sg13g2_decap_8 FILLER_51_531 ();
 sg13g2_decap_8 FILLER_51_538 ();
 sg13g2_decap_8 FILLER_51_545 ();
 sg13g2_decap_8 FILLER_51_552 ();
 sg13g2_decap_8 FILLER_51_559 ();
 sg13g2_fill_2 FILLER_51_566 ();
 sg13g2_fill_1 FILLER_51_568 ();
 sg13g2_fill_1 FILLER_51_587 ();
 sg13g2_decap_4 FILLER_51_592 ();
 sg13g2_fill_2 FILLER_51_596 ();
 sg13g2_fill_2 FILLER_51_624 ();
 sg13g2_decap_8 FILLER_51_634 ();
 sg13g2_decap_8 FILLER_51_641 ();
 sg13g2_decap_8 FILLER_51_648 ();
 sg13g2_decap_8 FILLER_51_655 ();
 sg13g2_decap_8 FILLER_51_662 ();
 sg13g2_decap_8 FILLER_51_669 ();
 sg13g2_decap_4 FILLER_51_676 ();
 sg13g2_fill_2 FILLER_51_685 ();
 sg13g2_decap_8 FILLER_51_691 ();
 sg13g2_decap_8 FILLER_51_698 ();
 sg13g2_decap_8 FILLER_51_705 ();
 sg13g2_decap_8 FILLER_51_716 ();
 sg13g2_decap_8 FILLER_51_723 ();
 sg13g2_decap_8 FILLER_51_730 ();
 sg13g2_fill_1 FILLER_51_737 ();
 sg13g2_fill_2 FILLER_51_746 ();
 sg13g2_fill_1 FILLER_51_748 ();
 sg13g2_fill_2 FILLER_51_753 ();
 sg13g2_fill_2 FILLER_51_763 ();
 sg13g2_decap_8 FILLER_51_782 ();
 sg13g2_fill_2 FILLER_51_789 ();
 sg13g2_decap_8 FILLER_51_801 ();
 sg13g2_decap_8 FILLER_51_808 ();
 sg13g2_decap_8 FILLER_51_815 ();
 sg13g2_decap_8 FILLER_51_822 ();
 sg13g2_decap_8 FILLER_51_829 ();
 sg13g2_decap_8 FILLER_51_836 ();
 sg13g2_decap_8 FILLER_51_843 ();
 sg13g2_decap_8 FILLER_51_850 ();
 sg13g2_decap_8 FILLER_51_857 ();
 sg13g2_decap_8 FILLER_51_864 ();
 sg13g2_decap_8 FILLER_51_871 ();
 sg13g2_decap_8 FILLER_51_878 ();
 sg13g2_fill_1 FILLER_51_885 ();
 sg13g2_decap_8 FILLER_51_895 ();
 sg13g2_decap_8 FILLER_51_902 ();
 sg13g2_fill_2 FILLER_51_909 ();
 sg13g2_fill_1 FILLER_51_911 ();
 sg13g2_decap_8 FILLER_51_920 ();
 sg13g2_fill_2 FILLER_51_927 ();
 sg13g2_decap_8 FILLER_51_933 ();
 sg13g2_decap_8 FILLER_51_955 ();
 sg13g2_decap_4 FILLER_51_969 ();
 sg13g2_fill_1 FILLER_51_973 ();
 sg13g2_decap_4 FILLER_51_979 ();
 sg13g2_fill_1 FILLER_51_983 ();
 sg13g2_decap_8 FILLER_51_992 ();
 sg13g2_decap_8 FILLER_51_999 ();
 sg13g2_fill_2 FILLER_51_1006 ();
 sg13g2_decap_8 FILLER_51_1017 ();
 sg13g2_decap_8 FILLER_51_1024 ();
 sg13g2_decap_8 FILLER_51_1031 ();
 sg13g2_decap_8 FILLER_51_1038 ();
 sg13g2_decap_8 FILLER_51_1045 ();
 sg13g2_decap_4 FILLER_51_1052 ();
 sg13g2_fill_2 FILLER_51_1056 ();
 sg13g2_decap_8 FILLER_51_1071 ();
 sg13g2_decap_4 FILLER_51_1078 ();
 sg13g2_decap_4 FILLER_51_1087 ();
 sg13g2_decap_4 FILLER_51_1100 ();
 sg13g2_fill_2 FILLER_51_1114 ();
 sg13g2_fill_2 FILLER_51_1129 ();
 sg13g2_fill_1 FILLER_51_1131 ();
 sg13g2_decap_4 FILLER_51_1144 ();
 sg13g2_decap_8 FILLER_51_1153 ();
 sg13g2_decap_8 FILLER_51_1165 ();
 sg13g2_fill_1 FILLER_51_1172 ();
 sg13g2_decap_8 FILLER_51_1177 ();
 sg13g2_decap_8 FILLER_51_1184 ();
 sg13g2_decap_8 FILLER_51_1191 ();
 sg13g2_fill_1 FILLER_51_1198 ();
 sg13g2_fill_2 FILLER_51_1207 ();
 sg13g2_fill_2 FILLER_51_1213 ();
 sg13g2_fill_1 FILLER_51_1215 ();
 sg13g2_fill_2 FILLER_51_1225 ();
 sg13g2_decap_4 FILLER_51_1231 ();
 sg13g2_decap_8 FILLER_51_1240 ();
 sg13g2_decap_8 FILLER_51_1247 ();
 sg13g2_decap_4 FILLER_51_1259 ();
 sg13g2_fill_1 FILLER_51_1263 ();
 sg13g2_fill_2 FILLER_51_1269 ();
 sg13g2_fill_1 FILLER_51_1271 ();
 sg13g2_decap_8 FILLER_51_1277 ();
 sg13g2_decap_8 FILLER_51_1284 ();
 sg13g2_decap_8 FILLER_51_1291 ();
 sg13g2_decap_8 FILLER_51_1298 ();
 sg13g2_decap_8 FILLER_51_1305 ();
 sg13g2_decap_8 FILLER_51_1312 ();
 sg13g2_decap_8 FILLER_51_1319 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_4 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_66 ();
 sg13g2_decap_8 FILLER_52_73 ();
 sg13g2_decap_8 FILLER_52_80 ();
 sg13g2_decap_4 FILLER_52_87 ();
 sg13g2_fill_2 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_fill_2 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_122 ();
 sg13g2_fill_2 FILLER_52_129 ();
 sg13g2_fill_1 FILLER_52_131 ();
 sg13g2_decap_8 FILLER_52_142 ();
 sg13g2_fill_2 FILLER_52_149 ();
 sg13g2_fill_1 FILLER_52_151 ();
 sg13g2_decap_8 FILLER_52_157 ();
 sg13g2_decap_8 FILLER_52_164 ();
 sg13g2_decap_8 FILLER_52_171 ();
 sg13g2_decap_8 FILLER_52_178 ();
 sg13g2_fill_2 FILLER_52_185 ();
 sg13g2_fill_1 FILLER_52_187 ();
 sg13g2_decap_8 FILLER_52_205 ();
 sg13g2_decap_8 FILLER_52_212 ();
 sg13g2_decap_8 FILLER_52_219 ();
 sg13g2_decap_8 FILLER_52_226 ();
 sg13g2_fill_2 FILLER_52_233 ();
 sg13g2_fill_2 FILLER_52_240 ();
 sg13g2_decap_8 FILLER_52_246 ();
 sg13g2_decap_8 FILLER_52_258 ();
 sg13g2_fill_1 FILLER_52_265 ();
 sg13g2_decap_8 FILLER_52_270 ();
 sg13g2_decap_8 FILLER_52_277 ();
 sg13g2_fill_2 FILLER_52_284 ();
 sg13g2_fill_1 FILLER_52_286 ();
 sg13g2_decap_8 FILLER_52_292 ();
 sg13g2_fill_1 FILLER_52_299 ();
 sg13g2_fill_2 FILLER_52_304 ();
 sg13g2_fill_1 FILLER_52_306 ();
 sg13g2_decap_8 FILLER_52_316 ();
 sg13g2_fill_2 FILLER_52_323 ();
 sg13g2_fill_1 FILLER_52_325 ();
 sg13g2_decap_8 FILLER_52_356 ();
 sg13g2_decap_8 FILLER_52_363 ();
 sg13g2_fill_2 FILLER_52_370 ();
 sg13g2_fill_1 FILLER_52_372 ();
 sg13g2_decap_8 FILLER_52_378 ();
 sg13g2_decap_8 FILLER_52_385 ();
 sg13g2_decap_8 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_decap_8 FILLER_52_406 ();
 sg13g2_decap_8 FILLER_52_413 ();
 sg13g2_decap_8 FILLER_52_420 ();
 sg13g2_decap_8 FILLER_52_427 ();
 sg13g2_decap_8 FILLER_52_434 ();
 sg13g2_decap_4 FILLER_52_441 ();
 sg13g2_fill_1 FILLER_52_445 ();
 sg13g2_decap_8 FILLER_52_451 ();
 sg13g2_decap_8 FILLER_52_458 ();
 sg13g2_decap_8 FILLER_52_465 ();
 sg13g2_decap_8 FILLER_52_472 ();
 sg13g2_decap_8 FILLER_52_479 ();
 sg13g2_decap_8 FILLER_52_486 ();
 sg13g2_fill_2 FILLER_52_493 ();
 sg13g2_fill_1 FILLER_52_495 ();
 sg13g2_fill_1 FILLER_52_500 ();
 sg13g2_fill_1 FILLER_52_510 ();
 sg13g2_decap_8 FILLER_52_516 ();
 sg13g2_decap_8 FILLER_52_523 ();
 sg13g2_decap_8 FILLER_52_530 ();
 sg13g2_decap_8 FILLER_52_537 ();
 sg13g2_decap_8 FILLER_52_544 ();
 sg13g2_decap_8 FILLER_52_551 ();
 sg13g2_decap_8 FILLER_52_558 ();
 sg13g2_decap_8 FILLER_52_565 ();
 sg13g2_decap_8 FILLER_52_572 ();
 sg13g2_decap_4 FILLER_52_579 ();
 sg13g2_fill_1 FILLER_52_583 ();
 sg13g2_decap_8 FILLER_52_590 ();
 sg13g2_decap_8 FILLER_52_597 ();
 sg13g2_decap_4 FILLER_52_617 ();
 sg13g2_fill_1 FILLER_52_621 ();
 sg13g2_decap_8 FILLER_52_626 ();
 sg13g2_decap_4 FILLER_52_633 ();
 sg13g2_decap_8 FILLER_52_663 ();
 sg13g2_decap_4 FILLER_52_674 ();
 sg13g2_fill_2 FILLER_52_678 ();
 sg13g2_decap_8 FILLER_52_706 ();
 sg13g2_decap_8 FILLER_52_713 ();
 sg13g2_decap_8 FILLER_52_720 ();
 sg13g2_decap_4 FILLER_52_727 ();
 sg13g2_decap_8 FILLER_52_736 ();
 sg13g2_decap_8 FILLER_52_743 ();
 sg13g2_fill_2 FILLER_52_750 ();
 sg13g2_fill_2 FILLER_52_756 ();
 sg13g2_fill_1 FILLER_52_758 ();
 sg13g2_fill_1 FILLER_52_763 ();
 sg13g2_decap_4 FILLER_52_768 ();
 sg13g2_decap_8 FILLER_52_780 ();
 sg13g2_decap_8 FILLER_52_787 ();
 sg13g2_decap_8 FILLER_52_794 ();
 sg13g2_fill_2 FILLER_52_801 ();
 sg13g2_fill_1 FILLER_52_803 ();
 sg13g2_decap_8 FILLER_52_809 ();
 sg13g2_decap_8 FILLER_52_816 ();
 sg13g2_decap_8 FILLER_52_823 ();
 sg13g2_decap_8 FILLER_52_830 ();
 sg13g2_decap_8 FILLER_52_837 ();
 sg13g2_decap_8 FILLER_52_844 ();
 sg13g2_decap_8 FILLER_52_851 ();
 sg13g2_decap_8 FILLER_52_858 ();
 sg13g2_decap_8 FILLER_52_865 ();
 sg13g2_decap_8 FILLER_52_872 ();
 sg13g2_decap_4 FILLER_52_879 ();
 sg13g2_decap_8 FILLER_52_887 ();
 sg13g2_decap_4 FILLER_52_894 ();
 sg13g2_decap_8 FILLER_52_907 ();
 sg13g2_decap_8 FILLER_52_914 ();
 sg13g2_fill_2 FILLER_52_921 ();
 sg13g2_fill_1 FILLER_52_923 ();
 sg13g2_fill_1 FILLER_52_934 ();
 sg13g2_fill_2 FILLER_52_944 ();
 sg13g2_fill_1 FILLER_52_946 ();
 sg13g2_fill_2 FILLER_52_952 ();
 sg13g2_fill_1 FILLER_52_954 ();
 sg13g2_fill_1 FILLER_52_963 ();
 sg13g2_decap_4 FILLER_52_969 ();
 sg13g2_decap_4 FILLER_52_978 ();
 sg13g2_fill_1 FILLER_52_982 ();
 sg13g2_decap_8 FILLER_52_988 ();
 sg13g2_decap_8 FILLER_52_995 ();
 sg13g2_fill_1 FILLER_52_1002 ();
 sg13g2_decap_8 FILLER_52_1013 ();
 sg13g2_decap_4 FILLER_52_1020 ();
 sg13g2_fill_1 FILLER_52_1024 ();
 sg13g2_decap_4 FILLER_52_1038 ();
 sg13g2_fill_1 FILLER_52_1042 ();
 sg13g2_decap_4 FILLER_52_1048 ();
 sg13g2_fill_2 FILLER_52_1052 ();
 sg13g2_fill_2 FILLER_52_1069 ();
 sg13g2_decap_8 FILLER_52_1080 ();
 sg13g2_decap_8 FILLER_52_1087 ();
 sg13g2_fill_2 FILLER_52_1094 ();
 sg13g2_decap_8 FILLER_52_1101 ();
 sg13g2_fill_2 FILLER_52_1108 ();
 sg13g2_fill_1 FILLER_52_1110 ();
 sg13g2_decap_8 FILLER_52_1116 ();
 sg13g2_decap_8 FILLER_52_1123 ();
 sg13g2_fill_1 FILLER_52_1130 ();
 sg13g2_fill_2 FILLER_52_1136 ();
 sg13g2_fill_1 FILLER_52_1138 ();
 sg13g2_fill_2 FILLER_52_1143 ();
 sg13g2_fill_1 FILLER_52_1145 ();
 sg13g2_fill_2 FILLER_52_1151 ();
 sg13g2_fill_1 FILLER_52_1153 ();
 sg13g2_decap_8 FILLER_52_1170 ();
 sg13g2_decap_8 FILLER_52_1182 ();
 sg13g2_fill_2 FILLER_52_1189 ();
 sg13g2_fill_1 FILLER_52_1191 ();
 sg13g2_decap_8 FILLER_52_1200 ();
 sg13g2_fill_1 FILLER_52_1207 ();
 sg13g2_decap_8 FILLER_52_1213 ();
 sg13g2_decap_8 FILLER_52_1220 ();
 sg13g2_decap_4 FILLER_52_1227 ();
 sg13g2_fill_1 FILLER_52_1231 ();
 sg13g2_decap_4 FILLER_52_1237 ();
 sg13g2_fill_1 FILLER_52_1241 ();
 sg13g2_fill_2 FILLER_52_1250 ();
 sg13g2_decap_8 FILLER_52_1260 ();
 sg13g2_fill_2 FILLER_52_1267 ();
 sg13g2_fill_2 FILLER_52_1273 ();
 sg13g2_decap_8 FILLER_52_1281 ();
 sg13g2_decap_8 FILLER_52_1288 ();
 sg13g2_decap_8 FILLER_52_1295 ();
 sg13g2_decap_8 FILLER_52_1302 ();
 sg13g2_decap_8 FILLER_52_1309 ();
 sg13g2_decap_8 FILLER_52_1316 ();
 sg13g2_fill_2 FILLER_52_1323 ();
 sg13g2_fill_1 FILLER_52_1325 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_4 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_4 FILLER_53_77 ();
 sg13g2_fill_2 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_99 ();
 sg13g2_decap_4 FILLER_53_106 ();
 sg13g2_fill_1 FILLER_53_110 ();
 sg13g2_decap_8 FILLER_53_137 ();
 sg13g2_decap_8 FILLER_53_144 ();
 sg13g2_decap_8 FILLER_53_151 ();
 sg13g2_decap_8 FILLER_53_158 ();
 sg13g2_decap_8 FILLER_53_165 ();
 sg13g2_decap_8 FILLER_53_172 ();
 sg13g2_decap_8 FILLER_53_179 ();
 sg13g2_decap_8 FILLER_53_186 ();
 sg13g2_decap_8 FILLER_53_193 ();
 sg13g2_decap_4 FILLER_53_200 ();
 sg13g2_fill_1 FILLER_53_204 ();
 sg13g2_decap_8 FILLER_53_211 ();
 sg13g2_decap_4 FILLER_53_218 ();
 sg13g2_fill_2 FILLER_53_222 ();
 sg13g2_decap_8 FILLER_53_229 ();
 sg13g2_fill_2 FILLER_53_236 ();
 sg13g2_fill_1 FILLER_53_238 ();
 sg13g2_fill_1 FILLER_53_243 ();
 sg13g2_fill_1 FILLER_53_249 ();
 sg13g2_fill_2 FILLER_53_255 ();
 sg13g2_fill_1 FILLER_53_257 ();
 sg13g2_decap_4 FILLER_53_284 ();
 sg13g2_decap_8 FILLER_53_292 ();
 sg13g2_decap_4 FILLER_53_299 ();
 sg13g2_fill_2 FILLER_53_312 ();
 sg13g2_fill_2 FILLER_53_318 ();
 sg13g2_decap_8 FILLER_53_344 ();
 sg13g2_decap_4 FILLER_53_351 ();
 sg13g2_fill_1 FILLER_53_355 ();
 sg13g2_decap_4 FILLER_53_361 ();
 sg13g2_decap_4 FILLER_53_369 ();
 sg13g2_fill_1 FILLER_53_382 ();
 sg13g2_fill_1 FILLER_53_388 ();
 sg13g2_fill_2 FILLER_53_393 ();
 sg13g2_fill_2 FILLER_53_400 ();
 sg13g2_fill_2 FILLER_53_405 ();
 sg13g2_fill_1 FILLER_53_407 ();
 sg13g2_fill_2 FILLER_53_418 ();
 sg13g2_fill_2 FILLER_53_432 ();
 sg13g2_decap_8 FILLER_53_439 ();
 sg13g2_fill_1 FILLER_53_446 ();
 sg13g2_decap_4 FILLER_53_480 ();
 sg13g2_fill_2 FILLER_53_497 ();
 sg13g2_fill_2 FILLER_53_510 ();
 sg13g2_fill_1 FILLER_53_512 ();
 sg13g2_decap_8 FILLER_53_543 ();
 sg13g2_decap_8 FILLER_53_550 ();
 sg13g2_decap_4 FILLER_53_557 ();
 sg13g2_fill_2 FILLER_53_561 ();
 sg13g2_decap_4 FILLER_53_573 ();
 sg13g2_fill_1 FILLER_53_577 ();
 sg13g2_decap_8 FILLER_53_586 ();
 sg13g2_decap_8 FILLER_53_593 ();
 sg13g2_decap_8 FILLER_53_600 ();
 sg13g2_decap_8 FILLER_53_607 ();
 sg13g2_decap_8 FILLER_53_614 ();
 sg13g2_decap_8 FILLER_53_621 ();
 sg13g2_decap_8 FILLER_53_628 ();
 sg13g2_decap_4 FILLER_53_635 ();
 sg13g2_fill_2 FILLER_53_639 ();
 sg13g2_decap_8 FILLER_53_657 ();
 sg13g2_decap_8 FILLER_53_664 ();
 sg13g2_decap_8 FILLER_53_671 ();
 sg13g2_decap_8 FILLER_53_678 ();
 sg13g2_decap_8 FILLER_53_685 ();
 sg13g2_decap_8 FILLER_53_692 ();
 sg13g2_decap_8 FILLER_53_699 ();
 sg13g2_fill_1 FILLER_53_706 ();
 sg13g2_decap_8 FILLER_53_722 ();
 sg13g2_decap_8 FILLER_53_729 ();
 sg13g2_decap_8 FILLER_53_736 ();
 sg13g2_decap_8 FILLER_53_743 ();
 sg13g2_fill_1 FILLER_53_750 ();
 sg13g2_decap_8 FILLER_53_759 ();
 sg13g2_fill_2 FILLER_53_766 ();
 sg13g2_decap_8 FILLER_53_778 ();
 sg13g2_decap_8 FILLER_53_785 ();
 sg13g2_decap_8 FILLER_53_792 ();
 sg13g2_fill_2 FILLER_53_799 ();
 sg13g2_fill_1 FILLER_53_808 ();
 sg13g2_fill_2 FILLER_53_835 ();
 sg13g2_fill_1 FILLER_53_837 ();
 sg13g2_decap_4 FILLER_53_842 ();
 sg13g2_fill_2 FILLER_53_846 ();
 sg13g2_decap_8 FILLER_53_852 ();
 sg13g2_decap_8 FILLER_53_859 ();
 sg13g2_decap_8 FILLER_53_866 ();
 sg13g2_decap_4 FILLER_53_873 ();
 sg13g2_decap_4 FILLER_53_884 ();
 sg13g2_fill_1 FILLER_53_888 ();
 sg13g2_decap_8 FILLER_53_898 ();
 sg13g2_decap_8 FILLER_53_905 ();
 sg13g2_decap_8 FILLER_53_912 ();
 sg13g2_fill_2 FILLER_53_919 ();
 sg13g2_fill_1 FILLER_53_921 ();
 sg13g2_decap_4 FILLER_53_940 ();
 sg13g2_fill_1 FILLER_53_948 ();
 sg13g2_fill_2 FILLER_53_953 ();
 sg13g2_fill_2 FILLER_53_959 ();
 sg13g2_fill_1 FILLER_53_968 ();
 sg13g2_fill_2 FILLER_53_972 ();
 sg13g2_fill_1 FILLER_53_974 ();
 sg13g2_decap_8 FILLER_53_980 ();
 sg13g2_decap_4 FILLER_53_987 ();
 sg13g2_fill_2 FILLER_53_1011 ();
 sg13g2_fill_1 FILLER_53_1013 ();
 sg13g2_decap_8 FILLER_53_1018 ();
 sg13g2_decap_8 FILLER_53_1025 ();
 sg13g2_decap_4 FILLER_53_1032 ();
 sg13g2_fill_2 FILLER_53_1036 ();
 sg13g2_fill_2 FILLER_53_1047 ();
 sg13g2_fill_2 FILLER_53_1058 ();
 sg13g2_decap_8 FILLER_53_1069 ();
 sg13g2_decap_8 FILLER_53_1076 ();
 sg13g2_decap_8 FILLER_53_1083 ();
 sg13g2_decap_8 FILLER_53_1090 ();
 sg13g2_decap_8 FILLER_53_1097 ();
 sg13g2_decap_4 FILLER_53_1104 ();
 sg13g2_fill_2 FILLER_53_1108 ();
 sg13g2_decap_8 FILLER_53_1114 ();
 sg13g2_decap_8 FILLER_53_1121 ();
 sg13g2_decap_8 FILLER_53_1128 ();
 sg13g2_decap_8 FILLER_53_1151 ();
 sg13g2_decap_8 FILLER_53_1158 ();
 sg13g2_fill_1 FILLER_53_1165 ();
 sg13g2_decap_8 FILLER_53_1172 ();
 sg13g2_decap_8 FILLER_53_1179 ();
 sg13g2_fill_2 FILLER_53_1191 ();
 sg13g2_fill_1 FILLER_53_1197 ();
 sg13g2_fill_2 FILLER_53_1209 ();
 sg13g2_fill_1 FILLER_53_1211 ();
 sg13g2_decap_4 FILLER_53_1217 ();
 sg13g2_fill_1 FILLER_53_1221 ();
 sg13g2_fill_1 FILLER_53_1235 ();
 sg13g2_fill_2 FILLER_53_1245 ();
 sg13g2_fill_1 FILLER_53_1247 ();
 sg13g2_decap_8 FILLER_53_1253 ();
 sg13g2_decap_4 FILLER_53_1260 ();
 sg13g2_fill_2 FILLER_53_1264 ();
 sg13g2_fill_1 FILLER_53_1274 ();
 sg13g2_decap_8 FILLER_53_1289 ();
 sg13g2_decap_8 FILLER_53_1296 ();
 sg13g2_decap_8 FILLER_53_1303 ();
 sg13g2_decap_8 FILLER_53_1310 ();
 sg13g2_decap_8 FILLER_53_1317 ();
 sg13g2_fill_2 FILLER_53_1324 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_61 ();
 sg13g2_decap_8 FILLER_54_68 ();
 sg13g2_decap_8 FILLER_54_75 ();
 sg13g2_decap_8 FILLER_54_82 ();
 sg13g2_fill_2 FILLER_54_89 ();
 sg13g2_decap_4 FILLER_54_95 ();
 sg13g2_fill_1 FILLER_54_108 ();
 sg13g2_decap_8 FILLER_54_114 ();
 sg13g2_decap_8 FILLER_54_121 ();
 sg13g2_decap_4 FILLER_54_128 ();
 sg13g2_fill_1 FILLER_54_132 ();
 sg13g2_decap_8 FILLER_54_138 ();
 sg13g2_decap_8 FILLER_54_145 ();
 sg13g2_decap_8 FILLER_54_152 ();
 sg13g2_decap_8 FILLER_54_159 ();
 sg13g2_decap_4 FILLER_54_166 ();
 sg13g2_decap_8 FILLER_54_178 ();
 sg13g2_fill_1 FILLER_54_185 ();
 sg13g2_fill_2 FILLER_54_201 ();
 sg13g2_fill_1 FILLER_54_203 ();
 sg13g2_decap_4 FILLER_54_208 ();
 sg13g2_fill_2 FILLER_54_212 ();
 sg13g2_decap_8 FILLER_54_222 ();
 sg13g2_decap_8 FILLER_54_229 ();
 sg13g2_fill_2 FILLER_54_236 ();
 sg13g2_fill_1 FILLER_54_243 ();
 sg13g2_decap_8 FILLER_54_253 ();
 sg13g2_decap_4 FILLER_54_260 ();
 sg13g2_fill_2 FILLER_54_264 ();
 sg13g2_decap_8 FILLER_54_271 ();
 sg13g2_decap_8 FILLER_54_278 ();
 sg13g2_decap_8 FILLER_54_285 ();
 sg13g2_decap_8 FILLER_54_292 ();
 sg13g2_decap_8 FILLER_54_299 ();
 sg13g2_fill_1 FILLER_54_306 ();
 sg13g2_fill_2 FILLER_54_319 ();
 sg13g2_decap_8 FILLER_54_330 ();
 sg13g2_decap_4 FILLER_54_337 ();
 sg13g2_fill_2 FILLER_54_346 ();
 sg13g2_fill_1 FILLER_54_348 ();
 sg13g2_decap_8 FILLER_54_353 ();
 sg13g2_decap_8 FILLER_54_360 ();
 sg13g2_decap_8 FILLER_54_367 ();
 sg13g2_decap_8 FILLER_54_445 ();
 sg13g2_decap_4 FILLER_54_452 ();
 sg13g2_fill_2 FILLER_54_456 ();
 sg13g2_decap_8 FILLER_54_462 ();
 sg13g2_decap_8 FILLER_54_469 ();
 sg13g2_decap_8 FILLER_54_476 ();
 sg13g2_decap_8 FILLER_54_483 ();
 sg13g2_decap_8 FILLER_54_495 ();
 sg13g2_fill_1 FILLER_54_507 ();
 sg13g2_decap_8 FILLER_54_512 ();
 sg13g2_fill_2 FILLER_54_519 ();
 sg13g2_fill_1 FILLER_54_521 ();
 sg13g2_decap_8 FILLER_54_526 ();
 sg13g2_fill_1 FILLER_54_533 ();
 sg13g2_decap_4 FILLER_54_539 ();
 sg13g2_fill_2 FILLER_54_543 ();
 sg13g2_decap_8 FILLER_54_549 ();
 sg13g2_decap_4 FILLER_54_556 ();
 sg13g2_fill_1 FILLER_54_560 ();
 sg13g2_decap_4 FILLER_54_566 ();
 sg13g2_decap_8 FILLER_54_574 ();
 sg13g2_fill_2 FILLER_54_581 ();
 sg13g2_fill_1 FILLER_54_583 ();
 sg13g2_decap_8 FILLER_54_588 ();
 sg13g2_decap_8 FILLER_54_595 ();
 sg13g2_decap_8 FILLER_54_602 ();
 sg13g2_decap_8 FILLER_54_609 ();
 sg13g2_decap_8 FILLER_54_616 ();
 sg13g2_decap_8 FILLER_54_623 ();
 sg13g2_decap_4 FILLER_54_630 ();
 sg13g2_fill_2 FILLER_54_634 ();
 sg13g2_decap_4 FILLER_54_643 ();
 sg13g2_decap_8 FILLER_54_658 ();
 sg13g2_decap_8 FILLER_54_665 ();
 sg13g2_decap_8 FILLER_54_672 ();
 sg13g2_decap_8 FILLER_54_679 ();
 sg13g2_decap_8 FILLER_54_690 ();
 sg13g2_decap_8 FILLER_54_697 ();
 sg13g2_fill_2 FILLER_54_704 ();
 sg13g2_fill_1 FILLER_54_706 ();
 sg13g2_decap_8 FILLER_54_711 ();
 sg13g2_decap_8 FILLER_54_718 ();
 sg13g2_decap_8 FILLER_54_725 ();
 sg13g2_fill_2 FILLER_54_732 ();
 sg13g2_fill_1 FILLER_54_734 ();
 sg13g2_decap_8 FILLER_54_744 ();
 sg13g2_decap_8 FILLER_54_751 ();
 sg13g2_decap_8 FILLER_54_758 ();
 sg13g2_decap_8 FILLER_54_765 ();
 sg13g2_fill_2 FILLER_54_772 ();
 sg13g2_fill_1 FILLER_54_774 ();
 sg13g2_decap_4 FILLER_54_780 ();
 sg13g2_fill_1 FILLER_54_784 ();
 sg13g2_decap_8 FILLER_54_788 ();
 sg13g2_decap_8 FILLER_54_795 ();
 sg13g2_fill_2 FILLER_54_802 ();
 sg13g2_decap_8 FILLER_54_809 ();
 sg13g2_fill_1 FILLER_54_816 ();
 sg13g2_decap_8 FILLER_54_821 ();
 sg13g2_decap_8 FILLER_54_828 ();
 sg13g2_decap_8 FILLER_54_835 ();
 sg13g2_decap_8 FILLER_54_842 ();
 sg13g2_decap_8 FILLER_54_849 ();
 sg13g2_fill_2 FILLER_54_860 ();
 sg13g2_decap_8 FILLER_54_866 ();
 sg13g2_decap_4 FILLER_54_873 ();
 sg13g2_fill_2 FILLER_54_877 ();
 sg13g2_fill_2 FILLER_54_883 ();
 sg13g2_decap_4 FILLER_54_889 ();
 sg13g2_decap_4 FILLER_54_897 ();
 sg13g2_decap_4 FILLER_54_905 ();
 sg13g2_decap_8 FILLER_54_914 ();
 sg13g2_fill_2 FILLER_54_921 ();
 sg13g2_fill_1 FILLER_54_923 ();
 sg13g2_decap_8 FILLER_54_934 ();
 sg13g2_decap_8 FILLER_54_941 ();
 sg13g2_decap_8 FILLER_54_948 ();
 sg13g2_decap_8 FILLER_54_955 ();
 sg13g2_decap_4 FILLER_54_962 ();
 sg13g2_fill_1 FILLER_54_966 ();
 sg13g2_decap_4 FILLER_54_982 ();
 sg13g2_fill_1 FILLER_54_986 ();
 sg13g2_decap_8 FILLER_54_993 ();
 sg13g2_decap_4 FILLER_54_1000 ();
 sg13g2_fill_1 FILLER_54_1004 ();
 sg13g2_decap_8 FILLER_54_1022 ();
 sg13g2_decap_8 FILLER_54_1029 ();
 sg13g2_decap_8 FILLER_54_1036 ();
 sg13g2_decap_8 FILLER_54_1043 ();
 sg13g2_decap_4 FILLER_54_1050 ();
 sg13g2_fill_1 FILLER_54_1054 ();
 sg13g2_decap_8 FILLER_54_1059 ();
 sg13g2_decap_8 FILLER_54_1066 ();
 sg13g2_decap_8 FILLER_54_1073 ();
 sg13g2_decap_8 FILLER_54_1080 ();
 sg13g2_decap_8 FILLER_54_1087 ();
 sg13g2_decap_4 FILLER_54_1094 ();
 sg13g2_fill_2 FILLER_54_1098 ();
 sg13g2_decap_4 FILLER_54_1116 ();
 sg13g2_fill_2 FILLER_54_1120 ();
 sg13g2_fill_2 FILLER_54_1146 ();
 sg13g2_fill_1 FILLER_54_1148 ();
 sg13g2_decap_8 FILLER_54_1153 ();
 sg13g2_fill_2 FILLER_54_1160 ();
 sg13g2_fill_1 FILLER_54_1162 ();
 sg13g2_decap_8 FILLER_54_1167 ();
 sg13g2_decap_4 FILLER_54_1174 ();
 sg13g2_decap_4 FILLER_54_1193 ();
 sg13g2_fill_2 FILLER_54_1197 ();
 sg13g2_fill_2 FILLER_54_1204 ();
 sg13g2_decap_8 FILLER_54_1214 ();
 sg13g2_decap_8 FILLER_54_1221 ();
 sg13g2_decap_4 FILLER_54_1228 ();
 sg13g2_decap_4 FILLER_54_1241 ();
 sg13g2_fill_1 FILLER_54_1245 ();
 sg13g2_decap_4 FILLER_54_1250 ();
 sg13g2_decap_4 FILLER_54_1263 ();
 sg13g2_fill_2 FILLER_54_1273 ();
 sg13g2_fill_1 FILLER_54_1280 ();
 sg13g2_fill_2 FILLER_54_1286 ();
 sg13g2_fill_1 FILLER_54_1288 ();
 sg13g2_decap_8 FILLER_54_1294 ();
 sg13g2_decap_8 FILLER_54_1301 ();
 sg13g2_decap_8 FILLER_54_1308 ();
 sg13g2_decap_8 FILLER_54_1315 ();
 sg13g2_decap_4 FILLER_54_1322 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_fill_2 FILLER_55_21 ();
 sg13g2_fill_1 FILLER_55_23 ();
 sg13g2_fill_2 FILLER_55_55 ();
 sg13g2_fill_1 FILLER_55_57 ();
 sg13g2_decap_8 FILLER_55_64 ();
 sg13g2_decap_8 FILLER_55_71 ();
 sg13g2_decap_8 FILLER_55_78 ();
 sg13g2_decap_8 FILLER_55_85 ();
 sg13g2_fill_2 FILLER_55_92 ();
 sg13g2_fill_1 FILLER_55_115 ();
 sg13g2_fill_1 FILLER_55_122 ();
 sg13g2_decap_8 FILLER_55_127 ();
 sg13g2_decap_8 FILLER_55_134 ();
 sg13g2_decap_8 FILLER_55_141 ();
 sg13g2_fill_1 FILLER_55_148 ();
 sg13g2_fill_2 FILLER_55_158 ();
 sg13g2_fill_1 FILLER_55_169 ();
 sg13g2_fill_2 FILLER_55_209 ();
 sg13g2_fill_2 FILLER_55_216 ();
 sg13g2_decap_4 FILLER_55_223 ();
 sg13g2_decap_4 FILLER_55_232 ();
 sg13g2_decap_4 FILLER_55_241 ();
 sg13g2_decap_8 FILLER_55_254 ();
 sg13g2_decap_4 FILLER_55_261 ();
 sg13g2_fill_1 FILLER_55_265 ();
 sg13g2_fill_2 FILLER_55_271 ();
 sg13g2_fill_1 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_279 ();
 sg13g2_decap_8 FILLER_55_286 ();
 sg13g2_decap_8 FILLER_55_293 ();
 sg13g2_decap_8 FILLER_55_300 ();
 sg13g2_decap_8 FILLER_55_307 ();
 sg13g2_decap_8 FILLER_55_314 ();
 sg13g2_decap_8 FILLER_55_326 ();
 sg13g2_decap_8 FILLER_55_333 ();
 sg13g2_decap_4 FILLER_55_340 ();
 sg13g2_decap_8 FILLER_55_349 ();
 sg13g2_fill_2 FILLER_55_356 ();
 sg13g2_fill_1 FILLER_55_358 ();
 sg13g2_decap_8 FILLER_55_364 ();
 sg13g2_fill_2 FILLER_55_371 ();
 sg13g2_fill_1 FILLER_55_373 ();
 sg13g2_decap_8 FILLER_55_379 ();
 sg13g2_fill_2 FILLER_55_386 ();
 sg13g2_fill_1 FILLER_55_388 ();
 sg13g2_fill_2 FILLER_55_393 ();
 sg13g2_decap_8 FILLER_55_399 ();
 sg13g2_decap_8 FILLER_55_406 ();
 sg13g2_decap_8 FILLER_55_413 ();
 sg13g2_decap_8 FILLER_55_420 ();
 sg13g2_decap_8 FILLER_55_427 ();
 sg13g2_decap_4 FILLER_55_434 ();
 sg13g2_decap_8 FILLER_55_447 ();
 sg13g2_decap_8 FILLER_55_454 ();
 sg13g2_decap_8 FILLER_55_461 ();
 sg13g2_decap_8 FILLER_55_468 ();
 sg13g2_fill_1 FILLER_55_475 ();
 sg13g2_decap_8 FILLER_55_491 ();
 sg13g2_decap_8 FILLER_55_498 ();
 sg13g2_decap_8 FILLER_55_505 ();
 sg13g2_decap_8 FILLER_55_512 ();
 sg13g2_decap_8 FILLER_55_519 ();
 sg13g2_decap_8 FILLER_55_526 ();
 sg13g2_decap_4 FILLER_55_533 ();
 sg13g2_fill_1 FILLER_55_537 ();
 sg13g2_fill_2 FILLER_55_590 ();
 sg13g2_fill_1 FILLER_55_592 ();
 sg13g2_fill_1 FILLER_55_645 ();
 sg13g2_fill_2 FILLER_55_667 ();
 sg13g2_fill_1 FILLER_55_669 ();
 sg13g2_decap_8 FILLER_55_703 ();
 sg13g2_decap_8 FILLER_55_710 ();
 sg13g2_decap_4 FILLER_55_717 ();
 sg13g2_fill_1 FILLER_55_721 ();
 sg13g2_decap_8 FILLER_55_730 ();
 sg13g2_fill_1 FILLER_55_742 ();
 sg13g2_decap_8 FILLER_55_751 ();
 sg13g2_decap_4 FILLER_55_758 ();
 sg13g2_fill_2 FILLER_55_762 ();
 sg13g2_decap_4 FILLER_55_773 ();
 sg13g2_fill_2 FILLER_55_781 ();
 sg13g2_fill_1 FILLER_55_783 ();
 sg13g2_decap_8 FILLER_55_794 ();
 sg13g2_decap_8 FILLER_55_801 ();
 sg13g2_decap_8 FILLER_55_808 ();
 sg13g2_decap_8 FILLER_55_815 ();
 sg13g2_decap_8 FILLER_55_822 ();
 sg13g2_decap_8 FILLER_55_829 ();
 sg13g2_decap_8 FILLER_55_836 ();
 sg13g2_decap_8 FILLER_55_843 ();
 sg13g2_decap_8 FILLER_55_850 ();
 sg13g2_decap_8 FILLER_55_857 ();
 sg13g2_decap_8 FILLER_55_864 ();
 sg13g2_decap_8 FILLER_55_871 ();
 sg13g2_decap_8 FILLER_55_878 ();
 sg13g2_decap_4 FILLER_55_885 ();
 sg13g2_fill_2 FILLER_55_889 ();
 sg13g2_fill_1 FILLER_55_896 ();
 sg13g2_decap_4 FILLER_55_902 ();
 sg13g2_fill_1 FILLER_55_906 ();
 sg13g2_decap_4 FILLER_55_920 ();
 sg13g2_fill_1 FILLER_55_938 ();
 sg13g2_decap_8 FILLER_55_953 ();
 sg13g2_decap_4 FILLER_55_960 ();
 sg13g2_decap_8 FILLER_55_983 ();
 sg13g2_decap_4 FILLER_55_990 ();
 sg13g2_decap_4 FILLER_55_999 ();
 sg13g2_fill_2 FILLER_55_1003 ();
 sg13g2_decap_8 FILLER_55_1009 ();
 sg13g2_fill_2 FILLER_55_1016 ();
 sg13g2_decap_8 FILLER_55_1023 ();
 sg13g2_decap_4 FILLER_55_1036 ();
 sg13g2_fill_2 FILLER_55_1040 ();
 sg13g2_fill_2 FILLER_55_1050 ();
 sg13g2_decap_8 FILLER_55_1057 ();
 sg13g2_fill_1 FILLER_55_1070 ();
 sg13g2_fill_2 FILLER_55_1081 ();
 sg13g2_decap_8 FILLER_55_1102 ();
 sg13g2_decap_8 FILLER_55_1109 ();
 sg13g2_decap_4 FILLER_55_1116 ();
 sg13g2_fill_2 FILLER_55_1120 ();
 sg13g2_decap_8 FILLER_55_1133 ();
 sg13g2_decap_4 FILLER_55_1140 ();
 sg13g2_decap_8 FILLER_55_1150 ();
 sg13g2_decap_4 FILLER_55_1157 ();
 sg13g2_fill_1 FILLER_55_1161 ();
 sg13g2_decap_8 FILLER_55_1167 ();
 sg13g2_decap_8 FILLER_55_1174 ();
 sg13g2_decap_4 FILLER_55_1181 ();
 sg13g2_fill_1 FILLER_55_1185 ();
 sg13g2_fill_2 FILLER_55_1194 ();
 sg13g2_fill_1 FILLER_55_1196 ();
 sg13g2_fill_2 FILLER_55_1202 ();
 sg13g2_decap_8 FILLER_55_1210 ();
 sg13g2_decap_8 FILLER_55_1217 ();
 sg13g2_fill_2 FILLER_55_1224 ();
 sg13g2_fill_1 FILLER_55_1226 ();
 sg13g2_decap_8 FILLER_55_1231 ();
 sg13g2_decap_8 FILLER_55_1238 ();
 sg13g2_decap_8 FILLER_55_1245 ();
 sg13g2_fill_2 FILLER_55_1252 ();
 sg13g2_decap_4 FILLER_55_1260 ();
 sg13g2_decap_4 FILLER_55_1269 ();
 sg13g2_fill_2 FILLER_55_1273 ();
 sg13g2_decap_8 FILLER_55_1279 ();
 sg13g2_decap_8 FILLER_55_1286 ();
 sg13g2_decap_8 FILLER_55_1293 ();
 sg13g2_decap_8 FILLER_55_1300 ();
 sg13g2_decap_8 FILLER_55_1307 ();
 sg13g2_decap_8 FILLER_55_1314 ();
 sg13g2_decap_4 FILLER_55_1321 ();
 sg13g2_fill_1 FILLER_55_1325 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_fill_2 FILLER_56_35 ();
 sg13g2_fill_1 FILLER_56_37 ();
 sg13g2_fill_2 FILLER_56_64 ();
 sg13g2_fill_1 FILLER_56_66 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_4 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_115 ();
 sg13g2_decap_8 FILLER_56_122 ();
 sg13g2_decap_8 FILLER_56_129 ();
 sg13g2_decap_8 FILLER_56_136 ();
 sg13g2_fill_2 FILLER_56_143 ();
 sg13g2_fill_1 FILLER_56_145 ();
 sg13g2_fill_2 FILLER_56_153 ();
 sg13g2_fill_1 FILLER_56_155 ();
 sg13g2_decap_8 FILLER_56_165 ();
 sg13g2_fill_2 FILLER_56_172 ();
 sg13g2_decap_8 FILLER_56_179 ();
 sg13g2_fill_1 FILLER_56_186 ();
 sg13g2_fill_1 FILLER_56_191 ();
 sg13g2_fill_1 FILLER_56_222 ();
 sg13g2_decap_8 FILLER_56_227 ();
 sg13g2_decap_8 FILLER_56_234 ();
 sg13g2_decap_8 FILLER_56_241 ();
 sg13g2_decap_8 FILLER_56_248 ();
 sg13g2_decap_8 FILLER_56_255 ();
 sg13g2_decap_8 FILLER_56_262 ();
 sg13g2_decap_8 FILLER_56_269 ();
 sg13g2_decap_8 FILLER_56_276 ();
 sg13g2_decap_8 FILLER_56_287 ();
 sg13g2_decap_8 FILLER_56_294 ();
 sg13g2_decap_8 FILLER_56_301 ();
 sg13g2_decap_4 FILLER_56_308 ();
 sg13g2_fill_2 FILLER_56_316 ();
 sg13g2_decap_8 FILLER_56_326 ();
 sg13g2_decap_8 FILLER_56_333 ();
 sg13g2_decap_8 FILLER_56_340 ();
 sg13g2_decap_8 FILLER_56_347 ();
 sg13g2_decap_8 FILLER_56_354 ();
 sg13g2_decap_8 FILLER_56_361 ();
 sg13g2_fill_2 FILLER_56_368 ();
 sg13g2_decap_8 FILLER_56_375 ();
 sg13g2_decap_8 FILLER_56_382 ();
 sg13g2_decap_8 FILLER_56_389 ();
 sg13g2_decap_8 FILLER_56_396 ();
 sg13g2_decap_8 FILLER_56_403 ();
 sg13g2_decap_4 FILLER_56_410 ();
 sg13g2_fill_1 FILLER_56_414 ();
 sg13g2_decap_4 FILLER_56_420 ();
 sg13g2_fill_2 FILLER_56_424 ();
 sg13g2_decap_8 FILLER_56_441 ();
 sg13g2_fill_2 FILLER_56_448 ();
 sg13g2_decap_8 FILLER_56_454 ();
 sg13g2_fill_2 FILLER_56_461 ();
 sg13g2_decap_4 FILLER_56_467 ();
 sg13g2_fill_1 FILLER_56_471 ();
 sg13g2_decap_8 FILLER_56_477 ();
 sg13g2_decap_4 FILLER_56_484 ();
 sg13g2_decap_8 FILLER_56_493 ();
 sg13g2_decap_8 FILLER_56_500 ();
 sg13g2_decap_8 FILLER_56_507 ();
 sg13g2_decap_8 FILLER_56_514 ();
 sg13g2_decap_8 FILLER_56_521 ();
 sg13g2_decap_8 FILLER_56_533 ();
 sg13g2_decap_8 FILLER_56_540 ();
 sg13g2_fill_2 FILLER_56_547 ();
 sg13g2_fill_1 FILLER_56_549 ();
 sg13g2_decap_8 FILLER_56_558 ();
 sg13g2_decap_8 FILLER_56_565 ();
 sg13g2_decap_8 FILLER_56_572 ();
 sg13g2_decap_8 FILLER_56_579 ();
 sg13g2_decap_8 FILLER_56_586 ();
 sg13g2_decap_8 FILLER_56_593 ();
 sg13g2_fill_2 FILLER_56_600 ();
 sg13g2_decap_4 FILLER_56_606 ();
 sg13g2_fill_2 FILLER_56_610 ();
 sg13g2_fill_2 FILLER_56_619 ();
 sg13g2_fill_1 FILLER_56_621 ();
 sg13g2_fill_1 FILLER_56_627 ();
 sg13g2_fill_2 FILLER_56_632 ();
 sg13g2_fill_1 FILLER_56_634 ();
 sg13g2_decap_8 FILLER_56_640 ();
 sg13g2_decap_8 FILLER_56_647 ();
 sg13g2_decap_8 FILLER_56_654 ();
 sg13g2_decap_8 FILLER_56_661 ();
 sg13g2_decap_8 FILLER_56_668 ();
 sg13g2_decap_8 FILLER_56_675 ();
 sg13g2_decap_4 FILLER_56_682 ();
 sg13g2_fill_2 FILLER_56_686 ();
 sg13g2_decap_4 FILLER_56_735 ();
 sg13g2_fill_2 FILLER_56_770 ();
 sg13g2_fill_1 FILLER_56_772 ();
 sg13g2_fill_1 FILLER_56_777 ();
 sg13g2_decap_8 FILLER_56_813 ();
 sg13g2_decap_8 FILLER_56_820 ();
 sg13g2_decap_8 FILLER_56_827 ();
 sg13g2_decap_8 FILLER_56_834 ();
 sg13g2_decap_8 FILLER_56_841 ();
 sg13g2_decap_8 FILLER_56_848 ();
 sg13g2_decap_8 FILLER_56_855 ();
 sg13g2_decap_8 FILLER_56_862 ();
 sg13g2_decap_8 FILLER_56_869 ();
 sg13g2_decap_8 FILLER_56_876 ();
 sg13g2_decap_8 FILLER_56_883 ();
 sg13g2_decap_8 FILLER_56_890 ();
 sg13g2_decap_8 FILLER_56_897 ();
 sg13g2_fill_2 FILLER_56_904 ();
 sg13g2_decap_4 FILLER_56_911 ();
 sg13g2_fill_1 FILLER_56_937 ();
 sg13g2_fill_2 FILLER_56_943 ();
 sg13g2_decap_8 FILLER_56_958 ();
 sg13g2_decap_4 FILLER_56_965 ();
 sg13g2_fill_1 FILLER_56_969 ();
 sg13g2_fill_1 FILLER_56_975 ();
 sg13g2_decap_4 FILLER_56_982 ();
 sg13g2_fill_2 FILLER_56_986 ();
 sg13g2_decap_8 FILLER_56_992 ();
 sg13g2_decap_8 FILLER_56_999 ();
 sg13g2_decap_8 FILLER_56_1006 ();
 sg13g2_fill_2 FILLER_56_1013 ();
 sg13g2_fill_1 FILLER_56_1015 ();
 sg13g2_decap_8 FILLER_56_1020 ();
 sg13g2_decap_8 FILLER_56_1032 ();
 sg13g2_decap_8 FILLER_56_1039 ();
 sg13g2_decap_4 FILLER_56_1046 ();
 sg13g2_fill_1 FILLER_56_1050 ();
 sg13g2_fill_2 FILLER_56_1056 ();
 sg13g2_decap_8 FILLER_56_1063 ();
 sg13g2_decap_8 FILLER_56_1070 ();
 sg13g2_decap_8 FILLER_56_1077 ();
 sg13g2_decap_8 FILLER_56_1084 ();
 sg13g2_decap_4 FILLER_56_1091 ();
 sg13g2_decap_8 FILLER_56_1100 ();
 sg13g2_decap_8 FILLER_56_1107 ();
 sg13g2_fill_2 FILLER_56_1114 ();
 sg13g2_decap_8 FILLER_56_1121 ();
 sg13g2_decap_8 FILLER_56_1128 ();
 sg13g2_fill_2 FILLER_56_1135 ();
 sg13g2_fill_1 FILLER_56_1137 ();
 sg13g2_fill_1 FILLER_56_1142 ();
 sg13g2_fill_2 FILLER_56_1148 ();
 sg13g2_decap_8 FILLER_56_1158 ();
 sg13g2_fill_1 FILLER_56_1170 ();
 sg13g2_decap_8 FILLER_56_1181 ();
 sg13g2_decap_8 FILLER_56_1188 ();
 sg13g2_fill_2 FILLER_56_1195 ();
 sg13g2_decap_8 FILLER_56_1204 ();
 sg13g2_decap_8 FILLER_56_1211 ();
 sg13g2_decap_8 FILLER_56_1218 ();
 sg13g2_decap_4 FILLER_56_1225 ();
 sg13g2_fill_1 FILLER_56_1229 ();
 sg13g2_decap_8 FILLER_56_1234 ();
 sg13g2_decap_4 FILLER_56_1241 ();
 sg13g2_fill_1 FILLER_56_1245 ();
 sg13g2_decap_8 FILLER_56_1254 ();
 sg13g2_decap_8 FILLER_56_1261 ();
 sg13g2_decap_8 FILLER_56_1268 ();
 sg13g2_decap_8 FILLER_56_1275 ();
 sg13g2_decap_8 FILLER_56_1282 ();
 sg13g2_decap_8 FILLER_56_1289 ();
 sg13g2_decap_8 FILLER_56_1296 ();
 sg13g2_decap_8 FILLER_56_1303 ();
 sg13g2_decap_8 FILLER_56_1310 ();
 sg13g2_decap_8 FILLER_56_1317 ();
 sg13g2_fill_2 FILLER_56_1324 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_fill_2 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_42 ();
 sg13g2_fill_1 FILLER_57_61 ();
 sg13g2_fill_2 FILLER_57_67 ();
 sg13g2_fill_1 FILLER_57_69 ();
 sg13g2_fill_1 FILLER_57_75 ();
 sg13g2_decap_8 FILLER_57_88 ();
 sg13g2_fill_2 FILLER_57_95 ();
 sg13g2_fill_1 FILLER_57_97 ();
 sg13g2_decap_4 FILLER_57_103 ();
 sg13g2_fill_2 FILLER_57_107 ();
 sg13g2_decap_8 FILLER_57_113 ();
 sg13g2_decap_8 FILLER_57_120 ();
 sg13g2_decap_8 FILLER_57_127 ();
 sg13g2_decap_8 FILLER_57_134 ();
 sg13g2_fill_2 FILLER_57_141 ();
 sg13g2_fill_1 FILLER_57_143 ();
 sg13g2_decap_8 FILLER_57_149 ();
 sg13g2_decap_8 FILLER_57_156 ();
 sg13g2_decap_8 FILLER_57_163 ();
 sg13g2_decap_8 FILLER_57_170 ();
 sg13g2_decap_4 FILLER_57_177 ();
 sg13g2_fill_1 FILLER_57_181 ();
 sg13g2_decap_8 FILLER_57_188 ();
 sg13g2_fill_1 FILLER_57_195 ();
 sg13g2_decap_4 FILLER_57_211 ();
 sg13g2_fill_1 FILLER_57_231 ();
 sg13g2_decap_8 FILLER_57_237 ();
 sg13g2_decap_8 FILLER_57_244 ();
 sg13g2_decap_8 FILLER_57_251 ();
 sg13g2_decap_4 FILLER_57_258 ();
 sg13g2_fill_1 FILLER_57_262 ();
 sg13g2_fill_1 FILLER_57_268 ();
 sg13g2_decap_8 FILLER_57_278 ();
 sg13g2_fill_2 FILLER_57_285 ();
 sg13g2_fill_1 FILLER_57_287 ();
 sg13g2_decap_8 FILLER_57_293 ();
 sg13g2_decap_8 FILLER_57_305 ();
 sg13g2_fill_1 FILLER_57_312 ();
 sg13g2_decap_8 FILLER_57_323 ();
 sg13g2_decap_4 FILLER_57_333 ();
 sg13g2_decap_8 FILLER_57_342 ();
 sg13g2_decap_8 FILLER_57_349 ();
 sg13g2_decap_8 FILLER_57_356 ();
 sg13g2_fill_2 FILLER_57_363 ();
 sg13g2_decap_8 FILLER_57_399 ();
 sg13g2_decap_4 FILLER_57_406 ();
 sg13g2_fill_1 FILLER_57_410 ();
 sg13g2_fill_1 FILLER_57_416 ();
 sg13g2_decap_8 FILLER_57_422 ();
 sg13g2_decap_8 FILLER_57_429 ();
 sg13g2_decap_8 FILLER_57_436 ();
 sg13g2_fill_2 FILLER_57_443 ();
 sg13g2_fill_1 FILLER_57_445 ();
 sg13g2_decap_4 FILLER_57_450 ();
 sg13g2_decap_8 FILLER_57_459 ();
 sg13g2_decap_8 FILLER_57_466 ();
 sg13g2_decap_8 FILLER_57_473 ();
 sg13g2_decap_4 FILLER_57_480 ();
 sg13g2_fill_1 FILLER_57_484 ();
 sg13g2_fill_2 FILLER_57_489 ();
 sg13g2_fill_1 FILLER_57_491 ();
 sg13g2_decap_4 FILLER_57_496 ();
 sg13g2_fill_2 FILLER_57_500 ();
 sg13g2_decap_8 FILLER_57_515 ();
 sg13g2_decap_8 FILLER_57_522 ();
 sg13g2_decap_8 FILLER_57_529 ();
 sg13g2_decap_8 FILLER_57_536 ();
 sg13g2_decap_8 FILLER_57_543 ();
 sg13g2_decap_8 FILLER_57_550 ();
 sg13g2_decap_8 FILLER_57_557 ();
 sg13g2_decap_8 FILLER_57_564 ();
 sg13g2_decap_8 FILLER_57_571 ();
 sg13g2_decap_4 FILLER_57_578 ();
 sg13g2_decap_8 FILLER_57_586 ();
 sg13g2_decap_8 FILLER_57_593 ();
 sg13g2_decap_8 FILLER_57_600 ();
 sg13g2_decap_8 FILLER_57_607 ();
 sg13g2_decap_8 FILLER_57_614 ();
 sg13g2_decap_4 FILLER_57_621 ();
 sg13g2_fill_1 FILLER_57_625 ();
 sg13g2_decap_8 FILLER_57_630 ();
 sg13g2_decap_8 FILLER_57_641 ();
 sg13g2_decap_8 FILLER_57_652 ();
 sg13g2_decap_8 FILLER_57_659 ();
 sg13g2_decap_8 FILLER_57_666 ();
 sg13g2_fill_2 FILLER_57_677 ();
 sg13g2_decap_4 FILLER_57_684 ();
 sg13g2_decap_8 FILLER_57_692 ();
 sg13g2_decap_8 FILLER_57_699 ();
 sg13g2_decap_8 FILLER_57_706 ();
 sg13g2_decap_8 FILLER_57_713 ();
 sg13g2_decap_8 FILLER_57_720 ();
 sg13g2_decap_4 FILLER_57_727 ();
 sg13g2_fill_2 FILLER_57_731 ();
 sg13g2_decap_8 FILLER_57_746 ();
 sg13g2_decap_8 FILLER_57_753 ();
 sg13g2_decap_8 FILLER_57_760 ();
 sg13g2_decap_4 FILLER_57_767 ();
 sg13g2_fill_1 FILLER_57_771 ();
 sg13g2_fill_2 FILLER_57_777 ();
 sg13g2_fill_1 FILLER_57_787 ();
 sg13g2_decap_8 FILLER_57_809 ();
 sg13g2_decap_4 FILLER_57_816 ();
 sg13g2_fill_1 FILLER_57_820 ();
 sg13g2_decap_4 FILLER_57_826 ();
 sg13g2_fill_2 FILLER_57_830 ();
 sg13g2_fill_1 FILLER_57_836 ();
 sg13g2_decap_8 FILLER_57_843 ();
 sg13g2_decap_8 FILLER_57_850 ();
 sg13g2_decap_4 FILLER_57_857 ();
 sg13g2_decap_8 FILLER_57_865 ();
 sg13g2_fill_1 FILLER_57_872 ();
 sg13g2_fill_2 FILLER_57_890 ();
 sg13g2_fill_1 FILLER_57_892 ();
 sg13g2_fill_2 FILLER_57_903 ();
 sg13g2_fill_1 FILLER_57_905 ();
 sg13g2_decap_8 FILLER_57_911 ();
 sg13g2_decap_4 FILLER_57_926 ();
 sg13g2_fill_1 FILLER_57_930 ();
 sg13g2_decap_8 FILLER_57_949 ();
 sg13g2_decap_8 FILLER_57_956 ();
 sg13g2_fill_2 FILLER_57_963 ();
 sg13g2_fill_1 FILLER_57_965 ();
 sg13g2_decap_8 FILLER_57_981 ();
 sg13g2_decap_4 FILLER_57_988 ();
 sg13g2_fill_2 FILLER_57_992 ();
 sg13g2_decap_8 FILLER_57_999 ();
 sg13g2_decap_8 FILLER_57_1006 ();
 sg13g2_fill_2 FILLER_57_1013 ();
 sg13g2_fill_1 FILLER_57_1015 ();
 sg13g2_decap_8 FILLER_57_1022 ();
 sg13g2_decap_8 FILLER_57_1029 ();
 sg13g2_decap_4 FILLER_57_1036 ();
 sg13g2_decap_8 FILLER_57_1045 ();
 sg13g2_decap_8 FILLER_57_1052 ();
 sg13g2_decap_8 FILLER_57_1059 ();
 sg13g2_decap_8 FILLER_57_1066 ();
 sg13g2_decap_8 FILLER_57_1073 ();
 sg13g2_decap_4 FILLER_57_1080 ();
 sg13g2_fill_1 FILLER_57_1084 ();
 sg13g2_decap_8 FILLER_57_1089 ();
 sg13g2_decap_8 FILLER_57_1096 ();
 sg13g2_decap_8 FILLER_57_1103 ();
 sg13g2_decap_4 FILLER_57_1110 ();
 sg13g2_fill_1 FILLER_57_1114 ();
 sg13g2_decap_8 FILLER_57_1125 ();
 sg13g2_decap_8 FILLER_57_1137 ();
 sg13g2_decap_8 FILLER_57_1144 ();
 sg13g2_fill_2 FILLER_57_1157 ();
 sg13g2_fill_1 FILLER_57_1159 ();
 sg13g2_fill_1 FILLER_57_1164 ();
 sg13g2_fill_2 FILLER_57_1177 ();
 sg13g2_fill_1 FILLER_57_1179 ();
 sg13g2_fill_1 FILLER_57_1186 ();
 sg13g2_fill_1 FILLER_57_1192 ();
 sg13g2_decap_8 FILLER_57_1202 ();
 sg13g2_decap_8 FILLER_57_1209 ();
 sg13g2_decap_8 FILLER_57_1216 ();
 sg13g2_decap_8 FILLER_57_1223 ();
 sg13g2_fill_1 FILLER_57_1230 ();
 sg13g2_decap_8 FILLER_57_1245 ();
 sg13g2_decap_8 FILLER_57_1260 ();
 sg13g2_decap_8 FILLER_57_1267 ();
 sg13g2_decap_8 FILLER_57_1274 ();
 sg13g2_decap_8 FILLER_57_1281 ();
 sg13g2_decap_8 FILLER_57_1288 ();
 sg13g2_decap_8 FILLER_57_1295 ();
 sg13g2_decap_8 FILLER_57_1302 ();
 sg13g2_decap_8 FILLER_57_1309 ();
 sg13g2_decap_8 FILLER_57_1316 ();
 sg13g2_fill_2 FILLER_57_1323 ();
 sg13g2_fill_1 FILLER_57_1325 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_fill_2 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_27 ();
 sg13g2_fill_1 FILLER_58_34 ();
 sg13g2_decap_4 FILLER_58_61 ();
 sg13g2_fill_2 FILLER_58_70 ();
 sg13g2_fill_1 FILLER_58_72 ();
 sg13g2_decap_8 FILLER_58_78 ();
 sg13g2_decap_8 FILLER_58_85 ();
 sg13g2_decap_8 FILLER_58_92 ();
 sg13g2_decap_8 FILLER_58_99 ();
 sg13g2_decap_4 FILLER_58_116 ();
 sg13g2_decap_4 FILLER_58_129 ();
 sg13g2_fill_1 FILLER_58_133 ();
 sg13g2_fill_1 FILLER_58_138 ();
 sg13g2_fill_2 FILLER_58_152 ();
 sg13g2_fill_1 FILLER_58_154 ();
 sg13g2_fill_1 FILLER_58_160 ();
 sg13g2_decap_8 FILLER_58_165 ();
 sg13g2_decap_8 FILLER_58_172 ();
 sg13g2_decap_8 FILLER_58_179 ();
 sg13g2_decap_8 FILLER_58_186 ();
 sg13g2_decap_4 FILLER_58_193 ();
 sg13g2_fill_1 FILLER_58_197 ();
 sg13g2_decap_8 FILLER_58_202 ();
 sg13g2_decap_8 FILLER_58_213 ();
 sg13g2_decap_8 FILLER_58_220 ();
 sg13g2_fill_1 FILLER_58_227 ();
 sg13g2_decap_8 FILLER_58_237 ();
 sg13g2_decap_8 FILLER_58_244 ();
 sg13g2_fill_2 FILLER_58_251 ();
 sg13g2_fill_1 FILLER_58_253 ();
 sg13g2_decap_8 FILLER_58_294 ();
 sg13g2_fill_2 FILLER_58_301 ();
 sg13g2_fill_1 FILLER_58_303 ();
 sg13g2_decap_8 FILLER_58_327 ();
 sg13g2_decap_8 FILLER_58_334 ();
 sg13g2_fill_2 FILLER_58_341 ();
 sg13g2_fill_1 FILLER_58_343 ();
 sg13g2_fill_1 FILLER_58_352 ();
 sg13g2_decap_8 FILLER_58_359 ();
 sg13g2_decap_8 FILLER_58_366 ();
 sg13g2_fill_1 FILLER_58_373 ();
 sg13g2_decap_8 FILLER_58_395 ();
 sg13g2_fill_1 FILLER_58_402 ();
 sg13g2_decap_4 FILLER_58_438 ();
 sg13g2_decap_8 FILLER_58_468 ();
 sg13g2_fill_1 FILLER_58_475 ();
 sg13g2_fill_2 FILLER_58_483 ();
 sg13g2_decap_8 FILLER_58_522 ();
 sg13g2_decap_8 FILLER_58_529 ();
 sg13g2_decap_8 FILLER_58_562 ();
 sg13g2_decap_4 FILLER_58_569 ();
 sg13g2_fill_2 FILLER_58_573 ();
 sg13g2_decap_8 FILLER_58_601 ();
 sg13g2_decap_8 FILLER_58_608 ();
 sg13g2_decap_8 FILLER_58_615 ();
 sg13g2_decap_8 FILLER_58_622 ();
 sg13g2_decap_8 FILLER_58_629 ();
 sg13g2_decap_8 FILLER_58_636 ();
 sg13g2_decap_8 FILLER_58_643 ();
 sg13g2_decap_8 FILLER_58_650 ();
 sg13g2_decap_8 FILLER_58_690 ();
 sg13g2_decap_4 FILLER_58_697 ();
 sg13g2_fill_2 FILLER_58_701 ();
 sg13g2_decap_4 FILLER_58_729 ();
 sg13g2_decap_8 FILLER_58_741 ();
 sg13g2_decap_8 FILLER_58_748 ();
 sg13g2_decap_8 FILLER_58_755 ();
 sg13g2_fill_2 FILLER_58_762 ();
 sg13g2_fill_1 FILLER_58_764 ();
 sg13g2_decap_8 FILLER_58_777 ();
 sg13g2_decap_4 FILLER_58_784 ();
 sg13g2_decap_8 FILLER_58_793 ();
 sg13g2_decap_8 FILLER_58_800 ();
 sg13g2_decap_4 FILLER_58_807 ();
 sg13g2_fill_2 FILLER_58_811 ();
 sg13g2_decap_8 FILLER_58_833 ();
 sg13g2_decap_4 FILLER_58_840 ();
 sg13g2_fill_2 FILLER_58_844 ();
 sg13g2_decap_4 FILLER_58_856 ();
 sg13g2_fill_1 FILLER_58_868 ();
 sg13g2_decap_8 FILLER_58_874 ();
 sg13g2_fill_1 FILLER_58_881 ();
 sg13g2_decap_4 FILLER_58_890 ();
 sg13g2_decap_8 FILLER_58_898 ();
 sg13g2_decap_8 FILLER_58_905 ();
 sg13g2_decap_8 FILLER_58_912 ();
 sg13g2_decap_8 FILLER_58_919 ();
 sg13g2_decap_8 FILLER_58_926 ();
 sg13g2_decap_8 FILLER_58_933 ();
 sg13g2_fill_2 FILLER_58_940 ();
 sg13g2_fill_1 FILLER_58_942 ();
 sg13g2_fill_2 FILLER_58_953 ();
 sg13g2_fill_1 FILLER_58_955 ();
 sg13g2_fill_1 FILLER_58_960 ();
 sg13g2_decap_4 FILLER_58_976 ();
 sg13g2_fill_1 FILLER_58_980 ();
 sg13g2_fill_2 FILLER_58_1009 ();
 sg13g2_decap_4 FILLER_58_1017 ();
 sg13g2_fill_2 FILLER_58_1021 ();
 sg13g2_decap_8 FILLER_58_1028 ();
 sg13g2_decap_8 FILLER_58_1035 ();
 sg13g2_decap_8 FILLER_58_1042 ();
 sg13g2_decap_8 FILLER_58_1049 ();
 sg13g2_fill_1 FILLER_58_1056 ();
 sg13g2_fill_1 FILLER_58_1066 ();
 sg13g2_decap_8 FILLER_58_1085 ();
 sg13g2_decap_8 FILLER_58_1092 ();
 sg13g2_fill_2 FILLER_58_1099 ();
 sg13g2_fill_1 FILLER_58_1101 ();
 sg13g2_decap_8 FILLER_58_1111 ();
 sg13g2_fill_1 FILLER_58_1118 ();
 sg13g2_decap_8 FILLER_58_1130 ();
 sg13g2_decap_8 FILLER_58_1145 ();
 sg13g2_decap_4 FILLER_58_1152 ();
 sg13g2_fill_2 FILLER_58_1156 ();
 sg13g2_fill_1 FILLER_58_1177 ();
 sg13g2_decap_8 FILLER_58_1193 ();
 sg13g2_decap_8 FILLER_58_1200 ();
 sg13g2_decap_8 FILLER_58_1207 ();
 sg13g2_decap_4 FILLER_58_1214 ();
 sg13g2_fill_2 FILLER_58_1228 ();
 sg13g2_fill_1 FILLER_58_1230 ();
 sg13g2_decap_4 FILLER_58_1236 ();
 sg13g2_fill_1 FILLER_58_1240 ();
 sg13g2_decap_4 FILLER_58_1254 ();
 sg13g2_decap_4 FILLER_58_1264 ();
 sg13g2_fill_2 FILLER_58_1268 ();
 sg13g2_decap_8 FILLER_58_1280 ();
 sg13g2_decap_8 FILLER_58_1287 ();
 sg13g2_decap_8 FILLER_58_1294 ();
 sg13g2_decap_8 FILLER_58_1301 ();
 sg13g2_decap_8 FILLER_58_1308 ();
 sg13g2_decap_8 FILLER_58_1315 ();
 sg13g2_decap_4 FILLER_58_1322 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_fill_2 FILLER_59_65 ();
 sg13g2_decap_8 FILLER_59_72 ();
 sg13g2_decap_4 FILLER_59_79 ();
 sg13g2_decap_4 FILLER_59_88 ();
 sg13g2_fill_1 FILLER_59_92 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_fill_2 FILLER_59_127 ();
 sg13g2_fill_1 FILLER_59_129 ();
 sg13g2_decap_8 FILLER_59_180 ();
 sg13g2_fill_2 FILLER_59_187 ();
 sg13g2_decap_4 FILLER_59_210 ();
 sg13g2_fill_1 FILLER_59_214 ();
 sg13g2_decap_8 FILLER_59_219 ();
 sg13g2_decap_4 FILLER_59_226 ();
 sg13g2_fill_1 FILLER_59_239 ();
 sg13g2_decap_8 FILLER_59_245 ();
 sg13g2_fill_2 FILLER_59_252 ();
 sg13g2_decap_8 FILLER_59_267 ();
 sg13g2_decap_8 FILLER_59_274 ();
 sg13g2_decap_8 FILLER_59_281 ();
 sg13g2_decap_8 FILLER_59_288 ();
 sg13g2_decap_4 FILLER_59_295 ();
 sg13g2_fill_1 FILLER_59_299 ();
 sg13g2_decap_4 FILLER_59_304 ();
 sg13g2_decap_8 FILLER_59_311 ();
 sg13g2_decap_8 FILLER_59_318 ();
 sg13g2_decap_8 FILLER_59_325 ();
 sg13g2_fill_2 FILLER_59_332 ();
 sg13g2_fill_1 FILLER_59_334 ();
 sg13g2_decap_8 FILLER_59_339 ();
 sg13g2_fill_1 FILLER_59_346 ();
 sg13g2_decap_8 FILLER_59_356 ();
 sg13g2_decap_8 FILLER_59_363 ();
 sg13g2_decap_8 FILLER_59_370 ();
 sg13g2_fill_1 FILLER_59_381 ();
 sg13g2_decap_4 FILLER_59_386 ();
 sg13g2_fill_1 FILLER_59_401 ();
 sg13g2_decap_4 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_410 ();
 sg13g2_decap_8 FILLER_59_416 ();
 sg13g2_decap_8 FILLER_59_423 ();
 sg13g2_decap_8 FILLER_59_430 ();
 sg13g2_decap_8 FILLER_59_437 ();
 sg13g2_decap_4 FILLER_59_444 ();
 sg13g2_decap_8 FILLER_59_452 ();
 sg13g2_fill_2 FILLER_59_459 ();
 sg13g2_decap_8 FILLER_59_466 ();
 sg13g2_decap_8 FILLER_59_473 ();
 sg13g2_decap_4 FILLER_59_480 ();
 sg13g2_decap_8 FILLER_59_487 ();
 sg13g2_fill_1 FILLER_59_494 ();
 sg13g2_decap_8 FILLER_59_499 ();
 sg13g2_fill_2 FILLER_59_506 ();
 sg13g2_decap_4 FILLER_59_511 ();
 sg13g2_decap_4 FILLER_59_549 ();
 sg13g2_decap_8 FILLER_59_579 ();
 sg13g2_decap_8 FILLER_59_586 ();
 sg13g2_decap_8 FILLER_59_597 ();
 sg13g2_fill_2 FILLER_59_604 ();
 sg13g2_decap_8 FILLER_59_628 ();
 sg13g2_decap_4 FILLER_59_653 ();
 sg13g2_fill_2 FILLER_59_657 ();
 sg13g2_decap_4 FILLER_59_663 ();
 sg13g2_decap_8 FILLER_59_676 ();
 sg13g2_decap_8 FILLER_59_683 ();
 sg13g2_decap_8 FILLER_59_690 ();
 sg13g2_fill_1 FILLER_59_697 ();
 sg13g2_fill_2 FILLER_59_716 ();
 sg13g2_fill_1 FILLER_59_718 ();
 sg13g2_decap_8 FILLER_59_722 ();
 sg13g2_decap_8 FILLER_59_729 ();
 sg13g2_fill_1 FILLER_59_736 ();
 sg13g2_fill_2 FILLER_59_770 ();
 sg13g2_decap_8 FILLER_59_776 ();
 sg13g2_decap_8 FILLER_59_783 ();
 sg13g2_decap_8 FILLER_59_790 ();
 sg13g2_decap_8 FILLER_59_797 ();
 sg13g2_decap_8 FILLER_59_804 ();
 sg13g2_decap_8 FILLER_59_811 ();
 sg13g2_decap_8 FILLER_59_818 ();
 sg13g2_decap_4 FILLER_59_825 ();
 sg13g2_fill_2 FILLER_59_829 ();
 sg13g2_decap_8 FILLER_59_836 ();
 sg13g2_fill_2 FILLER_59_843 ();
 sg13g2_decap_8 FILLER_59_856 ();
 sg13g2_decap_8 FILLER_59_863 ();
 sg13g2_fill_2 FILLER_59_870 ();
 sg13g2_fill_1 FILLER_59_872 ();
 sg13g2_decap_8 FILLER_59_879 ();
 sg13g2_fill_2 FILLER_59_886 ();
 sg13g2_fill_1 FILLER_59_888 ();
 sg13g2_decap_4 FILLER_59_915 ();
 sg13g2_fill_2 FILLER_59_919 ();
 sg13g2_fill_1 FILLER_59_927 ();
 sg13g2_fill_2 FILLER_59_937 ();
 sg13g2_fill_1 FILLER_59_939 ();
 sg13g2_fill_2 FILLER_59_949 ();
 sg13g2_fill_1 FILLER_59_951 ();
 sg13g2_decap_8 FILLER_59_964 ();
 sg13g2_decap_8 FILLER_59_976 ();
 sg13g2_decap_4 FILLER_59_983 ();
 sg13g2_fill_2 FILLER_59_987 ();
 sg13g2_fill_1 FILLER_59_999 ();
 sg13g2_decap_8 FILLER_59_1005 ();
 sg13g2_decap_8 FILLER_59_1012 ();
 sg13g2_fill_1 FILLER_59_1019 ();
 sg13g2_fill_1 FILLER_59_1026 ();
 sg13g2_decap_8 FILLER_59_1032 ();
 sg13g2_decap_4 FILLER_59_1055 ();
 sg13g2_fill_1 FILLER_59_1059 ();
 sg13g2_fill_1 FILLER_59_1072 ();
 sg13g2_decap_8 FILLER_59_1093 ();
 sg13g2_decap_4 FILLER_59_1100 ();
 sg13g2_decap_4 FILLER_59_1109 ();
 sg13g2_fill_1 FILLER_59_1113 ();
 sg13g2_decap_8 FILLER_59_1118 ();
 sg13g2_decap_8 FILLER_59_1125 ();
 sg13g2_decap_8 FILLER_59_1132 ();
 sg13g2_decap_8 FILLER_59_1139 ();
 sg13g2_decap_8 FILLER_59_1146 ();
 sg13g2_fill_2 FILLER_59_1153 ();
 sg13g2_decap_4 FILLER_59_1159 ();
 sg13g2_fill_1 FILLER_59_1163 ();
 sg13g2_decap_8 FILLER_59_1173 ();
 sg13g2_decap_8 FILLER_59_1180 ();
 sg13g2_fill_2 FILLER_59_1187 ();
 sg13g2_fill_1 FILLER_59_1189 ();
 sg13g2_fill_2 FILLER_59_1206 ();
 sg13g2_fill_1 FILLER_59_1208 ();
 sg13g2_decap_8 FILLER_59_1214 ();
 sg13g2_fill_1 FILLER_59_1234 ();
 sg13g2_decap_4 FILLER_59_1241 ();
 sg13g2_fill_2 FILLER_59_1245 ();
 sg13g2_decap_4 FILLER_59_1252 ();
 sg13g2_fill_2 FILLER_59_1271 ();
 sg13g2_decap_8 FILLER_59_1282 ();
 sg13g2_decap_8 FILLER_59_1289 ();
 sg13g2_decap_8 FILLER_59_1296 ();
 sg13g2_decap_8 FILLER_59_1303 ();
 sg13g2_decap_8 FILLER_59_1310 ();
 sg13g2_decap_8 FILLER_59_1317 ();
 sg13g2_fill_2 FILLER_59_1324 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_4 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_48 ();
 sg13g2_decap_8 FILLER_60_55 ();
 sg13g2_fill_2 FILLER_60_62 ();
 sg13g2_fill_1 FILLER_60_64 ();
 sg13g2_decap_8 FILLER_60_78 ();
 sg13g2_decap_8 FILLER_60_85 ();
 sg13g2_decap_8 FILLER_60_92 ();
 sg13g2_decap_8 FILLER_60_99 ();
 sg13g2_fill_2 FILLER_60_112 ();
 sg13g2_fill_1 FILLER_60_114 ();
 sg13g2_fill_2 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_decap_8 FILLER_60_133 ();
 sg13g2_fill_1 FILLER_60_140 ();
 sg13g2_decap_8 FILLER_60_146 ();
 sg13g2_decap_8 FILLER_60_153 ();
 sg13g2_decap_8 FILLER_60_160 ();
 sg13g2_decap_8 FILLER_60_167 ();
 sg13g2_decap_4 FILLER_60_174 ();
 sg13g2_fill_2 FILLER_60_178 ();
 sg13g2_decap_4 FILLER_60_184 ();
 sg13g2_decap_8 FILLER_60_193 ();
 sg13g2_decap_8 FILLER_60_200 ();
 sg13g2_fill_2 FILLER_60_207 ();
 sg13g2_fill_1 FILLER_60_218 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_decap_4 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_239 ();
 sg13g2_decap_8 FILLER_60_246 ();
 sg13g2_decap_8 FILLER_60_253 ();
 sg13g2_decap_8 FILLER_60_260 ();
 sg13g2_decap_8 FILLER_60_267 ();
 sg13g2_decap_8 FILLER_60_274 ();
 sg13g2_decap_8 FILLER_60_281 ();
 sg13g2_decap_8 FILLER_60_288 ();
 sg13g2_decap_8 FILLER_60_295 ();
 sg13g2_decap_8 FILLER_60_311 ();
 sg13g2_decap_8 FILLER_60_322 ();
 sg13g2_decap_4 FILLER_60_329 ();
 sg13g2_fill_2 FILLER_60_337 ();
 sg13g2_fill_1 FILLER_60_339 ();
 sg13g2_decap_8 FILLER_60_345 ();
 sg13g2_decap_8 FILLER_60_352 ();
 sg13g2_decap_8 FILLER_60_359 ();
 sg13g2_decap_8 FILLER_60_366 ();
 sg13g2_decap_8 FILLER_60_373 ();
 sg13g2_fill_2 FILLER_60_380 ();
 sg13g2_fill_1 FILLER_60_382 ();
 sg13g2_decap_8 FILLER_60_388 ();
 sg13g2_decap_8 FILLER_60_395 ();
 sg13g2_decap_8 FILLER_60_402 ();
 sg13g2_decap_8 FILLER_60_409 ();
 sg13g2_decap_8 FILLER_60_416 ();
 sg13g2_decap_8 FILLER_60_423 ();
 sg13g2_decap_8 FILLER_60_430 ();
 sg13g2_decap_8 FILLER_60_437 ();
 sg13g2_decap_8 FILLER_60_444 ();
 sg13g2_decap_8 FILLER_60_451 ();
 sg13g2_decap_8 FILLER_60_458 ();
 sg13g2_decap_4 FILLER_60_465 ();
 sg13g2_fill_1 FILLER_60_469 ();
 sg13g2_decap_8 FILLER_60_475 ();
 sg13g2_decap_8 FILLER_60_482 ();
 sg13g2_decap_8 FILLER_60_489 ();
 sg13g2_decap_8 FILLER_60_496 ();
 sg13g2_decap_8 FILLER_60_503 ();
 sg13g2_decap_8 FILLER_60_510 ();
 sg13g2_decap_8 FILLER_60_517 ();
 sg13g2_fill_2 FILLER_60_524 ();
 sg13g2_fill_1 FILLER_60_526 ();
 sg13g2_decap_8 FILLER_60_531 ();
 sg13g2_decap_8 FILLER_60_538 ();
 sg13g2_decap_8 FILLER_60_545 ();
 sg13g2_decap_8 FILLER_60_552 ();
 sg13g2_fill_2 FILLER_60_559 ();
 sg13g2_fill_2 FILLER_60_565 ();
 sg13g2_fill_1 FILLER_60_567 ();
 sg13g2_decap_8 FILLER_60_572 ();
 sg13g2_decap_8 FILLER_60_579 ();
 sg13g2_decap_8 FILLER_60_586 ();
 sg13g2_decap_8 FILLER_60_593 ();
 sg13g2_decap_8 FILLER_60_600 ();
 sg13g2_fill_2 FILLER_60_607 ();
 sg13g2_fill_1 FILLER_60_609 ();
 sg13g2_decap_4 FILLER_60_614 ();
 sg13g2_decap_8 FILLER_60_654 ();
 sg13g2_decap_8 FILLER_60_661 ();
 sg13g2_decap_8 FILLER_60_668 ();
 sg13g2_decap_8 FILLER_60_675 ();
 sg13g2_decap_8 FILLER_60_682 ();
 sg13g2_decap_8 FILLER_60_689 ();
 sg13g2_decap_8 FILLER_60_696 ();
 sg13g2_decap_8 FILLER_60_703 ();
 sg13g2_decap_8 FILLER_60_710 ();
 sg13g2_decap_8 FILLER_60_717 ();
 sg13g2_decap_8 FILLER_60_724 ();
 sg13g2_decap_8 FILLER_60_731 ();
 sg13g2_decap_4 FILLER_60_738 ();
 sg13g2_fill_1 FILLER_60_742 ();
 sg13g2_decap_8 FILLER_60_747 ();
 sg13g2_decap_8 FILLER_60_754 ();
 sg13g2_fill_1 FILLER_60_761 ();
 sg13g2_decap_8 FILLER_60_767 ();
 sg13g2_decap_4 FILLER_60_774 ();
 sg13g2_decap_4 FILLER_60_784 ();
 sg13g2_decap_8 FILLER_60_794 ();
 sg13g2_decap_8 FILLER_60_801 ();
 sg13g2_decap_8 FILLER_60_808 ();
 sg13g2_decap_8 FILLER_60_815 ();
 sg13g2_decap_8 FILLER_60_822 ();
 sg13g2_decap_8 FILLER_60_829 ();
 sg13g2_decap_8 FILLER_60_841 ();
 sg13g2_fill_2 FILLER_60_848 ();
 sg13g2_decap_8 FILLER_60_856 ();
 sg13g2_decap_8 FILLER_60_863 ();
 sg13g2_decap_8 FILLER_60_870 ();
 sg13g2_decap_8 FILLER_60_877 ();
 sg13g2_decap_8 FILLER_60_884 ();
 sg13g2_decap_8 FILLER_60_891 ();
 sg13g2_decap_8 FILLER_60_898 ();
 sg13g2_fill_2 FILLER_60_905 ();
 sg13g2_decap_4 FILLER_60_912 ();
 sg13g2_decap_8 FILLER_60_921 ();
 sg13g2_decap_8 FILLER_60_928 ();
 sg13g2_decap_8 FILLER_60_935 ();
 sg13g2_decap_8 FILLER_60_942 ();
 sg13g2_fill_1 FILLER_60_949 ();
 sg13g2_decap_4 FILLER_60_954 ();
 sg13g2_fill_1 FILLER_60_972 ();
 sg13g2_decap_8 FILLER_60_977 ();
 sg13g2_decap_8 FILLER_60_984 ();
 sg13g2_fill_2 FILLER_60_991 ();
 sg13g2_fill_2 FILLER_60_996 ();
 sg13g2_fill_1 FILLER_60_998 ();
 sg13g2_decap_8 FILLER_60_1003 ();
 sg13g2_decap_8 FILLER_60_1010 ();
 sg13g2_decap_8 FILLER_60_1017 ();
 sg13g2_decap_8 FILLER_60_1024 ();
 sg13g2_decap_8 FILLER_60_1031 ();
 sg13g2_fill_2 FILLER_60_1038 ();
 sg13g2_decap_4 FILLER_60_1045 ();
 sg13g2_decap_8 FILLER_60_1059 ();
 sg13g2_decap_8 FILLER_60_1066 ();
 sg13g2_decap_4 FILLER_60_1073 ();
 sg13g2_fill_2 FILLER_60_1077 ();
 sg13g2_decap_8 FILLER_60_1084 ();
 sg13g2_decap_8 FILLER_60_1091 ();
 sg13g2_decap_4 FILLER_60_1098 ();
 sg13g2_decap_8 FILLER_60_1117 ();
 sg13g2_decap_4 FILLER_60_1124 ();
 sg13g2_fill_1 FILLER_60_1128 ();
 sg13g2_decap_8 FILLER_60_1134 ();
 sg13g2_decap_8 FILLER_60_1141 ();
 sg13g2_decap_4 FILLER_60_1148 ();
 sg13g2_fill_2 FILLER_60_1152 ();
 sg13g2_decap_8 FILLER_60_1159 ();
 sg13g2_decap_8 FILLER_60_1166 ();
 sg13g2_decap_8 FILLER_60_1173 ();
 sg13g2_decap_8 FILLER_60_1180 ();
 sg13g2_decap_8 FILLER_60_1187 ();
 sg13g2_decap_8 FILLER_60_1194 ();
 sg13g2_fill_2 FILLER_60_1201 ();
 sg13g2_fill_1 FILLER_60_1203 ();
 sg13g2_fill_2 FILLER_60_1209 ();
 sg13g2_fill_2 FILLER_60_1221 ();
 sg13g2_decap_8 FILLER_60_1228 ();
 sg13g2_decap_8 FILLER_60_1235 ();
 sg13g2_decap_8 FILLER_60_1242 ();
 sg13g2_decap_8 FILLER_60_1249 ();
 sg13g2_decap_8 FILLER_60_1256 ();
 sg13g2_decap_8 FILLER_60_1263 ();
 sg13g2_fill_2 FILLER_60_1270 ();
 sg13g2_fill_2 FILLER_60_1277 ();
 sg13g2_decap_8 FILLER_60_1283 ();
 sg13g2_decap_8 FILLER_60_1290 ();
 sg13g2_decap_8 FILLER_60_1297 ();
 sg13g2_decap_8 FILLER_60_1304 ();
 sg13g2_decap_8 FILLER_60_1311 ();
 sg13g2_decap_8 FILLER_60_1318 ();
 sg13g2_fill_1 FILLER_60_1325 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_fill_2 FILLER_61_35 ();
 sg13g2_fill_1 FILLER_61_37 ();
 sg13g2_decap_8 FILLER_61_43 ();
 sg13g2_decap_8 FILLER_61_50 ();
 sg13g2_decap_8 FILLER_61_57 ();
 sg13g2_decap_8 FILLER_61_64 ();
 sg13g2_fill_2 FILLER_61_79 ();
 sg13g2_decap_8 FILLER_61_92 ();
 sg13g2_fill_2 FILLER_61_99 ();
 sg13g2_fill_1 FILLER_61_101 ();
 sg13g2_decap_4 FILLER_61_105 ();
 sg13g2_fill_1 FILLER_61_109 ();
 sg13g2_fill_2 FILLER_61_118 ();
 sg13g2_fill_1 FILLER_61_125 ();
 sg13g2_fill_2 FILLER_61_130 ();
 sg13g2_fill_2 FILLER_61_136 ();
 sg13g2_fill_2 FILLER_61_142 ();
 sg13g2_decap_8 FILLER_61_149 ();
 sg13g2_decap_8 FILLER_61_156 ();
 sg13g2_decap_8 FILLER_61_163 ();
 sg13g2_decap_8 FILLER_61_170 ();
 sg13g2_decap_8 FILLER_61_177 ();
 sg13g2_decap_8 FILLER_61_184 ();
 sg13g2_decap_8 FILLER_61_191 ();
 sg13g2_fill_1 FILLER_61_198 ();
 sg13g2_decap_4 FILLER_61_204 ();
 sg13g2_fill_1 FILLER_61_218 ();
 sg13g2_decap_8 FILLER_61_224 ();
 sg13g2_decap_8 FILLER_61_231 ();
 sg13g2_decap_8 FILLER_61_238 ();
 sg13g2_decap_8 FILLER_61_245 ();
 sg13g2_fill_2 FILLER_61_252 ();
 sg13g2_fill_1 FILLER_61_254 ();
 sg13g2_decap_8 FILLER_61_260 ();
 sg13g2_fill_1 FILLER_61_267 ();
 sg13g2_fill_2 FILLER_61_281 ();
 sg13g2_decap_8 FILLER_61_296 ();
 sg13g2_decap_8 FILLER_61_303 ();
 sg13g2_decap_8 FILLER_61_310 ();
 sg13g2_decap_8 FILLER_61_317 ();
 sg13g2_decap_8 FILLER_61_324 ();
 sg13g2_decap_4 FILLER_61_331 ();
 sg13g2_fill_1 FILLER_61_335 ();
 sg13g2_decap_8 FILLER_61_341 ();
 sg13g2_decap_8 FILLER_61_348 ();
 sg13g2_decap_8 FILLER_61_355 ();
 sg13g2_decap_8 FILLER_61_362 ();
 sg13g2_decap_8 FILLER_61_369 ();
 sg13g2_decap_4 FILLER_61_376 ();
 sg13g2_fill_1 FILLER_61_380 ();
 sg13g2_decap_8 FILLER_61_385 ();
 sg13g2_decap_8 FILLER_61_392 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_decap_8 FILLER_61_406 ();
 sg13g2_decap_4 FILLER_61_413 ();
 sg13g2_fill_1 FILLER_61_417 ();
 sg13g2_decap_4 FILLER_61_422 ();
 sg13g2_decap_8 FILLER_61_430 ();
 sg13g2_decap_8 FILLER_61_437 ();
 sg13g2_decap_8 FILLER_61_444 ();
 sg13g2_decap_4 FILLER_61_451 ();
 sg13g2_decap_8 FILLER_61_486 ();
 sg13g2_decap_8 FILLER_61_493 ();
 sg13g2_fill_2 FILLER_61_500 ();
 sg13g2_decap_8 FILLER_61_510 ();
 sg13g2_decap_8 FILLER_61_517 ();
 sg13g2_decap_8 FILLER_61_524 ();
 sg13g2_decap_8 FILLER_61_531 ();
 sg13g2_decap_4 FILLER_61_538 ();
 sg13g2_decap_8 FILLER_61_547 ();
 sg13g2_decap_8 FILLER_61_554 ();
 sg13g2_fill_2 FILLER_61_561 ();
 sg13g2_fill_1 FILLER_61_563 ();
 sg13g2_decap_8 FILLER_61_580 ();
 sg13g2_decap_8 FILLER_61_587 ();
 sg13g2_decap_8 FILLER_61_594 ();
 sg13g2_decap_8 FILLER_61_601 ();
 sg13g2_decap_8 FILLER_61_608 ();
 sg13g2_decap_8 FILLER_61_615 ();
 sg13g2_fill_2 FILLER_61_622 ();
 sg13g2_decap_4 FILLER_61_628 ();
 sg13g2_decap_4 FILLER_61_636 ();
 sg13g2_fill_2 FILLER_61_640 ();
 sg13g2_fill_1 FILLER_61_645 ();
 sg13g2_decap_8 FILLER_61_651 ();
 sg13g2_fill_1 FILLER_61_658 ();
 sg13g2_decap_4 FILLER_61_664 ();
 sg13g2_fill_1 FILLER_61_668 ();
 sg13g2_decap_8 FILLER_61_673 ();
 sg13g2_decap_8 FILLER_61_680 ();
 sg13g2_decap_8 FILLER_61_687 ();
 sg13g2_decap_4 FILLER_61_694 ();
 sg13g2_fill_1 FILLER_61_698 ();
 sg13g2_fill_1 FILLER_61_713 ();
 sg13g2_decap_8 FILLER_61_718 ();
 sg13g2_decap_8 FILLER_61_725 ();
 sg13g2_decap_8 FILLER_61_732 ();
 sg13g2_decap_8 FILLER_61_739 ();
 sg13g2_decap_8 FILLER_61_746 ();
 sg13g2_decap_8 FILLER_61_753 ();
 sg13g2_decap_8 FILLER_61_760 ();
 sg13g2_fill_1 FILLER_61_767 ();
 sg13g2_decap_8 FILLER_61_790 ();
 sg13g2_decap_8 FILLER_61_797 ();
 sg13g2_decap_8 FILLER_61_804 ();
 sg13g2_decap_8 FILLER_61_811 ();
 sg13g2_decap_8 FILLER_61_818 ();
 sg13g2_decap_8 FILLER_61_825 ();
 sg13g2_decap_8 FILLER_61_832 ();
 sg13g2_fill_2 FILLER_61_839 ();
 sg13g2_decap_8 FILLER_61_845 ();
 sg13g2_decap_8 FILLER_61_852 ();
 sg13g2_decap_4 FILLER_61_859 ();
 sg13g2_fill_2 FILLER_61_863 ();
 sg13g2_fill_2 FILLER_61_871 ();
 sg13g2_fill_1 FILLER_61_873 ();
 sg13g2_decap_8 FILLER_61_878 ();
 sg13g2_decap_4 FILLER_61_885 ();
 sg13g2_fill_2 FILLER_61_889 ();
 sg13g2_decap_8 FILLER_61_896 ();
 sg13g2_decap_4 FILLER_61_903 ();
 sg13g2_fill_1 FILLER_61_907 ();
 sg13g2_decap_8 FILLER_61_913 ();
 sg13g2_decap_8 FILLER_61_920 ();
 sg13g2_fill_1 FILLER_61_930 ();
 sg13g2_decap_8 FILLER_61_936 ();
 sg13g2_fill_1 FILLER_61_943 ();
 sg13g2_fill_1 FILLER_61_950 ();
 sg13g2_decap_8 FILLER_61_960 ();
 sg13g2_decap_8 FILLER_61_967 ();
 sg13g2_decap_4 FILLER_61_974 ();
 sg13g2_fill_2 FILLER_61_983 ();
 sg13g2_fill_1 FILLER_61_985 ();
 sg13g2_decap_8 FILLER_61_990 ();
 sg13g2_fill_1 FILLER_61_997 ();
 sg13g2_decap_4 FILLER_61_1009 ();
 sg13g2_fill_2 FILLER_61_1013 ();
 sg13g2_decap_8 FILLER_61_1022 ();
 sg13g2_decap_8 FILLER_61_1029 ();
 sg13g2_decap_4 FILLER_61_1036 ();
 sg13g2_decap_8 FILLER_61_1044 ();
 sg13g2_fill_1 FILLER_61_1051 ();
 sg13g2_decap_8 FILLER_61_1057 ();
 sg13g2_decap_8 FILLER_61_1067 ();
 sg13g2_fill_2 FILLER_61_1074 ();
 sg13g2_decap_4 FILLER_61_1080 ();
 sg13g2_decap_8 FILLER_61_1092 ();
 sg13g2_decap_8 FILLER_61_1099 ();
 sg13g2_decap_8 FILLER_61_1106 ();
 sg13g2_decap_8 FILLER_61_1113 ();
 sg13g2_decap_4 FILLER_61_1120 ();
 sg13g2_fill_1 FILLER_61_1129 ();
 sg13g2_decap_4 FILLER_61_1138 ();
 sg13g2_fill_2 FILLER_61_1142 ();
 sg13g2_decap_4 FILLER_61_1154 ();
 sg13g2_fill_2 FILLER_61_1163 ();
 sg13g2_fill_2 FILLER_61_1170 ();
 sg13g2_decap_8 FILLER_61_1188 ();
 sg13g2_decap_4 FILLER_61_1195 ();
 sg13g2_fill_2 FILLER_61_1199 ();
 sg13g2_fill_2 FILLER_61_1217 ();
 sg13g2_fill_1 FILLER_61_1219 ();
 sg13g2_decap_8 FILLER_61_1225 ();
 sg13g2_fill_2 FILLER_61_1232 ();
 sg13g2_fill_2 FILLER_61_1239 ();
 sg13g2_fill_1 FILLER_61_1241 ();
 sg13g2_fill_1 FILLER_61_1247 ();
 sg13g2_fill_2 FILLER_61_1254 ();
 sg13g2_fill_1 FILLER_61_1260 ();
 sg13g2_decap_8 FILLER_61_1280 ();
 sg13g2_decap_8 FILLER_61_1287 ();
 sg13g2_decap_8 FILLER_61_1294 ();
 sg13g2_decap_8 FILLER_61_1301 ();
 sg13g2_decap_8 FILLER_61_1308 ();
 sg13g2_decap_8 FILLER_61_1315 ();
 sg13g2_decap_4 FILLER_61_1322 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_12 ();
 sg13g2_decap_8 FILLER_62_19 ();
 sg13g2_decap_8 FILLER_62_26 ();
 sg13g2_fill_1 FILLER_62_33 ();
 sg13g2_decap_8 FILLER_62_39 ();
 sg13g2_fill_1 FILLER_62_46 ();
 sg13g2_decap_8 FILLER_62_52 ();
 sg13g2_decap_4 FILLER_62_59 ();
 sg13g2_fill_2 FILLER_62_63 ();
 sg13g2_fill_1 FILLER_62_70 ();
 sg13g2_fill_2 FILLER_62_81 ();
 sg13g2_fill_1 FILLER_62_87 ();
 sg13g2_decap_8 FILLER_62_93 ();
 sg13g2_fill_1 FILLER_62_100 ();
 sg13g2_fill_1 FILLER_62_106 ();
 sg13g2_decap_8 FILLER_62_150 ();
 sg13g2_decap_4 FILLER_62_157 ();
 sg13g2_decap_4 FILLER_62_167 ();
 sg13g2_fill_1 FILLER_62_171 ();
 sg13g2_decap_8 FILLER_62_184 ();
 sg13g2_decap_8 FILLER_62_191 ();
 sg13g2_decap_4 FILLER_62_198 ();
 sg13g2_fill_1 FILLER_62_202 ();
 sg13g2_decap_4 FILLER_62_208 ();
 sg13g2_fill_2 FILLER_62_212 ();
 sg13g2_fill_1 FILLER_62_224 ();
 sg13g2_fill_2 FILLER_62_234 ();
 sg13g2_fill_1 FILLER_62_236 ();
 sg13g2_decap_4 FILLER_62_262 ();
 sg13g2_fill_2 FILLER_62_272 ();
 sg13g2_fill_1 FILLER_62_274 ();
 sg13g2_decap_8 FILLER_62_280 ();
 sg13g2_fill_2 FILLER_62_287 ();
 sg13g2_fill_1 FILLER_62_307 ();
 sg13g2_decap_4 FILLER_62_313 ();
 sg13g2_fill_1 FILLER_62_317 ();
 sg13g2_decap_4 FILLER_62_348 ();
 sg13g2_decap_8 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_364 ();
 sg13g2_decap_8 FILLER_62_371 ();
 sg13g2_decap_8 FILLER_62_378 ();
 sg13g2_decap_8 FILLER_62_385 ();
 sg13g2_decap_8 FILLER_62_392 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_decap_8 FILLER_62_406 ();
 sg13g2_decap_4 FILLER_62_413 ();
 sg13g2_fill_1 FILLER_62_417 ();
 sg13g2_decap_8 FILLER_62_427 ();
 sg13g2_decap_8 FILLER_62_434 ();
 sg13g2_decap_8 FILLER_62_441 ();
 sg13g2_decap_8 FILLER_62_448 ();
 sg13g2_decap_8 FILLER_62_455 ();
 sg13g2_decap_4 FILLER_62_462 ();
 sg13g2_decap_8 FILLER_62_470 ();
 sg13g2_decap_4 FILLER_62_477 ();
 sg13g2_fill_1 FILLER_62_481 ();
 sg13g2_decap_8 FILLER_62_487 ();
 sg13g2_decap_8 FILLER_62_494 ();
 sg13g2_fill_1 FILLER_62_501 ();
 sg13g2_decap_8 FILLER_62_510 ();
 sg13g2_decap_8 FILLER_62_517 ();
 sg13g2_decap_4 FILLER_62_524 ();
 sg13g2_fill_2 FILLER_62_528 ();
 sg13g2_decap_8 FILLER_62_566 ();
 sg13g2_decap_8 FILLER_62_573 ();
 sg13g2_decap_8 FILLER_62_606 ();
 sg13g2_decap_8 FILLER_62_613 ();
 sg13g2_decap_8 FILLER_62_620 ();
 sg13g2_decap_8 FILLER_62_627 ();
 sg13g2_decap_8 FILLER_62_634 ();
 sg13g2_decap_8 FILLER_62_641 ();
 sg13g2_decap_8 FILLER_62_648 ();
 sg13g2_decap_8 FILLER_62_655 ();
 sg13g2_decap_8 FILLER_62_662 ();
 sg13g2_fill_2 FILLER_62_669 ();
 sg13g2_fill_1 FILLER_62_671 ();
 sg13g2_decap_4 FILLER_62_677 ();
 sg13g2_fill_1 FILLER_62_681 ();
 sg13g2_decap_8 FILLER_62_686 ();
 sg13g2_decap_4 FILLER_62_693 ();
 sg13g2_fill_1 FILLER_62_697 ();
 sg13g2_decap_4 FILLER_62_701 ();
 sg13g2_fill_2 FILLER_62_705 ();
 sg13g2_decap_8 FILLER_62_733 ();
 sg13g2_decap_8 FILLER_62_740 ();
 sg13g2_decap_8 FILLER_62_747 ();
 sg13g2_fill_2 FILLER_62_754 ();
 sg13g2_fill_2 FILLER_62_764 ();
 sg13g2_decap_8 FILLER_62_780 ();
 sg13g2_decap_8 FILLER_62_787 ();
 sg13g2_decap_8 FILLER_62_794 ();
 sg13g2_decap_4 FILLER_62_801 ();
 sg13g2_fill_2 FILLER_62_805 ();
 sg13g2_decap_4 FILLER_62_815 ();
 sg13g2_fill_1 FILLER_62_819 ();
 sg13g2_decap_8 FILLER_62_825 ();
 sg13g2_fill_1 FILLER_62_838 ();
 sg13g2_decap_4 FILLER_62_844 ();
 sg13g2_fill_2 FILLER_62_848 ();
 sg13g2_fill_2 FILLER_62_856 ();
 sg13g2_fill_1 FILLER_62_858 ();
 sg13g2_decap_8 FILLER_62_874 ();
 sg13g2_decap_8 FILLER_62_881 ();
 sg13g2_decap_8 FILLER_62_888 ();
 sg13g2_decap_4 FILLER_62_908 ();
 sg13g2_decap_8 FILLER_62_917 ();
 sg13g2_fill_2 FILLER_62_924 ();
 sg13g2_fill_1 FILLER_62_926 ();
 sg13g2_decap_8 FILLER_62_941 ();
 sg13g2_decap_4 FILLER_62_948 ();
 sg13g2_decap_8 FILLER_62_956 ();
 sg13g2_decap_4 FILLER_62_963 ();
 sg13g2_fill_1 FILLER_62_967 ();
 sg13g2_decap_8 FILLER_62_972 ();
 sg13g2_decap_8 FILLER_62_979 ();
 sg13g2_decap_4 FILLER_62_986 ();
 sg13g2_fill_2 FILLER_62_990 ();
 sg13g2_decap_8 FILLER_62_1005 ();
 sg13g2_decap_8 FILLER_62_1012 ();
 sg13g2_decap_8 FILLER_62_1019 ();
 sg13g2_decap_4 FILLER_62_1026 ();
 sg13g2_fill_1 FILLER_62_1030 ();
 sg13g2_decap_8 FILLER_62_1042 ();
 sg13g2_decap_8 FILLER_62_1049 ();
 sg13g2_decap_8 FILLER_62_1056 ();
 sg13g2_fill_2 FILLER_62_1063 ();
 sg13g2_decap_8 FILLER_62_1070 ();
 sg13g2_fill_2 FILLER_62_1077 ();
 sg13g2_fill_1 FILLER_62_1079 ();
 sg13g2_fill_1 FILLER_62_1089 ();
 sg13g2_decap_8 FILLER_62_1095 ();
 sg13g2_fill_1 FILLER_62_1102 ();
 sg13g2_decap_8 FILLER_62_1108 ();
 sg13g2_fill_1 FILLER_62_1115 ();
 sg13g2_fill_2 FILLER_62_1126 ();
 sg13g2_decap_8 FILLER_62_1134 ();
 sg13g2_decap_8 FILLER_62_1145 ();
 sg13g2_decap_8 FILLER_62_1152 ();
 sg13g2_fill_1 FILLER_62_1159 ();
 sg13g2_decap_8 FILLER_62_1166 ();
 sg13g2_decap_8 FILLER_62_1173 ();
 sg13g2_fill_1 FILLER_62_1180 ();
 sg13g2_decap_8 FILLER_62_1185 ();
 sg13g2_decap_8 FILLER_62_1192 ();
 sg13g2_fill_2 FILLER_62_1199 ();
 sg13g2_fill_1 FILLER_62_1201 ();
 sg13g2_fill_2 FILLER_62_1212 ();
 sg13g2_fill_1 FILLER_62_1214 ();
 sg13g2_decap_4 FILLER_62_1221 ();
 sg13g2_fill_2 FILLER_62_1225 ();
 sg13g2_decap_4 FILLER_62_1232 ();
 sg13g2_fill_2 FILLER_62_1250 ();
 sg13g2_fill_1 FILLER_62_1252 ();
 sg13g2_fill_2 FILLER_62_1273 ();
 sg13g2_fill_1 FILLER_62_1275 ();
 sg13g2_decap_8 FILLER_62_1281 ();
 sg13g2_decap_8 FILLER_62_1288 ();
 sg13g2_decap_8 FILLER_62_1295 ();
 sg13g2_decap_8 FILLER_62_1302 ();
 sg13g2_decap_8 FILLER_62_1309 ();
 sg13g2_decap_8 FILLER_62_1316 ();
 sg13g2_fill_2 FILLER_62_1323 ();
 sg13g2_fill_1 FILLER_62_1325 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_27 ();
 sg13g2_fill_2 FILLER_63_34 ();
 sg13g2_decap_8 FILLER_63_44 ();
 sg13g2_decap_8 FILLER_63_51 ();
 sg13g2_decap_8 FILLER_63_58 ();
 sg13g2_decap_4 FILLER_63_65 ();
 sg13g2_fill_1 FILLER_63_69 ();
 sg13g2_decap_4 FILLER_63_74 ();
 sg13g2_fill_2 FILLER_63_78 ();
 sg13g2_decap_8 FILLER_63_88 ();
 sg13g2_decap_8 FILLER_63_100 ();
 sg13g2_decap_8 FILLER_63_107 ();
 sg13g2_decap_4 FILLER_63_114 ();
 sg13g2_fill_2 FILLER_63_118 ();
 sg13g2_decap_8 FILLER_63_129 ();
 sg13g2_decap_8 FILLER_63_136 ();
 sg13g2_decap_8 FILLER_63_143 ();
 sg13g2_fill_2 FILLER_63_150 ();
 sg13g2_fill_1 FILLER_63_152 ();
 sg13g2_fill_1 FILLER_63_172 ();
 sg13g2_decap_8 FILLER_63_184 ();
 sg13g2_decap_8 FILLER_63_191 ();
 sg13g2_decap_8 FILLER_63_198 ();
 sg13g2_fill_2 FILLER_63_205 ();
 sg13g2_fill_1 FILLER_63_207 ();
 sg13g2_decap_8 FILLER_63_213 ();
 sg13g2_fill_2 FILLER_63_264 ();
 sg13g2_fill_2 FILLER_63_270 ();
 sg13g2_decap_8 FILLER_63_280 ();
 sg13g2_decap_8 FILLER_63_287 ();
 sg13g2_fill_1 FILLER_63_294 ();
 sg13g2_decap_8 FILLER_63_307 ();
 sg13g2_fill_2 FILLER_63_314 ();
 sg13g2_decap_4 FILLER_63_326 ();
 sg13g2_fill_1 FILLER_63_330 ();
 sg13g2_decap_8 FILLER_63_357 ();
 sg13g2_fill_2 FILLER_63_364 ();
 sg13g2_decap_8 FILLER_63_371 ();
 sg13g2_decap_8 FILLER_63_378 ();
 sg13g2_decap_8 FILLER_63_385 ();
 sg13g2_decap_4 FILLER_63_392 ();
 sg13g2_fill_2 FILLER_63_396 ();
 sg13g2_decap_4 FILLER_63_402 ();
 sg13g2_fill_1 FILLER_63_406 ();
 sg13g2_fill_2 FILLER_63_411 ();
 sg13g2_fill_1 FILLER_63_413 ();
 sg13g2_decap_8 FILLER_63_444 ();
 sg13g2_decap_8 FILLER_63_451 ();
 sg13g2_fill_2 FILLER_63_458 ();
 sg13g2_fill_1 FILLER_63_460 ();
 sg13g2_decap_4 FILLER_63_465 ();
 sg13g2_fill_2 FILLER_63_469 ();
 sg13g2_decap_8 FILLER_63_475 ();
 sg13g2_decap_8 FILLER_63_482 ();
 sg13g2_decap_8 FILLER_63_489 ();
 sg13g2_fill_2 FILLER_63_527 ();
 sg13g2_decap_8 FILLER_63_534 ();
 sg13g2_decap_8 FILLER_63_541 ();
 sg13g2_decap_8 FILLER_63_552 ();
 sg13g2_decap_8 FILLER_63_559 ();
 sg13g2_decap_8 FILLER_63_566 ();
 sg13g2_decap_8 FILLER_63_573 ();
 sg13g2_decap_8 FILLER_63_610 ();
 sg13g2_decap_8 FILLER_63_617 ();
 sg13g2_decap_8 FILLER_63_624 ();
 sg13g2_decap_4 FILLER_63_631 ();
 sg13g2_fill_1 FILLER_63_635 ();
 sg13g2_decap_8 FILLER_63_649 ();
 sg13g2_decap_8 FILLER_63_656 ();
 sg13g2_fill_2 FILLER_63_692 ();
 sg13g2_fill_1 FILLER_63_694 ();
 sg13g2_decap_4 FILLER_63_700 ();
 sg13g2_decap_8 FILLER_63_725 ();
 sg13g2_decap_8 FILLER_63_732 ();
 sg13g2_decap_8 FILLER_63_739 ();
 sg13g2_decap_8 FILLER_63_746 ();
 sg13g2_decap_4 FILLER_63_753 ();
 sg13g2_fill_1 FILLER_63_757 ();
 sg13g2_decap_8 FILLER_63_763 ();
 sg13g2_decap_4 FILLER_63_770 ();
 sg13g2_fill_1 FILLER_63_774 ();
 sg13g2_decap_8 FILLER_63_784 ();
 sg13g2_decap_8 FILLER_63_791 ();
 sg13g2_decap_8 FILLER_63_798 ();
 sg13g2_decap_8 FILLER_63_805 ();
 sg13g2_decap_8 FILLER_63_812 ();
 sg13g2_decap_8 FILLER_63_819 ();
 sg13g2_decap_8 FILLER_63_826 ();
 sg13g2_decap_8 FILLER_63_833 ();
 sg13g2_decap_4 FILLER_63_840 ();
 sg13g2_fill_2 FILLER_63_844 ();
 sg13g2_fill_2 FILLER_63_850 ();
 sg13g2_decap_4 FILLER_63_858 ();
 sg13g2_fill_1 FILLER_63_862 ();
 sg13g2_decap_8 FILLER_63_878 ();
 sg13g2_fill_1 FILLER_63_885 ();
 sg13g2_decap_8 FILLER_63_891 ();
 sg13g2_fill_1 FILLER_63_908 ();
 sg13g2_fill_1 FILLER_63_923 ();
 sg13g2_fill_1 FILLER_63_938 ();
 sg13g2_fill_2 FILLER_63_944 ();
 sg13g2_decap_8 FILLER_63_951 ();
 sg13g2_decap_8 FILLER_63_958 ();
 sg13g2_decap_8 FILLER_63_965 ();
 sg13g2_fill_2 FILLER_63_972 ();
 sg13g2_fill_1 FILLER_63_974 ();
 sg13g2_decap_8 FILLER_63_980 ();
 sg13g2_fill_2 FILLER_63_987 ();
 sg13g2_decap_8 FILLER_63_993 ();
 sg13g2_decap_8 FILLER_63_1000 ();
 sg13g2_decap_8 FILLER_63_1011 ();
 sg13g2_fill_2 FILLER_63_1018 ();
 sg13g2_fill_1 FILLER_63_1020 ();
 sg13g2_decap_8 FILLER_63_1026 ();
 sg13g2_fill_1 FILLER_63_1033 ();
 sg13g2_decap_8 FILLER_63_1039 ();
 sg13g2_decap_8 FILLER_63_1046 ();
 sg13g2_decap_4 FILLER_63_1057 ();
 sg13g2_fill_2 FILLER_63_1061 ();
 sg13g2_decap_8 FILLER_63_1067 ();
 sg13g2_fill_2 FILLER_63_1074 ();
 sg13g2_fill_1 FILLER_63_1076 ();
 sg13g2_fill_1 FILLER_63_1082 ();
 sg13g2_decap_4 FILLER_63_1088 ();
 sg13g2_fill_2 FILLER_63_1092 ();
 sg13g2_decap_8 FILLER_63_1098 ();
 sg13g2_decap_8 FILLER_63_1105 ();
 sg13g2_fill_1 FILLER_63_1112 ();
 sg13g2_fill_2 FILLER_63_1130 ();
 sg13g2_fill_1 FILLER_63_1137 ();
 sg13g2_fill_1 FILLER_63_1143 ();
 sg13g2_decap_8 FILLER_63_1149 ();
 sg13g2_decap_8 FILLER_63_1156 ();
 sg13g2_decap_4 FILLER_63_1163 ();
 sg13g2_fill_2 FILLER_63_1172 ();
 sg13g2_fill_1 FILLER_63_1174 ();
 sg13g2_fill_2 FILLER_63_1186 ();
 sg13g2_fill_1 FILLER_63_1188 ();
 sg13g2_fill_2 FILLER_63_1194 ();
 sg13g2_fill_1 FILLER_63_1196 ();
 sg13g2_fill_2 FILLER_63_1207 ();
 sg13g2_fill_1 FILLER_63_1209 ();
 sg13g2_decap_8 FILLER_63_1219 ();
 sg13g2_decap_8 FILLER_63_1226 ();
 sg13g2_decap_8 FILLER_63_1246 ();
 sg13g2_decap_4 FILLER_63_1258 ();
 sg13g2_fill_1 FILLER_63_1262 ();
 sg13g2_decap_8 FILLER_63_1289 ();
 sg13g2_decap_8 FILLER_63_1296 ();
 sg13g2_decap_8 FILLER_63_1303 ();
 sg13g2_decap_8 FILLER_63_1310 ();
 sg13g2_decap_8 FILLER_63_1317 ();
 sg13g2_fill_2 FILLER_63_1324 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_40 ();
 sg13g2_decap_8 FILLER_64_47 ();
 sg13g2_decap_8 FILLER_64_54 ();
 sg13g2_decap_4 FILLER_64_61 ();
 sg13g2_fill_1 FILLER_64_65 ();
 sg13g2_decap_8 FILLER_64_75 ();
 sg13g2_decap_8 FILLER_64_82 ();
 sg13g2_decap_8 FILLER_64_89 ();
 sg13g2_decap_8 FILLER_64_96 ();
 sg13g2_decap_8 FILLER_64_103 ();
 sg13g2_decap_4 FILLER_64_110 ();
 sg13g2_decap_8 FILLER_64_129 ();
 sg13g2_decap_8 FILLER_64_136 ();
 sg13g2_decap_8 FILLER_64_143 ();
 sg13g2_fill_1 FILLER_64_150 ();
 sg13g2_fill_2 FILLER_64_164 ();
 sg13g2_fill_1 FILLER_64_166 ();
 sg13g2_decap_4 FILLER_64_172 ();
 sg13g2_fill_2 FILLER_64_181 ();
 sg13g2_decap_8 FILLER_64_188 ();
 sg13g2_decap_8 FILLER_64_195 ();
 sg13g2_decap_8 FILLER_64_202 ();
 sg13g2_decap_8 FILLER_64_209 ();
 sg13g2_decap_4 FILLER_64_216 ();
 sg13g2_fill_2 FILLER_64_235 ();
 sg13g2_fill_2 FILLER_64_245 ();
 sg13g2_fill_1 FILLER_64_247 ();
 sg13g2_fill_2 FILLER_64_253 ();
 sg13g2_fill_1 FILLER_64_255 ();
 sg13g2_fill_2 FILLER_64_268 ();
 sg13g2_decap_8 FILLER_64_280 ();
 sg13g2_decap_4 FILLER_64_287 ();
 sg13g2_fill_1 FILLER_64_291 ();
 sg13g2_fill_1 FILLER_64_307 ();
 sg13g2_decap_8 FILLER_64_326 ();
 sg13g2_decap_4 FILLER_64_333 ();
 sg13g2_decap_4 FILLER_64_341 ();
 sg13g2_decap_8 FILLER_64_371 ();
 sg13g2_decap_8 FILLER_64_378 ();
 sg13g2_decap_4 FILLER_64_385 ();
 sg13g2_fill_2 FILLER_64_389 ();
 sg13g2_fill_2 FILLER_64_417 ();
 sg13g2_fill_1 FILLER_64_423 ();
 sg13g2_decap_8 FILLER_64_428 ();
 sg13g2_decap_8 FILLER_64_435 ();
 sg13g2_decap_8 FILLER_64_442 ();
 sg13g2_decap_8 FILLER_64_480 ();
 sg13g2_decap_8 FILLER_64_487 ();
 sg13g2_decap_8 FILLER_64_494 ();
 sg13g2_decap_8 FILLER_64_501 ();
 sg13g2_fill_2 FILLER_64_508 ();
 sg13g2_decap_8 FILLER_64_518 ();
 sg13g2_decap_8 FILLER_64_525 ();
 sg13g2_decap_4 FILLER_64_532 ();
 sg13g2_fill_2 FILLER_64_536 ();
 sg13g2_decap_4 FILLER_64_542 ();
 sg13g2_decap_8 FILLER_64_550 ();
 sg13g2_decap_8 FILLER_64_557 ();
 sg13g2_decap_8 FILLER_64_564 ();
 sg13g2_decap_8 FILLER_64_571 ();
 sg13g2_decap_8 FILLER_64_578 ();
 sg13g2_decap_8 FILLER_64_585 ();
 sg13g2_decap_8 FILLER_64_596 ();
 sg13g2_decap_8 FILLER_64_603 ();
 sg13g2_decap_8 FILLER_64_610 ();
 sg13g2_decap_4 FILLER_64_651 ();
 sg13g2_fill_1 FILLER_64_659 ();
 sg13g2_decap_4 FILLER_64_664 ();
 sg13g2_fill_2 FILLER_64_668 ();
 sg13g2_decap_4 FILLER_64_679 ();
 sg13g2_fill_2 FILLER_64_687 ();
 sg13g2_fill_1 FILLER_64_689 ();
 sg13g2_decap_4 FILLER_64_695 ();
 sg13g2_fill_1 FILLER_64_699 ();
 sg13g2_decap_8 FILLER_64_708 ();
 sg13g2_fill_1 FILLER_64_715 ();
 sg13g2_decap_8 FILLER_64_724 ();
 sg13g2_decap_8 FILLER_64_731 ();
 sg13g2_decap_8 FILLER_64_738 ();
 sg13g2_decap_8 FILLER_64_745 ();
 sg13g2_decap_4 FILLER_64_752 ();
 sg13g2_fill_2 FILLER_64_767 ();
 sg13g2_decap_8 FILLER_64_774 ();
 sg13g2_decap_8 FILLER_64_781 ();
 sg13g2_decap_8 FILLER_64_788 ();
 sg13g2_decap_8 FILLER_64_795 ();
 sg13g2_decap_8 FILLER_64_802 ();
 sg13g2_decap_8 FILLER_64_809 ();
 sg13g2_decap_8 FILLER_64_816 ();
 sg13g2_decap_8 FILLER_64_823 ();
 sg13g2_decap_8 FILLER_64_830 ();
 sg13g2_decap_8 FILLER_64_837 ();
 sg13g2_decap_8 FILLER_64_844 ();
 sg13g2_decap_8 FILLER_64_851 ();
 sg13g2_decap_8 FILLER_64_858 ();
 sg13g2_decap_8 FILLER_64_865 ();
 sg13g2_decap_4 FILLER_64_872 ();
 sg13g2_fill_2 FILLER_64_876 ();
 sg13g2_decap_8 FILLER_64_882 ();
 sg13g2_decap_8 FILLER_64_889 ();
 sg13g2_decap_4 FILLER_64_896 ();
 sg13g2_fill_2 FILLER_64_900 ();
 sg13g2_decap_4 FILLER_64_907 ();
 sg13g2_fill_1 FILLER_64_911 ();
 sg13g2_decap_8 FILLER_64_922 ();
 sg13g2_fill_2 FILLER_64_929 ();
 sg13g2_fill_1 FILLER_64_931 ();
 sg13g2_decap_4 FILLER_64_948 ();
 sg13g2_fill_1 FILLER_64_952 ();
 sg13g2_fill_2 FILLER_64_957 ();
 sg13g2_fill_1 FILLER_64_959 ();
 sg13g2_decap_8 FILLER_64_985 ();
 sg13g2_decap_8 FILLER_64_992 ();
 sg13g2_decap_8 FILLER_64_999 ();
 sg13g2_fill_1 FILLER_64_1019 ();
 sg13g2_decap_8 FILLER_64_1024 ();
 sg13g2_decap_8 FILLER_64_1031 ();
 sg13g2_fill_1 FILLER_64_1046 ();
 sg13g2_decap_4 FILLER_64_1058 ();
 sg13g2_fill_2 FILLER_64_1062 ();
 sg13g2_decap_8 FILLER_64_1069 ();
 sg13g2_decap_8 FILLER_64_1076 ();
 sg13g2_decap_8 FILLER_64_1083 ();
 sg13g2_decap_4 FILLER_64_1090 ();
 sg13g2_fill_1 FILLER_64_1094 ();
 sg13g2_decap_8 FILLER_64_1100 ();
 sg13g2_decap_4 FILLER_64_1107 ();
 sg13g2_fill_1 FILLER_64_1111 ();
 sg13g2_fill_1 FILLER_64_1121 ();
 sg13g2_fill_2 FILLER_64_1127 ();
 sg13g2_fill_1 FILLER_64_1129 ();
 sg13g2_decap_8 FILLER_64_1135 ();
 sg13g2_decap_4 FILLER_64_1142 ();
 sg13g2_fill_2 FILLER_64_1146 ();
 sg13g2_decap_8 FILLER_64_1159 ();
 sg13g2_decap_4 FILLER_64_1166 ();
 sg13g2_fill_1 FILLER_64_1170 ();
 sg13g2_decap_8 FILLER_64_1181 ();
 sg13g2_decap_8 FILLER_64_1188 ();
 sg13g2_fill_2 FILLER_64_1195 ();
 sg13g2_fill_1 FILLER_64_1197 ();
 sg13g2_decap_4 FILLER_64_1208 ();
 sg13g2_fill_1 FILLER_64_1212 ();
 sg13g2_decap_4 FILLER_64_1228 ();
 sg13g2_fill_2 FILLER_64_1232 ();
 sg13g2_fill_2 FILLER_64_1255 ();
 sg13g2_decap_8 FILLER_64_1261 ();
 sg13g2_fill_1 FILLER_64_1268 ();
 sg13g2_decap_4 FILLER_64_1276 ();
 sg13g2_fill_2 FILLER_64_1280 ();
 sg13g2_decap_8 FILLER_64_1286 ();
 sg13g2_decap_8 FILLER_64_1293 ();
 sg13g2_decap_8 FILLER_64_1300 ();
 sg13g2_decap_8 FILLER_64_1307 ();
 sg13g2_decap_8 FILLER_64_1314 ();
 sg13g2_decap_4 FILLER_64_1321 ();
 sg13g2_fill_1 FILLER_64_1325 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_4 FILLER_65_35 ();
 sg13g2_fill_1 FILLER_65_39 ();
 sg13g2_fill_2 FILLER_65_65 ();
 sg13g2_fill_1 FILLER_65_67 ();
 sg13g2_fill_1 FILLER_65_73 ();
 sg13g2_decap_4 FILLER_65_97 ();
 sg13g2_decap_8 FILLER_65_106 ();
 sg13g2_decap_8 FILLER_65_113 ();
 sg13g2_decap_4 FILLER_65_120 ();
 sg13g2_fill_2 FILLER_65_124 ();
 sg13g2_decap_4 FILLER_65_131 ();
 sg13g2_fill_1 FILLER_65_135 ();
 sg13g2_decap_8 FILLER_65_141 ();
 sg13g2_decap_8 FILLER_65_183 ();
 sg13g2_decap_8 FILLER_65_190 ();
 sg13g2_decap_8 FILLER_65_197 ();
 sg13g2_decap_8 FILLER_65_204 ();
 sg13g2_decap_8 FILLER_65_211 ();
 sg13g2_decap_8 FILLER_65_218 ();
 sg13g2_fill_2 FILLER_65_225 ();
 sg13g2_fill_1 FILLER_65_233 ();
 sg13g2_decap_8 FILLER_65_243 ();
 sg13g2_decap_8 FILLER_65_250 ();
 sg13g2_decap_8 FILLER_65_257 ();
 sg13g2_decap_8 FILLER_65_264 ();
 sg13g2_decap_8 FILLER_65_271 ();
 sg13g2_decap_8 FILLER_65_278 ();
 sg13g2_decap_8 FILLER_65_285 ();
 sg13g2_fill_2 FILLER_65_292 ();
 sg13g2_decap_8 FILLER_65_303 ();
 sg13g2_decap_8 FILLER_65_310 ();
 sg13g2_decap_8 FILLER_65_317 ();
 sg13g2_decap_8 FILLER_65_329 ();
 sg13g2_decap_8 FILLER_65_336 ();
 sg13g2_decap_8 FILLER_65_343 ();
 sg13g2_fill_1 FILLER_65_350 ();
 sg13g2_decap_4 FILLER_65_355 ();
 sg13g2_fill_2 FILLER_65_359 ();
 sg13g2_decap_8 FILLER_65_365 ();
 sg13g2_decap_8 FILLER_65_372 ();
 sg13g2_decap_8 FILLER_65_379 ();
 sg13g2_decap_8 FILLER_65_386 ();
 sg13g2_decap_8 FILLER_65_393 ();
 sg13g2_decap_4 FILLER_65_409 ();
 sg13g2_fill_2 FILLER_65_413 ();
 sg13g2_decap_8 FILLER_65_431 ();
 sg13g2_decap_8 FILLER_65_438 ();
 sg13g2_decap_8 FILLER_65_445 ();
 sg13g2_decap_8 FILLER_65_452 ();
 sg13g2_fill_1 FILLER_65_459 ();
 sg13g2_decap_8 FILLER_65_486 ();
 sg13g2_decap_4 FILLER_65_498 ();
 sg13g2_decap_8 FILLER_65_564 ();
 sg13g2_decap_8 FILLER_65_571 ();
 sg13g2_decap_8 FILLER_65_578 ();
 sg13g2_decap_8 FILLER_65_585 ();
 sg13g2_decap_8 FILLER_65_592 ();
 sg13g2_decap_8 FILLER_65_599 ();
 sg13g2_decap_8 FILLER_65_606 ();
 sg13g2_decap_8 FILLER_65_613 ();
 sg13g2_decap_4 FILLER_65_620 ();
 sg13g2_fill_1 FILLER_65_624 ();
 sg13g2_decap_8 FILLER_65_629 ();
 sg13g2_decap_8 FILLER_65_636 ();
 sg13g2_decap_8 FILLER_65_647 ();
 sg13g2_decap_8 FILLER_65_654 ();
 sg13g2_decap_8 FILLER_65_661 ();
 sg13g2_decap_8 FILLER_65_668 ();
 sg13g2_decap_8 FILLER_65_675 ();
 sg13g2_decap_8 FILLER_65_682 ();
 sg13g2_decap_8 FILLER_65_689 ();
 sg13g2_decap_4 FILLER_65_696 ();
 sg13g2_fill_1 FILLER_65_700 ();
 sg13g2_fill_1 FILLER_65_706 ();
 sg13g2_fill_2 FILLER_65_711 ();
 sg13g2_decap_8 FILLER_65_729 ();
 sg13g2_decap_8 FILLER_65_736 ();
 sg13g2_decap_8 FILLER_65_743 ();
 sg13g2_decap_8 FILLER_65_750 ();
 sg13g2_fill_2 FILLER_65_757 ();
 sg13g2_decap_4 FILLER_65_763 ();
 sg13g2_fill_1 FILLER_65_767 ();
 sg13g2_decap_8 FILLER_65_786 ();
 sg13g2_decap_4 FILLER_65_793 ();
 sg13g2_fill_1 FILLER_65_797 ();
 sg13g2_decap_8 FILLER_65_803 ();
 sg13g2_decap_8 FILLER_65_810 ();
 sg13g2_decap_8 FILLER_65_817 ();
 sg13g2_decap_8 FILLER_65_824 ();
 sg13g2_decap_8 FILLER_65_831 ();
 sg13g2_decap_8 FILLER_65_838 ();
 sg13g2_decap_8 FILLER_65_845 ();
 sg13g2_decap_8 FILLER_65_852 ();
 sg13g2_decap_8 FILLER_65_859 ();
 sg13g2_decap_8 FILLER_65_866 ();
 sg13g2_decap_8 FILLER_65_873 ();
 sg13g2_decap_8 FILLER_65_880 ();
 sg13g2_decap_8 FILLER_65_887 ();
 sg13g2_decap_8 FILLER_65_894 ();
 sg13g2_decap_8 FILLER_65_901 ();
 sg13g2_decap_8 FILLER_65_908 ();
 sg13g2_decap_4 FILLER_65_915 ();
 sg13g2_decap_8 FILLER_65_924 ();
 sg13g2_decap_8 FILLER_65_931 ();
 sg13g2_fill_1 FILLER_65_938 ();
 sg13g2_decap_8 FILLER_65_947 ();
 sg13g2_decap_4 FILLER_65_959 ();
 sg13g2_fill_2 FILLER_65_963 ();
 sg13g2_fill_1 FILLER_65_969 ();
 sg13g2_decap_4 FILLER_65_976 ();
 sg13g2_fill_2 FILLER_65_985 ();
 sg13g2_decap_8 FILLER_65_996 ();
 sg13g2_decap_4 FILLER_65_1003 ();
 sg13g2_fill_2 FILLER_65_1007 ();
 sg13g2_decap_8 FILLER_65_1021 ();
 sg13g2_decap_8 FILLER_65_1028 ();
 sg13g2_fill_1 FILLER_65_1040 ();
 sg13g2_decap_8 FILLER_65_1045 ();
 sg13g2_decap_4 FILLER_65_1057 ();
 sg13g2_fill_1 FILLER_65_1061 ();
 sg13g2_decap_4 FILLER_65_1074 ();
 sg13g2_decap_8 FILLER_65_1088 ();
 sg13g2_decap_4 FILLER_65_1095 ();
 sg13g2_decap_8 FILLER_65_1103 ();
 sg13g2_decap_4 FILLER_65_1110 ();
 sg13g2_fill_1 FILLER_65_1114 ();
 sg13g2_decap_4 FILLER_65_1131 ();
 sg13g2_fill_2 FILLER_65_1135 ();
 sg13g2_decap_8 FILLER_65_1144 ();
 sg13g2_fill_2 FILLER_65_1151 ();
 sg13g2_fill_1 FILLER_65_1153 ();
 sg13g2_fill_2 FILLER_65_1158 ();
 sg13g2_fill_1 FILLER_65_1160 ();
 sg13g2_decap_8 FILLER_65_1166 ();
 sg13g2_fill_2 FILLER_65_1173 ();
 sg13g2_fill_1 FILLER_65_1180 ();
 sg13g2_decap_8 FILLER_65_1186 ();
 sg13g2_decap_4 FILLER_65_1193 ();
 sg13g2_decap_8 FILLER_65_1201 ();
 sg13g2_decap_8 FILLER_65_1216 ();
 sg13g2_decap_8 FILLER_65_1223 ();
 sg13g2_decap_8 FILLER_65_1230 ();
 sg13g2_decap_8 FILLER_65_1237 ();
 sg13g2_decap_8 FILLER_65_1244 ();
 sg13g2_decap_8 FILLER_65_1251 ();
 sg13g2_decap_8 FILLER_65_1258 ();
 sg13g2_fill_2 FILLER_65_1265 ();
 sg13g2_fill_1 FILLER_65_1267 ();
 sg13g2_decap_8 FILLER_65_1277 ();
 sg13g2_decap_8 FILLER_65_1294 ();
 sg13g2_decap_8 FILLER_65_1301 ();
 sg13g2_decap_8 FILLER_65_1308 ();
 sg13g2_decap_8 FILLER_65_1315 ();
 sg13g2_decap_4 FILLER_65_1322 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_fill_2 FILLER_66_42 ();
 sg13g2_fill_1 FILLER_66_44 ();
 sg13g2_fill_2 FILLER_66_54 ();
 sg13g2_decap_8 FILLER_66_61 ();
 sg13g2_decap_8 FILLER_66_68 ();
 sg13g2_decap_8 FILLER_66_75 ();
 sg13g2_decap_8 FILLER_66_82 ();
 sg13g2_decap_4 FILLER_66_89 ();
 sg13g2_fill_2 FILLER_66_93 ();
 sg13g2_fill_1 FILLER_66_99 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_decap_4 FILLER_66_147 ();
 sg13g2_fill_1 FILLER_66_151 ();
 sg13g2_fill_2 FILLER_66_156 ();
 sg13g2_fill_1 FILLER_66_163 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_decap_4 FILLER_66_182 ();
 sg13g2_decap_8 FILLER_66_221 ();
 sg13g2_decap_8 FILLER_66_228 ();
 sg13g2_decap_8 FILLER_66_235 ();
 sg13g2_decap_8 FILLER_66_242 ();
 sg13g2_decap_8 FILLER_66_249 ();
 sg13g2_decap_8 FILLER_66_256 ();
 sg13g2_decap_8 FILLER_66_263 ();
 sg13g2_fill_2 FILLER_66_270 ();
 sg13g2_decap_8 FILLER_66_275 ();
 sg13g2_decap_8 FILLER_66_282 ();
 sg13g2_fill_2 FILLER_66_289 ();
 sg13g2_decap_4 FILLER_66_301 ();
 sg13g2_fill_1 FILLER_66_305 ();
 sg13g2_fill_2 FILLER_66_324 ();
 sg13g2_decap_8 FILLER_66_357 ();
 sg13g2_fill_2 FILLER_66_364 ();
 sg13g2_decap_8 FILLER_66_370 ();
 sg13g2_decap_8 FILLER_66_377 ();
 sg13g2_decap_8 FILLER_66_384 ();
 sg13g2_fill_2 FILLER_66_391 ();
 sg13g2_decap_4 FILLER_66_423 ();
 sg13g2_fill_2 FILLER_66_427 ();
 sg13g2_decap_8 FILLER_66_434 ();
 sg13g2_decap_8 FILLER_66_441 ();
 sg13g2_decap_8 FILLER_66_448 ();
 sg13g2_decap_4 FILLER_66_455 ();
 sg13g2_fill_1 FILLER_66_459 ();
 sg13g2_decap_8 FILLER_66_490 ();
 sg13g2_decap_8 FILLER_66_497 ();
 sg13g2_decap_8 FILLER_66_504 ();
 sg13g2_fill_2 FILLER_66_511 ();
 sg13g2_decap_8 FILLER_66_517 ();
 sg13g2_decap_8 FILLER_66_524 ();
 sg13g2_decap_8 FILLER_66_531 ();
 sg13g2_decap_8 FILLER_66_538 ();
 sg13g2_decap_8 FILLER_66_545 ();
 sg13g2_decap_8 FILLER_66_552 ();
 sg13g2_decap_8 FILLER_66_559 ();
 sg13g2_decap_8 FILLER_66_566 ();
 sg13g2_fill_2 FILLER_66_573 ();
 sg13g2_fill_1 FILLER_66_575 ();
 sg13g2_decap_4 FILLER_66_581 ();
 sg13g2_fill_2 FILLER_66_585 ();
 sg13g2_decap_8 FILLER_66_591 ();
 sg13g2_decap_8 FILLER_66_598 ();
 sg13g2_decap_8 FILLER_66_605 ();
 sg13g2_decap_8 FILLER_66_612 ();
 sg13g2_decap_8 FILLER_66_619 ();
 sg13g2_fill_1 FILLER_66_633 ();
 sg13g2_fill_2 FILLER_66_639 ();
 sg13g2_decap_8 FILLER_66_670 ();
 sg13g2_decap_8 FILLER_66_677 ();
 sg13g2_decap_4 FILLER_66_684 ();
 sg13g2_fill_2 FILLER_66_688 ();
 sg13g2_fill_1 FILLER_66_699 ();
 sg13g2_decap_8 FILLER_66_730 ();
 sg13g2_fill_2 FILLER_66_737 ();
 sg13g2_decap_8 FILLER_66_769 ();
 sg13g2_decap_8 FILLER_66_776 ();
 sg13g2_fill_2 FILLER_66_783 ();
 sg13g2_decap_8 FILLER_66_811 ();
 sg13g2_decap_8 FILLER_66_818 ();
 sg13g2_decap_8 FILLER_66_825 ();
 sg13g2_decap_8 FILLER_66_832 ();
 sg13g2_decap_8 FILLER_66_839 ();
 sg13g2_decap_8 FILLER_66_846 ();
 sg13g2_decap_8 FILLER_66_853 ();
 sg13g2_decap_8 FILLER_66_860 ();
 sg13g2_decap_8 FILLER_66_867 ();
 sg13g2_decap_4 FILLER_66_874 ();
 sg13g2_fill_2 FILLER_66_878 ();
 sg13g2_decap_8 FILLER_66_888 ();
 sg13g2_decap_4 FILLER_66_905 ();
 sg13g2_fill_1 FILLER_66_909 ();
 sg13g2_decap_8 FILLER_66_915 ();
 sg13g2_decap_8 FILLER_66_922 ();
 sg13g2_fill_2 FILLER_66_929 ();
 sg13g2_decap_8 FILLER_66_939 ();
 sg13g2_decap_4 FILLER_66_946 ();
 sg13g2_decap_8 FILLER_66_957 ();
 sg13g2_decap_8 FILLER_66_964 ();
 sg13g2_fill_1 FILLER_66_971 ();
 sg13g2_decap_8 FILLER_66_978 ();
 sg13g2_decap_4 FILLER_66_985 ();
 sg13g2_fill_2 FILLER_66_989 ();
 sg13g2_decap_8 FILLER_66_996 ();
 sg13g2_decap_8 FILLER_66_1003 ();
 sg13g2_fill_2 FILLER_66_1010 ();
 sg13g2_fill_1 FILLER_66_1012 ();
 sg13g2_decap_8 FILLER_66_1017 ();
 sg13g2_decap_8 FILLER_66_1024 ();
 sg13g2_decap_8 FILLER_66_1031 ();
 sg13g2_fill_1 FILLER_66_1038 ();
 sg13g2_fill_1 FILLER_66_1053 ();
 sg13g2_fill_1 FILLER_66_1064 ();
 sg13g2_decap_8 FILLER_66_1076 ();
 sg13g2_fill_2 FILLER_66_1083 ();
 sg13g2_decap_4 FILLER_66_1091 ();
 sg13g2_fill_1 FILLER_66_1095 ();
 sg13g2_decap_8 FILLER_66_1101 ();
 sg13g2_decap_8 FILLER_66_1108 ();
 sg13g2_decap_4 FILLER_66_1115 ();
 sg13g2_decap_8 FILLER_66_1124 ();
 sg13g2_decap_8 FILLER_66_1137 ();
 sg13g2_decap_8 FILLER_66_1144 ();
 sg13g2_decap_4 FILLER_66_1151 ();
 sg13g2_fill_2 FILLER_66_1160 ();
 sg13g2_fill_2 FILLER_66_1167 ();
 sg13g2_decap_8 FILLER_66_1177 ();
 sg13g2_decap_4 FILLER_66_1184 ();
 sg13g2_fill_2 FILLER_66_1188 ();
 sg13g2_decap_4 FILLER_66_1199 ();
 sg13g2_decap_4 FILLER_66_1227 ();
 sg13g2_fill_1 FILLER_66_1231 ();
 sg13g2_decap_8 FILLER_66_1236 ();
 sg13g2_fill_1 FILLER_66_1243 ();
 sg13g2_decap_8 FILLER_66_1257 ();
 sg13g2_fill_1 FILLER_66_1269 ();
 sg13g2_fill_1 FILLER_66_1274 ();
 sg13g2_decap_4 FILLER_66_1279 ();
 sg13g2_decap_8 FILLER_66_1288 ();
 sg13g2_decap_8 FILLER_66_1295 ();
 sg13g2_decap_8 FILLER_66_1302 ();
 sg13g2_decap_8 FILLER_66_1309 ();
 sg13g2_decap_8 FILLER_66_1316 ();
 sg13g2_fill_2 FILLER_66_1323 ();
 sg13g2_fill_1 FILLER_66_1325 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_fill_2 FILLER_67_35 ();
 sg13g2_fill_1 FILLER_67_37 ();
 sg13g2_decap_8 FILLER_67_64 ();
 sg13g2_decap_8 FILLER_67_71 ();
 sg13g2_fill_2 FILLER_67_78 ();
 sg13g2_fill_1 FILLER_67_80 ();
 sg13g2_fill_2 FILLER_67_85 ();
 sg13g2_decap_8 FILLER_67_127 ();
 sg13g2_decap_4 FILLER_67_134 ();
 sg13g2_decap_8 FILLER_67_156 ();
 sg13g2_decap_8 FILLER_67_163 ();
 sg13g2_decap_8 FILLER_67_170 ();
 sg13g2_decap_8 FILLER_67_177 ();
 sg13g2_decap_8 FILLER_67_184 ();
 sg13g2_fill_2 FILLER_67_191 ();
 sg13g2_fill_2 FILLER_67_200 ();
 sg13g2_decap_8 FILLER_67_206 ();
 sg13g2_fill_1 FILLER_67_213 ();
 sg13g2_decap_8 FILLER_67_219 ();
 sg13g2_decap_4 FILLER_67_226 ();
 sg13g2_fill_2 FILLER_67_230 ();
 sg13g2_fill_2 FILLER_67_240 ();
 sg13g2_decap_8 FILLER_67_247 ();
 sg13g2_decap_8 FILLER_67_254 ();
 sg13g2_fill_1 FILLER_67_261 ();
 sg13g2_decap_8 FILLER_67_275 ();
 sg13g2_decap_8 FILLER_67_282 ();
 sg13g2_decap_4 FILLER_67_289 ();
 sg13g2_fill_2 FILLER_67_293 ();
 sg13g2_decap_8 FILLER_67_300 ();
 sg13g2_decap_8 FILLER_67_307 ();
 sg13g2_fill_1 FILLER_67_314 ();
 sg13g2_decap_8 FILLER_67_320 ();
 sg13g2_decap_8 FILLER_67_327 ();
 sg13g2_fill_1 FILLER_67_334 ();
 sg13g2_decap_8 FILLER_67_339 ();
 sg13g2_decap_8 FILLER_67_346 ();
 sg13g2_decap_8 FILLER_67_353 ();
 sg13g2_decap_8 FILLER_67_360 ();
 sg13g2_fill_2 FILLER_67_367 ();
 sg13g2_decap_8 FILLER_67_373 ();
 sg13g2_decap_8 FILLER_67_380 ();
 sg13g2_decap_4 FILLER_67_387 ();
 sg13g2_fill_1 FILLER_67_391 ();
 sg13g2_decap_4 FILLER_67_397 ();
 sg13g2_fill_1 FILLER_67_401 ();
 sg13g2_fill_1 FILLER_67_407 ();
 sg13g2_fill_2 FILLER_67_412 ();
 sg13g2_fill_2 FILLER_67_420 ();
 sg13g2_decap_8 FILLER_67_438 ();
 sg13g2_decap_8 FILLER_67_445 ();
 sg13g2_decap_8 FILLER_67_452 ();
 sg13g2_decap_8 FILLER_67_459 ();
 sg13g2_decap_4 FILLER_67_466 ();
 sg13g2_fill_1 FILLER_67_470 ();
 sg13g2_decap_8 FILLER_67_475 ();
 sg13g2_decap_8 FILLER_67_482 ();
 sg13g2_decap_8 FILLER_67_489 ();
 sg13g2_decap_8 FILLER_67_496 ();
 sg13g2_decap_8 FILLER_67_503 ();
 sg13g2_decap_8 FILLER_67_510 ();
 sg13g2_decap_8 FILLER_67_517 ();
 sg13g2_decap_8 FILLER_67_524 ();
 sg13g2_decap_8 FILLER_67_539 ();
 sg13g2_decap_4 FILLER_67_546 ();
 sg13g2_fill_2 FILLER_67_576 ();
 sg13g2_decap_8 FILLER_67_604 ();
 sg13g2_decap_4 FILLER_67_611 ();
 sg13g2_fill_1 FILLER_67_615 ();
 sg13g2_fill_2 FILLER_67_642 ();
 sg13g2_fill_1 FILLER_67_644 ();
 sg13g2_fill_1 FILLER_67_652 ();
 sg13g2_fill_2 FILLER_67_658 ();
 sg13g2_fill_1 FILLER_67_660 ();
 sg13g2_decap_8 FILLER_67_666 ();
 sg13g2_decap_8 FILLER_67_673 ();
 sg13g2_decap_4 FILLER_67_680 ();
 sg13g2_decap_8 FILLER_67_714 ();
 sg13g2_decap_8 FILLER_67_721 ();
 sg13g2_fill_2 FILLER_67_728 ();
 sg13g2_fill_1 FILLER_67_730 ();
 sg13g2_decap_8 FILLER_67_735 ();
 sg13g2_decap_4 FILLER_67_742 ();
 sg13g2_decap_8 FILLER_67_750 ();
 sg13g2_fill_1 FILLER_67_786 ();
 sg13g2_decap_4 FILLER_67_824 ();
 sg13g2_fill_1 FILLER_67_828 ();
 sg13g2_decap_8 FILLER_67_834 ();
 sg13g2_decap_8 FILLER_67_841 ();
 sg13g2_decap_8 FILLER_67_848 ();
 sg13g2_decap_8 FILLER_67_855 ();
 sg13g2_decap_8 FILLER_67_862 ();
 sg13g2_fill_2 FILLER_67_869 ();
 sg13g2_decap_8 FILLER_67_876 ();
 sg13g2_fill_1 FILLER_67_893 ();
 sg13g2_decap_4 FILLER_67_898 ();
 sg13g2_decap_4 FILLER_67_906 ();
 sg13g2_fill_1 FILLER_67_910 ();
 sg13g2_fill_1 FILLER_67_916 ();
 sg13g2_fill_1 FILLER_67_922 ();
 sg13g2_decap_4 FILLER_67_938 ();
 sg13g2_fill_2 FILLER_67_942 ();
 sg13g2_decap_4 FILLER_67_949 ();
 sg13g2_fill_2 FILLER_67_953 ();
 sg13g2_decap_4 FILLER_67_959 ();
 sg13g2_fill_2 FILLER_67_963 ();
 sg13g2_fill_2 FILLER_67_975 ();
 sg13g2_decap_8 FILLER_67_982 ();
 sg13g2_decap_8 FILLER_67_989 ();
 sg13g2_fill_2 FILLER_67_996 ();
 sg13g2_fill_1 FILLER_67_998 ();
 sg13g2_fill_2 FILLER_67_1014 ();
 sg13g2_decap_8 FILLER_67_1021 ();
 sg13g2_fill_1 FILLER_67_1028 ();
 sg13g2_fill_2 FILLER_67_1034 ();
 sg13g2_fill_2 FILLER_67_1045 ();
 sg13g2_fill_1 FILLER_67_1052 ();
 sg13g2_decap_4 FILLER_67_1058 ();
 sg13g2_fill_1 FILLER_67_1062 ();
 sg13g2_fill_2 FILLER_67_1067 ();
 sg13g2_decap_4 FILLER_67_1075 ();
 sg13g2_fill_1 FILLER_67_1079 ();
 sg13g2_decap_4 FILLER_67_1087 ();
 sg13g2_fill_1 FILLER_67_1091 ();
 sg13g2_decap_8 FILLER_67_1097 ();
 sg13g2_decap_8 FILLER_67_1104 ();
 sg13g2_decap_8 FILLER_67_1111 ();
 sg13g2_fill_2 FILLER_67_1118 ();
 sg13g2_fill_1 FILLER_67_1120 ();
 sg13g2_fill_2 FILLER_67_1126 ();
 sg13g2_fill_1 FILLER_67_1128 ();
 sg13g2_decap_8 FILLER_67_1133 ();
 sg13g2_fill_2 FILLER_67_1140 ();
 sg13g2_fill_1 FILLER_67_1142 ();
 sg13g2_decap_8 FILLER_67_1148 ();
 sg13g2_fill_2 FILLER_67_1155 ();
 sg13g2_fill_2 FILLER_67_1162 ();
 sg13g2_fill_1 FILLER_67_1164 ();
 sg13g2_fill_2 FILLER_67_1172 ();
 sg13g2_decap_8 FILLER_67_1179 ();
 sg13g2_decap_8 FILLER_67_1186 ();
 sg13g2_decap_4 FILLER_67_1193 ();
 sg13g2_fill_1 FILLER_67_1197 ();
 sg13g2_fill_1 FILLER_67_1207 ();
 sg13g2_decap_4 FILLER_67_1213 ();
 sg13g2_fill_2 FILLER_67_1217 ();
 sg13g2_decap_8 FILLER_67_1223 ();
 sg13g2_fill_2 FILLER_67_1230 ();
 sg13g2_fill_2 FILLER_67_1249 ();
 sg13g2_decap_4 FILLER_67_1260 ();
 sg13g2_fill_2 FILLER_67_1269 ();
 sg13g2_decap_8 FILLER_67_1285 ();
 sg13g2_decap_8 FILLER_67_1292 ();
 sg13g2_decap_8 FILLER_67_1299 ();
 sg13g2_decap_8 FILLER_67_1306 ();
 sg13g2_decap_8 FILLER_67_1313 ();
 sg13g2_decap_4 FILLER_67_1320 ();
 sg13g2_fill_2 FILLER_67_1324 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_fill_2 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_82 ();
 sg13g2_fill_2 FILLER_68_89 ();
 sg13g2_fill_2 FILLER_68_103 ();
 sg13g2_decap_8 FILLER_68_109 ();
 sg13g2_decap_8 FILLER_68_120 ();
 sg13g2_fill_2 FILLER_68_127 ();
 sg13g2_fill_1 FILLER_68_129 ();
 sg13g2_fill_1 FILLER_68_139 ();
 sg13g2_decap_8 FILLER_68_150 ();
 sg13g2_decap_8 FILLER_68_157 ();
 sg13g2_decap_8 FILLER_68_164 ();
 sg13g2_decap_8 FILLER_68_176 ();
 sg13g2_decap_8 FILLER_68_183 ();
 sg13g2_decap_8 FILLER_68_190 ();
 sg13g2_decap_8 FILLER_68_197 ();
 sg13g2_decap_8 FILLER_68_204 ();
 sg13g2_decap_4 FILLER_68_211 ();
 sg13g2_fill_2 FILLER_68_215 ();
 sg13g2_fill_1 FILLER_68_221 ();
 sg13g2_fill_2 FILLER_68_245 ();
 sg13g2_fill_1 FILLER_68_254 ();
 sg13g2_fill_2 FILLER_68_273 ();
 sg13g2_decap_8 FILLER_68_301 ();
 sg13g2_decap_8 FILLER_68_308 ();
 sg13g2_decap_8 FILLER_68_315 ();
 sg13g2_decap_8 FILLER_68_322 ();
 sg13g2_decap_8 FILLER_68_329 ();
 sg13g2_fill_2 FILLER_68_336 ();
 sg13g2_decap_8 FILLER_68_346 ();
 sg13g2_decap_8 FILLER_68_353 ();
 sg13g2_decap_8 FILLER_68_360 ();
 sg13g2_fill_2 FILLER_68_367 ();
 sg13g2_decap_8 FILLER_68_374 ();
 sg13g2_decap_8 FILLER_68_381 ();
 sg13g2_decap_8 FILLER_68_388 ();
 sg13g2_decap_8 FILLER_68_395 ();
 sg13g2_decap_4 FILLER_68_402 ();
 sg13g2_fill_1 FILLER_68_406 ();
 sg13g2_fill_1 FILLER_68_421 ();
 sg13g2_fill_2 FILLER_68_427 ();
 sg13g2_decap_4 FILLER_68_459 ();
 sg13g2_fill_1 FILLER_68_463 ();
 sg13g2_decap_8 FILLER_68_469 ();
 sg13g2_decap_8 FILLER_68_476 ();
 sg13g2_decap_8 FILLER_68_483 ();
 sg13g2_decap_8 FILLER_68_490 ();
 sg13g2_decap_8 FILLER_68_497 ();
 sg13g2_decap_8 FILLER_68_504 ();
 sg13g2_decap_4 FILLER_68_511 ();
 sg13g2_fill_1 FILLER_68_515 ();
 sg13g2_decap_8 FILLER_68_550 ();
 sg13g2_decap_8 FILLER_68_561 ();
 sg13g2_decap_8 FILLER_68_568 ();
 sg13g2_decap_8 FILLER_68_575 ();
 sg13g2_decap_8 FILLER_68_582 ();
 sg13g2_decap_8 FILLER_68_589 ();
 sg13g2_decap_8 FILLER_68_596 ();
 sg13g2_decap_8 FILLER_68_603 ();
 sg13g2_decap_8 FILLER_68_610 ();
 sg13g2_decap_8 FILLER_68_617 ();
 sg13g2_decap_8 FILLER_68_628 ();
 sg13g2_fill_1 FILLER_68_635 ();
 sg13g2_decap_8 FILLER_68_662 ();
 sg13g2_decap_8 FILLER_68_669 ();
 sg13g2_decap_8 FILLER_68_676 ();
 sg13g2_decap_8 FILLER_68_683 ();
 sg13g2_decap_8 FILLER_68_690 ();
 sg13g2_decap_8 FILLER_68_697 ();
 sg13g2_decap_8 FILLER_68_704 ();
 sg13g2_decap_8 FILLER_68_711 ();
 sg13g2_decap_8 FILLER_68_718 ();
 sg13g2_decap_4 FILLER_68_751 ();
 sg13g2_fill_2 FILLER_68_755 ();
 sg13g2_fill_2 FILLER_68_769 ();
 sg13g2_fill_1 FILLER_68_771 ();
 sg13g2_decap_8 FILLER_68_777 ();
 sg13g2_decap_8 FILLER_68_784 ();
 sg13g2_decap_8 FILLER_68_791 ();
 sg13g2_fill_1 FILLER_68_798 ();
 sg13g2_decap_8 FILLER_68_834 ();
 sg13g2_decap_8 FILLER_68_841 ();
 sg13g2_decap_8 FILLER_68_848 ();
 sg13g2_decap_8 FILLER_68_855 ();
 sg13g2_decap_4 FILLER_68_862 ();
 sg13g2_fill_2 FILLER_68_866 ();
 sg13g2_decap_4 FILLER_68_877 ();
 sg13g2_fill_2 FILLER_68_886 ();
 sg13g2_fill_1 FILLER_68_909 ();
 sg13g2_decap_8 FILLER_68_914 ();
 sg13g2_fill_2 FILLER_68_921 ();
 sg13g2_fill_2 FILLER_68_932 ();
 sg13g2_fill_1 FILLER_68_944 ();
 sg13g2_decap_8 FILLER_68_950 ();
 sg13g2_decap_8 FILLER_68_957 ();
 sg13g2_decap_8 FILLER_68_964 ();
 sg13g2_decap_8 FILLER_68_971 ();
 sg13g2_decap_8 FILLER_68_978 ();
 sg13g2_decap_8 FILLER_68_985 ();
 sg13g2_decap_8 FILLER_68_992 ();
 sg13g2_fill_1 FILLER_68_999 ();
 sg13g2_decap_8 FILLER_68_1005 ();
 sg13g2_decap_8 FILLER_68_1012 ();
 sg13g2_decap_8 FILLER_68_1019 ();
 sg13g2_decap_8 FILLER_68_1026 ();
 sg13g2_decap_8 FILLER_68_1033 ();
 sg13g2_fill_2 FILLER_68_1040 ();
 sg13g2_fill_1 FILLER_68_1042 ();
 sg13g2_decap_4 FILLER_68_1048 ();
 sg13g2_fill_2 FILLER_68_1052 ();
 sg13g2_decap_8 FILLER_68_1058 ();
 sg13g2_decap_8 FILLER_68_1065 ();
 sg13g2_decap_4 FILLER_68_1072 ();
 sg13g2_fill_2 FILLER_68_1082 ();
 sg13g2_fill_1 FILLER_68_1084 ();
 sg13g2_decap_8 FILLER_68_1090 ();
 sg13g2_decap_8 FILLER_68_1097 ();
 sg13g2_decap_8 FILLER_68_1104 ();
 sg13g2_decap_4 FILLER_68_1111 ();
 sg13g2_decap_8 FILLER_68_1120 ();
 sg13g2_decap_8 FILLER_68_1127 ();
 sg13g2_decap_8 FILLER_68_1134 ();
 sg13g2_decap_8 FILLER_68_1141 ();
 sg13g2_decap_8 FILLER_68_1148 ();
 sg13g2_decap_4 FILLER_68_1155 ();
 sg13g2_decap_8 FILLER_68_1164 ();
 sg13g2_decap_8 FILLER_68_1179 ();
 sg13g2_decap_8 FILLER_68_1186 ();
 sg13g2_decap_8 FILLER_68_1193 ();
 sg13g2_decap_8 FILLER_68_1212 ();
 sg13g2_decap_4 FILLER_68_1219 ();
 sg13g2_fill_2 FILLER_68_1223 ();
 sg13g2_decap_8 FILLER_68_1236 ();
 sg13g2_decap_8 FILLER_68_1243 ();
 sg13g2_decap_4 FILLER_68_1250 ();
 sg13g2_decap_8 FILLER_68_1262 ();
 sg13g2_decap_8 FILLER_68_1269 ();
 sg13g2_decap_8 FILLER_68_1276 ();
 sg13g2_decap_8 FILLER_68_1283 ();
 sg13g2_decap_8 FILLER_68_1290 ();
 sg13g2_decap_8 FILLER_68_1297 ();
 sg13g2_decap_8 FILLER_68_1304 ();
 sg13g2_decap_8 FILLER_68_1311 ();
 sg13g2_decap_8 FILLER_68_1318 ();
 sg13g2_fill_1 FILLER_68_1325 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_4 FILLER_69_28 ();
 sg13g2_fill_1 FILLER_69_36 ();
 sg13g2_decap_8 FILLER_69_53 ();
 sg13g2_decap_4 FILLER_69_60 ();
 sg13g2_decap_4 FILLER_69_69 ();
 sg13g2_fill_2 FILLER_69_73 ();
 sg13g2_decap_8 FILLER_69_79 ();
 sg13g2_fill_2 FILLER_69_86 ();
 sg13g2_fill_1 FILLER_69_88 ();
 sg13g2_decap_4 FILLER_69_93 ();
 sg13g2_fill_1 FILLER_69_97 ();
 sg13g2_decap_8 FILLER_69_103 ();
 sg13g2_decap_8 FILLER_69_110 ();
 sg13g2_decap_8 FILLER_69_117 ();
 sg13g2_decap_8 FILLER_69_124 ();
 sg13g2_decap_4 FILLER_69_131 ();
 sg13g2_fill_2 FILLER_69_135 ();
 sg13g2_decap_4 FILLER_69_152 ();
 sg13g2_fill_2 FILLER_69_156 ();
 sg13g2_decap_4 FILLER_69_173 ();
 sg13g2_fill_1 FILLER_69_177 ();
 sg13g2_decap_4 FILLER_69_183 ();
 sg13g2_fill_2 FILLER_69_187 ();
 sg13g2_decap_8 FILLER_69_200 ();
 sg13g2_decap_8 FILLER_69_207 ();
 sg13g2_decap_8 FILLER_69_219 ();
 sg13g2_fill_1 FILLER_69_226 ();
 sg13g2_fill_1 FILLER_69_232 ();
 sg13g2_decap_8 FILLER_69_268 ();
 sg13g2_fill_2 FILLER_69_275 ();
 sg13g2_fill_1 FILLER_69_277 ();
 sg13g2_decap_8 FILLER_69_287 ();
 sg13g2_decap_4 FILLER_69_294 ();
 sg13g2_fill_2 FILLER_69_298 ();
 sg13g2_decap_8 FILLER_69_305 ();
 sg13g2_decap_8 FILLER_69_342 ();
 sg13g2_decap_8 FILLER_69_349 ();
 sg13g2_decap_8 FILLER_69_356 ();
 sg13g2_fill_2 FILLER_69_363 ();
 sg13g2_decap_8 FILLER_69_396 ();
 sg13g2_decap_8 FILLER_69_403 ();
 sg13g2_decap_4 FILLER_69_410 ();
 sg13g2_fill_1 FILLER_69_414 ();
 sg13g2_decap_8 FILLER_69_430 ();
 sg13g2_fill_2 FILLER_69_437 ();
 sg13g2_decap_8 FILLER_69_443 ();
 sg13g2_decap_8 FILLER_69_458 ();
 sg13g2_decap_8 FILLER_69_465 ();
 sg13g2_decap_8 FILLER_69_472 ();
 sg13g2_decap_8 FILLER_69_479 ();
 sg13g2_decap_8 FILLER_69_486 ();
 sg13g2_decap_8 FILLER_69_493 ();
 sg13g2_decap_8 FILLER_69_500 ();
 sg13g2_decap_4 FILLER_69_507 ();
 sg13g2_fill_1 FILLER_69_511 ();
 sg13g2_decap_4 FILLER_69_516 ();
 sg13g2_decap_4 FILLER_69_524 ();
 sg13g2_decap_8 FILLER_69_554 ();
 sg13g2_decap_8 FILLER_69_561 ();
 sg13g2_fill_2 FILLER_69_568 ();
 sg13g2_decap_8 FILLER_69_582 ();
 sg13g2_fill_1 FILLER_69_589 ();
 sg13g2_decap_8 FILLER_69_599 ();
 sg13g2_decap_8 FILLER_69_606 ();
 sg13g2_decap_8 FILLER_69_613 ();
 sg13g2_decap_8 FILLER_69_620 ();
 sg13g2_decap_8 FILLER_69_627 ();
 sg13g2_decap_8 FILLER_69_634 ();
 sg13g2_decap_8 FILLER_69_645 ();
 sg13g2_fill_2 FILLER_69_652 ();
 sg13g2_decap_8 FILLER_69_680 ();
 sg13g2_decap_8 FILLER_69_687 ();
 sg13g2_decap_8 FILLER_69_694 ();
 sg13g2_decap_8 FILLER_69_701 ();
 sg13g2_decap_8 FILLER_69_708 ();
 sg13g2_decap_8 FILLER_69_715 ();
 sg13g2_decap_8 FILLER_69_722 ();
 sg13g2_decap_8 FILLER_69_729 ();
 sg13g2_fill_1 FILLER_69_736 ();
 sg13g2_decap_8 FILLER_69_741 ();
 sg13g2_decap_8 FILLER_69_748 ();
 sg13g2_decap_4 FILLER_69_755 ();
 sg13g2_fill_1 FILLER_69_759 ();
 sg13g2_decap_8 FILLER_69_763 ();
 sg13g2_decap_8 FILLER_69_770 ();
 sg13g2_fill_2 FILLER_69_777 ();
 sg13g2_fill_1 FILLER_69_779 ();
 sg13g2_decap_8 FILLER_69_784 ();
 sg13g2_decap_8 FILLER_69_791 ();
 sg13g2_decap_8 FILLER_69_798 ();
 sg13g2_decap_4 FILLER_69_805 ();
 sg13g2_fill_2 FILLER_69_809 ();
 sg13g2_decap_8 FILLER_69_815 ();
 sg13g2_decap_8 FILLER_69_822 ();
 sg13g2_decap_8 FILLER_69_829 ();
 sg13g2_decap_8 FILLER_69_836 ();
 sg13g2_decap_8 FILLER_69_843 ();
 sg13g2_decap_8 FILLER_69_850 ();
 sg13g2_decap_8 FILLER_69_857 ();
 sg13g2_decap_8 FILLER_69_864 ();
 sg13g2_decap_8 FILLER_69_871 ();
 sg13g2_decap_4 FILLER_69_878 ();
 sg13g2_fill_1 FILLER_69_882 ();
 sg13g2_decap_8 FILLER_69_888 ();
 sg13g2_fill_2 FILLER_69_895 ();
 sg13g2_fill_1 FILLER_69_909 ();
 sg13g2_fill_2 FILLER_69_915 ();
 sg13g2_fill_1 FILLER_69_917 ();
 sg13g2_fill_1 FILLER_69_937 ();
 sg13g2_decap_8 FILLER_69_942 ();
 sg13g2_decap_8 FILLER_69_949 ();
 sg13g2_decap_8 FILLER_69_956 ();
 sg13g2_decap_8 FILLER_69_963 ();
 sg13g2_fill_1 FILLER_69_970 ();
 sg13g2_decap_4 FILLER_69_976 ();
 sg13g2_decap_8 FILLER_69_984 ();
 sg13g2_decap_8 FILLER_69_991 ();
 sg13g2_decap_8 FILLER_69_1003 ();
 sg13g2_decap_4 FILLER_69_1010 ();
 sg13g2_fill_1 FILLER_69_1014 ();
 sg13g2_decap_8 FILLER_69_1019 ();
 sg13g2_decap_8 FILLER_69_1026 ();
 sg13g2_decap_8 FILLER_69_1033 ();
 sg13g2_fill_2 FILLER_69_1040 ();
 sg13g2_fill_1 FILLER_69_1042 ();
 sg13g2_decap_8 FILLER_69_1049 ();
 sg13g2_decap_8 FILLER_69_1056 ();
 sg13g2_decap_8 FILLER_69_1063 ();
 sg13g2_decap_4 FILLER_69_1070 ();
 sg13g2_fill_2 FILLER_69_1074 ();
 sg13g2_decap_4 FILLER_69_1081 ();
 sg13g2_fill_2 FILLER_69_1085 ();
 sg13g2_decap_8 FILLER_69_1093 ();
 sg13g2_decap_8 FILLER_69_1100 ();
 sg13g2_decap_4 FILLER_69_1107 ();
 sg13g2_fill_2 FILLER_69_1111 ();
 sg13g2_decap_8 FILLER_69_1121 ();
 sg13g2_decap_4 FILLER_69_1128 ();
 sg13g2_fill_1 FILLER_69_1132 ();
 sg13g2_decap_8 FILLER_69_1136 ();
 sg13g2_decap_8 FILLER_69_1143 ();
 sg13g2_decap_8 FILLER_69_1150 ();
 sg13g2_decap_4 FILLER_69_1157 ();
 sg13g2_fill_1 FILLER_69_1161 ();
 sg13g2_decap_8 FILLER_69_1167 ();
 sg13g2_decap_4 FILLER_69_1174 ();
 sg13g2_fill_2 FILLER_69_1178 ();
 sg13g2_decap_8 FILLER_69_1184 ();
 sg13g2_decap_4 FILLER_69_1191 ();
 sg13g2_fill_2 FILLER_69_1209 ();
 sg13g2_fill_1 FILLER_69_1211 ();
 sg13g2_fill_2 FILLER_69_1217 ();
 sg13g2_fill_1 FILLER_69_1219 ();
 sg13g2_decap_4 FILLER_69_1224 ();
 sg13g2_fill_2 FILLER_69_1228 ();
 sg13g2_decap_8 FILLER_69_1248 ();
 sg13g2_fill_1 FILLER_69_1255 ();
 sg13g2_decap_4 FILLER_69_1266 ();
 sg13g2_fill_1 FILLER_69_1270 ();
 sg13g2_decap_8 FILLER_69_1276 ();
 sg13g2_decap_8 FILLER_69_1283 ();
 sg13g2_decap_8 FILLER_69_1290 ();
 sg13g2_decap_8 FILLER_69_1297 ();
 sg13g2_decap_8 FILLER_69_1304 ();
 sg13g2_decap_8 FILLER_69_1311 ();
 sg13g2_decap_8 FILLER_69_1318 ();
 sg13g2_fill_1 FILLER_69_1325 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_fill_2 FILLER_70_21 ();
 sg13g2_fill_1 FILLER_70_23 ();
 sg13g2_decap_4 FILLER_70_50 ();
 sg13g2_fill_1 FILLER_70_54 ();
 sg13g2_fill_1 FILLER_70_60 ();
 sg13g2_decap_8 FILLER_70_71 ();
 sg13g2_decap_8 FILLER_70_78 ();
 sg13g2_fill_1 FILLER_70_85 ();
 sg13g2_decap_4 FILLER_70_95 ();
 sg13g2_decap_8 FILLER_70_103 ();
 sg13g2_decap_8 FILLER_70_110 ();
 sg13g2_fill_2 FILLER_70_117 ();
 sg13g2_fill_1 FILLER_70_119 ();
 sg13g2_fill_2 FILLER_70_123 ();
 sg13g2_fill_1 FILLER_70_125 ();
 sg13g2_decap_8 FILLER_70_131 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_fill_1 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_211 ();
 sg13g2_decap_8 FILLER_70_218 ();
 sg13g2_fill_2 FILLER_70_225 ();
 sg13g2_fill_1 FILLER_70_227 ();
 sg13g2_fill_1 FILLER_70_237 ();
 sg13g2_fill_2 FILLER_70_247 ();
 sg13g2_fill_1 FILLER_70_249 ();
 sg13g2_decap_4 FILLER_70_255 ();
 sg13g2_fill_2 FILLER_70_259 ();
 sg13g2_decap_8 FILLER_70_268 ();
 sg13g2_decap_8 FILLER_70_275 ();
 sg13g2_decap_8 FILLER_70_282 ();
 sg13g2_decap_8 FILLER_70_289 ();
 sg13g2_decap_4 FILLER_70_296 ();
 sg13g2_fill_1 FILLER_70_300 ();
 sg13g2_decap_4 FILLER_70_306 ();
 sg13g2_fill_1 FILLER_70_310 ();
 sg13g2_fill_1 FILLER_70_320 ();
 sg13g2_fill_1 FILLER_70_326 ();
 sg13g2_decap_8 FILLER_70_332 ();
 sg13g2_decap_8 FILLER_70_339 ();
 sg13g2_decap_8 FILLER_70_346 ();
 sg13g2_decap_8 FILLER_70_353 ();
 sg13g2_fill_1 FILLER_70_369 ();
 sg13g2_decap_8 FILLER_70_379 ();
 sg13g2_decap_8 FILLER_70_386 ();
 sg13g2_decap_8 FILLER_70_393 ();
 sg13g2_decap_8 FILLER_70_400 ();
 sg13g2_fill_1 FILLER_70_407 ();
 sg13g2_fill_2 FILLER_70_413 ();
 sg13g2_fill_1 FILLER_70_415 ();
 sg13g2_decap_8 FILLER_70_420 ();
 sg13g2_decap_8 FILLER_70_427 ();
 sg13g2_decap_8 FILLER_70_434 ();
 sg13g2_decap_8 FILLER_70_441 ();
 sg13g2_decap_8 FILLER_70_448 ();
 sg13g2_decap_8 FILLER_70_455 ();
 sg13g2_decap_8 FILLER_70_462 ();
 sg13g2_decap_8 FILLER_70_469 ();
 sg13g2_decap_8 FILLER_70_476 ();
 sg13g2_decap_8 FILLER_70_483 ();
 sg13g2_decap_4 FILLER_70_490 ();
 sg13g2_fill_1 FILLER_70_494 ();
 sg13g2_fill_1 FILLER_70_499 ();
 sg13g2_decap_8 FILLER_70_531 ();
 sg13g2_decap_8 FILLER_70_538 ();
 sg13g2_decap_8 FILLER_70_545 ();
 sg13g2_decap_4 FILLER_70_552 ();
 sg13g2_fill_2 FILLER_70_556 ();
 sg13g2_fill_2 FILLER_70_579 ();
 sg13g2_fill_1 FILLER_70_581 ();
 sg13g2_decap_8 FILLER_70_608 ();
 sg13g2_decap_8 FILLER_70_615 ();
 sg13g2_decap_8 FILLER_70_622 ();
 sg13g2_decap_8 FILLER_70_629 ();
 sg13g2_decap_8 FILLER_70_636 ();
 sg13g2_decap_8 FILLER_70_643 ();
 sg13g2_decap_8 FILLER_70_683 ();
 sg13g2_decap_8 FILLER_70_690 ();
 sg13g2_decap_4 FILLER_70_697 ();
 sg13g2_fill_2 FILLER_70_701 ();
 sg13g2_decap_4 FILLER_70_708 ();
 sg13g2_fill_1 FILLER_70_712 ();
 sg13g2_decap_8 FILLER_70_717 ();
 sg13g2_decap_8 FILLER_70_724 ();
 sg13g2_decap_8 FILLER_70_731 ();
 sg13g2_fill_2 FILLER_70_738 ();
 sg13g2_fill_1 FILLER_70_740 ();
 sg13g2_decap_4 FILLER_70_746 ();
 sg13g2_fill_1 FILLER_70_750 ();
 sg13g2_decap_4 FILLER_70_756 ();
 sg13g2_decap_4 FILLER_70_769 ();
 sg13g2_fill_1 FILLER_70_773 ();
 sg13g2_decap_8 FILLER_70_778 ();
 sg13g2_decap_8 FILLER_70_785 ();
 sg13g2_decap_8 FILLER_70_792 ();
 sg13g2_decap_8 FILLER_70_799 ();
 sg13g2_decap_4 FILLER_70_806 ();
 sg13g2_fill_1 FILLER_70_810 ();
 sg13g2_decap_8 FILLER_70_815 ();
 sg13g2_decap_8 FILLER_70_822 ();
 sg13g2_decap_8 FILLER_70_829 ();
 sg13g2_fill_1 FILLER_70_836 ();
 sg13g2_decap_8 FILLER_70_841 ();
 sg13g2_decap_8 FILLER_70_848 ();
 sg13g2_decap_8 FILLER_70_855 ();
 sg13g2_decap_8 FILLER_70_862 ();
 sg13g2_decap_8 FILLER_70_869 ();
 sg13g2_decap_8 FILLER_70_876 ();
 sg13g2_decap_8 FILLER_70_883 ();
 sg13g2_fill_2 FILLER_70_890 ();
 sg13g2_fill_1 FILLER_70_892 ();
 sg13g2_decap_8 FILLER_70_903 ();
 sg13g2_decap_8 FILLER_70_910 ();
 sg13g2_fill_2 FILLER_70_928 ();
 sg13g2_decap_4 FILLER_70_939 ();
 sg13g2_fill_2 FILLER_70_943 ();
 sg13g2_decap_8 FILLER_70_962 ();
 sg13g2_fill_2 FILLER_70_969 ();
 sg13g2_decap_8 FILLER_70_977 ();
 sg13g2_decap_8 FILLER_70_984 ();
 sg13g2_decap_8 FILLER_70_991 ();
 sg13g2_decap_8 FILLER_70_998 ();
 sg13g2_decap_8 FILLER_70_1005 ();
 sg13g2_decap_8 FILLER_70_1017 ();
 sg13g2_decap_8 FILLER_70_1024 ();
 sg13g2_decap_8 FILLER_70_1036 ();
 sg13g2_decap_8 FILLER_70_1043 ();
 sg13g2_decap_8 FILLER_70_1050 ();
 sg13g2_fill_1 FILLER_70_1057 ();
 sg13g2_fill_2 FILLER_70_1073 ();
 sg13g2_fill_1 FILLER_70_1075 ();
 sg13g2_decap_8 FILLER_70_1080 ();
 sg13g2_decap_4 FILLER_70_1087 ();
 sg13g2_fill_2 FILLER_70_1091 ();
 sg13g2_decap_8 FILLER_70_1097 ();
 sg13g2_fill_2 FILLER_70_1104 ();
 sg13g2_fill_1 FILLER_70_1106 ();
 sg13g2_decap_8 FILLER_70_1110 ();
 sg13g2_decap_8 FILLER_70_1122 ();
 sg13g2_fill_1 FILLER_70_1129 ();
 sg13g2_fill_2 FILLER_70_1140 ();
 sg13g2_decap_8 FILLER_70_1147 ();
 sg13g2_decap_8 FILLER_70_1154 ();
 sg13g2_decap_4 FILLER_70_1161 ();
 sg13g2_fill_1 FILLER_70_1165 ();
 sg13g2_decap_4 FILLER_70_1169 ();
 sg13g2_fill_2 FILLER_70_1173 ();
 sg13g2_decap_4 FILLER_70_1188 ();
 sg13g2_fill_1 FILLER_70_1192 ();
 sg13g2_fill_2 FILLER_70_1207 ();
 sg13g2_decap_4 FILLER_70_1213 ();
 sg13g2_decap_8 FILLER_70_1222 ();
 sg13g2_decap_8 FILLER_70_1229 ();
 sg13g2_decap_8 FILLER_70_1236 ();
 sg13g2_fill_1 FILLER_70_1243 ();
 sg13g2_fill_2 FILLER_70_1248 ();
 sg13g2_fill_1 FILLER_70_1250 ();
 sg13g2_fill_2 FILLER_70_1256 ();
 sg13g2_decap_8 FILLER_70_1266 ();
 sg13g2_fill_1 FILLER_70_1273 ();
 sg13g2_decap_8 FILLER_70_1295 ();
 sg13g2_decap_8 FILLER_70_1302 ();
 sg13g2_decap_8 FILLER_70_1309 ();
 sg13g2_decap_8 FILLER_70_1316 ();
 sg13g2_fill_2 FILLER_70_1323 ();
 sg13g2_fill_1 FILLER_70_1325 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_fill_1 FILLER_71_35 ();
 sg13g2_decap_4 FILLER_71_40 ();
 sg13g2_fill_1 FILLER_71_44 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_fill_2 FILLER_71_56 ();
 sg13g2_decap_4 FILLER_71_68 ();
 sg13g2_fill_2 FILLER_71_72 ();
 sg13g2_fill_2 FILLER_71_83 ();
 sg13g2_fill_1 FILLER_71_85 ();
 sg13g2_decap_4 FILLER_71_96 ();
 sg13g2_fill_1 FILLER_71_100 ();
 sg13g2_decap_8 FILLER_71_110 ();
 sg13g2_decap_4 FILLER_71_122 ();
 sg13g2_fill_1 FILLER_71_126 ();
 sg13g2_fill_2 FILLER_71_131 ();
 sg13g2_fill_1 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_149 ();
 sg13g2_decap_8 FILLER_71_166 ();
 sg13g2_decap_8 FILLER_71_173 ();
 sg13g2_decap_8 FILLER_71_180 ();
 sg13g2_decap_8 FILLER_71_187 ();
 sg13g2_decap_8 FILLER_71_194 ();
 sg13g2_decap_8 FILLER_71_201 ();
 sg13g2_decap_4 FILLER_71_208 ();
 sg13g2_fill_2 FILLER_71_212 ();
 sg13g2_decap_8 FILLER_71_219 ();
 sg13g2_decap_8 FILLER_71_226 ();
 sg13g2_decap_8 FILLER_71_233 ();
 sg13g2_decap_8 FILLER_71_240 ();
 sg13g2_decap_8 FILLER_71_247 ();
 sg13g2_decap_8 FILLER_71_254 ();
 sg13g2_decap_8 FILLER_71_267 ();
 sg13g2_decap_8 FILLER_71_305 ();
 sg13g2_decap_8 FILLER_71_312 ();
 sg13g2_decap_8 FILLER_71_319 ();
 sg13g2_decap_8 FILLER_71_330 ();
 sg13g2_decap_8 FILLER_71_337 ();
 sg13g2_decap_8 FILLER_71_344 ();
 sg13g2_decap_8 FILLER_71_351 ();
 sg13g2_fill_2 FILLER_71_358 ();
 sg13g2_decap_8 FILLER_71_365 ();
 sg13g2_decap_8 FILLER_71_372 ();
 sg13g2_decap_8 FILLER_71_379 ();
 sg13g2_decap_8 FILLER_71_386 ();
 sg13g2_fill_1 FILLER_71_393 ();
 sg13g2_decap_8 FILLER_71_400 ();
 sg13g2_decap_4 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_71_420 ();
 sg13g2_fill_2 FILLER_71_427 ();
 sg13g2_fill_1 FILLER_71_429 ();
 sg13g2_decap_8 FILLER_71_435 ();
 sg13g2_decap_8 FILLER_71_442 ();
 sg13g2_fill_2 FILLER_71_449 ();
 sg13g2_fill_1 FILLER_71_451 ();
 sg13g2_decap_8 FILLER_71_478 ();
 sg13g2_decap_4 FILLER_71_485 ();
 sg13g2_fill_1 FILLER_71_489 ();
 sg13g2_fill_2 FILLER_71_521 ();
 sg13g2_decap_8 FILLER_71_544 ();
 sg13g2_decap_8 FILLER_71_551 ();
 sg13g2_decap_8 FILLER_71_558 ();
 sg13g2_fill_1 FILLER_71_565 ();
 sg13g2_decap_8 FILLER_71_587 ();
 sg13g2_decap_8 FILLER_71_599 ();
 sg13g2_decap_8 FILLER_71_606 ();
 sg13g2_decap_8 FILLER_71_613 ();
 sg13g2_decap_8 FILLER_71_620 ();
 sg13g2_decap_4 FILLER_71_627 ();
 sg13g2_decap_8 FILLER_71_635 ();
 sg13g2_decap_8 FILLER_71_642 ();
 sg13g2_decap_8 FILLER_71_649 ();
 sg13g2_decap_4 FILLER_71_656 ();
 sg13g2_fill_2 FILLER_71_660 ();
 sg13g2_decap_8 FILLER_71_666 ();
 sg13g2_decap_8 FILLER_71_676 ();
 sg13g2_decap_8 FILLER_71_688 ();
 sg13g2_decap_8 FILLER_71_695 ();
 sg13g2_fill_1 FILLER_71_702 ();
 sg13g2_decap_8 FILLER_71_712 ();
 sg13g2_decap_8 FILLER_71_719 ();
 sg13g2_decap_8 FILLER_71_726 ();
 sg13g2_decap_8 FILLER_71_733 ();
 sg13g2_decap_8 FILLER_71_740 ();
 sg13g2_fill_2 FILLER_71_760 ();
 sg13g2_fill_2 FILLER_71_806 ();
 sg13g2_decap_8 FILLER_71_812 ();
 sg13g2_fill_1 FILLER_71_819 ();
 sg13g2_fill_1 FILLER_71_826 ();
 sg13g2_decap_4 FILLER_71_842 ();
 sg13g2_decap_8 FILLER_71_851 ();
 sg13g2_decap_8 FILLER_71_858 ();
 sg13g2_decap_8 FILLER_71_865 ();
 sg13g2_decap_4 FILLER_71_872 ();
 sg13g2_fill_1 FILLER_71_876 ();
 sg13g2_decap_8 FILLER_71_898 ();
 sg13g2_fill_2 FILLER_71_905 ();
 sg13g2_fill_1 FILLER_71_907 ();
 sg13g2_fill_2 FILLER_71_929 ();
 sg13g2_decap_4 FILLER_71_941 ();
 sg13g2_decap_4 FILLER_71_961 ();
 sg13g2_fill_2 FILLER_71_965 ();
 sg13g2_fill_1 FILLER_71_975 ();
 sg13g2_decap_8 FILLER_71_981 ();
 sg13g2_fill_2 FILLER_71_1003 ();
 sg13g2_decap_8 FILLER_71_1024 ();
 sg13g2_decap_8 FILLER_71_1031 ();
 sg13g2_fill_1 FILLER_71_1038 ();
 sg13g2_fill_1 FILLER_71_1044 ();
 sg13g2_decap_4 FILLER_71_1058 ();
 sg13g2_fill_1 FILLER_71_1075 ();
 sg13g2_decap_8 FILLER_71_1085 ();
 sg13g2_decap_8 FILLER_71_1092 ();
 sg13g2_decap_8 FILLER_71_1099 ();
 sg13g2_decap_8 FILLER_71_1106 ();
 sg13g2_fill_2 FILLER_71_1113 ();
 sg13g2_fill_2 FILLER_71_1141 ();
 sg13g2_decap_8 FILLER_71_1156 ();
 sg13g2_decap_4 FILLER_71_1163 ();
 sg13g2_decap_8 FILLER_71_1172 ();
 sg13g2_fill_2 FILLER_71_1179 ();
 sg13g2_fill_1 FILLER_71_1186 ();
 sg13g2_fill_2 FILLER_71_1197 ();
 sg13g2_fill_2 FILLER_71_1214 ();
 sg13g2_fill_1 FILLER_71_1216 ();
 sg13g2_decap_4 FILLER_71_1222 ();
 sg13g2_fill_1 FILLER_71_1226 ();
 sg13g2_decap_8 FILLER_71_1231 ();
 sg13g2_decap_8 FILLER_71_1238 ();
 sg13g2_decap_8 FILLER_71_1245 ();
 sg13g2_fill_2 FILLER_71_1261 ();
 sg13g2_fill_1 FILLER_71_1263 ();
 sg13g2_decap_8 FILLER_71_1272 ();
 sg13g2_decap_8 FILLER_71_1279 ();
 sg13g2_decap_8 FILLER_71_1286 ();
 sg13g2_decap_8 FILLER_71_1293 ();
 sg13g2_decap_8 FILLER_71_1300 ();
 sg13g2_decap_8 FILLER_71_1307 ();
 sg13g2_decap_8 FILLER_71_1314 ();
 sg13g2_decap_4 FILLER_71_1321 ();
 sg13g2_fill_1 FILLER_71_1325 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_4 FILLER_72_28 ();
 sg13g2_fill_2 FILLER_72_32 ();
 sg13g2_fill_2 FILLER_72_46 ();
 sg13g2_decap_8 FILLER_72_53 ();
 sg13g2_fill_1 FILLER_72_60 ();
 sg13g2_decap_8 FILLER_72_80 ();
 sg13g2_decap_4 FILLER_72_87 ();
 sg13g2_decap_4 FILLER_72_96 ();
 sg13g2_fill_2 FILLER_72_100 ();
 sg13g2_decap_8 FILLER_72_107 ();
 sg13g2_decap_8 FILLER_72_114 ();
 sg13g2_decap_8 FILLER_72_121 ();
 sg13g2_decap_8 FILLER_72_132 ();
 sg13g2_decap_8 FILLER_72_139 ();
 sg13g2_fill_2 FILLER_72_149 ();
 sg13g2_decap_8 FILLER_72_164 ();
 sg13g2_decap_8 FILLER_72_171 ();
 sg13g2_fill_2 FILLER_72_178 ();
 sg13g2_fill_1 FILLER_72_180 ();
 sg13g2_decap_8 FILLER_72_185 ();
 sg13g2_fill_2 FILLER_72_192 ();
 sg13g2_fill_1 FILLER_72_194 ();
 sg13g2_decap_8 FILLER_72_214 ();
 sg13g2_decap_8 FILLER_72_221 ();
 sg13g2_decap_8 FILLER_72_228 ();
 sg13g2_decap_8 FILLER_72_235 ();
 sg13g2_decap_8 FILLER_72_242 ();
 sg13g2_decap_8 FILLER_72_249 ();
 sg13g2_decap_8 FILLER_72_256 ();
 sg13g2_decap_4 FILLER_72_263 ();
 sg13g2_fill_2 FILLER_72_267 ();
 sg13g2_decap_8 FILLER_72_273 ();
 sg13g2_decap_4 FILLER_72_280 ();
 sg13g2_fill_2 FILLER_72_284 ();
 sg13g2_decap_8 FILLER_72_290 ();
 sg13g2_decap_8 FILLER_72_297 ();
 sg13g2_decap_4 FILLER_72_304 ();
 sg13g2_decap_8 FILLER_72_313 ();
 sg13g2_decap_8 FILLER_72_320 ();
 sg13g2_decap_8 FILLER_72_327 ();
 sg13g2_decap_8 FILLER_72_334 ();
 sg13g2_decap_8 FILLER_72_341 ();
 sg13g2_decap_8 FILLER_72_348 ();
 sg13g2_decap_8 FILLER_72_386 ();
 sg13g2_fill_1 FILLER_72_393 ();
 sg13g2_fill_2 FILLER_72_399 ();
 sg13g2_fill_2 FILLER_72_410 ();
 sg13g2_decap_8 FILLER_72_423 ();
 sg13g2_decap_4 FILLER_72_430 ();
 sg13g2_fill_2 FILLER_72_434 ();
 sg13g2_decap_8 FILLER_72_440 ();
 sg13g2_decap_8 FILLER_72_447 ();
 sg13g2_decap_8 FILLER_72_454 ();
 sg13g2_decap_8 FILLER_72_465 ();
 sg13g2_decap_8 FILLER_72_472 ();
 sg13g2_decap_8 FILLER_72_479 ();
 sg13g2_decap_8 FILLER_72_486 ();
 sg13g2_decap_8 FILLER_72_493 ();
 sg13g2_decap_8 FILLER_72_500 ();
 sg13g2_decap_8 FILLER_72_538 ();
 sg13g2_decap_8 FILLER_72_545 ();
 sg13g2_decap_8 FILLER_72_552 ();
 sg13g2_decap_8 FILLER_72_559 ();
 sg13g2_decap_8 FILLER_72_566 ();
 sg13g2_decap_8 FILLER_72_573 ();
 sg13g2_decap_8 FILLER_72_580 ();
 sg13g2_fill_1 FILLER_72_587 ();
 sg13g2_fill_1 FILLER_72_596 ();
 sg13g2_decap_8 FILLER_72_639 ();
 sg13g2_fill_1 FILLER_72_646 ();
 sg13g2_decap_8 FILLER_72_655 ();
 sg13g2_fill_2 FILLER_72_662 ();
 sg13g2_fill_1 FILLER_72_664 ();
 sg13g2_decap_4 FILLER_72_669 ();
 sg13g2_decap_8 FILLER_72_677 ();
 sg13g2_decap_8 FILLER_72_684 ();
 sg13g2_decap_4 FILLER_72_691 ();
 sg13g2_fill_2 FILLER_72_695 ();
 sg13g2_decap_8 FILLER_72_728 ();
 sg13g2_decap_8 FILLER_72_735 ();
 sg13g2_fill_2 FILLER_72_742 ();
 sg13g2_decap_4 FILLER_72_761 ();
 sg13g2_fill_1 FILLER_72_765 ();
 sg13g2_fill_1 FILLER_72_778 ();
 sg13g2_fill_2 FILLER_72_787 ();
 sg13g2_fill_1 FILLER_72_801 ();
 sg13g2_decap_8 FILLER_72_807 ();
 sg13g2_decap_8 FILLER_72_814 ();
 sg13g2_decap_8 FILLER_72_821 ();
 sg13g2_decap_8 FILLER_72_828 ();
 sg13g2_decap_8 FILLER_72_835 ();
 sg13g2_decap_8 FILLER_72_842 ();
 sg13g2_decap_8 FILLER_72_849 ();
 sg13g2_decap_8 FILLER_72_856 ();
 sg13g2_decap_8 FILLER_72_863 ();
 sg13g2_decap_4 FILLER_72_870 ();
 sg13g2_decap_8 FILLER_72_888 ();
 sg13g2_decap_8 FILLER_72_895 ();
 sg13g2_decap_4 FILLER_72_902 ();
 sg13g2_fill_1 FILLER_72_906 ();
 sg13g2_fill_1 FILLER_72_912 ();
 sg13g2_decap_8 FILLER_72_922 ();
 sg13g2_fill_2 FILLER_72_929 ();
 sg13g2_fill_1 FILLER_72_931 ();
 sg13g2_decap_8 FILLER_72_946 ();
 sg13g2_decap_4 FILLER_72_953 ();
 sg13g2_fill_1 FILLER_72_957 ();
 sg13g2_fill_1 FILLER_72_964 ();
 sg13g2_decap_4 FILLER_72_972 ();
 sg13g2_fill_2 FILLER_72_976 ();
 sg13g2_decap_4 FILLER_72_982 ();
 sg13g2_fill_1 FILLER_72_986 ();
 sg13g2_fill_2 FILLER_72_1005 ();
 sg13g2_fill_1 FILLER_72_1007 ();
 sg13g2_fill_1 FILLER_72_1013 ();
 sg13g2_decap_8 FILLER_72_1019 ();
 sg13g2_decap_8 FILLER_72_1026 ();
 sg13g2_fill_2 FILLER_72_1033 ();
 sg13g2_decap_8 FILLER_72_1054 ();
 sg13g2_fill_1 FILLER_72_1061 ();
 sg13g2_decap_8 FILLER_72_1077 ();
 sg13g2_fill_2 FILLER_72_1084 ();
 sg13g2_fill_1 FILLER_72_1086 ();
 sg13g2_decap_8 FILLER_72_1091 ();
 sg13g2_decap_8 FILLER_72_1098 ();
 sg13g2_decap_4 FILLER_72_1105 ();
 sg13g2_decap_8 FILLER_72_1114 ();
 sg13g2_decap_8 FILLER_72_1121 ();
 sg13g2_fill_2 FILLER_72_1128 ();
 sg13g2_fill_1 FILLER_72_1130 ();
 sg13g2_fill_1 FILLER_72_1136 ();
 sg13g2_decap_8 FILLER_72_1141 ();
 sg13g2_decap_4 FILLER_72_1148 ();
 sg13g2_fill_2 FILLER_72_1152 ();
 sg13g2_decap_8 FILLER_72_1159 ();
 sg13g2_fill_1 FILLER_72_1166 ();
 sg13g2_decap_8 FILLER_72_1173 ();
 sg13g2_decap_4 FILLER_72_1180 ();
 sg13g2_fill_1 FILLER_72_1184 ();
 sg13g2_decap_4 FILLER_72_1189 ();
 sg13g2_fill_1 FILLER_72_1193 ();
 sg13g2_decap_4 FILLER_72_1204 ();
 sg13g2_fill_1 FILLER_72_1208 ();
 sg13g2_decap_4 FILLER_72_1214 ();
 sg13g2_fill_1 FILLER_72_1218 ();
 sg13g2_decap_8 FILLER_72_1223 ();
 sg13g2_decap_4 FILLER_72_1230 ();
 sg13g2_decap_4 FILLER_72_1238 ();
 sg13g2_fill_1 FILLER_72_1242 ();
 sg13g2_decap_8 FILLER_72_1263 ();
 sg13g2_decap_8 FILLER_72_1270 ();
 sg13g2_decap_8 FILLER_72_1277 ();
 sg13g2_decap_8 FILLER_72_1284 ();
 sg13g2_decap_8 FILLER_72_1291 ();
 sg13g2_decap_8 FILLER_72_1298 ();
 sg13g2_decap_8 FILLER_72_1305 ();
 sg13g2_decap_8 FILLER_72_1312 ();
 sg13g2_decap_8 FILLER_72_1319 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_fill_1 FILLER_73_28 ();
 sg13g2_fill_1 FILLER_73_37 ();
 sg13g2_fill_2 FILLER_73_51 ();
 sg13g2_fill_1 FILLER_73_66 ();
 sg13g2_fill_2 FILLER_73_82 ();
 sg13g2_fill_1 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_100 ();
 sg13g2_decap_8 FILLER_73_107 ();
 sg13g2_decap_4 FILLER_73_114 ();
 sg13g2_fill_1 FILLER_73_128 ();
 sg13g2_decap_8 FILLER_73_135 ();
 sg13g2_decap_8 FILLER_73_153 ();
 sg13g2_fill_2 FILLER_73_163 ();
 sg13g2_decap_8 FILLER_73_186 ();
 sg13g2_decap_8 FILLER_73_193 ();
 sg13g2_fill_2 FILLER_73_222 ();
 sg13g2_fill_1 FILLER_73_224 ();
 sg13g2_decap_8 FILLER_73_229 ();
 sg13g2_decap_8 FILLER_73_236 ();
 sg13g2_fill_2 FILLER_73_243 ();
 sg13g2_decap_8 FILLER_73_249 ();
 sg13g2_fill_1 FILLER_73_256 ();
 sg13g2_decap_8 FILLER_73_261 ();
 sg13g2_fill_1 FILLER_73_268 ();
 sg13g2_decap_8 FILLER_73_273 ();
 sg13g2_decap_8 FILLER_73_280 ();
 sg13g2_decap_8 FILLER_73_287 ();
 sg13g2_decap_4 FILLER_73_299 ();
 sg13g2_decap_8 FILLER_73_342 ();
 sg13g2_decap_8 FILLER_73_349 ();
 sg13g2_decap_8 FILLER_73_356 ();
 sg13g2_fill_2 FILLER_73_363 ();
 sg13g2_decap_8 FILLER_73_369 ();
 sg13g2_decap_8 FILLER_73_376 ();
 sg13g2_decap_8 FILLER_73_383 ();
 sg13g2_decap_4 FILLER_73_390 ();
 sg13g2_fill_2 FILLER_73_394 ();
 sg13g2_decap_4 FILLER_73_406 ();
 sg13g2_fill_1 FILLER_73_410 ();
 sg13g2_decap_8 FILLER_73_417 ();
 sg13g2_fill_1 FILLER_73_424 ();
 sg13g2_decap_8 FILLER_73_460 ();
 sg13g2_decap_8 FILLER_73_467 ();
 sg13g2_decap_8 FILLER_73_474 ();
 sg13g2_decap_4 FILLER_73_481 ();
 sg13g2_fill_1 FILLER_73_485 ();
 sg13g2_decap_8 FILLER_73_490 ();
 sg13g2_decap_8 FILLER_73_497 ();
 sg13g2_fill_2 FILLER_73_504 ();
 sg13g2_decap_8 FILLER_73_510 ();
 sg13g2_fill_2 FILLER_73_517 ();
 sg13g2_decap_8 FILLER_73_524 ();
 sg13g2_fill_2 FILLER_73_531 ();
 sg13g2_decap_8 FILLER_73_537 ();
 sg13g2_fill_1 FILLER_73_544 ();
 sg13g2_decap_8 FILLER_73_550 ();
 sg13g2_decap_8 FILLER_73_557 ();
 sg13g2_decap_8 FILLER_73_564 ();
 sg13g2_decap_8 FILLER_73_571 ();
 sg13g2_decap_8 FILLER_73_578 ();
 sg13g2_decap_8 FILLER_73_585 ();
 sg13g2_decap_4 FILLER_73_592 ();
 sg13g2_fill_2 FILLER_73_596 ();
 sg13g2_decap_8 FILLER_73_624 ();
 sg13g2_decap_8 FILLER_73_631 ();
 sg13g2_decap_8 FILLER_73_638 ();
 sg13g2_decap_8 FILLER_73_645 ();
 sg13g2_decap_8 FILLER_73_652 ();
 sg13g2_decap_8 FILLER_73_659 ();
 sg13g2_decap_8 FILLER_73_666 ();
 sg13g2_fill_2 FILLER_73_673 ();
 sg13g2_decap_8 FILLER_73_680 ();
 sg13g2_decap_8 FILLER_73_687 ();
 sg13g2_decap_8 FILLER_73_694 ();
 sg13g2_decap_8 FILLER_73_701 ();
 sg13g2_decap_8 FILLER_73_708 ();
 sg13g2_decap_8 FILLER_73_715 ();
 sg13g2_decap_8 FILLER_73_722 ();
 sg13g2_decap_8 FILLER_73_729 ();
 sg13g2_decap_8 FILLER_73_736 ();
 sg13g2_fill_1 FILLER_73_743 ();
 sg13g2_decap_4 FILLER_73_748 ();
 sg13g2_fill_2 FILLER_73_752 ();
 sg13g2_decap_8 FILLER_73_758 ();
 sg13g2_decap_8 FILLER_73_765 ();
 sg13g2_decap_8 FILLER_73_772 ();
 sg13g2_decap_4 FILLER_73_779 ();
 sg13g2_decap_4 FILLER_73_793 ();
 sg13g2_fill_2 FILLER_73_797 ();
 sg13g2_decap_8 FILLER_73_804 ();
 sg13g2_decap_8 FILLER_73_811 ();
 sg13g2_decap_8 FILLER_73_818 ();
 sg13g2_decap_8 FILLER_73_825 ();
 sg13g2_decap_8 FILLER_73_832 ();
 sg13g2_decap_8 FILLER_73_839 ();
 sg13g2_decap_4 FILLER_73_846 ();
 sg13g2_fill_2 FILLER_73_850 ();
 sg13g2_decap_8 FILLER_73_856 ();
 sg13g2_decap_8 FILLER_73_863 ();
 sg13g2_decap_8 FILLER_73_870 ();
 sg13g2_decap_8 FILLER_73_877 ();
 sg13g2_decap_8 FILLER_73_884 ();
 sg13g2_fill_1 FILLER_73_891 ();
 sg13g2_decap_8 FILLER_73_896 ();
 sg13g2_decap_8 FILLER_73_903 ();
 sg13g2_fill_2 FILLER_73_910 ();
 sg13g2_decap_8 FILLER_73_920 ();
 sg13g2_fill_1 FILLER_73_927 ();
 sg13g2_decap_4 FILLER_73_933 ();
 sg13g2_decap_4 FILLER_73_942 ();
 sg13g2_decap_8 FILLER_73_951 ();
 sg13g2_fill_2 FILLER_73_962 ();
 sg13g2_decap_8 FILLER_73_969 ();
 sg13g2_decap_8 FILLER_73_976 ();
 sg13g2_decap_4 FILLER_73_994 ();
 sg13g2_fill_1 FILLER_73_998 ();
 sg13g2_fill_2 FILLER_73_1003 ();
 sg13g2_fill_1 FILLER_73_1005 ();
 sg13g2_decap_8 FILLER_73_1011 ();
 sg13g2_decap_8 FILLER_73_1023 ();
 sg13g2_decap_4 FILLER_73_1030 ();
 sg13g2_fill_1 FILLER_73_1034 ();
 sg13g2_fill_1 FILLER_73_1043 ();
 sg13g2_decap_8 FILLER_73_1050 ();
 sg13g2_decap_8 FILLER_73_1057 ();
 sg13g2_decap_8 FILLER_73_1064 ();
 sg13g2_decap_8 FILLER_73_1071 ();
 sg13g2_decap_8 FILLER_73_1078 ();
 sg13g2_decap_8 FILLER_73_1085 ();
 sg13g2_fill_2 FILLER_73_1092 ();
 sg13g2_decap_8 FILLER_73_1107 ();
 sg13g2_decap_4 FILLER_73_1135 ();
 sg13g2_fill_2 FILLER_73_1139 ();
 sg13g2_decap_4 FILLER_73_1151 ();
 sg13g2_fill_1 FILLER_73_1155 ();
 sg13g2_decap_8 FILLER_73_1160 ();
 sg13g2_decap_8 FILLER_73_1167 ();
 sg13g2_fill_2 FILLER_73_1174 ();
 sg13g2_fill_1 FILLER_73_1176 ();
 sg13g2_decap_8 FILLER_73_1182 ();
 sg13g2_fill_2 FILLER_73_1189 ();
 sg13g2_fill_2 FILLER_73_1202 ();
 sg13g2_decap_4 FILLER_73_1209 ();
 sg13g2_fill_1 FILLER_73_1213 ();
 sg13g2_decap_8 FILLER_73_1237 ();
 sg13g2_decap_4 FILLER_73_1244 ();
 sg13g2_fill_1 FILLER_73_1248 ();
 sg13g2_decap_8 FILLER_73_1254 ();
 sg13g2_fill_2 FILLER_73_1261 ();
 sg13g2_decap_8 FILLER_73_1267 ();
 sg13g2_decap_8 FILLER_73_1274 ();
 sg13g2_decap_8 FILLER_73_1281 ();
 sg13g2_decap_8 FILLER_73_1288 ();
 sg13g2_decap_8 FILLER_73_1295 ();
 sg13g2_decap_8 FILLER_73_1302 ();
 sg13g2_decap_8 FILLER_73_1309 ();
 sg13g2_decap_8 FILLER_73_1316 ();
 sg13g2_fill_2 FILLER_73_1323 ();
 sg13g2_fill_1 FILLER_73_1325 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_4 FILLER_74_28 ();
 sg13g2_fill_2 FILLER_74_32 ();
 sg13g2_fill_2 FILLER_74_52 ();
 sg13g2_decap_4 FILLER_74_75 ();
 sg13g2_decap_4 FILLER_74_97 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_4 FILLER_74_119 ();
 sg13g2_fill_2 FILLER_74_123 ();
 sg13g2_decap_8 FILLER_74_129 ();
 sg13g2_decap_8 FILLER_74_136 ();
 sg13g2_decap_8 FILLER_74_143 ();
 sg13g2_fill_1 FILLER_74_150 ();
 sg13g2_decap_4 FILLER_74_156 ();
 sg13g2_fill_1 FILLER_74_160 ();
 sg13g2_fill_2 FILLER_74_169 ();
 sg13g2_fill_1 FILLER_74_171 ();
 sg13g2_fill_2 FILLER_74_177 ();
 sg13g2_fill_1 FILLER_74_179 ();
 sg13g2_fill_2 FILLER_74_205 ();
 sg13g2_fill_2 FILLER_74_216 ();
 sg13g2_fill_2 FILLER_74_222 ();
 sg13g2_fill_1 FILLER_74_224 ();
 sg13g2_decap_4 FILLER_74_230 ();
 sg13g2_fill_1 FILLER_74_234 ();
 sg13g2_decap_4 FILLER_74_239 ();
 sg13g2_fill_2 FILLER_74_255 ();
 sg13g2_decap_8 FILLER_74_282 ();
 sg13g2_decap_8 FILLER_74_289 ();
 sg13g2_decap_8 FILLER_74_296 ();
 sg13g2_decap_8 FILLER_74_303 ();
 sg13g2_decap_8 FILLER_74_310 ();
 sg13g2_fill_2 FILLER_74_317 ();
 sg13g2_fill_1 FILLER_74_319 ();
 sg13g2_decap_8 FILLER_74_324 ();
 sg13g2_decap_8 FILLER_74_331 ();
 sg13g2_decap_8 FILLER_74_338 ();
 sg13g2_fill_2 FILLER_74_345 ();
 sg13g2_fill_1 FILLER_74_347 ();
 sg13g2_decap_4 FILLER_74_353 ();
 sg13g2_decap_8 FILLER_74_365 ();
 sg13g2_decap_8 FILLER_74_372 ();
 sg13g2_decap_8 FILLER_74_379 ();
 sg13g2_decap_8 FILLER_74_386 ();
 sg13g2_fill_1 FILLER_74_393 ();
 sg13g2_decap_8 FILLER_74_398 ();
 sg13g2_decap_8 FILLER_74_405 ();
 sg13g2_decap_8 FILLER_74_412 ();
 sg13g2_decap_4 FILLER_74_419 ();
 sg13g2_decap_4 FILLER_74_427 ();
 sg13g2_decap_8 FILLER_74_435 ();
 sg13g2_fill_1 FILLER_74_442 ();
 sg13g2_fill_2 FILLER_74_447 ();
 sg13g2_decap_8 FILLER_74_453 ();
 sg13g2_decap_8 FILLER_74_460 ();
 sg13g2_decap_8 FILLER_74_467 ();
 sg13g2_decap_8 FILLER_74_505 ();
 sg13g2_decap_8 FILLER_74_512 ();
 sg13g2_fill_1 FILLER_74_519 ();
 sg13g2_decap_8 FILLER_74_572 ();
 sg13g2_decap_8 FILLER_74_579 ();
 sg13g2_decap_8 FILLER_74_586 ();
 sg13g2_decap_8 FILLER_74_593 ();
 sg13g2_fill_2 FILLER_74_600 ();
 sg13g2_fill_1 FILLER_74_602 ();
 sg13g2_decap_8 FILLER_74_607 ();
 sg13g2_decap_8 FILLER_74_614 ();
 sg13g2_decap_8 FILLER_74_621 ();
 sg13g2_decap_8 FILLER_74_628 ();
 sg13g2_decap_8 FILLER_74_635 ();
 sg13g2_decap_4 FILLER_74_642 ();
 sg13g2_fill_2 FILLER_74_646 ();
 sg13g2_decap_8 FILLER_74_679 ();
 sg13g2_decap_8 FILLER_74_686 ();
 sg13g2_decap_8 FILLER_74_693 ();
 sg13g2_decap_8 FILLER_74_700 ();
 sg13g2_decap_4 FILLER_74_707 ();
 sg13g2_fill_2 FILLER_74_711 ();
 sg13g2_decap_8 FILLER_74_717 ();
 sg13g2_fill_2 FILLER_74_724 ();
 sg13g2_decap_8 FILLER_74_752 ();
 sg13g2_decap_8 FILLER_74_759 ();
 sg13g2_decap_8 FILLER_74_766 ();
 sg13g2_decap_8 FILLER_74_773 ();
 sg13g2_decap_8 FILLER_74_780 ();
 sg13g2_decap_8 FILLER_74_787 ();
 sg13g2_decap_8 FILLER_74_794 ();
 sg13g2_decap_8 FILLER_74_801 ();
 sg13g2_decap_8 FILLER_74_808 ();
 sg13g2_decap_8 FILLER_74_815 ();
 sg13g2_decap_8 FILLER_74_822 ();
 sg13g2_decap_8 FILLER_74_829 ();
 sg13g2_fill_1 FILLER_74_836 ();
 sg13g2_decap_8 FILLER_74_841 ();
 sg13g2_fill_2 FILLER_74_848 ();
 sg13g2_fill_1 FILLER_74_850 ();
 sg13g2_decap_8 FILLER_74_856 ();
 sg13g2_decap_8 FILLER_74_863 ();
 sg13g2_decap_4 FILLER_74_870 ();
 sg13g2_decap_8 FILLER_74_879 ();
 sg13g2_decap_8 FILLER_74_886 ();
 sg13g2_decap_8 FILLER_74_893 ();
 sg13g2_decap_8 FILLER_74_900 ();
 sg13g2_decap_4 FILLER_74_907 ();
 sg13g2_fill_1 FILLER_74_911 ();
 sg13g2_fill_2 FILLER_74_930 ();
 sg13g2_fill_1 FILLER_74_932 ();
 sg13g2_decap_8 FILLER_74_950 ();
 sg13g2_decap_8 FILLER_74_957 ();
 sg13g2_decap_8 FILLER_74_964 ();
 sg13g2_fill_2 FILLER_74_971 ();
 sg13g2_fill_1 FILLER_74_973 ();
 sg13g2_fill_2 FILLER_74_979 ();
 sg13g2_fill_1 FILLER_74_981 ();
 sg13g2_decap_8 FILLER_74_987 ();
 sg13g2_decap_8 FILLER_74_994 ();
 sg13g2_decap_8 FILLER_74_1001 ();
 sg13g2_fill_1 FILLER_74_1008 ();
 sg13g2_decap_8 FILLER_74_1014 ();
 sg13g2_decap_8 FILLER_74_1021 ();
 sg13g2_decap_8 FILLER_74_1028 ();
 sg13g2_fill_1 FILLER_74_1035 ();
 sg13g2_decap_8 FILLER_74_1044 ();
 sg13g2_decap_8 FILLER_74_1051 ();
 sg13g2_decap_8 FILLER_74_1058 ();
 sg13g2_decap_8 FILLER_74_1065 ();
 sg13g2_fill_1 FILLER_74_1072 ();
 sg13g2_decap_4 FILLER_74_1078 ();
 sg13g2_decap_8 FILLER_74_1086 ();
 sg13g2_fill_1 FILLER_74_1093 ();
 sg13g2_decap_8 FILLER_74_1103 ();
 sg13g2_decap_8 FILLER_74_1110 ();
 sg13g2_fill_2 FILLER_74_1117 ();
 sg13g2_decap_8 FILLER_74_1123 ();
 sg13g2_fill_1 FILLER_74_1130 ();
 sg13g2_decap_4 FILLER_74_1145 ();
 sg13g2_decap_8 FILLER_74_1153 ();
 sg13g2_decap_8 FILLER_74_1160 ();
 sg13g2_fill_1 FILLER_74_1167 ();
 sg13g2_decap_4 FILLER_74_1173 ();
 sg13g2_decap_8 FILLER_74_1181 ();
 sg13g2_decap_4 FILLER_74_1188 ();
 sg13g2_fill_1 FILLER_74_1192 ();
 sg13g2_decap_4 FILLER_74_1198 ();
 sg13g2_fill_1 FILLER_74_1202 ();
 sg13g2_decap_4 FILLER_74_1209 ();
 sg13g2_fill_1 FILLER_74_1213 ();
 sg13g2_fill_2 FILLER_74_1223 ();
 sg13g2_fill_2 FILLER_74_1231 ();
 sg13g2_fill_1 FILLER_74_1237 ();
 sg13g2_decap_8 FILLER_74_1243 ();
 sg13g2_decap_4 FILLER_74_1250 ();
 sg13g2_fill_2 FILLER_74_1258 ();
 sg13g2_fill_1 FILLER_74_1260 ();
 sg13g2_decap_8 FILLER_74_1275 ();
 sg13g2_decap_8 FILLER_74_1282 ();
 sg13g2_decap_8 FILLER_74_1289 ();
 sg13g2_decap_8 FILLER_74_1296 ();
 sg13g2_decap_8 FILLER_74_1303 ();
 sg13g2_decap_8 FILLER_74_1310 ();
 sg13g2_decap_8 FILLER_74_1317 ();
 sg13g2_fill_2 FILLER_74_1324 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_4 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_51 ();
 sg13g2_fill_1 FILLER_75_58 ();
 sg13g2_fill_1 FILLER_75_64 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_fill_1 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_118 ();
 sg13g2_decap_8 FILLER_75_125 ();
 sg13g2_decap_8 FILLER_75_132 ();
 sg13g2_decap_8 FILLER_75_139 ();
 sg13g2_decap_4 FILLER_75_146 ();
 sg13g2_fill_2 FILLER_75_150 ();
 sg13g2_decap_8 FILLER_75_157 ();
 sg13g2_decap_8 FILLER_75_164 ();
 sg13g2_decap_8 FILLER_75_176 ();
 sg13g2_decap_8 FILLER_75_187 ();
 sg13g2_decap_4 FILLER_75_194 ();
 sg13g2_decap_8 FILLER_75_208 ();
 sg13g2_fill_2 FILLER_75_215 ();
 sg13g2_decap_8 FILLER_75_248 ();
 sg13g2_fill_1 FILLER_75_255 ();
 sg13g2_decap_4 FILLER_75_261 ();
 sg13g2_decap_8 FILLER_75_269 ();
 sg13g2_decap_8 FILLER_75_276 ();
 sg13g2_decap_8 FILLER_75_283 ();
 sg13g2_decap_8 FILLER_75_290 ();
 sg13g2_decap_4 FILLER_75_297 ();
 sg13g2_fill_1 FILLER_75_301 ();
 sg13g2_decap_8 FILLER_75_307 ();
 sg13g2_decap_8 FILLER_75_314 ();
 sg13g2_decap_8 FILLER_75_321 ();
 sg13g2_decap_8 FILLER_75_328 ();
 sg13g2_decap_8 FILLER_75_335 ();
 sg13g2_decap_8 FILLER_75_342 ();
 sg13g2_fill_1 FILLER_75_354 ();
 sg13g2_decap_8 FILLER_75_359 ();
 sg13g2_fill_2 FILLER_75_366 ();
 sg13g2_decap_4 FILLER_75_372 ();
 sg13g2_fill_1 FILLER_75_376 ();
 sg13g2_decap_4 FILLER_75_383 ();
 sg13g2_fill_2 FILLER_75_387 ();
 sg13g2_fill_1 FILLER_75_393 ();
 sg13g2_fill_1 FILLER_75_399 ();
 sg13g2_fill_1 FILLER_75_403 ();
 sg13g2_decap_8 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_75_415 ();
 sg13g2_decap_8 FILLER_75_422 ();
 sg13g2_decap_4 FILLER_75_433 ();
 sg13g2_fill_2 FILLER_75_437 ();
 sg13g2_decap_8 FILLER_75_448 ();
 sg13g2_decap_8 FILLER_75_455 ();
 sg13g2_decap_8 FILLER_75_462 ();
 sg13g2_decap_8 FILLER_75_469 ();
 sg13g2_decap_8 FILLER_75_476 ();
 sg13g2_decap_8 FILLER_75_483 ();
 sg13g2_decap_8 FILLER_75_490 ();
 sg13g2_decap_8 FILLER_75_497 ();
 sg13g2_decap_8 FILLER_75_504 ();
 sg13g2_decap_8 FILLER_75_511 ();
 sg13g2_decap_8 FILLER_75_518 ();
 sg13g2_decap_8 FILLER_75_525 ();
 sg13g2_decap_8 FILLER_75_532 ();
 sg13g2_decap_8 FILLER_75_539 ();
 sg13g2_decap_8 FILLER_75_546 ();
 sg13g2_decap_4 FILLER_75_557 ();
 sg13g2_fill_2 FILLER_75_569 ();
 sg13g2_decap_8 FILLER_75_597 ();
 sg13g2_decap_8 FILLER_75_604 ();
 sg13g2_decap_8 FILLER_75_611 ();
 sg13g2_decap_8 FILLER_75_618 ();
 sg13g2_decap_8 FILLER_75_625 ();
 sg13g2_fill_2 FILLER_75_632 ();
 sg13g2_decap_8 FILLER_75_642 ();
 sg13g2_decap_8 FILLER_75_649 ();
 sg13g2_decap_4 FILLER_75_656 ();
 sg13g2_fill_2 FILLER_75_660 ();
 sg13g2_decap_8 FILLER_75_666 ();
 sg13g2_fill_2 FILLER_75_673 ();
 sg13g2_fill_2 FILLER_75_680 ();
 sg13g2_fill_1 FILLER_75_682 ();
 sg13g2_decap_8 FILLER_75_687 ();
 sg13g2_decap_8 FILLER_75_694 ();
 sg13g2_decap_4 FILLER_75_701 ();
 sg13g2_fill_2 FILLER_75_705 ();
 sg13g2_fill_1 FILLER_75_733 ();
 sg13g2_decap_8 FILLER_75_738 ();
 sg13g2_decap_8 FILLER_75_745 ();
 sg13g2_decap_8 FILLER_75_752 ();
 sg13g2_decap_8 FILLER_75_759 ();
 sg13g2_decap_8 FILLER_75_766 ();
 sg13g2_decap_8 FILLER_75_773 ();
 sg13g2_decap_8 FILLER_75_780 ();
 sg13g2_decap_8 FILLER_75_787 ();
 sg13g2_decap_8 FILLER_75_794 ();
 sg13g2_decap_8 FILLER_75_801 ();
 sg13g2_decap_8 FILLER_75_808 ();
 sg13g2_decap_8 FILLER_75_815 ();
 sg13g2_decap_4 FILLER_75_822 ();
 sg13g2_decap_8 FILLER_75_830 ();
 sg13g2_decap_8 FILLER_75_837 ();
 sg13g2_decap_8 FILLER_75_844 ();
 sg13g2_decap_8 FILLER_75_851 ();
 sg13g2_decap_8 FILLER_75_858 ();
 sg13g2_decap_8 FILLER_75_865 ();
 sg13g2_fill_2 FILLER_75_872 ();
 sg13g2_decap_4 FILLER_75_879 ();
 sg13g2_fill_2 FILLER_75_901 ();
 sg13g2_fill_1 FILLER_75_908 ();
 sg13g2_decap_8 FILLER_75_913 ();
 sg13g2_decap_8 FILLER_75_920 ();
 sg13g2_decap_8 FILLER_75_927 ();
 sg13g2_decap_4 FILLER_75_934 ();
 sg13g2_fill_2 FILLER_75_938 ();
 sg13g2_decap_8 FILLER_75_950 ();
 sg13g2_decap_8 FILLER_75_957 ();
 sg13g2_decap_4 FILLER_75_974 ();
 sg13g2_decap_4 FILLER_75_983 ();
 sg13g2_fill_1 FILLER_75_987 ();
 sg13g2_decap_8 FILLER_75_993 ();
 sg13g2_fill_2 FILLER_75_1000 ();
 sg13g2_fill_1 FILLER_75_1002 ();
 sg13g2_decap_8 FILLER_75_1008 ();
 sg13g2_decap_8 FILLER_75_1015 ();
 sg13g2_decap_8 FILLER_75_1022 ();
 sg13g2_decap_4 FILLER_75_1029 ();
 sg13g2_decap_4 FILLER_75_1048 ();
 sg13g2_fill_2 FILLER_75_1052 ();
 sg13g2_decap_4 FILLER_75_1064 ();
 sg13g2_decap_8 FILLER_75_1072 ();
 sg13g2_decap_4 FILLER_75_1079 ();
 sg13g2_decap_8 FILLER_75_1088 ();
 sg13g2_decap_8 FILLER_75_1095 ();
 sg13g2_fill_1 FILLER_75_1102 ();
 sg13g2_decap_8 FILLER_75_1108 ();
 sg13g2_decap_8 FILLER_75_1115 ();
 sg13g2_decap_4 FILLER_75_1122 ();
 sg13g2_fill_1 FILLER_75_1126 ();
 sg13g2_fill_2 FILLER_75_1140 ();
 sg13g2_fill_1 FILLER_75_1142 ();
 sg13g2_fill_1 FILLER_75_1154 ();
 sg13g2_decap_8 FILLER_75_1165 ();
 sg13g2_fill_2 FILLER_75_1172 ();
 sg13g2_decap_8 FILLER_75_1179 ();
 sg13g2_decap_8 FILLER_75_1186 ();
 sg13g2_decap_4 FILLER_75_1193 ();
 sg13g2_fill_2 FILLER_75_1197 ();
 sg13g2_decap_8 FILLER_75_1207 ();
 sg13g2_fill_2 FILLER_75_1214 ();
 sg13g2_decap_8 FILLER_75_1234 ();
 sg13g2_decap_8 FILLER_75_1241 ();
 sg13g2_decap_8 FILLER_75_1248 ();
 sg13g2_decap_8 FILLER_75_1255 ();
 sg13g2_decap_8 FILLER_75_1262 ();
 sg13g2_decap_8 FILLER_75_1269 ();
 sg13g2_decap_8 FILLER_75_1276 ();
 sg13g2_decap_8 FILLER_75_1283 ();
 sg13g2_decap_8 FILLER_75_1290 ();
 sg13g2_decap_8 FILLER_75_1297 ();
 sg13g2_decap_8 FILLER_75_1304 ();
 sg13g2_decap_8 FILLER_75_1311 ();
 sg13g2_decap_8 FILLER_75_1318 ();
 sg13g2_fill_1 FILLER_75_1325 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_4 FILLER_76_49 ();
 sg13g2_fill_1 FILLER_76_61 ();
 sg13g2_decap_8 FILLER_76_67 ();
 sg13g2_decap_8 FILLER_76_74 ();
 sg13g2_decap_8 FILLER_76_81 ();
 sg13g2_decap_8 FILLER_76_88 ();
 sg13g2_decap_8 FILLER_76_95 ();
 sg13g2_decap_8 FILLER_76_102 ();
 sg13g2_decap_8 FILLER_76_109 ();
 sg13g2_decap_4 FILLER_76_116 ();
 sg13g2_fill_1 FILLER_76_120 ();
 sg13g2_decap_8 FILLER_76_125 ();
 sg13g2_decap_8 FILLER_76_132 ();
 sg13g2_fill_2 FILLER_76_139 ();
 sg13g2_decap_4 FILLER_76_145 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_fill_2 FILLER_76_189 ();
 sg13g2_fill_1 FILLER_76_191 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_4 FILLER_76_231 ();
 sg13g2_fill_2 FILLER_76_235 ();
 sg13g2_fill_2 FILLER_76_242 ();
 sg13g2_decap_8 FILLER_76_283 ();
 sg13g2_decap_4 FILLER_76_290 ();
 sg13g2_fill_1 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_299 ();
 sg13g2_fill_2 FILLER_76_306 ();
 sg13g2_decap_8 FILLER_76_313 ();
 sg13g2_decap_4 FILLER_76_320 ();
 sg13g2_decap_8 FILLER_76_328 ();
 sg13g2_decap_8 FILLER_76_335 ();
 sg13g2_fill_1 FILLER_76_342 ();
 sg13g2_decap_8 FILLER_76_373 ();
 sg13g2_decap_8 FILLER_76_380 ();
 sg13g2_decap_8 FILLER_76_387 ();
 sg13g2_fill_1 FILLER_76_394 ();
 sg13g2_decap_4 FILLER_76_399 ();
 sg13g2_fill_1 FILLER_76_403 ();
 sg13g2_decap_8 FILLER_76_409 ();
 sg13g2_decap_8 FILLER_76_416 ();
 sg13g2_decap_8 FILLER_76_423 ();
 sg13g2_fill_2 FILLER_76_430 ();
 sg13g2_fill_1 FILLER_76_437 ();
 sg13g2_decap_8 FILLER_76_469 ();
 sg13g2_decap_8 FILLER_76_476 ();
 sg13g2_decap_8 FILLER_76_483 ();
 sg13g2_decap_8 FILLER_76_490 ();
 sg13g2_decap_8 FILLER_76_497 ();
 sg13g2_decap_8 FILLER_76_504 ();
 sg13g2_decap_8 FILLER_76_511 ();
 sg13g2_decap_4 FILLER_76_518 ();
 sg13g2_fill_1 FILLER_76_522 ();
 sg13g2_decap_8 FILLER_76_531 ();
 sg13g2_fill_1 FILLER_76_538 ();
 sg13g2_decap_8 FILLER_76_544 ();
 sg13g2_decap_8 FILLER_76_551 ();
 sg13g2_decap_8 FILLER_76_558 ();
 sg13g2_fill_1 FILLER_76_565 ();
 sg13g2_decap_4 FILLER_76_571 ();
 sg13g2_decap_8 FILLER_76_610 ();
 sg13g2_decap_8 FILLER_76_617 ();
 sg13g2_decap_4 FILLER_76_624 ();
 sg13g2_fill_2 FILLER_76_628 ();
 sg13g2_decap_8 FILLER_76_656 ();
 sg13g2_decap_8 FILLER_76_663 ();
 sg13g2_decap_8 FILLER_76_670 ();
 sg13g2_decap_4 FILLER_76_712 ();
 sg13g2_fill_2 FILLER_76_716 ();
 sg13g2_decap_8 FILLER_76_726 ();
 sg13g2_decap_8 FILLER_76_733 ();
 sg13g2_decap_8 FILLER_76_740 ();
 sg13g2_decap_8 FILLER_76_747 ();
 sg13g2_decap_8 FILLER_76_754 ();
 sg13g2_decap_8 FILLER_76_761 ();
 sg13g2_fill_2 FILLER_76_768 ();
 sg13g2_decap_8 FILLER_76_796 ();
 sg13g2_decap_8 FILLER_76_803 ();
 sg13g2_decap_4 FILLER_76_810 ();
 sg13g2_fill_1 FILLER_76_814 ();
 sg13g2_fill_1 FILLER_76_823 ();
 sg13g2_decap_4 FILLER_76_832 ();
 sg13g2_fill_2 FILLER_76_836 ();
 sg13g2_decap_8 FILLER_76_842 ();
 sg13g2_decap_8 FILLER_76_849 ();
 sg13g2_decap_8 FILLER_76_856 ();
 sg13g2_decap_8 FILLER_76_863 ();
 sg13g2_fill_2 FILLER_76_870 ();
 sg13g2_fill_1 FILLER_76_872 ();
 sg13g2_fill_2 FILLER_76_877 ();
 sg13g2_fill_1 FILLER_76_879 ();
 sg13g2_fill_2 FILLER_76_891 ();
 sg13g2_fill_1 FILLER_76_893 ();
 sg13g2_fill_1 FILLER_76_903 ();
 sg13g2_fill_2 FILLER_76_929 ();
 sg13g2_decap_4 FILLER_76_935 ();
 sg13g2_fill_1 FILLER_76_939 ();
 sg13g2_fill_2 FILLER_76_945 ();
 sg13g2_fill_1 FILLER_76_957 ();
 sg13g2_fill_1 FILLER_76_972 ();
 sg13g2_fill_2 FILLER_76_978 ();
 sg13g2_fill_1 FILLER_76_980 ();
 sg13g2_fill_1 FILLER_76_991 ();
 sg13g2_fill_1 FILLER_76_998 ();
 sg13g2_fill_1 FILLER_76_1005 ();
 sg13g2_fill_2 FILLER_76_1010 ();
 sg13g2_decap_8 FILLER_76_1023 ();
 sg13g2_decap_8 FILLER_76_1030 ();
 sg13g2_fill_2 FILLER_76_1037 ();
 sg13g2_decap_4 FILLER_76_1045 ();
 sg13g2_fill_1 FILLER_76_1049 ();
 sg13g2_decap_4 FILLER_76_1055 ();
 sg13g2_fill_1 FILLER_76_1059 ();
 sg13g2_decap_8 FILLER_76_1064 ();
 sg13g2_decap_8 FILLER_76_1071 ();
 sg13g2_fill_2 FILLER_76_1078 ();
 sg13g2_fill_2 FILLER_76_1088 ();
 sg13g2_fill_2 FILLER_76_1096 ();
 sg13g2_fill_1 FILLER_76_1107 ();
 sg13g2_fill_2 FILLER_76_1123 ();
 sg13g2_fill_1 FILLER_76_1125 ();
 sg13g2_fill_1 FILLER_76_1145 ();
 sg13g2_fill_1 FILLER_76_1152 ();
 sg13g2_decap_4 FILLER_76_1157 ();
 sg13g2_decap_4 FILLER_76_1164 ();
 sg13g2_fill_2 FILLER_76_1168 ();
 sg13g2_decap_4 FILLER_76_1183 ();
 sg13g2_fill_1 FILLER_76_1196 ();
 sg13g2_fill_2 FILLER_76_1206 ();
 sg13g2_decap_4 FILLER_76_1216 ();
 sg13g2_fill_2 FILLER_76_1220 ();
 sg13g2_fill_1 FILLER_76_1231 ();
 sg13g2_decap_8 FILLER_76_1241 ();
 sg13g2_decap_8 FILLER_76_1252 ();
 sg13g2_decap_8 FILLER_76_1259 ();
 sg13g2_decap_8 FILLER_76_1266 ();
 sg13g2_decap_8 FILLER_76_1273 ();
 sg13g2_decap_8 FILLER_76_1280 ();
 sg13g2_decap_8 FILLER_76_1287 ();
 sg13g2_decap_8 FILLER_76_1294 ();
 sg13g2_decap_8 FILLER_76_1301 ();
 sg13g2_decap_8 FILLER_76_1308 ();
 sg13g2_decap_8 FILLER_76_1315 ();
 sg13g2_decap_4 FILLER_76_1322 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_fill_1 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_48 ();
 sg13g2_decap_8 FILLER_77_81 ();
 sg13g2_decap_8 FILLER_77_88 ();
 sg13g2_decap_8 FILLER_77_95 ();
 sg13g2_decap_8 FILLER_77_102 ();
 sg13g2_decap_4 FILLER_77_109 ();
 sg13g2_fill_1 FILLER_77_113 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_fill_1 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_177 ();
 sg13g2_fill_1 FILLER_77_184 ();
 sg13g2_decap_8 FILLER_77_216 ();
 sg13g2_decap_8 FILLER_77_223 ();
 sg13g2_decap_8 FILLER_77_230 ();
 sg13g2_decap_8 FILLER_77_237 ();
 sg13g2_decap_8 FILLER_77_244 ();
 sg13g2_decap_8 FILLER_77_263 ();
 sg13g2_decap_8 FILLER_77_270 ();
 sg13g2_fill_1 FILLER_77_277 ();
 sg13g2_fill_1 FILLER_77_294 ();
 sg13g2_decap_4 FILLER_77_300 ();
 sg13g2_fill_1 FILLER_77_304 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_fill_2 FILLER_77_322 ();
 sg13g2_fill_1 FILLER_77_324 ();
 sg13g2_decap_8 FILLER_77_330 ();
 sg13g2_decap_8 FILLER_77_337 ();
 sg13g2_decap_8 FILLER_77_344 ();
 sg13g2_decap_8 FILLER_77_351 ();
 sg13g2_fill_1 FILLER_77_358 ();
 sg13g2_decap_4 FILLER_77_363 ();
 sg13g2_fill_1 FILLER_77_372 ();
 sg13g2_decap_8 FILLER_77_377 ();
 sg13g2_decap_8 FILLER_77_384 ();
 sg13g2_decap_4 FILLER_77_391 ();
 sg13g2_fill_1 FILLER_77_395 ();
 sg13g2_decap_4 FILLER_77_401 ();
 sg13g2_fill_2 FILLER_77_405 ();
 sg13g2_fill_2 FILLER_77_412 ();
 sg13g2_decap_8 FILLER_77_419 ();
 sg13g2_decap_8 FILLER_77_426 ();
 sg13g2_decap_8 FILLER_77_433 ();
 sg13g2_decap_8 FILLER_77_440 ();
 sg13g2_decap_8 FILLER_77_447 ();
 sg13g2_decap_8 FILLER_77_454 ();
 sg13g2_decap_8 FILLER_77_461 ();
 sg13g2_decap_8 FILLER_77_468 ();
 sg13g2_decap_8 FILLER_77_475 ();
 sg13g2_decap_4 FILLER_77_482 ();
 sg13g2_fill_1 FILLER_77_494 ();
 sg13g2_decap_8 FILLER_77_521 ();
 sg13g2_decap_8 FILLER_77_528 ();
 sg13g2_fill_1 FILLER_77_535 ();
 sg13g2_decap_8 FILLER_77_583 ();
 sg13g2_fill_1 FILLER_77_590 ();
 sg13g2_decap_8 FILLER_77_595 ();
 sg13g2_decap_8 FILLER_77_602 ();
 sg13g2_decap_8 FILLER_77_609 ();
 sg13g2_decap_8 FILLER_77_616 ();
 sg13g2_decap_8 FILLER_77_623 ();
 sg13g2_decap_4 FILLER_77_630 ();
 sg13g2_fill_2 FILLER_77_634 ();
 sg13g2_decap_8 FILLER_77_640 ();
 sg13g2_decap_8 FILLER_77_647 ();
 sg13g2_decap_8 FILLER_77_654 ();
 sg13g2_decap_8 FILLER_77_661 ();
 sg13g2_decap_8 FILLER_77_668 ();
 sg13g2_decap_8 FILLER_77_675 ();
 sg13g2_decap_8 FILLER_77_682 ();
 sg13g2_decap_8 FILLER_77_689 ();
 sg13g2_decap_8 FILLER_77_727 ();
 sg13g2_decap_8 FILLER_77_734 ();
 sg13g2_decap_8 FILLER_77_741 ();
 sg13g2_decap_8 FILLER_77_748 ();
 sg13g2_decap_8 FILLER_77_755 ();
 sg13g2_decap_8 FILLER_77_762 ();
 sg13g2_decap_8 FILLER_77_769 ();
 sg13g2_decap_8 FILLER_77_780 ();
 sg13g2_decap_8 FILLER_77_787 ();
 sg13g2_decap_8 FILLER_77_794 ();
 sg13g2_decap_8 FILLER_77_801 ();
 sg13g2_fill_2 FILLER_77_808 ();
 sg13g2_fill_1 FILLER_77_810 ();
 sg13g2_decap_8 FILLER_77_841 ();
 sg13g2_decap_8 FILLER_77_848 ();
 sg13g2_decap_8 FILLER_77_855 ();
 sg13g2_decap_8 FILLER_77_862 ();
 sg13g2_decap_8 FILLER_77_869 ();
 sg13g2_decap_8 FILLER_77_876 ();
 sg13g2_fill_1 FILLER_77_892 ();
 sg13g2_fill_1 FILLER_77_917 ();
 sg13g2_fill_1 FILLER_77_927 ();
 sg13g2_fill_1 FILLER_77_933 ();
 sg13g2_fill_1 FILLER_77_939 ();
 sg13g2_fill_2 FILLER_77_950 ();
 sg13g2_fill_2 FILLER_77_958 ();
 sg13g2_fill_1 FILLER_77_980 ();
 sg13g2_fill_1 FILLER_77_986 ();
 sg13g2_fill_2 FILLER_77_993 ();
 sg13g2_fill_2 FILLER_77_1000 ();
 sg13g2_fill_1 FILLER_77_1002 ();
 sg13g2_decap_4 FILLER_77_1018 ();
 sg13g2_fill_1 FILLER_77_1022 ();
 sg13g2_fill_2 FILLER_77_1037 ();
 sg13g2_fill_1 FILLER_77_1071 ();
 sg13g2_fill_1 FILLER_77_1077 ();
 sg13g2_fill_2 FILLER_77_1084 ();
 sg13g2_decap_8 FILLER_77_1091 ();
 sg13g2_decap_8 FILLER_77_1098 ();
 sg13g2_decap_8 FILLER_77_1110 ();
 sg13g2_decap_8 FILLER_77_1117 ();
 sg13g2_fill_2 FILLER_77_1165 ();
 sg13g2_fill_1 FILLER_77_1167 ();
 sg13g2_fill_1 FILLER_77_1178 ();
 sg13g2_decap_8 FILLER_77_1187 ();
 sg13g2_fill_1 FILLER_77_1194 ();
 sg13g2_decap_4 FILLER_77_1200 ();
 sg13g2_decap_8 FILLER_77_1213 ();
 sg13g2_decap_4 FILLER_77_1224 ();
 sg13g2_fill_2 FILLER_77_1228 ();
 sg13g2_fill_1 FILLER_77_1234 ();
 sg13g2_decap_8 FILLER_77_1244 ();
 sg13g2_decap_8 FILLER_77_1251 ();
 sg13g2_decap_8 FILLER_77_1258 ();
 sg13g2_decap_8 FILLER_77_1265 ();
 sg13g2_decap_8 FILLER_77_1272 ();
 sg13g2_decap_8 FILLER_77_1279 ();
 sg13g2_decap_8 FILLER_77_1286 ();
 sg13g2_decap_8 FILLER_77_1293 ();
 sg13g2_decap_8 FILLER_77_1300 ();
 sg13g2_decap_8 FILLER_77_1307 ();
 sg13g2_decap_8 FILLER_77_1314 ();
 sg13g2_decap_4 FILLER_77_1321 ();
 sg13g2_fill_1 FILLER_77_1325 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_fill_1 FILLER_78_28 ();
 sg13g2_fill_2 FILLER_78_33 ();
 sg13g2_fill_1 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_66 ();
 sg13g2_decap_8 FILLER_78_73 ();
 sg13g2_fill_2 FILLER_78_80 ();
 sg13g2_fill_1 FILLER_78_82 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_4 FILLER_78_140 ();
 sg13g2_fill_1 FILLER_78_144 ();
 sg13g2_decap_8 FILLER_78_171 ();
 sg13g2_decap_8 FILLER_78_178 ();
 sg13g2_decap_8 FILLER_78_185 ();
 sg13g2_decap_8 FILLER_78_192 ();
 sg13g2_decap_8 FILLER_78_199 ();
 sg13g2_fill_2 FILLER_78_232 ();
 sg13g2_decap_4 FILLER_78_239 ();
 sg13g2_fill_1 FILLER_78_243 ();
 sg13g2_fill_2 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_283 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_fill_2 FILLER_78_336 ();
 sg13g2_fill_1 FILLER_78_338 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_4 FILLER_78_350 ();
 sg13g2_fill_2 FILLER_78_354 ();
 sg13g2_fill_2 FILLER_78_387 ();
 sg13g2_decap_8 FILLER_78_400 ();
 sg13g2_fill_1 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_78_418 ();
 sg13g2_fill_1 FILLER_78_435 ();
 sg13g2_fill_1 FILLER_78_441 ();
 sg13g2_fill_1 FILLER_78_447 ();
 sg13g2_decap_4 FILLER_78_474 ();
 sg13g2_decap_8 FILLER_78_483 ();
 sg13g2_fill_2 FILLER_78_490 ();
 sg13g2_fill_1 FILLER_78_492 ();
 sg13g2_decap_4 FILLER_78_497 ();
 sg13g2_decap_8 FILLER_78_531 ();
 sg13g2_decap_4 FILLER_78_538 ();
 sg13g2_decap_8 FILLER_78_572 ();
 sg13g2_fill_2 FILLER_78_579 ();
 sg13g2_fill_1 FILLER_78_581 ();
 sg13g2_decap_8 FILLER_78_586 ();
 sg13g2_decap_4 FILLER_78_593 ();
 sg13g2_fill_1 FILLER_78_597 ();
 sg13g2_decap_4 FILLER_78_603 ();
 sg13g2_fill_2 FILLER_78_607 ();
 sg13g2_decap_8 FILLER_78_613 ();
 sg13g2_decap_4 FILLER_78_620 ();
 sg13g2_fill_1 FILLER_78_624 ();
 sg13g2_fill_2 FILLER_78_630 ();
 sg13g2_fill_1 FILLER_78_632 ();
 sg13g2_decap_8 FILLER_78_637 ();
 sg13g2_decap_4 FILLER_78_644 ();
 sg13g2_fill_2 FILLER_78_648 ();
 sg13g2_decap_4 FILLER_78_655 ();
 sg13g2_fill_1 FILLER_78_659 ();
 sg13g2_decap_8 FILLER_78_669 ();
 sg13g2_fill_1 FILLER_78_676 ();
 sg13g2_decap_4 FILLER_78_682 ();
 sg13g2_decap_8 FILLER_78_690 ();
 sg13g2_decap_8 FILLER_78_697 ();
 sg13g2_decap_8 FILLER_78_704 ();
 sg13g2_decap_8 FILLER_78_711 ();
 sg13g2_fill_2 FILLER_78_718 ();
 sg13g2_fill_1 FILLER_78_720 ();
 sg13g2_decap_8 FILLER_78_725 ();
 sg13g2_decap_8 FILLER_78_732 ();
 sg13g2_fill_1 FILLER_78_739 ();
 sg13g2_decap_8 FILLER_78_766 ();
 sg13g2_decap_8 FILLER_78_773 ();
 sg13g2_fill_2 FILLER_78_780 ();
 sg13g2_decap_8 FILLER_78_808 ();
 sg13g2_decap_8 FILLER_78_815 ();
 sg13g2_fill_2 FILLER_78_830 ();
 sg13g2_fill_1 FILLER_78_832 ();
 sg13g2_decap_8 FILLER_78_837 ();
 sg13g2_fill_2 FILLER_78_844 ();
 sg13g2_fill_1 FILLER_78_846 ();
 sg13g2_decap_8 FILLER_78_852 ();
 sg13g2_decap_8 FILLER_78_859 ();
 sg13g2_decap_8 FILLER_78_866 ();
 sg13g2_decap_8 FILLER_78_873 ();
 sg13g2_decap_8 FILLER_78_880 ();
 sg13g2_decap_8 FILLER_78_887 ();
 sg13g2_decap_8 FILLER_78_894 ();
 sg13g2_decap_8 FILLER_78_901 ();
 sg13g2_decap_8 FILLER_78_908 ();
 sg13g2_decap_4 FILLER_78_915 ();
 sg13g2_decap_8 FILLER_78_923 ();
 sg13g2_decap_4 FILLER_78_930 ();
 sg13g2_fill_1 FILLER_78_934 ();
 sg13g2_decap_4 FILLER_78_940 ();
 sg13g2_fill_1 FILLER_78_944 ();
 sg13g2_fill_2 FILLER_78_949 ();
 sg13g2_fill_1 FILLER_78_956 ();
 sg13g2_fill_2 FILLER_78_962 ();
 sg13g2_decap_8 FILLER_78_969 ();
 sg13g2_decap_8 FILLER_78_976 ();
 sg13g2_decap_8 FILLER_78_983 ();
 sg13g2_fill_1 FILLER_78_990 ();
 sg13g2_decap_8 FILLER_78_1002 ();
 sg13g2_decap_8 FILLER_78_1009 ();
 sg13g2_decap_8 FILLER_78_1016 ();
 sg13g2_decap_8 FILLER_78_1023 ();
 sg13g2_decap_8 FILLER_78_1030 ();
 sg13g2_decap_8 FILLER_78_1037 ();
 sg13g2_decap_8 FILLER_78_1044 ();
 sg13g2_decap_8 FILLER_78_1051 ();
 sg13g2_fill_2 FILLER_78_1058 ();
 sg13g2_fill_1 FILLER_78_1072 ();
 sg13g2_fill_1 FILLER_78_1078 ();
 sg13g2_fill_2 FILLER_78_1083 ();
 sg13g2_decap_8 FILLER_78_1088 ();
 sg13g2_decap_8 FILLER_78_1095 ();
 sg13g2_decap_8 FILLER_78_1102 ();
 sg13g2_decap_8 FILLER_78_1109 ();
 sg13g2_fill_2 FILLER_78_1116 ();
 sg13g2_fill_1 FILLER_78_1122 ();
 sg13g2_fill_1 FILLER_78_1133 ();
 sg13g2_fill_1 FILLER_78_1142 ();
 sg13g2_fill_1 FILLER_78_1151 ();
 sg13g2_decap_8 FILLER_78_1162 ();
 sg13g2_decap_8 FILLER_78_1169 ();
 sg13g2_decap_4 FILLER_78_1176 ();
 sg13g2_fill_1 FILLER_78_1180 ();
 sg13g2_decap_8 FILLER_78_1186 ();
 sg13g2_decap_8 FILLER_78_1193 ();
 sg13g2_fill_1 FILLER_78_1200 ();
 sg13g2_decap_8 FILLER_78_1205 ();
 sg13g2_decap_8 FILLER_78_1212 ();
 sg13g2_decap_8 FILLER_78_1219 ();
 sg13g2_decap_8 FILLER_78_1226 ();
 sg13g2_decap_8 FILLER_78_1233 ();
 sg13g2_decap_8 FILLER_78_1240 ();
 sg13g2_decap_8 FILLER_78_1247 ();
 sg13g2_decap_8 FILLER_78_1254 ();
 sg13g2_decap_8 FILLER_78_1261 ();
 sg13g2_decap_8 FILLER_78_1268 ();
 sg13g2_decap_8 FILLER_78_1275 ();
 sg13g2_decap_8 FILLER_78_1282 ();
 sg13g2_decap_8 FILLER_78_1289 ();
 sg13g2_decap_8 FILLER_78_1296 ();
 sg13g2_decap_8 FILLER_78_1303 ();
 sg13g2_decap_8 FILLER_78_1310 ();
 sg13g2_decap_8 FILLER_78_1317 ();
 sg13g2_fill_2 FILLER_78_1324 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_4 FILLER_79_35 ();
 sg13g2_fill_2 FILLER_79_39 ();
 sg13g2_decap_8 FILLER_79_45 ();
 sg13g2_decap_8 FILLER_79_52 ();
 sg13g2_decap_4 FILLER_79_59 ();
 sg13g2_fill_2 FILLER_79_89 ();
 sg13g2_fill_1 FILLER_79_91 ();
 sg13g2_decap_4 FILLER_79_100 ();
 sg13g2_decap_8 FILLER_79_108 ();
 sg13g2_decap_8 FILLER_79_115 ();
 sg13g2_decap_8 FILLER_79_122 ();
 sg13g2_decap_8 FILLER_79_129 ();
 sg13g2_decap_8 FILLER_79_136 ();
 sg13g2_decap_8 FILLER_79_143 ();
 sg13g2_decap_8 FILLER_79_150 ();
 sg13g2_decap_8 FILLER_79_157 ();
 sg13g2_decap_8 FILLER_79_164 ();
 sg13g2_decap_8 FILLER_79_171 ();
 sg13g2_decap_8 FILLER_79_190 ();
 sg13g2_decap_8 FILLER_79_197 ();
 sg13g2_decap_8 FILLER_79_204 ();
 sg13g2_fill_2 FILLER_79_211 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_fill_1 FILLER_79_238 ();
 sg13g2_fill_1 FILLER_79_255 ();
 sg13g2_fill_1 FILLER_79_262 ();
 sg13g2_fill_1 FILLER_79_282 ();
 sg13g2_fill_1 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_311 ();
 sg13g2_fill_1 FILLER_79_318 ();
 sg13g2_decap_8 FILLER_79_349 ();
 sg13g2_decap_8 FILLER_79_356 ();
 sg13g2_decap_8 FILLER_79_363 ();
 sg13g2_decap_8 FILLER_79_374 ();
 sg13g2_decap_8 FILLER_79_381 ();
 sg13g2_decap_4 FILLER_79_388 ();
 sg13g2_decap_8 FILLER_79_418 ();
 sg13g2_decap_4 FILLER_79_451 ();
 sg13g2_decap_4 FILLER_79_459 ();
 sg13g2_fill_1 FILLER_79_463 ();
 sg13g2_decap_8 FILLER_79_469 ();
 sg13g2_decap_8 FILLER_79_476 ();
 sg13g2_decap_4 FILLER_79_509 ();
 sg13g2_fill_1 FILLER_79_513 ();
 sg13g2_fill_2 FILLER_79_518 ();
 sg13g2_decap_8 FILLER_79_525 ();
 sg13g2_decap_8 FILLER_79_532 ();
 sg13g2_decap_8 FILLER_79_539 ();
 sg13g2_decap_4 FILLER_79_546 ();
 sg13g2_fill_1 FILLER_79_550 ();
 sg13g2_decap_8 FILLER_79_555 ();
 sg13g2_decap_8 FILLER_79_562 ();
 sg13g2_fill_1 FILLER_79_569 ();
 sg13g2_decap_8 FILLER_79_705 ();
 sg13g2_fill_2 FILLER_79_712 ();
 sg13g2_fill_1 FILLER_79_740 ();
 sg13g2_fill_1 FILLER_79_745 ();
 sg13g2_decap_4 FILLER_79_772 ();
 sg13g2_fill_1 FILLER_79_776 ();
 sg13g2_decap_8 FILLER_79_811 ();
 sg13g2_decap_8 FILLER_79_818 ();
 sg13g2_fill_2 FILLER_79_825 ();
 sg13g2_decap_8 FILLER_79_853 ();
 sg13g2_decap_8 FILLER_79_860 ();
 sg13g2_decap_8 FILLER_79_867 ();
 sg13g2_decap_8 FILLER_79_874 ();
 sg13g2_decap_8 FILLER_79_881 ();
 sg13g2_decap_8 FILLER_79_888 ();
 sg13g2_decap_8 FILLER_79_895 ();
 sg13g2_decap_8 FILLER_79_902 ();
 sg13g2_decap_8 FILLER_79_909 ();
 sg13g2_decap_8 FILLER_79_916 ();
 sg13g2_decap_8 FILLER_79_923 ();
 sg13g2_decap_8 FILLER_79_930 ();
 sg13g2_decap_8 FILLER_79_937 ();
 sg13g2_decap_8 FILLER_79_944 ();
 sg13g2_decap_8 FILLER_79_951 ();
 sg13g2_decap_8 FILLER_79_958 ();
 sg13g2_decap_8 FILLER_79_965 ();
 sg13g2_decap_8 FILLER_79_972 ();
 sg13g2_decap_8 FILLER_79_979 ();
 sg13g2_decap_8 FILLER_79_986 ();
 sg13g2_decap_8 FILLER_79_993 ();
 sg13g2_decap_8 FILLER_79_1000 ();
 sg13g2_decap_8 FILLER_79_1007 ();
 sg13g2_decap_8 FILLER_79_1014 ();
 sg13g2_decap_8 FILLER_79_1021 ();
 sg13g2_decap_8 FILLER_79_1028 ();
 sg13g2_decap_8 FILLER_79_1035 ();
 sg13g2_decap_8 FILLER_79_1042 ();
 sg13g2_decap_8 FILLER_79_1049 ();
 sg13g2_decap_8 FILLER_79_1056 ();
 sg13g2_decap_8 FILLER_79_1063 ();
 sg13g2_decap_8 FILLER_79_1070 ();
 sg13g2_decap_8 FILLER_79_1077 ();
 sg13g2_decap_8 FILLER_79_1084 ();
 sg13g2_decap_8 FILLER_79_1091 ();
 sg13g2_decap_8 FILLER_79_1098 ();
 sg13g2_decap_8 FILLER_79_1105 ();
 sg13g2_decap_8 FILLER_79_1112 ();
 sg13g2_decap_8 FILLER_79_1119 ();
 sg13g2_fill_2 FILLER_79_1126 ();
 sg13g2_decap_8 FILLER_79_1133 ();
 sg13g2_decap_8 FILLER_79_1140 ();
 sg13g2_decap_8 FILLER_79_1147 ();
 sg13g2_decap_8 FILLER_79_1154 ();
 sg13g2_decap_8 FILLER_79_1161 ();
 sg13g2_decap_8 FILLER_79_1168 ();
 sg13g2_decap_8 FILLER_79_1175 ();
 sg13g2_decap_8 FILLER_79_1182 ();
 sg13g2_decap_8 FILLER_79_1189 ();
 sg13g2_decap_8 FILLER_79_1196 ();
 sg13g2_decap_8 FILLER_79_1203 ();
 sg13g2_decap_8 FILLER_79_1210 ();
 sg13g2_decap_8 FILLER_79_1217 ();
 sg13g2_decap_8 FILLER_79_1224 ();
 sg13g2_decap_8 FILLER_79_1231 ();
 sg13g2_decap_8 FILLER_79_1238 ();
 sg13g2_decap_8 FILLER_79_1245 ();
 sg13g2_decap_8 FILLER_79_1252 ();
 sg13g2_decap_8 FILLER_79_1259 ();
 sg13g2_decap_8 FILLER_79_1266 ();
 sg13g2_decap_8 FILLER_79_1273 ();
 sg13g2_decap_8 FILLER_79_1280 ();
 sg13g2_decap_8 FILLER_79_1287 ();
 sg13g2_decap_8 FILLER_79_1294 ();
 sg13g2_decap_8 FILLER_79_1301 ();
 sg13g2_decap_8 FILLER_79_1308 ();
 sg13g2_decap_8 FILLER_79_1315 ();
 sg13g2_decap_4 FILLER_79_1322 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_2 FILLER_80_70 ();
 sg13g2_decap_8 FILLER_80_76 ();
 sg13g2_fill_1 FILLER_80_83 ();
 sg13g2_decap_4 FILLER_80_96 ();
 sg13g2_fill_2 FILLER_80_104 ();
 sg13g2_fill_1 FILLER_80_118 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_decap_8 FILLER_80_136 ();
 sg13g2_decap_8 FILLER_80_143 ();
 sg13g2_decap_4 FILLER_80_150 ();
 sg13g2_fill_2 FILLER_80_154 ();
 sg13g2_decap_4 FILLER_80_160 ();
 sg13g2_fill_2 FILLER_80_180 ();
 sg13g2_fill_2 FILLER_80_190 ();
 sg13g2_decap_8 FILLER_80_200 ();
 sg13g2_decap_4 FILLER_80_207 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_4 FILLER_80_222 ();
 sg13g2_fill_1 FILLER_80_226 ();
 sg13g2_fill_2 FILLER_80_240 ();
 sg13g2_fill_1 FILLER_80_263 ();
 sg13g2_fill_2 FILLER_80_275 ();
 sg13g2_fill_2 FILLER_80_284 ();
 sg13g2_fill_2 FILLER_80_307 ();
 sg13g2_decap_4 FILLER_80_313 ();
 sg13g2_decap_8 FILLER_80_321 ();
 sg13g2_fill_2 FILLER_80_328 ();
 sg13g2_fill_1 FILLER_80_338 ();
 sg13g2_decap_8 FILLER_80_343 ();
 sg13g2_decap_8 FILLER_80_350 ();
 sg13g2_fill_2 FILLER_80_357 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_decap_4 FILLER_80_373 ();
 sg13g2_fill_2 FILLER_80_381 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_fill_1 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_403 ();
 sg13g2_fill_1 FILLER_80_410 ();
 sg13g2_decap_4 FILLER_80_415 ();
 sg13g2_fill_1 FILLER_80_419 ();
 sg13g2_decap_8 FILLER_80_424 ();
 sg13g2_fill_2 FILLER_80_431 ();
 sg13g2_fill_1 FILLER_80_433 ();
 sg13g2_decap_8 FILLER_80_438 ();
 sg13g2_decap_8 FILLER_80_445 ();
 sg13g2_decap_8 FILLER_80_452 ();
 sg13g2_decap_8 FILLER_80_459 ();
 sg13g2_decap_8 FILLER_80_466 ();
 sg13g2_decap_8 FILLER_80_473 ();
 sg13g2_decap_8 FILLER_80_480 ();
 sg13g2_decap_8 FILLER_80_487 ();
 sg13g2_decap_8 FILLER_80_494 ();
 sg13g2_decap_8 FILLER_80_501 ();
 sg13g2_decap_8 FILLER_80_508 ();
 sg13g2_decap_8 FILLER_80_515 ();
 sg13g2_decap_8 FILLER_80_522 ();
 sg13g2_decap_8 FILLER_80_529 ();
 sg13g2_decap_8 FILLER_80_536 ();
 sg13g2_decap_8 FILLER_80_543 ();
 sg13g2_decap_8 FILLER_80_550 ();
 sg13g2_decap_8 FILLER_80_557 ();
 sg13g2_decap_8 FILLER_80_564 ();
 sg13g2_decap_8 FILLER_80_571 ();
 sg13g2_decap_8 FILLER_80_578 ();
 sg13g2_decap_8 FILLER_80_585 ();
 sg13g2_decap_8 FILLER_80_592 ();
 sg13g2_decap_8 FILLER_80_599 ();
 sg13g2_decap_8 FILLER_80_606 ();
 sg13g2_decap_8 FILLER_80_613 ();
 sg13g2_decap_8 FILLER_80_620 ();
 sg13g2_decap_8 FILLER_80_627 ();
 sg13g2_decap_8 FILLER_80_634 ();
 sg13g2_decap_8 FILLER_80_641 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_669 ();
 sg13g2_decap_8 FILLER_80_676 ();
 sg13g2_decap_8 FILLER_80_683 ();
 sg13g2_decap_8 FILLER_80_690 ();
 sg13g2_decap_8 FILLER_80_697 ();
 sg13g2_decap_8 FILLER_80_704 ();
 sg13g2_decap_8 FILLER_80_711 ();
 sg13g2_decap_8 FILLER_80_718 ();
 sg13g2_decap_8 FILLER_80_725 ();
 sg13g2_decap_8 FILLER_80_732 ();
 sg13g2_decap_8 FILLER_80_739 ();
 sg13g2_decap_8 FILLER_80_746 ();
 sg13g2_fill_2 FILLER_80_753 ();
 sg13g2_decap_8 FILLER_80_759 ();
 sg13g2_decap_8 FILLER_80_766 ();
 sg13g2_decap_8 FILLER_80_773 ();
 sg13g2_decap_4 FILLER_80_780 ();
 sg13g2_fill_2 FILLER_80_788 ();
 sg13g2_decap_8 FILLER_80_798 ();
 sg13g2_decap_8 FILLER_80_805 ();
 sg13g2_decap_8 FILLER_80_812 ();
 sg13g2_decap_8 FILLER_80_819 ();
 sg13g2_decap_8 FILLER_80_826 ();
 sg13g2_decap_8 FILLER_80_833 ();
 sg13g2_decap_8 FILLER_80_840 ();
 sg13g2_decap_8 FILLER_80_847 ();
 sg13g2_decap_8 FILLER_80_854 ();
 sg13g2_decap_8 FILLER_80_861 ();
 sg13g2_decap_8 FILLER_80_868 ();
 sg13g2_decap_8 FILLER_80_875 ();
 sg13g2_decap_8 FILLER_80_882 ();
 sg13g2_decap_8 FILLER_80_889 ();
 sg13g2_decap_8 FILLER_80_896 ();
 sg13g2_decap_8 FILLER_80_903 ();
 sg13g2_decap_8 FILLER_80_910 ();
 sg13g2_decap_8 FILLER_80_917 ();
 sg13g2_decap_8 FILLER_80_924 ();
 sg13g2_decap_8 FILLER_80_931 ();
 sg13g2_decap_8 FILLER_80_938 ();
 sg13g2_decap_8 FILLER_80_945 ();
 sg13g2_decap_8 FILLER_80_952 ();
 sg13g2_decap_8 FILLER_80_959 ();
 sg13g2_decap_8 FILLER_80_966 ();
 sg13g2_decap_8 FILLER_80_973 ();
 sg13g2_decap_8 FILLER_80_980 ();
 sg13g2_decap_8 FILLER_80_987 ();
 sg13g2_decap_8 FILLER_80_994 ();
 sg13g2_decap_8 FILLER_80_1001 ();
 sg13g2_decap_8 FILLER_80_1008 ();
 sg13g2_decap_8 FILLER_80_1015 ();
 sg13g2_decap_8 FILLER_80_1022 ();
 sg13g2_decap_8 FILLER_80_1029 ();
 sg13g2_decap_8 FILLER_80_1036 ();
 sg13g2_decap_8 FILLER_80_1043 ();
 sg13g2_decap_8 FILLER_80_1050 ();
 sg13g2_decap_8 FILLER_80_1057 ();
 sg13g2_decap_8 FILLER_80_1064 ();
 sg13g2_decap_8 FILLER_80_1071 ();
 sg13g2_decap_8 FILLER_80_1078 ();
 sg13g2_decap_8 FILLER_80_1085 ();
 sg13g2_decap_8 FILLER_80_1092 ();
 sg13g2_decap_8 FILLER_80_1099 ();
 sg13g2_decap_8 FILLER_80_1106 ();
 sg13g2_decap_8 FILLER_80_1113 ();
 sg13g2_decap_8 FILLER_80_1120 ();
 sg13g2_decap_8 FILLER_80_1127 ();
 sg13g2_decap_8 FILLER_80_1134 ();
 sg13g2_decap_8 FILLER_80_1141 ();
 sg13g2_decap_8 FILLER_80_1148 ();
 sg13g2_decap_8 FILLER_80_1155 ();
 sg13g2_decap_8 FILLER_80_1162 ();
 sg13g2_decap_8 FILLER_80_1169 ();
 sg13g2_decap_8 FILLER_80_1176 ();
 sg13g2_decap_8 FILLER_80_1183 ();
 sg13g2_decap_8 FILLER_80_1190 ();
 sg13g2_decap_8 FILLER_80_1197 ();
 sg13g2_decap_8 FILLER_80_1204 ();
 sg13g2_decap_8 FILLER_80_1211 ();
 sg13g2_decap_8 FILLER_80_1218 ();
 sg13g2_decap_8 FILLER_80_1225 ();
 sg13g2_decap_8 FILLER_80_1232 ();
 sg13g2_decap_8 FILLER_80_1239 ();
 sg13g2_decap_8 FILLER_80_1246 ();
 sg13g2_decap_8 FILLER_80_1253 ();
 sg13g2_decap_8 FILLER_80_1260 ();
 sg13g2_decap_8 FILLER_80_1267 ();
 sg13g2_decap_8 FILLER_80_1274 ();
 sg13g2_decap_8 FILLER_80_1281 ();
 sg13g2_decap_8 FILLER_80_1288 ();
 sg13g2_decap_8 FILLER_80_1295 ();
 sg13g2_decap_8 FILLER_80_1302 ();
 sg13g2_decap_8 FILLER_80_1309 ();
 sg13g2_decap_8 FILLER_80_1316 ();
 sg13g2_fill_2 FILLER_80_1323 ();
 sg13g2_fill_1 FILLER_80_1325 ();
endmodule
