module tt_um_MichaelBell_rle_vga (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire clknet_leaf_0_clk;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire net300;
 wire net91;
 wire \addr[10] ;
 wire \addr[11] ;
 wire \addr[12] ;
 wire \addr[13] ;
 wire \addr[14] ;
 wire \addr[15] ;
 wire \addr[16] ;
 wire \addr[17] ;
 wire \addr[18] ;
 wire \addr[19] ;
 wire \addr[1] ;
 wire \addr[20] ;
 wire \addr[21] ;
 wire \addr[22] ;
 wire \addr[23] ;
 wire \addr[2] ;
 wire \addr[3] ;
 wire \addr[4] ;
 wire \addr[5] ;
 wire \addr[6] ;
 wire \addr[7] ;
 wire \addr[8] ;
 wire \addr[9] ;
 wire \addr_offset1[1] ;
 wire \addr_offset1[2] ;
 wire \addr_offset1[3] ;
 wire \addr_offset1[4] ;
 wire \addr_offset1[5] ;
 wire \addr_offset1[6] ;
 wire \addr_offset1[7] ;
 wire \addr_offset1[8] ;
 wire \addr_saved0[10] ;
 wire \addr_saved0[11] ;
 wire \addr_saved0[12] ;
 wire \addr_saved0[13] ;
 wire \addr_saved0[14] ;
 wire \addr_saved0[15] ;
 wire \addr_saved0[16] ;
 wire \addr_saved0[17] ;
 wire \addr_saved0[18] ;
 wire \addr_saved0[19] ;
 wire \addr_saved0[1] ;
 wire \addr_saved0[20] ;
 wire \addr_saved0[21] ;
 wire \addr_saved0[22] ;
 wire \addr_saved0[23] ;
 wire \addr_saved0[2] ;
 wire \addr_saved0[3] ;
 wire \addr_saved0[4] ;
 wire \addr_saved0[5] ;
 wire \addr_saved0[6] ;
 wire \addr_saved0[7] ;
 wire \addr_saved0[8] ;
 wire \addr_saved0[9] ;
 wire clear_addr;
 wire \i_spi.addr[10] ;
 wire \i_spi.addr[11] ;
 wire \i_spi.addr[12] ;
 wire \i_spi.addr[13] ;
 wire \i_spi.addr[14] ;
 wire \i_spi.addr[15] ;
 wire \i_spi.addr[16] ;
 wire \i_spi.addr[17] ;
 wire \i_spi.addr[18] ;
 wire \i_spi.addr[19] ;
 wire \i_spi.addr[1] ;
 wire \i_spi.addr[20] ;
 wire \i_spi.addr[21] ;
 wire \i_spi.addr[22] ;
 wire \i_spi.addr[23] ;
 wire \i_spi.addr[2] ;
 wire \i_spi.addr[3] ;
 wire \i_spi.addr[4] ;
 wire \i_spi.addr[5] ;
 wire \i_spi.addr[6] ;
 wire \i_spi.addr[7] ;
 wire \i_spi.addr[8] ;
 wire \i_spi.addr[9] ;
 wire \i_spi.bits_remaining[0] ;
 wire \i_spi.bits_remaining[1] ;
 wire \i_spi.bits_remaining[2] ;
 wire \i_spi.bits_remaining[3] ;
 wire \i_spi.bits_remaining[4] ;
 wire \i_spi.data[0] ;
 wire \i_spi.data[10] ;
 wire \i_spi.data[11] ;
 wire \i_spi.data[12] ;
 wire \i_spi.data[13] ;
 wire \i_spi.data[14] ;
 wire \i_spi.data[15] ;
 wire \i_spi.data[1] ;
 wire \i_spi.data[2] ;
 wire \i_spi.data[3] ;
 wire \i_spi.data[4] ;
 wire \i_spi.data[5] ;
 wire \i_spi.data[6] ;
 wire \i_spi.data[7] ;
 wire \i_spi.data[8] ;
 wire \i_spi.data[9] ;
 wire \i_spi.fsm_state[0] ;
 wire \i_spi.fsm_state[1] ;
 wire \i_spi.fsm_state[2] ;
 wire \i_spi.spi_clk_out ;
 wire \i_spi.spi_data_oe[0] ;
 wire \i_spi.spi_miso_buf_n[0] ;
 wire \i_spi.spi_miso_buf_n[1] ;
 wire \i_spi.spi_miso_buf_n[2] ;
 wire \i_spi.spi_miso_buf_n[3] ;
 wire \i_spi.spi_miso_buf_n[4] ;
 wire \i_spi.spi_miso_buf_n[5] ;
 wire \i_spi.spi_miso_buf_n[6] ;
 wire \i_spi.spi_miso_buf_n[7] ;
 wire \i_spi.spi_miso_buf_p[0] ;
 wire \i_spi.spi_miso_buf_p[1] ;
 wire \i_spi.spi_miso_buf_p[2] ;
 wire \i_spi.spi_miso_buf_p[3] ;
 wire \i_spi.spi_miso_buf_p[4] ;
 wire \i_spi.spi_miso_buf_p[5] ;
 wire \i_spi.spi_miso_buf_p[6] ;
 wire \i_spi.spi_miso_buf_p[7] ;
 wire \i_spi.spi_mosi ;
 wire \i_spi.spi_select ;
 wire \i_spi_buf.empty ;
 wire \i_spi_buf.fifo[0] ;
 wire \i_spi_buf.fifo[10] ;
 wire \i_spi_buf.fifo[11] ;
 wire \i_spi_buf.fifo[12] ;
 wire \i_spi_buf.fifo[13] ;
 wire \i_spi_buf.fifo[14] ;
 wire \i_spi_buf.fifo[15] ;
 wire \i_spi_buf.fifo[1] ;
 wire \i_spi_buf.fifo[2] ;
 wire \i_spi_buf.fifo[3] ;
 wire \i_spi_buf.fifo[4] ;
 wire \i_spi_buf.fifo[5] ;
 wire \i_spi_buf.fifo[6] ;
 wire \i_spi_buf.fifo[7] ;
 wire \i_spi_buf.fifo[8] ;
 wire \i_spi_buf.fifo[9] ;
 wire \i_spi_buf.prev_empty ;
 wire \i_spi_buf0.fifo[0] ;
 wire \i_spi_buf0.fifo[10] ;
 wire \i_spi_buf0.fifo[11] ;
 wire \i_spi_buf0.fifo[12] ;
 wire \i_spi_buf0.fifo[13] ;
 wire \i_spi_buf0.fifo[14] ;
 wire \i_spi_buf0.fifo[15] ;
 wire \i_spi_buf0.fifo[1] ;
 wire \i_spi_buf0.fifo[2] ;
 wire \i_spi_buf0.fifo[3] ;
 wire \i_spi_buf0.fifo[4] ;
 wire \i_spi_buf0.fifo[5] ;
 wire \i_spi_buf0.fifo[6] ;
 wire \i_spi_buf0.fifo[7] ;
 wire \i_spi_buf0.fifo[8] ;
 wire \i_spi_buf0.fifo[9] ;
 wire \i_vga.hsync ;
 wire \i_vga.timing_hor.counter[0] ;
 wire \i_vga.timing_hor.counter[10] ;
 wire \i_vga.timing_hor.counter[1] ;
 wire \i_vga.timing_hor.counter[2] ;
 wire \i_vga.timing_hor.counter[3] ;
 wire \i_vga.timing_hor.counter[4] ;
 wire \i_vga.timing_hor.counter[5] ;
 wire \i_vga.timing_hor.counter[6] ;
 wire \i_vga.timing_hor.counter[7] ;
 wire \i_vga.timing_hor.counter[8] ;
 wire \i_vga.timing_hor.counter[9] ;
 wire \i_vga.timing_ver.blank ;
 wire \i_vga.timing_ver.counter[0] ;
 wire \i_vga.timing_ver.counter[10] ;
 wire \i_vga.timing_ver.counter[1] ;
 wire \i_vga.timing_ver.counter[2] ;
 wire \i_vga.timing_ver.counter[3] ;
 wire \i_vga.timing_ver.counter[4] ;
 wire \i_vga.timing_ver.counter[5] ;
 wire \i_vga.timing_ver.counter[6] ;
 wire \i_vga.timing_ver.counter[7] ;
 wire \i_vga.timing_ver.counter[8] ;
 wire \i_vga.timing_ver.counter[9] ;
 wire \i_vga.timing_ver.sync ;
 wire \i_vga.vblank ;
 wire \i_video.colour[0] ;
 wire \i_video.colour[1] ;
 wire \i_video.colour[2] ;
 wire \i_video.colour[3] ;
 wire \i_video.colour[4] ;
 wire \i_video.colour[5] ;
 wire \i_video.frame_counter ;
 wire \i_video.read_next_r ;
 wire \i_video.repeat_count[0] ;
 wire \i_video.repeat_count[1] ;
 wire \i_video.repeat_count[2] ;
 wire \i_video.repeat_count[3] ;
 wire \i_video.repeat_count[4] ;
 wire \i_video.repeat_count[5] ;
 wire \i_video.repeat_count[6] ;
 wire \i_video.repeat_count[7] ;
 wire \i_video.repeat_count[8] ;
 wire \i_video.run_length[0] ;
 wire \i_video.run_length[1] ;
 wire \i_video.run_length[2] ;
 wire \i_video.run_length[3] ;
 wire \i_video.run_length[4] ;
 wire \i_video.run_length[5] ;
 wire \i_video.run_length[6] ;
 wire \i_video.run_length[7] ;
 wire \i_video.run_length[8] ;
 wire \i_video.run_length[9] ;
 wire \i_video.start ;
 wire spi_started;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_buf_2 _1661_ (.A(\i_spi.fsm_state[0] ),
    .X(_1015_));
 sg13g2_inv_1 _1662_ (.Y(_1016_),
    .A(_1015_));
 sg13g2_buf_1 _1663_ (.A(\i_spi.fsm_state[1] ),
    .X(_1017_));
 sg13g2_nand2_2 _1664_ (.Y(_1018_),
    .A(_1017_),
    .B(_0019_));
 sg13g2_nor2_2 _1665_ (.A(_1016_),
    .B(_1018_),
    .Y(\i_spi.spi_select ));
 sg13g2_buf_2 _1666_ (.A(_0017_),
    .X(_1019_));
 sg13g2_buf_1 _1667_ (.A(\i_vga.timing_ver.counter[1] ),
    .X(_1020_));
 sg13g2_inv_1 _1668_ (.Y(_1021_),
    .A(_1020_));
 sg13g2_inv_1 _1669_ (.Y(_1022_),
    .A(\i_vga.timing_ver.counter[4] ));
 sg13g2_nand2_1 _1670_ (.Y(_1023_),
    .A(\i_vga.timing_ver.counter[3] ),
    .B(\i_vga.timing_ver.counter[2] ));
 sg13g2_nor3_1 _1671_ (.A(_1021_),
    .B(_1022_),
    .C(_1023_),
    .Y(_1024_));
 sg13g2_inv_1 _1672_ (.Y(_1025_),
    .A(_1024_));
 sg13g2_buf_2 _1673_ (.A(\i_vga.timing_ver.counter[5] ),
    .X(_1026_));
 sg13g2_inv_1 _1674_ (.Y(_1027_),
    .A(\i_vga.timing_ver.counter[6] ));
 sg13g2_nor2_1 _1675_ (.A(_1026_),
    .B(_1027_),
    .Y(_1028_));
 sg13g2_nand2_1 _1676_ (.Y(_1029_),
    .A(_1025_),
    .B(_1028_));
 sg13g2_buf_1 _1677_ (.A(\i_vga.timing_ver.counter[10] ),
    .X(_1030_));
 sg13g2_nand2_1 _1678_ (.Y(_1031_),
    .A(\i_vga.timing_ver.counter[8] ),
    .B(\i_vga.timing_ver.counter[9] ));
 sg13g2_nand2_1 _1679_ (.Y(_1032_),
    .A(\i_vga.timing_ver.counter[7] ),
    .B(\i_vga.timing_ver.counter[6] ));
 sg13g2_nor2_1 _1680_ (.A(_1031_),
    .B(_1032_),
    .Y(_1033_));
 sg13g2_nand3_1 _1681_ (.B(_1030_),
    .C(_1033_),
    .A(_1029_),
    .Y(_1034_));
 sg13g2_xnor2_1 _1682_ (.Y(_1035_),
    .A(_1019_),
    .B(_1034_));
 sg13g2_nor3_2 _1683_ (.A(_1026_),
    .B(_1022_),
    .C(_1032_),
    .Y(_1036_));
 sg13g2_inv_1 _1684_ (.Y(_1037_),
    .A(\i_vga.timing_ver.counter[0] ));
 sg13g2_nor3_1 _1685_ (.A(_1020_),
    .B(_1037_),
    .C(_1023_),
    .Y(_1038_));
 sg13g2_nor2_1 _1686_ (.A(_1019_),
    .B(_1031_),
    .Y(_1039_));
 sg13g2_nand3_1 _1687_ (.B(_1038_),
    .C(_1039_),
    .A(_1036_),
    .Y(_1040_));
 sg13g2_inv_1 _1688_ (.Y(_1041_),
    .A(_1040_));
 sg13g2_nand3_1 _1689_ (.B(_1026_),
    .C(_1030_),
    .A(_1033_),
    .Y(_1042_));
 sg13g2_inv_1 _1690_ (.Y(_1043_),
    .A(_1031_));
 sg13g2_and3_1 _1691_ (.X(_1044_),
    .A(_1043_),
    .B(\i_vga.timing_ver.counter[0] ),
    .C(_1030_));
 sg13g2_inv_1 _1692_ (.Y(_1045_),
    .A(_1023_));
 sg13g2_nand4_1 _1693_ (.B(_1020_),
    .C(_1045_),
    .A(_1044_),
    .Y(_1046_),
    .D(_1036_));
 sg13g2_o21ai_1 _1694_ (.B1(_1046_),
    .Y(_1047_),
    .A1(_1019_),
    .A2(_1042_));
 sg13g2_a21oi_1 _1695_ (.A1(_1019_),
    .A2(_1042_),
    .Y(_1048_),
    .B1(_1047_));
 sg13g2_o21ai_1 _1696_ (.B1(_1048_),
    .Y(_0001_),
    .A1(_1035_),
    .A2(_1041_));
 sg13g2_inv_1 _1697_ (.Y(_1049_),
    .A(\i_vga.timing_hor.counter[5] ));
 sg13g2_inv_1 _1698_ (.Y(_1050_),
    .A(\i_vga.timing_hor.counter[10] ));
 sg13g2_a21oi_1 _1699_ (.A1(_1049_),
    .A2(_0014_),
    .Y(_1051_),
    .B1(_1050_));
 sg13g2_buf_2 _1700_ (.A(\i_vga.timing_hor.counter[7] ),
    .X(_1052_));
 sg13g2_nand2_1 _1701_ (.Y(_1053_),
    .A(\i_vga.timing_hor.counter[9] ),
    .B(\i_vga.timing_hor.counter[8] ));
 sg13g2_inv_1 _1702_ (.Y(_1054_),
    .A(_1053_));
 sg13g2_nand4_1 _1703_ (.B(\i_vga.timing_hor.counter[6] ),
    .C(_1052_),
    .A(_1051_),
    .Y(_1055_),
    .D(_1054_));
 sg13g2_nand2_1 _1704_ (.Y(_1056_),
    .A(\i_vga.timing_hor.counter[6] ),
    .B(_1052_));
 sg13g2_nor4_1 _1705_ (.A(\i_vga.timing_hor.counter[5] ),
    .B(_1050_),
    .C(_1053_),
    .D(_1056_),
    .Y(_1057_));
 sg13g2_inv_1 _1706_ (.Y(_1058_),
    .A(\i_vga.timing_hor.counter[0] ));
 sg13g2_and3_1 _1707_ (.X(_1059_),
    .A(\i_vga.timing_hor.counter[1] ),
    .B(\i_vga.timing_hor.counter[3] ),
    .C(\i_vga.timing_hor.counter[2] ));
 sg13g2_inv_2 _1708_ (.Y(_1060_),
    .A(_1059_));
 sg13g2_nor2_2 _1709_ (.A(_1058_),
    .B(_1060_),
    .Y(_1061_));
 sg13g2_inv_1 _1710_ (.Y(_1062_),
    .A(\i_vga.timing_hor.counter[4] ));
 sg13g2_nand3_1 _1711_ (.B(_1061_),
    .C(_1062_),
    .A(_1057_),
    .Y(_1063_));
 sg13g2_o21ai_1 _1712_ (.B1(_1063_),
    .Y(_1064_),
    .A1(_0015_),
    .A2(_1055_));
 sg13g2_nor2_1 _1713_ (.A(_0015_),
    .B(_1053_),
    .Y(_1065_));
 sg13g2_inv_2 _1714_ (.Y(_1066_),
    .A(\i_vga.timing_hor.counter[6] ));
 sg13g2_nor4_1 _1715_ (.A(\i_vga.timing_hor.counter[4] ),
    .B(_1052_),
    .C(_1049_),
    .D(_1066_),
    .Y(_1067_));
 sg13g2_nand3_1 _1716_ (.B(_1065_),
    .C(_1067_),
    .A(_1061_),
    .Y(_1068_));
 sg13g2_nor3_1 _1717_ (.A(_0014_),
    .B(_1049_),
    .C(_1066_),
    .Y(_1069_));
 sg13g2_o21ai_1 _1718_ (.B1(_1054_),
    .Y(_1070_),
    .A1(_1052_),
    .A2(_1069_));
 sg13g2_nand3_1 _1719_ (.B(\i_vga.timing_hor.counter[10] ),
    .C(_1070_),
    .A(_1068_),
    .Y(_1071_));
 sg13g2_nand2_1 _1720_ (.Y(_1072_),
    .A(_1055_),
    .B(_0015_));
 sg13g2_nand3b_1 _1721_ (.B(_1071_),
    .C(_1072_),
    .Y(_0000_),
    .A_N(_1064_));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_nor2_1 _1723_ (.A(\i_video.repeat_count[4] ),
    .B(\i_video.repeat_count[3] ),
    .Y(_1073_));
 sg13g2_nor2_1 _1724_ (.A(\i_video.repeat_count[2] ),
    .B(\i_video.repeat_count[1] ),
    .Y(_1074_));
 sg13g2_nand2_1 _1725_ (.Y(_1075_),
    .A(_1073_),
    .B(_1074_));
 sg13g2_nor2_1 _1726_ (.A(\i_video.repeat_count[7] ),
    .B(\i_video.repeat_count[8] ),
    .Y(_1076_));
 sg13g2_nor2_1 _1727_ (.A(\i_video.repeat_count[6] ),
    .B(\i_video.repeat_count[5] ),
    .Y(_1077_));
 sg13g2_nand2_1 _1728_ (.Y(_1078_),
    .A(_1076_),
    .B(_1077_));
 sg13g2_nor2_2 _1729_ (.A(_1075_),
    .B(_1078_),
    .Y(_1079_));
 sg13g2_buf_8 _1730_ (.A(\i_video.run_length[8] ),
    .X(_1080_));
 sg13g2_nand2_1 _1731_ (.Y(_1081_),
    .A(\i_video.run_length[6] ),
    .B(_1080_));
 sg13g2_buf_8 _1732_ (.A(\i_video.run_length[9] ),
    .X(_1082_));
 sg13g2_nand2_1 _1733_ (.Y(_1083_),
    .A(\i_video.run_length[7] ),
    .B(_1082_));
 sg13g2_inv_1 _1734_ (.Y(_1084_),
    .A(\i_video.run_length[4] ));
 sg13g2_nand2_1 _1735_ (.Y(_1085_),
    .A(_1084_),
    .B(\i_video.run_length[5] ));
 sg13g2_nor3_2 _1736_ (.A(_1081_),
    .B(_1083_),
    .C(_1085_),
    .Y(_1086_));
 sg13g2_inv_2 _1737_ (.Y(_1087_),
    .A(_1086_));
 sg13g2_a21oi_1 _1738_ (.A1(_1079_),
    .A2(\i_video.repeat_count[0] ),
    .Y(_1088_),
    .B1(_1087_));
 sg13g2_buf_8 _1739_ (.A(_1088_),
    .X(_1089_));
 sg13g2_nand2_1 _1740_ (.Y(_1090_),
    .A(\i_vga.timing_hor.counter[4] ),
    .B(\i_vga.timing_hor.counter[5] ));
 sg13g2_nor3_1 _1741_ (.A(_1066_),
    .B(_1052_),
    .C(_1090_),
    .Y(_1091_));
 sg13g2_inv_1 _1742_ (.Y(_1092_),
    .A(\i_vga.timing_hor.counter[9] ));
 sg13g2_nor3_1 _1743_ (.A(\i_vga.timing_hor.counter[8] ),
    .B(\i_vga.timing_hor.counter[10] ),
    .C(_1092_),
    .Y(_1093_));
 sg13g2_nand2_1 _1744_ (.Y(_1094_),
    .A(_1091_),
    .B(_1093_));
 sg13g2_inv_2 _1745_ (.Y(_1095_),
    .A(_1061_));
 sg13g2_nor2_1 _1746_ (.A(_1094_),
    .B(_1095_),
    .Y(_1096_));
 sg13g2_nand2_1 _1747_ (.Y(_1097_),
    .A(_1096_),
    .B(_1041_));
 sg13g2_nor2b_2 _1748_ (.A(_1097_),
    .B_N(_0016_),
    .Y(_1098_));
 sg13g2_nor2_2 _1749_ (.A(_1089_),
    .B(_1098_),
    .Y(_1099_));
 sg13g2_inv_1 _1750_ (.Y(_1100_),
    .A(\i_video.run_length[5] ));
 sg13g2_inv_1 _1751_ (.Y(_1101_),
    .A(\i_video.run_length[7] ));
 sg13g2_inv_1 _1752_ (.Y(_1102_),
    .A(_1082_));
 sg13g2_nor4_1 _1753_ (.A(_1100_),
    .B(_1101_),
    .C(_1102_),
    .D(_1081_),
    .Y(_1103_));
 sg13g2_inv_1 _1754_ (.Y(_1104_),
    .A(\i_video.run_length[3] ));
 sg13g2_inv_1 _1755_ (.Y(_1105_),
    .A(\i_video.run_length[2] ));
 sg13g2_buf_2 _1756_ (.A(\i_video.run_length[1] ),
    .X(_1106_));
 sg13g2_buf_1 _1757_ (.A(\i_video.run_length[0] ),
    .X(_1107_));
 sg13g2_nand2_1 _1758_ (.Y(_1108_),
    .A(_1106_),
    .B(net84));
 sg13g2_nor4_1 _1759_ (.A(_1104_),
    .B(_1105_),
    .C(_1084_),
    .D(_1108_),
    .Y(_1109_));
 sg13g2_nand2_2 _1760_ (.Y(_1110_),
    .A(_1103_),
    .B(_1109_));
 sg13g2_nand3_1 _1761_ (.B(\i_video.read_next_r ),
    .C(_1110_),
    .A(_1099_),
    .Y(_1111_));
 sg13g2_nor2b_1 _1762_ (.A(_1111_),
    .B_N(_0020_),
    .Y(_1112_));
 sg13g2_nand2_1 _1763_ (.Y(_1113_),
    .A(_1112_),
    .B(\i_spi.spi_select ));
 sg13g2_buf_1 _1764_ (.A(_1113_),
    .X(_1114_));
 sg13g2_buf_1 _1765_ (.A(_1114_),
    .X(_1115_));
 sg13g2_inv_1 _1766_ (.Y(_1116_),
    .A(\i_spi.fsm_state[2] ));
 sg13g2_nor2_1 _1767_ (.A(_1017_),
    .B(_1116_),
    .Y(_1117_));
 sg13g2_inv_1 _1768_ (.Y(_1118_),
    .A(_1117_));
 sg13g2_nor2_1 _1769_ (.A(_1016_),
    .B(_1118_),
    .Y(_1119_));
 sg13g2_buf_2 _1770_ (.A(_1119_),
    .X(_1120_));
 sg13g2_inv_1 _1771_ (.Y(_1121_),
    .A(_1120_));
 sg13g2_buf_1 _1772_ (.A(_1121_),
    .X(_1122_));
 sg13g2_inv_1 _1773_ (.Y(_1123_),
    .A(\i_spi.addr[9] ));
 sg13g2_nor2_1 _1774_ (.A(_1123_),
    .B(net54),
    .Y(_1124_));
 sg13g2_a21oi_1 _1775_ (.A1(\i_spi.addr[10] ),
    .A2(net54),
    .Y(_1125_),
    .B1(_1124_));
 sg13g2_buf_1 _1776_ (.A(_1114_),
    .X(_1126_));
 sg13g2_nor2_1 _1777_ (.A(\addr[10] ),
    .B(_1126_),
    .Y(_1127_));
 sg13g2_a21oi_1 _1778_ (.A1(_1115_),
    .A2(_1125_),
    .Y(_0093_),
    .B1(_1127_));
 sg13g2_buf_1 _1779_ (.A(_1120_),
    .X(_1128_));
 sg13g2_buf_1 _1780_ (.A(_1120_),
    .X(_1129_));
 sg13g2_nor2b_1 _1781_ (.A(net59),
    .B_N(\i_spi.addr[11] ),
    .Y(_1130_));
 sg13g2_a21oi_1 _1782_ (.A1(\i_spi.addr[10] ),
    .A2(net60),
    .Y(_1131_),
    .B1(_1130_));
 sg13g2_nor2_1 _1783_ (.A(\addr[11] ),
    .B(net40),
    .Y(_1132_));
 sg13g2_a21oi_1 _1784_ (.A1(_1115_),
    .A2(_1131_),
    .Y(_0094_),
    .B1(_1132_));
 sg13g2_nor2b_1 _1785_ (.A(net59),
    .B_N(\i_spi.addr[12] ),
    .Y(_1133_));
 sg13g2_a21oi_1 _1786_ (.A1(\i_spi.addr[11] ),
    .A2(net60),
    .Y(_1134_),
    .B1(_1133_));
 sg13g2_nor2_1 _1787_ (.A(\addr[12] ),
    .B(net40),
    .Y(_1135_));
 sg13g2_a21oi_1 _1788_ (.A1(net41),
    .A2(_1134_),
    .Y(_0095_),
    .B1(_1135_));
 sg13g2_buf_1 _1789_ (.A(_1120_),
    .X(_1136_));
 sg13g2_nor2b_1 _1790_ (.A(net58),
    .B_N(\i_spi.addr[13] ),
    .Y(_1137_));
 sg13g2_a21oi_1 _1791_ (.A1(\i_spi.addr[12] ),
    .A2(net60),
    .Y(_1138_),
    .B1(_1137_));
 sg13g2_buf_2 _1792_ (.A(\addr[13] ),
    .X(_1139_));
 sg13g2_nor2_1 _1793_ (.A(_1139_),
    .B(net40),
    .Y(_1140_));
 sg13g2_a21oi_1 _1794_ (.A1(net41),
    .A2(_1138_),
    .Y(_0096_),
    .B1(_1140_));
 sg13g2_nor2b_1 _1795_ (.A(net58),
    .B_N(\i_spi.addr[14] ),
    .Y(_1141_));
 sg13g2_a21oi_1 _1796_ (.A1(\i_spi.addr[13] ),
    .A2(net60),
    .Y(_1142_),
    .B1(_1141_));
 sg13g2_buf_2 _1797_ (.A(\addr[14] ),
    .X(_1143_));
 sg13g2_nor2_1 _1798_ (.A(_1143_),
    .B(net40),
    .Y(_1144_));
 sg13g2_a21oi_1 _1799_ (.A1(net41),
    .A2(_1142_),
    .Y(_0097_),
    .B1(_1144_));
 sg13g2_nor2b_1 _1800_ (.A(net58),
    .B_N(\i_spi.addr[15] ),
    .Y(_1145_));
 sg13g2_a21oi_1 _1801_ (.A1(\i_spi.addr[14] ),
    .A2(net60),
    .Y(_1146_),
    .B1(_1145_));
 sg13g2_nor2_1 _1802_ (.A(\addr[15] ),
    .B(net40),
    .Y(_1147_));
 sg13g2_a21oi_1 _1803_ (.A1(net41),
    .A2(_1146_),
    .Y(_0098_),
    .B1(_1147_));
 sg13g2_nor2b_1 _1804_ (.A(net58),
    .B_N(\i_spi.addr[16] ),
    .Y(_1148_));
 sg13g2_a21oi_1 _1805_ (.A1(\i_spi.addr[15] ),
    .A2(net60),
    .Y(_1149_),
    .B1(_1148_));
 sg13g2_nor2_1 _1806_ (.A(\addr[16] ),
    .B(net40),
    .Y(_1150_));
 sg13g2_a21oi_1 _1807_ (.A1(net41),
    .A2(_1149_),
    .Y(_0099_),
    .B1(_1150_));
 sg13g2_nor2b_1 _1808_ (.A(net58),
    .B_N(\i_spi.addr[17] ),
    .Y(_1151_));
 sg13g2_a21oi_1 _1809_ (.A1(\i_spi.addr[16] ),
    .A2(_1128_),
    .Y(_1152_),
    .B1(_1151_));
 sg13g2_buf_2 _1810_ (.A(\addr[17] ),
    .X(_1153_));
 sg13g2_nor2_1 _1811_ (.A(_1153_),
    .B(net40),
    .Y(_1154_));
 sg13g2_a21oi_1 _1812_ (.A1(net41),
    .A2(_1152_),
    .Y(_0100_),
    .B1(_1154_));
 sg13g2_nor2b_1 _1813_ (.A(net58),
    .B_N(\i_spi.addr[18] ),
    .Y(_1155_));
 sg13g2_a21oi_1 _1814_ (.A1(\i_spi.addr[17] ),
    .A2(_1128_),
    .Y(_1156_),
    .B1(_1155_));
 sg13g2_nor2_1 _1815_ (.A(\addr[18] ),
    .B(net40),
    .Y(_1157_));
 sg13g2_a21oi_1 _1816_ (.A1(net41),
    .A2(_1156_),
    .Y(_0101_),
    .B1(_1157_));
 sg13g2_nor2b_1 _1817_ (.A(net58),
    .B_N(\i_spi.addr[19] ),
    .Y(_1158_));
 sg13g2_a21oi_1 _1818_ (.A1(\i_spi.addr[18] ),
    .A2(net59),
    .Y(_1159_),
    .B1(_1158_));
 sg13g2_buf_1 _1819_ (.A(\addr[19] ),
    .X(_1160_));
 sg13g2_buf_1 _1820_ (.A(_1114_),
    .X(_1161_));
 sg13g2_nor2_1 _1821_ (.A(_1160_),
    .B(net39),
    .Y(_1162_));
 sg13g2_a21oi_1 _1822_ (.A1(net41),
    .A2(_1159_),
    .Y(_0102_),
    .B1(_1162_));
 sg13g2_inv_1 _1823_ (.Y(_1163_),
    .A(\i_spi.addr[1] ));
 sg13g2_nand2_1 _1824_ (.Y(_1164_),
    .A(_1114_),
    .B(net54));
 sg13g2_inv_1 _1825_ (.Y(_1165_),
    .A(_1114_));
 sg13g2_nand2_1 _1826_ (.Y(_1166_),
    .A(_1165_),
    .B(\addr[1] ));
 sg13g2_o21ai_1 _1827_ (.B1(_1166_),
    .Y(_0103_),
    .A1(_1163_),
    .A2(_1164_));
 sg13g2_buf_1 _1828_ (.A(_1114_),
    .X(_1167_));
 sg13g2_nor2b_1 _1829_ (.A(_1136_),
    .B_N(\i_spi.addr[20] ),
    .Y(_1168_));
 sg13g2_a21oi_1 _1830_ (.A1(\i_spi.addr[19] ),
    .A2(net59),
    .Y(_1169_),
    .B1(_1168_));
 sg13g2_buf_1 _1831_ (.A(\addr[20] ),
    .X(_1170_));
 sg13g2_nor2_1 _1832_ (.A(_1170_),
    .B(net39),
    .Y(_1171_));
 sg13g2_a21oi_1 _1833_ (.A1(net38),
    .A2(_1169_),
    .Y(_0104_),
    .B1(_1171_));
 sg13g2_inv_1 _1834_ (.Y(_1172_),
    .A(\i_spi.addr[21] ));
 sg13g2_nor2_1 _1835_ (.A(_1172_),
    .B(_1120_),
    .Y(_1173_));
 sg13g2_a21oi_1 _1836_ (.A1(\i_spi.addr[20] ),
    .A2(_1129_),
    .Y(_1174_),
    .B1(_1173_));
 sg13g2_buf_1 _1837_ (.A(\addr[21] ),
    .X(_1175_));
 sg13g2_nor2_1 _1838_ (.A(_1175_),
    .B(net39),
    .Y(_1176_));
 sg13g2_a21oi_1 _1839_ (.A1(net38),
    .A2(_1174_),
    .Y(_0105_),
    .B1(_1176_));
 sg13g2_nor2_1 _1840_ (.A(_1172_),
    .B(net54),
    .Y(_1177_));
 sg13g2_a21oi_1 _1841_ (.A1(\i_spi.addr[22] ),
    .A2(net54),
    .Y(_1178_),
    .B1(_1177_));
 sg13g2_nor2_1 _1842_ (.A(\addr[22] ),
    .B(net39),
    .Y(_1179_));
 sg13g2_a21oi_1 _1843_ (.A1(_1167_),
    .A2(_1178_),
    .Y(_0106_),
    .B1(_1179_));
 sg13g2_inv_1 _1844_ (.Y(_1180_),
    .A(\i_spi.addr[23] ));
 sg13g2_a22oi_1 _1845_ (.Y(_1181_),
    .B1(\addr[23] ),
    .B2(_1165_),
    .A2(net60),
    .A1(\i_spi.addr[22] ));
 sg13g2_o21ai_1 _1846_ (.B1(_1181_),
    .Y(_0107_),
    .A1(_1180_),
    .A2(_1164_));
 sg13g2_nor2_1 _1847_ (.A(_1163_),
    .B(net54),
    .Y(_1182_));
 sg13g2_a21oi_1 _1848_ (.A1(\i_spi.addr[2] ),
    .A2(net54),
    .Y(_1183_),
    .B1(_1182_));
 sg13g2_nor2_1 _1849_ (.A(\addr[2] ),
    .B(_1161_),
    .Y(_1184_));
 sg13g2_a21oi_1 _1850_ (.A1(net38),
    .A2(_1183_),
    .Y(_0108_),
    .B1(_1184_));
 sg13g2_nor2b_1 _1851_ (.A(_1136_),
    .B_N(\i_spi.addr[3] ),
    .Y(_1185_));
 sg13g2_a21oi_1 _1852_ (.A1(\i_spi.addr[2] ),
    .A2(net59),
    .Y(_1186_),
    .B1(_1185_));
 sg13g2_nor2_1 _1853_ (.A(\addr[3] ),
    .B(net39),
    .Y(_1187_));
 sg13g2_a21oi_1 _1854_ (.A1(net38),
    .A2(_1186_),
    .Y(_0109_),
    .B1(_1187_));
 sg13g2_nor2b_1 _1855_ (.A(net58),
    .B_N(\i_spi.addr[4] ),
    .Y(_1188_));
 sg13g2_a21oi_1 _1856_ (.A1(\i_spi.addr[3] ),
    .A2(net59),
    .Y(_1189_),
    .B1(_1188_));
 sg13g2_nor2_1 _1857_ (.A(\addr[4] ),
    .B(net39),
    .Y(_1190_));
 sg13g2_a21oi_1 _1858_ (.A1(net38),
    .A2(_1189_),
    .Y(_0110_),
    .B1(_1190_));
 sg13g2_nor2b_1 _1859_ (.A(_1120_),
    .B_N(\i_spi.addr[5] ),
    .Y(_1191_));
 sg13g2_a21oi_1 _1860_ (.A1(\i_spi.addr[4] ),
    .A2(net59),
    .Y(_1192_),
    .B1(_1191_));
 sg13g2_buf_2 _1861_ (.A(\addr[5] ),
    .X(_1193_));
 sg13g2_nor2_1 _1862_ (.A(_1193_),
    .B(net39),
    .Y(_1194_));
 sg13g2_a21oi_1 _1863_ (.A1(_1167_),
    .A2(_1192_),
    .Y(_0111_),
    .B1(_1194_));
 sg13g2_nor2b_1 _1864_ (.A(_1120_),
    .B_N(\i_spi.addr[6] ),
    .Y(_1195_));
 sg13g2_a21oi_1 _1865_ (.A1(\i_spi.addr[5] ),
    .A2(_1129_),
    .Y(_1196_),
    .B1(_1195_));
 sg13g2_nor2_1 _1866_ (.A(\addr[6] ),
    .B(net39),
    .Y(_1197_));
 sg13g2_a21oi_1 _1867_ (.A1(net38),
    .A2(_1196_),
    .Y(_0112_),
    .B1(_1197_));
 sg13g2_inv_1 _1868_ (.Y(_1198_),
    .A(\i_spi.addr[7] ));
 sg13g2_nor2_1 _1869_ (.A(_1198_),
    .B(_1120_),
    .Y(_1199_));
 sg13g2_a21oi_1 _1870_ (.A1(\i_spi.addr[6] ),
    .A2(net59),
    .Y(_1200_),
    .B1(_1199_));
 sg13g2_nor2_1 _1871_ (.A(\addr[7] ),
    .B(_1161_),
    .Y(_1201_));
 sg13g2_a21oi_1 _1872_ (.A1(net38),
    .A2(_1200_),
    .Y(_0113_),
    .B1(_1201_));
 sg13g2_nor2_1 _1873_ (.A(_1198_),
    .B(_1122_),
    .Y(_1202_));
 sg13g2_a21oi_1 _1874_ (.A1(\i_spi.addr[8] ),
    .A2(net54),
    .Y(_1203_),
    .B1(_1202_));
 sg13g2_nor2_1 _1875_ (.A(\addr[8] ),
    .B(_1114_),
    .Y(_1204_));
 sg13g2_a21oi_1 _1876_ (.A1(net38),
    .A2(_1203_),
    .Y(_0114_),
    .B1(_1204_));
 sg13g2_a22oi_1 _1877_ (.Y(_1205_),
    .B1(\addr[9] ),
    .B2(_1165_),
    .A2(net60),
    .A1(\i_spi.addr[8] ));
 sg13g2_o21ai_1 _1878_ (.B1(_1205_),
    .Y(_0115_),
    .A1(_1123_),
    .A2(_1164_));
 sg13g2_inv_1 _1879_ (.Y(_1206_),
    .A(\i_spi_buf.fifo[0] ));
 sg13g2_buf_1 _1880_ (.A(\i_spi_buf.empty ),
    .X(_1207_));
 sg13g2_inv_1 _1881_ (.Y(_1208_),
    .A(spi_started));
 sg13g2_nor2_2 _1882_ (.A(_1208_),
    .B(_1111_),
    .Y(_1209_));
 sg13g2_inv_1 _1883_ (.Y(_1210_),
    .A(_1209_));
 sg13g2_nor2_1 _1884_ (.A(_1207_),
    .B(_1210_),
    .Y(_1211_));
 sg13g2_inv_1 _1885_ (.Y(_1212_),
    .A(_1207_));
 sg13g2_inv_1 _1886_ (.Y(_1213_),
    .A(_1017_));
 sg13g2_nor2_1 _1887_ (.A(\i_spi.fsm_state[2] ),
    .B(_1213_),
    .Y(_1214_));
 sg13g2_buf_1 _1888_ (.A(_1214_),
    .X(_1215_));
 sg13g2_inv_1 _1889_ (.Y(_1216_),
    .A(net66));
 sg13g2_nor3_1 _1890_ (.A(_1212_),
    .B(_1216_),
    .C(_1209_),
    .Y(_1217_));
 sg13g2_buf_1 _1891_ (.A(rst_n),
    .X(_1218_));
 sg13g2_o21ai_1 _1892_ (.B1(_1218_),
    .Y(_1219_),
    .A1(_1211_),
    .A2(_1217_));
 sg13g2_buf_2 _1893_ (.A(\i_spi_buf.prev_empty ),
    .X(_1220_));
 sg13g2_inv_1 _1894_ (.Y(_1221_),
    .A(_1220_));
 sg13g2_nor2_1 _1895_ (.A(_1221_),
    .B(net66),
    .Y(_1222_));
 sg13g2_a21oi_1 _1896_ (.A1(_1211_),
    .A2(_1222_),
    .Y(_1223_),
    .B1(_1112_));
 sg13g2_nor2b_1 _1897_ (.A(_1219_),
    .B_N(_1223_),
    .Y(_1224_));
 sg13g2_buf_1 _1898_ (.A(_1224_),
    .X(_1225_));
 sg13g2_buf_1 _1899_ (.A(_1225_),
    .X(_1226_));
 sg13g2_buf_1 _1900_ (.A(_1220_),
    .X(_1227_));
 sg13g2_buf_1 _1901_ (.A(net80),
    .X(_1228_));
 sg13g2_inv_1 _1902_ (.Y(_1229_),
    .A(\i_spi.data[0] ));
 sg13g2_nor2_1 _1903_ (.A(net73),
    .B(\i_spi_buf0.fifo[0] ),
    .Y(_1230_));
 sg13g2_a21oi_1 _1904_ (.A1(net73),
    .A2(_1229_),
    .Y(_1231_),
    .B1(_1230_));
 sg13g2_nand2_1 _1905_ (.Y(_1232_),
    .A(net31),
    .B(_1231_));
 sg13g2_o21ai_1 _1906_ (.B1(_1232_),
    .Y(_0142_),
    .A1(_1206_),
    .A2(net31));
 sg13g2_inv_1 _1907_ (.Y(_1233_),
    .A(\i_spi.data[10] ));
 sg13g2_buf_1 _1908_ (.A(_1220_),
    .X(_1234_));
 sg13g2_nor2_1 _1909_ (.A(net79),
    .B(\i_spi_buf0.fifo[10] ),
    .Y(_1235_));
 sg13g2_a21oi_1 _1910_ (.A1(net80),
    .A2(_1233_),
    .Y(_1236_),
    .B1(_1235_));
 sg13g2_buf_1 _1911_ (.A(_1225_),
    .X(_1237_));
 sg13g2_mux2_1 _1912_ (.A0(\i_spi_buf.fifo[10] ),
    .A1(_1236_),
    .S(net30),
    .X(_0143_));
 sg13g2_inv_1 _1913_ (.Y(_1238_),
    .A(\i_spi.data[11] ));
 sg13g2_nor2_1 _1914_ (.A(net79),
    .B(\i_spi_buf0.fifo[11] ),
    .Y(_1239_));
 sg13g2_a21oi_1 _1915_ (.A1(net80),
    .A2(_1238_),
    .Y(_1240_),
    .B1(_1239_));
 sg13g2_mux2_1 _1916_ (.A0(\i_spi_buf.fifo[11] ),
    .A1(_1240_),
    .S(net30),
    .X(_0144_));
 sg13g2_inv_1 _1917_ (.Y(_1241_),
    .A(\i_spi.data[12] ));
 sg13g2_nor2_1 _1918_ (.A(net80),
    .B(\i_spi_buf0.fifo[12] ),
    .Y(_1242_));
 sg13g2_a21oi_1 _1919_ (.A1(_1227_),
    .A2(_1241_),
    .Y(_1243_),
    .B1(_1242_));
 sg13g2_mux2_1 _1920_ (.A0(\i_spi_buf.fifo[12] ),
    .A1(_1243_),
    .S(net30),
    .X(_0145_));
 sg13g2_inv_1 _1921_ (.Y(_1244_),
    .A(\i_spi.data[13] ));
 sg13g2_nor2_1 _1922_ (.A(net79),
    .B(\i_spi_buf0.fifo[13] ),
    .Y(_1245_));
 sg13g2_a21oi_1 _1923_ (.A1(_1227_),
    .A2(_1244_),
    .Y(_1246_),
    .B1(_1245_));
 sg13g2_mux2_1 _1924_ (.A0(\i_spi_buf.fifo[13] ),
    .A1(_1246_),
    .S(net30),
    .X(_0146_));
 sg13g2_inv_1 _1925_ (.Y(_1247_),
    .A(\i_spi.data[14] ));
 sg13g2_nor2_1 _1926_ (.A(net79),
    .B(\i_spi_buf0.fifo[14] ),
    .Y(_1248_));
 sg13g2_a21oi_1 _1927_ (.A1(net79),
    .A2(_1247_),
    .Y(_1249_),
    .B1(_1248_));
 sg13g2_mux2_1 _1928_ (.A0(\i_spi_buf.fifo[14] ),
    .A1(_1249_),
    .S(net30),
    .X(_0147_));
 sg13g2_inv_1 _1929_ (.Y(_1250_),
    .A(\i_spi.data[15] ));
 sg13g2_nor2_1 _1930_ (.A(_1220_),
    .B(\i_spi_buf0.fifo[15] ),
    .Y(_1251_));
 sg13g2_a21oi_1 _1931_ (.A1(net79),
    .A2(_1250_),
    .Y(_1252_),
    .B1(_1251_));
 sg13g2_mux2_1 _1932_ (.A0(\i_spi_buf.fifo[15] ),
    .A1(_1252_),
    .S(net30),
    .X(_0148_));
 sg13g2_inv_1 _1933_ (.Y(_1253_),
    .A(\i_spi_buf.fifo[1] ));
 sg13g2_inv_1 _1934_ (.Y(_1254_),
    .A(\i_spi.data[1] ));
 sg13g2_nor2_1 _1935_ (.A(net73),
    .B(\i_spi_buf0.fifo[1] ),
    .Y(_1255_));
 sg13g2_a21oi_1 _1936_ (.A1(_1228_),
    .A2(_1254_),
    .Y(_1256_),
    .B1(_1255_));
 sg13g2_nand2_1 _1937_ (.Y(_1257_),
    .A(_1226_),
    .B(_1256_));
 sg13g2_o21ai_1 _1938_ (.B1(_1257_),
    .Y(_0149_),
    .A1(_1253_),
    .A2(net31));
 sg13g2_inv_1 _1939_ (.Y(_1258_),
    .A(\i_spi_buf.fifo[2] ));
 sg13g2_inv_1 _1940_ (.Y(_1259_),
    .A(\i_spi.data[2] ));
 sg13g2_nor2_1 _1941_ (.A(net73),
    .B(\i_spi_buf0.fifo[2] ),
    .Y(_1260_));
 sg13g2_a21oi_1 _1942_ (.A1(net73),
    .A2(_1259_),
    .Y(_1261_),
    .B1(_1260_));
 sg13g2_nand2_1 _1943_ (.Y(_1262_),
    .A(net31),
    .B(_1261_));
 sg13g2_o21ai_1 _1944_ (.B1(_1262_),
    .Y(_0150_),
    .A1(_1258_),
    .A2(net31));
 sg13g2_inv_1 _1945_ (.Y(_1263_),
    .A(\i_spi_buf.fifo[3] ));
 sg13g2_inv_1 _1946_ (.Y(_1264_),
    .A(\i_spi.data[3] ));
 sg13g2_nor2_1 _1947_ (.A(net73),
    .B(\i_spi_buf0.fifo[3] ),
    .Y(_1265_));
 sg13g2_a21oi_1 _1948_ (.A1(net73),
    .A2(_1264_),
    .Y(_1266_),
    .B1(_1265_));
 sg13g2_nand2_1 _1949_ (.Y(_1267_),
    .A(net31),
    .B(_1266_));
 sg13g2_o21ai_1 _1950_ (.B1(_1267_),
    .Y(_0151_),
    .A1(_1263_),
    .A2(net31));
 sg13g2_inv_1 _1951_ (.Y(_1268_),
    .A(\i_spi_buf.fifo[4] ));
 sg13g2_inv_1 _1952_ (.Y(_1269_),
    .A(\i_spi.data[4] ));
 sg13g2_nor2_1 _1953_ (.A(net80),
    .B(\i_spi_buf0.fifo[4] ),
    .Y(_1270_));
 sg13g2_a21oi_1 _1954_ (.A1(_1228_),
    .A2(_1269_),
    .Y(_1271_),
    .B1(_1270_));
 sg13g2_nand2_1 _1955_ (.Y(_1272_),
    .A(net30),
    .B(_1271_));
 sg13g2_o21ai_1 _1956_ (.B1(_1272_),
    .Y(_0152_),
    .A1(_1268_),
    .A2(_1226_));
 sg13g2_inv_1 _1957_ (.Y(_1273_),
    .A(\i_spi_buf.fifo[5] ));
 sg13g2_inv_1 _1958_ (.Y(_1274_),
    .A(\i_spi.data[5] ));
 sg13g2_nor2_1 _1959_ (.A(net80),
    .B(\i_spi_buf0.fifo[5] ),
    .Y(_1275_));
 sg13g2_a21oi_1 _1960_ (.A1(net73),
    .A2(_1274_),
    .Y(_1276_),
    .B1(_1275_));
 sg13g2_nand2_1 _1961_ (.Y(_1277_),
    .A(net30),
    .B(_1276_));
 sg13g2_o21ai_1 _1962_ (.B1(_1277_),
    .Y(_0153_),
    .A1(_1273_),
    .A2(net31));
 sg13g2_inv_1 _1963_ (.Y(_1278_),
    .A(\i_spi.data[6] ));
 sg13g2_nor2_1 _1964_ (.A(_1220_),
    .B(\i_spi_buf0.fifo[6] ),
    .Y(_1279_));
 sg13g2_a21oi_1 _1965_ (.A1(net79),
    .A2(_1278_),
    .Y(_1280_),
    .B1(_1279_));
 sg13g2_mux2_1 _1966_ (.A0(\i_spi_buf.fifo[6] ),
    .A1(_1280_),
    .S(_1237_),
    .X(_0154_));
 sg13g2_inv_1 _1967_ (.Y(_1281_),
    .A(\i_spi.data[7] ));
 sg13g2_nor2_1 _1968_ (.A(_1220_),
    .B(\i_spi_buf0.fifo[7] ),
    .Y(_1282_));
 sg13g2_a21oi_1 _1969_ (.A1(net79),
    .A2(_1281_),
    .Y(_1283_),
    .B1(_1282_));
 sg13g2_mux2_1 _1970_ (.A0(\i_spi_buf.fifo[7] ),
    .A1(_1283_),
    .S(_1237_),
    .X(_0155_));
 sg13g2_inv_1 _1971_ (.Y(_1284_),
    .A(\i_spi.data[8] ));
 sg13g2_nor2_1 _1972_ (.A(_1220_),
    .B(\i_spi_buf0.fifo[8] ),
    .Y(_1285_));
 sg13g2_a21oi_1 _1973_ (.A1(_1234_),
    .A2(_1284_),
    .Y(_1286_),
    .B1(_1285_));
 sg13g2_mux2_1 _1974_ (.A0(\i_spi_buf.fifo[8] ),
    .A1(_1286_),
    .S(_1225_),
    .X(_0156_));
 sg13g2_inv_1 _1975_ (.Y(_1287_),
    .A(\i_spi.data[9] ));
 sg13g2_nor2_1 _1976_ (.A(_1220_),
    .B(\i_spi_buf0.fifo[9] ),
    .Y(_1288_));
 sg13g2_a21oi_1 _1977_ (.A1(_1234_),
    .A2(_1287_),
    .Y(_1289_),
    .B1(_1288_));
 sg13g2_mux2_1 _1978_ (.A0(\i_spi_buf.fifo[9] ),
    .A1(_1289_),
    .S(_1225_),
    .X(_0157_));
 sg13g2_nand2_1 _1979_ (.Y(_1290_),
    .A(_1210_),
    .B(_1212_));
 sg13g2_a21oi_1 _1980_ (.A1(_1290_),
    .A2(net80),
    .Y(_1291_),
    .B1(_1112_));
 sg13g2_nor2_1 _1981_ (.A(net80),
    .B(_1290_),
    .Y(_1292_));
 sg13g2_inv_1 _1982_ (.Y(_1293_),
    .A(_1292_));
 sg13g2_nand4_1 _1983_ (.B(_1218_),
    .C(net66),
    .A(_1291_),
    .Y(_1294_),
    .D(_1293_));
 sg13g2_buf_1 _1984_ (.A(_1294_),
    .X(_1295_));
 sg13g2_buf_1 _1985_ (.A(_1295_),
    .X(_1296_));
 sg13g2_buf_1 _1986_ (.A(_1295_),
    .X(_1297_));
 sg13g2_nand2_1 _1987_ (.Y(_1298_),
    .A(_1297_),
    .B(\i_spi_buf0.fifo[0] ));
 sg13g2_o21ai_1 _1988_ (.B1(_1298_),
    .Y(_0159_),
    .A1(_1229_),
    .A2(net27));
 sg13g2_nand2_1 _1989_ (.Y(_1299_),
    .A(net26),
    .B(\i_spi_buf0.fifo[10] ));
 sg13g2_o21ai_1 _1990_ (.B1(_1299_),
    .Y(_0160_),
    .A1(_1233_),
    .A2(net27));
 sg13g2_nand2_1 _1991_ (.Y(_1300_),
    .A(net26),
    .B(\i_spi_buf0.fifo[11] ));
 sg13g2_o21ai_1 _1992_ (.B1(_1300_),
    .Y(_0161_),
    .A1(_1238_),
    .A2(net27));
 sg13g2_nand2_1 _1993_ (.Y(_1301_),
    .A(net26),
    .B(\i_spi_buf0.fifo[12] ));
 sg13g2_o21ai_1 _1994_ (.B1(_1301_),
    .Y(_0162_),
    .A1(_1241_),
    .A2(net27));
 sg13g2_buf_1 _1995_ (.A(_1295_),
    .X(_1302_));
 sg13g2_nand2_1 _1996_ (.Y(_1303_),
    .A(net25),
    .B(\i_spi_buf0.fifo[13] ));
 sg13g2_o21ai_1 _1997_ (.B1(_1303_),
    .Y(_0163_),
    .A1(_1244_),
    .A2(net27));
 sg13g2_nand2_1 _1998_ (.Y(_1304_),
    .A(net25),
    .B(\i_spi_buf0.fifo[14] ));
 sg13g2_o21ai_1 _1999_ (.B1(_1304_),
    .Y(_0164_),
    .A1(_1247_),
    .A2(net27));
 sg13g2_nand2_1 _2000_ (.Y(_1305_),
    .A(net25),
    .B(\i_spi_buf0.fifo[15] ));
 sg13g2_o21ai_1 _2001_ (.B1(_1305_),
    .Y(_0165_),
    .A1(_1250_),
    .A2(net27));
 sg13g2_nand2_1 _2002_ (.Y(_1306_),
    .A(net25),
    .B(\i_spi_buf0.fifo[1] ));
 sg13g2_o21ai_1 _2003_ (.B1(_1306_),
    .Y(_0166_),
    .A1(_1254_),
    .A2(net27));
 sg13g2_nand2_1 _2004_ (.Y(_1307_),
    .A(net25),
    .B(\i_spi_buf0.fifo[2] ));
 sg13g2_o21ai_1 _2005_ (.B1(_1307_),
    .Y(_0167_),
    .A1(_1259_),
    .A2(_1296_));
 sg13g2_nand2_1 _2006_ (.Y(_1308_),
    .A(net25),
    .B(\i_spi_buf0.fifo[3] ));
 sg13g2_o21ai_1 _2007_ (.B1(_1308_),
    .Y(_0168_),
    .A1(_1264_),
    .A2(_1296_));
 sg13g2_nand2_1 _2008_ (.Y(_1309_),
    .A(_1302_),
    .B(\i_spi_buf0.fifo[4] ));
 sg13g2_o21ai_1 _2009_ (.B1(_1309_),
    .Y(_0169_),
    .A1(_1269_),
    .A2(_1297_));
 sg13g2_nand2_1 _2010_ (.Y(_1310_),
    .A(net25),
    .B(\i_spi_buf0.fifo[5] ));
 sg13g2_o21ai_1 _2011_ (.B1(_1310_),
    .Y(_0170_),
    .A1(_1274_),
    .A2(net26));
 sg13g2_nand2_1 _2012_ (.Y(_1311_),
    .A(_1302_),
    .B(\i_spi_buf0.fifo[6] ));
 sg13g2_o21ai_1 _2013_ (.B1(_1311_),
    .Y(_0171_),
    .A1(_1278_),
    .A2(net26));
 sg13g2_nand2_1 _2014_ (.Y(_1312_),
    .A(net25),
    .B(\i_spi_buf0.fifo[7] ));
 sg13g2_o21ai_1 _2015_ (.B1(_1312_),
    .Y(_0172_),
    .A1(_1281_),
    .A2(net26));
 sg13g2_nand2_1 _2016_ (.Y(_1313_),
    .A(_1295_),
    .B(\i_spi_buf0.fifo[8] ));
 sg13g2_o21ai_1 _2017_ (.B1(_1313_),
    .Y(_0173_),
    .A1(_1284_),
    .A2(net26));
 sg13g2_nand2_1 _2018_ (.Y(_1314_),
    .A(_1295_),
    .B(\i_spi_buf0.fifo[9] ));
 sg13g2_o21ai_1 _2019_ (.B1(_1314_),
    .Y(_0174_),
    .A1(_1287_),
    .A2(net26));
 sg13g2_buf_1 _2020_ (.A(net66),
    .X(_1315_));
 sg13g2_inv_1 _2021_ (.Y(_1316_),
    .A(net2));
 sg13g2_nand2_1 _2022_ (.Y(_1317_),
    .A(_1316_),
    .B(\i_spi.spi_miso_buf_n[4] ));
 sg13g2_nand2_1 _2023_ (.Y(_1318_),
    .A(\i_spi.spi_miso_buf_n[0] ),
    .B(net2));
 sg13g2_buf_2 _2024_ (.A(ui_in[0]),
    .X(_1319_));
 sg13g2_a21o_1 _2025_ (.A2(_1318_),
    .A1(_1317_),
    .B1(_1319_),
    .X(_1320_));
 sg13g2_mux2_1 _2026_ (.A0(\i_spi.spi_miso_buf_p[4] ),
    .A1(\i_spi.spi_miso_buf_p[0] ),
    .S(net1),
    .X(_1321_));
 sg13g2_buf_1 _2027_ (.A(net66),
    .X(_1322_));
 sg13g2_a21oi_1 _2028_ (.A1(_1321_),
    .A2(_1319_),
    .Y(_1323_),
    .B1(net63));
 sg13g2_a22oi_1 _2029_ (.Y(_0121_),
    .B1(_1320_),
    .B2(_1323_),
    .A2(net64),
    .A1(_1229_));
 sg13g2_buf_1 _2030_ (.A(net66),
    .X(_1324_));
 sg13g2_nor2_1 _2031_ (.A(\i_spi.data[6] ),
    .B(net64),
    .Y(_1325_));
 sg13g2_a21oi_1 _2032_ (.A1(_1233_),
    .A2(net62),
    .Y(_0122_),
    .B1(_1325_));
 sg13g2_nor2_1 _2033_ (.A(\i_spi.data[7] ),
    .B(net64),
    .Y(_1326_));
 sg13g2_a21oi_1 _2034_ (.A1(_1238_),
    .A2(net62),
    .Y(_0123_),
    .B1(_1326_));
 sg13g2_nor2_1 _2035_ (.A(\i_spi.data[8] ),
    .B(net64),
    .Y(_1327_));
 sg13g2_a21oi_1 _2036_ (.A1(_1241_),
    .A2(net62),
    .Y(_0124_),
    .B1(_1327_));
 sg13g2_nor2_1 _2037_ (.A(\i_spi.data[9] ),
    .B(net64),
    .Y(_1328_));
 sg13g2_a21oi_1 _2038_ (.A1(_1244_),
    .A2(net62),
    .Y(_0125_),
    .B1(_1328_));
 sg13g2_nor2_1 _2039_ (.A(\i_spi.data[10] ),
    .B(net63),
    .Y(_1329_));
 sg13g2_a21oi_1 _2040_ (.A1(_1247_),
    .A2(net62),
    .Y(_0126_),
    .B1(_1329_));
 sg13g2_nor2_1 _2041_ (.A(\i_spi.data[11] ),
    .B(net63),
    .Y(_1330_));
 sg13g2_a21oi_1 _2042_ (.A1(_1250_),
    .A2(net62),
    .Y(_0127_),
    .B1(_1330_));
 sg13g2_nand2_1 _2043_ (.Y(_1331_),
    .A(_1316_),
    .B(\i_spi.spi_miso_buf_n[5] ));
 sg13g2_nand2_1 _2044_ (.Y(_1332_),
    .A(net2),
    .B(\i_spi.spi_miso_buf_n[1] ));
 sg13g2_a21o_1 _2045_ (.A2(_1332_),
    .A1(_1331_),
    .B1(_1319_),
    .X(_1333_));
 sg13g2_mux2_1 _2046_ (.A0(\i_spi.spi_miso_buf_p[5] ),
    .A1(\i_spi.spi_miso_buf_p[1] ),
    .S(net1),
    .X(_1334_));
 sg13g2_a21oi_1 _2047_ (.A1(_1334_),
    .A2(_1319_),
    .Y(_1335_),
    .B1(_1322_));
 sg13g2_a22oi_1 _2048_ (.Y(_0128_),
    .B1(_1333_),
    .B2(_1335_),
    .A2(net64),
    .A1(_1254_));
 sg13g2_nand2_1 _2049_ (.Y(_1336_),
    .A(_1316_),
    .B(\i_spi.spi_miso_buf_n[6] ));
 sg13g2_nand2_1 _2050_ (.Y(_1337_),
    .A(net2),
    .B(\i_spi.spi_miso_buf_n[2] ));
 sg13g2_a21o_1 _2051_ (.A2(_1337_),
    .A1(_1336_),
    .B1(_1319_),
    .X(_1338_));
 sg13g2_mux2_1 _2052_ (.A0(\i_spi.spi_miso_buf_p[6] ),
    .A1(\i_spi.spi_miso_buf_p[2] ),
    .S(net1),
    .X(_1339_));
 sg13g2_a21oi_1 _2053_ (.A1(_1339_),
    .A2(_1319_),
    .Y(_1340_),
    .B1(net66));
 sg13g2_a22oi_1 _2054_ (.Y(_0129_),
    .B1(_1338_),
    .B2(_1340_),
    .A2(_1315_),
    .A1(_1259_));
 sg13g2_nand2_1 _2055_ (.Y(_1341_),
    .A(_1316_),
    .B(\i_spi.spi_miso_buf_n[7] ));
 sg13g2_nand2_1 _2056_ (.Y(_1342_),
    .A(net2),
    .B(\i_spi.spi_miso_buf_n[3] ));
 sg13g2_a21o_1 _2057_ (.A2(_1342_),
    .A1(_1341_),
    .B1(_1319_),
    .X(_1343_));
 sg13g2_mux2_1 _2058_ (.A0(\i_spi.spi_miso_buf_p[7] ),
    .A1(\i_spi.spi_miso_buf_p[3] ),
    .S(net1),
    .X(_1344_));
 sg13g2_a21oi_1 _2059_ (.A1(_1344_),
    .A2(_1319_),
    .Y(_1345_),
    .B1(_1215_));
 sg13g2_a22oi_1 _2060_ (.Y(_0130_),
    .B1(_1343_),
    .B2(_1345_),
    .A2(_1315_),
    .A1(_1264_));
 sg13g2_nor2_1 _2061_ (.A(\i_spi.data[0] ),
    .B(net63),
    .Y(_1346_));
 sg13g2_a21oi_1 _2062_ (.A1(_1269_),
    .A2(_1324_),
    .Y(_0131_),
    .B1(_1346_));
 sg13g2_nor2_1 _2063_ (.A(\i_spi.data[1] ),
    .B(net63),
    .Y(_1347_));
 sg13g2_a21oi_1 _2064_ (.A1(_1274_),
    .A2(net62),
    .Y(_0132_),
    .B1(_1347_));
 sg13g2_nor2_1 _2065_ (.A(\i_spi.data[2] ),
    .B(net63),
    .Y(_1348_));
 sg13g2_a21oi_1 _2066_ (.A1(_1278_),
    .A2(_1324_),
    .Y(_0133_),
    .B1(_1348_));
 sg13g2_nor2_1 _2067_ (.A(\i_spi.data[3] ),
    .B(net63),
    .Y(_1349_));
 sg13g2_a21oi_1 _2068_ (.A1(_1281_),
    .A2(net62),
    .Y(_0134_),
    .B1(_1349_));
 sg13g2_nor2_1 _2069_ (.A(\i_spi.data[4] ),
    .B(net63),
    .Y(_1350_));
 sg13g2_a21oi_1 _2070_ (.A1(_1284_),
    .A2(net64),
    .Y(_0135_),
    .B1(_1350_));
 sg13g2_nor2_1 _2071_ (.A(\i_spi.data[5] ),
    .B(_1322_),
    .Y(_1351_));
 sg13g2_a21oi_1 _2072_ (.A1(_1287_),
    .A2(net64),
    .Y(_0136_),
    .B1(_1351_));
 sg13g2_inv_1 _2073_ (.Y(_1352_),
    .A(_1218_));
 sg13g2_nor2_1 _2074_ (.A(clear_addr),
    .B(_1352_),
    .Y(_1353_));
 sg13g2_inv_1 _2075_ (.Y(_1354_),
    .A(_1353_));
 sg13g2_buf_1 _2076_ (.A(net72),
    .X(_1355_));
 sg13g2_nand2_2 _2077_ (.Y(_1356_),
    .A(_1210_),
    .B(_1099_));
 sg13g2_inv_1 _2078_ (.Y(_1357_),
    .A(_1356_));
 sg13g2_buf_1 _2079_ (.A(_1357_),
    .X(_1358_));
 sg13g2_nand2_2 _2080_ (.Y(_1359_),
    .A(_1079_),
    .B(\i_video.repeat_count[0] ));
 sg13g2_nand2_2 _2081_ (.Y(_1360_),
    .A(_1359_),
    .B(_1086_));
 sg13g2_buf_8 _2082_ (.A(_1360_),
    .X(_1361_));
 sg13g2_buf_8 _2083_ (.A(net57),
    .X(_1362_));
 sg13g2_buf_1 _2084_ (.A(net53),
    .X(_1363_));
 sg13g2_nor3_1 _2085_ (.A(\addr_offset1[1] ),
    .B(_0037_),
    .C(net50),
    .Y(_1364_));
 sg13g2_o21ai_1 _2086_ (.B1(_0037_),
    .Y(_1365_),
    .A1(\addr_offset1[1] ),
    .A2(_1360_));
 sg13g2_inv_1 _2087_ (.Y(_1366_),
    .A(_1365_));
 sg13g2_nor3_1 _2088_ (.A(_1020_),
    .B(_1019_),
    .C(_1037_),
    .Y(_1367_));
 sg13g2_nand4_1 _2089_ (.B(_1043_),
    .C(_1045_),
    .A(_1036_),
    .Y(_1368_),
    .D(_1367_));
 sg13g2_inv_1 _2090_ (.Y(_1369_),
    .A(_1096_));
 sg13g2_nor2_1 _2091_ (.A(_1368_),
    .B(_1369_),
    .Y(_1370_));
 sg13g2_nand2_1 _2092_ (.Y(_1371_),
    .A(_1370_),
    .B(_0016_));
 sg13g2_buf_1 _2093_ (.A(_1371_),
    .X(_1372_));
 sg13g2_o21ai_1 _2094_ (.B1(net49),
    .Y(_1373_),
    .A1(_1364_),
    .A2(_1366_));
 sg13g2_nand2_1 _2095_ (.Y(_1374_),
    .A(_1098_),
    .B(\addr_saved0[1] ));
 sg13g2_a21oi_1 _2096_ (.A1(_1373_),
    .A2(_1374_),
    .Y(_1375_),
    .B1(_1357_));
 sg13g2_a21oi_1 _2097_ (.A1(\addr[1] ),
    .A2(net34),
    .Y(_1376_),
    .B1(_1375_));
 sg13g2_nor2_1 _2098_ (.A(net65),
    .B(_1376_),
    .Y(_0039_));
 sg13g2_xnor2_1 _2099_ (.Y(_1377_),
    .A(_0026_),
    .B(net53));
 sg13g2_nor2_1 _2100_ (.A(\addr_offset1[5] ),
    .B(_1360_),
    .Y(_1378_));
 sg13g2_nand2_1 _2101_ (.Y(_1379_),
    .A(_1378_),
    .B(_1193_));
 sg13g2_inv_1 _2102_ (.Y(_1380_),
    .A(\addr_offset1[6] ));
 sg13g2_nand3_1 _2103_ (.B(_1380_),
    .C(\addr[6] ),
    .A(_1089_),
    .Y(_1381_));
 sg13g2_inv_1 _2104_ (.Y(_1382_),
    .A(\addr[6] ));
 sg13g2_o21ai_1 _2105_ (.B1(_1382_),
    .Y(_1383_),
    .A1(\addr_offset1[6] ),
    .A2(net57));
 sg13g2_inv_1 _2106_ (.Y(_1384_),
    .A(_1383_));
 sg13g2_a21oi_1 _2107_ (.A1(_1379_),
    .A2(_1381_),
    .Y(_1385_),
    .B1(_1384_));
 sg13g2_inv_1 _2108_ (.Y(_1386_),
    .A(\addr_offset1[5] ));
 sg13g2_nand2_1 _2109_ (.Y(_1387_),
    .A(_1089_),
    .B(_1386_));
 sg13g2_inv_1 _2110_ (.Y(_1388_),
    .A(_1193_));
 sg13g2_nand2_1 _2111_ (.Y(_1389_),
    .A(_1387_),
    .B(_1388_));
 sg13g2_nand2_1 _2112_ (.Y(_1390_),
    .A(_1379_),
    .B(_1389_));
 sg13g2_nand2_1 _2113_ (.Y(_1391_),
    .A(_1383_),
    .B(_1381_));
 sg13g2_nor2_1 _2114_ (.A(_1390_),
    .B(_1391_),
    .Y(_1392_));
 sg13g2_inv_1 _2115_ (.Y(_1393_),
    .A(\addr[3] ));
 sg13g2_inv_1 _2116_ (.Y(_1394_),
    .A(\addr_offset1[3] ));
 sg13g2_nand3_1 _2117_ (.B(_1394_),
    .C(_1086_),
    .A(_1359_),
    .Y(_1395_));
 sg13g2_nor2_1 _2118_ (.A(_1393_),
    .B(_1395_),
    .Y(_1396_));
 sg13g2_inv_1 _2119_ (.Y(_1397_),
    .A(_1396_));
 sg13g2_inv_1 _2120_ (.Y(_1398_),
    .A(\addr_offset1[4] ));
 sg13g2_nand3_1 _2121_ (.B(_1398_),
    .C(\addr[4] ),
    .A(_1089_),
    .Y(_1399_));
 sg13g2_nand2_1 _2122_ (.Y(_1400_),
    .A(_1089_),
    .B(_1398_));
 sg13g2_inv_1 _2123_ (.Y(_1401_),
    .A(\addr[4] ));
 sg13g2_nand2_1 _2124_ (.Y(_1402_),
    .A(_1400_),
    .B(_1401_));
 sg13g2_inv_1 _2125_ (.Y(_1403_),
    .A(_1402_));
 sg13g2_a21oi_1 _2126_ (.A1(_1397_),
    .A2(_1399_),
    .Y(_1404_),
    .B1(_1403_));
 sg13g2_nand2_1 _2127_ (.Y(_1405_),
    .A(_1392_),
    .B(_1404_));
 sg13g2_nand2b_1 _2128_ (.Y(_1406_),
    .B(_1405_),
    .A_N(_1385_));
 sg13g2_nand2_1 _2129_ (.Y(_1407_),
    .A(_1402_),
    .B(_1399_));
 sg13g2_nand2_1 _2130_ (.Y(_1408_),
    .A(_1395_),
    .B(_1393_));
 sg13g2_nand2_1 _2131_ (.Y(_1409_),
    .A(_1397_),
    .B(_1408_));
 sg13g2_nor2_1 _2132_ (.A(_1407_),
    .B(_1409_),
    .Y(_1410_));
 sg13g2_and2_1 _2133_ (.A(_1392_),
    .B(_1410_),
    .X(_1411_));
 sg13g2_inv_1 _2134_ (.Y(_1412_),
    .A(\addr[2] ));
 sg13g2_o21ai_1 _2135_ (.B1(_1412_),
    .Y(_1413_),
    .A1(\addr_offset1[2] ),
    .A2(_1361_));
 sg13g2_nor3_1 _2136_ (.A(\addr_offset1[2] ),
    .B(_1412_),
    .C(_1360_),
    .Y(_1414_));
 sg13g2_a21oi_1 _2137_ (.A1(_1365_),
    .A2(_1413_),
    .Y(_1415_),
    .B1(_1414_));
 sg13g2_inv_1 _2138_ (.Y(_1416_),
    .A(_1415_));
 sg13g2_nand2_1 _2139_ (.Y(_1417_),
    .A(_1411_),
    .B(_1416_));
 sg13g2_nand2b_1 _2140_ (.Y(_1418_),
    .B(_1417_),
    .A_N(_1406_));
 sg13g2_inv_1 _2141_ (.Y(_1419_),
    .A(\addr[8] ));
 sg13g2_o21ai_1 _2142_ (.B1(_1419_),
    .Y(_1420_),
    .A1(\addr_offset1[8] ),
    .A2(_1361_));
 sg13g2_nor3_1 _2143_ (.A(\addr_offset1[8] ),
    .B(_1419_),
    .C(_1360_),
    .Y(_1421_));
 sg13g2_inv_1 _2144_ (.Y(_1422_),
    .A(_1421_));
 sg13g2_nand2_2 _2145_ (.Y(_1423_),
    .A(_1420_),
    .B(_1422_));
 sg13g2_inv_1 _2146_ (.Y(_1424_),
    .A(\addr_offset1[7] ));
 sg13g2_nand3_1 _2147_ (.B(_1424_),
    .C(_1086_),
    .A(_1359_),
    .Y(_1425_));
 sg13g2_nand2_1 _2148_ (.Y(_1426_),
    .A(_1425_),
    .B(_0023_));
 sg13g2_inv_1 _2149_ (.Y(_1427_),
    .A(_0023_));
 sg13g2_nand4_1 _2150_ (.B(_1424_),
    .C(_1427_),
    .A(_1359_),
    .Y(_1428_),
    .D(_1086_));
 sg13g2_nand2_2 _2151_ (.Y(_1429_),
    .A(_1426_),
    .B(_1428_));
 sg13g2_xnor2_1 _2152_ (.Y(_1430_),
    .A(_0025_),
    .B(net57));
 sg13g2_xnor2_1 _2153_ (.Y(_1431_),
    .A(_0024_),
    .B(net57));
 sg13g2_nor2_1 _2154_ (.A(_1430_),
    .B(_1431_),
    .Y(_1432_));
 sg13g2_inv_1 _2155_ (.Y(_1433_),
    .A(_1432_));
 sg13g2_nor3_2 _2156_ (.A(_1423_),
    .B(_1429_),
    .C(_1433_),
    .Y(_1434_));
 sg13g2_inv_1 _2157_ (.Y(_1435_),
    .A(\addr[7] ));
 sg13g2_nor2_1 _2158_ (.A(_1435_),
    .B(_1425_),
    .Y(_1436_));
 sg13g2_nand2_1 _2159_ (.Y(_1437_),
    .A(_1420_),
    .B(_1436_));
 sg13g2_nand2_1 _2160_ (.Y(_1438_),
    .A(_1437_),
    .B(_1422_));
 sg13g2_buf_1 _2161_ (.A(_1089_),
    .X(_1439_));
 sg13g2_nand2_1 _2162_ (.Y(_1440_),
    .A(net52),
    .B(\addr[9] ));
 sg13g2_inv_1 _2163_ (.Y(_1441_),
    .A(_1440_));
 sg13g2_inv_1 _2164_ (.Y(_1442_),
    .A(\addr[10] ));
 sg13g2_nor2_1 _2165_ (.A(_1442_),
    .B(net50),
    .Y(_1443_));
 sg13g2_a21o_1 _2166_ (.A2(_0025_),
    .A1(_1441_),
    .B1(_1443_),
    .X(_1444_));
 sg13g2_a21oi_1 _2167_ (.A1(_1438_),
    .A2(_1432_),
    .Y(_1445_),
    .B1(_1444_));
 sg13g2_inv_1 _2168_ (.Y(_1446_),
    .A(_1445_));
 sg13g2_a21oi_1 _2169_ (.A1(_1418_),
    .A2(_1434_),
    .Y(_1447_),
    .B1(_1446_));
 sg13g2_xor2_1 _2170_ (.B(_1447_),
    .A(_1377_),
    .X(_1448_));
 sg13g2_buf_1 _2171_ (.A(_1371_),
    .X(_1449_));
 sg13g2_nand2_1 _2172_ (.Y(_1450_),
    .A(_1448_),
    .B(net48));
 sg13g2_inv_1 _2173_ (.Y(_1451_),
    .A(_1371_));
 sg13g2_buf_1 _2174_ (.A(net47),
    .X(_1452_));
 sg13g2_a21oi_1 _2175_ (.A1(\addr_saved0[11] ),
    .A2(net45),
    .Y(_1453_),
    .B1(net34));
 sg13g2_buf_1 _2176_ (.A(_1356_),
    .X(_1454_));
 sg13g2_buf_1 _2177_ (.A(_1353_),
    .X(_1455_));
 sg13g2_o21ai_1 _2178_ (.B1(net71),
    .Y(_1456_),
    .A1(\addr[11] ),
    .A2(net37));
 sg13g2_a21oi_1 _2179_ (.A1(_1450_),
    .A2(_1453_),
    .Y(_0040_),
    .B1(_1456_));
 sg13g2_xnor2_1 _2180_ (.Y(_1457_),
    .A(_0027_),
    .B(net53));
 sg13g2_inv_1 _2181_ (.Y(_1458_),
    .A(_1457_));
 sg13g2_inv_1 _2182_ (.Y(_1459_),
    .A(_1414_));
 sg13g2_nand2_1 _2183_ (.Y(_1460_),
    .A(_1413_),
    .B(_1459_));
 sg13g2_nor2_1 _2184_ (.A(_1409_),
    .B(_1460_),
    .Y(_1461_));
 sg13g2_nand2_1 _2185_ (.Y(_1462_),
    .A(_1461_),
    .B(_1365_));
 sg13g2_a21oi_1 _2186_ (.A1(_1414_),
    .A2(_1408_),
    .Y(_1463_),
    .B1(_1396_));
 sg13g2_nand2_2 _2187_ (.Y(_1464_),
    .A(_1462_),
    .B(_1463_));
 sg13g2_nor2_1 _2188_ (.A(_1429_),
    .B(_1391_),
    .Y(_1465_));
 sg13g2_nor2_1 _2189_ (.A(_1407_),
    .B(_1390_),
    .Y(_1466_));
 sg13g2_nand2_1 _2190_ (.Y(_1467_),
    .A(_1465_),
    .B(_1466_));
 sg13g2_nor2_1 _2191_ (.A(_1431_),
    .B(_1423_),
    .Y(_1468_));
 sg13g2_nor2_1 _2192_ (.A(_1430_),
    .B(_1377_),
    .Y(_1469_));
 sg13g2_nand2_1 _2193_ (.Y(_1470_),
    .A(_1468_),
    .B(_1469_));
 sg13g2_nor2_1 _2194_ (.A(_1467_),
    .B(_1470_),
    .Y(_1471_));
 sg13g2_nor3_1 _2195_ (.A(\addr_offset1[6] ),
    .B(_1382_),
    .C(net53),
    .Y(_1472_));
 sg13g2_nand3_1 _2196_ (.B(_1426_),
    .C(_1428_),
    .A(_1472_),
    .Y(_1473_));
 sg13g2_inv_1 _2197_ (.Y(_1474_),
    .A(_1436_));
 sg13g2_nand2_1 _2198_ (.Y(_1475_),
    .A(_1473_),
    .B(_1474_));
 sg13g2_nor2_1 _2199_ (.A(_1193_),
    .B(_1378_),
    .Y(_1476_));
 sg13g2_o21ai_1 _2200_ (.B1(_1379_),
    .Y(_1477_),
    .A1(_1399_),
    .A2(_1476_));
 sg13g2_nand2_1 _2201_ (.Y(_1478_),
    .A(_1477_),
    .B(_1465_));
 sg13g2_nand2b_1 _2202_ (.Y(_1479_),
    .B(_1478_),
    .A_N(_1475_));
 sg13g2_nand2b_1 _2203_ (.Y(_1480_),
    .B(_1479_),
    .A_N(_1470_));
 sg13g2_a21oi_1 _2204_ (.A1(_1421_),
    .A2(_0024_),
    .Y(_1481_),
    .B1(_1441_));
 sg13g2_inv_1 _2205_ (.Y(_1482_),
    .A(_1481_));
 sg13g2_inv_1 _2206_ (.Y(_1483_),
    .A(\addr[11] ));
 sg13g2_nor2_1 _2207_ (.A(_1483_),
    .B(net53),
    .Y(_1484_));
 sg13g2_a21oi_1 _2208_ (.A1(_1443_),
    .A2(_0026_),
    .Y(_1485_),
    .B1(_1484_));
 sg13g2_inv_1 _2209_ (.Y(_1486_),
    .A(_1485_));
 sg13g2_a21oi_1 _2210_ (.A1(_1482_),
    .A2(_1469_),
    .Y(_1487_),
    .B1(_1486_));
 sg13g2_nand2_1 _2211_ (.Y(_0227_),
    .A(_1480_),
    .B(_1487_));
 sg13g2_a21oi_1 _2212_ (.A1(_1464_),
    .A2(_1471_),
    .Y(_0228_),
    .B1(_0227_));
 sg13g2_xnor2_1 _2213_ (.Y(_0229_),
    .A(_1458_),
    .B(_0228_));
 sg13g2_nand2_1 _2214_ (.Y(_0230_),
    .A(_0229_),
    .B(net48));
 sg13g2_a21oi_1 _2215_ (.A1(\addr_saved0[12] ),
    .A2(net45),
    .Y(_0231_),
    .B1(net34));
 sg13g2_o21ai_1 _2216_ (.B1(net71),
    .Y(_0232_),
    .A1(\addr[12] ),
    .A2(net37));
 sg13g2_a21oi_1 _2217_ (.A1(_0230_),
    .A2(_0231_),
    .Y(_0041_),
    .B1(_0232_));
 sg13g2_nand2_1 _2218_ (.Y(_0233_),
    .A(_1416_),
    .B(_1410_));
 sg13g2_nand2b_2 _2219_ (.Y(_0234_),
    .B(_0233_),
    .A_N(_1404_));
 sg13g2_nor2_1 _2220_ (.A(_1377_),
    .B(_1457_),
    .Y(_0235_));
 sg13g2_nand2_1 _2221_ (.Y(_0236_),
    .A(_1432_),
    .B(_0235_));
 sg13g2_nor2_1 _2222_ (.A(_1429_),
    .B(_1423_),
    .Y(_0237_));
 sg13g2_nand2_1 _2223_ (.Y(_0238_),
    .A(_0237_),
    .B(_1392_));
 sg13g2_nor2_1 _2224_ (.A(_0236_),
    .B(_0238_),
    .Y(_0239_));
 sg13g2_nand2_1 _2225_ (.Y(_0240_),
    .A(_0237_),
    .B(_1385_));
 sg13g2_nand2b_1 _2226_ (.Y(_0241_),
    .B(_0240_),
    .A_N(_1438_));
 sg13g2_nand2b_1 _2227_ (.Y(_0242_),
    .B(_0241_),
    .A_N(_0236_));
 sg13g2_inv_1 _2228_ (.Y(_0243_),
    .A(\addr[12] ));
 sg13g2_nor2_1 _2229_ (.A(_0243_),
    .B(net53),
    .Y(_0244_));
 sg13g2_a21oi_1 _2230_ (.A1(_1484_),
    .A2(_0027_),
    .Y(_0245_),
    .B1(_0244_));
 sg13g2_inv_1 _2231_ (.Y(_0246_),
    .A(_0245_));
 sg13g2_a21oi_1 _2232_ (.A1(_1444_),
    .A2(_0235_),
    .Y(_0247_),
    .B1(_0246_));
 sg13g2_nand2_1 _2233_ (.Y(_0248_),
    .A(_0242_),
    .B(_0247_));
 sg13g2_a21o_1 _2234_ (.A2(_0239_),
    .A1(_0234_),
    .B1(_0248_),
    .X(_0249_));
 sg13g2_inv_1 _2235_ (.Y(_0250_),
    .A(_0028_));
 sg13g2_xnor2_1 _2236_ (.Y(_0251_),
    .A(_0250_),
    .B(net57));
 sg13g2_a21oi_1 _2237_ (.A1(_0249_),
    .A2(_0251_),
    .Y(_0252_),
    .B1(_1451_));
 sg13g2_o21ai_1 _2238_ (.B1(_0252_),
    .Y(_0253_),
    .A1(_0249_),
    .A2(_0251_));
 sg13g2_a21oi_1 _2239_ (.A1(\addr_saved0[13] ),
    .A2(net45),
    .Y(_0254_),
    .B1(net34));
 sg13g2_o21ai_1 _2240_ (.B1(net71),
    .Y(_0255_),
    .A1(_1139_),
    .A2(net37));
 sg13g2_a21oi_1 _2241_ (.A1(_0253_),
    .A2(_0254_),
    .Y(_0042_),
    .B1(_0255_));
 sg13g2_xnor2_1 _2242_ (.Y(_0256_),
    .A(_0029_),
    .B(net57));
 sg13g2_inv_1 _2243_ (.Y(_0257_),
    .A(_0256_));
 sg13g2_nand2_1 _2244_ (.Y(_0258_),
    .A(_1475_),
    .B(_1468_));
 sg13g2_nand2_1 _2245_ (.Y(_0259_),
    .A(_0258_),
    .B(_1481_));
 sg13g2_nand2_1 _2246_ (.Y(_0260_),
    .A(_1458_),
    .B(_0251_));
 sg13g2_nor2b_1 _2247_ (.A(_0260_),
    .B_N(_1469_),
    .Y(_0261_));
 sg13g2_nand2_1 _2248_ (.Y(_0262_),
    .A(_0259_),
    .B(_0261_));
 sg13g2_nor2_1 _2249_ (.A(_1485_),
    .B(_0260_),
    .Y(_0263_));
 sg13g2_a22oi_1 _2250_ (.Y(_0264_),
    .B1(_0244_),
    .B2(_0251_),
    .A2(net52),
    .A1(_1139_));
 sg13g2_nor2b_1 _2251_ (.A(_0263_),
    .B_N(_0264_),
    .Y(_0265_));
 sg13g2_nand2_1 _2252_ (.Y(_0266_),
    .A(_0262_),
    .B(_0265_));
 sg13g2_and2_1 _2253_ (.A(_1468_),
    .B(_1465_),
    .X(_0267_));
 sg13g2_nand2_1 _2254_ (.Y(_0268_),
    .A(_0267_),
    .B(_0261_));
 sg13g2_xnor2_1 _2255_ (.Y(_0269_),
    .A(_1193_),
    .B(_1387_));
 sg13g2_xnor2_1 _2256_ (.Y(_0270_),
    .A(\addr[4] ),
    .B(_1400_));
 sg13g2_nand2_1 _2257_ (.Y(_0271_),
    .A(_0269_),
    .B(_0270_));
 sg13g2_nor2_1 _2258_ (.A(_1463_),
    .B(_0271_),
    .Y(_0272_));
 sg13g2_nor2_1 _2259_ (.A(_1477_),
    .B(_0272_),
    .Y(_0273_));
 sg13g2_nand3_1 _2260_ (.B(_1466_),
    .C(_1365_),
    .A(_1461_),
    .Y(_0274_));
 sg13g2_nand2_1 _2261_ (.Y(_0275_),
    .A(_0273_),
    .B(_0274_));
 sg13g2_inv_1 _2262_ (.Y(_0276_),
    .A(_0275_));
 sg13g2_nor2_1 _2263_ (.A(_0268_),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_nor2_1 _2264_ (.A(_0266_),
    .B(_0277_),
    .Y(_0278_));
 sg13g2_xnor2_1 _2265_ (.Y(_0279_),
    .A(_0257_),
    .B(_0278_));
 sg13g2_inv_1 _2266_ (.Y(_0280_),
    .A(_1098_));
 sg13g2_nand2_1 _2267_ (.Y(_0281_),
    .A(_0279_),
    .B(_0280_));
 sg13g2_buf_1 _2268_ (.A(_1357_),
    .X(_0282_));
 sg13g2_a21oi_1 _2269_ (.A1(\addr_saved0[14] ),
    .A2(net45),
    .Y(_0283_),
    .B1(net33));
 sg13g2_o21ai_1 _2270_ (.B1(_1455_),
    .Y(_0284_),
    .A1(_1143_),
    .A2(net37));
 sg13g2_a21oi_1 _2271_ (.A1(_0281_),
    .A2(_0283_),
    .Y(_0043_),
    .B1(_0284_));
 sg13g2_nand2_1 _2272_ (.Y(_0285_),
    .A(_0257_),
    .B(_0251_));
 sg13g2_inv_1 _2273_ (.Y(_0286_),
    .A(_0285_));
 sg13g2_nand2_1 _2274_ (.Y(_0287_),
    .A(_0286_),
    .B(_0235_));
 sg13g2_inv_1 _2275_ (.Y(_0288_),
    .A(_0029_));
 sg13g2_nor2_1 _2276_ (.A(_0288_),
    .B(net50),
    .Y(_0289_));
 sg13g2_a22oi_1 _2277_ (.Y(_0290_),
    .B1(_1139_),
    .B2(_0289_),
    .A2(_1143_),
    .A1(net52));
 sg13g2_inv_1 _2278_ (.Y(_0291_),
    .A(_0290_));
 sg13g2_a21oi_1 _2279_ (.A1(_0286_),
    .A2(_0246_),
    .Y(_0292_),
    .B1(_0291_));
 sg13g2_o21ai_1 _2280_ (.B1(_0292_),
    .Y(_0293_),
    .A1(_0287_),
    .A2(_1445_));
 sg13g2_nand2b_1 _2281_ (.Y(_0294_),
    .B(_1434_),
    .A_N(_0287_));
 sg13g2_nand2b_1 _2282_ (.Y(_0295_),
    .B(_1418_),
    .A_N(_0294_));
 sg13g2_nand2b_1 _2283_ (.Y(_0296_),
    .B(_0295_),
    .A_N(_0293_));
 sg13g2_inv_1 _2284_ (.Y(_0297_),
    .A(_0030_));
 sg13g2_nor2_1 _2285_ (.A(_0297_),
    .B(net57),
    .Y(_0298_));
 sg13g2_inv_1 _2286_ (.Y(_0299_),
    .A(_0298_));
 sg13g2_nand2_1 _2287_ (.Y(_0300_),
    .A(net57),
    .B(_0297_));
 sg13g2_nand2_1 _2288_ (.Y(_0301_),
    .A(_0299_),
    .B(_0300_));
 sg13g2_o21ai_1 _2289_ (.B1(net49),
    .Y(_0302_),
    .A1(_0301_),
    .A2(_0296_));
 sg13g2_a21o_1 _2290_ (.A2(_0301_),
    .A1(_0296_),
    .B1(_0302_),
    .X(_0303_));
 sg13g2_a21oi_1 _2291_ (.A1(\addr_saved0[15] ),
    .A2(net45),
    .Y(_0304_),
    .B1(net33));
 sg13g2_o21ai_1 _2292_ (.B1(_1455_),
    .Y(_0305_),
    .A1(\addr[15] ),
    .A2(net37));
 sg13g2_a21oi_1 _2293_ (.A1(_0303_),
    .A2(_0304_),
    .Y(_0044_),
    .B1(_0305_));
 sg13g2_o21ai_1 _2294_ (.B1(_1454_),
    .Y(_0306_),
    .A1(\addr_saved0[16] ),
    .A2(net49));
 sg13g2_inv_1 _2295_ (.Y(_0307_),
    .A(_1467_));
 sg13g2_a21o_1 _2296_ (.A2(_0307_),
    .A1(_1464_),
    .B1(_1479_),
    .X(_0308_));
 sg13g2_nand2_1 _2297_ (.Y(_0309_),
    .A(_0257_),
    .B(_0301_));
 sg13g2_inv_1 _2298_ (.Y(_0310_),
    .A(_0309_));
 sg13g2_nand2b_1 _2299_ (.Y(_0311_),
    .B(_0310_),
    .A_N(_0260_));
 sg13g2_nor2_1 _2300_ (.A(_0311_),
    .B(_1470_),
    .Y(_0312_));
 sg13g2_nand2_1 _2301_ (.Y(_0313_),
    .A(_0308_),
    .B(_0312_));
 sg13g2_nor2_1 _2302_ (.A(_0311_),
    .B(_1487_),
    .Y(_0314_));
 sg13g2_inv_1 _2303_ (.Y(_0315_),
    .A(_1139_));
 sg13g2_o21ai_1 _2304_ (.B1(_0315_),
    .Y(_0316_),
    .A1(_0250_),
    .A2(_0243_));
 sg13g2_nor2b_1 _2305_ (.A(net50),
    .B_N(_0316_),
    .Y(_0317_));
 sg13g2_inv_1 _2306_ (.Y(_0318_),
    .A(\addr[15] ));
 sg13g2_nor2_1 _2307_ (.A(_0318_),
    .B(net50),
    .Y(_0319_));
 sg13g2_a21oi_1 _2308_ (.A1(_0298_),
    .A2(_1143_),
    .Y(_0320_),
    .B1(_0319_));
 sg13g2_inv_1 _2309_ (.Y(_0321_),
    .A(_0320_));
 sg13g2_a21oi_1 _2310_ (.A1(_0310_),
    .A2(_0317_),
    .Y(_0322_),
    .B1(_0321_));
 sg13g2_nor2b_1 _2311_ (.A(_0314_),
    .B_N(_0322_),
    .Y(_0323_));
 sg13g2_nand2_1 _2312_ (.Y(_0324_),
    .A(_0313_),
    .B(_0323_));
 sg13g2_xnor2_1 _2313_ (.Y(_0325_),
    .A(_0031_),
    .B(_1089_));
 sg13g2_inv_1 _2314_ (.Y(_0326_),
    .A(_0325_));
 sg13g2_nand2_1 _2315_ (.Y(_0327_),
    .A(_0324_),
    .B(_0326_));
 sg13g2_nand3_1 _2316_ (.B(_0323_),
    .C(_0325_),
    .A(_0313_),
    .Y(_0328_));
 sg13g2_nand3_1 _2317_ (.B(_0328_),
    .C(_1449_),
    .A(_0327_),
    .Y(_0329_));
 sg13g2_nand2b_1 _2318_ (.Y(_0330_),
    .B(_0329_),
    .A_N(_0306_));
 sg13g2_buf_1 _2319_ (.A(_1357_),
    .X(_0331_));
 sg13g2_nand2_1 _2320_ (.Y(_0332_),
    .A(net32),
    .B(\addr[16] ));
 sg13g2_a21oi_1 _2321_ (.A1(_0330_),
    .A2(_0332_),
    .Y(_0045_),
    .B1(net65));
 sg13g2_o21ai_1 _2322_ (.B1(_1454_),
    .Y(_0333_),
    .A1(\addr_saved0[17] ),
    .A2(net49));
 sg13g2_xnor2_1 _2323_ (.Y(_0334_),
    .A(_0032_),
    .B(_1089_));
 sg13g2_nand2b_1 _2324_ (.Y(_0335_),
    .B(_0234_),
    .A_N(_0238_));
 sg13g2_nand2b_1 _2325_ (.Y(_0336_),
    .B(_0335_),
    .A_N(_0241_));
 sg13g2_nand2_1 _2326_ (.Y(_0337_),
    .A(_0301_),
    .B(_0325_));
 sg13g2_nand2b_1 _2327_ (.Y(_0338_),
    .B(_0286_),
    .A_N(_0337_));
 sg13g2_nor2_1 _2328_ (.A(_0236_),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_nand2_1 _2329_ (.Y(_0340_),
    .A(_0336_),
    .B(_0339_));
 sg13g2_nor2b_1 _2330_ (.A(net50),
    .B_N(\addr[16] ),
    .Y(_0341_));
 sg13g2_a21oi_1 _2331_ (.A1(_0319_),
    .A2(_0031_),
    .Y(_0342_),
    .B1(_0341_));
 sg13g2_o21ai_1 _2332_ (.B1(_0342_),
    .Y(_0343_),
    .A1(_0337_),
    .A2(_0290_));
 sg13g2_nor2_1 _2333_ (.A(_0338_),
    .B(_0247_),
    .Y(_0344_));
 sg13g2_nor2_1 _2334_ (.A(_0343_),
    .B(_0344_),
    .Y(_0345_));
 sg13g2_nand2_1 _2335_ (.Y(_0346_),
    .A(_0340_),
    .B(_0345_));
 sg13g2_xnor2_1 _2336_ (.Y(_0347_),
    .A(_0334_),
    .B(_0346_));
 sg13g2_nand2_1 _2337_ (.Y(_0348_),
    .A(_0347_),
    .B(net48));
 sg13g2_nand2b_1 _2338_ (.Y(_0349_),
    .B(_0348_),
    .A_N(_0333_));
 sg13g2_nand2_1 _2339_ (.Y(_0350_),
    .A(net32),
    .B(_1153_));
 sg13g2_a21oi_1 _2340_ (.A1(_0349_),
    .A2(_0350_),
    .Y(_0046_),
    .B1(net65));
 sg13g2_o21ai_1 _2341_ (.B1(net37),
    .Y(_0351_),
    .A1(\addr_saved0[18] ),
    .A2(net49));
 sg13g2_nand2_1 _2342_ (.Y(_0352_),
    .A(_0275_),
    .B(_0267_));
 sg13g2_nand2b_1 _2343_ (.Y(_0353_),
    .B(_0352_),
    .A_N(_0259_));
 sg13g2_nand2_1 _2344_ (.Y(_0354_),
    .A(_0325_),
    .B(_0334_));
 sg13g2_nor2_1 _2345_ (.A(_0354_),
    .B(_0309_),
    .Y(_0355_));
 sg13g2_inv_1 _2346_ (.Y(_0356_),
    .A(_0355_));
 sg13g2_nor2b_1 _2347_ (.A(_0356_),
    .B_N(_0261_),
    .Y(_0357_));
 sg13g2_nand2_1 _2348_ (.Y(_0358_),
    .A(_0353_),
    .B(_0357_));
 sg13g2_a22oi_1 _2349_ (.Y(_0359_),
    .B1(_0032_),
    .B2(_0341_),
    .A2(_1153_),
    .A1(net52));
 sg13g2_o21ai_1 _2350_ (.B1(_0359_),
    .Y(_0360_),
    .A1(_0320_),
    .A2(_0354_));
 sg13g2_nor2_1 _2351_ (.A(_0356_),
    .B(_0265_),
    .Y(_0361_));
 sg13g2_nor2_1 _2352_ (.A(_0360_),
    .B(_0361_),
    .Y(_0362_));
 sg13g2_nand2_1 _2353_ (.Y(_0363_),
    .A(_0358_),
    .B(_0362_));
 sg13g2_inv_1 _2354_ (.Y(_0364_),
    .A(_0033_));
 sg13g2_xnor2_1 _2355_ (.Y(_0365_),
    .A(_0364_),
    .B(net53));
 sg13g2_inv_1 _2356_ (.Y(_0366_),
    .A(_0365_));
 sg13g2_nand2_1 _2357_ (.Y(_0367_),
    .A(_0363_),
    .B(_0366_));
 sg13g2_nand3_1 _2358_ (.B(_0362_),
    .C(_0365_),
    .A(_0358_),
    .Y(_0368_));
 sg13g2_nand3_1 _2359_ (.B(_0368_),
    .C(net48),
    .A(_0367_),
    .Y(_0369_));
 sg13g2_nand2b_1 _2360_ (.Y(_0370_),
    .B(_0369_),
    .A_N(_0351_));
 sg13g2_nand2_1 _2361_ (.Y(_0371_),
    .A(net34),
    .B(\addr[18] ));
 sg13g2_a21oi_1 _2362_ (.A1(_0370_),
    .A2(_0371_),
    .Y(_0047_),
    .B1(net65));
 sg13g2_o21ai_1 _2363_ (.B1(_1356_),
    .Y(_0372_),
    .A1(\addr_saved0[19] ),
    .A2(_1372_));
 sg13g2_xnor2_1 _2364_ (.Y(_0373_),
    .A(_1160_),
    .B(net53));
 sg13g2_nand2_1 _2365_ (.Y(_0374_),
    .A(_1406_),
    .B(_1434_));
 sg13g2_nand2_1 _2366_ (.Y(_0375_),
    .A(_0374_),
    .B(_1445_));
 sg13g2_nand2_1 _2367_ (.Y(_0376_),
    .A(_0334_),
    .B(_0365_));
 sg13g2_nor2_1 _2368_ (.A(_0376_),
    .B(_0337_),
    .Y(_0377_));
 sg13g2_inv_1 _2369_ (.Y(_0378_),
    .A(_0377_));
 sg13g2_nor2_1 _2370_ (.A(_0378_),
    .B(_0287_),
    .Y(_0379_));
 sg13g2_nand2_1 _2371_ (.Y(_0380_),
    .A(_0375_),
    .B(_0379_));
 sg13g2_inv_1 _2372_ (.Y(_0381_),
    .A(_1153_));
 sg13g2_inv_1 _2373_ (.Y(_0382_),
    .A(\addr[18] ));
 sg13g2_o21ai_1 _2374_ (.B1(_0382_),
    .Y(_0383_),
    .A1(_0364_),
    .A2(_0381_));
 sg13g2_nand2_1 _2375_ (.Y(_0384_),
    .A(net52),
    .B(_0383_));
 sg13g2_o21ai_1 _2376_ (.B1(_0384_),
    .Y(_0385_),
    .A1(_0342_),
    .A2(_0376_));
 sg13g2_nor2_1 _2377_ (.A(_0378_),
    .B(_0292_),
    .Y(_0386_));
 sg13g2_nor2_1 _2378_ (.A(_0385_),
    .B(_0386_),
    .Y(_0387_));
 sg13g2_nand4_1 _2379_ (.B(_1411_),
    .C(_1434_),
    .A(_0379_),
    .Y(_0388_),
    .D(_1416_));
 sg13g2_nand3_1 _2380_ (.B(_0387_),
    .C(_0388_),
    .A(_0380_),
    .Y(_0389_));
 sg13g2_nand2b_1 _2381_ (.Y(_0390_),
    .B(_0389_),
    .A_N(_0373_));
 sg13g2_nand4_1 _2382_ (.B(_0388_),
    .C(_0387_),
    .A(_0380_),
    .Y(_0391_),
    .D(_0373_));
 sg13g2_nand3_1 _2383_ (.B(_0391_),
    .C(net48),
    .A(_0390_),
    .Y(_0392_));
 sg13g2_nand2b_1 _2384_ (.Y(_0393_),
    .B(_0392_),
    .A_N(_0372_));
 sg13g2_nand2_1 _2385_ (.Y(_0394_),
    .A(net34),
    .B(_1160_));
 sg13g2_a21oi_1 _2386_ (.A1(_0393_),
    .A2(_0394_),
    .Y(_0048_),
    .B1(net65));
 sg13g2_o21ai_1 _2387_ (.B1(_1356_),
    .Y(_0395_),
    .A1(\addr_saved0[20] ),
    .A2(net49));
 sg13g2_nand2_1 _2388_ (.Y(_0396_),
    .A(_0365_),
    .B(_0373_));
 sg13g2_or2_1 _2389_ (.X(_0397_),
    .B(_0354_),
    .A(_0396_));
 sg13g2_nor2_1 _2390_ (.A(_0397_),
    .B(_0311_),
    .Y(_0398_));
 sg13g2_nand2_1 _2391_ (.Y(_0399_),
    .A(_0227_),
    .B(_0398_));
 sg13g2_inv_1 _2392_ (.Y(_0400_),
    .A(_1160_));
 sg13g2_a21oi_1 _2393_ (.A1(_0400_),
    .A2(_0382_),
    .Y(_0401_),
    .B1(net50));
 sg13g2_nor2_1 _2394_ (.A(_0396_),
    .B(_0359_),
    .Y(_0402_));
 sg13g2_nor2_1 _2395_ (.A(_0397_),
    .B(_0322_),
    .Y(_0403_));
 sg13g2_nor3_1 _2396_ (.A(_0401_),
    .B(_0402_),
    .C(_0403_),
    .Y(_0404_));
 sg13g2_nand3_1 _2397_ (.B(_1464_),
    .C(_0398_),
    .A(_1471_),
    .Y(_0405_));
 sg13g2_nand3_1 _2398_ (.B(_0404_),
    .C(_0405_),
    .A(_0399_),
    .Y(_0406_));
 sg13g2_xnor2_1 _2399_ (.Y(_0407_),
    .A(_1170_),
    .B(_1362_));
 sg13g2_inv_1 _2400_ (.Y(_0408_),
    .A(_0407_));
 sg13g2_nand2_1 _2401_ (.Y(_0409_),
    .A(_0406_),
    .B(_0408_));
 sg13g2_nand4_1 _2402_ (.B(_0404_),
    .C(_0405_),
    .A(_0399_),
    .Y(_0410_),
    .D(_0407_));
 sg13g2_nand3_1 _2403_ (.B(_0410_),
    .C(_1449_),
    .A(_0409_),
    .Y(_0411_));
 sg13g2_nand2b_1 _2404_ (.Y(_0412_),
    .B(_0411_),
    .A_N(_0395_));
 sg13g2_nand2_1 _2405_ (.Y(_0413_),
    .A(_1358_),
    .B(_1170_));
 sg13g2_a21oi_1 _2406_ (.A1(_0412_),
    .A2(_0413_),
    .Y(_0049_),
    .B1(net65));
 sg13g2_o21ai_1 _2407_ (.B1(net49),
    .Y(_0414_),
    .A1(_1366_),
    .A2(_1460_));
 sg13g2_a21oi_1 _2408_ (.A1(_1366_),
    .A2(_1460_),
    .Y(_0415_),
    .B1(_0414_));
 sg13g2_a21oi_1 _2409_ (.A1(\addr_saved0[2] ),
    .A2(_1098_),
    .Y(_0416_),
    .B1(_0415_));
 sg13g2_o21ai_1 _2410_ (.B1(net71),
    .Y(_0417_),
    .A1(\addr[2] ),
    .A2(net37));
 sg13g2_a21oi_1 _2411_ (.A1(net37),
    .A2(_0416_),
    .Y(_0050_),
    .B1(_0417_));
 sg13g2_o21ai_1 _2412_ (.B1(_1356_),
    .Y(_0418_),
    .A1(\addr_saved0[21] ),
    .A2(_1372_));
 sg13g2_nand2_1 _2413_ (.Y(_0419_),
    .A(_0373_),
    .B(_0407_));
 sg13g2_or2_1 _2414_ (.X(_0420_),
    .B(_0419_),
    .A(_0376_));
 sg13g2_nor2_1 _2415_ (.A(_0338_),
    .B(_0420_),
    .Y(_0421_));
 sg13g2_nand2_1 _2416_ (.Y(_0422_),
    .A(_0248_),
    .B(_0421_));
 sg13g2_nor2b_1 _2417_ (.A(_0420_),
    .B_N(_0343_),
    .Y(_0423_));
 sg13g2_nand2b_1 _2418_ (.Y(_0424_),
    .B(_0400_),
    .A_N(_1170_));
 sg13g2_o21ai_1 _2419_ (.B1(net52),
    .Y(_0425_),
    .A1(_0383_),
    .A2(_0424_));
 sg13g2_nor2b_1 _2420_ (.A(_0423_),
    .B_N(_0425_),
    .Y(_0426_));
 sg13g2_nand3_1 _2421_ (.B(_0239_),
    .C(_0421_),
    .A(_0234_),
    .Y(_0427_));
 sg13g2_nand3_1 _2422_ (.B(_0426_),
    .C(_0427_),
    .A(_0422_),
    .Y(_0428_));
 sg13g2_xnor2_1 _2423_ (.Y(_0429_),
    .A(_0034_),
    .B(_1362_));
 sg13g2_nand2_1 _2424_ (.Y(_0430_),
    .A(_0428_),
    .B(_0429_));
 sg13g2_inv_1 _2425_ (.Y(_0431_),
    .A(_0429_));
 sg13g2_nand4_1 _2426_ (.B(_0426_),
    .C(_0427_),
    .A(_0422_),
    .Y(_0432_),
    .D(_0431_));
 sg13g2_nand3_1 _2427_ (.B(_0432_),
    .C(net48),
    .A(_0430_),
    .Y(_0433_));
 sg13g2_nand2b_1 _2428_ (.Y(_0434_),
    .B(_0433_),
    .A_N(_0418_));
 sg13g2_nand2_1 _2429_ (.Y(_0435_),
    .A(_1358_),
    .B(_1175_));
 sg13g2_a21oi_1 _2430_ (.A1(_0434_),
    .A2(_0435_),
    .Y(_0051_),
    .B1(_1355_));
 sg13g2_nor3_1 _2431_ (.A(_0408_),
    .B(_0429_),
    .C(_0396_),
    .Y(_0436_));
 sg13g2_nand2_1 _2432_ (.Y(_0437_),
    .A(_0436_),
    .B(_0355_));
 sg13g2_inv_1 _2433_ (.Y(_0438_),
    .A(_0437_));
 sg13g2_nand2_1 _2434_ (.Y(_0439_),
    .A(_0266_),
    .B(_0438_));
 sg13g2_nor2b_1 _2435_ (.A(net50),
    .B_N(_1175_),
    .Y(_0440_));
 sg13g2_nand3_1 _2436_ (.B(_0401_),
    .C(_0407_),
    .A(_0431_),
    .Y(_0441_));
 sg13g2_nand3_1 _2437_ (.B(_1170_),
    .C(_0034_),
    .A(net52),
    .Y(_0442_));
 sg13g2_nand3b_1 _2438_ (.B(_0441_),
    .C(_0442_),
    .Y(_0443_),
    .A_N(_0440_));
 sg13g2_a21oi_1 _2439_ (.A1(_0360_),
    .A2(_0436_),
    .Y(_0444_),
    .B1(_0443_));
 sg13g2_nor2_1 _2440_ (.A(_0437_),
    .B(_0268_),
    .Y(_0445_));
 sg13g2_nand2_1 _2441_ (.Y(_0446_),
    .A(_0445_),
    .B(_0275_));
 sg13g2_nand3_1 _2442_ (.B(_0444_),
    .C(_0446_),
    .A(_0439_),
    .Y(_0447_));
 sg13g2_xnor2_1 _2443_ (.Y(_0448_),
    .A(_0035_),
    .B(_1363_));
 sg13g2_nand2_1 _2444_ (.Y(_0449_),
    .A(_0447_),
    .B(_0448_));
 sg13g2_inv_1 _2445_ (.Y(_0450_),
    .A(_0448_));
 sg13g2_nand4_1 _2446_ (.B(_0444_),
    .C(_0446_),
    .A(_0439_),
    .Y(_0451_),
    .D(_0450_));
 sg13g2_nand3_1 _2447_ (.B(_0451_),
    .C(net48),
    .A(_0449_),
    .Y(_0452_));
 sg13g2_inv_1 _2448_ (.Y(_0453_),
    .A(\addr_saved0[22] ));
 sg13g2_a21oi_1 _2449_ (.A1(_0453_),
    .A2(net47),
    .Y(_0454_),
    .B1(_1357_));
 sg13g2_nand2_1 _2450_ (.Y(_0455_),
    .A(_0452_),
    .B(_0454_));
 sg13g2_nand2_1 _2451_ (.Y(_0456_),
    .A(net34),
    .B(\addr[22] ));
 sg13g2_a21oi_1 _2452_ (.A1(_0455_),
    .A2(_0456_),
    .Y(_0052_),
    .B1(_1355_));
 sg13g2_xnor2_1 _2453_ (.Y(_0457_),
    .A(\addr[23] ),
    .B(_1363_));
 sg13g2_nor3_1 _2454_ (.A(_0429_),
    .B(_0448_),
    .C(_0419_),
    .Y(_0458_));
 sg13g2_nand2_1 _2455_ (.Y(_0459_),
    .A(_0458_),
    .B(_0377_));
 sg13g2_inv_1 _2456_ (.Y(_0460_),
    .A(_0459_));
 sg13g2_nand2_1 _2457_ (.Y(_0461_),
    .A(_0293_),
    .B(_0460_));
 sg13g2_a22oi_1 _2458_ (.Y(_0462_),
    .B1(_0035_),
    .B2(_0440_),
    .A2(\addr[22] ),
    .A1(net52));
 sg13g2_nand4_1 _2459_ (.B(_0034_),
    .C(_0035_),
    .A(_1439_),
    .Y(_0463_),
    .D(_0424_));
 sg13g2_nand2_1 _2460_ (.Y(_0464_),
    .A(_0462_),
    .B(_0463_));
 sg13g2_a21oi_1 _2461_ (.A1(_0385_),
    .A2(_0458_),
    .Y(_0465_),
    .B1(_0464_));
 sg13g2_nor2_1 _2462_ (.A(_0459_),
    .B(_0294_),
    .Y(_0466_));
 sg13g2_nand2_1 _2463_ (.Y(_0467_),
    .A(_1418_),
    .B(_0466_));
 sg13g2_nand3_1 _2464_ (.B(_0465_),
    .C(_0467_),
    .A(_0461_),
    .Y(_0468_));
 sg13g2_nand2b_1 _2465_ (.Y(_0469_),
    .B(_0468_),
    .A_N(_0457_));
 sg13g2_nand4_1 _2466_ (.B(_0465_),
    .C(_0467_),
    .A(_0461_),
    .Y(_0470_),
    .D(_0457_));
 sg13g2_nand3_1 _2467_ (.B(_0470_),
    .C(net48),
    .A(_0469_),
    .Y(_0471_));
 sg13g2_inv_1 _2468_ (.Y(_0472_),
    .A(\addr_saved0[23] ));
 sg13g2_a21oi_1 _2469_ (.A1(_0472_),
    .A2(net47),
    .Y(_0473_),
    .B1(_1357_));
 sg13g2_nand2_1 _2470_ (.Y(_0474_),
    .A(_0471_),
    .B(_0473_));
 sg13g2_nand2_1 _2471_ (.Y(_0475_),
    .A(net34),
    .B(\addr[23] ));
 sg13g2_a21oi_1 _2472_ (.A1(_0474_),
    .A2(_0475_),
    .Y(_0053_),
    .B1(net65));
 sg13g2_a21oi_1 _2473_ (.A1(\addr_saved0[3] ),
    .A2(net45),
    .Y(_0476_),
    .B1(net33));
 sg13g2_a21oi_1 _2474_ (.A1(_1415_),
    .A2(_1409_),
    .Y(_0477_),
    .B1(net47));
 sg13g2_o21ai_1 _2475_ (.B1(_0477_),
    .Y(_0478_),
    .A1(_1415_),
    .A2(_1409_));
 sg13g2_a221oi_1 _2476_ (.B2(_0478_),
    .C1(net72),
    .B1(_0476_),
    .A1(_1393_),
    .Y(_0054_),
    .A2(net32));
 sg13g2_a21oi_1 _2477_ (.A1(_1464_),
    .A2(_0270_),
    .Y(_0479_),
    .B1(_1451_));
 sg13g2_o21ai_1 _2478_ (.B1(_0479_),
    .Y(_0480_),
    .A1(_0270_),
    .A2(_1464_));
 sg13g2_a21oi_1 _2479_ (.A1(\addr_saved0[4] ),
    .A2(net45),
    .Y(_0481_),
    .B1(net33));
 sg13g2_a221oi_1 _2480_ (.B2(_0481_),
    .C1(net72),
    .B1(_0480_),
    .A1(_1401_),
    .Y(_0055_),
    .A2(net32));
 sg13g2_o21ai_1 _2481_ (.B1(net49),
    .Y(_0482_),
    .A1(_0269_),
    .A2(_0234_));
 sg13g2_a21o_1 _2482_ (.A2(_0234_),
    .A1(_0269_),
    .B1(_0482_),
    .X(_0483_));
 sg13g2_a21oi_1 _2483_ (.A1(\addr_saved0[5] ),
    .A2(net45),
    .Y(_0484_),
    .B1(net33));
 sg13g2_a221oi_1 _2484_ (.B2(_0484_),
    .C1(net72),
    .B1(_0483_),
    .A1(_1388_),
    .Y(_0056_),
    .A2(net32));
 sg13g2_a21oi_1 _2485_ (.A1(_0276_),
    .A2(_1391_),
    .Y(_0485_),
    .B1(net47));
 sg13g2_o21ai_1 _2486_ (.B1(_0485_),
    .Y(_0486_),
    .A1(_1391_),
    .A2(_0276_));
 sg13g2_a21oi_1 _2487_ (.A1(\addr_saved0[6] ),
    .A2(_1452_),
    .Y(_0487_),
    .B1(net33));
 sg13g2_a221oi_1 _2488_ (.B2(_0487_),
    .C1(net72),
    .B1(_0486_),
    .A1(_1382_),
    .Y(_0057_),
    .A2(_0331_));
 sg13g2_xnor2_1 _2489_ (.Y(_0488_),
    .A(_1429_),
    .B(_1418_));
 sg13g2_nand2_1 _2490_ (.Y(_0489_),
    .A(_0488_),
    .B(_0280_));
 sg13g2_a21oi_1 _2491_ (.A1(\addr_saved0[7] ),
    .A2(_1452_),
    .Y(_0490_),
    .B1(_0282_));
 sg13g2_a221oi_1 _2492_ (.B2(_0490_),
    .C1(net72),
    .B1(_0489_),
    .A1(_1435_),
    .Y(_0058_),
    .A2(net32));
 sg13g2_xnor2_1 _2493_ (.Y(_0491_),
    .A(_1423_),
    .B(_0308_));
 sg13g2_nand2_1 _2494_ (.Y(_0492_),
    .A(_0491_),
    .B(_0280_));
 sg13g2_a21oi_1 _2495_ (.A1(\addr_saved0[8] ),
    .A2(net47),
    .Y(_0493_),
    .B1(_0282_));
 sg13g2_a221oi_1 _2496_ (.B2(_0493_),
    .C1(_1354_),
    .B1(_0492_),
    .A1(_1419_),
    .Y(_0059_),
    .A2(_0331_));
 sg13g2_inv_1 _2497_ (.Y(_0494_),
    .A(\addr[9] ));
 sg13g2_xnor2_1 _2498_ (.Y(_0495_),
    .A(_1431_),
    .B(_0336_));
 sg13g2_nand2_1 _2499_ (.Y(_0496_),
    .A(_0495_),
    .B(_0280_));
 sg13g2_a21oi_1 _2500_ (.A1(\addr_saved0[9] ),
    .A2(net47),
    .Y(_0497_),
    .B1(net33));
 sg13g2_a221oi_1 _2501_ (.B2(_0497_),
    .C1(net72),
    .B1(_0496_),
    .A1(_0494_),
    .Y(_0060_),
    .A2(net32));
 sg13g2_xnor2_1 _2502_ (.Y(_0498_),
    .A(_1430_),
    .B(_0353_));
 sg13g2_nand2_1 _2503_ (.Y(_0499_),
    .A(_0498_),
    .B(_0280_));
 sg13g2_a21oi_1 _2504_ (.A1(\addr_saved0[10] ),
    .A2(net47),
    .Y(_0500_),
    .B1(net33));
 sg13g2_a221oi_1 _2505_ (.B2(_0500_),
    .C1(net72),
    .B1(_0499_),
    .A1(_1442_),
    .Y(_0061_),
    .A2(net32));
 sg13g2_xnor2_1 _2506_ (.Y(_0501_),
    .A(\addr_offset1[1] ),
    .B(_1209_));
 sg13g2_nor3_1 _2507_ (.A(_1062_),
    .B(\i_vga.timing_hor.counter[5] ),
    .C(_1056_),
    .Y(_0502_));
 sg13g2_nor2_1 _2508_ (.A(\i_vga.timing_hor.counter[3] ),
    .B(\i_vga.timing_hor.counter[2] ),
    .Y(_0503_));
 sg13g2_nor2_1 _2509_ (.A(\i_vga.timing_hor.counter[1] ),
    .B(\i_vga.timing_hor.counter[0] ),
    .Y(_0504_));
 sg13g2_nand4_1 _2510_ (.B(_1065_),
    .C(_0503_),
    .A(_0502_),
    .Y(_0505_),
    .D(_0504_));
 sg13g2_a21oi_1 _2511_ (.A1(_0501_),
    .A2(_0505_),
    .Y(_0062_),
    .B1(net65));
 sg13g2_buf_1 _2512_ (.A(_1353_),
    .X(_0506_));
 sg13g2_nand2_2 _2513_ (.Y(_0507_),
    .A(_0505_),
    .B(_0506_));
 sg13g2_nand2_1 _2514_ (.Y(_0508_),
    .A(\addr_offset1[1] ),
    .B(\addr_offset1[2] ));
 sg13g2_nand2b_1 _2515_ (.Y(_0509_),
    .B(_1209_),
    .A_N(_0508_));
 sg13g2_inv_1 _2516_ (.Y(_0510_),
    .A(_0509_));
 sg13g2_a21oi_1 _2517_ (.A1(_1209_),
    .A2(\addr_offset1[1] ),
    .Y(_0511_),
    .B1(\addr_offset1[2] ));
 sg13g2_nor3_1 _2518_ (.A(_0507_),
    .B(_0510_),
    .C(_0511_),
    .Y(_0063_));
 sg13g2_nor2_1 _2519_ (.A(_1394_),
    .B(_0509_),
    .Y(_0512_));
 sg13g2_nor2_1 _2520_ (.A(\addr_offset1[3] ),
    .B(_0510_),
    .Y(_0513_));
 sg13g2_nor3_1 _2521_ (.A(_0507_),
    .B(_0512_),
    .C(_0513_),
    .Y(_0064_));
 sg13g2_nor3_2 _2522_ (.A(_1394_),
    .B(_1398_),
    .C(_0509_),
    .Y(_0514_));
 sg13g2_nor2_1 _2523_ (.A(\addr_offset1[4] ),
    .B(_0512_),
    .Y(_0515_));
 sg13g2_nor3_1 _2524_ (.A(_0507_),
    .B(_0514_),
    .C(_0515_),
    .Y(_0065_));
 sg13g2_nor2_1 _2525_ (.A(\addr_offset1[5] ),
    .B(_0514_),
    .Y(_0516_));
 sg13g2_nor2b_1 _2526_ (.A(_1386_),
    .B_N(_0514_),
    .Y(_0517_));
 sg13g2_nor3_1 _2527_ (.A(_0507_),
    .B(_0516_),
    .C(_0517_),
    .Y(_0066_));
 sg13g2_and3_1 _2528_ (.X(_0518_),
    .A(_0514_),
    .B(\addr_offset1[5] ),
    .C(\addr_offset1[6] ));
 sg13g2_nor2_1 _2529_ (.A(\addr_offset1[6] ),
    .B(_0517_),
    .Y(_0519_));
 sg13g2_nor3_1 _2530_ (.A(_0507_),
    .B(_0518_),
    .C(_0519_),
    .Y(_0067_));
 sg13g2_nor2_1 _2531_ (.A(\addr_offset1[7] ),
    .B(_0518_),
    .Y(_0520_));
 sg13g2_nand2_1 _2532_ (.Y(_0521_),
    .A(_0518_),
    .B(\addr_offset1[7] ));
 sg13g2_inv_1 _2533_ (.Y(_0522_),
    .A(_0521_));
 sg13g2_nor3_1 _2534_ (.A(_0507_),
    .B(_0520_),
    .C(_0522_),
    .Y(_0068_));
 sg13g2_nor2b_1 _2535_ (.A(_0521_),
    .B_N(\addr_offset1[8] ),
    .Y(_0523_));
 sg13g2_nor2_1 _2536_ (.A(\addr_offset1[8] ),
    .B(_0522_),
    .Y(_0524_));
 sg13g2_nor3_1 _2537_ (.A(_0507_),
    .B(_0523_),
    .C(_0524_),
    .Y(_0069_));
 sg13g2_inv_1 _2538_ (.Y(_0525_),
    .A(_0037_));
 sg13g2_nand2_1 _2539_ (.Y(_0526_),
    .A(_1370_),
    .B(\i_video.frame_counter ));
 sg13g2_buf_1 _2540_ (.A(_0526_),
    .X(_0527_));
 sg13g2_inv_1 _2541_ (.Y(_0528_),
    .A(net46));
 sg13g2_buf_1 _2542_ (.A(_0528_),
    .X(_0529_));
 sg13g2_o21ai_1 _2543_ (.B1(net71),
    .Y(_0530_),
    .A1(\addr_saved0[1] ),
    .A2(net44));
 sg13g2_a21oi_1 _2544_ (.A1(_0525_),
    .A2(net44),
    .Y(_0070_),
    .B1(_0530_));
 sg13g2_buf_1 _2545_ (.A(_0528_),
    .X(_0531_));
 sg13g2_o21ai_1 _2546_ (.B1(net71),
    .Y(_0532_),
    .A1(\addr_saved0[11] ),
    .A2(net43));
 sg13g2_nor2_1 _2547_ (.A(\addr[2] ),
    .B(\addr[1] ),
    .Y(_0533_));
 sg13g2_nand2_1 _2548_ (.Y(_0534_),
    .A(_0533_),
    .B(_1393_));
 sg13g2_nor2_1 _2549_ (.A(\addr[4] ),
    .B(_0534_),
    .Y(_0535_));
 sg13g2_nand2_1 _2550_ (.Y(_0536_),
    .A(_0535_),
    .B(_1388_));
 sg13g2_nor2_1 _2551_ (.A(\addr[6] ),
    .B(_0536_),
    .Y(_0537_));
 sg13g2_nand2_1 _2552_ (.Y(_0538_),
    .A(_0537_),
    .B(_1435_));
 sg13g2_nor2_1 _2553_ (.A(\addr[8] ),
    .B(_0538_),
    .Y(_0539_));
 sg13g2_nand2_1 _2554_ (.Y(_0540_),
    .A(_0539_),
    .B(_0494_));
 sg13g2_nor2_1 _2555_ (.A(\addr[10] ),
    .B(_0540_),
    .Y(_0541_));
 sg13g2_nor2_1 _2556_ (.A(_1483_),
    .B(_0541_),
    .Y(_0542_));
 sg13g2_nand2_1 _2557_ (.Y(_0543_),
    .A(_0541_),
    .B(_1483_));
 sg13g2_inv_1 _2558_ (.Y(_0544_),
    .A(_0543_));
 sg13g2_nor3_1 _2559_ (.A(net46),
    .B(_0542_),
    .C(_0544_),
    .Y(_0545_));
 sg13g2_nor2_1 _2560_ (.A(_0532_),
    .B(_0545_),
    .Y(_0071_));
 sg13g2_nor2_1 _2561_ (.A(\addr[12] ),
    .B(_0543_),
    .Y(_0546_));
 sg13g2_nor2_1 _2562_ (.A(net46),
    .B(_0546_),
    .Y(_0547_));
 sg13g2_nand2_1 _2563_ (.Y(_0548_),
    .A(_0543_),
    .B(\addr[12] ));
 sg13g2_o21ai_1 _2564_ (.B1(net71),
    .Y(_0549_),
    .A1(\addr_saved0[12] ),
    .A2(net44));
 sg13g2_a21oi_1 _2565_ (.A1(_0547_),
    .A2(_0548_),
    .Y(_0072_),
    .B1(_0549_));
 sg13g2_xnor2_1 _2566_ (.Y(_0550_),
    .A(_1139_),
    .B(_0546_));
 sg13g2_nand3_1 _2567_ (.B(_1045_),
    .C(_1367_),
    .A(_1036_),
    .Y(_0551_));
 sg13g2_nor3_1 _2568_ (.A(_1031_),
    .B(_0551_),
    .C(_1369_),
    .Y(_0552_));
 sg13g2_nand2_1 _2569_ (.Y(_0553_),
    .A(_0552_),
    .B(\i_video.frame_counter ));
 sg13g2_inv_2 _2570_ (.Y(_0554_),
    .A(_0553_));
 sg13g2_buf_1 _2571_ (.A(_0528_),
    .X(_0555_));
 sg13g2_buf_1 _2572_ (.A(_1353_),
    .X(_0556_));
 sg13g2_o21ai_1 _2573_ (.B1(net69),
    .Y(_0557_),
    .A1(\addr_saved0[13] ),
    .A2(net42));
 sg13g2_a21oi_1 _2574_ (.A1(_0550_),
    .A2(_0554_),
    .Y(_0073_),
    .B1(_0557_));
 sg13g2_nand2_1 _2575_ (.Y(_0558_),
    .A(_0546_),
    .B(_0315_));
 sg13g2_xor2_1 _2576_ (.B(_0558_),
    .A(_1143_),
    .X(_0559_));
 sg13g2_o21ai_1 _2577_ (.B1(net69),
    .Y(_0560_),
    .A1(\addr_saved0[14] ),
    .A2(net42));
 sg13g2_a21oi_1 _2578_ (.A1(_0559_),
    .A2(_0554_),
    .Y(_0074_),
    .B1(_0560_));
 sg13g2_nor2_1 _2579_ (.A(_1143_),
    .B(_0558_),
    .Y(_0561_));
 sg13g2_nor2_1 _2580_ (.A(_0318_),
    .B(_0561_),
    .Y(_0562_));
 sg13g2_nor2_1 _2581_ (.A(net46),
    .B(_0562_),
    .Y(_0563_));
 sg13g2_nand2_1 _2582_ (.Y(_0564_),
    .A(_0561_),
    .B(_0318_));
 sg13g2_o21ai_1 _2583_ (.B1(net69),
    .Y(_0565_),
    .A1(\addr_saved0[15] ),
    .A2(net42));
 sg13g2_a21oi_1 _2584_ (.A1(_0563_),
    .A2(_0564_),
    .Y(_0075_),
    .B1(_0565_));
 sg13g2_nor2_2 _2585_ (.A(\addr[16] ),
    .B(_0564_),
    .Y(_0566_));
 sg13g2_nor2_1 _2586_ (.A(_0527_),
    .B(_0566_),
    .Y(_0567_));
 sg13g2_nand2_1 _2587_ (.Y(_0568_),
    .A(_0564_),
    .B(\addr[16] ));
 sg13g2_o21ai_1 _2588_ (.B1(net69),
    .Y(_0569_),
    .A1(\addr_saved0[16] ),
    .A2(net42));
 sg13g2_a21oi_1 _2589_ (.A1(_0567_),
    .A2(_0568_),
    .Y(_0076_),
    .B1(_0569_));
 sg13g2_xnor2_1 _2590_ (.Y(_0570_),
    .A(_1153_),
    .B(_0566_));
 sg13g2_o21ai_1 _2591_ (.B1(net69),
    .Y(_0571_),
    .A1(\addr_saved0[17] ),
    .A2(net42));
 sg13g2_a21oi_1 _2592_ (.A1(_0570_),
    .A2(_0554_),
    .Y(_0077_),
    .B1(_0571_));
 sg13g2_nand2_1 _2593_ (.Y(_0572_),
    .A(_0566_),
    .B(_0381_));
 sg13g2_xnor2_1 _2594_ (.Y(_0573_),
    .A(_0382_),
    .B(_0572_));
 sg13g2_o21ai_1 _2595_ (.B1(_0556_),
    .Y(_0574_),
    .A1(\addr_saved0[18] ),
    .A2(_0555_));
 sg13g2_a21oi_1 _2596_ (.A1(_0573_),
    .A2(_0554_),
    .Y(_0078_),
    .B1(_0574_));
 sg13g2_nor2_1 _2597_ (.A(\addr[18] ),
    .B(_0572_),
    .Y(_0575_));
 sg13g2_xnor2_1 _2598_ (.Y(_0576_),
    .A(_1160_),
    .B(_0575_));
 sg13g2_o21ai_1 _2599_ (.B1(net69),
    .Y(_0577_),
    .A1(\addr_saved0[19] ),
    .A2(net42));
 sg13g2_a21oi_1 _2600_ (.A1(_0576_),
    .A2(_0554_),
    .Y(_0079_),
    .B1(_0577_));
 sg13g2_nand2_1 _2601_ (.Y(_0578_),
    .A(_0575_),
    .B(_0400_));
 sg13g2_nand2_1 _2602_ (.Y(_0579_),
    .A(_0578_),
    .B(_1170_));
 sg13g2_nor3_1 _2603_ (.A(_1153_),
    .B(\addr[18] ),
    .C(_0424_),
    .Y(_0580_));
 sg13g2_a21oi_1 _2604_ (.A1(_0566_),
    .A2(_0580_),
    .Y(_0581_),
    .B1(_0527_));
 sg13g2_o21ai_1 _2605_ (.B1(_0556_),
    .Y(_0582_),
    .A1(\addr_saved0[20] ),
    .A2(_0555_));
 sg13g2_a21oi_1 _2606_ (.A1(_0579_),
    .A2(_0581_),
    .Y(_0080_),
    .B1(_0582_));
 sg13g2_xor2_1 _2607_ (.B(\addr[1] ),
    .A(\addr[2] ),
    .X(_0583_));
 sg13g2_o21ai_1 _2608_ (.B1(net69),
    .Y(_0584_),
    .A1(\addr_saved0[2] ),
    .A2(net42));
 sg13g2_a21oi_1 _2609_ (.A1(net44),
    .A2(_0583_),
    .Y(_0081_),
    .B1(_0584_));
 sg13g2_nand2_1 _2610_ (.Y(_0585_),
    .A(_0566_),
    .B(_0580_));
 sg13g2_nor2_1 _2611_ (.A(_1175_),
    .B(_0585_),
    .Y(_0586_));
 sg13g2_nor2_1 _2612_ (.A(net46),
    .B(_0586_),
    .Y(_0587_));
 sg13g2_nand2_1 _2613_ (.Y(_0588_),
    .A(_0585_),
    .B(_1175_));
 sg13g2_o21ai_1 _2614_ (.B1(net69),
    .Y(_0589_),
    .A1(\addr_saved0[21] ),
    .A2(net42));
 sg13g2_a21oi_1 _2615_ (.A1(_0587_),
    .A2(_0588_),
    .Y(_0082_),
    .B1(_0589_));
 sg13g2_xnor2_1 _2616_ (.Y(_0590_),
    .A(\addr[22] ),
    .B(_0586_));
 sg13g2_o21ai_1 _2617_ (.B1(net70),
    .Y(_0591_),
    .A1(\addr_saved0[22] ),
    .A2(net43));
 sg13g2_a21oi_1 _2618_ (.A1(_0590_),
    .A2(_0554_),
    .Y(_0083_),
    .B1(_0591_));
 sg13g2_nor3_1 _2619_ (.A(_1175_),
    .B(\addr[22] ),
    .C(_0585_),
    .Y(_0592_));
 sg13g2_xnor2_1 _2620_ (.Y(_0593_),
    .A(\addr[23] ),
    .B(_0592_));
 sg13g2_o21ai_1 _2621_ (.B1(net70),
    .Y(_0594_),
    .A1(\addr_saved0[23] ),
    .A2(_0531_));
 sg13g2_a21oi_1 _2622_ (.A1(_0593_),
    .A2(_0554_),
    .Y(_0084_),
    .B1(_0594_));
 sg13g2_xnor2_1 _2623_ (.Y(_0595_),
    .A(\addr[3] ),
    .B(_0533_));
 sg13g2_o21ai_1 _2624_ (.B1(net70),
    .Y(_0596_),
    .A1(\addr_saved0[3] ),
    .A2(net43));
 sg13g2_a21oi_1 _2625_ (.A1(net44),
    .A2(_0595_),
    .Y(_0085_),
    .B1(_0596_));
 sg13g2_xnor2_1 _2626_ (.Y(_0597_),
    .A(_1401_),
    .B(_0534_));
 sg13g2_o21ai_1 _2627_ (.B1(net70),
    .Y(_0598_),
    .A1(\addr_saved0[4] ),
    .A2(net43));
 sg13g2_a21oi_1 _2628_ (.A1(net44),
    .A2(_0597_),
    .Y(_0086_),
    .B1(_0598_));
 sg13g2_xnor2_1 _2629_ (.Y(_0599_),
    .A(_1193_),
    .B(_0535_));
 sg13g2_o21ai_1 _2630_ (.B1(net70),
    .Y(_0600_),
    .A1(\addr_saved0[5] ),
    .A2(net43));
 sg13g2_a21oi_1 _2631_ (.A1(net44),
    .A2(_0599_),
    .Y(_0087_),
    .B1(_0600_));
 sg13g2_xnor2_1 _2632_ (.Y(_0601_),
    .A(_1382_),
    .B(_0536_));
 sg13g2_o21ai_1 _2633_ (.B1(net70),
    .Y(_0602_),
    .A1(\addr_saved0[6] ),
    .A2(net43));
 sg13g2_a21oi_1 _2634_ (.A1(_0529_),
    .A2(_0601_),
    .Y(_0088_),
    .B1(_0602_));
 sg13g2_xnor2_1 _2635_ (.Y(_0603_),
    .A(_1427_),
    .B(_0537_));
 sg13g2_o21ai_1 _2636_ (.B1(_0506_),
    .Y(_0604_),
    .A1(\addr_saved0[7] ),
    .A2(_0531_));
 sg13g2_a21oi_1 _2637_ (.A1(_0529_),
    .A2(_0603_),
    .Y(_0089_),
    .B1(_0604_));
 sg13g2_nand2_1 _2638_ (.Y(_0605_),
    .A(_0538_),
    .B(\addr[8] ));
 sg13g2_nor2_1 _2639_ (.A(_0539_),
    .B(net46),
    .Y(_0606_));
 sg13g2_o21ai_1 _2640_ (.B1(net70),
    .Y(_0607_),
    .A1(\addr_saved0[8] ),
    .A2(net43));
 sg13g2_a21oi_1 _2641_ (.A1(_0605_),
    .A2(_0606_),
    .Y(_0090_),
    .B1(_0607_));
 sg13g2_nor2_1 _2642_ (.A(_0494_),
    .B(_0539_),
    .Y(_0608_));
 sg13g2_inv_1 _2643_ (.Y(_0609_),
    .A(_0540_));
 sg13g2_nor3_1 _2644_ (.A(net46),
    .B(_0608_),
    .C(_0609_),
    .Y(_0610_));
 sg13g2_o21ai_1 _2645_ (.B1(net71),
    .Y(_0611_),
    .A1(\addr_saved0[9] ),
    .A2(net44));
 sg13g2_nor2_1 _2646_ (.A(_0610_),
    .B(_0611_),
    .Y(_0091_));
 sg13g2_nand2_1 _2647_ (.Y(_0612_),
    .A(_0540_),
    .B(\addr[10] ));
 sg13g2_nor2_1 _2648_ (.A(net46),
    .B(_0541_),
    .Y(_0613_));
 sg13g2_o21ai_1 _2649_ (.B1(net70),
    .Y(_0614_),
    .A1(\addr_saved0[10] ),
    .A2(net43));
 sg13g2_a21oi_1 _2650_ (.A1(_0612_),
    .A2(_0613_),
    .Y(_0092_),
    .B1(_0614_));
 sg13g2_inv_1 _2651_ (.Y(_0615_),
    .A(_1018_));
 sg13g2_nor2_1 _2652_ (.A(\i_spi.bits_remaining[0] ),
    .B(\i_spi.bits_remaining[1] ),
    .Y(_0616_));
 sg13g2_inv_1 _2653_ (.Y(_0617_),
    .A(_0616_));
 sg13g2_nor2_1 _2654_ (.A(\i_spi.bits_remaining[2] ),
    .B(_0617_),
    .Y(_0618_));
 sg13g2_inv_1 _2655_ (.Y(_0619_),
    .A(_0618_));
 sg13g2_nor2_1 _2656_ (.A(\i_spi.bits_remaining[3] ),
    .B(_0619_),
    .Y(_0620_));
 sg13g2_nand2_1 _2657_ (.Y(_0621_),
    .A(_0620_),
    .B(_0021_));
 sg13g2_inv_1 _2658_ (.Y(_0622_),
    .A(_0621_));
 sg13g2_nor2_1 _2659_ (.A(_0615_),
    .B(_0622_),
    .Y(_0623_));
 sg13g2_nor2_1 _2660_ (.A(_1015_),
    .B(_1018_),
    .Y(_0624_));
 sg13g2_nand2_1 _2661_ (.Y(_0625_),
    .A(_1292_),
    .B(_0624_));
 sg13g2_nand2b_1 _2662_ (.Y(_0626_),
    .B(\i_spi.spi_select ),
    .A_N(_1112_));
 sg13g2_nand2_1 _2663_ (.Y(_0627_),
    .A(_0625_),
    .B(_0626_));
 sg13g2_nor2_1 _2664_ (.A(_0623_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_buf_1 _2665_ (.A(_1352_),
    .X(_0629_));
 sg13g2_nand2_1 _2666_ (.Y(_0630_),
    .A(_1099_),
    .B(_1110_));
 sg13g2_nor2_1 _2667_ (.A(net78),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_inv_1 _2668_ (.Y(_0632_),
    .A(_0631_));
 sg13g2_nand3_1 _2669_ (.B(_1016_),
    .C(_1018_),
    .A(_0622_),
    .Y(_0633_));
 sg13g2_nor2b_1 _2670_ (.A(_0632_),
    .B_N(_0633_),
    .Y(_0634_));
 sg13g2_o21ai_1 _2671_ (.B1(_0634_),
    .Y(_0137_),
    .A1(_1016_),
    .A2(_0628_));
 sg13g2_nand2_1 _2672_ (.Y(_0635_),
    .A(_0628_),
    .B(_1015_));
 sg13g2_a21oi_1 _2673_ (.A1(_0635_),
    .A2(_1017_),
    .Y(_0636_),
    .B1(_0632_));
 sg13g2_o21ai_1 _2674_ (.B1(_0636_),
    .Y(_0138_),
    .A1(_1017_),
    .A2(_0635_));
 sg13g2_a21oi_1 _2675_ (.A1(_1017_),
    .A2(_1015_),
    .Y(_0637_),
    .B1(_0019_));
 sg13g2_nor2_1 _2676_ (.A(_0615_),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_o21ai_1 _2677_ (.B1(_0631_),
    .Y(_0639_),
    .A1(\i_spi.fsm_state[2] ),
    .A2(_0628_));
 sg13g2_a21oi_1 _2678_ (.A1(_0628_),
    .A2(_0638_),
    .Y(_0139_),
    .B1(_0639_));
 sg13g2_nor2_2 _2679_ (.A(net78),
    .B(_1096_),
    .Y(_0640_));
 sg13g2_inv_1 _2680_ (.Y(_0641_),
    .A(_0640_));
 sg13g2_nor2b_1 _2681_ (.A(_0641_),
    .B_N(_0036_),
    .Y(_0175_));
 sg13g2_nand2b_1 _2682_ (.Y(_0642_),
    .B(_1061_),
    .A_N(_1090_));
 sg13g2_nor2_2 _2683_ (.A(_1056_),
    .B(_0642_),
    .Y(_0643_));
 sg13g2_inv_1 _2684_ (.Y(_0644_),
    .A(_0643_));
 sg13g2_nor2_1 _2685_ (.A(_1053_),
    .B(_0644_),
    .Y(_0645_));
 sg13g2_a21oi_1 _2686_ (.A1(_0645_),
    .A2(_1050_),
    .Y(_0646_),
    .B1(_0641_));
 sg13g2_o21ai_1 _2687_ (.B1(_0646_),
    .Y(_0176_),
    .A1(_1050_),
    .A2(_0645_));
 sg13g2_nand2_1 _2688_ (.Y(_0647_),
    .A(\i_vga.timing_hor.counter[1] ),
    .B(\i_vga.timing_hor.counter[0] ));
 sg13g2_inv_1 _2689_ (.Y(_0648_),
    .A(_0647_));
 sg13g2_nor3_1 _2690_ (.A(_0648_),
    .B(_0504_),
    .C(_0641_),
    .Y(_0177_));
 sg13g2_inv_1 _2691_ (.Y(_0649_),
    .A(\i_vga.timing_hor.counter[2] ));
 sg13g2_nor2_1 _2692_ (.A(_0649_),
    .B(_0647_),
    .Y(_0650_));
 sg13g2_nor2_1 _2693_ (.A(\i_vga.timing_hor.counter[2] ),
    .B(_0648_),
    .Y(_0651_));
 sg13g2_nor3_1 _2694_ (.A(net78),
    .B(_0650_),
    .C(_0651_),
    .Y(_0178_));
 sg13g2_nor2_1 _2695_ (.A(\i_vga.timing_hor.counter[3] ),
    .B(_0650_),
    .Y(_0652_));
 sg13g2_nor3_1 _2696_ (.A(net78),
    .B(_0652_),
    .C(_1061_),
    .Y(_0179_));
 sg13g2_nor2_1 _2697_ (.A(_1062_),
    .B(_1095_),
    .Y(_0653_));
 sg13g2_nor2_1 _2698_ (.A(\i_vga.timing_hor.counter[4] ),
    .B(_1061_),
    .Y(_0654_));
 sg13g2_nor3_1 _2699_ (.A(_0653_),
    .B(_0654_),
    .C(_0641_),
    .Y(_0180_));
 sg13g2_inv_1 _2700_ (.Y(_0655_),
    .A(_0642_));
 sg13g2_nor2_1 _2701_ (.A(\i_vga.timing_hor.counter[5] ),
    .B(_0653_),
    .Y(_0656_));
 sg13g2_o21ai_1 _2702_ (.B1(_0640_),
    .Y(_0181_),
    .A1(_0655_),
    .A2(_0656_));
 sg13g2_nor2_1 _2703_ (.A(_1066_),
    .B(_0642_),
    .Y(_0657_));
 sg13g2_nor2_1 _2704_ (.A(\i_vga.timing_hor.counter[6] ),
    .B(_0655_),
    .Y(_0658_));
 sg13g2_o21ai_1 _2705_ (.B1(_0640_),
    .Y(_0182_),
    .A1(_0657_),
    .A2(_0658_));
 sg13g2_nor2_1 _2706_ (.A(_1052_),
    .B(_0657_),
    .Y(_0659_));
 sg13g2_nor3_1 _2707_ (.A(_0643_),
    .B(_0641_),
    .C(_0659_),
    .Y(_0183_));
 sg13g2_xnor2_1 _2708_ (.Y(_0660_),
    .A(\i_vga.timing_hor.counter[8] ),
    .B(_0643_));
 sg13g2_nand2_1 _2709_ (.Y(_0184_),
    .A(_0660_),
    .B(_0640_));
 sg13g2_a21oi_1 _2710_ (.A1(_0643_),
    .A2(\i_vga.timing_hor.counter[8] ),
    .Y(_0661_),
    .B1(\i_vga.timing_hor.counter[9] ));
 sg13g2_o21ai_1 _2711_ (.B1(_0640_),
    .Y(_0185_),
    .A1(_0645_),
    .A2(_0661_));
 sg13g2_buf_1 _2712_ (.A(_1207_),
    .X(_0662_));
 sg13g2_buf_1 _2713_ (.A(net77),
    .X(_0663_));
 sg13g2_nor2_1 _2714_ (.A(net68),
    .B(_1206_),
    .Y(_0664_));
 sg13g2_a21o_1 _2715_ (.A2(net68),
    .A1(_1231_),
    .B1(_0664_),
    .X(_0665_));
 sg13g2_nand2b_1 _2716_ (.Y(_0666_),
    .B(_1105_),
    .A_N(_1106_));
 sg13g2_nor2_1 _2717_ (.A(net84),
    .B(_0666_),
    .Y(_0667_));
 sg13g2_nand2_2 _2718_ (.Y(_0668_),
    .A(_0667_),
    .B(_1104_));
 sg13g2_nor2_1 _2719_ (.A(\i_video.run_length[5] ),
    .B(\i_video.run_length[4] ),
    .Y(_0669_));
 sg13g2_nor2_1 _2720_ (.A(_1080_),
    .B(_1082_),
    .Y(_0670_));
 sg13g2_inv_1 _2721_ (.Y(_0671_),
    .A(\i_video.run_length[6] ));
 sg13g2_nand4_1 _2722_ (.B(_0670_),
    .C(_1101_),
    .A(_0669_),
    .Y(_0672_),
    .D(_0671_));
 sg13g2_nor2_2 _2723_ (.A(_0668_),
    .B(_0672_),
    .Y(_0673_));
 sg13g2_inv_1 _2724_ (.Y(_0674_),
    .A(_0673_));
 sg13g2_nor2_1 _2725_ (.A(\i_vga.timing_hor.counter[10] ),
    .B(\i_vga.vblank ),
    .Y(_0675_));
 sg13g2_nand2_1 _2726_ (.Y(_0676_),
    .A(_0674_),
    .B(_0675_));
 sg13g2_inv_1 _2727_ (.Y(_0677_),
    .A(_0022_));
 sg13g2_a21oi_1 _2728_ (.A1(_1222_),
    .A2(_0677_),
    .Y(_0678_),
    .B1(_0020_));
 sg13g2_nor2b_1 _2729_ (.A(_1209_),
    .B_N(_0678_),
    .Y(_0679_));
 sg13g2_inv_1 _2730_ (.Y(_0680_),
    .A(net84));
 sg13g2_nor4_1 _2731_ (.A(_0680_),
    .B(\i_video.run_length[3] ),
    .C(_0666_),
    .D(_0672_),
    .Y(_0681_));
 sg13g2_nand2_1 _2732_ (.Y(_0682_),
    .A(_0679_),
    .B(_0681_));
 sg13g2_inv_2 _2733_ (.Y(_0683_),
    .A(_0682_));
 sg13g2_o21ai_1 _2734_ (.B1(_1087_),
    .Y(_0684_),
    .A1(_0676_),
    .A2(net36));
 sg13g2_inv_1 _2735_ (.Y(_0685_),
    .A(_0018_));
 sg13g2_inv_1 _2736_ (.Y(_0686_),
    .A(_1097_));
 sg13g2_nand2_1 _2737_ (.Y(_0687_),
    .A(_0686_),
    .B(net3));
 sg13g2_inv_1 _2738_ (.Y(_0688_),
    .A(_0687_));
 sg13g2_nor2_1 _2739_ (.A(_0685_),
    .B(_0688_),
    .Y(_0689_));
 sg13g2_nand2_1 _2740_ (.Y(_0690_),
    .A(_0684_),
    .B(_0689_));
 sg13g2_buf_1 _2741_ (.A(\i_video.start ),
    .X(_0691_));
 sg13g2_nand2_1 _2742_ (.Y(_0692_),
    .A(_1370_),
    .B(net3));
 sg13g2_nor2_1 _2743_ (.A(net83),
    .B(_0692_),
    .Y(_0693_));
 sg13g2_inv_1 _2744_ (.Y(_0694_),
    .A(_0679_));
 sg13g2_nor2_1 _2745_ (.A(_0674_),
    .B(_0688_),
    .Y(_0695_));
 sg13g2_nand3_1 _2746_ (.B(_0018_),
    .C(_0695_),
    .A(_0694_),
    .Y(_0696_));
 sg13g2_nor2_1 _2747_ (.A(_0673_),
    .B(_0688_),
    .Y(_0697_));
 sg13g2_inv_2 _2748_ (.Y(_0698_),
    .A(_0675_));
 sg13g2_nand4_1 _2749_ (.B(_0018_),
    .C(_1087_),
    .A(_0697_),
    .Y(_0699_),
    .D(_0698_));
 sg13g2_nand2_1 _2750_ (.Y(_0700_),
    .A(_0696_),
    .B(_0699_));
 sg13g2_nor2_1 _2751_ (.A(_0693_),
    .B(_0700_),
    .Y(_0701_));
 sg13g2_nand2_1 _2752_ (.Y(_0702_),
    .A(_0679_),
    .B(_0686_));
 sg13g2_o21ai_1 _2753_ (.B1(net83),
    .Y(_0703_),
    .A1(net84),
    .A2(_0702_));
 sg13g2_buf_2 _2754_ (.A(_0703_),
    .X(_0704_));
 sg13g2_nand3_1 _2755_ (.B(_0701_),
    .C(_0704_),
    .A(_0690_),
    .Y(_0705_));
 sg13g2_buf_1 _2756_ (.A(_0705_),
    .X(_0706_));
 sg13g2_inv_1 _2757_ (.Y(_0707_),
    .A(_1110_));
 sg13g2_nor2_1 _2758_ (.A(net78),
    .B(_0707_),
    .Y(_0708_));
 sg13g2_o21ai_1 _2759_ (.B1(net56),
    .Y(_0709_),
    .A1(_0665_),
    .A2(net24));
 sg13g2_inv_1 _2760_ (.Y(_0710_),
    .A(\i_video.colour[0] ));
 sg13g2_nand2_1 _2761_ (.Y(_0711_),
    .A(net24),
    .B(_0710_));
 sg13g2_nor2b_1 _2762_ (.A(_0709_),
    .B_N(_0711_),
    .Y(_0198_));
 sg13g2_nor2_1 _2763_ (.A(net68),
    .B(_1253_),
    .Y(_0712_));
 sg13g2_a21o_1 _2764_ (.A2(net68),
    .A1(_1256_),
    .B1(_0712_),
    .X(_0713_));
 sg13g2_o21ai_1 _2765_ (.B1(net56),
    .Y(_0714_),
    .A1(_0713_),
    .A2(net24));
 sg13g2_inv_1 _2766_ (.Y(_0715_),
    .A(\i_video.colour[1] ));
 sg13g2_nand2_1 _2767_ (.Y(_0716_),
    .A(net24),
    .B(_0715_));
 sg13g2_nor2b_1 _2768_ (.A(_0714_),
    .B_N(_0716_),
    .Y(_0199_));
 sg13g2_nor2_1 _2769_ (.A(net68),
    .B(_1258_),
    .Y(_0717_));
 sg13g2_a21o_1 _2770_ (.A2(_0663_),
    .A1(_1261_),
    .B1(_0717_),
    .X(_0718_));
 sg13g2_o21ai_1 _2771_ (.B1(net56),
    .Y(_0719_),
    .A1(_0718_),
    .A2(net24));
 sg13g2_inv_1 _2772_ (.Y(_0720_),
    .A(\i_video.colour[2] ));
 sg13g2_nand2_1 _2773_ (.Y(_0721_),
    .A(_0706_),
    .B(_0720_));
 sg13g2_nor2b_1 _2774_ (.A(_0719_),
    .B_N(_0721_),
    .Y(_0200_));
 sg13g2_nor2_1 _2775_ (.A(net77),
    .B(_1263_),
    .Y(_0722_));
 sg13g2_a21o_1 _2776_ (.A2(_0663_),
    .A1(_1266_),
    .B1(_0722_),
    .X(_0723_));
 sg13g2_o21ai_1 _2777_ (.B1(net56),
    .Y(_0724_),
    .A1(_0723_),
    .A2(net24));
 sg13g2_inv_1 _2778_ (.Y(_0725_),
    .A(\i_video.colour[3] ));
 sg13g2_nand2_1 _2779_ (.Y(_0726_),
    .A(_0706_),
    .B(_0725_));
 sg13g2_nor2b_1 _2780_ (.A(_0724_),
    .B_N(_0726_),
    .Y(_0201_));
 sg13g2_nor2_1 _2781_ (.A(_0662_),
    .B(_1268_),
    .Y(_0727_));
 sg13g2_a21o_1 _2782_ (.A2(net68),
    .A1(_1271_),
    .B1(_0727_),
    .X(_0728_));
 sg13g2_o21ai_1 _2783_ (.B1(net56),
    .Y(_0729_),
    .A1(_0728_),
    .A2(net24));
 sg13g2_inv_1 _2784_ (.Y(_0730_),
    .A(\i_video.colour[4] ));
 sg13g2_nand2_1 _2785_ (.Y(_0731_),
    .A(_0705_),
    .B(_0730_));
 sg13g2_nor2b_1 _2786_ (.A(_0729_),
    .B_N(_0731_),
    .Y(_0202_));
 sg13g2_nor2_1 _2787_ (.A(_0662_),
    .B(_1273_),
    .Y(_0732_));
 sg13g2_a21o_1 _2788_ (.A2(net68),
    .A1(_1276_),
    .B1(_0732_),
    .X(_0733_));
 sg13g2_o21ai_1 _2789_ (.B1(_0708_),
    .Y(_0734_),
    .A1(_0733_),
    .A2(net24));
 sg13g2_inv_1 _2790_ (.Y(_0735_),
    .A(\i_video.colour[5] ));
 sg13g2_nand2_1 _2791_ (.Y(_0736_),
    .A(_0705_),
    .B(_0735_));
 sg13g2_nor2b_1 _2792_ (.A(_0734_),
    .B_N(_0736_),
    .Y(_0203_));
 sg13g2_inv_1 _2793_ (.Y(_0737_),
    .A(_0704_));
 sg13g2_o21ai_1 _2794_ (.B1(\i_video.frame_counter ),
    .Y(_0738_),
    .A1(_0689_),
    .A2(_0737_));
 sg13g2_buf_1 _2795_ (.A(net83),
    .X(_0739_));
 sg13g2_nor2_1 _2796_ (.A(_0016_),
    .B(net83),
    .Y(_0740_));
 sg13g2_a21oi_1 _2797_ (.A1(net3),
    .A2(net76),
    .Y(_0741_),
    .B1(_0740_));
 sg13g2_nand3b_1 _2798_ (.B(_0704_),
    .C(_0741_),
    .Y(_0742_),
    .A_N(_0689_));
 sg13g2_nand3_1 _2799_ (.B(_0742_),
    .C(net56),
    .A(_0738_),
    .Y(_0204_));
 sg13g2_nand2_1 _2800_ (.Y(_0743_),
    .A(_1087_),
    .B(_0675_));
 sg13g2_buf_1 _2801_ (.A(_0682_),
    .X(_0744_));
 sg13g2_buf_1 _2802_ (.A(_0673_),
    .X(_0745_));
 sg13g2_nor2_1 _2803_ (.A(net55),
    .B(_1439_),
    .Y(_0746_));
 sg13g2_o21ai_1 _2804_ (.B1(_0746_),
    .Y(_0747_),
    .A1(_0743_),
    .A2(_0744_));
 sg13g2_inv_1 _2805_ (.Y(_0748_),
    .A(_0692_));
 sg13g2_a21oi_1 _2806_ (.A1(_0694_),
    .A2(net55),
    .Y(_0749_),
    .B1(_0748_));
 sg13g2_nand2_1 _2807_ (.Y(_0750_),
    .A(_0747_),
    .B(_0749_));
 sg13g2_buf_1 _2808_ (.A(net83),
    .X(_0751_));
 sg13g2_a21oi_1 _2809_ (.A1(_0748_),
    .A2(_0016_),
    .Y(_0752_),
    .B1(_0751_));
 sg13g2_nand3_1 _2810_ (.B(_0680_),
    .C(net83),
    .A(_0702_),
    .Y(_0753_));
 sg13g2_nand2_1 _2811_ (.Y(_0754_),
    .A(_0753_),
    .B(net56));
 sg13g2_a21oi_1 _2812_ (.A1(_0750_),
    .A2(_0752_),
    .Y(_0205_),
    .B1(_0754_));
 sg13g2_nand3b_1 _2813_ (.B(_0688_),
    .C(\i_video.frame_counter ),
    .Y(_0755_),
    .A_N(net83));
 sg13g2_nand3_1 _2814_ (.B(_0699_),
    .C(_0755_),
    .A(_0696_),
    .Y(_0756_));
 sg13g2_nor2_1 _2815_ (.A(_1212_),
    .B(_1280_),
    .Y(_0757_));
 sg13g2_a21oi_1 _2816_ (.A1(_1212_),
    .A2(_0004_),
    .Y(_0758_),
    .B1(_0757_));
 sg13g2_nor2_1 _2817_ (.A(_1086_),
    .B(_0673_),
    .Y(_0759_));
 sg13g2_buf_1 _2818_ (.A(_0759_),
    .X(_0760_));
 sg13g2_nand2_1 _2819_ (.Y(_0761_),
    .A(net35),
    .B(net84));
 sg13g2_a22oi_1 _2820_ (.Y(_0762_),
    .B1(net51),
    .B2(_0761_),
    .A2(_0758_),
    .A1(_0673_));
 sg13g2_nor4_1 _2821_ (.A(_1106_),
    .B(\i_video.run_length[3] ),
    .C(_0680_),
    .D(\i_video.run_length[2] ),
    .Y(_0763_));
 sg13g2_nor3_1 _2822_ (.A(\i_video.run_length[7] ),
    .B(_1080_),
    .C(_1082_),
    .Y(_0764_));
 sg13g2_nand4_1 _2823_ (.B(_0671_),
    .C(_0669_),
    .A(_0763_),
    .Y(_0765_),
    .D(_0764_));
 sg13g2_nor3_1 _2824_ (.A(_0765_),
    .B(_0758_),
    .C(_0694_),
    .Y(_0766_));
 sg13g2_nor3_1 _2825_ (.A(net83),
    .B(_0748_),
    .C(_0766_),
    .Y(_0767_));
 sg13g2_nor2b_1 _2826_ (.A(_0762_),
    .B_N(_0767_),
    .Y(_0768_));
 sg13g2_inv_1 _2827_ (.Y(_0769_),
    .A(_0702_));
 sg13g2_nand4_1 _2828_ (.B(_0680_),
    .C(net76),
    .A(_0769_),
    .Y(_0770_),
    .D(_0758_));
 sg13g2_nor2b_1 _2829_ (.A(_0768_),
    .B_N(_0770_),
    .Y(_0771_));
 sg13g2_inv_1 _2830_ (.Y(_0772_),
    .A(net56));
 sg13g2_a21oi_1 _2831_ (.A1(_0756_),
    .A2(net84),
    .Y(_0773_),
    .B1(_0772_));
 sg13g2_o21ai_1 _2832_ (.B1(_0773_),
    .Y(_0215_),
    .A1(_0756_),
    .A2(_0771_));
 sg13g2_a21oi_1 _2833_ (.A1(_1208_),
    .A2(_1111_),
    .Y(_0226_),
    .B1(_0632_));
 sg13g2_nor2_1 _2834_ (.A(_1015_),
    .B(net66),
    .Y(_0774_));
 sg13g2_nor3_1 _2835_ (.A(_0019_),
    .B(_1117_),
    .C(_0774_),
    .Y(_0775_));
 sg13g2_a21oi_1 _2836_ (.A1(_0622_),
    .A2(_0775_),
    .Y(_0776_),
    .B1(_0630_));
 sg13g2_nand3_1 _2837_ (.B(_0626_),
    .C(_0776_),
    .A(_0625_),
    .Y(_0777_));
 sg13g2_inv_2 _2838_ (.Y(_0778_),
    .A(_0777_));
 sg13g2_nor2_1 _2839_ (.A(_1015_),
    .B(_1118_),
    .Y(_0779_));
 sg13g2_inv_1 _2840_ (.Y(_0780_),
    .A(_0779_));
 sg13g2_a21oi_1 _2841_ (.A1(_0622_),
    .A2(_0780_),
    .Y(_0781_),
    .B1(_0624_));
 sg13g2_inv_1 _2842_ (.Y(_0782_),
    .A(\i_spi.bits_remaining[0] ));
 sg13g2_a21oi_1 _2843_ (.A1(_0781_),
    .A2(_0782_),
    .Y(_0783_),
    .B1(\i_spi.spi_select ));
 sg13g2_buf_1 _2844_ (.A(_1218_),
    .X(_0784_));
 sg13g2_o21ai_1 _2845_ (.B1(_0784_),
    .Y(_0785_),
    .A1(\i_spi.bits_remaining[0] ),
    .A2(_0778_));
 sg13g2_a21oi_1 _2846_ (.A1(_0778_),
    .A2(_0783_),
    .Y(_0116_),
    .B1(_0785_));
 sg13g2_xnor2_1 _2847_ (.Y(_0786_),
    .A(\i_spi.bits_remaining[0] ),
    .B(\i_spi.bits_remaining[1] ));
 sg13g2_o21ai_1 _2848_ (.B1(_1018_),
    .Y(_0787_),
    .A1(_1118_),
    .A2(_0621_));
 sg13g2_a21oi_1 _2849_ (.A1(_0621_),
    .A2(_0786_),
    .Y(_0788_),
    .B1(_0787_));
 sg13g2_o21ai_1 _2850_ (.B1(_0784_),
    .Y(_0789_),
    .A1(\i_spi.bits_remaining[1] ),
    .A2(_0778_));
 sg13g2_a21oi_1 _2851_ (.A1(_0778_),
    .A2(_0788_),
    .Y(_0117_),
    .B1(_0789_));
 sg13g2_a21oi_1 _2852_ (.A1(_0002_),
    .A2(_0616_),
    .Y(_0790_),
    .B1(_0622_));
 sg13g2_o21ai_1 _2853_ (.B1(_0790_),
    .Y(_0791_),
    .A1(_0002_),
    .A2(_0616_));
 sg13g2_a21oi_1 _2854_ (.A1(_0791_),
    .A2(_0781_),
    .Y(_0792_),
    .B1(\i_spi.spi_select ));
 sg13g2_o21ai_1 _2855_ (.B1(net82),
    .Y(_0793_),
    .A1(\i_spi.bits_remaining[2] ),
    .A2(_0778_));
 sg13g2_a21oi_1 _2856_ (.A1(_0778_),
    .A2(_0792_),
    .Y(_0118_),
    .B1(_0793_));
 sg13g2_inv_1 _2857_ (.Y(_0794_),
    .A(\i_spi.bits_remaining[3] ));
 sg13g2_inv_1 _2858_ (.Y(_0795_),
    .A(_0620_));
 sg13g2_nand2_1 _2859_ (.Y(_0796_),
    .A(_0619_),
    .B(\i_spi.bits_remaining[3] ));
 sg13g2_a221oi_1 _2860_ (.B2(_1121_),
    .C1(_0615_),
    .B1(_0622_),
    .A1(_0795_),
    .Y(_0797_),
    .A2(_0796_));
 sg13g2_o21ai_1 _2861_ (.B1(net82),
    .Y(_0798_),
    .A1(_0797_),
    .A2(_0777_));
 sg13g2_a21oi_1 _2862_ (.A1(_0794_),
    .A2(_0777_),
    .Y(_0119_),
    .B1(_0798_));
 sg13g2_nor2_1 _2863_ (.A(_0021_),
    .B(_0620_),
    .Y(_0799_));
 sg13g2_a21o_1 _2864_ (.A2(_0779_),
    .A1(_0622_),
    .B1(_0799_),
    .X(_0800_));
 sg13g2_nand3_1 _2865_ (.B(_1018_),
    .C(_0800_),
    .A(_0778_),
    .Y(_0801_));
 sg13g2_nand2_1 _2866_ (.Y(_0802_),
    .A(_0777_),
    .B(\i_spi.bits_remaining[4] ));
 sg13g2_buf_1 _2867_ (.A(net78),
    .X(_0803_));
 sg13g2_a21oi_1 _2868_ (.A1(_0801_),
    .A2(_0802_),
    .Y(_0120_),
    .B1(net67));
 sg13g2_nand4_1 _2869_ (.B(_1015_),
    .C(_1110_),
    .A(_1099_),
    .Y(_0804_),
    .D(_0787_));
 sg13g2_nand2b_1 _2870_ (.Y(_0805_),
    .B(_0626_),
    .A_N(_0804_));
 sg13g2_nand2_1 _2871_ (.Y(_0806_),
    .A(_0805_),
    .B(\i_spi.spi_data_oe[0] ));
 sg13g2_a21oi_1 _2872_ (.A1(_0806_),
    .A2(_1126_),
    .Y(_0140_),
    .B1(net67));
 sg13g2_o21ai_1 _2873_ (.B1(net68),
    .Y(_0807_),
    .A1(_1216_),
    .A2(_1209_));
 sg13g2_a21oi_1 _2874_ (.A1(_1223_),
    .A2(_0807_),
    .Y(_0141_),
    .B1(net67));
 sg13g2_nand2_1 _2875_ (.Y(_0808_),
    .A(_1293_),
    .B(_1216_));
 sg13g2_a21oi_1 _2876_ (.A1(_0808_),
    .A2(_1291_),
    .Y(_0158_),
    .B1(net67));
 sg13g2_nand3_1 _2877_ (.B(\i_vga.timing_hor.counter[1] ),
    .C(\i_vga.timing_hor.counter[2] ),
    .A(_1058_),
    .Y(_0809_));
 sg13g2_nor2_1 _2878_ (.A(\i_vga.timing_hor.counter[8] ),
    .B(\i_vga.timing_hor.counter[10] ),
    .Y(_0810_));
 sg13g2_nand4_1 _2879_ (.B(\i_vga.timing_hor.counter[3] ),
    .C(\i_vga.timing_hor.counter[9] ),
    .A(_1091_),
    .Y(_0811_),
    .D(_0810_));
 sg13g2_nor2_1 _2880_ (.A(_0809_),
    .B(_0811_),
    .Y(_0812_));
 sg13g2_nand2_1 _2881_ (.Y(_0813_),
    .A(_0812_),
    .B(\i_vga.timing_ver.counter[0] ));
 sg13g2_inv_1 _2882_ (.Y(_0814_),
    .A(_0813_));
 sg13g2_nor2_1 _2883_ (.A(\i_vga.timing_ver.counter[0] ),
    .B(_0812_),
    .Y(_0815_));
 sg13g2_nand2_1 _2884_ (.Y(_0816_),
    .A(_1020_),
    .B(\i_vga.timing_ver.counter[0] ));
 sg13g2_nor4_2 _2885_ (.A(\i_vga.timing_hor.counter[0] ),
    .B(_0816_),
    .C(_1060_),
    .Y(_0817_),
    .D(_1094_));
 sg13g2_nand2_1 _2886_ (.Y(_0818_),
    .A(_0817_),
    .B(_1045_));
 sg13g2_inv_1 _2887_ (.Y(_0819_),
    .A(_0818_));
 sg13g2_nand2_1 _2888_ (.Y(_0820_),
    .A(\i_vga.timing_ver.counter[7] ),
    .B(\i_vga.timing_ver.counter[8] ));
 sg13g2_nand2_1 _2889_ (.Y(_0821_),
    .A(_1028_),
    .B(\i_vga.timing_ver.counter[4] ));
 sg13g2_nor4_1 _2890_ (.A(\i_vga.timing_ver.counter[9] ),
    .B(_1030_),
    .C(_0820_),
    .D(_0821_),
    .Y(_0822_));
 sg13g2_a21oi_2 _2891_ (.B1(net78),
    .Y(_0823_),
    .A2(_0822_),
    .A1(_0819_));
 sg13g2_o21ai_1 _2892_ (.B1(_0823_),
    .Y(_0186_),
    .A1(_0814_),
    .A2(_0815_));
 sg13g2_nand3_1 _2893_ (.B(_1026_),
    .C(\i_vga.timing_ver.counter[4] ),
    .A(_0819_),
    .Y(_0824_));
 sg13g2_nor2b_1 _2894_ (.A(_0824_),
    .B_N(_1033_),
    .Y(_0825_));
 sg13g2_xnor2_1 _2895_ (.Y(_0826_),
    .A(_1030_),
    .B(_0825_));
 sg13g2_nand2_1 _2896_ (.Y(_0187_),
    .A(_0826_),
    .B(_0823_));
 sg13g2_nor2_1 _2897_ (.A(_1021_),
    .B(_0813_),
    .Y(_0827_));
 sg13g2_nor2_1 _2898_ (.A(_1020_),
    .B(_0814_),
    .Y(_0828_));
 sg13g2_o21ai_1 _2899_ (.B1(_0823_),
    .Y(_0188_),
    .A1(_0827_),
    .A2(_0828_));
 sg13g2_xnor2_1 _2900_ (.Y(_0829_),
    .A(\i_vga.timing_ver.counter[2] ),
    .B(_0817_));
 sg13g2_nor2_1 _2901_ (.A(net67),
    .B(_0829_),
    .Y(_0189_));
 sg13g2_a21oi_1 _2902_ (.A1(_0817_),
    .A2(\i_vga.timing_ver.counter[2] ),
    .Y(_0830_),
    .B1(\i_vga.timing_ver.counter[3] ));
 sg13g2_nor3_1 _2903_ (.A(net78),
    .B(_0819_),
    .C(_0830_),
    .Y(_0190_));
 sg13g2_nor2_1 _2904_ (.A(\i_vga.timing_ver.counter[4] ),
    .B(_0819_),
    .Y(_0831_));
 sg13g2_nor2_1 _2905_ (.A(_1025_),
    .B(_0813_),
    .Y(_0832_));
 sg13g2_o21ai_1 _2906_ (.B1(_0823_),
    .Y(_0191_),
    .A1(_0831_),
    .A2(_0832_));
 sg13g2_or2_1 _2907_ (.X(_0833_),
    .B(_0832_),
    .A(_1026_));
 sg13g2_nand2_1 _2908_ (.Y(_0834_),
    .A(_0832_),
    .B(_1026_));
 sg13g2_and3_1 _2909_ (.X(_0192_),
    .A(_0833_),
    .B(_0823_),
    .C(_0834_));
 sg13g2_a21oi_1 _2910_ (.A1(_0832_),
    .A2(_1026_),
    .Y(_0835_),
    .B1(\i_vga.timing_ver.counter[6] ));
 sg13g2_nor2_2 _2911_ (.A(_1027_),
    .B(_0834_),
    .Y(_0836_));
 sg13g2_o21ai_1 _2912_ (.B1(_0823_),
    .Y(_0193_),
    .A1(_0835_),
    .A2(_0836_));
 sg13g2_xnor2_1 _2913_ (.Y(_0837_),
    .A(\i_vga.timing_ver.counter[7] ),
    .B(_0836_));
 sg13g2_buf_1 _2914_ (.A(_1218_),
    .X(_0838_));
 sg13g2_nand2_1 _2915_ (.Y(_0194_),
    .A(_0837_),
    .B(net81));
 sg13g2_a21oi_1 _2916_ (.A1(_0836_),
    .A2(\i_vga.timing_ver.counter[7] ),
    .Y(_0839_),
    .B1(\i_vga.timing_ver.counter[8] ));
 sg13g2_nand2b_1 _2917_ (.Y(_0840_),
    .B(_0836_),
    .A_N(_0820_));
 sg13g2_nand2b_1 _2918_ (.Y(_0841_),
    .B(_0840_),
    .A_N(_0839_));
 sg13g2_nand2_1 _2919_ (.Y(_0195_),
    .A(_0841_),
    .B(net81));
 sg13g2_xor2_1 _2920_ (.B(_0840_),
    .A(\i_vga.timing_ver.counter[9] ),
    .X(_0842_));
 sg13g2_nand2_1 _2921_ (.Y(_0196_),
    .A(_0842_),
    .B(_0823_));
 sg13g2_nand2_2 _2922_ (.Y(_0843_),
    .A(_1110_),
    .B(_0018_));
 sg13g2_nand2_1 _2923_ (.Y(_0844_),
    .A(_0753_),
    .B(_0843_));
 sg13g2_nand2_1 _2924_ (.Y(_0845_),
    .A(_0844_),
    .B(clear_addr));
 sg13g2_nand2_1 _2925_ (.Y(_0846_),
    .A(_0843_),
    .B(net84));
 sg13g2_a21oi_1 _2926_ (.A1(_0845_),
    .A2(_0846_),
    .Y(_0197_),
    .B1(net67));
 sg13g2_inv_1 _2927_ (.Y(_0847_),
    .A(\i_video.repeat_count[0] ));
 sg13g2_nor3_2 _2928_ (.A(_1087_),
    .B(_0843_),
    .C(_0748_),
    .Y(_0848_));
 sg13g2_inv_2 _2929_ (.Y(_0849_),
    .A(_0848_));
 sg13g2_inv_1 _2930_ (.Y(_0850_),
    .A(_0003_));
 sg13g2_a21oi_1 _2931_ (.A1(_1079_),
    .A2(_0710_),
    .Y(_0851_),
    .B1(_0850_));
 sg13g2_o21ai_1 _2932_ (.B1(net82),
    .Y(_0852_),
    .A1(_0851_),
    .A2(_0849_));
 sg13g2_a21oi_1 _2933_ (.A1(_0847_),
    .A2(_0849_),
    .Y(_0206_),
    .B1(_0852_));
 sg13g2_nor4_1 _2934_ (.A(_1087_),
    .B(net55),
    .C(_0843_),
    .D(_0688_),
    .Y(_0853_));
 sg13g2_nand2_1 _2935_ (.Y(_0854_),
    .A(_1079_),
    .B(_0003_));
 sg13g2_buf_1 _2936_ (.A(_0854_),
    .X(_0855_));
 sg13g2_inv_2 _2937_ (.Y(_0856_),
    .A(_0855_));
 sg13g2_nand2_1 _2938_ (.Y(_0857_),
    .A(\i_video.repeat_count[1] ),
    .B(\i_video.repeat_count[0] ));
 sg13g2_nor2_1 _2939_ (.A(\i_video.repeat_count[1] ),
    .B(\i_video.repeat_count[0] ),
    .Y(_0858_));
 sg13g2_inv_1 _2940_ (.Y(_0859_),
    .A(_0858_));
 sg13g2_a21oi_1 _2941_ (.A1(_0857_),
    .A2(_0859_),
    .Y(_0860_),
    .B1(_0856_));
 sg13g2_a21oi_1 _2942_ (.A1(\i_video.colour[1] ),
    .A2(_0856_),
    .Y(_0861_),
    .B1(_0860_));
 sg13g2_o21ai_1 _2943_ (.B1(net82),
    .Y(_0862_),
    .A1(\i_video.repeat_count[1] ),
    .A2(_0848_));
 sg13g2_a21oi_1 _2944_ (.A1(_0853_),
    .A2(_0861_),
    .Y(_0207_),
    .B1(_0862_));
 sg13g2_xor2_1 _2945_ (.B(_0858_),
    .A(\i_video.repeat_count[2] ),
    .X(_0863_));
 sg13g2_nor2_1 _2946_ (.A(_0720_),
    .B(net61),
    .Y(_0864_));
 sg13g2_a21oi_1 _2947_ (.A1(net61),
    .A2(_0863_),
    .Y(_0865_),
    .B1(_0864_));
 sg13g2_o21ai_1 _2948_ (.B1(net82),
    .Y(_0866_),
    .A1(\i_video.repeat_count[2] ),
    .A2(_0848_));
 sg13g2_a21oi_1 _2949_ (.A1(_0853_),
    .A2(_0865_),
    .Y(_0208_),
    .B1(_0866_));
 sg13g2_inv_1 _2950_ (.Y(_0867_),
    .A(\i_video.repeat_count[3] ));
 sg13g2_o21ai_1 _2951_ (.B1(\i_video.repeat_count[3] ),
    .Y(_0868_),
    .A1(\i_video.repeat_count[2] ),
    .A2(_0859_));
 sg13g2_nor3_1 _2952_ (.A(\i_video.repeat_count[3] ),
    .B(\i_video.repeat_count[2] ),
    .C(_0859_),
    .Y(_0869_));
 sg13g2_nor2_1 _2953_ (.A(_0869_),
    .B(_0856_),
    .Y(_0870_));
 sg13g2_a22oi_1 _2954_ (.Y(_0871_),
    .B1(_0868_),
    .B2(_0870_),
    .A2(_0856_),
    .A1(_0725_));
 sg13g2_o21ai_1 _2955_ (.B1(net82),
    .Y(_0872_),
    .A1(_0871_),
    .A2(_0849_));
 sg13g2_a21oi_1 _2956_ (.A1(_0867_),
    .A2(_0849_),
    .Y(_0209_),
    .B1(_0872_));
 sg13g2_nand3_1 _2957_ (.B(_1074_),
    .C(_0847_),
    .A(_1073_),
    .Y(_0873_));
 sg13g2_a21oi_1 _2958_ (.A1(net61),
    .A2(_0873_),
    .Y(_0874_),
    .B1(_0849_));
 sg13g2_o21ai_1 _2959_ (.B1(_0874_),
    .Y(_0875_),
    .A1(\i_video.colour[4] ),
    .A2(net61));
 sg13g2_o21ai_1 _2960_ (.B1(\i_video.repeat_count[4] ),
    .Y(_0876_),
    .A1(_0870_),
    .A2(_0849_));
 sg13g2_a21oi_1 _2961_ (.A1(_0875_),
    .A2(_0876_),
    .Y(_0210_),
    .B1(net67));
 sg13g2_nand2b_1 _2962_ (.Y(_0877_),
    .B(\i_video.repeat_count[5] ),
    .A_N(_0874_));
 sg13g2_nor2_1 _2963_ (.A(\i_video.repeat_count[5] ),
    .B(_0873_),
    .Y(_0878_));
 sg13g2_nand2_1 _2964_ (.Y(_0879_),
    .A(net61),
    .B(_0878_));
 sg13g2_o21ai_1 _2965_ (.B1(_0879_),
    .Y(_0880_),
    .A1(_0735_),
    .A2(net61));
 sg13g2_nand2_1 _2966_ (.Y(_0881_),
    .A(_0848_),
    .B(_0880_));
 sg13g2_a21oi_1 _2967_ (.A1(_0877_),
    .A2(_0881_),
    .Y(_0211_),
    .B1(_0803_));
 sg13g2_inv_1 _2968_ (.Y(_0882_),
    .A(\i_video.repeat_count[6] ));
 sg13g2_nand2_1 _2969_ (.Y(_0883_),
    .A(_0856_),
    .B(_0680_));
 sg13g2_o21ai_1 _2970_ (.B1(_0883_),
    .Y(_0884_),
    .A1(_0882_),
    .A2(_0879_));
 sg13g2_nand2_1 _2971_ (.Y(_0885_),
    .A(_0878_),
    .B(_0882_));
 sg13g2_a21oi_1 _2972_ (.A1(net61),
    .A2(_0885_),
    .Y(_0886_),
    .B1(_0849_));
 sg13g2_inv_1 _2973_ (.Y(_0887_),
    .A(_0886_));
 sg13g2_a221oi_1 _2974_ (.B2(_0882_),
    .C1(_0629_),
    .B1(_0887_),
    .A1(_0848_),
    .Y(_0212_),
    .A2(_0884_));
 sg13g2_nor2_1 _2975_ (.A(\i_video.repeat_count[7] ),
    .B(_0887_),
    .Y(_0888_));
 sg13g2_o21ai_1 _2976_ (.B1(_0888_),
    .Y(_0889_),
    .A1(_1106_),
    .A2(net61));
 sg13g2_nand2_1 _2977_ (.Y(_0890_),
    .A(_0887_),
    .B(\i_video.repeat_count[7] ));
 sg13g2_a21oi_1 _2978_ (.A1(_0889_),
    .A2(_0890_),
    .Y(_0213_),
    .B1(_0803_));
 sg13g2_nor2_1 _2979_ (.A(\i_video.repeat_count[8] ),
    .B(_0888_),
    .Y(_0891_));
 sg13g2_nor2_1 _2980_ (.A(\i_video.repeat_count[8] ),
    .B(_0856_),
    .Y(_0892_));
 sg13g2_a21oi_1 _2981_ (.A1(\i_video.run_length[2] ),
    .A2(_0856_),
    .Y(_0893_),
    .B1(_0892_));
 sg13g2_a21oi_1 _2982_ (.A1(_0888_),
    .A2(_0893_),
    .Y(_0894_),
    .B1(_0629_));
 sg13g2_nor2b_1 _2983_ (.A(_0891_),
    .B_N(_0894_),
    .Y(_0214_));
 sg13g2_buf_1 _2984_ (.A(_1207_),
    .X(_0895_));
 sg13g2_nor2_1 _2985_ (.A(_1207_),
    .B(_0005_),
    .Y(_0896_));
 sg13g2_a21o_1 _2986_ (.A2(net74),
    .A1(_1283_),
    .B1(_0896_),
    .X(_0897_));
 sg13g2_inv_1 _2987_ (.Y(_0898_),
    .A(_0897_));
 sg13g2_a21oi_1 _2988_ (.A1(_0897_),
    .A2(_0745_),
    .Y(_0899_),
    .B1(_0739_));
 sg13g2_nor2_1 _2989_ (.A(_1106_),
    .B(net84),
    .Y(_0900_));
 sg13g2_nand3b_1 _2990_ (.B(_0682_),
    .C(_1108_),
    .Y(_0901_),
    .A_N(_0900_));
 sg13g2_nand2_1 _2991_ (.Y(_0902_),
    .A(net36),
    .B(_0898_));
 sg13g2_nand3_1 _2992_ (.B(net51),
    .C(_0902_),
    .A(_0901_),
    .Y(_0903_));
 sg13g2_a22oi_1 _2993_ (.Y(_0904_),
    .B1(_0899_),
    .B2(_0903_),
    .A2(_0898_),
    .A1(net75));
 sg13g2_nand3b_1 _2994_ (.B(_0704_),
    .C(_1110_),
    .Y(_0905_),
    .A_N(_0693_));
 sg13g2_nor2_1 _2995_ (.A(_0756_),
    .B(_0905_),
    .Y(_0906_));
 sg13g2_nand2_1 _2996_ (.Y(_0907_),
    .A(_0904_),
    .B(net29));
 sg13g2_inv_1 _2997_ (.Y(_0908_),
    .A(_0756_));
 sg13g2_a21oi_1 _2998_ (.A1(_0908_),
    .A2(_0704_),
    .Y(_0909_),
    .B1(_0707_));
 sg13g2_nand2_1 _2999_ (.Y(_0910_),
    .A(net28),
    .B(_1106_));
 sg13g2_nand3_1 _3000_ (.B(_0910_),
    .C(net81),
    .A(_0907_),
    .Y(_0216_));
 sg13g2_nor2_1 _3001_ (.A(net74),
    .B(_0006_),
    .Y(_0911_));
 sg13g2_a21o_1 _3002_ (.A2(net77),
    .A1(_1286_),
    .B1(_0911_),
    .X(_0912_));
 sg13g2_inv_1 _3003_ (.Y(_0913_),
    .A(_0912_));
 sg13g2_a21oi_1 _3004_ (.A1(_0912_),
    .A2(_0745_),
    .Y(_0914_),
    .B1(net76));
 sg13g2_inv_1 _3005_ (.Y(_0915_),
    .A(_0667_));
 sg13g2_o21ai_1 _3006_ (.B1(\i_video.run_length[2] ),
    .Y(_0916_),
    .A1(_1106_),
    .A2(_1107_));
 sg13g2_nand3_1 _3007_ (.B(_0915_),
    .C(_0916_),
    .A(net35),
    .Y(_0917_));
 sg13g2_nand2_1 _3008_ (.Y(_0918_),
    .A(net36),
    .B(_0913_));
 sg13g2_nand3_1 _3009_ (.B(_0918_),
    .C(net51),
    .A(_0917_),
    .Y(_0919_));
 sg13g2_a22oi_1 _3010_ (.Y(_0920_),
    .B1(_0914_),
    .B2(_0919_),
    .A2(_0913_),
    .A1(net75));
 sg13g2_nand2_1 _3011_ (.Y(_0921_),
    .A(_0920_),
    .B(net29));
 sg13g2_nand2_1 _3012_ (.Y(_0922_),
    .A(net28),
    .B(\i_video.run_length[2] ));
 sg13g2_nand3_1 _3013_ (.B(_0922_),
    .C(net81),
    .A(_0921_),
    .Y(_0217_));
 sg13g2_nor2_1 _3014_ (.A(_0895_),
    .B(_0007_),
    .Y(_0923_));
 sg13g2_a21o_1 _3015_ (.A2(net77),
    .A1(_1289_),
    .B1(_0923_),
    .X(_0924_));
 sg13g2_inv_1 _3016_ (.Y(_0925_),
    .A(_0924_));
 sg13g2_a21oi_1 _3017_ (.A1(_0924_),
    .A2(net55),
    .Y(_0926_),
    .B1(_0739_));
 sg13g2_nand2_1 _3018_ (.Y(_0927_),
    .A(_0915_),
    .B(\i_video.run_length[3] ));
 sg13g2_nand3_1 _3019_ (.B(_0668_),
    .C(_0927_),
    .A(_0744_),
    .Y(_0928_));
 sg13g2_nand2_1 _3020_ (.Y(_0929_),
    .A(net36),
    .B(_0925_));
 sg13g2_nand3_1 _3021_ (.B(_0929_),
    .C(_0760_),
    .A(_0928_),
    .Y(_0930_));
 sg13g2_a22oi_1 _3022_ (.Y(_0931_),
    .B1(_0926_),
    .B2(_0930_),
    .A2(_0925_),
    .A1(net75));
 sg13g2_nand2_1 _3023_ (.Y(_0932_),
    .A(_0931_),
    .B(net29));
 sg13g2_nand2_1 _3024_ (.Y(_0933_),
    .A(net28),
    .B(\i_video.run_length[3] ));
 sg13g2_nand3_1 _3025_ (.B(_0933_),
    .C(net81),
    .A(_0932_),
    .Y(_0218_));
 sg13g2_nor2_1 _3026_ (.A(net74),
    .B(_0008_),
    .Y(_0934_));
 sg13g2_a21o_1 _3027_ (.A2(net77),
    .A1(_1236_),
    .B1(_0934_),
    .X(_0935_));
 sg13g2_inv_1 _3028_ (.Y(_0936_),
    .A(_0935_));
 sg13g2_a21oi_1 _3029_ (.A1(_0935_),
    .A2(net55),
    .Y(_0937_),
    .B1(net76));
 sg13g2_nor2_1 _3030_ (.A(\i_video.run_length[4] ),
    .B(_0668_),
    .Y(_0938_));
 sg13g2_inv_1 _3031_ (.Y(_0939_),
    .A(_0938_));
 sg13g2_nand2_1 _3032_ (.Y(_0940_),
    .A(_0668_),
    .B(\i_video.run_length[4] ));
 sg13g2_nand3_1 _3033_ (.B(_0939_),
    .C(_0940_),
    .A(net35),
    .Y(_0941_));
 sg13g2_nand2_1 _3034_ (.Y(_0942_),
    .A(net36),
    .B(_0936_));
 sg13g2_nand3_1 _3035_ (.B(_0942_),
    .C(net51),
    .A(_0941_),
    .Y(_0943_));
 sg13g2_a22oi_1 _3036_ (.Y(_0944_),
    .B1(_0937_),
    .B2(_0943_),
    .A2(_0936_),
    .A1(net75));
 sg13g2_nand2_1 _3037_ (.Y(_0945_),
    .A(_0944_),
    .B(net29));
 sg13g2_nand2_1 _3038_ (.Y(_0946_),
    .A(net28),
    .B(\i_video.run_length[4] ));
 sg13g2_nand3_1 _3039_ (.B(_0946_),
    .C(net81),
    .A(_0945_),
    .Y(_0219_));
 sg13g2_nor2_1 _3040_ (.A(net74),
    .B(_0009_),
    .Y(_0947_));
 sg13g2_a21o_1 _3041_ (.A2(net77),
    .A1(_1240_),
    .B1(_0947_),
    .X(_0948_));
 sg13g2_inv_1 _3042_ (.Y(_0949_),
    .A(_0948_));
 sg13g2_a21oi_1 _3043_ (.A1(_0948_),
    .A2(net55),
    .Y(_0950_),
    .B1(net76));
 sg13g2_nand2_1 _3044_ (.Y(_0951_),
    .A(_0938_),
    .B(_1100_));
 sg13g2_nand2_1 _3045_ (.Y(_0952_),
    .A(_0939_),
    .B(\i_video.run_length[5] ));
 sg13g2_nand3_1 _3046_ (.B(_0951_),
    .C(_0952_),
    .A(net35),
    .Y(_0953_));
 sg13g2_nand2_1 _3047_ (.Y(_0954_),
    .A(net36),
    .B(_0949_));
 sg13g2_nand3_1 _3048_ (.B(_0954_),
    .C(net51),
    .A(_0953_),
    .Y(_0955_));
 sg13g2_a22oi_1 _3049_ (.Y(_0956_),
    .B1(_0950_),
    .B2(_0955_),
    .A2(_0949_),
    .A1(net75));
 sg13g2_nand2_1 _3050_ (.Y(_0957_),
    .A(_0956_),
    .B(net29));
 sg13g2_nand2_1 _3051_ (.Y(_0958_),
    .A(net28),
    .B(\i_video.run_length[5] ));
 sg13g2_nand3_1 _3052_ (.B(_0958_),
    .C(net81),
    .A(_0957_),
    .Y(_0220_));
 sg13g2_nor2_1 _3053_ (.A(net77),
    .B(_0010_),
    .Y(_0959_));
 sg13g2_a21o_1 _3054_ (.A2(net77),
    .A1(_1243_),
    .B1(_0959_),
    .X(_0960_));
 sg13g2_inv_1 _3055_ (.Y(_0961_),
    .A(_0960_));
 sg13g2_nand2_1 _3056_ (.Y(_0962_),
    .A(_0961_),
    .B(net75));
 sg13g2_nor2_1 _3057_ (.A(\i_video.run_length[6] ),
    .B(_0951_),
    .Y(_0963_));
 sg13g2_a21oi_1 _3058_ (.A1(_0938_),
    .A2(_1100_),
    .Y(_0964_),
    .B1(_0671_));
 sg13g2_nor3_1 _3059_ (.A(_0963_),
    .B(_0964_),
    .C(net36),
    .Y(_0965_));
 sg13g2_o21ai_1 _3060_ (.B1(net51),
    .Y(_0966_),
    .A1(_0960_),
    .A2(net35));
 sg13g2_a21oi_1 _3061_ (.A1(_0960_),
    .A2(_0673_),
    .Y(_0967_),
    .B1(_0691_));
 sg13g2_o21ai_1 _3062_ (.B1(_0967_),
    .Y(_0968_),
    .A1(_0965_),
    .A2(_0966_));
 sg13g2_nand3_1 _3063_ (.B(_0962_),
    .C(_0968_),
    .A(net29),
    .Y(_0969_));
 sg13g2_nand2_1 _3064_ (.Y(_0970_),
    .A(_0909_),
    .B(\i_video.run_length[6] ));
 sg13g2_nand3_1 _3065_ (.B(_0970_),
    .C(net81),
    .A(_0969_),
    .Y(_0221_));
 sg13g2_nor2_1 _3066_ (.A(net74),
    .B(_0011_),
    .Y(_0971_));
 sg13g2_a21o_1 _3067_ (.A2(net74),
    .A1(_1246_),
    .B1(_0971_),
    .X(_0972_));
 sg13g2_inv_1 _3068_ (.Y(_0973_),
    .A(_0972_));
 sg13g2_a21oi_1 _3069_ (.A1(_0972_),
    .A2(net55),
    .Y(_0974_),
    .B1(net76));
 sg13g2_nand2_1 _3070_ (.Y(_0975_),
    .A(_0963_),
    .B(_1101_));
 sg13g2_o21ai_1 _3071_ (.B1(\i_video.run_length[7] ),
    .Y(_0976_),
    .A1(\i_video.run_length[6] ),
    .A2(_0951_));
 sg13g2_nand3_1 _3072_ (.B(_0975_),
    .C(_0976_),
    .A(net35),
    .Y(_0977_));
 sg13g2_nand2_1 _3073_ (.Y(_0978_),
    .A(net36),
    .B(_0973_));
 sg13g2_nand3_1 _3074_ (.B(_0978_),
    .C(net51),
    .A(_0977_),
    .Y(_0979_));
 sg13g2_a22oi_1 _3075_ (.Y(_0980_),
    .B1(_0974_),
    .B2(_0979_),
    .A2(_0973_),
    .A1(net75));
 sg13g2_nand2_1 _3076_ (.Y(_0981_),
    .A(_0980_),
    .B(net29));
 sg13g2_nand2_1 _3077_ (.Y(_0982_),
    .A(net28),
    .B(\i_video.run_length[7] ));
 sg13g2_nand3_1 _3078_ (.B(_0982_),
    .C(_0838_),
    .A(_0981_),
    .Y(_0222_));
 sg13g2_nor2_1 _3079_ (.A(net74),
    .B(_0012_),
    .Y(_0983_));
 sg13g2_a21o_1 _3080_ (.A2(net74),
    .A1(_1249_),
    .B1(_0983_),
    .X(_0984_));
 sg13g2_inv_1 _3081_ (.Y(_0985_),
    .A(_0984_));
 sg13g2_a21oi_1 _3082_ (.A1(_0984_),
    .A2(net55),
    .Y(_0986_),
    .B1(net76));
 sg13g2_nor2_1 _3083_ (.A(_1080_),
    .B(_0975_),
    .Y(_0987_));
 sg13g2_inv_1 _3084_ (.Y(_0988_),
    .A(_0987_));
 sg13g2_nand2_1 _3085_ (.Y(_0989_),
    .A(_0975_),
    .B(_1080_));
 sg13g2_nand3_1 _3086_ (.B(_0988_),
    .C(_0989_),
    .A(net35),
    .Y(_0990_));
 sg13g2_nand2_1 _3087_ (.Y(_0991_),
    .A(_0683_),
    .B(_0985_));
 sg13g2_nand3_1 _3088_ (.B(_0991_),
    .C(net51),
    .A(_0990_),
    .Y(_0992_));
 sg13g2_a22oi_1 _3089_ (.Y(_0993_),
    .B1(_0986_),
    .B2(_0992_),
    .A2(_0985_),
    .A1(net75));
 sg13g2_nand2_1 _3090_ (.Y(_0994_),
    .A(_0993_),
    .B(net29));
 sg13g2_nand2_1 _3091_ (.Y(_0995_),
    .A(net28),
    .B(_1080_));
 sg13g2_nand3_1 _3092_ (.B(_0995_),
    .C(_0838_),
    .A(_0994_),
    .Y(_0223_));
 sg13g2_nor2_1 _3093_ (.A(_1207_),
    .B(_0013_),
    .Y(_0996_));
 sg13g2_a21o_1 _3094_ (.A2(_0895_),
    .A1(_1252_),
    .B1(_0996_),
    .X(_0997_));
 sg13g2_inv_1 _3095_ (.Y(_0998_),
    .A(_0997_));
 sg13g2_a21oi_1 _3096_ (.A1(_0997_),
    .A2(_0673_),
    .Y(_0999_),
    .B1(net76));
 sg13g2_nand2_1 _3097_ (.Y(_1000_),
    .A(_0988_),
    .B(_1082_));
 sg13g2_nand3_1 _3098_ (.B(_0674_),
    .C(_1000_),
    .A(net35),
    .Y(_1001_));
 sg13g2_nand2_1 _3099_ (.Y(_1002_),
    .A(_0683_),
    .B(_0998_));
 sg13g2_nand3_1 _3100_ (.B(_1002_),
    .C(_0760_),
    .A(_1001_),
    .Y(_1003_));
 sg13g2_a22oi_1 _3101_ (.Y(_1004_),
    .B1(_0999_),
    .B2(_1003_),
    .A2(_0998_),
    .A1(_0751_));
 sg13g2_nand2_1 _3102_ (.Y(_1005_),
    .A(_1004_),
    .B(_0906_));
 sg13g2_nand2_1 _3103_ (.Y(_1006_),
    .A(net28),
    .B(_1082_));
 sg13g2_nand3_1 _3104_ (.B(_1006_),
    .C(net82),
    .A(_1005_),
    .Y(_0224_));
 sg13g2_a21oi_1 _3105_ (.A1(_0704_),
    .A2(_1110_),
    .Y(_0225_),
    .B1(net67));
 sg13g2_nor2_1 _3106_ (.A(clknet_leaf_7_clk),
    .B(_1116_),
    .Y(\i_spi.spi_clk_out ));
 sg13g2_a21oi_1 _3107_ (.A1(_0782_),
    .A2(\i_spi.bits_remaining[1] ),
    .Y(_1007_),
    .B1(\i_spi.bits_remaining[2] ));
 sg13g2_nor2b_1 _3108_ (.A(_0786_),
    .B_N(\i_spi.bits_remaining[2] ),
    .Y(_1008_));
 sg13g2_o21ai_1 _3109_ (.B1(_0779_),
    .Y(_1009_),
    .A1(_1007_),
    .A2(_1008_));
 sg13g2_o21ai_1 _3110_ (.B1(_1009_),
    .Y(\i_spi.spi_mosi ),
    .A1(_1180_),
    .A2(_1122_));
 sg13g2_nor4_1 _3111_ (.A(_1026_),
    .B(\i_vga.timing_ver.counter[4] ),
    .C(\i_vga.timing_ver.counter[8] ),
    .D(\i_vga.timing_ver.counter[9] ),
    .Y(_1010_));
 sg13g2_nor4_1 _3112_ (.A(\i_vga.timing_ver.counter[3] ),
    .B(\i_vga.timing_ver.counter[2] ),
    .C(\i_vga.timing_ver.counter[7] ),
    .D(\i_vga.timing_ver.counter[6] ),
    .Y(_1011_));
 sg13g2_nand4_1 _3113_ (.B(_1011_),
    .C(_1021_),
    .A(_1010_),
    .Y(_1012_),
    .D(_1037_));
 sg13g2_nand2_1 _3114_ (.Y(_1013_),
    .A(_1012_),
    .B(_1030_));
 sg13g2_o21ai_1 _3115_ (.B1(_1013_),
    .Y(\i_vga.timing_ver.blank ),
    .A1(_1019_),
    .A2(_1012_));
 sg13g2_nand2_1 _3116_ (.Y(_1014_),
    .A(net82),
    .B(\i_spi.spi_data_oe[0] ));
 sg13g2_inv_1 _3117_ (.Y(net9),
    .A(_1014_));
 sg13g2_nor2_1 _3118_ (.A(_0735_),
    .B(_0698_),
    .Y(net16));
 sg13g2_nor2_1 _3119_ (.A(_0725_),
    .B(_0698_),
    .Y(net17));
 sg13g2_nor2_1 _3120_ (.A(_0715_),
    .B(_0698_),
    .Y(net18));
 sg13g2_nor2_1 _3121_ (.A(_0730_),
    .B(_0698_),
    .Y(net20));
 sg13g2_nor2_1 _3122_ (.A(_0720_),
    .B(_0698_),
    .Y(net21));
 sg13g2_nor2_1 _3123_ (.A(_0710_),
    .B(_0698_),
    .Y(net22));
 sg13g2_inv_1 _1722__1 (.Y(net300),
    .A(clknet_leaf_13_clk));
 sg13g2_tiehi _3139__91 (.L_HI(net91));
 sg13g2_buf_1 _3126_ (.A(rst_n),
    .X(net8));
 sg13g2_buf_1 _3127_ (.A(net85),
    .X(uio_oe[2]));
 sg13g2_buf_1 _3128_ (.A(rst_n),
    .X(net10));
 sg13g2_buf_1 _3129_ (.A(net86),
    .X(uio_oe[4]));
 sg13g2_buf_1 _3130_ (.A(net87),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3131_ (.A(rst_n),
    .X(net11));
 sg13g2_buf_1 _3132_ (.A(rst_n),
    .X(net12));
 sg13g2_buf_1 _3133_ (.A(\i_spi.spi_select ),
    .X(net13));
 sg13g2_buf_1 _3134_ (.A(\i_spi.spi_mosi ),
    .X(net14));
 sg13g2_buf_1 _3135_ (.A(net88),
    .X(uio_out[2]));
 sg13g2_buf_1 _3136_ (.A(\i_spi.spi_clk_out ),
    .X(net15));
 sg13g2_buf_1 _3137_ (.A(net89),
    .X(uio_out[4]));
 sg13g2_buf_1 _3138_ (.A(net90),
    .X(uio_out[5]));
 sg13g2_buf_1 _3139_ (.A(net91),
    .X(uio_out[6]));
 sg13g2_buf_1 _3140_ (.A(net92),
    .X(uio_out[7]));
 sg13g2_buf_1 _3141_ (.A(\i_vga.timing_ver.sync ),
    .X(net19));
 sg13g2_buf_1 _3142_ (.A(\i_vga.hsync ),
    .X(net23));
 sg13g2_dfrbp_1 \addr[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net93),
    .D(_0039_),
    .Q_N(_0037_),
    .Q(\addr[1] ));
 sg13g2_dfrbp_1 \addr[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net94),
    .D(_0040_),
    .Q_N(_0026_),
    .Q(\addr[11] ));
 sg13g2_dfrbp_1 \addr[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net95),
    .D(_0041_),
    .Q_N(_0027_),
    .Q(\addr[12] ));
 sg13g2_dfrbp_1 \addr[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net96),
    .D(_0042_),
    .Q_N(_0028_),
    .Q(\addr[13] ));
 sg13g2_dfrbp_1 \addr[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net97),
    .D(_0043_),
    .Q_N(_0029_),
    .Q(\addr[14] ));
 sg13g2_dfrbp_1 \addr[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net98),
    .D(_0044_),
    .Q_N(_0030_),
    .Q(\addr[15] ));
 sg13g2_dfrbp_1 \addr[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net99),
    .D(_0045_),
    .Q_N(_0031_),
    .Q(\addr[16] ));
 sg13g2_dfrbp_1 \addr[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net100),
    .D(_0046_),
    .Q_N(_0032_),
    .Q(\addr[17] ));
 sg13g2_dfrbp_1 \addr[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net101),
    .D(_0047_),
    .Q_N(_0033_),
    .Q(\addr[18] ));
 sg13g2_dfrbp_1 \addr[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net102),
    .D(_0048_),
    .Q_N(_1647_),
    .Q(\addr[19] ));
 sg13g2_dfrbp_1 \addr[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net103),
    .D(_0049_),
    .Q_N(_1646_),
    .Q(\addr[20] ));
 sg13g2_dfrbp_1 \addr[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net104),
    .D(_0050_),
    .Q_N(_1645_),
    .Q(\addr[2] ));
 sg13g2_dfrbp_1 \addr[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net105),
    .D(_0051_),
    .Q_N(_0034_),
    .Q(\addr[21] ));
 sg13g2_dfrbp_1 \addr[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net106),
    .D(_0052_),
    .Q_N(_0035_),
    .Q(\addr[22] ));
 sg13g2_dfrbp_1 \addr[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net107),
    .D(_0053_),
    .Q_N(_1644_),
    .Q(\addr[23] ));
 sg13g2_dfrbp_1 \addr[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net108),
    .D(_0054_),
    .Q_N(_1643_),
    .Q(\addr[3] ));
 sg13g2_dfrbp_1 \addr[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net109),
    .D(_0055_),
    .Q_N(_1642_),
    .Q(\addr[4] ));
 sg13g2_dfrbp_1 \addr[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net110),
    .D(_0056_),
    .Q_N(_1641_),
    .Q(\addr[5] ));
 sg13g2_dfrbp_1 \addr[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net111),
    .D(_0057_),
    .Q_N(_1640_),
    .Q(\addr[6] ));
 sg13g2_dfrbp_1 \addr[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net112),
    .D(_0058_),
    .Q_N(_0023_),
    .Q(\addr[7] ));
 sg13g2_dfrbp_1 \addr[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net113),
    .D(_0059_),
    .Q_N(_1639_),
    .Q(\addr[8] ));
 sg13g2_dfrbp_1 \addr[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net114),
    .D(_0060_),
    .Q_N(_0024_),
    .Q(\addr[9] ));
 sg13g2_dfrbp_1 \addr[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net115),
    .D(_0061_),
    .Q_N(_0025_),
    .Q(\addr[10] ));
 sg13g2_dfrbp_1 \addr_offset1[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net116),
    .D(_0062_),
    .Q_N(_1638_),
    .Q(\addr_offset1[1] ));
 sg13g2_dfrbp_1 \addr_offset1[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net117),
    .D(_0063_),
    .Q_N(_1637_),
    .Q(\addr_offset1[2] ));
 sg13g2_dfrbp_1 \addr_offset1[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net118),
    .D(_0064_),
    .Q_N(_1636_),
    .Q(\addr_offset1[3] ));
 sg13g2_dfrbp_1 \addr_offset1[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net119),
    .D(_0065_),
    .Q_N(_1635_),
    .Q(\addr_offset1[4] ));
 sg13g2_dfrbp_1 \addr_offset1[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net120),
    .D(_0066_),
    .Q_N(_1634_),
    .Q(\addr_offset1[5] ));
 sg13g2_dfrbp_1 \addr_offset1[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net121),
    .D(_0067_),
    .Q_N(_1633_),
    .Q(\addr_offset1[6] ));
 sg13g2_dfrbp_1 \addr_offset1[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net122),
    .D(_0068_),
    .Q_N(_1632_),
    .Q(\addr_offset1[7] ));
 sg13g2_dfrbp_1 \addr_offset1[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net123),
    .D(_0069_),
    .Q_N(_1631_),
    .Q(\addr_offset1[8] ));
 sg13g2_dfrbp_1 \addr_saved0[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net124),
    .D(_0070_),
    .Q_N(_1630_),
    .Q(\addr_saved0[1] ));
 sg13g2_dfrbp_1 \addr_saved0[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net125),
    .D(_0071_),
    .Q_N(_1629_),
    .Q(\addr_saved0[11] ));
 sg13g2_dfrbp_1 \addr_saved0[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net126),
    .D(_0072_),
    .Q_N(_1628_),
    .Q(\addr_saved0[12] ));
 sg13g2_dfrbp_1 \addr_saved0[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net127),
    .D(_0073_),
    .Q_N(_1627_),
    .Q(\addr_saved0[13] ));
 sg13g2_dfrbp_1 \addr_saved0[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net128),
    .D(_0074_),
    .Q_N(_1626_),
    .Q(\addr_saved0[14] ));
 sg13g2_dfrbp_1 \addr_saved0[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net129),
    .D(_0075_),
    .Q_N(_1625_),
    .Q(\addr_saved0[15] ));
 sg13g2_dfrbp_1 \addr_saved0[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net130),
    .D(_0076_),
    .Q_N(_1624_),
    .Q(\addr_saved0[16] ));
 sg13g2_dfrbp_1 \addr_saved0[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net131),
    .D(_0077_),
    .Q_N(_1623_),
    .Q(\addr_saved0[17] ));
 sg13g2_dfrbp_1 \addr_saved0[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net132),
    .D(_0078_),
    .Q_N(_1622_),
    .Q(\addr_saved0[18] ));
 sg13g2_dfrbp_1 \addr_saved0[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net133),
    .D(_0079_),
    .Q_N(_1621_),
    .Q(\addr_saved0[19] ));
 sg13g2_dfrbp_1 \addr_saved0[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net134),
    .D(_0080_),
    .Q_N(_1620_),
    .Q(\addr_saved0[20] ));
 sg13g2_dfrbp_1 \addr_saved0[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net135),
    .D(_0081_),
    .Q_N(_1619_),
    .Q(\addr_saved0[2] ));
 sg13g2_dfrbp_1 \addr_saved0[20]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net136),
    .D(_0082_),
    .Q_N(_1618_),
    .Q(\addr_saved0[21] ));
 sg13g2_dfrbp_1 \addr_saved0[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net137),
    .D(_0083_),
    .Q_N(_1617_),
    .Q(\addr_saved0[22] ));
 sg13g2_dfrbp_1 \addr_saved0[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net138),
    .D(_0084_),
    .Q_N(_1616_),
    .Q(\addr_saved0[23] ));
 sg13g2_dfrbp_1 \addr_saved0[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net139),
    .D(_0085_),
    .Q_N(_1615_),
    .Q(\addr_saved0[3] ));
 sg13g2_dfrbp_1 \addr_saved0[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net140),
    .D(_0086_),
    .Q_N(_1614_),
    .Q(\addr_saved0[4] ));
 sg13g2_dfrbp_1 \addr_saved0[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net141),
    .D(_0087_),
    .Q_N(_1613_),
    .Q(\addr_saved0[5] ));
 sg13g2_dfrbp_1 \addr_saved0[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net142),
    .D(_0088_),
    .Q_N(_1612_),
    .Q(\addr_saved0[6] ));
 sg13g2_dfrbp_1 \addr_saved0[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net143),
    .D(_0089_),
    .Q_N(_1611_),
    .Q(\addr_saved0[7] ));
 sg13g2_dfrbp_1 \addr_saved0[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net144),
    .D(_0090_),
    .Q_N(_1610_),
    .Q(\addr_saved0[8] ));
 sg13g2_dfrbp_1 \addr_saved0[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net145),
    .D(_0091_),
    .Q_N(_1609_),
    .Q(\addr_saved0[9] ));
 sg13g2_dfrbp_1 \addr_saved0[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net146),
    .D(_0092_),
    .Q_N(_1608_),
    .Q(\addr_saved0[10] ));
 sg13g2_dfrbp_1 \i_spi.addr[10]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net147),
    .D(_0093_),
    .Q_N(_1607_),
    .Q(\i_spi.addr[10] ));
 sg13g2_dfrbp_1 \i_spi.addr[11]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net148),
    .D(_0094_),
    .Q_N(_1606_),
    .Q(\i_spi.addr[11] ));
 sg13g2_dfrbp_1 \i_spi.addr[12]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net149),
    .D(_0095_),
    .Q_N(_1605_),
    .Q(\i_spi.addr[12] ));
 sg13g2_dfrbp_1 \i_spi.addr[13]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net150),
    .D(_0096_),
    .Q_N(_1604_),
    .Q(\i_spi.addr[13] ));
 sg13g2_dfrbp_1 \i_spi.addr[14]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net151),
    .D(_0097_),
    .Q_N(_1603_),
    .Q(\i_spi.addr[14] ));
 sg13g2_dfrbp_1 \i_spi.addr[15]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net152),
    .D(_0098_),
    .Q_N(_1602_),
    .Q(\i_spi.addr[15] ));
 sg13g2_dfrbp_1 \i_spi.addr[16]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net153),
    .D(_0099_),
    .Q_N(_1601_),
    .Q(\i_spi.addr[16] ));
 sg13g2_dfrbp_1 \i_spi.addr[17]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net154),
    .D(_0100_),
    .Q_N(_1600_),
    .Q(\i_spi.addr[17] ));
 sg13g2_dfrbp_1 \i_spi.addr[18]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net155),
    .D(_0101_),
    .Q_N(_1599_),
    .Q(\i_spi.addr[18] ));
 sg13g2_dfrbp_1 \i_spi.addr[19]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net156),
    .D(_0102_),
    .Q_N(_1598_),
    .Q(\i_spi.addr[19] ));
 sg13g2_dfrbp_1 \i_spi.addr[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net157),
    .D(_0103_),
    .Q_N(_1597_),
    .Q(\i_spi.addr[1] ));
 sg13g2_dfrbp_1 \i_spi.addr[20]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net158),
    .D(_0104_),
    .Q_N(_1596_),
    .Q(\i_spi.addr[20] ));
 sg13g2_dfrbp_1 \i_spi.addr[21]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net159),
    .D(_0105_),
    .Q_N(_1595_),
    .Q(\i_spi.addr[21] ));
 sg13g2_dfrbp_1 \i_spi.addr[22]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net160),
    .D(_0106_),
    .Q_N(_1594_),
    .Q(\i_spi.addr[22] ));
 sg13g2_dfrbp_1 \i_spi.addr[23]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net161),
    .D(_0107_),
    .Q_N(_1593_),
    .Q(\i_spi.addr[23] ));
 sg13g2_dfrbp_1 \i_spi.addr[2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net162),
    .D(_0108_),
    .Q_N(_1592_),
    .Q(\i_spi.addr[2] ));
 sg13g2_dfrbp_1 \i_spi.addr[3]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net163),
    .D(_0109_),
    .Q_N(_1591_),
    .Q(\i_spi.addr[3] ));
 sg13g2_dfrbp_1 \i_spi.addr[4]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net164),
    .D(_0110_),
    .Q_N(_1590_),
    .Q(\i_spi.addr[4] ));
 sg13g2_dfrbp_1 \i_spi.addr[5]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net165),
    .D(_0111_),
    .Q_N(_1589_),
    .Q(\i_spi.addr[5] ));
 sg13g2_dfrbp_1 \i_spi.addr[6]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net166),
    .D(_0112_),
    .Q_N(_1588_),
    .Q(\i_spi.addr[6] ));
 sg13g2_dfrbp_1 \i_spi.addr[7]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net167),
    .D(_0113_),
    .Q_N(_1587_),
    .Q(\i_spi.addr[7] ));
 sg13g2_dfrbp_1 \i_spi.addr[8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net168),
    .D(_0114_),
    .Q_N(_1586_),
    .Q(\i_spi.addr[8] ));
 sg13g2_dfrbp_1 \i_spi.addr[9]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net169),
    .D(_0115_),
    .Q_N(_1585_),
    .Q(\i_spi.addr[9] ));
 sg13g2_dfrbp_1 \i_spi.bits_remaining[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net170),
    .D(_0116_),
    .Q_N(_1584_),
    .Q(\i_spi.bits_remaining[0] ));
 sg13g2_dfrbp_1 \i_spi.bits_remaining[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net171),
    .D(_0117_),
    .Q_N(_1583_),
    .Q(\i_spi.bits_remaining[1] ));
 sg13g2_dfrbp_1 \i_spi.bits_remaining[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net172),
    .D(_0118_),
    .Q_N(_0002_),
    .Q(\i_spi.bits_remaining[2] ));
 sg13g2_dfrbp_1 \i_spi.bits_remaining[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net173),
    .D(_0119_),
    .Q_N(_1582_),
    .Q(\i_spi.bits_remaining[3] ));
 sg13g2_dfrbp_1 \i_spi.bits_remaining[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net174),
    .D(_0120_),
    .Q_N(_0021_),
    .Q(\i_spi.bits_remaining[4] ));
 sg13g2_dfrbp_1 \i_spi.data[0]$_DFFE_PN_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net175),
    .D(_0121_),
    .Q_N(_1581_),
    .Q(\i_spi.data[0] ));
 sg13g2_dfrbp_1 \i_spi.data[10]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net176),
    .D(_0122_),
    .Q_N(_1580_),
    .Q(\i_spi.data[10] ));
 sg13g2_dfrbp_1 \i_spi.data[11]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net177),
    .D(_0123_),
    .Q_N(_1579_),
    .Q(\i_spi.data[11] ));
 sg13g2_dfrbp_1 \i_spi.data[12]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net178),
    .D(_0124_),
    .Q_N(_1578_),
    .Q(\i_spi.data[12] ));
 sg13g2_dfrbp_1 \i_spi.data[13]$_DFFE_PN_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net179),
    .D(_0125_),
    .Q_N(_1577_),
    .Q(\i_spi.data[13] ));
 sg13g2_dfrbp_1 \i_spi.data[14]$_DFFE_PN_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net180),
    .D(_0126_),
    .Q_N(_1576_),
    .Q(\i_spi.data[14] ));
 sg13g2_dfrbp_1 \i_spi.data[15]$_DFFE_PN_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net181),
    .D(_0127_),
    .Q_N(_1575_),
    .Q(\i_spi.data[15] ));
 sg13g2_dfrbp_1 \i_spi.data[1]$_DFFE_PN_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net182),
    .D(_0128_),
    .Q_N(_1574_),
    .Q(\i_spi.data[1] ));
 sg13g2_dfrbp_1 \i_spi.data[2]$_DFFE_PN_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net183),
    .D(_0129_),
    .Q_N(_1573_),
    .Q(\i_spi.data[2] ));
 sg13g2_dfrbp_1 \i_spi.data[3]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net184),
    .D(_0130_),
    .Q_N(_1572_),
    .Q(\i_spi.data[3] ));
 sg13g2_dfrbp_1 \i_spi.data[4]$_DFFE_PN_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net185),
    .D(_0131_),
    .Q_N(_1571_),
    .Q(\i_spi.data[4] ));
 sg13g2_dfrbp_1 \i_spi.data[5]$_DFFE_PN_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net186),
    .D(_0132_),
    .Q_N(_1570_),
    .Q(\i_spi.data[5] ));
 sg13g2_dfrbp_1 \i_spi.data[6]$_DFFE_PN_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net187),
    .D(_0133_),
    .Q_N(_1569_),
    .Q(\i_spi.data[6] ));
 sg13g2_dfrbp_1 \i_spi.data[7]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net188),
    .D(_0134_),
    .Q_N(_1568_),
    .Q(\i_spi.data[7] ));
 sg13g2_dfrbp_1 \i_spi.data[8]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net189),
    .D(_0135_),
    .Q_N(_1567_),
    .Q(\i_spi.data[8] ));
 sg13g2_dfrbp_1 \i_spi.data[9]$_DFFE_PN_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net190),
    .D(_0136_),
    .Q_N(_1566_),
    .Q(\i_spi.data[9] ));
 sg13g2_dfrbp_1 \i_spi.fsm_state[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net191),
    .D(_0137_),
    .Q_N(_1565_),
    .Q(\i_spi.fsm_state[0] ));
 sg13g2_dfrbp_1 \i_spi.fsm_state[1]$_SDFFE_PP1P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net192),
    .D(_0138_),
    .Q_N(_1564_),
    .Q(\i_spi.fsm_state[1] ));
 sg13g2_dfrbp_1 \i_spi.fsm_state[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net193),
    .D(_0139_),
    .Q_N(_0019_),
    .Q(\i_spi.fsm_state[2] ));
 sg13g2_dfrbp_1 \i_spi.spi_data_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net194),
    .D(_0140_),
    .Q_N(_1563_),
    .Q(\i_spi.spi_data_oe[0] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_n[0]$_DFF_N_  (.CLK(net307),
    .RESET_B(net195),
    .D(net4),
    .Q_N(_1562_),
    .Q(\i_spi.spi_miso_buf_n[0] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_n[1]$_DFF_N_  (.CLK(net306),
    .RESET_B(net196),
    .D(net5),
    .Q_N(_1561_),
    .Q(\i_spi.spi_miso_buf_n[1] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_n[2]$_DFF_N_  (.CLK(net305),
    .RESET_B(net197),
    .D(net6),
    .Q_N(_1560_),
    .Q(\i_spi.spi_miso_buf_n[2] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_n[3]$_DFF_N_  (.CLK(net304),
    .RESET_B(net198),
    .D(net7),
    .Q_N(_1559_),
    .Q(\i_spi.spi_miso_buf_n[3] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_n[4]$_DFF_N_  (.CLK(net303),
    .RESET_B(net199),
    .D(\i_spi.spi_miso_buf_n[0] ),
    .Q_N(_1558_),
    .Q(\i_spi.spi_miso_buf_n[4] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_n[5]$_DFF_N_  (.CLK(net302),
    .RESET_B(net200),
    .D(\i_spi.spi_miso_buf_n[1] ),
    .Q_N(_1557_),
    .Q(\i_spi.spi_miso_buf_n[5] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_n[6]$_DFF_N_  (.CLK(net301),
    .RESET_B(net201),
    .D(\i_spi.spi_miso_buf_n[2] ),
    .Q_N(_1556_),
    .Q(\i_spi.spi_miso_buf_n[6] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_n[7]$_DFF_N_  (.CLK(net300),
    .RESET_B(net202),
    .D(\i_spi.spi_miso_buf_n[3] ),
    .Q_N(_1648_),
    .Q(\i_spi.spi_miso_buf_n[7] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_p[0]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net203),
    .D(net4),
    .Q_N(_1649_),
    .Q(\i_spi.spi_miso_buf_p[0] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_p[1]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net204),
    .D(net5),
    .Q_N(_1650_),
    .Q(\i_spi.spi_miso_buf_p[1] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_p[2]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net205),
    .D(net6),
    .Q_N(_1651_),
    .Q(\i_spi.spi_miso_buf_p[2] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_p[3]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net206),
    .D(net7),
    .Q_N(_1652_),
    .Q(\i_spi.spi_miso_buf_p[3] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_p[4]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net207),
    .D(\i_spi.spi_miso_buf_p[0] ),
    .Q_N(_1653_),
    .Q(\i_spi.spi_miso_buf_p[4] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_p[5]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net208),
    .D(\i_spi.spi_miso_buf_p[1] ),
    .Q_N(_1654_),
    .Q(\i_spi.spi_miso_buf_p[5] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_p[6]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net209),
    .D(\i_spi.spi_miso_buf_p[2] ),
    .Q_N(_1655_),
    .Q(\i_spi.spi_miso_buf_p[6] ));
 sg13g2_dfrbp_1 \i_spi.spi_miso_buf_p[7]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net210),
    .D(\i_spi.spi_miso_buf_p[3] ),
    .Q_N(_1555_),
    .Q(\i_spi.spi_miso_buf_p[7] ));
 sg13g2_dfrbp_1 \i_spi_buf.empty$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net211),
    .D(_0141_),
    .Q_N(_0022_),
    .Q(\i_spi_buf.empty ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[0]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net212),
    .D(_0142_),
    .Q_N(_1554_),
    .Q(\i_spi_buf.fifo[0] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[10]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net213),
    .D(_0143_),
    .Q_N(_0008_),
    .Q(\i_spi_buf.fifo[10] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[11]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net214),
    .D(_0144_),
    .Q_N(_0009_),
    .Q(\i_spi_buf.fifo[11] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[12]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net215),
    .D(_0145_),
    .Q_N(_0010_),
    .Q(\i_spi_buf.fifo[12] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[13]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net216),
    .D(_0146_),
    .Q_N(_0011_),
    .Q(\i_spi_buf.fifo[13] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[14]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net217),
    .D(_0147_),
    .Q_N(_0012_),
    .Q(\i_spi_buf.fifo[14] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[15]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net218),
    .D(_0148_),
    .Q_N(_0013_),
    .Q(\i_spi_buf.fifo[15] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net219),
    .D(_0149_),
    .Q_N(_1553_),
    .Q(\i_spi_buf.fifo[1] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[2]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net220),
    .D(_0150_),
    .Q_N(_1552_),
    .Q(\i_spi_buf.fifo[2] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net221),
    .D(_0151_),
    .Q_N(_1551_),
    .Q(\i_spi_buf.fifo[3] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[4]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net222),
    .D(_0152_),
    .Q_N(_1550_),
    .Q(\i_spi_buf.fifo[4] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[5]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net223),
    .D(_0153_),
    .Q_N(_1549_),
    .Q(\i_spi_buf.fifo[5] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[6]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net224),
    .D(_0154_),
    .Q_N(_0004_),
    .Q(\i_spi_buf.fifo[6] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[7]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net225),
    .D(_0155_),
    .Q_N(_0005_),
    .Q(\i_spi_buf.fifo[7] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[8]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net226),
    .D(_0156_),
    .Q_N(_0006_),
    .Q(\i_spi_buf.fifo[8] ));
 sg13g2_dfrbp_1 \i_spi_buf.fifo[9]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net227),
    .D(_0157_),
    .Q_N(_0007_),
    .Q(\i_spi_buf.fifo[9] ));
 sg13g2_dfrbp_1 \i_spi_buf0.empty$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net228),
    .D(_0158_),
    .Q_N(_1548_),
    .Q(\i_spi_buf.prev_empty ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net229),
    .D(_0159_),
    .Q_N(_1547_),
    .Q(\i_spi_buf0.fifo[0] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[10]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net230),
    .D(_0160_),
    .Q_N(_1546_),
    .Q(\i_spi_buf0.fifo[10] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[11]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net231),
    .D(_0161_),
    .Q_N(_1545_),
    .Q(\i_spi_buf0.fifo[11] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[12]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net232),
    .D(_0162_),
    .Q_N(_1544_),
    .Q(\i_spi_buf0.fifo[12] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[13]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net233),
    .D(_0163_),
    .Q_N(_1543_),
    .Q(\i_spi_buf0.fifo[13] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[14]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net234),
    .D(_0164_),
    .Q_N(_1542_),
    .Q(\i_spi_buf0.fifo[14] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[15]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net235),
    .D(_0165_),
    .Q_N(_1541_),
    .Q(\i_spi_buf0.fifo[15] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[1]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net236),
    .D(_0166_),
    .Q_N(_1540_),
    .Q(\i_spi_buf0.fifo[1] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[2]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net237),
    .D(_0167_),
    .Q_N(_1539_),
    .Q(\i_spi_buf0.fifo[2] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[3]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net238),
    .D(_0168_),
    .Q_N(_1538_),
    .Q(\i_spi_buf0.fifo[3] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[4]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net239),
    .D(_0169_),
    .Q_N(_1537_),
    .Q(\i_spi_buf0.fifo[4] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[5]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net240),
    .D(_0170_),
    .Q_N(_1536_),
    .Q(\i_spi_buf0.fifo[5] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[6]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net241),
    .D(_0171_),
    .Q_N(_1535_),
    .Q(\i_spi_buf0.fifo[6] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[7]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net242),
    .D(_0172_),
    .Q_N(_1534_),
    .Q(\i_spi_buf0.fifo[7] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[8]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net243),
    .D(_0173_),
    .Q_N(_1533_),
    .Q(\i_spi_buf0.fifo[8] ));
 sg13g2_dfrbp_1 \i_spi_buf0.fifo[9]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net244),
    .D(_0174_),
    .Q_N(_1532_),
    .Q(\i_spi_buf0.fifo[9] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[0]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net245),
    .D(_0175_),
    .Q_N(_0036_),
    .Q(\i_vga.timing_hor.counter[0] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[10]$_SDFF_PP1_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net246),
    .D(_0176_),
    .Q_N(_0015_),
    .Q(\i_vga.timing_hor.counter[10] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[1]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net247),
    .D(_0177_),
    .Q_N(_1531_),
    .Q(\i_vga.timing_hor.counter[1] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[2]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net248),
    .D(_0178_),
    .Q_N(_1530_),
    .Q(\i_vga.timing_hor.counter[2] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[3]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net249),
    .D(_0179_),
    .Q_N(_1529_),
    .Q(\i_vga.timing_hor.counter[3] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[4]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net250),
    .D(_0180_),
    .Q_N(_0014_),
    .Q(\i_vga.timing_hor.counter[4] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[5]$_SDFF_PP1_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net251),
    .D(_0181_),
    .Q_N(_1528_),
    .Q(\i_vga.timing_hor.counter[5] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[6]$_SDFF_PP1_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net252),
    .D(_0182_),
    .Q_N(_1527_),
    .Q(\i_vga.timing_hor.counter[6] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[7]$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net253),
    .D(_0183_),
    .Q_N(_1526_),
    .Q(\i_vga.timing_hor.counter[7] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[8]$_SDFF_PP1_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net254),
    .D(_0184_),
    .Q_N(_1525_),
    .Q(\i_vga.timing_hor.counter[8] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[9]$_SDFF_PP1_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net255),
    .D(_0185_),
    .Q_N(_1656_),
    .Q(\i_vga.timing_hor.counter[9] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.sync$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net256),
    .D(_0000_),
    .Q_N(_1524_),
    .Q(\i_vga.hsync ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[0]$_SDFFE_PN1N_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net257),
    .D(_0186_),
    .Q_N(_1523_),
    .Q(\i_vga.timing_ver.counter[0] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[10]$_SDFFE_PN1N_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net258),
    .D(_0187_),
    .Q_N(_0017_),
    .Q(\i_vga.timing_ver.counter[10] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[1]$_SDFFE_PN1N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net259),
    .D(_0188_),
    .Q_N(_1522_),
    .Q(\i_vga.timing_ver.counter[1] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[2]$_SDFFE_PN0N_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net260),
    .D(_0189_),
    .Q_N(_1521_),
    .Q(\i_vga.timing_ver.counter[2] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[3]$_SDFFE_PN0N_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net261),
    .D(_0190_),
    .Q_N(_1520_),
    .Q(\i_vga.timing_ver.counter[3] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[4]$_SDFFE_PN1N_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net262),
    .D(_0191_),
    .Q_N(_1519_),
    .Q(\i_vga.timing_ver.counter[4] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[5]$_SDFFE_PN0N_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net263),
    .D(_0192_),
    .Q_N(_1518_),
    .Q(\i_vga.timing_ver.counter[5] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[6]$_SDFFE_PN1N_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net264),
    .D(_0193_),
    .Q_N(_1517_),
    .Q(\i_vga.timing_ver.counter[6] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[7]$_SDFFE_PN1N_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net265),
    .D(_0194_),
    .Q_N(_1516_),
    .Q(\i_vga.timing_ver.counter[7] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[8]$_SDFFE_PN1N_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net266),
    .D(_0195_),
    .Q_N(_1515_),
    .Q(\i_vga.timing_ver.counter[8] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[9]$_SDFFE_PN1N_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net267),
    .D(_0196_),
    .Q_N(_1657_),
    .Q(\i_vga.timing_ver.counter[9] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.sync$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net268),
    .D(_0001_),
    .Q_N(_1658_),
    .Q(\i_vga.timing_ver.sync ));
 sg13g2_dfrbp_1 \i_vga.vblank$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net269),
    .D(\i_vga.timing_ver.blank ),
    .Q_N(_1514_),
    .Q(\i_vga.vblank ));
 sg13g2_dfrbp_1 \i_video.clear_addr$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net270),
    .D(_0197_),
    .Q_N(_1513_),
    .Q(clear_addr));
 sg13g2_dfrbp_1 \i_video.colour[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net271),
    .D(_0198_),
    .Q_N(_1512_),
    .Q(\i_video.colour[0] ));
 sg13g2_dfrbp_1 \i_video.colour[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net272),
    .D(_0199_),
    .Q_N(_1511_),
    .Q(\i_video.colour[1] ));
 sg13g2_dfrbp_1 \i_video.colour[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net273),
    .D(_0200_),
    .Q_N(_1510_),
    .Q(\i_video.colour[2] ));
 sg13g2_dfrbp_1 \i_video.colour[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net274),
    .D(_0201_),
    .Q_N(_1509_),
    .Q(\i_video.colour[3] ));
 sg13g2_dfrbp_1 \i_video.colour[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net275),
    .D(_0202_),
    .Q_N(_1508_),
    .Q(\i_video.colour[4] ));
 sg13g2_dfrbp_1 \i_video.colour[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net276),
    .D(_0203_),
    .Q_N(_1507_),
    .Q(\i_video.colour[5] ));
 sg13g2_dfrbp_1 \i_video.frame_counter$_SDFFE_PP1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net277),
    .D(_0204_),
    .Q_N(_0016_),
    .Q(\i_video.frame_counter ));
 sg13g2_dfrbp_1 \i_video.read_next_r$_SDFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net278),
    .D(_0205_),
    .Q_N(_1506_),
    .Q(\i_video.read_next_r ));
 sg13g2_dfrbp_1 \i_video.repeat_count[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net279),
    .D(_0206_),
    .Q_N(_0003_),
    .Q(\i_video.repeat_count[0] ));
 sg13g2_dfrbp_1 \i_video.repeat_count[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net280),
    .D(_0207_),
    .Q_N(_1505_),
    .Q(\i_video.repeat_count[1] ));
 sg13g2_dfrbp_1 \i_video.repeat_count[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net281),
    .D(_0208_),
    .Q_N(_1504_),
    .Q(\i_video.repeat_count[2] ));
 sg13g2_dfrbp_1 \i_video.repeat_count[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net282),
    .D(_0209_),
    .Q_N(_1503_),
    .Q(\i_video.repeat_count[3] ));
 sg13g2_dfrbp_1 \i_video.repeat_count[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net283),
    .D(_0210_),
    .Q_N(_1502_),
    .Q(\i_video.repeat_count[4] ));
 sg13g2_dfrbp_1 \i_video.repeat_count[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net284),
    .D(_0211_),
    .Q_N(_1501_),
    .Q(\i_video.repeat_count[5] ));
 sg13g2_dfrbp_1 \i_video.repeat_count[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net285),
    .D(_0212_),
    .Q_N(_1500_),
    .Q(\i_video.repeat_count[6] ));
 sg13g2_dfrbp_1 \i_video.repeat_count[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net286),
    .D(_0213_),
    .Q_N(_1499_),
    .Q(\i_video.repeat_count[7] ));
 sg13g2_dfrbp_1 \i_video.repeat_count[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net287),
    .D(_0214_),
    .Q_N(_1498_),
    .Q(\i_video.repeat_count[8] ));
 sg13g2_dfrbp_1 \i_video.run_length[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net288),
    .D(_0215_),
    .Q_N(_1497_),
    .Q(\i_video.run_length[0] ));
 sg13g2_dfrbp_1 \i_video.run_length[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net289),
    .D(_0216_),
    .Q_N(_1496_),
    .Q(\i_video.run_length[1] ));
 sg13g2_dfrbp_1 \i_video.run_length[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net290),
    .D(_0217_),
    .Q_N(_1495_),
    .Q(\i_video.run_length[2] ));
 sg13g2_dfrbp_1 \i_video.run_length[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net291),
    .D(_0218_),
    .Q_N(_1494_),
    .Q(\i_video.run_length[3] ));
 sg13g2_dfrbp_1 \i_video.run_length[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net292),
    .D(_0219_),
    .Q_N(_1493_),
    .Q(\i_video.run_length[4] ));
 sg13g2_dfrbp_1 \i_video.run_length[5]$_SDFFE_PN1P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net293),
    .D(_0220_),
    .Q_N(_1492_),
    .Q(\i_video.run_length[5] ));
 sg13g2_dfrbp_1 \i_video.run_length[6]$_SDFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net294),
    .D(_0221_),
    .Q_N(_1491_),
    .Q(\i_video.run_length[6] ));
 sg13g2_dfrbp_1 \i_video.run_length[7]$_SDFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net295),
    .D(_0222_),
    .Q_N(_1490_),
    .Q(\i_video.run_length[7] ));
 sg13g2_dfrbp_1 \i_video.run_length[8]$_SDFFE_PN1P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net296),
    .D(_0223_),
    .Q_N(_1489_),
    .Q(\i_video.run_length[8] ));
 sg13g2_dfrbp_1 \i_video.run_length[9]$_SDFFE_PN1P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net297),
    .D(_0224_),
    .Q_N(_1488_),
    .Q(\i_video.run_length[9] ));
 sg13g2_dfrbp_1 \i_video.start$_SDFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net298),
    .D(_0225_),
    .Q_N(_0018_),
    .Q(\i_video.start ));
 sg13g2_dfrbp_1 \spi_started$_SDFFE_PP0N_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net299),
    .D(_0226_),
    .Q_N(_0020_),
    .Q(spi_started));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[1]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[2]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[5]),
    .X(net7));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[0]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[1]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[3]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[6]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_oe[7]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[0]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[1]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[3]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[0]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[1]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[2]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[3]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[4]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[5]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[6]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout24 (.A(_0706_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1302_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_1297_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1296_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0909_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0906_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1237_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1226_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0331_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0282_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1358_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0744_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0683_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1454_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1167_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1161_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1126_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1115_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0555_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0531_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0529_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1452_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0527_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1451_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1449_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1372_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1363_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0760_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_1439_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1362_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1122_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0745_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0708_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1361_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1136_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1129_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1128_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0855_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1324_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1322_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1315_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1355_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1215_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0803_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0663_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0556_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0506_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_1455_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_1354_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_1228_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0895_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0751_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0739_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0662_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0629_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1234_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1227_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0838_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0784_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0691_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_1107_),
    .X(net84));
 sg13g2_tielo _3127__85 (.L_LO(net85));
 sg13g2_tielo _3129__86 (.L_LO(net86));
 sg13g2_tielo _3130__87 (.L_LO(net87));
 sg13g2_tielo _3135__88 (.L_LO(net88));
 sg13g2_tielo _3137__89 (.L_LO(net89));
 sg13g2_tielo _3138__90 (.L_LO(net90));
 sg13g2_tiehi _3140__92 (.L_HI(net92));
 sg13g2_tiehi \addr[0]$_SDFFE_PP0P__93  (.L_HI(net93));
 sg13g2_tiehi \addr[10]$_SDFFE_PP0P__94  (.L_HI(net94));
 sg13g2_tiehi \addr[11]$_SDFFE_PP0P__95  (.L_HI(net95));
 sg13g2_tiehi \addr[12]$_SDFFE_PP0P__96  (.L_HI(net96));
 sg13g2_tiehi \addr[13]$_SDFFE_PP0P__97  (.L_HI(net97));
 sg13g2_tiehi \addr[14]$_SDFFE_PP0P__98  (.L_HI(net98));
 sg13g2_tiehi \addr[15]$_SDFFE_PP0P__99  (.L_HI(net99));
 sg13g2_tiehi \addr[16]$_SDFFE_PP0P__100  (.L_HI(net100));
 sg13g2_tiehi \addr[17]$_SDFFE_PP0P__101  (.L_HI(net101));
 sg13g2_tiehi \addr[18]$_SDFFE_PP0P__102  (.L_HI(net102));
 sg13g2_tiehi \addr[19]$_SDFFE_PP0P__103  (.L_HI(net103));
 sg13g2_tiehi \addr[1]$_SDFFE_PP0P__104  (.L_HI(net104));
 sg13g2_tiehi \addr[20]$_SDFFE_PP0P__105  (.L_HI(net105));
 sg13g2_tiehi \addr[21]$_SDFFE_PP0P__106  (.L_HI(net106));
 sg13g2_tiehi \addr[22]$_SDFFE_PP0P__107  (.L_HI(net107));
 sg13g2_tiehi \addr[2]$_SDFFE_PP0P__108  (.L_HI(net108));
 sg13g2_tiehi \addr[3]$_SDFFE_PP0P__109  (.L_HI(net109));
 sg13g2_tiehi \addr[4]$_SDFFE_PP0P__110  (.L_HI(net110));
 sg13g2_tiehi \addr[5]$_SDFFE_PP0P__111  (.L_HI(net111));
 sg13g2_tiehi \addr[6]$_SDFFE_PP0P__112  (.L_HI(net112));
 sg13g2_tiehi \addr[7]$_SDFFE_PP0P__113  (.L_HI(net113));
 sg13g2_tiehi \addr[8]$_SDFFE_PP0P__114  (.L_HI(net114));
 sg13g2_tiehi \addr[9]$_SDFFE_PP0P__115  (.L_HI(net115));
 sg13g2_tiehi \addr_offset1[0]$_SDFFE_PP0P__116  (.L_HI(net116));
 sg13g2_tiehi \addr_offset1[1]$_SDFFE_PP0P__117  (.L_HI(net117));
 sg13g2_tiehi \addr_offset1[2]$_SDFFE_PP0P__118  (.L_HI(net118));
 sg13g2_tiehi \addr_offset1[3]$_SDFFE_PP0P__119  (.L_HI(net119));
 sg13g2_tiehi \addr_offset1[4]$_SDFFE_PP0P__120  (.L_HI(net120));
 sg13g2_tiehi \addr_offset1[5]$_SDFFE_PP0P__121  (.L_HI(net121));
 sg13g2_tiehi \addr_offset1[6]$_SDFFE_PP0P__122  (.L_HI(net122));
 sg13g2_tiehi \addr_offset1[7]$_SDFFE_PP0P__123  (.L_HI(net123));
 sg13g2_tiehi \addr_saved0[0]$_SDFFE_PP0P__124  (.L_HI(net124));
 sg13g2_tiehi \addr_saved0[10]$_SDFFE_PP0P__125  (.L_HI(net125));
 sg13g2_tiehi \addr_saved0[11]$_SDFFE_PP0P__126  (.L_HI(net126));
 sg13g2_tiehi \addr_saved0[12]$_SDFFE_PP0P__127  (.L_HI(net127));
 sg13g2_tiehi \addr_saved0[13]$_SDFFE_PP0P__128  (.L_HI(net128));
 sg13g2_tiehi \addr_saved0[14]$_SDFFE_PP0P__129  (.L_HI(net129));
 sg13g2_tiehi \addr_saved0[15]$_SDFFE_PP0P__130  (.L_HI(net130));
 sg13g2_tiehi \addr_saved0[16]$_SDFFE_PP0P__131  (.L_HI(net131));
 sg13g2_tiehi \addr_saved0[17]$_SDFFE_PP0P__132  (.L_HI(net132));
 sg13g2_tiehi \addr_saved0[18]$_SDFFE_PP0P__133  (.L_HI(net133));
 sg13g2_tiehi \addr_saved0[19]$_SDFFE_PP0P__134  (.L_HI(net134));
 sg13g2_tiehi \addr_saved0[1]$_SDFFE_PP0P__135  (.L_HI(net135));
 sg13g2_tiehi \addr_saved0[20]$_SDFFE_PP0P__136  (.L_HI(net136));
 sg13g2_tiehi \addr_saved0[21]$_SDFFE_PP0P__137  (.L_HI(net137));
 sg13g2_tiehi \addr_saved0[22]$_SDFFE_PP0P__138  (.L_HI(net138));
 sg13g2_tiehi \addr_saved0[2]$_SDFFE_PP0P__139  (.L_HI(net139));
 sg13g2_tiehi \addr_saved0[3]$_SDFFE_PP0P__140  (.L_HI(net140));
 sg13g2_tiehi \addr_saved0[4]$_SDFFE_PP0P__141  (.L_HI(net141));
 sg13g2_tiehi \addr_saved0[5]$_SDFFE_PP0P__142  (.L_HI(net142));
 sg13g2_tiehi \addr_saved0[6]$_SDFFE_PP0P__143  (.L_HI(net143));
 sg13g2_tiehi \addr_saved0[7]$_SDFFE_PP0P__144  (.L_HI(net144));
 sg13g2_tiehi \addr_saved0[8]$_SDFFE_PP0P__145  (.L_HI(net145));
 sg13g2_tiehi \addr_saved0[9]$_SDFFE_PP0P__146  (.L_HI(net146));
 sg13g2_tiehi \i_spi.addr[10]$_DFFE_PP__147  (.L_HI(net147));
 sg13g2_tiehi \i_spi.addr[11]$_DFFE_PP__148  (.L_HI(net148));
 sg13g2_tiehi \i_spi.addr[12]$_DFFE_PP__149  (.L_HI(net149));
 sg13g2_tiehi \i_spi.addr[13]$_DFFE_PP__150  (.L_HI(net150));
 sg13g2_tiehi \i_spi.addr[14]$_DFFE_PP__151  (.L_HI(net151));
 sg13g2_tiehi \i_spi.addr[15]$_DFFE_PP__152  (.L_HI(net152));
 sg13g2_tiehi \i_spi.addr[16]$_DFFE_PP__153  (.L_HI(net153));
 sg13g2_tiehi \i_spi.addr[17]$_DFFE_PP__154  (.L_HI(net154));
 sg13g2_tiehi \i_spi.addr[18]$_DFFE_PP__155  (.L_HI(net155));
 sg13g2_tiehi \i_spi.addr[19]$_DFFE_PP__156  (.L_HI(net156));
 sg13g2_tiehi \i_spi.addr[1]$_SDFFCE_PN0P__157  (.L_HI(net157));
 sg13g2_tiehi \i_spi.addr[20]$_DFFE_PP__158  (.L_HI(net158));
 sg13g2_tiehi \i_spi.addr[21]$_DFFE_PP__159  (.L_HI(net159));
 sg13g2_tiehi \i_spi.addr[22]$_DFFE_PP__160  (.L_HI(net160));
 sg13g2_tiehi \i_spi.addr[23]$_DFFE_PP__161  (.L_HI(net161));
 sg13g2_tiehi \i_spi.addr[2]$_DFFE_PP__162  (.L_HI(net162));
 sg13g2_tiehi \i_spi.addr[3]$_DFFE_PP__163  (.L_HI(net163));
 sg13g2_tiehi \i_spi.addr[4]$_DFFE_PP__164  (.L_HI(net164));
 sg13g2_tiehi \i_spi.addr[5]$_DFFE_PP__165  (.L_HI(net165));
 sg13g2_tiehi \i_spi.addr[6]$_DFFE_PP__166  (.L_HI(net166));
 sg13g2_tiehi \i_spi.addr[7]$_DFFE_PP__167  (.L_HI(net167));
 sg13g2_tiehi \i_spi.addr[8]$_DFFE_PP__168  (.L_HI(net168));
 sg13g2_tiehi \i_spi.addr[9]$_DFFE_PP__169  (.L_HI(net169));
 sg13g2_tiehi \i_spi.bits_remaining[0]$_SDFFE_PN0P__170  (.L_HI(net170));
 sg13g2_tiehi \i_spi.bits_remaining[1]$_SDFFE_PN0P__171  (.L_HI(net171));
 sg13g2_tiehi \i_spi.bits_remaining[2]$_SDFFE_PN0P__172  (.L_HI(net172));
 sg13g2_tiehi \i_spi.bits_remaining[3]$_SDFFE_PN0P__173  (.L_HI(net173));
 sg13g2_tiehi \i_spi.bits_remaining[4]$_SDFFE_PN0P__174  (.L_HI(net174));
 sg13g2_tiehi \i_spi.data[0]$_DFFE_PN__175  (.L_HI(net175));
 sg13g2_tiehi \i_spi.data[10]$_DFFE_PN__176  (.L_HI(net176));
 sg13g2_tiehi \i_spi.data[11]$_DFFE_PN__177  (.L_HI(net177));
 sg13g2_tiehi \i_spi.data[12]$_DFFE_PN__178  (.L_HI(net178));
 sg13g2_tiehi \i_spi.data[13]$_DFFE_PN__179  (.L_HI(net179));
 sg13g2_tiehi \i_spi.data[14]$_DFFE_PN__180  (.L_HI(net180));
 sg13g2_tiehi \i_spi.data[15]$_DFFE_PN__181  (.L_HI(net181));
 sg13g2_tiehi \i_spi.data[1]$_DFFE_PN__182  (.L_HI(net182));
 sg13g2_tiehi \i_spi.data[2]$_DFFE_PN__183  (.L_HI(net183));
 sg13g2_tiehi \i_spi.data[3]$_DFFE_PN__184  (.L_HI(net184));
 sg13g2_tiehi \i_spi.data[4]$_DFFE_PN__185  (.L_HI(net185));
 sg13g2_tiehi \i_spi.data[5]$_DFFE_PN__186  (.L_HI(net186));
 sg13g2_tiehi \i_spi.data[6]$_DFFE_PN__187  (.L_HI(net187));
 sg13g2_tiehi \i_spi.data[7]$_DFFE_PN__188  (.L_HI(net188));
 sg13g2_tiehi \i_spi.data[8]$_DFFE_PN__189  (.L_HI(net189));
 sg13g2_tiehi \i_spi.data[9]$_DFFE_PN__190  (.L_HI(net190));
 sg13g2_tiehi \i_spi.fsm_state[0]$_SDFFE_PP1P__191  (.L_HI(net191));
 sg13g2_tiehi \i_spi.fsm_state[1]$_SDFFE_PP1P__192  (.L_HI(net192));
 sg13g2_tiehi \i_spi.fsm_state[2]$_SDFFE_PP0P__193  (.L_HI(net193));
 sg13g2_tiehi \i_spi.spi_data_oe[0]$_SDFFE_PN0P__194  (.L_HI(net194));
 sg13g2_tiehi \i_spi.spi_miso_buf_n[0]$_DFF_N__195  (.L_HI(net195));
 sg13g2_tiehi \i_spi.spi_miso_buf_n[1]$_DFF_N__196  (.L_HI(net196));
 sg13g2_tiehi \i_spi.spi_miso_buf_n[2]$_DFF_N__197  (.L_HI(net197));
 sg13g2_tiehi \i_spi.spi_miso_buf_n[3]$_DFF_N__198  (.L_HI(net198));
 sg13g2_tiehi \i_spi.spi_miso_buf_n[4]$_DFF_N__199  (.L_HI(net199));
 sg13g2_tiehi \i_spi.spi_miso_buf_n[5]$_DFF_N__200  (.L_HI(net200));
 sg13g2_tiehi \i_spi.spi_miso_buf_n[6]$_DFF_N__201  (.L_HI(net201));
 sg13g2_tiehi \i_spi.spi_miso_buf_n[7]$_DFF_N__202  (.L_HI(net202));
 sg13g2_tiehi \i_spi.spi_miso_buf_p[0]$_DFF_P__203  (.L_HI(net203));
 sg13g2_tiehi \i_spi.spi_miso_buf_p[1]$_DFF_P__204  (.L_HI(net204));
 sg13g2_tiehi \i_spi.spi_miso_buf_p[2]$_DFF_P__205  (.L_HI(net205));
 sg13g2_tiehi \i_spi.spi_miso_buf_p[3]$_DFF_P__206  (.L_HI(net206));
 sg13g2_tiehi \i_spi.spi_miso_buf_p[4]$_DFF_P__207  (.L_HI(net207));
 sg13g2_tiehi \i_spi.spi_miso_buf_p[5]$_DFF_P__208  (.L_HI(net208));
 sg13g2_tiehi \i_spi.spi_miso_buf_p[6]$_DFF_P__209  (.L_HI(net209));
 sg13g2_tiehi \i_spi.spi_miso_buf_p[7]$_DFF_P__210  (.L_HI(net210));
 sg13g2_tiehi \i_spi_buf.empty$_SDFFE_PN0P__211  (.L_HI(net211));
 sg13g2_tiehi \i_spi_buf.fifo[0]$_DFFE_PP__212  (.L_HI(net212));
 sg13g2_tiehi \i_spi_buf.fifo[10]$_DFFE_PP__213  (.L_HI(net213));
 sg13g2_tiehi \i_spi_buf.fifo[11]$_DFFE_PP__214  (.L_HI(net214));
 sg13g2_tiehi \i_spi_buf.fifo[12]$_DFFE_PP__215  (.L_HI(net215));
 sg13g2_tiehi \i_spi_buf.fifo[13]$_DFFE_PP__216  (.L_HI(net216));
 sg13g2_tiehi \i_spi_buf.fifo[14]$_DFFE_PP__217  (.L_HI(net217));
 sg13g2_tiehi \i_spi_buf.fifo[15]$_DFFE_PP__218  (.L_HI(net218));
 sg13g2_tiehi \i_spi_buf.fifo[1]$_DFFE_PP__219  (.L_HI(net219));
 sg13g2_tiehi \i_spi_buf.fifo[2]$_DFFE_PP__220  (.L_HI(net220));
 sg13g2_tiehi \i_spi_buf.fifo[3]$_DFFE_PP__221  (.L_HI(net221));
 sg13g2_tiehi \i_spi_buf.fifo[4]$_DFFE_PP__222  (.L_HI(net222));
 sg13g2_tiehi \i_spi_buf.fifo[5]$_DFFE_PP__223  (.L_HI(net223));
 sg13g2_tiehi \i_spi_buf.fifo[6]$_DFFE_PP__224  (.L_HI(net224));
 sg13g2_tiehi \i_spi_buf.fifo[7]$_DFFE_PP__225  (.L_HI(net225));
 sg13g2_tiehi \i_spi_buf.fifo[8]$_DFFE_PP__226  (.L_HI(net226));
 sg13g2_tiehi \i_spi_buf.fifo[9]$_DFFE_PP__227  (.L_HI(net227));
 sg13g2_tiehi \i_spi_buf0.empty$_SDFFE_PN0P__228  (.L_HI(net228));
 sg13g2_tiehi \i_spi_buf0.fifo[0]$_DFFE_PP__229  (.L_HI(net229));
 sg13g2_tiehi \i_spi_buf0.fifo[10]$_DFFE_PP__230  (.L_HI(net230));
 sg13g2_tiehi \i_spi_buf0.fifo[11]$_DFFE_PP__231  (.L_HI(net231));
 sg13g2_tiehi \i_spi_buf0.fifo[12]$_DFFE_PP__232  (.L_HI(net232));
 sg13g2_tiehi \i_spi_buf0.fifo[13]$_DFFE_PP__233  (.L_HI(net233));
 sg13g2_tiehi \i_spi_buf0.fifo[14]$_DFFE_PP__234  (.L_HI(net234));
 sg13g2_tiehi \i_spi_buf0.fifo[15]$_DFFE_PP__235  (.L_HI(net235));
 sg13g2_tiehi \i_spi_buf0.fifo[1]$_DFFE_PP__236  (.L_HI(net236));
 sg13g2_tiehi \i_spi_buf0.fifo[2]$_DFFE_PP__237  (.L_HI(net237));
 sg13g2_tiehi \i_spi_buf0.fifo[3]$_DFFE_PP__238  (.L_HI(net238));
 sg13g2_tiehi \i_spi_buf0.fifo[4]$_DFFE_PP__239  (.L_HI(net239));
 sg13g2_tiehi \i_spi_buf0.fifo[5]$_DFFE_PP__240  (.L_HI(net240));
 sg13g2_tiehi \i_spi_buf0.fifo[6]$_DFFE_PP__241  (.L_HI(net241));
 sg13g2_tiehi \i_spi_buf0.fifo[7]$_DFFE_PP__242  (.L_HI(net242));
 sg13g2_tiehi \i_spi_buf0.fifo[8]$_DFFE_PP__243  (.L_HI(net243));
 sg13g2_tiehi \i_spi_buf0.fifo[9]$_DFFE_PP__244  (.L_HI(net244));
 sg13g2_tiehi \i_vga.timing_hor.counter[0]$_SDFF_PP0__245  (.L_HI(net245));
 sg13g2_tiehi \i_vga.timing_hor.counter[10]$_SDFF_PP1__246  (.L_HI(net246));
 sg13g2_tiehi \i_vga.timing_hor.counter[1]$_SDFF_PP0__247  (.L_HI(net247));
 sg13g2_tiehi \i_vga.timing_hor.counter[2]$_SDFF_PP0__248  (.L_HI(net248));
 sg13g2_tiehi \i_vga.timing_hor.counter[3]$_SDFF_PP0__249  (.L_HI(net249));
 sg13g2_tiehi \i_vga.timing_hor.counter[4]$_SDFF_PP0__250  (.L_HI(net250));
 sg13g2_tiehi \i_vga.timing_hor.counter[5]$_SDFF_PP1__251  (.L_HI(net251));
 sg13g2_tiehi \i_vga.timing_hor.counter[6]$_SDFF_PP1__252  (.L_HI(net252));
 sg13g2_tiehi \i_vga.timing_hor.counter[7]$_SDFF_PP0__253  (.L_HI(net253));
 sg13g2_tiehi \i_vga.timing_hor.counter[8]$_SDFF_PP1__254  (.L_HI(net254));
 sg13g2_tiehi \i_vga.timing_hor.counter[9]$_SDFF_PP1__255  (.L_HI(net255));
 sg13g2_tiehi \i_vga.timing_hor.sync$_DFF_P__256  (.L_HI(net256));
 sg13g2_tiehi \i_vga.timing_ver.counter[0]$_SDFFE_PN1N__257  (.L_HI(net257));
 sg13g2_tiehi \i_vga.timing_ver.counter[10]$_SDFFE_PN1N__258  (.L_HI(net258));
 sg13g2_tiehi \i_vga.timing_ver.counter[1]$_SDFFE_PN1N__259  (.L_HI(net259));
 sg13g2_tiehi \i_vga.timing_ver.counter[2]$_SDFFE_PN0N__260  (.L_HI(net260));
 sg13g2_tiehi \i_vga.timing_ver.counter[3]$_SDFFE_PN0N__261  (.L_HI(net261));
 sg13g2_tiehi \i_vga.timing_ver.counter[4]$_SDFFE_PN1N__262  (.L_HI(net262));
 sg13g2_tiehi \i_vga.timing_ver.counter[5]$_SDFFE_PN0N__263  (.L_HI(net263));
 sg13g2_tiehi \i_vga.timing_ver.counter[6]$_SDFFE_PN1N__264  (.L_HI(net264));
 sg13g2_tiehi \i_vga.timing_ver.counter[7]$_SDFFE_PN1N__265  (.L_HI(net265));
 sg13g2_tiehi \i_vga.timing_ver.counter[8]$_SDFFE_PN1N__266  (.L_HI(net266));
 sg13g2_tiehi \i_vga.timing_ver.counter[9]$_SDFFE_PN1N__267  (.L_HI(net267));
 sg13g2_tiehi \i_vga.timing_ver.sync$_DFF_P__268  (.L_HI(net268));
 sg13g2_tiehi \i_vga.vblank$_DFF_P__269  (.L_HI(net269));
 sg13g2_tiehi \i_video.clear_addr$_SDFFE_PN0P__270  (.L_HI(net270));
 sg13g2_tiehi \i_video.colour[0]$_SDFFE_PP0P__271  (.L_HI(net271));
 sg13g2_tiehi \i_video.colour[1]$_SDFFE_PP0P__272  (.L_HI(net272));
 sg13g2_tiehi \i_video.colour[2]$_SDFFE_PP0P__273  (.L_HI(net273));
 sg13g2_tiehi \i_video.colour[3]$_SDFFE_PP0P__274  (.L_HI(net274));
 sg13g2_tiehi \i_video.colour[4]$_SDFFE_PP0P__275  (.L_HI(net275));
 sg13g2_tiehi \i_video.colour[5]$_SDFFE_PP0P__276  (.L_HI(net276));
 sg13g2_tiehi \i_video.frame_counter$_SDFFE_PP1P__277  (.L_HI(net277));
 sg13g2_tiehi \i_video.read_next_r$_SDFF_PP0__278  (.L_HI(net278));
 sg13g2_tiehi \i_video.repeat_count[0]$_SDFFE_PN0P__279  (.L_HI(net279));
 sg13g2_tiehi \i_video.repeat_count[1]$_SDFFE_PN0P__280  (.L_HI(net280));
 sg13g2_tiehi \i_video.repeat_count[2]$_SDFFE_PN0P__281  (.L_HI(net281));
 sg13g2_tiehi \i_video.repeat_count[3]$_SDFFE_PN0P__282  (.L_HI(net282));
 sg13g2_tiehi \i_video.repeat_count[4]$_SDFFE_PN0P__283  (.L_HI(net283));
 sg13g2_tiehi \i_video.repeat_count[5]$_SDFFE_PN0P__284  (.L_HI(net284));
 sg13g2_tiehi \i_video.repeat_count[6]$_SDFFE_PN0P__285  (.L_HI(net285));
 sg13g2_tiehi \i_video.repeat_count[7]$_SDFFE_PN0P__286  (.L_HI(net286));
 sg13g2_tiehi \i_video.repeat_count[8]$_SDFFE_PN0P__287  (.L_HI(net287));
 sg13g2_tiehi \i_video.run_length[0]$_SDFFE_PP1P__288  (.L_HI(net288));
 sg13g2_tiehi \i_video.run_length[1]$_SDFFE_PN1P__289  (.L_HI(net289));
 sg13g2_tiehi \i_video.run_length[2]$_SDFFE_PN1P__290  (.L_HI(net290));
 sg13g2_tiehi \i_video.run_length[3]$_SDFFE_PN1P__291  (.L_HI(net291));
 sg13g2_tiehi \i_video.run_length[4]$_SDFFE_PN1P__292  (.L_HI(net292));
 sg13g2_tiehi \i_video.run_length[5]$_SDFFE_PN1P__293  (.L_HI(net293));
 sg13g2_tiehi \i_video.run_length[6]$_SDFFE_PN1P__294  (.L_HI(net294));
 sg13g2_tiehi \i_video.run_length[7]$_SDFFE_PN1P__295  (.L_HI(net295));
 sg13g2_tiehi \i_video.run_length[8]$_SDFFE_PN1P__296  (.L_HI(net296));
 sg13g2_tiehi \i_video.run_length[9]$_SDFFE_PN1P__297  (.L_HI(net297));
 sg13g2_tiehi \i_video.start$_SDFF_PN0__298  (.L_HI(net298));
 sg13g2_tiehi \spi_started$_SDFFE_PP0N__299  (.L_HI(net299));
 sg13g2_inv_1 net255_2 (.Y(net301),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 net255_3 (.Y(net302),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 net255_4 (.Y(net303),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 net255_5 (.Y(net304),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 net255_6 (.Y(net305),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 net255_7 (.Y(net306),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 net255_8 (.Y(net307),
    .A(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_7__leaf_clk));
 sg13g2_buf_16 clkload3 (.A(clknet_leaf_28_clk));
 sg13g2_buf_16 clkload4 (.A(clknet_leaf_25_clk));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_5_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_leaf_8_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_23_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_18_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_20_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_4 FILLER_0_63 ();
 sg13g2_fill_2 FILLER_0_67 ();
 sg13g2_fill_2 FILLER_0_95 ();
 sg13g2_fill_1 FILLER_0_97 ();
 sg13g2_fill_2 FILLER_0_124 ();
 sg13g2_fill_1 FILLER_0_126 ();
 sg13g2_fill_2 FILLER_0_130 ();
 sg13g2_decap_4 FILLER_0_144 ();
 sg13g2_fill_1 FILLER_0_148 ();
 sg13g2_decap_8 FILLER_0_158 ();
 sg13g2_fill_1 FILLER_0_165 ();
 sg13g2_fill_2 FILLER_0_174 ();
 sg13g2_fill_1 FILLER_0_202 ();
 sg13g2_fill_2 FILLER_0_210 ();
 sg13g2_fill_1 FILLER_0_212 ();
 sg13g2_fill_2 FILLER_0_244 ();
 sg13g2_decap_4 FILLER_0_251 ();
 sg13g2_fill_1 FILLER_0_255 ();
 sg13g2_fill_2 FILLER_0_291 ();
 sg13g2_decap_4 FILLER_0_319 ();
 sg13g2_fill_1 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_0_332 ();
 sg13g2_decap_8 FILLER_0_339 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_8 FILLER_0_403 ();
 sg13g2_decap_8 FILLER_0_410 ();
 sg13g2_decap_8 FILLER_0_417 ();
 sg13g2_decap_4 FILLER_0_424 ();
 sg13g2_fill_2 FILLER_0_428 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_4 FILLER_1_56 ();
 sg13g2_fill_1 FILLER_1_60 ();
 sg13g2_decap_8 FILLER_1_65 ();
 sg13g2_fill_2 FILLER_1_72 ();
 sg13g2_fill_1 FILLER_1_74 ();
 sg13g2_fill_2 FILLER_1_98 ();
 sg13g2_fill_2 FILLER_1_105 ();
 sg13g2_fill_1 FILLER_1_107 ();
 sg13g2_fill_2 FILLER_1_112 ();
 sg13g2_fill_1 FILLER_1_114 ();
 sg13g2_fill_2 FILLER_1_120 ();
 sg13g2_fill_1 FILLER_1_127 ();
 sg13g2_fill_1 FILLER_1_182 ();
 sg13g2_fill_1 FILLER_1_187 ();
 sg13g2_fill_1 FILLER_1_228 ();
 sg13g2_fill_1 FILLER_1_234 ();
 sg13g2_fill_1 FILLER_1_239 ();
 sg13g2_fill_1 FILLER_1_266 ();
 sg13g2_fill_1 FILLER_1_271 ();
 sg13g2_fill_1 FILLER_1_278 ();
 sg13g2_fill_2 FILLER_1_314 ();
 sg13g2_decap_8 FILLER_1_397 ();
 sg13g2_decap_8 FILLER_1_404 ();
 sg13g2_decap_8 FILLER_1_411 ();
 sg13g2_decap_8 FILLER_1_418 ();
 sg13g2_decap_4 FILLER_1_425 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_4 FILLER_2_49 ();
 sg13g2_fill_1 FILLER_2_53 ();
 sg13g2_fill_2 FILLER_2_90 ();
 sg13g2_fill_1 FILLER_2_92 ();
 sg13g2_fill_1 FILLER_2_127 ();
 sg13g2_fill_1 FILLER_2_148 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_fill_2 FILLER_2_161 ();
 sg13g2_fill_1 FILLER_2_193 ();
 sg13g2_decap_4 FILLER_2_199 ();
 sg13g2_fill_1 FILLER_2_208 ();
 sg13g2_fill_1 FILLER_2_213 ();
 sg13g2_fill_2 FILLER_2_222 ();
 sg13g2_fill_1 FILLER_2_224 ();
 sg13g2_fill_2 FILLER_2_230 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_fill_2 FILLER_2_245 ();
 sg13g2_fill_1 FILLER_2_251 ();
 sg13g2_fill_2 FILLER_2_257 ();
 sg13g2_fill_1 FILLER_2_324 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_8 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_2_412 ();
 sg13g2_decap_8 FILLER_2_419 ();
 sg13g2_decap_4 FILLER_2_426 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_4 FILLER_3_42 ();
 sg13g2_fill_1 FILLER_3_46 ();
 sg13g2_decap_4 FILLER_3_117 ();
 sg13g2_fill_1 FILLER_3_121 ();
 sg13g2_fill_2 FILLER_3_127 ();
 sg13g2_fill_1 FILLER_3_150 ();
 sg13g2_fill_1 FILLER_3_166 ();
 sg13g2_fill_1 FILLER_3_188 ();
 sg13g2_fill_1 FILLER_3_197 ();
 sg13g2_decap_4 FILLER_3_217 ();
 sg13g2_fill_2 FILLER_3_221 ();
 sg13g2_fill_1 FILLER_3_243 ();
 sg13g2_decap_4 FILLER_3_260 ();
 sg13g2_fill_2 FILLER_3_264 ();
 sg13g2_fill_2 FILLER_3_296 ();
 sg13g2_fill_1 FILLER_3_328 ();
 sg13g2_fill_2 FILLER_3_334 ();
 sg13g2_fill_2 FILLER_3_341 ();
 sg13g2_fill_2 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_fill_2 FILLER_4_35 ();
 sg13g2_fill_1 FILLER_4_37 ();
 sg13g2_fill_2 FILLER_4_63 ();
 sg13g2_fill_1 FILLER_4_77 ();
 sg13g2_fill_2 FILLER_4_144 ();
 sg13g2_fill_2 FILLER_4_166 ();
 sg13g2_fill_1 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_181 ();
 sg13g2_fill_2 FILLER_4_201 ();
 sg13g2_fill_2 FILLER_4_222 ();
 sg13g2_fill_1 FILLER_4_224 ();
 sg13g2_fill_2 FILLER_4_243 ();
 sg13g2_decap_4 FILLER_4_266 ();
 sg13g2_fill_1 FILLER_4_270 ();
 sg13g2_fill_1 FILLER_4_274 ();
 sg13g2_fill_1 FILLER_4_280 ();
 sg13g2_fill_1 FILLER_4_285 ();
 sg13g2_fill_2 FILLER_4_309 ();
 sg13g2_fill_2 FILLER_4_315 ();
 sg13g2_fill_2 FILLER_4_356 ();
 sg13g2_fill_1 FILLER_4_358 ();
 sg13g2_fill_2 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_4 FILLER_5_35 ();
 sg13g2_fill_1 FILLER_5_70 ();
 sg13g2_fill_1 FILLER_5_85 ();
 sg13g2_fill_2 FILLER_5_90 ();
 sg13g2_fill_2 FILLER_5_97 ();
 sg13g2_fill_2 FILLER_5_125 ();
 sg13g2_decap_4 FILLER_5_151 ();
 sg13g2_fill_1 FILLER_5_158 ();
 sg13g2_fill_1 FILLER_5_198 ();
 sg13g2_fill_2 FILLER_5_204 ();
 sg13g2_fill_1 FILLER_5_211 ();
 sg13g2_decap_4 FILLER_5_247 ();
 sg13g2_fill_2 FILLER_5_256 ();
 sg13g2_fill_2 FILLER_5_263 ();
 sg13g2_fill_1 FILLER_5_265 ();
 sg13g2_fill_2 FILLER_5_271 ();
 sg13g2_fill_1 FILLER_5_273 ();
 sg13g2_fill_1 FILLER_5_279 ();
 sg13g2_fill_1 FILLER_5_324 ();
 sg13g2_decap_4 FILLER_5_329 ();
 sg13g2_fill_1 FILLER_5_333 ();
 sg13g2_fill_1 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_decap_8 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_5_415 ();
 sg13g2_decap_8 FILLER_5_422 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_4 FILLER_6_21 ();
 sg13g2_fill_2 FILLER_6_25 ();
 sg13g2_fill_1 FILLER_6_53 ();
 sg13g2_fill_1 FILLER_6_59 ();
 sg13g2_fill_1 FILLER_6_93 ();
 sg13g2_fill_1 FILLER_6_99 ();
 sg13g2_fill_1 FILLER_6_105 ();
 sg13g2_fill_2 FILLER_6_110 ();
 sg13g2_decap_4 FILLER_6_116 ();
 sg13g2_fill_1 FILLER_6_127 ();
 sg13g2_fill_2 FILLER_6_135 ();
 sg13g2_fill_1 FILLER_6_137 ();
 sg13g2_fill_2 FILLER_6_150 ();
 sg13g2_fill_1 FILLER_6_165 ();
 sg13g2_fill_1 FILLER_6_175 ();
 sg13g2_decap_4 FILLER_6_184 ();
 sg13g2_fill_1 FILLER_6_188 ();
 sg13g2_fill_1 FILLER_6_209 ();
 sg13g2_decap_4 FILLER_6_214 ();
 sg13g2_fill_2 FILLER_6_222 ();
 sg13g2_fill_1 FILLER_6_252 ();
 sg13g2_fill_1 FILLER_6_266 ();
 sg13g2_fill_2 FILLER_6_272 ();
 sg13g2_fill_1 FILLER_6_274 ();
 sg13g2_fill_2 FILLER_6_377 ();
 sg13g2_fill_1 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_4 FILLER_7_21 ();
 sg13g2_fill_2 FILLER_7_25 ();
 sg13g2_decap_4 FILLER_7_100 ();
 sg13g2_fill_2 FILLER_7_150 ();
 sg13g2_fill_2 FILLER_7_163 ();
 sg13g2_fill_1 FILLER_7_165 ();
 sg13g2_fill_2 FILLER_7_171 ();
 sg13g2_fill_2 FILLER_7_188 ();
 sg13g2_fill_1 FILLER_7_203 ();
 sg13g2_decap_4 FILLER_7_221 ();
 sg13g2_fill_1 FILLER_7_225 ();
 sg13g2_fill_2 FILLER_7_231 ();
 sg13g2_fill_2 FILLER_7_236 ();
 sg13g2_fill_1 FILLER_7_247 ();
 sg13g2_fill_1 FILLER_7_282 ();
 sg13g2_fill_2 FILLER_7_310 ();
 sg13g2_fill_2 FILLER_7_316 ();
 sg13g2_fill_1 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_323 ();
 sg13g2_fill_1 FILLER_7_330 ();
 sg13g2_fill_1 FILLER_7_340 ();
 sg13g2_fill_2 FILLER_7_345 ();
 sg13g2_fill_2 FILLER_7_351 ();
 sg13g2_fill_2 FILLER_7_358 ();
 sg13g2_fill_1 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_391 ();
 sg13g2_decap_8 FILLER_7_398 ();
 sg13g2_decap_8 FILLER_7_405 ();
 sg13g2_decap_8 FILLER_7_412 ();
 sg13g2_decap_8 FILLER_7_419 ();
 sg13g2_decap_4 FILLER_7_426 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_4 FILLER_8_14 ();
 sg13g2_decap_4 FILLER_8_99 ();
 sg13g2_fill_1 FILLER_8_111 ();
 sg13g2_fill_1 FILLER_8_116 ();
 sg13g2_fill_2 FILLER_8_127 ();
 sg13g2_fill_1 FILLER_8_129 ();
 sg13g2_fill_1 FILLER_8_135 ();
 sg13g2_decap_4 FILLER_8_143 ();
 sg13g2_fill_2 FILLER_8_163 ();
 sg13g2_fill_1 FILLER_8_165 ();
 sg13g2_fill_1 FILLER_8_179 ();
 sg13g2_decap_8 FILLER_8_192 ();
 sg13g2_decap_8 FILLER_8_209 ();
 sg13g2_decap_8 FILLER_8_216 ();
 sg13g2_fill_1 FILLER_8_223 ();
 sg13g2_decap_8 FILLER_8_263 ();
 sg13g2_decap_4 FILLER_8_275 ();
 sg13g2_fill_2 FILLER_8_279 ();
 sg13g2_fill_2 FILLER_8_285 ();
 sg13g2_fill_1 FILLER_8_287 ();
 sg13g2_fill_1 FILLER_8_328 ();
 sg13g2_fill_2 FILLER_8_359 ();
 sg13g2_fill_1 FILLER_8_361 ();
 sg13g2_fill_1 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_4 FILLER_8_424 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_4 FILLER_9_14 ();
 sg13g2_fill_2 FILLER_9_18 ();
 sg13g2_fill_1 FILLER_9_98 ();
 sg13g2_fill_1 FILLER_9_104 ();
 sg13g2_fill_1 FILLER_9_182 ();
 sg13g2_fill_2 FILLER_9_186 ();
 sg13g2_fill_1 FILLER_9_188 ();
 sg13g2_fill_1 FILLER_9_198 ();
 sg13g2_fill_1 FILLER_9_218 ();
 sg13g2_fill_2 FILLER_9_226 ();
 sg13g2_fill_1 FILLER_9_246 ();
 sg13g2_fill_1 FILLER_9_255 ();
 sg13g2_fill_1 FILLER_9_262 ();
 sg13g2_fill_1 FILLER_9_267 ();
 sg13g2_fill_1 FILLER_9_274 ();
 sg13g2_fill_1 FILLER_9_280 ();
 sg13g2_fill_2 FILLER_9_286 ();
 sg13g2_fill_1 FILLER_9_288 ();
 sg13g2_fill_1 FILLER_9_304 ();
 sg13g2_fill_2 FILLER_9_309 ();
 sg13g2_fill_1 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_8 FILLER_9_404 ();
 sg13g2_decap_8 FILLER_9_411 ();
 sg13g2_decap_8 FILLER_9_418 ();
 sg13g2_decap_4 FILLER_9_425 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_67 ();
 sg13g2_fill_1 FILLER_10_84 ();
 sg13g2_fill_1 FILLER_10_95 ();
 sg13g2_fill_1 FILLER_10_101 ();
 sg13g2_fill_1 FILLER_10_107 ();
 sg13g2_fill_2 FILLER_10_124 ();
 sg13g2_fill_2 FILLER_10_154 ();
 sg13g2_fill_1 FILLER_10_192 ();
 sg13g2_fill_1 FILLER_10_196 ();
 sg13g2_fill_2 FILLER_10_201 ();
 sg13g2_fill_2 FILLER_10_207 ();
 sg13g2_fill_1 FILLER_10_218 ();
 sg13g2_fill_1 FILLER_10_279 ();
 sg13g2_fill_2 FILLER_10_319 ();
 sg13g2_fill_1 FILLER_10_321 ();
 sg13g2_fill_1 FILLER_10_334 ();
 sg13g2_fill_2 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_10_409 ();
 sg13g2_decap_8 FILLER_10_416 ();
 sg13g2_decap_8 FILLER_10_423 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_66 ();
 sg13g2_fill_1 FILLER_11_75 ();
 sg13g2_fill_1 FILLER_11_81 ();
 sg13g2_fill_1 FILLER_11_91 ();
 sg13g2_fill_1 FILLER_11_126 ();
 sg13g2_decap_4 FILLER_11_142 ();
 sg13g2_fill_2 FILLER_11_162 ();
 sg13g2_fill_2 FILLER_11_168 ();
 sg13g2_fill_1 FILLER_11_174 ();
 sg13g2_fill_1 FILLER_11_205 ();
 sg13g2_fill_1 FILLER_11_216 ();
 sg13g2_fill_1 FILLER_11_221 ();
 sg13g2_fill_2 FILLER_11_232 ();
 sg13g2_fill_1 FILLER_11_234 ();
 sg13g2_fill_1 FILLER_11_273 ();
 sg13g2_fill_2 FILLER_11_295 ();
 sg13g2_fill_1 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_302 ();
 sg13g2_decap_4 FILLER_11_312 ();
 sg13g2_fill_1 FILLER_11_316 ();
 sg13g2_fill_1 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_8 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_11_412 ();
 sg13g2_decap_8 FILLER_11_419 ();
 sg13g2_decap_4 FILLER_11_426 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_110 ();
 sg13g2_fill_2 FILLER_12_174 ();
 sg13g2_fill_2 FILLER_12_194 ();
 sg13g2_fill_2 FILLER_12_217 ();
 sg13g2_decap_4 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_233 ();
 sg13g2_decap_8 FILLER_12_240 ();
 sg13g2_fill_2 FILLER_12_247 ();
 sg13g2_fill_1 FILLER_12_249 ();
 sg13g2_fill_1 FILLER_12_254 ();
 sg13g2_decap_4 FILLER_12_264 ();
 sg13g2_fill_2 FILLER_12_268 ();
 sg13g2_fill_1 FILLER_12_275 ();
 sg13g2_fill_1 FILLER_12_338 ();
 sg13g2_fill_1 FILLER_12_349 ();
 sg13g2_fill_2 FILLER_12_354 ();
 sg13g2_fill_1 FILLER_12_361 ();
 sg13g2_fill_2 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_8 FILLER_12_404 ();
 sg13g2_decap_8 FILLER_12_411 ();
 sg13g2_decap_8 FILLER_12_418 ();
 sg13g2_decap_4 FILLER_12_425 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_4 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_32 ();
 sg13g2_fill_1 FILLER_13_59 ();
 sg13g2_fill_1 FILLER_13_98 ();
 sg13g2_fill_2 FILLER_13_103 ();
 sg13g2_fill_2 FILLER_13_110 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_fill_2 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_13_170 ();
 sg13g2_fill_1 FILLER_13_180 ();
 sg13g2_decap_4 FILLER_13_190 ();
 sg13g2_fill_1 FILLER_13_194 ();
 sg13g2_fill_2 FILLER_13_215 ();
 sg13g2_fill_1 FILLER_13_217 ();
 sg13g2_fill_1 FILLER_13_244 ();
 sg13g2_fill_1 FILLER_13_274 ();
 sg13g2_fill_1 FILLER_13_311 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_13_409 ();
 sg13g2_decap_8 FILLER_13_416 ();
 sg13g2_decap_8 FILLER_13_423 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_35 ();
 sg13g2_fill_1 FILLER_14_37 ();
 sg13g2_fill_1 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_47 ();
 sg13g2_decap_8 FILLER_14_54 ();
 sg13g2_decap_4 FILLER_14_61 ();
 sg13g2_fill_1 FILLER_14_65 ();
 sg13g2_fill_2 FILLER_14_81 ();
 sg13g2_fill_2 FILLER_14_125 ();
 sg13g2_fill_1 FILLER_14_146 ();
 sg13g2_fill_1 FILLER_14_152 ();
 sg13g2_fill_1 FILLER_14_160 ();
 sg13g2_fill_1 FILLER_14_165 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_185 ();
 sg13g2_fill_2 FILLER_14_191 ();
 sg13g2_fill_2 FILLER_14_205 ();
 sg13g2_fill_2 FILLER_14_220 ();
 sg13g2_fill_1 FILLER_14_222 ();
 sg13g2_fill_2 FILLER_14_249 ();
 sg13g2_fill_1 FILLER_14_251 ();
 sg13g2_fill_2 FILLER_14_256 ();
 sg13g2_fill_1 FILLER_14_262 ();
 sg13g2_fill_1 FILLER_14_294 ();
 sg13g2_fill_2 FILLER_14_304 ();
 sg13g2_fill_2 FILLER_14_323 ();
 sg13g2_fill_1 FILLER_14_329 ();
 sg13g2_fill_1 FILLER_14_335 ();
 sg13g2_fill_2 FILLER_14_340 ();
 sg13g2_fill_2 FILLER_14_384 ();
 sg13g2_decap_4 FILLER_14_390 ();
 sg13g2_fill_1 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_fill_2 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_23 ();
 sg13g2_fill_1 FILLER_15_28 ();
 sg13g2_fill_1 FILLER_15_80 ();
 sg13g2_fill_1 FILLER_15_86 ();
 sg13g2_fill_1 FILLER_15_92 ();
 sg13g2_fill_2 FILLER_15_110 ();
 sg13g2_fill_2 FILLER_15_124 ();
 sg13g2_fill_1 FILLER_15_126 ();
 sg13g2_fill_1 FILLER_15_138 ();
 sg13g2_fill_1 FILLER_15_144 ();
 sg13g2_fill_2 FILLER_15_152 ();
 sg13g2_fill_1 FILLER_15_157 ();
 sg13g2_fill_2 FILLER_15_195 ();
 sg13g2_fill_1 FILLER_15_197 ();
 sg13g2_fill_1 FILLER_15_206 ();
 sg13g2_fill_1 FILLER_15_264 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_293 ();
 sg13g2_fill_2 FILLER_15_298 ();
 sg13g2_fill_1 FILLER_15_393 ();
 sg13g2_decap_4 FILLER_15_425 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_fill_1 FILLER_16_28 ();
 sg13g2_fill_1 FILLER_16_64 ();
 sg13g2_fill_1 FILLER_16_70 ();
 sg13g2_fill_2 FILLER_16_86 ();
 sg13g2_fill_1 FILLER_16_88 ();
 sg13g2_fill_1 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_103 ();
 sg13g2_fill_2 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_117 ();
 sg13g2_decap_4 FILLER_16_135 ();
 sg13g2_fill_1 FILLER_16_139 ();
 sg13g2_fill_2 FILLER_16_156 ();
 sg13g2_fill_1 FILLER_16_158 ();
 sg13g2_fill_1 FILLER_16_163 ();
 sg13g2_fill_1 FILLER_16_188 ();
 sg13g2_fill_2 FILLER_16_267 ();
 sg13g2_fill_2 FILLER_16_298 ();
 sg13g2_fill_2 FILLER_16_327 ();
 sg13g2_fill_2 FILLER_16_332 ();
 sg13g2_fill_1 FILLER_16_334 ();
 sg13g2_fill_2 FILLER_16_339 ();
 sg13g2_fill_1 FILLER_16_341 ();
 sg13g2_fill_2 FILLER_16_352 ();
 sg13g2_fill_1 FILLER_16_354 ();
 sg13g2_decap_4 FILLER_16_426 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_4 FILLER_17_35 ();
 sg13g2_fill_1 FILLER_17_39 ();
 sg13g2_fill_2 FILLER_17_66 ();
 sg13g2_fill_2 FILLER_17_94 ();
 sg13g2_fill_2 FILLER_17_122 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_145 ();
 sg13g2_fill_2 FILLER_17_162 ();
 sg13g2_decap_4 FILLER_17_184 ();
 sg13g2_fill_2 FILLER_17_188 ();
 sg13g2_fill_2 FILLER_17_209 ();
 sg13g2_fill_1 FILLER_17_220 ();
 sg13g2_fill_2 FILLER_17_238 ();
 sg13g2_fill_2 FILLER_17_245 ();
 sg13g2_fill_2 FILLER_17_251 ();
 sg13g2_fill_1 FILLER_17_271 ();
 sg13g2_fill_1 FILLER_17_276 ();
 sg13g2_fill_2 FILLER_17_281 ();
 sg13g2_fill_1 FILLER_17_296 ();
 sg13g2_fill_2 FILLER_17_323 ();
 sg13g2_fill_1 FILLER_17_329 ();
 sg13g2_fill_2 FILLER_17_356 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_4 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_50 ();
 sg13g2_decap_8 FILLER_18_57 ();
 sg13g2_fill_2 FILLER_18_64 ();
 sg13g2_fill_2 FILLER_18_70 ();
 sg13g2_fill_1 FILLER_18_107 ();
 sg13g2_fill_1 FILLER_18_116 ();
 sg13g2_decap_4 FILLER_18_121 ();
 sg13g2_fill_1 FILLER_18_160 ();
 sg13g2_decap_8 FILLER_18_192 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_fill_1 FILLER_18_222 ();
 sg13g2_fill_2 FILLER_18_235 ();
 sg13g2_fill_2 FILLER_18_246 ();
 sg13g2_fill_2 FILLER_18_265 ();
 sg13g2_fill_1 FILLER_18_288 ();
 sg13g2_fill_2 FILLER_18_294 ();
 sg13g2_fill_1 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_318 ();
 sg13g2_fill_1 FILLER_18_326 ();
 sg13g2_fill_2 FILLER_18_347 ();
 sg13g2_fill_1 FILLER_18_349 ();
 sg13g2_fill_1 FILLER_18_354 ();
 sg13g2_fill_2 FILLER_18_360 ();
 sg13g2_fill_2 FILLER_18_366 ();
 sg13g2_fill_2 FILLER_18_394 ();
 sg13g2_fill_1 FILLER_18_396 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_4 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_32 ();
 sg13g2_decap_8 FILLER_19_38 ();
 sg13g2_decap_4 FILLER_19_45 ();
 sg13g2_fill_2 FILLER_19_49 ();
 sg13g2_decap_4 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_64 ();
 sg13g2_fill_2 FILLER_19_71 ();
 sg13g2_fill_2 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_163 ();
 sg13g2_fill_2 FILLER_19_168 ();
 sg13g2_fill_1 FILLER_19_170 ();
 sg13g2_fill_1 FILLER_19_174 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_decap_8 FILLER_19_185 ();
 sg13g2_decap_4 FILLER_19_192 ();
 sg13g2_fill_2 FILLER_19_229 ();
 sg13g2_fill_1 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_250 ();
 sg13g2_fill_1 FILLER_19_287 ();
 sg13g2_fill_1 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_341 ();
 sg13g2_fill_2 FILLER_19_368 ();
 sg13g2_fill_1 FILLER_19_383 ();
 sg13g2_fill_1 FILLER_19_389 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_11 ();
 sg13g2_decap_8 FILLER_20_16 ();
 sg13g2_decap_4 FILLER_20_79 ();
 sg13g2_fill_1 FILLER_20_83 ();
 sg13g2_fill_2 FILLER_20_135 ();
 sg13g2_fill_1 FILLER_20_137 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_224 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_fill_1 FILLER_20_242 ();
 sg13g2_fill_2 FILLER_20_251 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_fill_2 FILLER_20_264 ();
 sg13g2_fill_1 FILLER_20_271 ();
 sg13g2_decap_4 FILLER_20_286 ();
 sg13g2_fill_2 FILLER_20_293 ();
 sg13g2_fill_1 FILLER_20_295 ();
 sg13g2_fill_2 FILLER_20_304 ();
 sg13g2_decap_4 FILLER_20_316 ();
 sg13g2_fill_1 FILLER_20_324 ();
 sg13g2_fill_1 FILLER_20_332 ();
 sg13g2_fill_1 FILLER_20_337 ();
 sg13g2_fill_2 FILLER_20_348 ();
 sg13g2_decap_4 FILLER_20_367 ();
 sg13g2_fill_2 FILLER_20_371 ();
 sg13g2_fill_1 FILLER_20_390 ();
 sg13g2_fill_2 FILLER_20_413 ();
 sg13g2_fill_1 FILLER_20_415 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_fill_2 FILLER_20_427 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_fill_1 FILLER_21_39 ();
 sg13g2_fill_2 FILLER_21_68 ();
 sg13g2_fill_2 FILLER_21_83 ();
 sg13g2_fill_1 FILLER_21_85 ();
 sg13g2_decap_4 FILLER_21_90 ();
 sg13g2_fill_1 FILLER_21_94 ();
 sg13g2_decap_8 FILLER_21_99 ();
 sg13g2_fill_2 FILLER_21_106 ();
 sg13g2_fill_1 FILLER_21_199 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_fill_1 FILLER_21_208 ();
 sg13g2_fill_1 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_222 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_fill_2 FILLER_21_233 ();
 sg13g2_fill_2 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_280 ();
 sg13g2_fill_2 FILLER_21_323 ();
 sg13g2_fill_1 FILLER_21_325 ();
 sg13g2_fill_1 FILLER_21_330 ();
 sg13g2_fill_2 FILLER_21_341 ();
 sg13g2_fill_1 FILLER_22_26 ();
 sg13g2_fill_1 FILLER_22_39 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_fill_1 FILLER_22_55 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_fill_2 FILLER_22_112 ();
 sg13g2_fill_1 FILLER_22_114 ();
 sg13g2_decap_8 FILLER_22_122 ();
 sg13g2_decap_4 FILLER_22_129 ();
 sg13g2_fill_2 FILLER_22_137 ();
 sg13g2_fill_1 FILLER_22_139 ();
 sg13g2_fill_1 FILLER_22_144 ();
 sg13g2_fill_2 FILLER_22_180 ();
 sg13g2_fill_1 FILLER_22_214 ();
 sg13g2_fill_1 FILLER_22_225 ();
 sg13g2_fill_1 FILLER_22_230 ();
 sg13g2_fill_1 FILLER_22_236 ();
 sg13g2_fill_1 FILLER_22_242 ();
 sg13g2_fill_2 FILLER_22_284 ();
 sg13g2_fill_1 FILLER_22_303 ();
 sg13g2_fill_2 FILLER_22_342 ();
 sg13g2_fill_1 FILLER_22_348 ();
 sg13g2_fill_1 FILLER_22_375 ();
 sg13g2_decap_4 FILLER_22_420 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_11 ();
 sg13g2_decap_4 FILLER_23_18 ();
 sg13g2_fill_1 FILLER_23_25 ();
 sg13g2_fill_1 FILLER_23_35 ();
 sg13g2_fill_2 FILLER_23_41 ();
 sg13g2_fill_2 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_66 ();
 sg13g2_fill_2 FILLER_23_72 ();
 sg13g2_fill_2 FILLER_23_123 ();
 sg13g2_fill_1 FILLER_23_125 ();
 sg13g2_fill_2 FILLER_23_156 ();
 sg13g2_fill_2 FILLER_23_177 ();
 sg13g2_fill_1 FILLER_23_196 ();
 sg13g2_fill_2 FILLER_23_206 ();
 sg13g2_fill_2 FILLER_23_238 ();
 sg13g2_fill_2 FILLER_23_257 ();
 sg13g2_decap_4 FILLER_23_281 ();
 sg13g2_fill_2 FILLER_23_315 ();
 sg13g2_fill_1 FILLER_23_332 ();
 sg13g2_fill_1 FILLER_23_344 ();
 sg13g2_fill_2 FILLER_23_363 ();
 sg13g2_fill_1 FILLER_23_365 ();
 sg13g2_fill_1 FILLER_23_371 ();
 sg13g2_fill_2 FILLER_23_402 ();
 sg13g2_fill_1 FILLER_24_31 ();
 sg13g2_fill_2 FILLER_24_48 ();
 sg13g2_decap_4 FILLER_24_69 ();
 sg13g2_decap_8 FILLER_24_96 ();
 sg13g2_decap_4 FILLER_24_103 ();
 sg13g2_fill_1 FILLER_24_107 ();
 sg13g2_decap_4 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_143 ();
 sg13g2_fill_1 FILLER_24_150 ();
 sg13g2_fill_2 FILLER_24_158 ();
 sg13g2_fill_2 FILLER_24_173 ();
 sg13g2_fill_2 FILLER_24_180 ();
 sg13g2_fill_1 FILLER_24_182 ();
 sg13g2_fill_2 FILLER_24_193 ();
 sg13g2_fill_1 FILLER_24_195 ();
 sg13g2_fill_1 FILLER_24_200 ();
 sg13g2_fill_1 FILLER_24_214 ();
 sg13g2_fill_1 FILLER_24_233 ();
 sg13g2_fill_1 FILLER_24_247 ();
 sg13g2_fill_1 FILLER_24_253 ();
 sg13g2_fill_1 FILLER_24_259 ();
 sg13g2_fill_1 FILLER_24_289 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_fill_2 FILLER_24_393 ();
 sg13g2_fill_2 FILLER_24_398 ();
 sg13g2_fill_1 FILLER_25_31 ();
 sg13g2_fill_1 FILLER_25_36 ();
 sg13g2_fill_1 FILLER_25_47 ();
 sg13g2_decap_4 FILLER_25_52 ();
 sg13g2_fill_1 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_98 ();
 sg13g2_fill_1 FILLER_25_100 ();
 sg13g2_decap_4 FILLER_25_131 ();
 sg13g2_fill_1 FILLER_25_135 ();
 sg13g2_fill_2 FILLER_25_162 ();
 sg13g2_fill_1 FILLER_25_164 ();
 sg13g2_fill_2 FILLER_25_168 ();
 sg13g2_fill_1 FILLER_25_183 ();
 sg13g2_fill_1 FILLER_25_196 ();
 sg13g2_decap_4 FILLER_25_201 ();
 sg13g2_fill_1 FILLER_25_234 ();
 sg13g2_decap_4 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_258 ();
 sg13g2_fill_2 FILLER_25_290 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_fill_1 FILLER_25_345 ();
 sg13g2_fill_1 FILLER_25_351 ();
 sg13g2_fill_1 FILLER_25_362 ();
 sg13g2_fill_1 FILLER_25_371 ();
 sg13g2_fill_1 FILLER_25_378 ();
 sg13g2_fill_2 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_15 ();
 sg13g2_fill_2 FILLER_26_30 ();
 sg13g2_fill_1 FILLER_26_47 ();
 sg13g2_fill_1 FILLER_26_52 ();
 sg13g2_fill_2 FILLER_26_92 ();
 sg13g2_fill_1 FILLER_26_94 ();
 sg13g2_fill_2 FILLER_26_99 ();
 sg13g2_fill_2 FILLER_26_116 ();
 sg13g2_fill_2 FILLER_26_131 ();
 sg13g2_fill_1 FILLER_26_133 ();
 sg13g2_fill_1 FILLER_26_139 ();
 sg13g2_decap_4 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_153 ();
 sg13g2_decap_8 FILLER_26_160 ();
 sg13g2_fill_2 FILLER_26_167 ();
 sg13g2_fill_1 FILLER_26_192 ();
 sg13g2_fill_1 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_fill_1 FILLER_26_235 ();
 sg13g2_decap_4 FILLER_26_246 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_fill_1 FILLER_26_274 ();
 sg13g2_fill_2 FILLER_26_278 ();
 sg13g2_decap_4 FILLER_26_320 ();
 sg13g2_fill_1 FILLER_26_324 ();
 sg13g2_decap_4 FILLER_26_339 ();
 sg13g2_fill_1 FILLER_26_343 ();
 sg13g2_fill_1 FILLER_26_357 ();
 sg13g2_fill_1 FILLER_26_384 ();
 sg13g2_decap_4 FILLER_26_425 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_fill_2 FILLER_27_48 ();
 sg13g2_fill_2 FILLER_27_67 ();
 sg13g2_decap_4 FILLER_27_73 ();
 sg13g2_fill_2 FILLER_27_132 ();
 sg13g2_decap_4 FILLER_27_165 ();
 sg13g2_decap_4 FILLER_27_176 ();
 sg13g2_fill_1 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_207 ();
 sg13g2_fill_1 FILLER_27_211 ();
 sg13g2_fill_2 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_225 ();
 sg13g2_fill_2 FILLER_27_234 ();
 sg13g2_fill_2 FILLER_27_245 ();
 sg13g2_fill_1 FILLER_27_261 ();
 sg13g2_fill_1 FILLER_27_265 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_fill_1 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_302 ();
 sg13g2_fill_2 FILLER_27_307 ();
 sg13g2_fill_2 FILLER_27_313 ();
 sg13g2_fill_2 FILLER_27_318 ();
 sg13g2_fill_2 FILLER_27_325 ();
 sg13g2_fill_1 FILLER_27_327 ();
 sg13g2_fill_2 FILLER_27_376 ();
 sg13g2_fill_1 FILLER_27_382 ();
 sg13g2_fill_1 FILLER_27_388 ();
 sg13g2_fill_1 FILLER_27_392 ();
 sg13g2_fill_2 FILLER_27_410 ();
 sg13g2_fill_1 FILLER_28_30 ();
 sg13g2_fill_1 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_74 ();
 sg13g2_decap_8 FILLER_28_80 ();
 sg13g2_fill_1 FILLER_28_87 ();
 sg13g2_fill_1 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_148 ();
 sg13g2_decap_8 FILLER_28_157 ();
 sg13g2_decap_4 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_172 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_fill_1 FILLER_28_211 ();
 sg13g2_fill_2 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_242 ();
 sg13g2_fill_2 FILLER_28_295 ();
 sg13g2_decap_8 FILLER_28_323 ();
 sg13g2_decap_8 FILLER_28_330 ();
 sg13g2_fill_1 FILLER_28_341 ();
 sg13g2_fill_2 FILLER_28_347 ();
 sg13g2_fill_2 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_28_381 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_41 ();
 sg13g2_fill_1 FILLER_29_64 ();
 sg13g2_fill_1 FILLER_29_101 ();
 sg13g2_fill_2 FILLER_29_204 ();
 sg13g2_fill_1 FILLER_29_232 ();
 sg13g2_fill_1 FILLER_29_263 ();
 sg13g2_fill_1 FILLER_29_316 ();
 sg13g2_fill_2 FILLER_29_322 ();
 sg13g2_fill_2 FILLER_29_328 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_fill_2 FILLER_29_396 ();
 sg13g2_fill_1 FILLER_29_403 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_41 ();
 sg13g2_decap_4 FILLER_30_68 ();
 sg13g2_decap_8 FILLER_30_76 ();
 sg13g2_decap_4 FILLER_30_83 ();
 sg13g2_fill_2 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_146 ();
 sg13g2_decap_4 FILLER_30_151 ();
 sg13g2_decap_4 FILLER_30_160 ();
 sg13g2_fill_1 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_211 ();
 sg13g2_fill_1 FILLER_30_215 ();
 sg13g2_fill_1 FILLER_30_220 ();
 sg13g2_fill_2 FILLER_30_233 ();
 sg13g2_fill_2 FILLER_30_244 ();
 sg13g2_fill_1 FILLER_30_272 ();
 sg13g2_fill_1 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_305 ();
 sg13g2_fill_1 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_91 ();
 sg13g2_fill_2 FILLER_31_113 ();
 sg13g2_decap_4 FILLER_31_167 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_fill_1 FILLER_31_193 ();
 sg13g2_fill_1 FILLER_31_198 ();
 sg13g2_decap_4 FILLER_31_233 ();
 sg13g2_fill_2 FILLER_31_246 ();
 sg13g2_fill_1 FILLER_31_252 ();
 sg13g2_fill_1 FILLER_31_257 ();
 sg13g2_fill_2 FILLER_31_271 ();
 sg13g2_fill_1 FILLER_31_281 ();
 sg13g2_fill_1 FILLER_31_291 ();
 sg13g2_fill_1 FILLER_31_295 ();
 sg13g2_fill_2 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_31_381 ();
 sg13g2_fill_2 FILLER_31_391 ();
 sg13g2_fill_2 FILLER_31_428 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_68 ();
 sg13g2_fill_1 FILLER_32_75 ();
 sg13g2_fill_2 FILLER_32_107 ();
 sg13g2_fill_1 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_144 ();
 sg13g2_fill_1 FILLER_32_149 ();
 sg13g2_fill_1 FILLER_32_181 ();
 sg13g2_fill_2 FILLER_32_185 ();
 sg13g2_fill_2 FILLER_32_203 ();
 sg13g2_decap_4 FILLER_32_218 ();
 sg13g2_fill_1 FILLER_32_294 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_fill_2 FILLER_32_340 ();
 sg13g2_fill_1 FILLER_32_347 ();
 sg13g2_fill_2 FILLER_32_352 ();
 sg13g2_fill_1 FILLER_32_403 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_14 ();
 sg13g2_fill_2 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_32 ();
 sg13g2_fill_2 FILLER_33_53 ();
 sg13g2_fill_2 FILLER_33_59 ();
 sg13g2_fill_1 FILLER_33_66 ();
 sg13g2_fill_1 FILLER_33_70 ();
 sg13g2_decap_4 FILLER_33_79 ();
 sg13g2_fill_1 FILLER_33_83 ();
 sg13g2_decap_4 FILLER_33_88 ();
 sg13g2_fill_2 FILLER_33_97 ();
 sg13g2_fill_1 FILLER_33_99 ();
 sg13g2_fill_1 FILLER_33_169 ();
 sg13g2_fill_1 FILLER_33_176 ();
 sg13g2_decap_8 FILLER_33_212 ();
 sg13g2_fill_1 FILLER_33_219 ();
 sg13g2_fill_2 FILLER_33_232 ();
 sg13g2_fill_1 FILLER_33_244 ();
 sg13g2_fill_1 FILLER_33_268 ();
 sg13g2_fill_1 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_fill_1 FILLER_33_314 ();
 sg13g2_fill_2 FILLER_33_319 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_fill_1 FILLER_33_361 ();
 sg13g2_fill_1 FILLER_33_366 ();
 sg13g2_fill_2 FILLER_33_378 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_fill_1 FILLER_34_31 ();
 sg13g2_fill_2 FILLER_34_40 ();
 sg13g2_fill_1 FILLER_34_51 ();
 sg13g2_fill_2 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_142 ();
 sg13g2_fill_1 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_152 ();
 sg13g2_fill_2 FILLER_34_157 ();
 sg13g2_fill_1 FILLER_34_163 ();
 sg13g2_fill_1 FILLER_34_169 ();
 sg13g2_fill_2 FILLER_34_199 ();
 sg13g2_fill_1 FILLER_34_245 ();
 sg13g2_decap_4 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_258 ();
 sg13g2_fill_2 FILLER_34_267 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_6 ();
 sg13g2_fill_1 FILLER_35_20 ();
 sg13g2_fill_2 FILLER_35_60 ();
 sg13g2_fill_2 FILLER_35_66 ();
 sg13g2_fill_2 FILLER_35_120 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_178 ();
 sg13g2_fill_1 FILLER_35_190 ();
 sg13g2_fill_1 FILLER_35_200 ();
 sg13g2_fill_1 FILLER_35_210 ();
 sg13g2_fill_2 FILLER_35_227 ();
 sg13g2_fill_1 FILLER_35_233 ();
 sg13g2_fill_2 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_291 ();
 sg13g2_fill_1 FILLER_35_318 ();
 sg13g2_fill_1 FILLER_35_323 ();
 sg13g2_fill_1 FILLER_35_328 ();
 sg13g2_fill_1 FILLER_35_340 ();
 sg13g2_fill_1 FILLER_35_395 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_89 ();
 sg13g2_fill_1 FILLER_36_110 ();
 sg13g2_fill_1 FILLER_36_163 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_197 ();
 sg13g2_fill_2 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_232 ();
 sg13g2_fill_1 FILLER_36_234 ();
 sg13g2_fill_1 FILLER_36_239 ();
 sg13g2_fill_2 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_282 ();
 sg13g2_fill_2 FILLER_36_397 ();
 sg13g2_fill_2 FILLER_36_417 ();
 sg13g2_fill_1 FILLER_37_16 ();
 sg13g2_fill_2 FILLER_37_60 ();
 sg13g2_fill_1 FILLER_37_172 ();
 sg13g2_fill_1 FILLER_37_211 ();
 sg13g2_fill_2 FILLER_37_238 ();
 sg13g2_fill_1 FILLER_37_280 ();
 sg13g2_fill_2 FILLER_37_314 ();
 sg13g2_fill_2 FILLER_37_424 ();
 sg13g2_fill_2 FILLER_38_26 ();
 sg13g2_fill_2 FILLER_38_54 ();
 sg13g2_fill_1 FILLER_38_56 ();
 sg13g2_fill_1 FILLER_38_83 ();
 sg13g2_fill_2 FILLER_38_118 ();
 sg13g2_fill_2 FILLER_38_177 ();
 sg13g2_fill_1 FILLER_38_257 ();
 sg13g2_fill_2 FILLER_38_366 ();
endmodule
