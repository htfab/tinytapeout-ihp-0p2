module tt_um_rejunity_z80 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire clknet_leaf_0_clk;
 wire \addr_bus[0] ;
 wire \addr_bus[10] ;
 wire \addr_bus[11] ;
 wire \addr_bus[12] ;
 wire \addr_bus[13] ;
 wire \addr_bus[14] ;
 wire \addr_bus[15] ;
 wire \addr_bus[1] ;
 wire \addr_bus[2] ;
 wire \addr_bus[3] ;
 wire \addr_bus[4] ;
 wire \addr_bus[5] ;
 wire \addr_bus[6] ;
 wire \addr_bus[7] ;
 wire \addr_bus[8] ;
 wire \addr_bus[9] ;
 wire doe;
 wire \z80.iorq_n ;
 wire \z80.m1_n ;
 wire \z80.mreq_n ;
 wire \z80.rd_n ;
 wire \z80.rfsh_n ;
 wire \z80.tv80s.di_reg[0] ;
 wire \z80.tv80s.di_reg[1] ;
 wire \z80.tv80s.di_reg[2] ;
 wire \z80.tv80s.di_reg[3] ;
 wire \z80.tv80s.di_reg[4] ;
 wire \z80.tv80s.di_reg[5] ;
 wire \z80.tv80s.di_reg[6] ;
 wire \z80.tv80s.di_reg[7] ;
 wire \z80.tv80s.i_tv80_core.ACC[0] ;
 wire \z80.tv80s.i_tv80_core.ACC[1] ;
 wire \z80.tv80s.i_tv80_core.ACC[2] ;
 wire \z80.tv80s.i_tv80_core.ACC[3] ;
 wire \z80.tv80s.i_tv80_core.ACC[4] ;
 wire \z80.tv80s.i_tv80_core.ACC[5] ;
 wire \z80.tv80s.i_tv80_core.ACC[6] ;
 wire \z80.tv80s.i_tv80_core.ACC[7] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[0] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[1] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[2] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[3] ;
 wire \z80.tv80s.i_tv80_core.Alternate ;
 wire \z80.tv80s.i_tv80_core.Ap[0] ;
 wire \z80.tv80s.i_tv80_core.Ap[1] ;
 wire \z80.tv80s.i_tv80_core.Ap[2] ;
 wire \z80.tv80s.i_tv80_core.Ap[3] ;
 wire \z80.tv80s.i_tv80_core.Ap[4] ;
 wire \z80.tv80s.i_tv80_core.Ap[5] ;
 wire \z80.tv80s.i_tv80_core.Ap[6] ;
 wire \z80.tv80s.i_tv80_core.Ap[7] ;
 wire \z80.tv80s.i_tv80_core.Arith16_r ;
 wire \z80.tv80s.i_tv80_core.Auto_Wait_t1 ;
 wire \z80.tv80s.i_tv80_core.Auto_Wait_t2 ;
 wire \z80.tv80s.i_tv80_core.BTR_r ;
 wire \z80.tv80s.i_tv80_core.BusA[0] ;
 wire \z80.tv80s.i_tv80_core.BusA[1] ;
 wire \z80.tv80s.i_tv80_core.BusA[2] ;
 wire \z80.tv80s.i_tv80_core.BusA[3] ;
 wire \z80.tv80s.i_tv80_core.BusA[4] ;
 wire \z80.tv80s.i_tv80_core.BusA[5] ;
 wire \z80.tv80s.i_tv80_core.BusA[6] ;
 wire \z80.tv80s.i_tv80_core.BusA[7] ;
 wire \z80.tv80s.i_tv80_core.BusAck ;
 wire \z80.tv80s.i_tv80_core.BusB[0] ;
 wire \z80.tv80s.i_tv80_core.BusB[1] ;
 wire \z80.tv80s.i_tv80_core.BusB[2] ;
 wire \z80.tv80s.i_tv80_core.BusB[3] ;
 wire \z80.tv80s.i_tv80_core.BusB[4] ;
 wire \z80.tv80s.i_tv80_core.BusB[5] ;
 wire \z80.tv80s.i_tv80_core.BusB[6] ;
 wire \z80.tv80s.i_tv80_core.BusB[7] ;
 wire \z80.tv80s.i_tv80_core.BusReq_s ;
 wire \z80.tv80s.i_tv80_core.F[0] ;
 wire \z80.tv80s.i_tv80_core.F[1] ;
 wire \z80.tv80s.i_tv80_core.F[2] ;
 wire \z80.tv80s.i_tv80_core.F[3] ;
 wire \z80.tv80s.i_tv80_core.F[4] ;
 wire \z80.tv80s.i_tv80_core.F[5] ;
 wire \z80.tv80s.i_tv80_core.F[6] ;
 wire \z80.tv80s.i_tv80_core.F[7] ;
 wire \z80.tv80s.i_tv80_core.Fp[0] ;
 wire \z80.tv80s.i_tv80_core.Fp[1] ;
 wire \z80.tv80s.i_tv80_core.Fp[2] ;
 wire \z80.tv80s.i_tv80_core.Fp[3] ;
 wire \z80.tv80s.i_tv80_core.Fp[4] ;
 wire \z80.tv80s.i_tv80_core.Fp[5] ;
 wire \z80.tv80s.i_tv80_core.Fp[6] ;
 wire \z80.tv80s.i_tv80_core.Fp[7] ;
 wire \z80.tv80s.i_tv80_core.Halt_FF ;
 wire \z80.tv80s.i_tv80_core.INT_s ;
 wire \z80.tv80s.i_tv80_core.IR[0] ;
 wire \z80.tv80s.i_tv80_core.IR[1] ;
 wire \z80.tv80s.i_tv80_core.IR[2] ;
 wire \z80.tv80s.i_tv80_core.IR[3] ;
 wire \z80.tv80s.i_tv80_core.IR[4] ;
 wire \z80.tv80s.i_tv80_core.IR[5] ;
 wire \z80.tv80s.i_tv80_core.IR[6] ;
 wire \z80.tv80s.i_tv80_core.IR[7] ;
 wire \z80.tv80s.i_tv80_core.ISet[0] ;
 wire \z80.tv80s.i_tv80_core.ISet[1] ;
 wire \z80.tv80s.i_tv80_core.ISet[2] ;
 wire \z80.tv80s.i_tv80_core.ISet[3] ;
 wire \z80.tv80s.i_tv80_core.IStatus[1] ;
 wire \z80.tv80s.i_tv80_core.IStatus[2] ;
 wire \z80.tv80s.i_tv80_core.I[0] ;
 wire \z80.tv80s.i_tv80_core.I[1] ;
 wire \z80.tv80s.i_tv80_core.I[2] ;
 wire \z80.tv80s.i_tv80_core.I[3] ;
 wire \z80.tv80s.i_tv80_core.I[4] ;
 wire \z80.tv80s.i_tv80_core.I[5] ;
 wire \z80.tv80s.i_tv80_core.I[6] ;
 wire \z80.tv80s.i_tv80_core.I[7] ;
 wire \z80.tv80s.i_tv80_core.IncDecZ ;
 wire \z80.tv80s.i_tv80_core.IntCycle ;
 wire \z80.tv80s.i_tv80_core.IntE ;
 wire \z80.tv80s.i_tv80_core.IntE_FF2 ;
 wire \z80.tv80s.i_tv80_core.NMICycle ;
 wire \z80.tv80s.i_tv80_core.NMI_s ;
 wire \z80.tv80s.i_tv80_core.No_BTR ;
 wire \z80.tv80s.i_tv80_core.Oldnmi_n ;
 wire \z80.tv80s.i_tv80_core.PC[0] ;
 wire \z80.tv80s.i_tv80_core.PC[10] ;
 wire \z80.tv80s.i_tv80_core.PC[11] ;
 wire \z80.tv80s.i_tv80_core.PC[12] ;
 wire \z80.tv80s.i_tv80_core.PC[13] ;
 wire \z80.tv80s.i_tv80_core.PC[14] ;
 wire \z80.tv80s.i_tv80_core.PC[15] ;
 wire \z80.tv80s.i_tv80_core.PC[1] ;
 wire \z80.tv80s.i_tv80_core.PC[2] ;
 wire \z80.tv80s.i_tv80_core.PC[3] ;
 wire \z80.tv80s.i_tv80_core.PC[4] ;
 wire \z80.tv80s.i_tv80_core.PC[5] ;
 wire \z80.tv80s.i_tv80_core.PC[6] ;
 wire \z80.tv80s.i_tv80_core.PC[7] ;
 wire \z80.tv80s.i_tv80_core.PC[8] ;
 wire \z80.tv80s.i_tv80_core.PC[9] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ;
 wire \z80.tv80s.i_tv80_core.PreserveC_r ;
 wire \z80.tv80s.i_tv80_core.R[0] ;
 wire \z80.tv80s.i_tv80_core.R[1] ;
 wire \z80.tv80s.i_tv80_core.R[2] ;
 wire \z80.tv80s.i_tv80_core.R[3] ;
 wire \z80.tv80s.i_tv80_core.R[4] ;
 wire \z80.tv80s.i_tv80_core.R[5] ;
 wire \z80.tv80s.i_tv80_core.R[6] ;
 wire \z80.tv80s.i_tv80_core.R[7] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[2] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[10] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[11] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[12] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[13] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[14] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[15] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[3] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[4] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[5] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[6] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[7] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[8] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[9] ;
 wire \z80.tv80s.i_tv80_core.SP[0] ;
 wire \z80.tv80s.i_tv80_core.SP[10] ;
 wire \z80.tv80s.i_tv80_core.SP[11] ;
 wire \z80.tv80s.i_tv80_core.SP[12] ;
 wire \z80.tv80s.i_tv80_core.SP[13] ;
 wire \z80.tv80s.i_tv80_core.SP[14] ;
 wire \z80.tv80s.i_tv80_core.SP[15] ;
 wire \z80.tv80s.i_tv80_core.SP[1] ;
 wire \z80.tv80s.i_tv80_core.SP[2] ;
 wire \z80.tv80s.i_tv80_core.SP[3] ;
 wire \z80.tv80s.i_tv80_core.SP[4] ;
 wire \z80.tv80s.i_tv80_core.SP[5] ;
 wire \z80.tv80s.i_tv80_core.SP[6] ;
 wire \z80.tv80s.i_tv80_core.SP[7] ;
 wire \z80.tv80s.i_tv80_core.SP[8] ;
 wire \z80.tv80s.i_tv80_core.SP[9] ;
 wire \z80.tv80s.i_tv80_core.Save_ALU_r ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[0] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[10] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[11] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[12] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[13] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[14] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[15] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[1] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[2] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[3] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[4] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[5] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[6] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[7] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[8] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[9] ;
 wire \z80.tv80s.i_tv80_core.XY_Ind ;
 wire \z80.tv80s.i_tv80_core.XY_State[0] ;
 wire \z80.tv80s.i_tv80_core.XY_State[1] ;
 wire \z80.tv80s.i_tv80_core.Z16_r ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ;
 wire \z80.tv80s.i_tv80_core.mcycles[1] ;
 wire \z80.tv80s.i_tv80_core.mcycles[2] ;
 wire \z80.tv80s.i_tv80_core.mcycles[4] ;
 wire \z80.tv80s.i_tv80_core.mcycles[5] ;
 wire \z80.tv80s.i_tv80_core.ts[0] ;
 wire \z80.tv80s.i_tv80_core.ts[1] ;
 wire \z80.tv80s.i_tv80_core.ts[2] ;
 wire \z80.tv80s.i_tv80_core.ts[3] ;
 wire \z80.tv80s.i_tv80_core.ts[4] ;
 wire \z80.tv80s.i_tv80_core.ts[5] ;
 wire \z80.tv80s.i_tv80_core.ts[6] ;
 wire \z80.tv80s.wr_n ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_1 _05694_ (.A(ena),
    .X(_00635_));
 sg13g2_buf_1 _05695_ (.A(_00635_),
    .X(_00636_));
 sg13g2_buf_1 _05696_ (.A(\z80.tv80s.i_tv80_core.ts[2] ),
    .X(_00637_));
 sg13g2_buf_2 _05697_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ),
    .X(_00638_));
 sg13g2_buf_1 _05698_ (.A(_00638_),
    .X(_00639_));
 sg13g2_buf_1 _05699_ (.A(net369),
    .X(_00640_));
 sg13g2_buf_8 _05700_ (.A(\z80.tv80s.i_tv80_core.IR[2] ),
    .X(_00641_));
 sg13g2_buf_8 _05701_ (.A(_00641_),
    .X(_00642_));
 sg13g2_buf_1 _05702_ (.A(net368),
    .X(_00643_));
 sg13g2_buf_8 _05703_ (.A(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_00644_));
 sg13g2_buf_8 _05704_ (.A(_00644_),
    .X(_00645_));
 sg13g2_buf_8 _05705_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .X(_00646_));
 sg13g2_and2_1 _05706_ (.A(net367),
    .B(_00646_),
    .X(_00647_));
 sg13g2_buf_2 _05707_ (.A(_00647_),
    .X(_00648_));
 sg13g2_buf_8 _05708_ (.A(_00648_),
    .X(_00649_));
 sg13g2_buf_8 _05709_ (.A(\z80.tv80s.i_tv80_core.IR[1] ),
    .X(_00650_));
 sg13g2_buf_8 _05710_ (.A(_00650_),
    .X(_00651_));
 sg13g2_buf_8 _05711_ (.A(\z80.tv80s.i_tv80_core.IR[0] ),
    .X(_00652_));
 sg13g2_buf_8 _05712_ (.A(_00652_),
    .X(_00653_));
 sg13g2_nor2_1 _05713_ (.A(_00651_),
    .B(net365),
    .Y(_00654_));
 sg13g2_buf_2 _05714_ (.A(_00654_),
    .X(_00655_));
 sg13g2_nand3_1 _05715_ (.B(_00649_),
    .C(_00655_),
    .A(net323),
    .Y(_00656_));
 sg13g2_buf_2 _05716_ (.A(_00656_),
    .X(_00657_));
 sg13g2_nand2_1 _05717_ (.Y(_00658_),
    .A(_00644_),
    .B(_00646_));
 sg13g2_buf_8 _05718_ (.A(_00658_),
    .X(_00659_));
 sg13g2_buf_8 _05719_ (.A(_00659_),
    .X(_00660_));
 sg13g2_buf_8 _05720_ (.A(\z80.tv80s.i_tv80_core.IR[5] ),
    .X(_00661_));
 sg13g2_buf_8 _05721_ (.A(\z80.tv80s.i_tv80_core.IR[4] ),
    .X(_00662_));
 sg13g2_or2_1 _05722_ (.X(_00663_),
    .B(_00662_),
    .A(_00661_));
 sg13g2_buf_1 _05723_ (.A(_00663_),
    .X(_00664_));
 sg13g2_nor2_1 _05724_ (.A(net286),
    .B(_00664_),
    .Y(_00665_));
 sg13g2_nand2b_1 _05725_ (.Y(_00666_),
    .B(_00652_),
    .A_N(_00650_));
 sg13g2_buf_2 _05726_ (.A(_00666_),
    .X(_00667_));
 sg13g2_buf_8 _05727_ (.A(_00667_),
    .X(_00668_));
 sg13g2_buf_8 _05728_ (.A(net368),
    .X(_00669_));
 sg13g2_buf_8 _05729_ (.A(\z80.tv80s.i_tv80_core.IR[3] ),
    .X(_00670_));
 sg13g2_nand2_2 _05730_ (.Y(_00671_),
    .A(net321),
    .B(_00670_));
 sg13g2_nor2_2 _05731_ (.A(_00668_),
    .B(_00671_),
    .Y(_00672_));
 sg13g2_nand2_1 _05732_ (.Y(_00673_),
    .A(_00665_),
    .B(_00672_));
 sg13g2_buf_1 _05733_ (.A(_00673_),
    .X(_00674_));
 sg13g2_nand2_1 _05734_ (.Y(_00675_),
    .A(_00657_),
    .B(_00674_));
 sg13g2_inv_2 _05735_ (.Y(_00676_),
    .A(net368));
 sg13g2_or2_1 _05736_ (.X(_00677_),
    .B(net365),
    .A(_00650_));
 sg13g2_buf_8 _05737_ (.A(_00677_),
    .X(_00678_));
 sg13g2_nor3_1 _05738_ (.A(_00676_),
    .B(net286),
    .C(net284),
    .Y(_00679_));
 sg13g2_buf_8 _05739_ (.A(_00679_),
    .X(_00680_));
 sg13g2_buf_1 _05740_ (.A(_00662_),
    .X(_00681_));
 sg13g2_nor2b_1 _05741_ (.A(net364),
    .B_N(_00670_),
    .Y(_00682_));
 sg13g2_buf_2 _05742_ (.A(_00682_),
    .X(_00683_));
 sg13g2_buf_1 _05743_ (.A(\z80.tv80s.i_tv80_core.F[6] ),
    .X(_00684_));
 sg13g2_buf_2 _05744_ (.A(\z80.tv80s.i_tv80_core.F[2] ),
    .X(_00685_));
 sg13g2_buf_8 _05745_ (.A(_00661_),
    .X(_00686_));
 sg13g2_mux2_1 _05746_ (.A0(net397),
    .A1(_00685_),
    .S(net363),
    .X(_00687_));
 sg13g2_buf_1 _05747_ (.A(_00021_),
    .X(_00688_));
 sg13g2_inv_1 _05748_ (.Y(_00689_),
    .A(net396));
 sg13g2_and2_1 _05749_ (.A(net396),
    .B(net397),
    .X(_00690_));
 sg13g2_a21oi_1 _05750_ (.A1(_00689_),
    .A2(_00685_),
    .Y(_00691_),
    .B1(_00690_));
 sg13g2_buf_8 _05751_ (.A(_00670_),
    .X(_00692_));
 sg13g2_nor2_1 _05752_ (.A(net362),
    .B(net364),
    .Y(_00693_));
 sg13g2_nor2b_2 _05753_ (.A(_00692_),
    .B_N(_00662_),
    .Y(_00694_));
 sg13g2_and2_1 _05754_ (.A(_00670_),
    .B(_00662_),
    .X(_00695_));
 sg13g2_buf_1 _05755_ (.A(_00695_),
    .X(_00696_));
 sg13g2_buf_1 _05756_ (.A(\z80.tv80s.i_tv80_core.F[7] ),
    .X(_00697_));
 sg13g2_mux2_1 _05757_ (.A0(_00697_),
    .A1(\z80.tv80s.i_tv80_core.F[0] ),
    .S(net396),
    .X(_00698_));
 sg13g2_mux2_1 _05758_ (.A0(_00694_),
    .A1(_00696_),
    .S(_00698_),
    .X(_00699_));
 sg13g2_a221oi_1 _05759_ (.B2(_00693_),
    .C1(_00699_),
    .B1(_00691_),
    .A1(_00683_),
    .Y(_00700_),
    .A2(_00687_));
 sg13g2_buf_1 _05760_ (.A(_00700_),
    .X(_00701_));
 sg13g2_buf_2 _05761_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .X(_00702_));
 sg13g2_inv_2 _05762_ (.Y(_00703_),
    .A(_00702_));
 sg13g2_buf_1 _05763_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .X(_00704_));
 sg13g2_nand2_2 _05764_ (.Y(_00705_),
    .A(_00703_),
    .B(net395));
 sg13g2_a21o_1 _05765_ (.A2(net210),
    .A1(_00680_),
    .B1(_00705_),
    .X(_00706_));
 sg13g2_or2_1 _05766_ (.X(_00707_),
    .B(_00646_),
    .A(_00644_));
 sg13g2_buf_1 _05767_ (.A(_00707_),
    .X(_00708_));
 sg13g2_nand2b_1 _05768_ (.Y(_00709_),
    .B(_00670_),
    .A_N(_00641_));
 sg13g2_buf_8 _05769_ (.A(_00709_),
    .X(_00710_));
 sg13g2_nor3_1 _05770_ (.A(net320),
    .B(net285),
    .C(net319),
    .Y(_00711_));
 sg13g2_buf_1 _05771_ (.A(_00711_),
    .X(_00712_));
 sg13g2_buf_8 _05772_ (.A(net367),
    .X(_00713_));
 sg13g2_nor2b_1 _05773_ (.A(_00216_),
    .B_N(_00653_),
    .Y(_00714_));
 sg13g2_buf_8 _05774_ (.A(_00646_),
    .X(_00715_));
 sg13g2_nor2b_1 _05775_ (.A(net365),
    .B_N(net361),
    .Y(_00716_));
 sg13g2_nand2b_1 _05776_ (.Y(_00717_),
    .B(net321),
    .A_N(net366));
 sg13g2_nor4_1 _05777_ (.A(net318),
    .B(_00714_),
    .C(_00716_),
    .D(_00717_),
    .Y(_00718_));
 sg13g2_buf_1 _05778_ (.A(_00718_),
    .X(_00719_));
 sg13g2_nor2_2 _05779_ (.A(net209),
    .B(net208),
    .Y(_00720_));
 sg13g2_buf_1 _05780_ (.A(_00689_),
    .X(_00721_));
 sg13g2_nand2_1 _05781_ (.Y(_00722_),
    .A(net317),
    .B(_00694_));
 sg13g2_buf_1 _05782_ (.A(_00722_),
    .X(_00723_));
 sg13g2_a21oi_1 _05783_ (.A1(net208),
    .A2(net244),
    .Y(_00724_),
    .B1(_00703_));
 sg13g2_nor2_1 _05784_ (.A(_00720_),
    .B(_00724_),
    .Y(_00725_));
 sg13g2_a21oi_1 _05785_ (.A1(_00675_),
    .A2(_00706_),
    .Y(_00726_),
    .B1(_00725_));
 sg13g2_and2_1 _05786_ (.A(net366),
    .B(net365),
    .X(_00727_));
 sg13g2_buf_2 _05787_ (.A(_00727_),
    .X(_00728_));
 sg13g2_nor3_1 _05788_ (.A(_00642_),
    .B(_00645_),
    .C(net361),
    .Y(_00729_));
 sg13g2_buf_2 _05789_ (.A(_00729_),
    .X(_00730_));
 sg13g2_and2_1 _05790_ (.A(_00728_),
    .B(_00730_),
    .X(_00731_));
 sg13g2_buf_1 _05791_ (.A(_00731_),
    .X(_00732_));
 sg13g2_nand4_1 _05792_ (.B(_00662_),
    .C(net367),
    .A(net363),
    .Y(_00733_),
    .D(net361));
 sg13g2_buf_2 _05793_ (.A(_00733_),
    .X(_00734_));
 sg13g2_nor3_2 _05794_ (.A(net285),
    .B(net319),
    .C(_00734_),
    .Y(_00735_));
 sg13g2_nor2_1 _05795_ (.A(_00732_),
    .B(_00735_),
    .Y(_00736_));
 sg13g2_o21ai_1 _05796_ (.B1(_00736_),
    .Y(_00737_),
    .A1(net324),
    .A2(_00726_));
 sg13g2_buf_8 _05797_ (.A(net366),
    .X(_00738_));
 sg13g2_inv_1 _05798_ (.Y(_00739_),
    .A(net316));
 sg13g2_nor2_1 _05799_ (.A(net321),
    .B(net362),
    .Y(_00740_));
 sg13g2_nand2_1 _05800_ (.Y(_00741_),
    .A(net316),
    .B(net323));
 sg13g2_buf_1 _05801_ (.A(net363),
    .X(_00742_));
 sg13g2_buf_8 _05802_ (.A(net362),
    .X(_00743_));
 sg13g2_nand2b_1 _05803_ (.Y(_00744_),
    .B(net314),
    .A_N(net315));
 sg13g2_nor2_1 _05804_ (.A(_00741_),
    .B(_00744_),
    .Y(_00745_));
 sg13g2_a21o_1 _05805_ (.A2(_00740_),
    .A1(net283),
    .B1(_00745_),
    .X(_00746_));
 sg13g2_buf_1 _05806_ (.A(net365),
    .X(_00747_));
 sg13g2_inv_1 _05807_ (.Y(_00748_),
    .A(net313));
 sg13g2_buf_1 _05808_ (.A(_00748_),
    .X(_00749_));
 sg13g2_nor2_1 _05809_ (.A(net243),
    .B(net361),
    .Y(_00750_));
 sg13g2_buf_1 _05810_ (.A(net313),
    .X(_00751_));
 sg13g2_buf_1 _05811_ (.A(net316),
    .X(_00752_));
 sg13g2_nand2b_1 _05812_ (.Y(_00753_),
    .B(net363),
    .A_N(_00662_));
 sg13g2_buf_1 _05813_ (.A(_00753_),
    .X(_00754_));
 sg13g2_nor2_1 _05814_ (.A(_00686_),
    .B(net364),
    .Y(_00755_));
 sg13g2_buf_1 _05815_ (.A(_00755_),
    .X(_00756_));
 sg13g2_a22oi_1 _05816_ (.Y(_00757_),
    .B1(_00756_),
    .B2(net314),
    .A2(net280),
    .A1(net281));
 sg13g2_nor4_1 _05817_ (.A(_00751_),
    .B(net323),
    .C(net361),
    .D(_00757_),
    .Y(_00758_));
 sg13g2_a21o_1 _05818_ (.A2(_00750_),
    .A1(_00746_),
    .B1(_00758_),
    .X(_00759_));
 sg13g2_inv_1 _05819_ (.Y(_00760_),
    .A(net364));
 sg13g2_or2_1 _05820_ (.X(_00761_),
    .B(net363),
    .A(net362));
 sg13g2_nand3_1 _05821_ (.B(_00760_),
    .C(_00761_),
    .A(net313),
    .Y(_00762_));
 sg13g2_nor2b_1 _05822_ (.A(_00642_),
    .B_N(_00651_),
    .Y(_00763_));
 sg13g2_buf_1 _05823_ (.A(_00763_),
    .X(_00764_));
 sg13g2_and2_1 _05824_ (.A(_00764_),
    .B(_00648_),
    .X(_00765_));
 sg13g2_buf_1 _05825_ (.A(_00765_),
    .X(_00766_));
 sg13g2_nand2b_1 _05826_ (.Y(_00767_),
    .B(net366),
    .A_N(_00652_));
 sg13g2_buf_2 _05827_ (.A(_00767_),
    .X(_00768_));
 sg13g2_nor4_2 _05828_ (.A(net323),
    .B(_00754_),
    .C(net320),
    .Y(_00769_),
    .D(_00768_));
 sg13g2_a21oi_1 _05829_ (.A1(_00762_),
    .A2(_00766_),
    .Y(_00770_),
    .B1(_00769_));
 sg13g2_nor4_2 _05830_ (.A(_00659_),
    .B(net280),
    .C(_00667_),
    .Y(_00771_),
    .D(_00710_));
 sg13g2_or3_1 _05831_ (.A(net363),
    .B(net367),
    .C(_00646_),
    .X(_00772_));
 sg13g2_buf_8 _05832_ (.A(_00772_),
    .X(_00773_));
 sg13g2_nand3_1 _05833_ (.B(net365),
    .C(net368),
    .A(net366),
    .Y(_00774_));
 sg13g2_buf_2 _05834_ (.A(_00774_),
    .X(_00775_));
 sg13g2_nor3_1 _05835_ (.A(net362),
    .B(net279),
    .C(_00775_),
    .Y(_00776_));
 sg13g2_nand2_1 _05836_ (.Y(_00777_),
    .A(_00650_),
    .B(_00652_));
 sg13g2_nor4_1 _05837_ (.A(_00659_),
    .B(_00709_),
    .C(_00777_),
    .D(net322),
    .Y(_00778_));
 sg13g2_buf_1 _05838_ (.A(_00778_),
    .X(_00779_));
 sg13g2_inv_2 _05839_ (.Y(_00780_),
    .A(net363));
 sg13g2_nor3_1 _05840_ (.A(_00780_),
    .B(net320),
    .C(_00775_),
    .Y(_00781_));
 sg13g2_nor4_1 _05841_ (.A(_00771_),
    .B(_00776_),
    .C(net242),
    .D(_00781_),
    .Y(_00782_));
 sg13g2_nand3b_1 _05842_ (.B(_00216_),
    .C(net368),
    .Y(_00783_),
    .A_N(_00644_));
 sg13g2_buf_2 _05843_ (.A(_00783_),
    .X(_00784_));
 sg13g2_or2_1 _05844_ (.X(_00785_),
    .B(_00784_),
    .A(_00768_));
 sg13g2_buf_2 _05845_ (.A(_00785_),
    .X(_00786_));
 sg13g2_nand2b_1 _05846_ (.Y(_00787_),
    .B(net367),
    .A_N(net361));
 sg13g2_buf_1 _05847_ (.A(_00787_),
    .X(_00788_));
 sg13g2_nor2b_1 _05848_ (.A(net366),
    .B_N(net365),
    .Y(_00789_));
 sg13g2_buf_1 _05849_ (.A(_00789_),
    .X(_00790_));
 sg13g2_and2_1 _05850_ (.A(net368),
    .B(_00670_),
    .X(_00791_));
 sg13g2_buf_1 _05851_ (.A(_00791_),
    .X(_00792_));
 sg13g2_nand4_1 _05852_ (.B(_00790_),
    .C(net322),
    .A(net367),
    .Y(_00793_),
    .D(_00792_));
 sg13g2_and3_1 _05853_ (.X(_00794_),
    .A(_00786_),
    .B(net278),
    .C(_00793_));
 sg13g2_or2_1 _05854_ (.X(_00795_),
    .B(_00670_),
    .A(net368));
 sg13g2_buf_2 _05855_ (.A(_00795_),
    .X(_00796_));
 sg13g2_nor3_1 _05856_ (.A(_00659_),
    .B(net285),
    .C(_00796_),
    .Y(_00797_));
 sg13g2_nand3b_1 _05857_ (.B(_00641_),
    .C(_00650_),
    .Y(_00798_),
    .A_N(_00652_));
 sg13g2_buf_2 _05858_ (.A(_00798_),
    .X(_00799_));
 sg13g2_inv_1 _05859_ (.Y(_00800_),
    .A(_00646_));
 sg13g2_a21oi_1 _05860_ (.A1(net367),
    .A2(_00799_),
    .Y(_00801_),
    .B1(_00800_));
 sg13g2_buf_2 _05861_ (.A(_00801_),
    .X(_00802_));
 sg13g2_nor4_2 _05862_ (.A(_00659_),
    .B(_00753_),
    .C(net319),
    .Y(_00803_),
    .D(_00777_));
 sg13g2_nand2b_1 _05863_ (.Y(_00804_),
    .B(_00662_),
    .A_N(_00661_));
 sg13g2_buf_2 _05864_ (.A(_00804_),
    .X(_00805_));
 sg13g2_nor4_1 _05865_ (.A(_00659_),
    .B(_00667_),
    .C(net319),
    .D(_00805_),
    .Y(_00806_));
 sg13g2_buf_2 _05866_ (.A(_00806_),
    .X(_00807_));
 sg13g2_nor4_2 _05867_ (.A(_00797_),
    .B(_00802_),
    .C(_00803_),
    .Y(_00808_),
    .D(_00807_));
 sg13g2_nand4_1 _05868_ (.B(_00782_),
    .C(_00794_),
    .A(_00770_),
    .Y(_00809_),
    .D(_00808_));
 sg13g2_nor2_1 _05869_ (.A(net366),
    .B(net321),
    .Y(_00810_));
 sg13g2_buf_2 _05870_ (.A(_00810_),
    .X(_00811_));
 sg13g2_nand3_1 _05871_ (.B(_00756_),
    .C(_00811_),
    .A(net314),
    .Y(_00812_));
 sg13g2_nand2b_1 _05872_ (.Y(_00813_),
    .B(net362),
    .A_N(net316));
 sg13g2_and2_1 _05873_ (.A(net313),
    .B(_00669_),
    .X(_00814_));
 sg13g2_nor3_2 _05874_ (.A(_00738_),
    .B(_00747_),
    .C(_00669_),
    .Y(_00815_));
 sg13g2_a21oi_1 _05875_ (.A1(_00813_),
    .A2(_00814_),
    .Y(_00816_),
    .B1(_00815_));
 sg13g2_a21oi_2 _05876_ (.B1(net286),
    .Y(_00817_),
    .A2(_00816_),
    .A1(_00812_));
 sg13g2_nand3_1 _05877_ (.B(_00655_),
    .C(_00730_),
    .A(net322),
    .Y(_00818_));
 sg13g2_buf_2 _05878_ (.A(_00818_),
    .X(_00819_));
 sg13g2_buf_8 _05879_ (.A(_00702_),
    .X(_00820_));
 sg13g2_inv_1 _05880_ (.Y(_00821_),
    .A(net395));
 sg13g2_nor2_1 _05881_ (.A(net360),
    .B(_00821_),
    .Y(_00822_));
 sg13g2_buf_1 _05882_ (.A(_00822_),
    .X(_00823_));
 sg13g2_buf_1 _05883_ (.A(_00823_),
    .X(_00824_));
 sg13g2_buf_2 _05884_ (.A(\z80.tv80s.i_tv80_core.IntCycle ),
    .X(_00825_));
 sg13g2_buf_1 _05885_ (.A(\z80.tv80s.i_tv80_core.NMICycle ),
    .X(_00826_));
 sg13g2_nor2_1 _05886_ (.A(_00825_),
    .B(net394),
    .Y(_00827_));
 sg13g2_nor2_1 _05887_ (.A(net360),
    .B(net395),
    .Y(_00828_));
 sg13g2_buf_1 _05888_ (.A(_00828_),
    .X(_00829_));
 sg13g2_or4_1 _05889_ (.A(net368),
    .B(_00670_),
    .C(_00644_),
    .D(_00646_),
    .X(_00830_));
 sg13g2_buf_8 _05890_ (.A(_00830_),
    .X(_00831_));
 sg13g2_nor3_1 _05891_ (.A(net322),
    .B(net284),
    .C(_00831_),
    .Y(_00832_));
 sg13g2_buf_8 _05892_ (.A(_00832_),
    .X(_00833_));
 sg13g2_o21ai_1 _05893_ (.B1(_00833_),
    .Y(_00834_),
    .A1(_00827_),
    .A2(net277));
 sg13g2_o21ai_1 _05894_ (.B1(_00834_),
    .Y(_00835_),
    .A1(_00819_),
    .A2(net241));
 sg13g2_nor4_1 _05895_ (.A(_00759_),
    .B(_00809_),
    .C(_00817_),
    .D(_00835_),
    .Y(_00836_));
 sg13g2_a21oi_1 _05896_ (.A1(_00746_),
    .A2(_00750_),
    .Y(_00837_),
    .B1(_00758_));
 sg13g2_and4_1 _05897_ (.A(_00770_),
    .B(_00782_),
    .C(_00794_),
    .D(_00808_),
    .X(_00838_));
 sg13g2_buf_1 _05898_ (.A(_00838_),
    .X(_00839_));
 sg13g2_or2_1 _05899_ (.X(_00840_),
    .B(_00735_),
    .A(_00732_));
 sg13g2_nor2_1 _05900_ (.A(net367),
    .B(_00715_),
    .Y(_00841_));
 sg13g2_buf_2 _05901_ (.A(_00841_),
    .X(_00842_));
 sg13g2_nor2b_1 _05902_ (.A(net321),
    .B_N(net362),
    .Y(_00843_));
 sg13g2_nand3_1 _05903_ (.B(_00790_),
    .C(_00843_),
    .A(_00842_),
    .Y(_00844_));
 sg13g2_buf_2 _05904_ (.A(_00844_),
    .X(_00845_));
 sg13g2_nand2_1 _05905_ (.Y(_00846_),
    .A(_00845_),
    .B(_00819_));
 sg13g2_nor4_2 _05906_ (.A(net286),
    .B(net285),
    .C(net322),
    .Y(_00847_),
    .D(_00671_));
 sg13g2_or4_1 _05907_ (.A(_00680_),
    .B(_00847_),
    .C(_00833_),
    .D(_00718_),
    .X(_00848_));
 sg13g2_nor4_2 _05908_ (.A(_00840_),
    .B(_00846_),
    .C(_00817_),
    .Y(_00849_),
    .D(_00848_));
 sg13g2_buf_2 _05909_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .X(_00850_));
 sg13g2_inv_2 _05910_ (.Y(_00851_),
    .A(_00850_));
 sg13g2_buf_2 _05911_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .X(_00852_));
 sg13g2_nand2_1 _05912_ (.Y(_00853_),
    .A(_00851_),
    .B(_00852_));
 sg13g2_buf_1 _05913_ (.A(net360),
    .X(_00854_));
 sg13g2_a21oi_1 _05914_ (.A1(_00821_),
    .A2(_00853_),
    .Y(_00855_),
    .B1(net312));
 sg13g2_nor2_1 _05915_ (.A(net369),
    .B(_00855_),
    .Y(_00856_));
 sg13g2_nand4_1 _05916_ (.B(_00839_),
    .C(_00849_),
    .A(_00837_),
    .Y(_00857_),
    .D(_00856_));
 sg13g2_o21ai_1 _05917_ (.B1(_00857_),
    .Y(_00858_),
    .A1(net324),
    .A2(_00836_));
 sg13g2_buf_2 _05918_ (.A(\z80.tv80s.i_tv80_core.ISet[0] ),
    .X(_00859_));
 sg13g2_buf_1 _05919_ (.A(_00859_),
    .X(_00860_));
 sg13g2_o21ai_1 _05920_ (.B1(net359),
    .Y(_00861_),
    .A1(_00737_),
    .A2(_00858_));
 sg13g2_buf_1 _05921_ (.A(\z80.tv80s.i_tv80_core.ISet[2] ),
    .X(_00862_));
 sg13g2_buf_1 _05922_ (.A(_00862_),
    .X(_00863_));
 sg13g2_o21ai_1 _05923_ (.B1(_00786_),
    .Y(_00864_),
    .A1(_00842_),
    .A2(_00799_));
 sg13g2_buf_1 _05924_ (.A(_00864_),
    .X(_00865_));
 sg13g2_buf_2 _05925_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ),
    .X(_00866_));
 sg13g2_nor2_1 _05926_ (.A(_00703_),
    .B(_00866_),
    .Y(_00867_));
 sg13g2_a21oi_1 _05927_ (.A1(_00865_),
    .A2(_00867_),
    .Y(_00868_),
    .B1(net324));
 sg13g2_nor2_1 _05928_ (.A(_00862_),
    .B(_00859_),
    .Y(_00869_));
 sg13g2_buf_1 _05929_ (.A(_00869_),
    .X(_00870_));
 sg13g2_buf_1 _05930_ (.A(_00870_),
    .X(_00871_));
 sg13g2_a21oi_1 _05931_ (.A1(net358),
    .A2(_00868_),
    .Y(_00872_),
    .B1(net276));
 sg13g2_or2_1 _05932_ (.X(_00873_),
    .B(_00859_),
    .A(_00862_));
 sg13g2_buf_1 _05933_ (.A(_00873_),
    .X(_00874_));
 sg13g2_buf_1 _05934_ (.A(_00676_),
    .X(_00875_));
 sg13g2_nor2b_1 _05935_ (.A(net313),
    .B_N(net316),
    .Y(_00876_));
 sg13g2_buf_2 _05936_ (.A(_00876_),
    .X(_00877_));
 sg13g2_nand2_2 _05937_ (.Y(_00878_),
    .A(net275),
    .B(_00877_));
 sg13g2_nor2_1 _05938_ (.A(_00878_),
    .B(net278),
    .Y(_00879_));
 sg13g2_buf_1 _05939_ (.A(_00879_),
    .X(_00880_));
 sg13g2_inv_1 _05940_ (.Y(_00881_),
    .A(_00638_));
 sg13g2_buf_1 _05941_ (.A(_00881_),
    .X(_00882_));
 sg13g2_buf_1 _05942_ (.A(_00775_),
    .X(_00883_));
 sg13g2_nor3_1 _05943_ (.A(net280),
    .B(net240),
    .C(net278),
    .Y(_00884_));
 sg13g2_buf_2 _05944_ (.A(_00884_),
    .X(_00885_));
 sg13g2_nand2_2 _05945_ (.Y(_00886_),
    .A(_00823_),
    .B(_00885_));
 sg13g2_and3_1 _05946_ (.X(_00887_),
    .A(net316),
    .B(net313),
    .C(net321));
 sg13g2_buf_2 _05947_ (.A(_00887_),
    .X(_00888_));
 sg13g2_nand2_1 _05948_ (.Y(_00889_),
    .A(_00780_),
    .B(_00888_));
 sg13g2_or2_1 _05949_ (.X(_00890_),
    .B(_00889_),
    .A(net278));
 sg13g2_buf_1 _05950_ (.A(net395),
    .X(_00891_));
 sg13g2_nand2_1 _05951_ (.Y(_00892_),
    .A(net357),
    .B(_00728_));
 sg13g2_nand2b_1 _05952_ (.Y(_00893_),
    .B(_00715_),
    .A_N(_00645_));
 sg13g2_buf_2 _05953_ (.A(_00893_),
    .X(_00894_));
 sg13g2_nor3_1 _05954_ (.A(_00643_),
    .B(_00780_),
    .C(_00894_),
    .Y(_00895_));
 sg13g2_buf_1 _05955_ (.A(_00895_),
    .X(_00896_));
 sg13g2_a21oi_1 _05956_ (.A1(_00821_),
    .A2(_00851_),
    .Y(_00897_),
    .B1(net312));
 sg13g2_nand3_1 _05957_ (.B(net207),
    .C(_00897_),
    .A(_00892_),
    .Y(_00898_));
 sg13g2_nand4_1 _05958_ (.B(_00886_),
    .C(_00890_),
    .A(net311),
    .Y(_00899_),
    .D(_00898_));
 sg13g2_a21oi_1 _05959_ (.A1(net312),
    .A2(net170),
    .Y(_00900_),
    .B1(_00899_));
 sg13g2_inv_1 _05960_ (.Y(_00901_),
    .A(_00866_));
 sg13g2_o21ai_1 _05961_ (.B1(_00901_),
    .Y(_00902_),
    .A1(_00874_),
    .A2(_00900_));
 sg13g2_a21oi_2 _05962_ (.B1(_00902_),
    .Y(_00903_),
    .A2(_00872_),
    .A1(_00861_));
 sg13g2_mux2_1 _05963_ (.A0(\z80.tv80s.i_tv80_core.ts[0] ),
    .A1(net398),
    .S(_00903_),
    .X(_00904_));
 sg13g2_buf_1 _05964_ (.A(\z80.tv80s.i_tv80_core.ts[4] ),
    .X(_00905_));
 sg13g2_inv_1 _05965_ (.Y(_00906_),
    .A(_00030_));
 sg13g2_mux2_1 _05966_ (.A0(net393),
    .A1(_00906_),
    .S(_00903_),
    .X(_00907_));
 sg13g2_buf_1 _05967_ (.A(\z80.tv80s.i_tv80_core.ts[3] ),
    .X(_00908_));
 sg13g2_buf_1 _05968_ (.A(_00908_),
    .X(_00909_));
 sg13g2_mux2_1 _05969_ (.A0(\z80.tv80s.i_tv80_core.ts[1] ),
    .A1(_00909_),
    .S(_00903_),
    .X(_00910_));
 sg13g2_mux2_1 _05970_ (.A0(\z80.tv80s.i_tv80_core.ts[5] ),
    .A1(\z80.tv80s.i_tv80_core.ts[0] ),
    .S(_00903_),
    .X(_00911_));
 sg13g2_nand3_1 _05971_ (.B(_00839_),
    .C(_00849_),
    .A(_00837_),
    .Y(_00912_));
 sg13g2_buf_2 _05972_ (.A(_00912_),
    .X(_00913_));
 sg13g2_buf_1 _05973_ (.A(_00756_),
    .X(_00914_));
 sg13g2_buf_1 _05974_ (.A(_00643_),
    .X(_00915_));
 sg13g2_buf_1 _05975_ (.A(net314),
    .X(_00916_));
 sg13g2_buf_1 _05976_ (.A(net361),
    .X(_00917_));
 sg13g2_nor4_2 _05977_ (.A(net274),
    .B(net273),
    .C(net318),
    .Y(_00918_),
    .D(_00917_));
 sg13g2_nand3_1 _05978_ (.B(_00655_),
    .C(_00918_),
    .A(net239),
    .Y(_00919_));
 sg13g2_buf_1 _05979_ (.A(_00919_),
    .X(_00920_));
 sg13g2_or2_1 _05980_ (.X(_00921_),
    .B(_00826_),
    .A(_00825_));
 sg13g2_buf_1 _05981_ (.A(_00921_),
    .X(_00922_));
 sg13g2_buf_2 _05982_ (.A(_00217_),
    .X(_00923_));
 sg13g2_buf_1 _05983_ (.A(_00821_),
    .X(_00924_));
 sg13g2_nand2_1 _05984_ (.Y(_00925_),
    .A(_00923_),
    .B(net309));
 sg13g2_a21oi_1 _05985_ (.A1(_00922_),
    .A2(_00925_),
    .Y(_00926_),
    .B1(net324));
 sg13g2_o21ai_1 _05986_ (.B1(_00736_),
    .Y(_00927_),
    .A1(net185),
    .A2(_00926_));
 sg13g2_nor3_2 _05987_ (.A(_00657_),
    .B(net210),
    .C(_00705_),
    .Y(_00928_));
 sg13g2_a22oi_1 _05988_ (.Y(_00929_),
    .B1(_00705_),
    .B2(net311),
    .A2(_00674_),
    .A1(_00819_));
 sg13g2_inv_2 _05989_ (.Y(_00930_),
    .A(_00692_));
 sg13g2_buf_1 _05990_ (.A(net364),
    .X(_00931_));
 sg13g2_nand2_1 _05991_ (.Y(_00932_),
    .A(net308),
    .B(net307));
 sg13g2_buf_1 _05992_ (.A(_00932_),
    .X(_00933_));
 sg13g2_nor2_1 _05993_ (.A(net396),
    .B(_00933_),
    .Y(_00934_));
 sg13g2_buf_1 _05994_ (.A(_00934_),
    .X(_00935_));
 sg13g2_o21ai_1 _05995_ (.B1(net312),
    .Y(_00936_),
    .A1(net209),
    .A2(net184));
 sg13g2_a21oi_1 _05996_ (.A1(_00882_),
    .A2(_00936_),
    .Y(_00937_),
    .B1(_00720_));
 sg13g2_nor4_1 _05997_ (.A(_00927_),
    .B(_00928_),
    .C(_00929_),
    .D(_00937_),
    .Y(_00938_));
 sg13g2_nor2_1 _05998_ (.A(_00759_),
    .B(_00809_),
    .Y(_00939_));
 sg13g2_buf_2 _05999_ (.A(_00939_),
    .X(_00940_));
 sg13g2_nand2b_1 _06000_ (.Y(_00941_),
    .B(_00940_),
    .A_N(_00817_));
 sg13g2_buf_1 _06001_ (.A(net324),
    .X(_00942_));
 sg13g2_o21ai_1 _06002_ (.B1(net272),
    .Y(_00943_),
    .A1(_00680_),
    .A2(_00941_));
 sg13g2_and3_1 _06003_ (.X(_00944_),
    .A(_00913_),
    .B(_00938_),
    .C(_00943_));
 sg13g2_nand2_1 _06004_ (.Y(_00945_),
    .A(net359),
    .B(_00857_));
 sg13g2_inv_1 _06005_ (.Y(_00946_),
    .A(_00868_));
 sg13g2_a21oi_1 _06006_ (.A1(net358),
    .A2(_00946_),
    .Y(_00947_),
    .B1(_00902_));
 sg13g2_o21ai_1 _06007_ (.B1(_00947_),
    .Y(_00948_),
    .A1(_00944_),
    .A2(_00945_));
 sg13g2_nor2_1 _06008_ (.A(net272),
    .B(_00726_),
    .Y(_00949_));
 sg13g2_buf_1 _06009_ (.A(_00703_),
    .X(_00950_));
 sg13g2_buf_1 _06010_ (.A(net315),
    .X(_00951_));
 sg13g2_and2_1 _06011_ (.A(_00655_),
    .B(_00730_),
    .X(_00952_));
 sg13g2_buf_1 _06012_ (.A(_00952_),
    .X(_00953_));
 sg13g2_o21ai_1 _06013_ (.B1(_00953_),
    .Y(_00954_),
    .A1(net271),
    .A2(_00696_));
 sg13g2_buf_1 _06014_ (.A(_00954_),
    .X(_00955_));
 sg13g2_nand3_1 _06015_ (.B(net309),
    .C(_00833_),
    .A(net311),
    .Y(_00956_));
 sg13g2_o21ai_1 _06016_ (.B1(_00956_),
    .Y(_00957_),
    .A1(net309),
    .A2(_00955_));
 sg13g2_and2_1 _06017_ (.A(net306),
    .B(_00957_),
    .X(_00958_));
 sg13g2_nor3_2 _06018_ (.A(_00805_),
    .B(net284),
    .C(_00831_),
    .Y(_00959_));
 sg13g2_nor4_1 _06019_ (.A(_00817_),
    .B(_00949_),
    .C(_00958_),
    .D(_00959_),
    .Y(_00960_));
 sg13g2_buf_1 _06020_ (.A(net272),
    .X(_00961_));
 sg13g2_nor2_1 _06021_ (.A(net185),
    .B(_00827_),
    .Y(_00962_));
 sg13g2_o21ai_1 _06022_ (.B1(_00955_),
    .Y(_00963_),
    .A1(net185),
    .A2(_00922_));
 sg13g2_a21oi_1 _06023_ (.A1(_00849_),
    .A2(_00705_),
    .Y(_00964_),
    .B1(_00963_));
 sg13g2_a21oi_1 _06024_ (.A1(_00940_),
    .A2(_00964_),
    .Y(_00965_),
    .B1(net272));
 sg13g2_a21oi_1 _06025_ (.A1(net238),
    .A2(_00962_),
    .Y(_00966_),
    .B1(_00965_));
 sg13g2_inv_2 _06026_ (.Y(_00967_),
    .A(_00859_));
 sg13g2_buf_1 _06027_ (.A(net355),
    .X(_00968_));
 sg13g2_a21oi_1 _06028_ (.A1(_00960_),
    .A2(_00966_),
    .Y(_00969_),
    .B1(net305));
 sg13g2_buf_1 _06029_ (.A(net312),
    .X(_00970_));
 sg13g2_buf_2 _06030_ (.A(_00022_),
    .X(_00971_));
 sg13g2_a21oi_1 _06031_ (.A1(net243),
    .A2(_00971_),
    .Y(_00972_),
    .B1(net283));
 sg13g2_buf_1 _06032_ (.A(net207),
    .X(_00973_));
 sg13g2_a22oi_1 _06033_ (.Y(_00974_),
    .B1(_00972_),
    .B2(net183),
    .A2(net170),
    .A1(net270));
 sg13g2_nand2_1 _06034_ (.Y(_00975_),
    .A(net312),
    .B(net183));
 sg13g2_nor2b_1 _06035_ (.A(_00681_),
    .B_N(net363),
    .Y(_00976_));
 sg13g2_buf_1 _06036_ (.A(_00976_),
    .X(_00977_));
 sg13g2_inv_1 _06037_ (.Y(_00978_),
    .A(_00713_));
 sg13g2_nor2_1 _06038_ (.A(_00978_),
    .B(net310),
    .Y(_00979_));
 sg13g2_nand3_1 _06039_ (.B(_00888_),
    .C(_00979_),
    .A(net269),
    .Y(_00980_));
 sg13g2_buf_2 _06040_ (.A(_00980_),
    .X(_00981_));
 sg13g2_nand2_1 _06041_ (.Y(_00982_),
    .A(net282),
    .B(_00981_));
 sg13g2_o21ai_1 _06042_ (.B1(_00982_),
    .Y(_00983_),
    .A1(net282),
    .A2(_00975_));
 sg13g2_buf_1 _06043_ (.A(net281),
    .X(_00984_));
 sg13g2_a22oi_1 _06044_ (.Y(_00985_),
    .B1(_00983_),
    .B2(net237),
    .A2(_00974_),
    .A1(_00886_));
 sg13g2_buf_1 _06045_ (.A(_00788_),
    .X(_00986_));
 sg13g2_nor2_1 _06046_ (.A(net236),
    .B(_00889_),
    .Y(_00987_));
 sg13g2_a21oi_1 _06047_ (.A1(_00728_),
    .A2(net183),
    .Y(_00988_),
    .B1(_00987_));
 sg13g2_o21ai_1 _06048_ (.B1(_00988_),
    .Y(_00989_),
    .A1(net238),
    .A2(_00985_));
 sg13g2_buf_1 _06049_ (.A(_00212_),
    .X(_00990_));
 sg13g2_inv_1 _06050_ (.Y(_00991_),
    .A(_00990_));
 sg13g2_a221oi_1 _06051_ (.B2(net276),
    .C1(_00991_),
    .B1(_00989_),
    .A1(net358),
    .Y(_00992_),
    .A2(_00868_));
 sg13g2_nand2b_1 _06052_ (.Y(_00993_),
    .B(_00992_),
    .A_N(_00969_));
 sg13g2_mux4_1 _06053_ (.S0(_00948_),
    .A0(_00904_),
    .A1(_00907_),
    .A2(_00910_),
    .A3(_00911_),
    .S1(_00993_),
    .X(_00994_));
 sg13g2_buf_2 _06054_ (.A(_00994_),
    .X(_00995_));
 sg13g2_nand2b_1 _06055_ (.Y(_00996_),
    .B(net398),
    .A_N(net2));
 sg13g2_buf_1 _06056_ (.A(_00996_),
    .X(_00997_));
 sg13g2_buf_1 _06057_ (.A(\z80.tv80s.i_tv80_core.BusAck ),
    .X(_00998_));
 sg13g2_nand2_1 _06058_ (.Y(_00999_),
    .A(_00998_),
    .B(\z80.tv80s.i_tv80_core.BusReq_s ));
 sg13g2_and4_1 _06059_ (.A(net399),
    .B(_00995_),
    .C(_00997_),
    .D(_00999_),
    .X(_01000_));
 sg13g2_and2_1 _06060_ (.A(_00031_),
    .B(_01000_),
    .X(_01001_));
 sg13g2_buf_1 _06061_ (.A(_01001_),
    .X(_01002_));
 sg13g2_buf_1 _06062_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .X(_01003_));
 sg13g2_nor2b_1 _06063_ (.A(_01003_),
    .B_N(_00990_),
    .Y(_01004_));
 sg13g2_nor2_2 _06064_ (.A(_00850_),
    .B(_00852_),
    .Y(_01005_));
 sg13g2_nand3_1 _06065_ (.B(_01004_),
    .C(_01005_),
    .A(net357),
    .Y(_01006_));
 sg13g2_buf_1 _06066_ (.A(_01006_),
    .X(_01007_));
 sg13g2_buf_1 _06067_ (.A(_01003_),
    .X(_01008_));
 sg13g2_nand2b_1 _06068_ (.Y(_01009_),
    .B(_00852_),
    .A_N(net354));
 sg13g2_nand3_1 _06069_ (.B(_01007_),
    .C(_01009_),
    .A(_00990_),
    .Y(_01010_));
 sg13g2_nand2b_1 _06070_ (.Y(_01011_),
    .B(_00636_),
    .A_N(\z80.tv80s.i_tv80_core.BusReq_s ));
 sg13g2_nand3b_1 _06071_ (.B(_00997_),
    .C(_00995_),
    .Y(_01012_),
    .A_N(_01011_));
 sg13g2_buf_1 _06072_ (.A(_01012_),
    .X(_01013_));
 sg13g2_buf_1 _06073_ (.A(_00866_),
    .X(_01014_));
 sg13g2_nor2_1 _06074_ (.A(net354),
    .B(net353),
    .Y(_01015_));
 sg13g2_buf_1 _06075_ (.A(net270),
    .X(_01016_));
 sg13g2_buf_1 _06076_ (.A(net235),
    .X(_01017_));
 sg13g2_nand4_1 _06077_ (.B(net309),
    .C(_01015_),
    .A(_01017_),
    .Y(_01018_),
    .D(_01005_));
 sg13g2_nor2_1 _06078_ (.A(_00851_),
    .B(_00852_),
    .Y(_01019_));
 sg13g2_a21oi_1 _06079_ (.A1(_00852_),
    .A2(_00990_),
    .Y(_01020_),
    .B1(_01019_));
 sg13g2_nand4_1 _06080_ (.B(_01007_),
    .C(_01018_),
    .A(_01015_),
    .Y(_01021_),
    .D(_01020_));
 sg13g2_nor2_1 _06081_ (.A(_01013_),
    .B(_01021_),
    .Y(_01022_));
 sg13g2_a21o_1 _06082_ (.A2(_01010_),
    .A1(_01002_),
    .B1(_01022_),
    .X(_01023_));
 sg13g2_buf_1 _06083_ (.A(net320),
    .X(_01024_));
 sg13g2_nand2_1 _06084_ (.Y(_01025_),
    .A(_00686_),
    .B(_00662_));
 sg13g2_buf_2 _06085_ (.A(_01025_),
    .X(_01026_));
 sg13g2_nor4_1 _06086_ (.A(net273),
    .B(net268),
    .C(_00799_),
    .D(_01026_),
    .Y(_01027_));
 sg13g2_buf_2 _06087_ (.A(_01027_),
    .X(_01028_));
 sg13g2_buf_1 _06088_ (.A(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_01029_));
 sg13g2_buf_1 _06089_ (.A(_01029_),
    .X(_01030_));
 sg13g2_buf_1 _06090_ (.A(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .X(_01031_));
 sg13g2_or2_1 _06091_ (.X(_01032_),
    .B(\z80.tv80s.i_tv80_core.XY_State[0] ),
    .A(_01031_));
 sg13g2_buf_1 _06092_ (.A(_01032_),
    .X(_01033_));
 sg13g2_nand2b_2 _06093_ (.Y(_01034_),
    .B(net304),
    .A_N(_01030_));
 sg13g2_o21ai_1 _06094_ (.B1(_01003_),
    .Y(_01035_),
    .A1(net242),
    .A2(_01028_));
 sg13g2_nor4_1 _06095_ (.A(_00680_),
    .B(_00847_),
    .C(_00833_),
    .D(net208),
    .Y(_01036_));
 sg13g2_a21oi_1 _06096_ (.A1(net282),
    .A2(net322),
    .Y(_01037_),
    .B1(net274));
 sg13g2_buf_1 _06097_ (.A(_00660_),
    .X(_01038_));
 sg13g2_nor2b_1 _06098_ (.A(_00751_),
    .B_N(net274),
    .Y(_01039_));
 sg13g2_nor3_1 _06099_ (.A(_00764_),
    .B(net234),
    .C(_01039_),
    .Y(_01040_));
 sg13g2_o21ai_1 _06100_ (.B1(_01040_),
    .Y(_01041_),
    .A1(_00813_),
    .A2(_01037_));
 sg13g2_buf_1 _06101_ (.A(_00768_),
    .X(_01042_));
 sg13g2_nor2_1 _06102_ (.A(net274),
    .B(net233),
    .Y(_01043_));
 sg13g2_buf_2 _06103_ (.A(_01043_),
    .X(_01044_));
 sg13g2_buf_1 _06104_ (.A(_00777_),
    .X(_01045_));
 sg13g2_nor4_1 _06105_ (.A(net286),
    .B(_00754_),
    .C(net303),
    .D(_00796_),
    .Y(_01046_));
 sg13g2_buf_1 _06106_ (.A(_01046_),
    .X(_01047_));
 sg13g2_a21oi_1 _06107_ (.A1(_00842_),
    .A2(_01044_),
    .Y(_01048_),
    .B1(net205));
 sg13g2_inv_1 _06108_ (.Y(_01049_),
    .A(_00216_));
 sg13g2_o21ai_1 _06109_ (.B1(_00800_),
    .Y(_01050_),
    .A1(_01049_),
    .A2(_00799_));
 sg13g2_nand2_1 _06110_ (.Y(_01051_),
    .A(_00978_),
    .B(_01050_));
 sg13g2_nand4_1 _06111_ (.B(_01041_),
    .C(_01048_),
    .A(_01036_),
    .Y(_01052_),
    .D(_01051_));
 sg13g2_nor2_1 _06112_ (.A(_00771_),
    .B(_00776_),
    .Y(_01053_));
 sg13g2_nor2_2 _06113_ (.A(_01024_),
    .B(_01026_),
    .Y(_01054_));
 sg13g2_a21oi_1 _06114_ (.A1(_01024_),
    .A2(_00734_),
    .Y(_01055_),
    .B1(net274));
 sg13g2_o21ai_1 _06115_ (.B1(_00728_),
    .Y(_01056_),
    .A1(_01054_),
    .A2(_01055_));
 sg13g2_buf_1 _06116_ (.A(_01056_),
    .X(_01057_));
 sg13g2_nand4_1 _06117_ (.B(net365),
    .C(net321),
    .A(net366),
    .Y(_01058_),
    .D(net362));
 sg13g2_buf_2 _06118_ (.A(_01058_),
    .X(_01059_));
 sg13g2_or2_1 _06119_ (.X(_01060_),
    .B(_01059_),
    .A(net279));
 sg13g2_nand4_1 _06120_ (.B(_00819_),
    .C(_01057_),
    .A(_01053_),
    .Y(_01061_),
    .D(_01060_));
 sg13g2_buf_1 _06121_ (.A(net285),
    .X(_01062_));
 sg13g2_nor3_1 _06122_ (.A(net232),
    .B(net239),
    .C(_00671_),
    .Y(_01063_));
 sg13g2_buf_1 _06123_ (.A(_00790_),
    .X(_01064_));
 sg13g2_a221oi_1 _06124_ (.B2(net231),
    .C1(_00807_),
    .B1(_00730_),
    .A1(net245),
    .Y(_01065_),
    .A2(_01063_));
 sg13g2_nor2_1 _06125_ (.A(net275),
    .B(net233),
    .Y(_01066_));
 sg13g2_nor3_1 _06126_ (.A(net274),
    .B(net303),
    .C(_00805_),
    .Y(_01067_));
 sg13g2_o21ai_1 _06127_ (.B1(net245),
    .Y(_01068_),
    .A1(_01066_),
    .A2(_01067_));
 sg13g2_nor2_2 _06128_ (.A(net234),
    .B(net280),
    .Y(_01069_));
 sg13g2_nor2_1 _06129_ (.A(net319),
    .B(_01045_),
    .Y(_01070_));
 sg13g2_buf_2 _06130_ (.A(_01070_),
    .X(_01071_));
 sg13g2_or3_1 _06131_ (.A(net273),
    .B(net315),
    .C(net364),
    .X(_01072_));
 sg13g2_buf_1 _06132_ (.A(_01072_),
    .X(_01073_));
 sg13g2_nand2_1 _06133_ (.Y(_01074_),
    .A(net282),
    .B(_01073_));
 sg13g2_nor4_2 _06134_ (.A(net268),
    .B(net319),
    .C(net322),
    .Y(_01075_),
    .D(net284));
 sg13g2_a221oi_1 _06135_ (.B2(_00766_),
    .C1(_01075_),
    .B1(_01074_),
    .A1(_01069_),
    .Y(_01076_),
    .A2(_01071_));
 sg13g2_nor2_2 _06136_ (.A(net280),
    .B(net268),
    .Y(_01077_));
 sg13g2_nor2_1 _06137_ (.A(_01038_),
    .B(_01026_),
    .Y(_01078_));
 sg13g2_nor2_1 _06138_ (.A(net285),
    .B(net319),
    .Y(_01079_));
 sg13g2_a221oi_1 _06139_ (.B2(_01079_),
    .C1(net242),
    .B1(_01078_),
    .A1(_01077_),
    .Y(_01080_),
    .A2(_00888_));
 sg13g2_buf_1 _06140_ (.A(_01080_),
    .X(_01081_));
 sg13g2_nand4_1 _06141_ (.B(_01068_),
    .C(_01076_),
    .A(_01065_),
    .Y(_01082_),
    .D(_01081_));
 sg13g2_nor3_1 _06142_ (.A(_01052_),
    .B(_01061_),
    .C(_01082_),
    .Y(_01083_));
 sg13g2_buf_1 _06143_ (.A(_01026_),
    .X(_01084_));
 sg13g2_nor3_1 _06144_ (.A(_00916_),
    .B(_00799_),
    .C(net230),
    .Y(_01085_));
 sg13g2_a21oi_1 _06145_ (.A1(_00799_),
    .A2(net244),
    .Y(_01086_),
    .B1(_01085_));
 sg13g2_and2_1 _06146_ (.A(net369),
    .B(_01086_),
    .X(_01087_));
 sg13g2_nor2_1 _06147_ (.A(net271),
    .B(net311),
    .Y(_01088_));
 sg13g2_nor3_1 _06148_ (.A(net268),
    .B(_00878_),
    .C(_01088_),
    .Y(_01089_));
 sg13g2_inv_1 _06149_ (.Y(_01090_),
    .A(_01089_));
 sg13g2_and3_1 _06150_ (.X(_01091_),
    .A(_01036_),
    .B(_01048_),
    .C(_01051_));
 sg13g2_nor2_2 _06151_ (.A(net303),
    .B(_00796_),
    .Y(_01092_));
 sg13g2_nand2_1 _06152_ (.Y(_01093_),
    .A(_01069_),
    .B(_01092_));
 sg13g2_a22oi_1 _06153_ (.Y(_01094_),
    .B1(_00894_),
    .B2(_01093_),
    .A2(_01066_),
    .A1(net369));
 sg13g2_nand3_1 _06154_ (.B(_00674_),
    .C(net185),
    .A(_00657_),
    .Y(_01095_));
 sg13g2_nand3_1 _06155_ (.B(net317),
    .C(_00694_),
    .A(_00638_),
    .Y(_01096_));
 sg13g2_nand2_1 _06156_ (.Y(_01097_),
    .A(net208),
    .B(_01096_));
 sg13g2_a22oi_1 _06157_ (.Y(_01098_),
    .B1(_01097_),
    .B2(_00786_),
    .A2(_00934_),
    .A1(net312));
 sg13g2_nor4_1 _06158_ (.A(_01091_),
    .B(_01094_),
    .C(_01095_),
    .D(_01098_),
    .Y(_01099_));
 sg13g2_a221oi_1 _06159_ (.B2(_01099_),
    .C1(_00967_),
    .B1(_01090_),
    .A1(_01083_),
    .Y(_01100_),
    .A2(_01087_));
 sg13g2_buf_1 _06160_ (.A(_00799_),
    .X(_01101_));
 sg13g2_nand2_1 _06161_ (.Y(_01102_),
    .A(net274),
    .B(net310));
 sg13g2_a21oi_2 _06162_ (.B1(net233),
    .Y(_01103_),
    .A2(_01102_),
    .A1(_00784_));
 sg13g2_nor2_1 _06163_ (.A(net369),
    .B(_00866_),
    .Y(_01104_));
 sg13g2_inv_1 _06164_ (.Y(_01105_),
    .A(_01104_));
 sg13g2_a21oi_1 _06165_ (.A1(net312),
    .A2(_01103_),
    .Y(_01106_),
    .B1(_01105_));
 sg13g2_o21ai_1 _06166_ (.B1(net358),
    .Y(_01107_),
    .A1(net267),
    .A2(_01106_));
 sg13g2_nand2_1 _06167_ (.Y(_01108_),
    .A(_00874_),
    .B(_01107_));
 sg13g2_nor2_1 _06168_ (.A(_00885_),
    .B(net207),
    .Y(_01109_));
 sg13g2_o21ai_1 _06169_ (.B1(net281),
    .Y(_01110_),
    .A1(net243),
    .A2(_00915_));
 sg13g2_buf_1 _06170_ (.A(_00979_),
    .X(_01111_));
 sg13g2_nand3b_1 _06171_ (.B(_01110_),
    .C(net204),
    .Y(_01112_),
    .A_N(_01039_));
 sg13g2_nor2b_1 _06172_ (.A(net278),
    .B_N(_00811_),
    .Y(_01113_));
 sg13g2_a22oi_1 _06173_ (.Y(_01114_),
    .B1(_01113_),
    .B2(net311),
    .A2(_01112_),
    .A1(_01109_));
 sg13g2_nor2_2 _06174_ (.A(net360),
    .B(_00638_),
    .Y(_01115_));
 sg13g2_nor2b_1 _06175_ (.A(net318),
    .B_N(net310),
    .Y(_01116_));
 sg13g2_buf_1 _06176_ (.A(_01116_),
    .X(_01117_));
 sg13g2_nand3_1 _06177_ (.B(net271),
    .C(_01117_),
    .A(net275),
    .Y(_01118_));
 sg13g2_buf_1 _06178_ (.A(_01118_),
    .X(_01119_));
 sg13g2_nor2_2 _06179_ (.A(net283),
    .B(net182),
    .Y(_01120_));
 sg13g2_nor3_1 _06180_ (.A(net275),
    .B(net285),
    .C(net278),
    .Y(_01121_));
 sg13g2_a221oi_1 _06181_ (.B2(_01120_),
    .C1(_01121_),
    .B1(_01115_),
    .A1(_00885_),
    .Y(_01122_),
    .A2(_00829_));
 sg13g2_buf_1 _06182_ (.A(_00915_),
    .X(_01123_));
 sg13g2_nor3_2 _06183_ (.A(net229),
    .B(net303),
    .C(net278),
    .Y(_01124_));
 sg13g2_nor2_1 _06184_ (.A(_00874_),
    .B(_01124_),
    .Y(_01125_));
 sg13g2_nand2_1 _06185_ (.Y(_01126_),
    .A(net231),
    .B(net207));
 sg13g2_nand3_1 _06186_ (.B(_00655_),
    .C(net207),
    .A(_00703_),
    .Y(_01127_));
 sg13g2_buf_1 _06187_ (.A(_01127_),
    .X(_01128_));
 sg13g2_a21o_1 _06188_ (.A2(_01128_),
    .A1(_01126_),
    .B1(net324),
    .X(_01129_));
 sg13g2_nand4_1 _06189_ (.B(_01122_),
    .C(_01125_),
    .A(_01114_),
    .Y(_01130_),
    .D(_01129_));
 sg13g2_o21ai_1 _06190_ (.B1(_01130_),
    .Y(_01131_),
    .A1(_01100_),
    .A2(_01108_));
 sg13g2_or2_1 _06191_ (.X(_01132_),
    .B(\z80.tv80s.i_tv80_core.ISet[3] ),
    .A(\z80.tv80s.i_tv80_core.ISet[1] ));
 sg13g2_o21ai_1 _06192_ (.B1(_00866_),
    .Y(_01133_),
    .A1(net359),
    .A2(_01132_));
 sg13g2_buf_1 _06193_ (.A(_01133_),
    .X(_01134_));
 sg13g2_inv_1 _06194_ (.Y(_01135_),
    .A(_01134_));
 sg13g2_a21oi_1 _06195_ (.A1(_01035_),
    .A2(_01131_),
    .Y(_01136_),
    .B1(_01135_));
 sg13g2_buf_1 _06196_ (.A(_01136_),
    .X(_01137_));
 sg13g2_nor4_2 _06197_ (.A(net323),
    .B(net286),
    .C(_01045_),
    .Y(_01138_),
    .D(_00805_));
 sg13g2_nand2_1 _06198_ (.Y(_01139_),
    .A(_00923_),
    .B(_01138_));
 sg13g2_o21ai_1 _06199_ (.B1(_01139_),
    .Y(_01140_),
    .A1(_01052_),
    .A2(_01138_));
 sg13g2_buf_1 _06200_ (.A(net245),
    .X(_01141_));
 sg13g2_nand2_1 _06201_ (.Y(_01142_),
    .A(net203),
    .B(_00815_));
 sg13g2_a21oi_1 _06202_ (.A1(_00639_),
    .A2(net210),
    .Y(_01143_),
    .B1(_01115_));
 sg13g2_nor2_1 _06203_ (.A(_01142_),
    .B(_01143_),
    .Y(_01144_));
 sg13g2_o21ai_1 _06204_ (.B1(_00923_),
    .Y(_01145_),
    .A1(net395),
    .A2(_00850_));
 sg13g2_buf_1 _06205_ (.A(_01145_),
    .X(_01146_));
 sg13g2_nand2_1 _06206_ (.Y(_01147_),
    .A(net311),
    .B(_00923_));
 sg13g2_o21ai_1 _06207_ (.B1(_00674_),
    .Y(_01148_),
    .A1(_01093_),
    .A2(_01147_));
 sg13g2_and2_1 _06208_ (.A(_01146_),
    .B(_01148_),
    .X(_01149_));
 sg13g2_nor3_1 _06209_ (.A(net314),
    .B(net286),
    .C(_00668_),
    .Y(_01150_));
 sg13g2_buf_2 _06210_ (.A(_01150_),
    .X(_01151_));
 sg13g2_nand3_1 _06211_ (.B(_00843_),
    .C(net239),
    .A(net231),
    .Y(_01152_));
 sg13g2_a21oi_2 _06212_ (.B1(net234),
    .Y(_01153_),
    .A2(_01152_),
    .A1(net240));
 sg13g2_o21ai_1 _06213_ (.B1(_01115_),
    .Y(_01154_),
    .A1(_01151_),
    .A2(_01153_));
 sg13g2_nand2_1 _06214_ (.Y(_01155_),
    .A(_00703_),
    .B(_00881_));
 sg13g2_buf_2 _06215_ (.A(_01155_),
    .X(_01156_));
 sg13g2_a21oi_1 _06216_ (.A1(_00922_),
    .A2(_01156_),
    .Y(_01157_),
    .B1(net185));
 sg13g2_nor4_1 _06217_ (.A(_00862_),
    .B(net355),
    .C(net208),
    .D(_01157_),
    .Y(_01158_));
 sg13g2_nand4_1 _06218_ (.B(_01090_),
    .C(_01154_),
    .A(_01051_),
    .Y(_01159_),
    .D(_01158_));
 sg13g2_or4_1 _06219_ (.A(_01140_),
    .B(_01144_),
    .C(_01149_),
    .D(_01159_),
    .X(_01160_));
 sg13g2_buf_1 _06220_ (.A(_00923_),
    .X(_01161_));
 sg13g2_nor2b_1 _06221_ (.A(net395),
    .B_N(_00023_),
    .Y(_01162_));
 sg13g2_a21oi_1 _06222_ (.A1(net357),
    .A2(_00701_),
    .Y(_01163_),
    .B1(_01162_));
 sg13g2_a21oi_1 _06223_ (.A1(net351),
    .A2(_01163_),
    .Y(_01164_),
    .B1(_00657_));
 sg13g2_nand3_1 _06224_ (.B(net231),
    .C(_00979_),
    .A(net323),
    .Y(_01165_));
 sg13g2_buf_1 _06225_ (.A(_01165_),
    .X(_01166_));
 sg13g2_nor2_1 _06226_ (.A(net369),
    .B(_01166_),
    .Y(_01167_));
 sg13g2_xnor2_1 _06227_ (.Y(_01168_),
    .A(net316),
    .B(net313));
 sg13g2_and2_1 _06228_ (.A(_00896_),
    .B(_01168_),
    .X(_01169_));
 sg13g2_nand2b_1 _06229_ (.Y(_01170_),
    .B(net360),
    .A_N(_00638_));
 sg13g2_buf_1 _06230_ (.A(_01170_),
    .X(_01171_));
 sg13g2_buf_1 _06231_ (.A(_01171_),
    .X(_01172_));
 sg13g2_o21ai_1 _06232_ (.B1(net228),
    .Y(_01173_),
    .A1(_01167_),
    .A2(_01169_));
 sg13g2_o21ai_1 _06233_ (.B1(net232),
    .Y(_01174_),
    .A1(net369),
    .A2(net233));
 sg13g2_nand2_1 _06234_ (.Y(_01175_),
    .A(_00981_),
    .B(_01125_));
 sg13g2_a21oi_1 _06235_ (.A1(net183),
    .A2(_01174_),
    .Y(_01176_),
    .B1(_01175_));
 sg13g2_nand3_1 _06236_ (.B(_01173_),
    .C(_01176_),
    .A(_01114_),
    .Y(_01177_));
 sg13g2_o21ai_1 _06237_ (.B1(_01177_),
    .Y(_01178_),
    .A1(_01160_),
    .A2(_01164_));
 sg13g2_buf_1 _06238_ (.A(_01178_),
    .X(_01179_));
 sg13g2_a21o_1 _06239_ (.A2(_01087_),
    .A1(_01083_),
    .B1(net355),
    .X(_01180_));
 sg13g2_nor2_1 _06240_ (.A(_00813_),
    .B(_01037_),
    .Y(_01181_));
 sg13g2_nor2b_1 _06241_ (.A(_01181_),
    .B_N(_01040_),
    .Y(_01182_));
 sg13g2_or3_1 _06242_ (.A(_01094_),
    .B(_01095_),
    .C(_01098_),
    .X(_01183_));
 sg13g2_inv_1 _06243_ (.Y(_01184_),
    .A(_01146_));
 sg13g2_nor2_2 _06244_ (.A(_01042_),
    .B(_00796_),
    .Y(_01185_));
 sg13g2_a21oi_1 _06245_ (.A1(_00820_),
    .A2(_01185_),
    .Y(_01186_),
    .B1(_00821_));
 sg13g2_mux2_1 _06246_ (.A0(_01184_),
    .A1(_01186_),
    .S(net307),
    .X(_01187_));
 sg13g2_nand2_1 _06247_ (.Y(_01188_),
    .A(_00842_),
    .B(_01044_));
 sg13g2_a221oi_1 _06248_ (.B2(net271),
    .C1(_01188_),
    .B1(_01187_),
    .A1(net369),
    .Y(_01189_),
    .A2(net239));
 sg13g2_nor4_1 _06249_ (.A(_01182_),
    .B(_01183_),
    .C(_01140_),
    .D(_01189_),
    .Y(_01190_));
 sg13g2_nor2_2 _06250_ (.A(net281),
    .B(net182),
    .Y(_01191_));
 sg13g2_a22oi_1 _06251_ (.Y(_01192_),
    .B1(_01191_),
    .B2(net311),
    .A2(_01146_),
    .A1(_01124_));
 sg13g2_nand3_1 _06252_ (.B(_01122_),
    .C(_01192_),
    .A(_01114_),
    .Y(_01193_));
 sg13g2_nand2_1 _06253_ (.Y(_01194_),
    .A(_01035_),
    .B(_01107_));
 sg13g2_a21oi_1 _06254_ (.A1(_00870_),
    .A2(_01193_),
    .Y(_01195_),
    .B1(_01194_));
 sg13g2_o21ai_1 _06255_ (.B1(_01195_),
    .Y(_01196_),
    .A1(_01180_),
    .A2(_01190_));
 sg13g2_buf_1 _06256_ (.A(_01196_),
    .X(_01197_));
 sg13g2_o21ai_1 _06257_ (.B1(_01134_),
    .Y(_01198_),
    .A1(_01179_),
    .A2(_01197_));
 sg13g2_buf_1 _06258_ (.A(_01198_),
    .X(_01199_));
 sg13g2_nor2b_1 _06259_ (.A(_01137_),
    .B_N(_01199_),
    .Y(_01200_));
 sg13g2_buf_2 _06260_ (.A(_01200_),
    .X(_01201_));
 sg13g2_o21ai_1 _06261_ (.B1(net238),
    .Y(_01202_),
    .A1(net242),
    .A2(_01028_));
 sg13g2_nor2b_1 _06262_ (.A(_01201_),
    .B_N(_01202_),
    .Y(_01203_));
 sg13g2_nor3_1 _06263_ (.A(_01028_),
    .B(_01034_),
    .C(_01203_),
    .Y(_01204_));
 sg13g2_nor2_1 _06264_ (.A(_01034_),
    .B(_01203_),
    .Y(_01205_));
 sg13g2_buf_1 _06265_ (.A(_01205_),
    .X(_01206_));
 sg13g2_o21ai_1 _06266_ (.B1(_01002_),
    .Y(_01207_),
    .A1(_01013_),
    .A2(net72));
 sg13g2_buf_1 _06267_ (.A(_01207_),
    .X(_01208_));
 sg13g2_or4_1 _06268_ (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ),
    .B(\z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ),
    .C(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ),
    .D(\z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ),
    .X(_01209_));
 sg13g2_a22oi_1 _06269_ (.Y(_01210_),
    .B1(net58),
    .B2(_01209_),
    .A2(_01204_),
    .A1(_01023_));
 sg13g2_inv_1 _06270_ (.Y(_00017_),
    .A(_01210_));
 sg13g2_inv_1 _06271_ (.Y(_01211_),
    .A(_01013_));
 sg13g2_nor2_1 _06272_ (.A(_01018_),
    .B(_01028_),
    .Y(_01212_));
 sg13g2_a22oi_1 _06273_ (.Y(_01213_),
    .B1(_01212_),
    .B2(_01002_),
    .A2(_01028_),
    .A1(_01211_));
 sg13g2_nor2b_1 _06274_ (.A(_01213_),
    .B_N(net72),
    .Y(_01214_));
 sg13g2_or4_1 _06275_ (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ),
    .B(\z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ),
    .C(\z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ),
    .D(\z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ),
    .X(_01215_));
 sg13g2_buf_1 _06276_ (.A(_00901_),
    .X(_01216_));
 sg13g2_nand2_1 _06277_ (.Y(_01217_),
    .A(net354),
    .B(net302));
 sg13g2_and2_1 _06278_ (.A(_00990_),
    .B(_01217_),
    .X(_01218_));
 sg13g2_nand2_1 _06279_ (.Y(_01219_),
    .A(_01002_),
    .B(_01204_));
 sg13g2_buf_2 _06280_ (.A(_01219_),
    .X(_01220_));
 sg13g2_a21oi_1 _06281_ (.A1(_01007_),
    .A2(_01218_),
    .Y(_01221_),
    .B1(_01220_));
 sg13g2_a21oi_1 _06282_ (.A1(_01208_),
    .A2(_01215_),
    .Y(_01222_),
    .B1(_01221_));
 sg13g2_nand2b_1 _06283_ (.Y(_00018_),
    .B(_01222_),
    .A_N(_01214_));
 sg13g2_nand2_1 _06284_ (.Y(_01223_),
    .A(_00852_),
    .B(_01004_));
 sg13g2_nand2_1 _06285_ (.Y(_01224_),
    .A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ),
    .B(net58));
 sg13g2_o21ai_1 _06286_ (.B1(_01224_),
    .Y(_00009_),
    .A1(_01223_),
    .A2(_01220_));
 sg13g2_or3_1 _06287_ (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ),
    .B(\z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ),
    .C(\z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ),
    .X(_01225_));
 sg13g2_nand2_1 _06288_ (.Y(_01226_),
    .A(_01015_),
    .B(_01019_));
 sg13g2_a21oi_1 _06289_ (.A1(_01226_),
    .A2(_01218_),
    .Y(_01227_),
    .B1(_01220_));
 sg13g2_a21oi_1 _06290_ (.A1(_01208_),
    .A2(_01225_),
    .Y(_01228_),
    .B1(_01227_));
 sg13g2_nand2b_1 _06291_ (.Y(_00019_),
    .B(_01228_),
    .A_N(_00009_));
 sg13g2_buf_1 _06292_ (.A(_00874_),
    .X(_01229_));
 sg13g2_buf_1 _06293_ (.A(net359),
    .X(_01230_));
 sg13g2_buf_1 _06294_ (.A(net301),
    .X(_01231_));
 sg13g2_nand3_1 _06295_ (.B(_01044_),
    .C(_01054_),
    .A(net265),
    .Y(_01232_));
 sg13g2_o21ai_1 _06296_ (.B1(_01232_),
    .Y(_01233_),
    .A1(net266),
    .A2(_01109_));
 sg13g2_nor2b_1 _06297_ (.A(_00998_),
    .B_N(net399),
    .Y(_01234_));
 sg13g2_buf_1 _06298_ (.A(_01234_),
    .X(_01235_));
 sg13g2_buf_1 _06299_ (.A(_01235_),
    .X(_01236_));
 sg13g2_buf_1 _06300_ (.A(net264),
    .X(_01237_));
 sg13g2_mux2_1 _06301_ (.A0(\z80.tv80s.i_tv80_core.mcycles[1] ),
    .A1(_01233_),
    .S(net227),
    .X(_00012_));
 sg13g2_buf_1 _06302_ (.A(net264),
    .X(_01238_));
 sg13g2_nand2_1 _06303_ (.Y(_01239_),
    .A(net265),
    .B(net226));
 sg13g2_o21ai_1 _06304_ (.B1(_01102_),
    .Y(_01240_),
    .A1(net229),
    .A2(net279));
 sg13g2_nor2_1 _06305_ (.A(_00786_),
    .B(net184),
    .Y(_01241_));
 sg13g2_a221oi_1 _06306_ (.B2(_00877_),
    .C1(_01241_),
    .B1(_01240_),
    .A1(net204),
    .Y(_01242_),
    .A2(_01086_));
 sg13g2_nand2b_1 _06307_ (.Y(_01243_),
    .B(_00635_),
    .A_N(_00998_));
 sg13g2_buf_1 _06308_ (.A(_01243_),
    .X(_01244_));
 sg13g2_buf_1 _06309_ (.A(_01244_),
    .X(_01245_));
 sg13g2_buf_1 _06310_ (.A(net263),
    .X(_01246_));
 sg13g2_buf_1 _06311_ (.A(net276),
    .X(_01247_));
 sg13g2_and2_1 _06312_ (.A(net229),
    .B(net358),
    .X(_01248_));
 sg13g2_a22oi_1 _06313_ (.Y(_01249_),
    .B1(_01248_),
    .B2(_00877_),
    .A2(_01247_),
    .A1(_00811_));
 sg13g2_nor3_1 _06314_ (.A(net236),
    .B(net225),
    .C(_01249_),
    .Y(_01250_));
 sg13g2_and2_1 _06315_ (.A(\z80.tv80s.i_tv80_core.mcycles[2] ),
    .B(net225),
    .X(_01251_));
 sg13g2_buf_1 _06316_ (.A(net308),
    .X(_01252_));
 sg13g2_buf_1 _06317_ (.A(_00760_),
    .X(_01253_));
 sg13g2_buf_1 _06318_ (.A(\z80.tv80s.i_tv80_core.F[0] ),
    .X(_01254_));
 sg13g2_inv_1 _06319_ (.Y(_01255_),
    .A(net391));
 sg13g2_nor2_1 _06320_ (.A(net261),
    .B(_01255_),
    .Y(_01256_));
 sg13g2_a21oi_1 _06321_ (.A1(net261),
    .A2(net397),
    .Y(_01257_),
    .B1(_01256_));
 sg13g2_xnor2_1 _06322_ (.Y(_01258_),
    .A(net262),
    .B(_01257_));
 sg13g2_buf_1 _06323_ (.A(net271),
    .X(_01259_));
 sg13g2_buf_1 _06324_ (.A(net305),
    .X(_01260_));
 sg13g2_nor2_2 _06325_ (.A(net260),
    .B(net263),
    .Y(_01261_));
 sg13g2_and4_1 _06326_ (.A(net223),
    .B(net206),
    .C(_00953_),
    .D(_01261_),
    .X(_01262_));
 sg13g2_nor2b_1 _06327_ (.A(_01258_),
    .B_N(_01262_),
    .Y(_01263_));
 sg13g2_nor3_1 _06328_ (.A(_01250_),
    .B(_01251_),
    .C(_01263_),
    .Y(_01264_));
 sg13g2_o21ai_1 _06329_ (.B1(_01264_),
    .Y(_00013_),
    .A1(_01239_),
    .A2(_01242_));
 sg13g2_nor2_1 _06330_ (.A(\z80.tv80s.i_tv80_core.mcycles[4] ),
    .B(net226),
    .Y(_01265_));
 sg13g2_buf_1 _06331_ (.A(_01245_),
    .X(_01266_));
 sg13g2_buf_1 _06332_ (.A(net222),
    .X(_01267_));
 sg13g2_inv_1 _06333_ (.Y(_01268_),
    .A(_00825_));
 sg13g2_nor3_1 _06334_ (.A(_01268_),
    .B(net394),
    .C(net185),
    .Y(_01269_));
 sg13g2_nor3_1 _06335_ (.A(_00769_),
    .B(net205),
    .C(_01269_),
    .Y(_01270_));
 sg13g2_a21oi_1 _06336_ (.A1(_00674_),
    .A2(_01270_),
    .Y(_01271_),
    .B1(net260));
 sg13g2_and2_1 _06337_ (.A(net276),
    .B(_01124_),
    .X(_01272_));
 sg13g2_buf_1 _06338_ (.A(_01272_),
    .X(_01273_));
 sg13g2_nor3_1 _06339_ (.A(net202),
    .B(_01271_),
    .C(_01273_),
    .Y(_01274_));
 sg13g2_o21ai_1 _06340_ (.B1(net241),
    .Y(_01275_),
    .A1(_00971_),
    .A2(net210));
 sg13g2_nand3_1 _06341_ (.B(_01261_),
    .C(_01275_),
    .A(_00680_),
    .Y(_01276_));
 sg13g2_o21ai_1 _06342_ (.B1(_01276_),
    .Y(_00014_),
    .A1(_01265_),
    .A2(_01274_));
 sg13g2_buf_1 _06343_ (.A(net202),
    .X(_01277_));
 sg13g2_buf_1 _06344_ (.A(net358),
    .X(_01278_));
 sg13g2_nand2_2 _06345_ (.Y(_01279_),
    .A(_01044_),
    .B(net204));
 sg13g2_nand2_1 _06346_ (.Y(_01280_),
    .A(_01279_),
    .B(_01166_));
 sg13g2_inv_1 _06347_ (.Y(_01281_),
    .A(_00971_));
 sg13g2_nand3b_1 _06348_ (.B(net361),
    .C(net318),
    .Y(_01282_),
    .A_N(_00702_));
 sg13g2_nor3_2 _06349_ (.A(net275),
    .B(_00678_),
    .C(_01282_),
    .Y(_01283_));
 sg13g2_nand3_1 _06350_ (.B(net210),
    .C(_01283_),
    .A(_01281_),
    .Y(_01284_));
 sg13g2_buf_1 _06351_ (.A(net238),
    .X(_01285_));
 sg13g2_buf_1 _06352_ (.A(_01285_),
    .X(_01286_));
 sg13g2_a21oi_1 _06353_ (.A1(_01286_),
    .A2(net210),
    .Y(_01287_),
    .B1(_01142_));
 sg13g2_or4_1 _06354_ (.A(net318),
    .B(_00714_),
    .C(_00716_),
    .D(_00717_),
    .X(_01288_));
 sg13g2_buf_1 _06355_ (.A(_01288_),
    .X(_01289_));
 sg13g2_buf_1 _06356_ (.A(net244),
    .X(_01290_));
 sg13g2_a21oi_1 _06357_ (.A1(_00786_),
    .A2(_01289_),
    .Y(_01291_),
    .B1(net200));
 sg13g2_nor2_1 _06358_ (.A(net209),
    .B(_01138_),
    .Y(_01292_));
 sg13g2_o21ai_1 _06359_ (.B1(_00831_),
    .Y(_01293_),
    .A1(_00916_),
    .A2(_01038_));
 sg13g2_nand2_1 _06360_ (.Y(_01294_),
    .A(net231),
    .B(_01293_));
 sg13g2_buf_1 _06361_ (.A(_00780_),
    .X(_01295_));
 sg13g2_inv_1 _06362_ (.Y(_01296_),
    .A(net351));
 sg13g2_o21ai_1 _06363_ (.B1(_00805_),
    .Y(_01297_),
    .A1(net259),
    .A2(_01296_));
 sg13g2_and2_1 _06364_ (.A(_00766_),
    .B(_01074_),
    .X(_01298_));
 sg13g2_a21oi_1 _06365_ (.A1(_00953_),
    .A2(_01297_),
    .Y(_01299_),
    .B1(_01298_));
 sg13g2_nand3_1 _06366_ (.B(_01294_),
    .C(_01299_),
    .A(_01292_),
    .Y(_01300_));
 sg13g2_nor4_1 _06367_ (.A(_01153_),
    .B(_01287_),
    .C(_01291_),
    .D(_01300_),
    .Y(_01301_));
 sg13g2_a21oi_1 _06368_ (.A1(_01284_),
    .A2(_01301_),
    .Y(_01302_),
    .B1(net260));
 sg13g2_a221oi_1 _06369_ (.B2(net224),
    .C1(_01302_),
    .B1(_01280_),
    .A1(net300),
    .Y(_01303_),
    .A2(_01103_));
 sg13g2_and3_1 _06370_ (.X(_01304_),
    .A(net394),
    .B(_00833_),
    .C(_01261_));
 sg13g2_a221oi_1 _06371_ (.B2(_01258_),
    .C1(_01304_),
    .B1(_01262_),
    .A1(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .Y(_01305_),
    .A2(net202));
 sg13g2_o21ai_1 _06372_ (.B1(_01305_),
    .Y(_00015_),
    .A1(_01277_),
    .A2(_01303_));
 sg13g2_inv_1 _06373_ (.Y(_01306_),
    .A(\z80.tv80s.i_tv80_core.ISet[1] ));
 sg13g2_buf_2 _06374_ (.A(_00024_),
    .X(_01307_));
 sg13g2_nor2_1 _06375_ (.A(\z80.tv80s.i_tv80_core.ts[1] ),
    .B(net398),
    .Y(_01308_));
 sg13g2_buf_1 _06376_ (.A(net311),
    .X(_01309_));
 sg13g2_a21oi_1 _06377_ (.A1(_01307_),
    .A2(_01308_),
    .Y(_01310_),
    .B1(net258));
 sg13g2_and2_1 _06378_ (.A(net398),
    .B(net2),
    .X(_01311_));
 sg13g2_buf_1 _06379_ (.A(_01311_),
    .X(_01312_));
 sg13g2_nand2_1 _06380_ (.Y(_01313_),
    .A(_00635_),
    .B(_01312_));
 sg13g2_buf_1 _06381_ (.A(_01313_),
    .X(_01314_));
 sg13g2_nor2_1 _06382_ (.A(_00998_),
    .B(_01314_),
    .Y(_01315_));
 sg13g2_and2_1 _06383_ (.A(_01310_),
    .B(_01315_),
    .X(_01316_));
 sg13g2_buf_1 _06384_ (.A(_01316_),
    .X(_01317_));
 sg13g2_nand2_1 _06385_ (.Y(_01318_),
    .A(net398),
    .B(net2));
 sg13g2_buf_2 _06386_ (.A(_01318_),
    .X(_01319_));
 sg13g2_nor2_2 _06387_ (.A(net258),
    .B(_01319_),
    .Y(_01320_));
 sg13g2_nand4_1 _06388_ (.B(_00672_),
    .C(_01261_),
    .A(_01069_),
    .Y(_01321_),
    .D(_01320_));
 sg13g2_o21ai_1 _06389_ (.B1(_01321_),
    .Y(_00000_),
    .A1(_01306_),
    .A2(_01317_));
 sg13g2_nand2_1 _06390_ (.Y(_01322_),
    .A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ),
    .B(net58));
 sg13g2_o21ai_1 _06391_ (.B1(_01322_),
    .Y(_00005_),
    .A1(_01226_),
    .A2(_01220_));
 sg13g2_a21o_1 _06392_ (.A2(net58),
    .A1(\z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ),
    .B1(_01214_),
    .X(_00006_));
 sg13g2_nand2_1 _06393_ (.Y(_01323_),
    .A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ),
    .B(net58));
 sg13g2_o21ai_1 _06394_ (.B1(_01323_),
    .Y(_00007_),
    .A1(_01220_),
    .A2(_01217_));
 sg13g2_a22oi_1 _06395_ (.Y(_01324_),
    .B1(net58),
    .B2(\z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ),
    .A2(_01204_),
    .A1(_01022_));
 sg13g2_inv_1 _06396_ (.Y(_00008_),
    .A(_01324_));
 sg13g2_nand2_1 _06397_ (.Y(_01325_),
    .A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ),
    .B(net58));
 sg13g2_o21ai_1 _06398_ (.B1(_01325_),
    .Y(_00010_),
    .A1(_01007_),
    .A2(_01220_));
 sg13g2_nand2_1 _06399_ (.Y(_01326_),
    .A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ),
    .B(net58));
 sg13g2_o21ai_1 _06400_ (.B1(_01326_),
    .Y(_00011_),
    .A1(_00990_),
    .A2(_01220_));
 sg13g2_nor2b_2 _06401_ (.A(_00743_),
    .B_N(net313),
    .Y(_01327_));
 sg13g2_and2_1 _06402_ (.A(net315),
    .B(_00681_),
    .X(_01328_));
 sg13g2_buf_2 _06403_ (.A(_01328_),
    .X(_01329_));
 sg13g2_buf_1 _06404_ (.A(_01329_),
    .X(_01330_));
 sg13g2_buf_1 _06405_ (.A(_00931_),
    .X(_01331_));
 sg13g2_buf_1 _06406_ (.A(net257),
    .X(_01332_));
 sg13g2_nand2_1 _06407_ (.Y(_01333_),
    .A(net220),
    .B(_00744_));
 sg13g2_a22oi_1 _06408_ (.Y(_01334_),
    .B1(_01333_),
    .B2(net243),
    .A2(net199),
    .A1(_01327_));
 sg13g2_nand2_1 _06409_ (.Y(_01335_),
    .A(net204),
    .B(net276));
 sg13g2_nor4_1 _06410_ (.A(_00741_),
    .B(net222),
    .C(_01334_),
    .D(_01335_),
    .Y(_01336_));
 sg13g2_nor4_1 _06411_ (.A(net267),
    .B(_00696_),
    .C(net222),
    .D(_01335_),
    .Y(_01337_));
 sg13g2_nor2_1 _06412_ (.A(\z80.tv80s.i_tv80_core.IStatus[2] ),
    .B(_01337_),
    .Y(_01338_));
 sg13g2_nor2_1 _06413_ (.A(_01336_),
    .B(_01338_),
    .Y(_00004_));
 sg13g2_nor2_1 _06414_ (.A(\z80.tv80s.i_tv80_core.IStatus[1] ),
    .B(_01336_),
    .Y(_01339_));
 sg13g2_nor2_1 _06415_ (.A(_01337_),
    .B(_01339_),
    .Y(_00003_));
 sg13g2_buf_1 _06416_ (.A(_01310_),
    .X(_01340_));
 sg13g2_buf_1 _06417_ (.A(_01340_),
    .X(_01341_));
 sg13g2_nand2_1 _06418_ (.Y(_01342_),
    .A(net179),
    .B(_01315_));
 sg13g2_and2_1 _06419_ (.A(\z80.tv80s.i_tv80_core.ISet[3] ),
    .B(_01342_),
    .X(_00002_));
 sg13g2_nand4_1 _06420_ (.B(net203),
    .C(_01071_),
    .A(net265),
    .Y(_01343_),
    .D(net239));
 sg13g2_buf_1 _06421_ (.A(_01343_),
    .X(_01344_));
 sg13g2_nor2_1 _06422_ (.A(_01244_),
    .B(_01310_),
    .Y(_01345_));
 sg13g2_buf_2 _06423_ (.A(_01345_),
    .X(_01346_));
 sg13g2_nand2_1 _06424_ (.Y(_01347_),
    .A(net354),
    .B(_01346_));
 sg13g2_nand2_1 _06425_ (.Y(_01348_),
    .A(_00843_),
    .B(_00728_));
 sg13g2_nand2_1 _06426_ (.Y(_01349_),
    .A(net245),
    .B(_00756_));
 sg13g2_nor4_1 _06427_ (.A(net260),
    .B(_01348_),
    .C(_01349_),
    .D(_01342_),
    .Y(_01350_));
 sg13g2_a21oi_1 _06428_ (.A1(net300),
    .A2(_01342_),
    .Y(_01351_),
    .B1(_01350_));
 sg13g2_o21ai_1 _06429_ (.B1(_01351_),
    .Y(_00001_),
    .A1(_01344_),
    .A2(_01347_));
 sg13g2_nor2_2 _06430_ (.A(net233),
    .B(_00784_),
    .Y(_01352_));
 sg13g2_nor2_1 _06431_ (.A(net309),
    .B(_01156_),
    .Y(_01353_));
 sg13g2_buf_2 _06432_ (.A(_01353_),
    .X(_01354_));
 sg13g2_a22oi_1 _06433_ (.Y(_01355_),
    .B1(_00719_),
    .B2(_01354_),
    .A2(_01352_),
    .A1(_01281_));
 sg13g2_nor2_1 _06434_ (.A(net200),
    .B(_01355_),
    .Y(_01356_));
 sg13g2_nand2_2 _06435_ (.Y(_01357_),
    .A(_00728_),
    .B(_00740_));
 sg13g2_nor2_1 _06436_ (.A(_00660_),
    .B(_00805_),
    .Y(_01358_));
 sg13g2_buf_2 _06437_ (.A(_01358_),
    .X(_01359_));
 sg13g2_a21oi_1 _06438_ (.A1(_00971_),
    .A2(_00853_),
    .Y(_01360_),
    .B1(_01156_));
 sg13g2_a22oi_1 _06439_ (.Y(_01361_),
    .B1(_01360_),
    .B2(_01069_),
    .A2(_00824_),
    .A1(_01359_));
 sg13g2_nand2_1 _06440_ (.Y(_01362_),
    .A(_01077_),
    .B(_01185_));
 sg13g2_nand2_1 _06441_ (.Y(_01363_),
    .A(_00674_),
    .B(_01362_));
 sg13g2_nor2_2 _06442_ (.A(_00925_),
    .B(_01005_),
    .Y(_01364_));
 sg13g2_o21ai_1 _06443_ (.B1(_01364_),
    .Y(_01365_),
    .A1(_00680_),
    .A2(_01363_));
 sg13g2_o21ai_1 _06444_ (.B1(_01365_),
    .Y(_01366_),
    .A1(_01357_),
    .A2(_01361_));
 sg13g2_nand2_1 _06445_ (.Y(_01367_),
    .A(_00842_),
    .B(_01185_));
 sg13g2_nand2_1 _06446_ (.Y(_01368_),
    .A(net306),
    .B(net309));
 sg13g2_nor2_2 _06447_ (.A(_00851_),
    .B(_01368_),
    .Y(_01369_));
 sg13g2_nor2_1 _06448_ (.A(_00950_),
    .B(net272),
    .Y(_01370_));
 sg13g2_buf_2 _06449_ (.A(_01370_),
    .X(_01371_));
 sg13g2_nand2_1 _06450_ (.Y(_01372_),
    .A(net257),
    .B(_01371_));
 sg13g2_o21ai_1 _06451_ (.B1(_01372_),
    .Y(_01373_),
    .A1(net257),
    .A2(net351));
 sg13g2_a22oi_1 _06452_ (.Y(_01374_),
    .B1(_01373_),
    .B2(net259),
    .A2(_01369_),
    .A1(net199));
 sg13g2_nor2b_1 _06453_ (.A(_00738_),
    .B_N(_00743_),
    .Y(_01375_));
 sg13g2_nor4_2 _06454_ (.A(_00748_),
    .B(_00676_),
    .C(net286),
    .Y(_01376_),
    .D(_01375_));
 sg13g2_nor2_1 _06455_ (.A(_00638_),
    .B(net277),
    .Y(_01377_));
 sg13g2_o21ai_1 _06456_ (.B1(_01377_),
    .Y(_01378_),
    .A1(_00962_),
    .A2(_01376_));
 sg13g2_o21ai_1 _06457_ (.B1(_01378_),
    .Y(_01379_),
    .A1(_01367_),
    .A2(_01374_));
 sg13g2_nand2_1 _06458_ (.Y(_01380_),
    .A(net267),
    .B(_01083_));
 sg13g2_nor3_1 _06459_ (.A(_01161_),
    .B(net200),
    .C(_01380_),
    .Y(_01381_));
 sg13g2_nor4_1 _06460_ (.A(_01356_),
    .B(_01366_),
    .C(_01379_),
    .D(_01381_),
    .Y(_01382_));
 sg13g2_nor2_1 _06461_ (.A(net229),
    .B(net232),
    .Y(_01383_));
 sg13g2_a22oi_1 _06462_ (.Y(_01384_),
    .B1(_01364_),
    .B2(_01092_),
    .A2(_01371_),
    .A1(_01383_));
 sg13g2_nand3_1 _06463_ (.B(_00973_),
    .C(_01354_),
    .A(net232),
    .Y(_01385_));
 sg13g2_o21ai_1 _06464_ (.B1(_01385_),
    .Y(_01386_),
    .A1(net236),
    .A2(_01384_));
 sg13g2_and3_1 _06465_ (.X(_01387_),
    .A(net300),
    .B(net241),
    .C(_01104_));
 sg13g2_buf_1 _06466_ (.A(_01368_),
    .X(_01388_));
 sg13g2_nor4_1 _06467_ (.A(_00851_),
    .B(net266),
    .C(_00981_),
    .D(net219),
    .Y(_01389_));
 sg13g2_buf_2 _06468_ (.A(_01389_),
    .X(_01390_));
 sg13g2_a221oi_1 _06469_ (.B2(_01103_),
    .C1(_01390_),
    .B1(_01387_),
    .A1(_01247_),
    .Y(_01391_),
    .A2(_01386_));
 sg13g2_o21ai_1 _06470_ (.B1(_01391_),
    .Y(doe),
    .A1(_00968_),
    .A2(_01382_));
 sg13g2_buf_1 _06471_ (.A(\z80.tv80s.di_reg[0] ),
    .X(_01392_));
 sg13g2_buf_1 _06472_ (.A(_01392_),
    .X(_01393_));
 sg13g2_mux2_1 _06473_ (.A0(net6),
    .A1(net350),
    .S(net221),
    .X(_00278_));
 sg13g2_buf_1 _06474_ (.A(\z80.tv80s.di_reg[1] ),
    .X(_01394_));
 sg13g2_mux2_1 _06475_ (.A0(net7),
    .A1(net390),
    .S(net221),
    .X(_00279_));
 sg13g2_buf_1 _06476_ (.A(\z80.tv80s.di_reg[2] ),
    .X(_01395_));
 sg13g2_mux2_1 _06477_ (.A0(net8),
    .A1(_01395_),
    .S(net221),
    .X(_00280_));
 sg13g2_buf_1 _06478_ (.A(\z80.tv80s.di_reg[3] ),
    .X(_01396_));
 sg13g2_mux2_1 _06479_ (.A0(net9),
    .A1(_01396_),
    .S(net221),
    .X(_00281_));
 sg13g2_buf_1 _06480_ (.A(\z80.tv80s.di_reg[4] ),
    .X(_01397_));
 sg13g2_mux2_1 _06481_ (.A0(net10),
    .A1(_01397_),
    .S(net221),
    .X(_00282_));
 sg13g2_buf_1 _06482_ (.A(\z80.tv80s.di_reg[5] ),
    .X(_01398_));
 sg13g2_mux2_1 _06483_ (.A0(net11),
    .A1(net386),
    .S(net221),
    .X(_00283_));
 sg13g2_buf_1 _06484_ (.A(\z80.tv80s.di_reg[6] ),
    .X(_01399_));
 sg13g2_mux2_1 _06485_ (.A0(net12),
    .A1(net385),
    .S(net221),
    .X(_00284_));
 sg13g2_buf_1 _06486_ (.A(\z80.tv80s.di_reg[7] ),
    .X(_01400_));
 sg13g2_buf_1 _06487_ (.A(_01400_),
    .X(_01401_));
 sg13g2_mux2_1 _06488_ (.A0(net13),
    .A1(net349),
    .S(net221),
    .X(_00285_));
 sg13g2_buf_1 _06489_ (.A(\z80.tv80s.i_tv80_core.BusB[0] ),
    .X(_01402_));
 sg13g2_buf_1 _06490_ (.A(_01402_),
    .X(_01403_));
 sg13g2_or2_1 _06491_ (.X(_01404_),
    .B(_01138_),
    .A(net209));
 sg13g2_xnor2_1 _06492_ (.Y(_01405_),
    .A(net364),
    .B(net318));
 sg13g2_nor2_1 _06493_ (.A(net314),
    .B(net280),
    .Y(_01406_));
 sg13g2_nand3_1 _06494_ (.B(_00894_),
    .C(_00815_),
    .A(_00788_),
    .Y(_01407_));
 sg13g2_a221oi_1 _06495_ (.B2(net318),
    .C1(_01407_),
    .B1(_01406_),
    .A1(_00780_),
    .Y(_01408_),
    .A2(_01405_));
 sg13g2_nand2_1 _06496_ (.Y(_01409_),
    .A(net308),
    .B(net269));
 sg13g2_nor2b_2 _06497_ (.A(_00742_),
    .B_N(net364),
    .Y(_01410_));
 sg13g2_nor2_1 _06498_ (.A(net316),
    .B(_01410_),
    .Y(_01411_));
 sg13g2_nor2_1 _06499_ (.A(_00653_),
    .B(net321),
    .Y(_01412_));
 sg13g2_nand2_1 _06500_ (.Y(_01413_),
    .A(_00648_),
    .B(_01412_));
 sg13g2_a21oi_1 _06501_ (.A1(_01409_),
    .A2(_01411_),
    .Y(_01414_),
    .B1(_01413_));
 sg13g2_nand2_1 _06502_ (.Y(_01415_),
    .A(_00790_),
    .B(_00792_));
 sg13g2_a21oi_1 _06503_ (.A1(_01415_),
    .A2(_01357_),
    .Y(_01416_),
    .B1(_01349_));
 sg13g2_nor4_1 _06504_ (.A(_01404_),
    .B(_01408_),
    .C(_01414_),
    .D(_01416_),
    .Y(_01417_));
 sg13g2_buf_2 _06505_ (.A(_01417_),
    .X(_01418_));
 sg13g2_nand3_1 _06506_ (.B(_01289_),
    .C(_01418_),
    .A(net185),
    .Y(_01419_));
 sg13g2_buf_1 _06507_ (.A(_01419_),
    .X(_01420_));
 sg13g2_nor4_2 _06508_ (.A(net314),
    .B(net280),
    .C(net320),
    .Y(_01421_),
    .D(_00775_));
 sg13g2_nor4_2 _06509_ (.A(net355),
    .B(net242),
    .C(_00735_),
    .Y(_01422_),
    .D(_01421_));
 sg13g2_nor2_1 _06510_ (.A(_00732_),
    .B(_00680_),
    .Y(_01423_));
 sg13g2_nor2_1 _06511_ (.A(net279),
    .B(_01059_),
    .Y(_01424_));
 sg13g2_nor3_1 _06512_ (.A(net319),
    .B(net303),
    .C(_00734_),
    .Y(_01425_));
 sg13g2_nor4_2 _06513_ (.A(net314),
    .B(net320),
    .C(_00775_),
    .Y(_01426_),
    .D(_01026_));
 sg13g2_nor3_1 _06514_ (.A(net303),
    .B(_00796_),
    .C(_00734_),
    .Y(_01427_));
 sg13g2_nor4_1 _06515_ (.A(_01424_),
    .B(_01425_),
    .C(_01426_),
    .D(_01427_),
    .Y(_01428_));
 sg13g2_nor2_1 _06516_ (.A(_00708_),
    .B(_00775_),
    .Y(_01429_));
 sg13g2_nand2_1 _06517_ (.Y(_01430_),
    .A(net308),
    .B(net315));
 sg13g2_nand3_1 _06518_ (.B(_00744_),
    .C(_01430_),
    .A(_01429_),
    .Y(_01431_));
 sg13g2_nand4_1 _06519_ (.B(_01423_),
    .C(_01428_),
    .A(_01422_),
    .Y(_01432_),
    .D(_01431_));
 sg13g2_buf_2 _06520_ (.A(_01432_),
    .X(_01433_));
 sg13g2_nor2_1 _06521_ (.A(_00803_),
    .B(_01075_),
    .Y(_01434_));
 sg13g2_nor2_1 _06522_ (.A(_00807_),
    .B(net205),
    .Y(_01435_));
 sg13g2_nand2_1 _06523_ (.Y(_01436_),
    .A(_01434_),
    .B(_01435_));
 sg13g2_nor2_1 _06524_ (.A(net229),
    .B(_00713_),
    .Y(_01437_));
 sg13g2_a21oi_1 _06525_ (.A1(net229),
    .A2(net310),
    .Y(_01438_),
    .B1(_01437_));
 sg13g2_and2_1 _06526_ (.A(net283),
    .B(_01327_),
    .X(_01439_));
 sg13g2_o21ai_1 _06527_ (.B1(_01439_),
    .Y(_01440_),
    .A1(net310),
    .A2(_01437_));
 sg13g2_o21ai_1 _06528_ (.B1(_01440_),
    .Y(_01441_),
    .A1(_01042_),
    .A2(_01438_));
 sg13g2_nor3_1 _06529_ (.A(_01117_),
    .B(_01436_),
    .C(_01441_),
    .Y(_01442_));
 sg13g2_nand3_1 _06530_ (.B(net203),
    .C(_01079_),
    .A(_00760_),
    .Y(_01443_));
 sg13g2_buf_1 _06531_ (.A(_01443_),
    .X(_01444_));
 sg13g2_o21ai_1 _06532_ (.B1(net203),
    .Y(_01445_),
    .A1(_00888_),
    .A2(_01063_));
 sg13g2_nand4_1 _06533_ (.B(_01442_),
    .C(_01444_),
    .A(_00786_),
    .Y(_01446_),
    .D(_01445_));
 sg13g2_nor3_1 _06534_ (.A(_01420_),
    .B(_01433_),
    .C(_01446_),
    .Y(_01447_));
 sg13g2_and3_1 _06535_ (.X(_01448_),
    .A(net267),
    .B(net200),
    .C(_01447_));
 sg13g2_buf_2 _06536_ (.A(_01448_),
    .X(_01449_));
 sg13g2_buf_1 _06537_ (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_01450_));
 sg13g2_inv_1 _06538_ (.Y(_01451_),
    .A(_01450_));
 sg13g2_inv_1 _06539_ (.Y(_01452_),
    .A(_01392_));
 sg13g2_buf_2 _06540_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_01453_));
 sg13g2_buf_1 _06541_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .X(_01454_));
 sg13g2_buf_1 _06542_ (.A(_01454_),
    .X(_01455_));
 sg13g2_buf_1 _06543_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(_01456_));
 sg13g2_buf_1 _06544_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .X(_01457_));
 sg13g2_buf_1 _06545_ (.A(_01457_),
    .X(_01458_));
 sg13g2_nand3_1 _06546_ (.B(net384),
    .C(net345),
    .A(net346),
    .Y(_01459_));
 sg13g2_nand2_1 _06547_ (.Y(_01460_),
    .A(_01453_),
    .B(_01459_));
 sg13g2_buf_1 _06548_ (.A(_01460_),
    .X(_01461_));
 sg13g2_buf_1 _06549_ (.A(net384),
    .X(_01462_));
 sg13g2_nand2_1 _06550_ (.Y(_01463_),
    .A(net346),
    .B(net345));
 sg13g2_buf_1 _06551_ (.A(_00194_),
    .X(_01464_));
 sg13g2_xor2_1 _06552_ (.B(net348),
    .A(net382),
    .X(_01465_));
 sg13g2_nor2_1 _06553_ (.A(net345),
    .B(_00208_),
    .Y(_01466_));
 sg13g2_buf_1 _06554_ (.A(_01466_),
    .X(_01467_));
 sg13g2_buf_2 _06555_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .X(_01468_));
 sg13g2_xor2_1 _06556_ (.B(net348),
    .A(_01468_),
    .X(_01469_));
 sg13g2_nor2_1 _06557_ (.A(_01255_),
    .B(net346),
    .Y(_01470_));
 sg13g2_a22oi_1 _06558_ (.Y(_01471_),
    .B1(_01465_),
    .B2(_01470_),
    .A2(_01469_),
    .A1(net256));
 sg13g2_o21ai_1 _06559_ (.B1(_01471_),
    .Y(_01472_),
    .A1(_01463_),
    .A2(_01465_));
 sg13g2_a21oi_1 _06560_ (.A1(net391),
    .A2(net344),
    .Y(_01473_),
    .B1(_01465_));
 sg13g2_inv_1 _06561_ (.Y(_01474_),
    .A(_01454_));
 sg13g2_inv_1 _06562_ (.Y(_01475_),
    .A(net384));
 sg13g2_buf_1 _06563_ (.A(_01475_),
    .X(_01476_));
 sg13g2_inv_1 _06564_ (.Y(_01477_),
    .A(_01468_));
 sg13g2_buf_1 _06565_ (.A(net345),
    .X(_01478_));
 sg13g2_a22oi_1 _06566_ (.Y(_01479_),
    .B1(net348),
    .B2(_01467_),
    .A2(net298),
    .A1(_01455_));
 sg13g2_nand3_1 _06567_ (.B(_01478_),
    .C(net348),
    .A(_01455_),
    .Y(_01480_));
 sg13g2_o21ai_1 _06568_ (.B1(_01480_),
    .Y(_01481_),
    .A1(_01477_),
    .A2(_01479_));
 sg13g2_and2_1 _06569_ (.A(_01476_),
    .B(_01481_),
    .X(_01482_));
 sg13g2_a221oi_1 _06570_ (.B2(_01474_),
    .C1(_01482_),
    .B1(_01473_),
    .A1(net344),
    .Y(_01483_),
    .A2(_01472_));
 sg13g2_inv_1 _06571_ (.Y(_01484_),
    .A(_01483_));
 sg13g2_nand2_1 _06572_ (.Y(_01485_),
    .A(net218),
    .B(_01484_));
 sg13g2_nor2_1 _06573_ (.A(net384),
    .B(_01458_),
    .Y(_01486_));
 sg13g2_inv_1 _06574_ (.Y(_01487_),
    .A(_01453_));
 sg13g2_nor2_1 _06575_ (.A(_01487_),
    .B(net346),
    .Y(_01488_));
 sg13g2_and2_1 _06576_ (.A(_01486_),
    .B(_01488_),
    .X(_01489_));
 sg13g2_buf_2 _06577_ (.A(_01489_),
    .X(_01490_));
 sg13g2_buf_1 _06578_ (.A(net273),
    .X(_01491_));
 sg13g2_buf_1 _06579_ (.A(_00192_),
    .X(_01492_));
 sg13g2_buf_1 _06580_ (.A(_00193_),
    .X(_01493_));
 sg13g2_inv_2 _06581_ (.Y(_01494_),
    .A(net381));
 sg13g2_nand2_1 _06582_ (.Y(_01495_),
    .A(net396),
    .B(_01255_));
 sg13g2_a221oi_1 _06583_ (.B2(net307),
    .C1(net217),
    .B1(_01495_),
    .A1(_01494_),
    .Y(_01496_),
    .A2(net239));
 sg13g2_a21oi_1 _06584_ (.A1(net217),
    .A2(_01492_),
    .Y(_01497_),
    .B1(_01496_));
 sg13g2_and2_1 _06585_ (.A(_01490_),
    .B(_01497_),
    .X(_01498_));
 sg13g2_buf_1 _06586_ (.A(_00204_),
    .X(_01499_));
 sg13g2_nand2_1 _06587_ (.Y(_01500_),
    .A(_01475_),
    .B(net345));
 sg13g2_inv_1 _06588_ (.Y(_01501_),
    .A(net383));
 sg13g2_buf_1 _06589_ (.A(_01501_),
    .X(_01502_));
 sg13g2_nand2_1 _06590_ (.Y(_01503_),
    .A(net384),
    .B(_01502_));
 sg13g2_buf_1 _06591_ (.A(_01503_),
    .X(_01504_));
 sg13g2_nand2_1 _06592_ (.Y(_01505_),
    .A(_01453_),
    .B(net346));
 sg13g2_a21oi_1 _06593_ (.A1(_01500_),
    .A2(_01504_),
    .Y(_01506_),
    .B1(_01505_));
 sg13g2_buf_2 _06594_ (.A(_01506_),
    .X(_01507_));
 sg13g2_inv_1 _06595_ (.Y(_01508_),
    .A(_01507_));
 sg13g2_nor3_1 _06596_ (.A(_01476_),
    .B(_01499_),
    .C(_01508_),
    .Y(_01509_));
 sg13g2_nand3_1 _06597_ (.B(net346),
    .C(_01486_),
    .A(_01453_),
    .Y(_01510_));
 sg13g2_buf_2 _06598_ (.A(_01510_),
    .X(_01511_));
 sg13g2_buf_1 _06599_ (.A(_01450_),
    .X(_01512_));
 sg13g2_o21ai_1 _06600_ (.B1(_01512_),
    .Y(_01513_),
    .A1(net382),
    .A2(_01511_));
 sg13g2_buf_1 _06601_ (.A(_01462_),
    .X(_01514_));
 sg13g2_nand2_1 _06602_ (.Y(_01515_),
    .A(_01458_),
    .B(_01488_));
 sg13g2_buf_2 _06603_ (.A(_01515_),
    .X(_01516_));
 sg13g2_nor3_1 _06604_ (.A(_01514_),
    .B(_01073_),
    .C(_01516_),
    .Y(_01517_));
 sg13g2_or3_1 _06605_ (.A(_01509_),
    .B(_01513_),
    .C(_01517_),
    .X(_01518_));
 sg13g2_buf_1 _06606_ (.A(_00200_),
    .X(_01519_));
 sg13g2_nand2_1 _06607_ (.Y(_01520_),
    .A(_01478_),
    .B(_01073_));
 sg13g2_o21ai_1 _06608_ (.B1(_01520_),
    .Y(_01521_),
    .A1(_01073_),
    .A2(_01504_));
 sg13g2_nor2_1 _06609_ (.A(net384),
    .B(_01463_),
    .Y(_01522_));
 sg13g2_buf_2 _06610_ (.A(_01522_),
    .X(_01523_));
 sg13g2_a21oi_1 _06611_ (.A1(_01474_),
    .A2(_01521_),
    .Y(_01524_),
    .B1(_01523_));
 sg13g2_nor3_1 _06612_ (.A(_01487_),
    .B(_01519_),
    .C(_01524_),
    .Y(_01525_));
 sg13g2_nor3_1 _06613_ (.A(_01498_),
    .B(_01518_),
    .C(_01525_),
    .Y(_01526_));
 sg13g2_a221oi_1 _06614_ (.B2(_01526_),
    .C1(_01449_),
    .B1(_01485_),
    .A1(_01451_),
    .Y(_01527_),
    .A2(_01452_));
 sg13g2_a21oi_2 _06615_ (.B1(_01527_),
    .Y(_01528_),
    .A2(_01449_),
    .A1(net348));
 sg13g2_inv_1 _06616_ (.Y(_01529_),
    .A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ));
 sg13g2_buf_1 _06617_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ),
    .X(_01530_));
 sg13g2_nor3_1 _06618_ (.A(net347),
    .B(_01453_),
    .C(_01459_),
    .Y(_01531_));
 sg13g2_a21oi_1 _06619_ (.A1(\z80.tv80s.i_tv80_core.ts[1] ),
    .A2(_00209_),
    .Y(_01532_),
    .B1(net343));
 sg13g2_nor2_1 _06620_ (.A(_01531_),
    .B(_01532_),
    .Y(_01533_));
 sg13g2_nand2_1 _06621_ (.Y(_01534_),
    .A(_01530_),
    .B(_01533_));
 sg13g2_inv_1 _06622_ (.Y(_01535_),
    .A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ));
 sg13g2_nand2_1 _06623_ (.Y(_01536_),
    .A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ),
    .B(_01535_));
 sg13g2_or4_1 _06624_ (.A(_01529_),
    .B(_00210_),
    .C(_01534_),
    .D(_01536_),
    .X(_01537_));
 sg13g2_buf_1 _06625_ (.A(_01537_),
    .X(_01538_));
 sg13g2_buf_1 _06626_ (.A(_01538_),
    .X(_01539_));
 sg13g2_buf_1 _06627_ (.A(_00909_),
    .X(_01540_));
 sg13g2_nand4_1 _06628_ (.B(_01540_),
    .C(net276),
    .A(net257),
    .Y(_01541_),
    .D(_00987_));
 sg13g2_buf_1 _06629_ (.A(_01541_),
    .X(_01542_));
 sg13g2_buf_1 _06630_ (.A(_01542_),
    .X(_01543_));
 sg13g2_buf_1 _06631_ (.A(net155),
    .X(_01544_));
 sg13g2_buf_2 _06632_ (.A(\z80.tv80s.i_tv80_core.ACC[0] ),
    .X(_01545_));
 sg13g2_or2_1 _06633_ (.X(_01546_),
    .B(net205),
    .A(_00807_));
 sg13g2_buf_1 _06634_ (.A(_01546_),
    .X(_01547_));
 sg13g2_nor3_1 _06635_ (.A(_00802_),
    .B(_01420_),
    .C(_01547_),
    .Y(_01548_));
 sg13g2_nand2_1 _06636_ (.Y(_01549_),
    .A(_01069_),
    .B(_01071_));
 sg13g2_nand3_1 _06637_ (.B(net231),
    .C(_00792_),
    .A(net315),
    .Y(_01550_));
 sg13g2_nand3_1 _06638_ (.B(_00889_),
    .C(_01550_),
    .A(_00917_),
    .Y(_01551_));
 sg13g2_and2_1 _06639_ (.A(net318),
    .B(_01551_),
    .X(_01552_));
 sg13g2_buf_1 _06640_ (.A(_01552_),
    .X(_01553_));
 sg13g2_nor2_2 _06641_ (.A(_00768_),
    .B(_00710_),
    .Y(_01554_));
 sg13g2_nor2_1 _06642_ (.A(net269),
    .B(net320),
    .Y(_01555_));
 sg13g2_nor3_1 _06643_ (.A(net233),
    .B(_00773_),
    .C(_00796_),
    .Y(_01556_));
 sg13g2_a221oi_1 _06644_ (.B2(_01555_),
    .C1(_01556_),
    .B1(_01554_),
    .A1(_00672_),
    .Y(_01557_),
    .A2(_01359_));
 sg13g2_buf_1 _06645_ (.A(_01557_),
    .X(_01558_));
 sg13g2_inv_1 _06646_ (.Y(_01559_),
    .A(_01558_));
 sg13g2_nor2_1 _06647_ (.A(_00875_),
    .B(_00780_),
    .Y(_01560_));
 sg13g2_a22oi_1 _06648_ (.Y(_01561_),
    .B1(_01560_),
    .B2(net281),
    .A2(_00811_),
    .A1(_00683_));
 sg13g2_nand2_1 _06649_ (.Y(_01562_),
    .A(net282),
    .B(net245));
 sg13g2_nor4_1 _06650_ (.A(net268),
    .B(_00796_),
    .C(_01026_),
    .D(_01168_),
    .Y(_01563_));
 sg13g2_nor2_1 _06651_ (.A(_01352_),
    .B(_01563_),
    .Y(_01564_));
 sg13g2_o21ai_1 _06652_ (.B1(_01564_),
    .Y(_01565_),
    .A1(_01561_),
    .A2(_01562_));
 sg13g2_nor4_2 _06653_ (.A(_01433_),
    .B(_01553_),
    .C(_01559_),
    .Y(_01566_),
    .D(_01565_));
 sg13g2_buf_8 _06654_ (.A(_01566_),
    .X(_01567_));
 sg13g2_a22oi_1 _06655_ (.Y(_01568_),
    .B1(_01327_),
    .B2(net283),
    .A2(_00877_),
    .A1(net315));
 sg13g2_nor4_1 _06656_ (.A(net323),
    .B(net320),
    .C(_01329_),
    .D(_01568_),
    .Y(_01569_));
 sg13g2_nor2_1 _06657_ (.A(_01151_),
    .B(_01569_),
    .Y(_01570_));
 sg13g2_buf_1 _06658_ (.A(_01570_),
    .X(_01571_));
 sg13g2_and3_1 _06659_ (.X(_01572_),
    .A(_01549_),
    .B(_01567_),
    .C(_01571_));
 sg13g2_buf_1 _06660_ (.A(_01572_),
    .X(_01573_));
 sg13g2_and2_1 _06661_ (.A(_01548_),
    .B(_01573_),
    .X(_01574_));
 sg13g2_buf_1 _06662_ (.A(_01574_),
    .X(_01575_));
 sg13g2_buf_1 _06663_ (.A(_01575_),
    .X(_01576_));
 sg13g2_nand3_1 _06664_ (.B(net278),
    .C(_00793_),
    .A(_00786_),
    .Y(_01577_));
 sg13g2_buf_1 _06665_ (.A(_01577_),
    .X(_01578_));
 sg13g2_or4_1 _06666_ (.A(_01578_),
    .B(_01117_),
    .C(_01436_),
    .D(_01441_),
    .X(_01579_));
 sg13g2_or2_1 _06667_ (.X(_01580_),
    .B(_01579_),
    .A(_01420_));
 sg13g2_buf_1 _06668_ (.A(_01580_),
    .X(_01581_));
 sg13g2_nand2_1 _06669_ (.Y(_01582_),
    .A(net203),
    .B(_00888_));
 sg13g2_nand3_1 _06670_ (.B(_01444_),
    .C(_01582_),
    .A(_00657_),
    .Y(_01583_));
 sg13g2_buf_1 _06671_ (.A(_01583_),
    .X(_01584_));
 sg13g2_nand2_1 _06672_ (.Y(_01585_),
    .A(_00728_),
    .B(_00730_));
 sg13g2_o21ai_1 _06673_ (.B1(_01585_),
    .Y(_01586_),
    .A1(net279),
    .A2(net240));
 sg13g2_nor3_1 _06674_ (.A(net229),
    .B(net303),
    .C(_00734_),
    .Y(_01587_));
 sg13g2_nor4_1 _06675_ (.A(_01581_),
    .B(_01584_),
    .C(_01586_),
    .D(_01587_),
    .Y(_01588_));
 sg13g2_nand2_1 _06676_ (.Y(_01589_),
    .A(_00888_),
    .B(_01054_));
 sg13g2_nand3_1 _06677_ (.B(_01588_),
    .C(_01589_),
    .A(_01422_),
    .Y(_01590_));
 sg13g2_buf_1 _06678_ (.A(_01590_),
    .X(_01591_));
 sg13g2_nor2b_1 _06679_ (.A(_01591_),
    .B_N(_00995_),
    .Y(_01592_));
 sg13g2_nand2_2 _06680_ (.Y(_01593_),
    .A(_01307_),
    .B(_01308_));
 sg13g2_nand2_2 _06681_ (.Y(_01594_),
    .A(net238),
    .B(_01593_));
 sg13g2_buf_1 _06682_ (.A(_01594_),
    .X(_01595_));
 sg13g2_o21ai_1 _06683_ (.B1(net178),
    .Y(_01596_),
    .A1(net130),
    .A2(_01592_));
 sg13g2_buf_2 _06684_ (.A(_01596_),
    .X(_01597_));
 sg13g2_nand2b_1 _06685_ (.Y(_01598_),
    .B(_01592_),
    .A_N(_01575_));
 sg13g2_buf_2 _06686_ (.A(_01598_),
    .X(_01599_));
 sg13g2_buf_1 _06687_ (.A(_01575_),
    .X(_01600_));
 sg13g2_nand2_1 _06688_ (.Y(_01601_),
    .A(\z80.tv80s.i_tv80_core.Ap[0] ),
    .B(net129));
 sg13g2_o21ai_1 _06689_ (.B1(_01601_),
    .Y(_01602_),
    .A1(_01545_),
    .A2(_01599_));
 sg13g2_buf_1 _06690_ (.A(net178),
    .X(_01603_));
 sg13g2_a22oi_1 _06691_ (.Y(_01604_),
    .B1(_01602_),
    .B2(_01603_),
    .A2(_01597_),
    .A1(_01545_));
 sg13g2_buf_1 _06692_ (.A(\z80.tv80s.i_tv80_core.I[0] ),
    .X(_01605_));
 sg13g2_buf_1 _06693_ (.A(\z80.tv80s.i_tv80_core.R[0] ),
    .X(_01606_));
 sg13g2_nor3_1 _06694_ (.A(net223),
    .B(_01059_),
    .C(_01335_),
    .Y(_01607_));
 sg13g2_buf_1 _06695_ (.A(_01607_),
    .X(_01608_));
 sg13g2_mux2_1 _06696_ (.A0(_01605_),
    .A1(_01606_),
    .S(_01608_),
    .X(_01609_));
 sg13g2_nor2_1 _06697_ (.A(net155),
    .B(_01609_),
    .Y(_01610_));
 sg13g2_a21oi_1 _06698_ (.A1(net152),
    .A2(_01604_),
    .Y(_01611_),
    .B1(_01610_));
 sg13g2_nand2_1 _06699_ (.Y(_01612_),
    .A(_01539_),
    .B(_01611_));
 sg13g2_o21ai_1 _06700_ (.B1(_01612_),
    .Y(_01613_),
    .A1(_01528_),
    .A2(_01539_));
 sg13g2_buf_1 _06701_ (.A(_01245_),
    .X(_01614_));
 sg13g2_buf_1 _06702_ (.A(net216),
    .X(_01615_));
 sg13g2_nand2_1 _06703_ (.Y(_01616_),
    .A(_00221_),
    .B(net197));
 sg13g2_o21ai_1 _06704_ (.B1(_01616_),
    .Y(_00286_),
    .A1(net181),
    .A2(_01613_));
 sg13g2_and2_1 _06705_ (.A(_01453_),
    .B(_01459_),
    .X(_01617_));
 sg13g2_buf_1 _06706_ (.A(_01617_),
    .X(_01618_));
 sg13g2_nand2_2 _06707_ (.Y(_01619_),
    .A(net384),
    .B(net298));
 sg13g2_and2_1 _06708_ (.A(net346),
    .B(_01619_),
    .X(_01620_));
 sg13g2_buf_1 _06709_ (.A(_01620_),
    .X(_01621_));
 sg13g2_nor2b_1 _06710_ (.A(net383),
    .B_N(_01402_),
    .Y(_01622_));
 sg13g2_nor2b_1 _06711_ (.A(_01403_),
    .B_N(net383),
    .Y(_01623_));
 sg13g2_nand3b_1 _06712_ (.B(_01456_),
    .C(net391),
    .Y(_01624_),
    .A_N(_01454_));
 sg13g2_buf_1 _06713_ (.A(_01624_),
    .X(_01625_));
 sg13g2_mux2_1 _06714_ (.A0(_01622_),
    .A1(_01623_),
    .S(_01625_),
    .X(_01626_));
 sg13g2_and2_1 _06715_ (.A(net382),
    .B(_01626_),
    .X(_01627_));
 sg13g2_nor2b_1 _06716_ (.A(net382),
    .B_N(_01402_),
    .Y(_01628_));
 sg13g2_nor2b_1 _06717_ (.A(_01402_),
    .B_N(_01468_),
    .Y(_01629_));
 sg13g2_a21o_1 _06718_ (.A2(_01625_),
    .A1(_01628_),
    .B1(_01629_),
    .X(_01630_));
 sg13g2_or2_1 _06719_ (.X(_01631_),
    .B(_01402_),
    .A(net382));
 sg13g2_nand2_1 _06720_ (.Y(_01632_),
    .A(_01468_),
    .B(_01403_));
 sg13g2_o21ai_1 _06721_ (.B1(_01632_),
    .Y(_01633_),
    .A1(_01625_),
    .A2(_01631_));
 sg13g2_mux2_1 _06722_ (.A0(_01630_),
    .A1(_01633_),
    .S(_01501_),
    .X(_01634_));
 sg13g2_buf_1 _06723_ (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .X(_01635_));
 sg13g2_buf_2 _06724_ (.A(\z80.tv80s.i_tv80_core.BusB[1] ),
    .X(_01636_));
 sg13g2_xnor2_1 _06725_ (.Y(_01637_),
    .A(_01635_),
    .B(_01636_));
 sg13g2_xnor2_1 _06726_ (.Y(_01638_),
    .A(net383),
    .B(_01637_));
 sg13g2_o21ai_1 _06727_ (.B1(_01638_),
    .Y(_01639_),
    .A1(_01627_),
    .A2(_01634_));
 sg13g2_or3_1 _06728_ (.A(_01627_),
    .B(_01634_),
    .C(_01638_),
    .X(_01640_));
 sg13g2_nand2_1 _06729_ (.Y(_01641_),
    .A(_01639_),
    .B(_01640_));
 sg13g2_buf_1 _06730_ (.A(_01635_),
    .X(_01642_));
 sg13g2_nand3_1 _06731_ (.B(net342),
    .C(_01636_),
    .A(_01475_),
    .Y(_01643_));
 sg13g2_o21ai_1 _06732_ (.B1(_01643_),
    .Y(_01644_),
    .A1(net299),
    .A2(_01637_));
 sg13g2_or2_1 _06733_ (.X(_01645_),
    .B(_01636_),
    .A(net342));
 sg13g2_a22oi_1 _06734_ (.Y(_01646_),
    .B1(_01645_),
    .B2(_01523_),
    .A2(_01644_),
    .A1(net256));
 sg13g2_o21ai_1 _06735_ (.B1(_01646_),
    .Y(_01647_),
    .A1(_01621_),
    .A2(_01641_));
 sg13g2_buf_1 _06736_ (.A(_00201_),
    .X(_01648_));
 sg13g2_nor2b_1 _06737_ (.A(net344),
    .B_N(_01648_),
    .Y(_01649_));
 sg13g2_buf_2 _06738_ (.A(_00205_),
    .X(_01650_));
 sg13g2_and2_1 _06739_ (.A(net344),
    .B(_01650_),
    .X(_01651_));
 sg13g2_nor2_1 _06740_ (.A(_01649_),
    .B(_01651_),
    .Y(_01652_));
 sg13g2_buf_2 _06741_ (.A(\z80.tv80s.i_tv80_core.F[4] ),
    .X(_01653_));
 sg13g2_inv_1 _06742_ (.Y(_01654_),
    .A(_01653_));
 sg13g2_buf_1 _06743_ (.A(\z80.tv80s.i_tv80_core.BusA[2] ),
    .X(_01655_));
 sg13g2_buf_1 _06744_ (.A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(_01656_));
 sg13g2_o21ai_1 _06745_ (.B1(_01656_),
    .Y(_01657_),
    .A1(_01655_),
    .A2(_01635_));
 sg13g2_buf_2 _06746_ (.A(_01657_),
    .X(_01658_));
 sg13g2_nand2_1 _06747_ (.Y(_01659_),
    .A(_01654_),
    .B(_01658_));
 sg13g2_buf_2 _06748_ (.A(_01659_),
    .X(_01660_));
 sg13g2_xor2_1 _06749_ (.B(_01660_),
    .A(net342),
    .X(_01661_));
 sg13g2_nor3_2 _06750_ (.A(net344),
    .B(net298),
    .C(_01505_),
    .Y(_01662_));
 sg13g2_nand2_1 _06751_ (.Y(_01663_),
    .A(_01453_),
    .B(_01474_));
 sg13g2_or2_1 _06752_ (.X(_01664_),
    .B(_01504_),
    .A(_01663_));
 sg13g2_buf_1 _06753_ (.A(_01664_),
    .X(_01665_));
 sg13g2_nand2_1 _06754_ (.Y(_01666_),
    .A(net396),
    .B(_00683_));
 sg13g2_inv_1 _06755_ (.Y(_01667_),
    .A(_01666_));
 sg13g2_mux2_1 _06756_ (.A0(_01516_),
    .A1(_01665_),
    .S(_01667_),
    .X(_01668_));
 sg13g2_nor2_1 _06757_ (.A(_01462_),
    .B(_01516_),
    .Y(_01669_));
 sg13g2_buf_2 _06758_ (.A(_00195_),
    .X(_01670_));
 sg13g2_nand2b_1 _06759_ (.Y(_01671_),
    .B(net273),
    .A_N(_01670_));
 sg13g2_o21ai_1 _06760_ (.B1(_01671_),
    .Y(_01672_),
    .A1(net273),
    .A2(_01464_));
 sg13g2_a221oi_1 _06761_ (.B2(_01490_),
    .C1(net218),
    .B1(_01672_),
    .A1(_01669_),
    .Y(_01673_),
    .A2(_01667_));
 sg13g2_o21ai_1 _06762_ (.B1(_01673_),
    .Y(_01674_),
    .A1(_01648_),
    .A2(_01668_));
 sg13g2_a221oi_1 _06763_ (.B2(_01662_),
    .C1(_01674_),
    .B1(_01661_),
    .A1(_01507_),
    .Y(_01675_),
    .A2(_01652_));
 sg13g2_inv_1 _06764_ (.Y(_01676_),
    .A(_01675_));
 sg13g2_o21ai_1 _06765_ (.B1(_01676_),
    .Y(_01677_),
    .A1(_01618_),
    .A2(_01647_));
 sg13g2_nand2_1 _06766_ (.Y(_01678_),
    .A(net347),
    .B(net390));
 sg13g2_o21ai_1 _06767_ (.B1(_01678_),
    .Y(_01679_),
    .A1(net347),
    .A2(_01677_));
 sg13g2_mux2_1 _06768_ (.A0(_01679_),
    .A1(_01636_),
    .S(_01449_),
    .X(_01680_));
 sg13g2_buf_1 _06769_ (.A(_01680_),
    .X(_01681_));
 sg13g2_inv_1 _06770_ (.Y(_01682_),
    .A(_01681_));
 sg13g2_buf_2 _06771_ (.A(\z80.tv80s.i_tv80_core.ACC[1] ),
    .X(_01683_));
 sg13g2_nand2_1 _06772_ (.Y(_01684_),
    .A(\z80.tv80s.i_tv80_core.Ap[1] ),
    .B(net130));
 sg13g2_o21ai_1 _06773_ (.B1(_01684_),
    .Y(_01685_),
    .A1(_01683_),
    .A2(_01599_));
 sg13g2_a22oi_1 _06774_ (.Y(_01686_),
    .B1(_01685_),
    .B2(net169),
    .A2(_01597_),
    .A1(_01683_));
 sg13g2_inv_1 _06775_ (.Y(_01687_),
    .A(\z80.tv80s.i_tv80_core.I[1] ));
 sg13g2_nand2_1 _06776_ (.Y(_01688_),
    .A(\z80.tv80s.i_tv80_core.R[1] ),
    .B(net160));
 sg13g2_o21ai_1 _06777_ (.B1(_01688_),
    .Y(_01689_),
    .A1(_01687_),
    .A2(net160));
 sg13g2_nor2_1 _06778_ (.A(net155),
    .B(_01689_),
    .Y(_01690_));
 sg13g2_a21oi_1 _06779_ (.A1(net152),
    .A2(_01686_),
    .Y(_01691_),
    .B1(_01690_));
 sg13g2_nand2_1 _06780_ (.Y(_01692_),
    .A(net161),
    .B(_01691_));
 sg13g2_o21ai_1 _06781_ (.B1(_01692_),
    .Y(_01693_),
    .A1(net161),
    .A2(_01682_));
 sg13g2_nand2_1 _06782_ (.Y(_01694_),
    .A(_00222_),
    .B(net197));
 sg13g2_o21ai_1 _06783_ (.B1(_01694_),
    .Y(_00287_),
    .A1(net181),
    .A2(_01693_));
 sg13g2_buf_1 _06784_ (.A(_01449_),
    .X(_01695_));
 sg13g2_buf_1 _06785_ (.A(_01655_),
    .X(_01696_));
 sg13g2_buf_1 _06786_ (.A(\z80.tv80s.i_tv80_core.BusB[2] ),
    .X(_01697_));
 sg13g2_nand2_1 _06787_ (.Y(_01698_),
    .A(net341),
    .B(net380));
 sg13g2_xor2_1 _06788_ (.B(net380),
    .A(_01655_),
    .X(_01699_));
 sg13g2_nand2_1 _06789_ (.Y(_01700_),
    .A(net344),
    .B(_01699_));
 sg13g2_o21ai_1 _06790_ (.B1(_01700_),
    .Y(_01701_),
    .A1(net296),
    .A2(_01698_));
 sg13g2_or2_1 _06791_ (.X(_01702_),
    .B(net380),
    .A(net341));
 sg13g2_xor2_1 _06792_ (.B(_01636_),
    .A(net383),
    .X(_01703_));
 sg13g2_nand2b_1 _06793_ (.Y(_01704_),
    .B(_01703_),
    .A_N(_01492_));
 sg13g2_xnor2_1 _06794_ (.Y(_01705_),
    .A(net383),
    .B(_01699_));
 sg13g2_a21oi_1 _06795_ (.A1(_01639_),
    .A2(_01704_),
    .Y(_01706_),
    .B1(_01705_));
 sg13g2_and3_1 _06796_ (.X(_01707_),
    .A(_01639_),
    .B(_01704_),
    .C(_01705_));
 sg13g2_nor3_1 _06797_ (.A(_01621_),
    .B(_01706_),
    .C(_01707_),
    .Y(_01708_));
 sg13g2_a221oi_1 _06798_ (.B2(_01523_),
    .C1(_01708_),
    .B1(_01702_),
    .A1(net256),
    .Y(_01709_),
    .A2(_01701_));
 sg13g2_buf_1 _06799_ (.A(_01709_),
    .X(_01710_));
 sg13g2_nor2_1 _06800_ (.A(_01663_),
    .B(_01504_),
    .Y(_01711_));
 sg13g2_buf_2 _06801_ (.A(_01711_),
    .X(_01712_));
 sg13g2_nor2_1 _06802_ (.A(net317),
    .B(_00933_),
    .Y(_01713_));
 sg13g2_nor2_1 _06803_ (.A(_01516_),
    .B(_01713_),
    .Y(_01714_));
 sg13g2_a21oi_1 _06804_ (.A1(_01712_),
    .A2(_01713_),
    .Y(_01715_),
    .B1(_01714_));
 sg13g2_nor2_1 _06805_ (.A(_00202_),
    .B(_01715_),
    .Y(_01716_));
 sg13g2_buf_2 _06806_ (.A(\z80.tv80s.i_tv80_core.F[1] ),
    .X(_01717_));
 sg13g2_xnor2_1 _06807_ (.Y(_01718_),
    .A(net342),
    .B(_01717_));
 sg13g2_xnor2_1 _06808_ (.Y(_01719_),
    .A(net341),
    .B(_01718_));
 sg13g2_mux2_1 _06809_ (.A0(_01670_),
    .A1(_01719_),
    .S(_01660_),
    .X(_01720_));
 sg13g2_nor2_1 _06810_ (.A(_01511_),
    .B(_01720_),
    .Y(_01721_));
 sg13g2_mux2_1 _06811_ (.A0(_00202_),
    .A1(_00206_),
    .S(net296),
    .X(_01722_));
 sg13g2_buf_2 _06812_ (.A(_00196_),
    .X(_01723_));
 sg13g2_nor2b_1 _06813_ (.A(_01491_),
    .B_N(_01492_),
    .Y(_01724_));
 sg13g2_a21oi_1 _06814_ (.A1(_01491_),
    .A2(_01723_),
    .Y(_01725_),
    .B1(_01724_));
 sg13g2_a221oi_1 _06815_ (.B2(_01490_),
    .C1(net218),
    .B1(_01725_),
    .A1(_01669_),
    .Y(_01726_),
    .A2(_01713_));
 sg13g2_o21ai_1 _06816_ (.B1(_01726_),
    .Y(_01727_),
    .A1(_01508_),
    .A2(_01722_));
 sg13g2_nor3_1 _06817_ (.A(_01716_),
    .B(_01721_),
    .C(_01727_),
    .Y(_01728_));
 sg13g2_a21oi_1 _06818_ (.A1(net218),
    .A2(_01710_),
    .Y(_01729_),
    .B1(_01728_));
 sg13g2_nor2b_1 _06819_ (.A(net343),
    .B_N(\z80.tv80s.di_reg[2] ),
    .Y(_01730_));
 sg13g2_a21oi_1 _06820_ (.A1(net343),
    .A2(_01729_),
    .Y(_01731_),
    .B1(_01730_));
 sg13g2_nand2_1 _06821_ (.Y(_01732_),
    .A(net380),
    .B(_01449_));
 sg13g2_o21ai_1 _06822_ (.B1(_01732_),
    .Y(_01733_),
    .A1(net139),
    .A2(_01731_));
 sg13g2_buf_1 _06823_ (.A(_01733_),
    .X(_01734_));
 sg13g2_inv_1 _06824_ (.Y(_01735_),
    .A(_01734_));
 sg13g2_buf_2 _06825_ (.A(\z80.tv80s.i_tv80_core.ACC[2] ),
    .X(_01736_));
 sg13g2_nand2_1 _06826_ (.Y(_01737_),
    .A(\z80.tv80s.i_tv80_core.Ap[2] ),
    .B(net130));
 sg13g2_o21ai_1 _06827_ (.B1(_01737_),
    .Y(_01738_),
    .A1(_01736_),
    .A2(_01599_));
 sg13g2_a22oi_1 _06828_ (.Y(_01739_),
    .B1(_01738_),
    .B2(net169),
    .A2(_01597_),
    .A1(_01736_));
 sg13g2_buf_1 _06829_ (.A(\z80.tv80s.i_tv80_core.I[2] ),
    .X(_01740_));
 sg13g2_buf_1 _06830_ (.A(\z80.tv80s.i_tv80_core.R[2] ),
    .X(_01741_));
 sg13g2_mux2_1 _06831_ (.A0(_01740_),
    .A1(_01741_),
    .S(net160),
    .X(_01742_));
 sg13g2_nor2_1 _06832_ (.A(net155),
    .B(_01742_),
    .Y(_01743_));
 sg13g2_a21oi_1 _06833_ (.A1(net152),
    .A2(_01739_),
    .Y(_01744_),
    .B1(_01743_));
 sg13g2_nand2_1 _06834_ (.Y(_01745_),
    .A(_01538_),
    .B(_01744_));
 sg13g2_o21ai_1 _06835_ (.B1(_01745_),
    .Y(_01746_),
    .A1(net161),
    .A2(_01735_));
 sg13g2_buf_1 _06836_ (.A(net216),
    .X(_01747_));
 sg13g2_nand2_1 _06837_ (.Y(_01748_),
    .A(_00223_),
    .B(net196));
 sg13g2_o21ai_1 _06838_ (.B1(_01748_),
    .Y(_00288_),
    .A1(net181),
    .A2(_01746_));
 sg13g2_buf_1 _06839_ (.A(net346),
    .X(_01749_));
 sg13g2_nand2_1 _06840_ (.Y(_01750_),
    .A(net294),
    .B(_01619_));
 sg13g2_nor2_1 _06841_ (.A(_01670_),
    .B(net380),
    .Y(_01751_));
 sg13g2_or2_1 _06842_ (.X(_01752_),
    .B(_01751_),
    .A(_01706_));
 sg13g2_nand2b_1 _06843_ (.Y(_01753_),
    .B(_01697_),
    .A_N(_01670_));
 sg13g2_nand2b_1 _06844_ (.Y(_01754_),
    .B(_01753_),
    .A_N(_01706_));
 sg13g2_nor2_1 _06845_ (.A(net298),
    .B(_01754_),
    .Y(_01755_));
 sg13g2_a21oi_1 _06846_ (.A1(net298),
    .A2(_01752_),
    .Y(_01756_),
    .B1(_01755_));
 sg13g2_buf_2 _06847_ (.A(\z80.tv80s.i_tv80_core.BusB[3] ),
    .X(_01757_));
 sg13g2_xnor2_1 _06848_ (.Y(_01758_),
    .A(_01656_),
    .B(_01757_));
 sg13g2_xnor2_1 _06849_ (.Y(_01759_),
    .A(_01756_),
    .B(_01758_));
 sg13g2_buf_1 _06850_ (.A(_01656_),
    .X(_01760_));
 sg13g2_nand3_1 _06851_ (.B(net340),
    .C(_01757_),
    .A(net299),
    .Y(_01761_));
 sg13g2_o21ai_1 _06852_ (.B1(_01761_),
    .Y(_01762_),
    .A1(net299),
    .A2(_01758_));
 sg13g2_o21ai_1 _06853_ (.B1(_01523_),
    .Y(_01763_),
    .A1(net340),
    .A2(_01757_));
 sg13g2_inv_1 _06854_ (.Y(_01764_),
    .A(_01763_));
 sg13g2_a221oi_1 _06855_ (.B2(net256),
    .C1(_01764_),
    .B1(_01762_),
    .A1(_01750_),
    .Y(_01765_),
    .A2(_01759_));
 sg13g2_buf_1 _06856_ (.A(_01765_),
    .X(_01766_));
 sg13g2_inv_1 _06857_ (.Y(_01767_),
    .A(_01656_));
 sg13g2_or2_1 _06858_ (.X(_01768_),
    .B(net342),
    .A(_01655_));
 sg13g2_buf_1 _06859_ (.A(_01768_),
    .X(_01769_));
 sg13g2_nand3_1 _06860_ (.B(_01642_),
    .C(_01717_),
    .A(net341),
    .Y(_01770_));
 sg13g2_o21ai_1 _06861_ (.B1(_01770_),
    .Y(_01771_),
    .A1(_01717_),
    .A2(_01769_));
 sg13g2_nor2_1 _06862_ (.A(_01767_),
    .B(net341),
    .Y(_01772_));
 sg13g2_a22oi_1 _06863_ (.Y(_01773_),
    .B1(_01772_),
    .B2(_01717_),
    .A2(_01771_),
    .A1(_01767_));
 sg13g2_a22oi_1 _06864_ (.Y(_01774_),
    .B1(_01769_),
    .B2(net340),
    .A2(_01654_),
    .A1(_01723_));
 sg13g2_nand4_1 _06865_ (.B(_01696_),
    .C(_01642_),
    .A(net340),
    .Y(_01775_),
    .D(_01717_));
 sg13g2_nand2b_1 _06866_ (.Y(_01776_),
    .B(_01775_),
    .A_N(_01774_));
 sg13g2_o21ai_1 _06867_ (.B1(_01776_),
    .Y(_01777_),
    .A1(_01654_),
    .A2(_01773_));
 sg13g2_buf_1 _06868_ (.A(_00203_),
    .X(_01778_));
 sg13g2_buf_1 _06869_ (.A(_00207_),
    .X(_01779_));
 sg13g2_mux2_1 _06870_ (.A0(_01778_),
    .A1(_01779_),
    .S(net344),
    .X(_01780_));
 sg13g2_inv_1 _06871_ (.Y(_01781_),
    .A(_01780_));
 sg13g2_buf_2 _06872_ (.A(_00197_),
    .X(_01782_));
 sg13g2_inv_1 _06873_ (.Y(_01783_),
    .A(_01782_));
 sg13g2_nand2_1 _06874_ (.Y(_01784_),
    .A(net217),
    .B(_01783_));
 sg13g2_o21ai_1 _06875_ (.B1(_01784_),
    .Y(_01785_),
    .A1(net217),
    .A2(_01670_));
 sg13g2_a22oi_1 _06876_ (.Y(_01786_),
    .B1(_01785_),
    .B2(_01490_),
    .A2(_01781_),
    .A1(_01507_));
 sg13g2_o21ai_1 _06877_ (.B1(_01786_),
    .Y(_01787_),
    .A1(_01511_),
    .A2(_01777_));
 sg13g2_buf_1 _06878_ (.A(net396),
    .X(_01788_));
 sg13g2_nand2_1 _06879_ (.Y(_01789_),
    .A(net339),
    .B(_00696_));
 sg13g2_o21ai_1 _06880_ (.B1(_01500_),
    .Y(_01790_),
    .A1(_01778_),
    .A2(_01504_));
 sg13g2_nand2b_1 _06881_ (.Y(_01791_),
    .B(_01790_),
    .A_N(_01789_));
 sg13g2_nand3b_1 _06882_ (.B(_01789_),
    .C(net298),
    .Y(_01792_),
    .A_N(_01778_));
 sg13g2_a21oi_1 _06883_ (.A1(_01791_),
    .A2(_01792_),
    .Y(_01793_),
    .B1(net294));
 sg13g2_nor3_1 _06884_ (.A(net218),
    .B(_01787_),
    .C(_01793_),
    .Y(_01794_));
 sg13g2_a21oi_1 _06885_ (.A1(net218),
    .A2(_01766_),
    .Y(_01795_),
    .B1(_01794_));
 sg13g2_inv_1 _06886_ (.Y(_01796_),
    .A(net388));
 sg13g2_nor2_1 _06887_ (.A(net343),
    .B(_01796_),
    .Y(_01797_));
 sg13g2_a21oi_1 _06888_ (.A1(net343),
    .A2(_01795_),
    .Y(_01798_),
    .B1(_01797_));
 sg13g2_nand2_1 _06889_ (.Y(_01799_),
    .A(_01757_),
    .B(_01449_));
 sg13g2_o21ai_1 _06890_ (.B1(_01799_),
    .Y(_01800_),
    .A1(net139),
    .A2(_01798_));
 sg13g2_buf_1 _06891_ (.A(_01800_),
    .X(_01801_));
 sg13g2_inv_1 _06892_ (.Y(_01802_),
    .A(_01801_));
 sg13g2_buf_1 _06893_ (.A(\z80.tv80s.i_tv80_core.ACC[3] ),
    .X(_01803_));
 sg13g2_nand2_1 _06894_ (.Y(_01804_),
    .A(\z80.tv80s.i_tv80_core.Ap[3] ),
    .B(net130));
 sg13g2_o21ai_1 _06895_ (.B1(_01804_),
    .Y(_01805_),
    .A1(net379),
    .A2(_01599_));
 sg13g2_a22oi_1 _06896_ (.Y(_01806_),
    .B1(_01805_),
    .B2(net169),
    .A2(_01597_),
    .A1(net379));
 sg13g2_buf_1 _06897_ (.A(\z80.tv80s.i_tv80_core.I[3] ),
    .X(_01807_));
 sg13g2_mux2_1 _06898_ (.A0(_01807_),
    .A1(\z80.tv80s.i_tv80_core.R[3] ),
    .S(net160),
    .X(_01808_));
 sg13g2_nor2_1 _06899_ (.A(net155),
    .B(_01808_),
    .Y(_01809_));
 sg13g2_a21oi_1 _06900_ (.A1(net152),
    .A2(_01806_),
    .Y(_01810_),
    .B1(_01809_));
 sg13g2_nand2_1 _06901_ (.Y(_01811_),
    .A(_01538_),
    .B(_01810_));
 sg13g2_o21ai_1 _06902_ (.B1(_01811_),
    .Y(_01812_),
    .A1(net161),
    .A2(_01802_));
 sg13g2_nand2_1 _06903_ (.Y(_01813_),
    .A(_00224_),
    .B(net196));
 sg13g2_o21ai_1 _06904_ (.B1(_01813_),
    .Y(_00289_),
    .A1(net181),
    .A2(_01812_));
 sg13g2_and2_1 _06905_ (.A(net383),
    .B(_01758_),
    .X(_01814_));
 sg13g2_nor2_1 _06906_ (.A(net345),
    .B(_01758_),
    .Y(_01815_));
 sg13g2_xnor2_1 _06907_ (.Y(_01816_),
    .A(net383),
    .B(_01757_));
 sg13g2_nor2_1 _06908_ (.A(_01723_),
    .B(_01816_),
    .Y(_01817_));
 sg13g2_a221oi_1 _06909_ (.B2(_01754_),
    .C1(_01817_),
    .B1(_01815_),
    .A1(_01752_),
    .Y(_01818_),
    .A2(_01814_));
 sg13g2_buf_2 _06910_ (.A(_01818_),
    .X(_01819_));
 sg13g2_buf_1 _06911_ (.A(\z80.tv80s.i_tv80_core.BusB[4] ),
    .X(_01820_));
 sg13g2_xnor2_1 _06912_ (.Y(_01821_),
    .A(_01782_),
    .B(net378));
 sg13g2_xnor2_1 _06913_ (.Y(_01822_),
    .A(net298),
    .B(_01821_));
 sg13g2_xnor2_1 _06914_ (.Y(_01823_),
    .A(_01819_),
    .B(_01822_));
 sg13g2_buf_1 _06915_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .X(_01824_));
 sg13g2_buf_1 _06916_ (.A(_01824_),
    .X(_01825_));
 sg13g2_xnor2_1 _06917_ (.Y(_01826_),
    .A(net338),
    .B(net378));
 sg13g2_nand3_1 _06918_ (.B(net338),
    .C(net378),
    .A(net299),
    .Y(_01827_));
 sg13g2_o21ai_1 _06919_ (.B1(_01827_),
    .Y(_01828_),
    .A1(net299),
    .A2(_01826_));
 sg13g2_inv_2 _06920_ (.Y(_01829_),
    .A(_01824_));
 sg13g2_inv_2 _06921_ (.Y(_01830_),
    .A(net378));
 sg13g2_nand2_1 _06922_ (.Y(_01831_),
    .A(_01829_),
    .B(_01830_));
 sg13g2_a22oi_1 _06923_ (.Y(_01832_),
    .B1(_01831_),
    .B2(_01523_),
    .A2(_01828_),
    .A1(net256));
 sg13g2_o21ai_1 _06924_ (.B1(_01832_),
    .Y(_01833_),
    .A1(_01621_),
    .A2(_01823_));
 sg13g2_inv_2 _06925_ (.Y(_01834_),
    .A(_01717_));
 sg13g2_nand3_1 _06926_ (.B(_01653_),
    .C(_01658_),
    .A(net338),
    .Y(_01835_));
 sg13g2_o21ai_1 _06927_ (.B1(_01835_),
    .Y(_01836_),
    .A1(net338),
    .A2(_01658_));
 sg13g2_nand2_1 _06928_ (.Y(_01837_),
    .A(_01655_),
    .B(_01635_));
 sg13g2_o21ai_1 _06929_ (.B1(_01723_),
    .Y(_01838_),
    .A1(net340),
    .A2(_01837_));
 sg13g2_and2_1 _06930_ (.A(_01783_),
    .B(_01838_),
    .X(_01839_));
 sg13g2_nand2_1 _06931_ (.Y(_01840_),
    .A(_01653_),
    .B(_01837_));
 sg13g2_nand2_1 _06932_ (.Y(_01841_),
    .A(_01723_),
    .B(_01782_));
 sg13g2_a21oi_1 _06933_ (.A1(_01658_),
    .A2(_01840_),
    .Y(_01842_),
    .B1(_01841_));
 sg13g2_buf_1 _06934_ (.A(_01717_),
    .X(_01843_));
 sg13g2_o21ai_1 _06935_ (.B1(net337),
    .Y(_01844_),
    .A1(_01839_),
    .A2(_01842_));
 sg13g2_o21ai_1 _06936_ (.B1(_01844_),
    .Y(_01845_),
    .A1(_01782_),
    .A2(_01660_));
 sg13g2_a21oi_2 _06937_ (.B1(_01845_),
    .Y(_01846_),
    .A2(_01836_),
    .A1(_01834_));
 sg13g2_nor3_2 _06938_ (.A(net217),
    .B(net307),
    .C(net339),
    .Y(_01847_));
 sg13g2_nor2_1 _06939_ (.A(_01516_),
    .B(_01847_),
    .Y(_01848_));
 sg13g2_a21oi_1 _06940_ (.A1(_01712_),
    .A2(_01847_),
    .Y(_01849_),
    .B1(_01848_));
 sg13g2_buf_1 _06941_ (.A(_00198_),
    .X(_01850_));
 sg13g2_inv_1 _06942_ (.Y(_01851_),
    .A(net377));
 sg13g2_nor2_1 _06943_ (.A(net308),
    .B(_01851_),
    .Y(_01852_));
 sg13g2_a21oi_1 _06944_ (.A1(net308),
    .A2(_01723_),
    .Y(_01853_),
    .B1(_01852_));
 sg13g2_a221oi_1 _06945_ (.B2(_01490_),
    .C1(net218),
    .B1(_01853_),
    .A1(_01825_),
    .Y(_01854_),
    .A2(_01507_));
 sg13g2_o21ai_1 _06946_ (.B1(_01854_),
    .Y(_01855_),
    .A1(_01499_),
    .A2(_01849_));
 sg13g2_a21oi_1 _06947_ (.A1(_01669_),
    .A2(_01847_),
    .Y(_01856_),
    .B1(_01855_));
 sg13g2_o21ai_1 _06948_ (.B1(_01856_),
    .Y(_01857_),
    .A1(_01511_),
    .A2(_01846_));
 sg13g2_o21ai_1 _06949_ (.B1(_01857_),
    .Y(_01858_),
    .A1(_01618_),
    .A2(_01833_));
 sg13g2_nand2_1 _06950_ (.Y(_01859_),
    .A(net347),
    .B(\z80.tv80s.di_reg[4] ));
 sg13g2_o21ai_1 _06951_ (.B1(_01859_),
    .Y(_01860_),
    .A1(net347),
    .A2(_01858_));
 sg13g2_nand2_1 _06952_ (.Y(_01861_),
    .A(_01830_),
    .B(net139));
 sg13g2_o21ai_1 _06953_ (.B1(_01861_),
    .Y(_01862_),
    .A1(net139),
    .A2(_01860_));
 sg13g2_buf_1 _06954_ (.A(_01862_),
    .X(_01863_));
 sg13g2_buf_2 _06955_ (.A(\z80.tv80s.i_tv80_core.ACC[4] ),
    .X(_01864_));
 sg13g2_nand2_1 _06956_ (.Y(_01865_),
    .A(\z80.tv80s.i_tv80_core.Ap[4] ),
    .B(_01576_));
 sg13g2_o21ai_1 _06957_ (.B1(_01865_),
    .Y(_01866_),
    .A1(_01864_),
    .A2(_01599_));
 sg13g2_a22oi_1 _06958_ (.Y(_01867_),
    .B1(_01866_),
    .B2(net169),
    .A2(_01597_),
    .A1(_01864_));
 sg13g2_buf_1 _06959_ (.A(\z80.tv80s.i_tv80_core.I[4] ),
    .X(_01868_));
 sg13g2_mux2_1 _06960_ (.A0(_01868_),
    .A1(\z80.tv80s.i_tv80_core.R[4] ),
    .S(net160),
    .X(_01869_));
 sg13g2_nor2_1 _06961_ (.A(net155),
    .B(_01869_),
    .Y(_01870_));
 sg13g2_a21oi_1 _06962_ (.A1(_01544_),
    .A2(_01867_),
    .Y(_01871_),
    .B1(_01870_));
 sg13g2_nand2_1 _06963_ (.Y(_01872_),
    .A(_01538_),
    .B(_01871_));
 sg13g2_o21ai_1 _06964_ (.B1(_01872_),
    .Y(_01873_),
    .A1(net161),
    .A2(_01863_));
 sg13g2_nand2_1 _06965_ (.Y(_01874_),
    .A(_00225_),
    .B(net196));
 sg13g2_o21ai_1 _06966_ (.B1(_01874_),
    .Y(_00290_),
    .A1(net181),
    .A2(_01873_));
 sg13g2_buf_1 _06967_ (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .X(_01875_));
 sg13g2_buf_2 _06968_ (.A(\z80.tv80s.i_tv80_core.BusB[5] ),
    .X(_01876_));
 sg13g2_xor2_1 _06969_ (.B(_01876_),
    .A(_01875_),
    .X(_01877_));
 sg13g2_buf_2 _06970_ (.A(_01877_),
    .X(_01878_));
 sg13g2_buf_1 _06971_ (.A(net298),
    .X(_01879_));
 sg13g2_nand2_1 _06972_ (.Y(_01880_),
    .A(_01783_),
    .B(net378));
 sg13g2_nand2b_1 _06973_ (.Y(_01881_),
    .B(_01880_),
    .A_N(_01819_));
 sg13g2_a22oi_1 _06974_ (.Y(_01882_),
    .B1(_01881_),
    .B2(_01829_),
    .A2(_01819_),
    .A1(_01830_));
 sg13g2_nand2_1 _06975_ (.Y(_01883_),
    .A(net338),
    .B(_01830_));
 sg13g2_o21ai_1 _06976_ (.B1(_01883_),
    .Y(_01884_),
    .A1(_01819_),
    .A2(_01880_));
 sg13g2_nor3_1 _06977_ (.A(_01783_),
    .B(net378),
    .C(_01819_),
    .Y(_01885_));
 sg13g2_a21oi_1 _06978_ (.A1(net255),
    .A2(_01884_),
    .Y(_01886_),
    .B1(_01885_));
 sg13g2_o21ai_1 _06979_ (.B1(_01886_),
    .Y(_01887_),
    .A1(net255),
    .A2(_01882_));
 sg13g2_xor2_1 _06980_ (.B(_01887_),
    .A(_01878_),
    .X(_01888_));
 sg13g2_buf_1 _06981_ (.A(_01875_),
    .X(_01889_));
 sg13g2_nand2_1 _06982_ (.Y(_01890_),
    .A(net336),
    .B(_01876_));
 sg13g2_nand2_1 _06983_ (.Y(_01891_),
    .A(net384),
    .B(_01878_));
 sg13g2_o21ai_1 _06984_ (.B1(_01891_),
    .Y(_01892_),
    .A1(net344),
    .A2(_01890_));
 sg13g2_or2_1 _06985_ (.X(_01893_),
    .B(_01876_),
    .A(_01889_));
 sg13g2_a22oi_1 _06986_ (.Y(_01894_),
    .B1(_01893_),
    .B2(_01523_),
    .A2(_01892_),
    .A1(net256));
 sg13g2_o21ai_1 _06987_ (.B1(_01894_),
    .Y(_01895_),
    .A1(_01621_),
    .A2(_01888_));
 sg13g2_buf_1 _06988_ (.A(net217),
    .X(_01896_));
 sg13g2_nand2_1 _06989_ (.Y(_01897_),
    .A(net195),
    .B(net269));
 sg13g2_o21ai_1 _06990_ (.B1(_01500_),
    .Y(_01898_),
    .A1(_01650_),
    .A2(_01504_));
 sg13g2_nand2b_1 _06991_ (.Y(_01899_),
    .B(_01898_),
    .A_N(_01897_));
 sg13g2_nand3b_1 _06992_ (.B(_01897_),
    .C(_01879_),
    .Y(_01900_),
    .A_N(_01650_));
 sg13g2_a21oi_1 _06993_ (.A1(_01899_),
    .A2(_01900_),
    .Y(_01901_),
    .B1(_01749_));
 sg13g2_nor2_1 _06994_ (.A(_01829_),
    .B(_01658_),
    .Y(_01902_));
 sg13g2_buf_2 _06995_ (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .X(_01903_));
 sg13g2_inv_1 _06996_ (.Y(_01904_),
    .A(_01875_));
 sg13g2_nor3_1 _06997_ (.A(_01829_),
    .B(_01904_),
    .C(_01658_),
    .Y(_01905_));
 sg13g2_and2_1 _06998_ (.A(_01903_),
    .B(_01905_),
    .X(_01906_));
 sg13g2_buf_1 _06999_ (.A(_01906_),
    .X(_01907_));
 sg13g2_xor2_1 _07000_ (.B(_01905_),
    .A(_01903_),
    .X(_01908_));
 sg13g2_o21ai_1 _07001_ (.B1(net377),
    .Y(_01909_),
    .A1(_01829_),
    .A2(_01658_));
 sg13g2_nand2_1 _07002_ (.Y(_01910_),
    .A(_01851_),
    .B(_01902_));
 sg13g2_buf_2 _07003_ (.A(_00199_),
    .X(_01911_));
 sg13g2_nor2_1 _07004_ (.A(_01911_),
    .B(_01660_),
    .Y(_01912_));
 sg13g2_a221oi_1 _07005_ (.B2(_01910_),
    .C1(_01912_),
    .B1(_01909_),
    .A1(_01660_),
    .Y(_01913_),
    .A2(_01908_));
 sg13g2_buf_1 _07006_ (.A(\z80.tv80s.i_tv80_core.BusA[7] ),
    .X(_01914_));
 sg13g2_inv_1 _07007_ (.Y(_01915_),
    .A(net376));
 sg13g2_o21ai_1 _07008_ (.B1(_01915_),
    .Y(_01916_),
    .A1(_01494_),
    .A2(_01913_));
 sg13g2_nor2_1 _07009_ (.A(net381),
    .B(_01907_),
    .Y(_01917_));
 sg13g2_and2_1 _07010_ (.A(_01909_),
    .B(_01910_),
    .X(_01918_));
 sg13g2_a21oi_1 _07011_ (.A1(_01660_),
    .A2(_01908_),
    .Y(_01919_),
    .B1(_01912_));
 sg13g2_nand2b_1 _07012_ (.Y(_01920_),
    .B(_01919_),
    .A_N(_01918_));
 sg13g2_buf_1 _07013_ (.A(_01920_),
    .X(_01921_));
 sg13g2_a221oi_1 _07014_ (.B2(_01921_),
    .C1(net391),
    .B1(_01917_),
    .A1(_01907_),
    .Y(_01922_),
    .A2(_01916_));
 sg13g2_buf_1 _07015_ (.A(_01922_),
    .X(_01923_));
 sg13g2_xor2_1 _07016_ (.B(_01923_),
    .A(_01902_),
    .X(_01924_));
 sg13g2_nor2_1 _07017_ (.A(_01903_),
    .B(net336),
    .Y(_01925_));
 sg13g2_o21ai_1 _07018_ (.B1(_01925_),
    .Y(_01926_),
    .A1(_01829_),
    .A2(_01658_));
 sg13g2_a21oi_2 _07019_ (.B1(_01254_),
    .Y(_01927_),
    .A2(_01926_),
    .A1(net376));
 sg13g2_or3_1 _07020_ (.A(_01824_),
    .B(_01656_),
    .C(_01840_),
    .X(_01928_));
 sg13g2_buf_2 _07021_ (.A(_01928_),
    .X(_01929_));
 sg13g2_or2_1 _07022_ (.X(_01930_),
    .B(_01929_),
    .A(_01927_));
 sg13g2_nand2_1 _07023_ (.Y(_01931_),
    .A(_01927_),
    .B(_01929_));
 sg13g2_a21oi_1 _07024_ (.A1(_01930_),
    .A2(_01931_),
    .Y(_01932_),
    .B1(_01834_));
 sg13g2_a21oi_1 _07025_ (.A1(_01834_),
    .A2(_01924_),
    .Y(_01933_),
    .B1(_01932_));
 sg13g2_xnor2_1 _07026_ (.Y(_01934_),
    .A(net377),
    .B(_01933_));
 sg13g2_nand2_1 _07027_ (.Y(_01935_),
    .A(_01486_),
    .B(_01488_));
 sg13g2_nand2_1 _07028_ (.Y(_01936_),
    .A(net195),
    .B(_01911_));
 sg13g2_o21ai_1 _07029_ (.B1(_01936_),
    .Y(_01937_),
    .A1(net195),
    .A2(_01783_));
 sg13g2_nor2_1 _07030_ (.A(_01935_),
    .B(_01937_),
    .Y(_01938_));
 sg13g2_a221oi_1 _07031_ (.B2(_01934_),
    .C1(_01938_),
    .B1(_01662_),
    .A1(net336),
    .Y(_01939_),
    .A2(_01507_));
 sg13g2_nor2b_1 _07032_ (.A(_01901_),
    .B_N(_01939_),
    .Y(_01940_));
 sg13g2_nand2b_1 _07033_ (.Y(_01941_),
    .B(_01512_),
    .A_N(_01449_));
 sg13g2_a21oi_1 _07034_ (.A1(_01618_),
    .A2(_01940_),
    .Y(_01942_),
    .B1(_01941_));
 sg13g2_o21ai_1 _07035_ (.B1(_01942_),
    .Y(_01943_),
    .A1(_01618_),
    .A2(_01895_));
 sg13g2_inv_1 _07036_ (.Y(_01944_),
    .A(net386));
 sg13g2_nor3_1 _07037_ (.A(net343),
    .B(_01944_),
    .C(net139),
    .Y(_01945_));
 sg13g2_a21oi_2 _07038_ (.B1(_01945_),
    .Y(_01946_),
    .A2(net139),
    .A1(_01876_));
 sg13g2_nand2_2 _07039_ (.Y(_01947_),
    .A(_01943_),
    .B(_01946_));
 sg13g2_buf_1 _07040_ (.A(\z80.tv80s.i_tv80_core.ACC[5] ),
    .X(_01948_));
 sg13g2_nand2_1 _07041_ (.Y(_01949_),
    .A(\z80.tv80s.i_tv80_core.Ap[5] ),
    .B(net129));
 sg13g2_o21ai_1 _07042_ (.B1(_01949_),
    .Y(_01950_),
    .A1(net375),
    .A2(_01599_));
 sg13g2_buf_1 _07043_ (.A(_01595_),
    .X(_01951_));
 sg13g2_a22oi_1 _07044_ (.Y(_01952_),
    .B1(_01950_),
    .B2(net168),
    .A2(_01597_),
    .A1(net375));
 sg13g2_buf_1 _07045_ (.A(\z80.tv80s.i_tv80_core.I[5] ),
    .X(_01953_));
 sg13g2_buf_1 _07046_ (.A(\z80.tv80s.i_tv80_core.R[5] ),
    .X(_01954_));
 sg13g2_mux2_1 _07047_ (.A0(_01953_),
    .A1(_01954_),
    .S(net160),
    .X(_01955_));
 sg13g2_nor2_1 _07048_ (.A(net152),
    .B(_01955_),
    .Y(_01956_));
 sg13g2_a21oi_1 _07049_ (.A1(net152),
    .A2(_01952_),
    .Y(_01957_),
    .B1(_01956_));
 sg13g2_mux2_1 _07050_ (.A0(_01947_),
    .A1(_01957_),
    .S(net161),
    .X(_01958_));
 sg13g2_nand2_1 _07051_ (.Y(_01959_),
    .A(_00226_),
    .B(net196));
 sg13g2_o21ai_1 _07052_ (.B1(_01959_),
    .Y(_00291_),
    .A1(net181),
    .A2(_01958_));
 sg13g2_buf_1 _07053_ (.A(net202),
    .X(_01960_));
 sg13g2_buf_1 _07054_ (.A(\z80.tv80s.i_tv80_core.BusB[6] ),
    .X(_01961_));
 sg13g2_inv_1 _07055_ (.Y(_01962_),
    .A(net374));
 sg13g2_nor3_1 _07056_ (.A(net297),
    .B(_01821_),
    .C(_01878_),
    .Y(_01963_));
 sg13g2_nand3_1 _07057_ (.B(_01821_),
    .C(_01878_),
    .A(net297),
    .Y(_01964_));
 sg13g2_nand2b_1 _07058_ (.Y(_01965_),
    .B(_01964_),
    .A_N(_01963_));
 sg13g2_inv_1 _07059_ (.Y(_01966_),
    .A(_01965_));
 sg13g2_nand2_1 _07060_ (.Y(_01967_),
    .A(net345),
    .B(_01830_));
 sg13g2_nand3_1 _07061_ (.B(_01820_),
    .C(_01878_),
    .A(_01502_),
    .Y(_01968_));
 sg13g2_o21ai_1 _07062_ (.B1(_01968_),
    .Y(_01969_),
    .A1(_01878_),
    .A2(_01967_));
 sg13g2_xor2_1 _07063_ (.B(_01876_),
    .A(net345),
    .X(_01970_));
 sg13g2_a22oi_1 _07064_ (.Y(_01971_),
    .B1(_01970_),
    .B2(_01851_),
    .A2(_01969_),
    .A1(net338));
 sg13g2_o21ai_1 _07065_ (.B1(_01971_),
    .Y(_01972_),
    .A1(_01819_),
    .A2(_01966_));
 sg13g2_buf_1 _07066_ (.A(_01972_),
    .X(_01973_));
 sg13g2_xor2_1 _07067_ (.B(net374),
    .A(_01903_),
    .X(_01974_));
 sg13g2_xnor2_1 _07068_ (.Y(_01975_),
    .A(net297),
    .B(_01974_));
 sg13g2_xnor2_1 _07069_ (.Y(_01976_),
    .A(net149),
    .B(_01975_));
 sg13g2_and2_1 _07070_ (.A(_01903_),
    .B(net374),
    .X(_01977_));
 sg13g2_mux2_1 _07071_ (.A0(_01974_),
    .A1(_01977_),
    .S(net299),
    .X(_01978_));
 sg13g2_or2_1 _07072_ (.X(_01979_),
    .B(\z80.tv80s.i_tv80_core.BusB[6] ),
    .A(_01903_));
 sg13g2_a22oi_1 _07073_ (.Y(_01980_),
    .B1(_01979_),
    .B2(_01523_),
    .A2(_01978_),
    .A1(net256));
 sg13g2_o21ai_1 _07074_ (.B1(_01980_),
    .Y(_01981_),
    .A1(_01621_),
    .A2(_01976_));
 sg13g2_nor2_1 _07075_ (.A(_01918_),
    .B(_01923_),
    .Y(_01982_));
 sg13g2_xnor2_1 _07076_ (.Y(_01983_),
    .A(_01919_),
    .B(_01982_));
 sg13g2_o21ai_1 _07077_ (.B1(_01931_),
    .Y(_01984_),
    .A1(_01904_),
    .A2(_01929_));
 sg13g2_nand2_1 _07078_ (.Y(_01985_),
    .A(net377),
    .B(net336));
 sg13g2_mux2_1 _07079_ (.A0(_01985_),
    .A1(net336),
    .S(_01927_),
    .X(_01986_));
 sg13g2_or2_1 _07080_ (.X(_01987_),
    .B(_01986_),
    .A(_01929_));
 sg13g2_o21ai_1 _07081_ (.B1(_01987_),
    .Y(_01988_),
    .A1(net377),
    .A2(_01984_));
 sg13g2_xor2_1 _07082_ (.B(_01988_),
    .A(_01911_),
    .X(_01989_));
 sg13g2_nand2_1 _07083_ (.Y(_01990_),
    .A(net337),
    .B(_01989_));
 sg13g2_o21ai_1 _07084_ (.B1(_01990_),
    .Y(_01991_),
    .A1(net337),
    .A2(_01983_));
 sg13g2_nor2_1 _07085_ (.A(net184),
    .B(_01516_),
    .Y(_01992_));
 sg13g2_a21oi_1 _07086_ (.A1(net184),
    .A2(_01712_),
    .Y(_01993_),
    .B1(_01992_));
 sg13g2_buf_1 _07087_ (.A(_01903_),
    .X(_01994_));
 sg13g2_nor2_1 _07088_ (.A(net308),
    .B(_01494_),
    .Y(_01995_));
 sg13g2_a21oi_1 _07089_ (.A1(net262),
    .A2(_01850_),
    .Y(_01996_),
    .B1(_01995_));
 sg13g2_a221oi_1 _07090_ (.B2(_01490_),
    .C1(_01461_),
    .B1(_01996_),
    .A1(_01994_),
    .Y(_01997_),
    .A2(_01507_));
 sg13g2_o21ai_1 _07091_ (.B1(_01997_),
    .Y(_01998_),
    .A1(_00206_),
    .A2(_01993_));
 sg13g2_a21oi_1 _07092_ (.A1(net184),
    .A2(_01669_),
    .Y(_01999_),
    .B1(_01998_));
 sg13g2_o21ai_1 _07093_ (.B1(_01999_),
    .Y(_02000_),
    .A1(_01511_),
    .A2(_01991_));
 sg13g2_o21ai_1 _07094_ (.B1(_02000_),
    .Y(_02001_),
    .A1(_01618_),
    .A2(_01981_));
 sg13g2_nand2_1 _07095_ (.Y(_02002_),
    .A(net347),
    .B(net385));
 sg13g2_o21ai_1 _07096_ (.B1(_02002_),
    .Y(_02003_),
    .A1(net347),
    .A2(_02001_));
 sg13g2_nor2_1 _07097_ (.A(_01695_),
    .B(_02003_),
    .Y(_02004_));
 sg13g2_a21oi_1 _07098_ (.A1(_01962_),
    .A2(_01695_),
    .Y(_02005_),
    .B1(_02004_));
 sg13g2_buf_2 _07099_ (.A(_02005_),
    .X(_02006_));
 sg13g2_buf_2 _07100_ (.A(\z80.tv80s.i_tv80_core.ACC[6] ),
    .X(_02007_));
 sg13g2_nand2_1 _07101_ (.Y(_02008_),
    .A(\z80.tv80s.i_tv80_core.Ap[6] ),
    .B(net129));
 sg13g2_o21ai_1 _07102_ (.B1(_02008_),
    .Y(_02009_),
    .A1(_02007_),
    .A2(_01599_));
 sg13g2_a22oi_1 _07103_ (.Y(_02010_),
    .B1(_02009_),
    .B2(net168),
    .A2(_01597_),
    .A1(_02007_));
 sg13g2_buf_1 _07104_ (.A(\z80.tv80s.i_tv80_core.I[6] ),
    .X(_02011_));
 sg13g2_mux2_1 _07105_ (.A0(_02011_),
    .A1(\z80.tv80s.i_tv80_core.R[6] ),
    .S(net160),
    .X(_02012_));
 sg13g2_nor2_1 _07106_ (.A(net152),
    .B(_02012_),
    .Y(_02013_));
 sg13g2_a21oi_1 _07107_ (.A1(net152),
    .A2(_02010_),
    .Y(_02014_),
    .B1(_02013_));
 sg13g2_mux2_1 _07108_ (.A0(_02006_),
    .A1(_02014_),
    .S(net161),
    .X(_02015_));
 sg13g2_nand2_1 _07109_ (.Y(_02016_),
    .A(_00227_),
    .B(net196));
 sg13g2_o21ai_1 _07110_ (.B1(_02016_),
    .Y(_00292_),
    .A1(net177),
    .A2(_02015_));
 sg13g2_buf_1 _07111_ (.A(\z80.tv80s.i_tv80_core.BusB[7] ),
    .X(_02017_));
 sg13g2_buf_1 _07112_ (.A(_02017_),
    .X(_02018_));
 sg13g2_inv_1 _07113_ (.Y(_02019_),
    .A(_01400_));
 sg13g2_nor3_1 _07114_ (.A(_01903_),
    .B(net336),
    .C(_01929_),
    .Y(_02020_));
 sg13g2_xnor2_1 _07115_ (.Y(_02021_),
    .A(_01493_),
    .B(_02020_));
 sg13g2_xnor2_1 _07116_ (.Y(_02022_),
    .A(_01911_),
    .B(net336));
 sg13g2_nor2_1 _07117_ (.A(_01929_),
    .B(_02022_),
    .Y(_02023_));
 sg13g2_nor2_1 _07118_ (.A(net377),
    .B(_01911_),
    .Y(_02024_));
 sg13g2_a22oi_1 _07119_ (.Y(_02025_),
    .B1(_02024_),
    .B2(_01929_),
    .A2(_02023_),
    .A1(net377));
 sg13g2_nor2b_1 _07120_ (.A(_01927_),
    .B_N(_02025_),
    .Y(_02026_));
 sg13g2_xnor2_1 _07121_ (.Y(_02027_),
    .A(_02021_),
    .B(_02026_));
 sg13g2_xnor2_1 _07122_ (.Y(_02028_),
    .A(_01494_),
    .B(_01907_));
 sg13g2_nand2_1 _07123_ (.Y(_02029_),
    .A(_01921_),
    .B(_02028_));
 sg13g2_nor2_1 _07124_ (.A(_01923_),
    .B(_02029_),
    .Y(_02030_));
 sg13g2_nor2_1 _07125_ (.A(_01921_),
    .B(_02028_),
    .Y(_02031_));
 sg13g2_nor3_1 _07126_ (.A(_01717_),
    .B(_02030_),
    .C(_02031_),
    .Y(_02032_));
 sg13g2_a21o_1 _07127_ (.A2(_02027_),
    .A1(net337),
    .B1(_02032_),
    .X(_02033_));
 sg13g2_buf_1 _07128_ (.A(_02033_),
    .X(_02034_));
 sg13g2_nor2_1 _07129_ (.A(net261),
    .B(net339),
    .Y(_02035_));
 sg13g2_a22oi_1 _07130_ (.Y(_02036_),
    .B1(_02035_),
    .B2(net217),
    .A2(_01406_),
    .A1(net339));
 sg13g2_nor2_1 _07131_ (.A(_01779_),
    .B(_02036_),
    .Y(_02037_));
 sg13g2_a22oi_1 _07132_ (.Y(_02038_),
    .B1(_01712_),
    .B2(_02037_),
    .A2(_01507_),
    .A1(net376));
 sg13g2_o21ai_1 _07133_ (.B1(_02038_),
    .Y(_02039_),
    .A1(_01511_),
    .A2(_02034_));
 sg13g2_nand3_1 _07134_ (.B(_00688_),
    .C(_01254_),
    .A(net307),
    .Y(_02040_));
 sg13g2_o21ai_1 _07135_ (.B1(_02040_),
    .Y(_02041_),
    .A1(_00931_),
    .A2(_01477_));
 sg13g2_a22oi_1 _07136_ (.Y(_02042_),
    .B1(_02041_),
    .B2(net259),
    .A2(net269),
    .A1(_01494_));
 sg13g2_nand2_1 _07137_ (.Y(_02043_),
    .A(net195),
    .B(_02042_));
 sg13g2_o21ai_1 _07138_ (.B1(_02043_),
    .Y(_02044_),
    .A1(net195),
    .A2(net335));
 sg13g2_nor2_1 _07139_ (.A(_01935_),
    .B(_02044_),
    .Y(_02045_));
 sg13g2_nand2_1 _07140_ (.Y(_02046_),
    .A(net257),
    .B(_01779_));
 sg13g2_nand4_1 _07141_ (.B(net261),
    .C(net339),
    .A(net271),
    .Y(_02047_),
    .D(net296));
 sg13g2_buf_1 _07142_ (.A(_01896_),
    .X(_02048_));
 sg13g2_a21oi_1 _07143_ (.A1(_02046_),
    .A2(_02047_),
    .Y(_02049_),
    .B1(net176));
 sg13g2_nor2_1 _07144_ (.A(_01788_),
    .B(net296),
    .Y(_02050_));
 sg13g2_o21ai_1 _07145_ (.B1(_01779_),
    .Y(_02051_),
    .A1(net259),
    .A2(_00721_));
 sg13g2_nor2_1 _07146_ (.A(_01779_),
    .B(_02035_),
    .Y(_02052_));
 sg13g2_a221oi_1 _07147_ (.B2(net262),
    .C1(_02052_),
    .B1(_02051_),
    .A1(_00696_),
    .Y(_02053_),
    .A2(_02050_));
 sg13g2_nor3_1 _07148_ (.A(_01516_),
    .B(_02049_),
    .C(_02053_),
    .Y(_02054_));
 sg13g2_nor4_1 _07149_ (.A(_01451_),
    .B(_02039_),
    .C(_02045_),
    .D(_02054_),
    .Y(_02055_));
 sg13g2_nand2b_1 _07150_ (.Y(_02056_),
    .B(net374),
    .A_N(net335));
 sg13g2_a21o_1 _07151_ (.A2(_01962_),
    .A1(net335),
    .B1(net297),
    .X(_02057_));
 sg13g2_a21o_1 _07152_ (.A2(_02056_),
    .A1(net149),
    .B1(_02057_),
    .X(_02058_));
 sg13g2_and2_1 _07153_ (.A(net297),
    .B(_01979_),
    .X(_02059_));
 sg13g2_o21ai_1 _07154_ (.B1(_02059_),
    .Y(_02060_),
    .A1(_01973_),
    .A2(_01977_));
 sg13g2_nor2b_1 _07155_ (.A(net381),
    .B_N(net334),
    .Y(_02061_));
 sg13g2_nor2_1 _07156_ (.A(_01494_),
    .B(net334),
    .Y(_02062_));
 sg13g2_nor2_1 _07157_ (.A(_02061_),
    .B(_02062_),
    .Y(_02063_));
 sg13g2_a221oi_1 _07158_ (.B2(_02060_),
    .C1(_02063_),
    .B1(_02058_),
    .A1(net294),
    .Y(_02064_),
    .A2(_01619_));
 sg13g2_nand4_1 _07159_ (.B(_02058_),
    .C(_02060_),
    .A(_01750_),
    .Y(_02065_),
    .D(_02063_));
 sg13g2_xnor2_1 _07160_ (.Y(_02066_),
    .A(net376),
    .B(_02017_));
 sg13g2_nand3_1 _07161_ (.B(net376),
    .C(_02017_),
    .A(_01475_),
    .Y(_02067_));
 sg13g2_o21ai_1 _07162_ (.B1(_02067_),
    .Y(_02068_),
    .A1(_01475_),
    .A2(_02066_));
 sg13g2_or2_1 _07163_ (.X(_02069_),
    .B(net334),
    .A(net376));
 sg13g2_a22oi_1 _07164_ (.Y(_02070_),
    .B1(_02069_),
    .B2(_01523_),
    .A2(_02068_),
    .A1(net256));
 sg13g2_nand3b_1 _07165_ (.B(_02065_),
    .C(_02070_),
    .Y(_02071_),
    .A_N(_02064_));
 sg13g2_nand2_1 _07166_ (.Y(_02072_),
    .A(net218),
    .B(_02071_));
 sg13g2_a221oi_1 _07167_ (.B2(_02072_),
    .C1(net139),
    .B1(_02055_),
    .A1(net347),
    .Y(_02073_),
    .A2(_02019_));
 sg13g2_a21oi_1 _07168_ (.A1(net334),
    .A2(net139),
    .Y(_02074_),
    .B1(_02073_));
 sg13g2_buf_2 _07169_ (.A(_02074_),
    .X(_02075_));
 sg13g2_buf_2 _07170_ (.A(\z80.tv80s.i_tv80_core.ACC[7] ),
    .X(_02076_));
 sg13g2_nand2_1 _07171_ (.Y(_02077_),
    .A(\z80.tv80s.i_tv80_core.Ap[7] ),
    .B(_01576_));
 sg13g2_o21ai_1 _07172_ (.B1(_02077_),
    .Y(_02078_),
    .A1(_02076_),
    .A2(_01599_));
 sg13g2_a22oi_1 _07173_ (.Y(_02079_),
    .B1(_02078_),
    .B2(net169),
    .A2(_01597_),
    .A1(_02076_));
 sg13g2_buf_2 _07174_ (.A(\z80.tv80s.i_tv80_core.I[7] ),
    .X(_02080_));
 sg13g2_mux2_1 _07175_ (.A0(_02080_),
    .A1(\z80.tv80s.i_tv80_core.R[7] ),
    .S(net160),
    .X(_02081_));
 sg13g2_nor2_1 _07176_ (.A(net155),
    .B(_02081_),
    .Y(_02082_));
 sg13g2_a21oi_1 _07177_ (.A1(_01544_),
    .A2(_02079_),
    .Y(_02083_),
    .B1(_02082_));
 sg13g2_nand2_1 _07178_ (.Y(_02084_),
    .A(_01538_),
    .B(_02083_));
 sg13g2_o21ai_1 _07179_ (.B1(_02084_),
    .Y(_02085_),
    .A1(net161),
    .A2(_02075_));
 sg13g2_nand2_1 _07180_ (.Y(_02086_),
    .A(_00228_),
    .B(net196));
 sg13g2_o21ai_1 _07181_ (.B1(_02086_),
    .Y(_00293_),
    .A1(net177),
    .A2(_02085_));
 sg13g2_buf_1 _07182_ (.A(net226),
    .X(_02087_));
 sg13g2_buf_1 _07183_ (.A(_00995_),
    .X(_02088_));
 sg13g2_buf_1 _07184_ (.A(net115),
    .X(_02089_));
 sg13g2_nand2_2 _07185_ (.Y(_02090_),
    .A(net281),
    .B(net183));
 sg13g2_nor3_1 _07186_ (.A(net280),
    .B(net236),
    .C(_01059_),
    .Y(_02091_));
 sg13g2_buf_1 _07187_ (.A(_00033_),
    .X(_02092_));
 sg13g2_nand2_1 _07188_ (.Y(_02093_),
    .A(net235),
    .B(_02092_));
 sg13g2_a21oi_1 _07189_ (.A1(_02091_),
    .A2(_02093_),
    .Y(_02094_),
    .B1(net170));
 sg13g2_o21ai_1 _07190_ (.B1(_02094_),
    .Y(_02095_),
    .A1(net180),
    .A2(_02090_));
 sg13g2_o21ai_1 _07191_ (.B1(net262),
    .Y(_02096_),
    .A1(net277),
    .A2(_02094_));
 sg13g2_nand3_1 _07192_ (.B(net231),
    .C(_00973_),
    .A(net206),
    .Y(_02097_));
 sg13g2_nor2_1 _07193_ (.A(net308),
    .B(net360),
    .Y(_02098_));
 sg13g2_nor2_1 _07194_ (.A(net180),
    .B(_02098_),
    .Y(_02099_));
 sg13g2_a22oi_1 _07195_ (.Y(_02100_),
    .B1(_02097_),
    .B2(_02099_),
    .A2(_02092_),
    .A1(net180));
 sg13g2_buf_1 _07196_ (.A(net176),
    .X(_02101_));
 sg13g2_nor2_1 _07197_ (.A(net167),
    .B(_00981_),
    .Y(_02102_));
 sg13g2_nor3_1 _07198_ (.A(_00875_),
    .B(_00986_),
    .C(_00678_),
    .Y(_02103_));
 sg13g2_buf_1 _07199_ (.A(_02103_),
    .X(_02104_));
 sg13g2_nor4_2 _07200_ (.A(_00885_),
    .B(net183),
    .C(net170),
    .Y(_02105_),
    .D(_02104_));
 sg13g2_a21oi_1 _07201_ (.A1(net206),
    .A2(_02102_),
    .Y(_02106_),
    .B1(_02105_));
 sg13g2_o21ai_1 _07202_ (.B1(net224),
    .Y(_02107_),
    .A1(_02092_),
    .A2(_02106_));
 sg13g2_a221oi_1 _07203_ (.B2(_01191_),
    .C1(_02107_),
    .B1(_02100_),
    .A1(_02095_),
    .Y(_02108_),
    .A2(_02096_));
 sg13g2_nand2_1 _07204_ (.Y(_02109_),
    .A(net300),
    .B(net260));
 sg13g2_nor2_1 _07205_ (.A(_00779_),
    .B(_00735_),
    .Y(_02110_));
 sg13g2_nand2_1 _07206_ (.Y(_02111_),
    .A(_01057_),
    .B(_02110_));
 sg13g2_nor2_1 _07207_ (.A(_00749_),
    .B(net315),
    .Y(_02112_));
 sg13g2_nor2b_1 _07208_ (.A(net281),
    .B_N(net323),
    .Y(_02113_));
 sg13g2_mux2_1 _07209_ (.A0(_00764_),
    .A1(_02113_),
    .S(_00683_),
    .X(_02114_));
 sg13g2_nand3_1 _07210_ (.B(_02112_),
    .C(_02114_),
    .A(_00649_),
    .Y(_02115_));
 sg13g2_nand3_1 _07211_ (.B(_01413_),
    .C(_02115_),
    .A(_00955_),
    .Y(_02116_));
 sg13g2_nand2_1 _07212_ (.Y(_02117_),
    .A(net269),
    .B(_00842_));
 sg13g2_o21ai_1 _07213_ (.B1(_00920_),
    .Y(_02118_),
    .A1(_02117_),
    .A2(_01059_));
 sg13g2_or3_1 _07214_ (.A(_02111_),
    .B(_02116_),
    .C(_02118_),
    .X(_02119_));
 sg13g2_nor3_2 _07215_ (.A(_01579_),
    .B(_01584_),
    .C(_02119_),
    .Y(_02120_));
 sg13g2_nand2_1 _07216_ (.Y(_02121_),
    .A(net262),
    .B(_01077_));
 sg13g2_a21oi_2 _07217_ (.B1(net240),
    .Y(_02122_),
    .A2(_02121_),
    .A1(net279));
 sg13g2_nor3_1 _07218_ (.A(_00712_),
    .B(_00959_),
    .C(_02122_),
    .Y(_02123_));
 sg13g2_nand2b_1 _07219_ (.Y(_02124_),
    .B(_02123_),
    .A_N(_01096_));
 sg13g2_a21oi_1 _07220_ (.A1(_02120_),
    .A2(_02124_),
    .Y(_02125_),
    .B1(_02092_));
 sg13g2_a21oi_1 _07221_ (.A1(net306),
    .A2(net209),
    .Y(_02126_),
    .B1(_01260_));
 sg13g2_nand2b_1 _07222_ (.Y(_02127_),
    .B(_02126_),
    .A_N(_02125_));
 sg13g2_buf_1 _07223_ (.A(net258),
    .X(_02128_));
 sg13g2_nand2_1 _07224_ (.Y(_02129_),
    .A(net236),
    .B(_00894_));
 sg13g2_and3_1 _07225_ (.X(_02130_),
    .A(net201),
    .B(net267),
    .C(_02129_));
 sg13g2_a21oi_1 _07226_ (.A1(_02101_),
    .A2(net215),
    .Y(_02131_),
    .B1(_02130_));
 sg13g2_nand2_1 _07227_ (.Y(_02132_),
    .A(_02092_),
    .B(_01105_));
 sg13g2_buf_1 _07228_ (.A(_01066_),
    .X(_02133_));
 sg13g2_nand3_1 _07229_ (.B(net175),
    .C(_02129_),
    .A(net235),
    .Y(_02134_));
 sg13g2_nand3b_1 _07230_ (.B(_02134_),
    .C(_01104_),
    .Y(_02135_),
    .A_N(_02098_));
 sg13g2_nand3_1 _07231_ (.B(_02132_),
    .C(_02135_),
    .A(net171),
    .Y(_02136_));
 sg13g2_o21ai_1 _07232_ (.B1(_02136_),
    .Y(_02137_),
    .A1(net171),
    .A2(_02131_));
 sg13g2_inv_1 _07233_ (.Y(_02138_),
    .A(_00034_));
 sg13g2_a22oi_1 _07234_ (.Y(_02139_),
    .B1(_02137_),
    .B2(_02138_),
    .A2(_02127_),
    .A1(_02109_));
 sg13g2_nor2_1 _07235_ (.A(_02108_),
    .B(_02139_),
    .Y(_02140_));
 sg13g2_nand3_1 _07236_ (.B(_01346_),
    .C(_02140_),
    .A(net100),
    .Y(_02141_));
 sg13g2_o21ai_1 _07237_ (.B1(_02141_),
    .Y(_00294_),
    .A1(net299),
    .A2(net194));
 sg13g2_nand2_2 _07238_ (.Y(_02142_),
    .A(_02088_),
    .B(_01346_));
 sg13g2_nand2_1 _07239_ (.Y(_02143_),
    .A(net195),
    .B(net261));
 sg13g2_buf_1 _07240_ (.A(net282),
    .X(_02144_));
 sg13g2_a21oi_1 _07241_ (.A1(_02143_),
    .A2(_00933_),
    .Y(_02145_),
    .B1(net214));
 sg13g2_a221oi_1 _07242_ (.B2(_02112_),
    .C1(_02145_),
    .B1(_02143_),
    .A1(net176),
    .Y(_02146_),
    .A2(net269));
 sg13g2_nor2b_1 _07243_ (.A(_02146_),
    .B_N(_00764_),
    .Y(_02147_));
 sg13g2_nand3b_1 _07244_ (.B(_01327_),
    .C(net257),
    .Y(_02148_),
    .A_N(_01560_));
 sg13g2_nand2_1 _07245_ (.Y(_02149_),
    .A(net214),
    .B(net223));
 sg13g2_nand3_1 _07246_ (.B(_00683_),
    .C(_02149_),
    .A(_01123_),
    .Y(_02150_));
 sg13g2_a21oi_1 _07247_ (.A1(_02148_),
    .A2(_02150_),
    .Y(_02151_),
    .B1(net237));
 sg13g2_o21ai_1 _07248_ (.B1(net203),
    .Y(_02152_),
    .A1(_02147_),
    .A2(_02151_));
 sg13g2_nor2_1 _07249_ (.A(net237),
    .B(_01412_),
    .Y(_02153_));
 sg13g2_nor2_1 _07250_ (.A(net176),
    .B(_01349_),
    .Y(_02154_));
 sg13g2_a21oi_1 _07251_ (.A1(net176),
    .A2(_01078_),
    .Y(_02155_),
    .B1(_02154_));
 sg13g2_nand2_1 _07252_ (.Y(_02156_),
    .A(_01252_),
    .B(_01069_));
 sg13g2_o21ai_1 _07253_ (.B1(_02156_),
    .Y(_02157_),
    .A1(net214),
    .A2(_02155_));
 sg13g2_o21ai_1 _07254_ (.B1(_02157_),
    .Y(_02158_),
    .A1(_01044_),
    .A2(_02153_));
 sg13g2_nand2_1 _07255_ (.Y(_02159_),
    .A(net243),
    .B(_00811_));
 sg13g2_a22oi_1 _07256_ (.Y(_02160_),
    .B1(_01375_),
    .B2(_00742_),
    .A2(_01026_),
    .A1(_00752_));
 sg13g2_nand2b_1 _07257_ (.Y(_02161_),
    .B(_00814_),
    .A_N(_02160_));
 sg13g2_a21oi_2 _07258_ (.B1(net234),
    .Y(_02162_),
    .A2(_02161_),
    .A1(_02159_));
 sg13g2_a21oi_1 _07259_ (.A1(_00749_),
    .A2(_01359_),
    .Y(_02163_),
    .B1(_01078_));
 sg13g2_nor3_1 _07260_ (.A(_02048_),
    .B(_00717_),
    .C(_02163_),
    .Y(_02164_));
 sg13g2_a22oi_1 _07261_ (.Y(_02165_),
    .B1(_01078_),
    .B2(_02144_),
    .A2(_01359_),
    .A1(_02048_));
 sg13g2_nor2b_1 _07262_ (.A(_02165_),
    .B_N(_00764_),
    .Y(_02166_));
 sg13g2_nor2_1 _07263_ (.A(_00671_),
    .B(net284),
    .Y(_02167_));
 sg13g2_a22oi_1 _07264_ (.Y(_02168_),
    .B1(_02167_),
    .B2(_01359_),
    .A2(_01151_),
    .A1(_00914_));
 sg13g2_o21ai_1 _07265_ (.B1(_02168_),
    .Y(_02169_),
    .A1(net175),
    .A2(_00894_));
 sg13g2_nor4_1 _07266_ (.A(_02162_),
    .B(_02164_),
    .C(_02166_),
    .D(_02169_),
    .Y(_02170_));
 sg13g2_nand3_1 _07267_ (.B(_02158_),
    .C(_02170_),
    .A(_02152_),
    .Y(_02171_));
 sg13g2_nand2_1 _07268_ (.Y(_02172_),
    .A(_00672_),
    .B(_01359_));
 sg13g2_o21ai_1 _07269_ (.B1(_02172_),
    .Y(_02173_),
    .A1(net240),
    .A2(_00734_));
 sg13g2_nand3_1 _07270_ (.B(_02110_),
    .C(_01444_),
    .A(net201),
    .Y(_02174_));
 sg13g2_or4_1 _07271_ (.A(_01547_),
    .B(_02171_),
    .C(_02173_),
    .D(_02174_),
    .X(_02175_));
 sg13g2_o21ai_1 _07272_ (.B1(_02175_),
    .Y(_02176_),
    .A1(net220),
    .A2(net180));
 sg13g2_buf_2 _07273_ (.A(_00029_),
    .X(_02177_));
 sg13g2_nand2_1 _07274_ (.Y(_02178_),
    .A(_02177_),
    .B(_01105_));
 sg13g2_nand2_1 _07275_ (.Y(_02179_),
    .A(net220),
    .B(net306));
 sg13g2_nand3_1 _07276_ (.B(net235),
    .C(net175),
    .A(net310),
    .Y(_02180_));
 sg13g2_nand3_1 _07277_ (.B(_02179_),
    .C(_02180_),
    .A(_01104_),
    .Y(_02181_));
 sg13g2_nand3_1 _07278_ (.B(_02178_),
    .C(_02181_),
    .A(net171),
    .Y(_02182_));
 sg13g2_o21ai_1 _07279_ (.B1(_02182_),
    .Y(_02183_),
    .A1(net171),
    .A2(_02176_));
 sg13g2_nand2_1 _07280_ (.Y(_02184_),
    .A(net220),
    .B(_01115_));
 sg13g2_o21ai_1 _07281_ (.B1(_02184_),
    .Y(_02185_),
    .A1(net215),
    .A2(_02177_));
 sg13g2_nand3_1 _07282_ (.B(_02123_),
    .C(_02185_),
    .A(net184),
    .Y(_02186_));
 sg13g2_nor2_1 _07283_ (.A(net232),
    .B(_00784_),
    .Y(_02187_));
 sg13g2_nor2b_1 _07284_ (.A(_02187_),
    .B_N(_02120_),
    .Y(_02188_));
 sg13g2_mux2_1 _07285_ (.A0(_02177_),
    .A1(_02186_),
    .S(_02188_),
    .X(_02189_));
 sg13g2_nor2_1 _07286_ (.A(_00845_),
    .B(net219),
    .Y(_02190_));
 sg13g2_a221oi_1 _07287_ (.B2(net220),
    .C1(_00959_),
    .B1(_02190_),
    .A1(_01096_),
    .Y(_02191_),
    .A2(_02187_));
 sg13g2_nand3_1 _07288_ (.B(_02189_),
    .C(_02191_),
    .A(net265),
    .Y(_02192_));
 sg13g2_a22oi_1 _07289_ (.Y(_02193_),
    .B1(_02192_),
    .B2(_02109_),
    .A2(_02183_),
    .A1(_02138_));
 sg13g2_nand2_1 _07290_ (.Y(_02194_),
    .A(net206),
    .B(_02177_));
 sg13g2_a22oi_1 _07291_ (.Y(_02195_),
    .B1(_02102_),
    .B2(_02194_),
    .A2(_01185_),
    .A1(net204));
 sg13g2_nand4_1 _07292_ (.B(net204),
    .C(net277),
    .A(_01332_),
    .Y(_02196_),
    .D(_01554_));
 sg13g2_o21ai_1 _07293_ (.B1(_02196_),
    .Y(_02197_),
    .A1(net277),
    .A2(_02195_));
 sg13g2_a21oi_1 _07294_ (.A1(_01332_),
    .A2(net306),
    .Y(_02198_),
    .B1(net180));
 sg13g2_a22oi_1 _07295_ (.Y(_02199_),
    .B1(_02097_),
    .B2(_02198_),
    .A2(_02177_),
    .A1(net180));
 sg13g2_and2_1 _07296_ (.A(_01191_),
    .B(_02199_),
    .X(_02200_));
 sg13g2_a21oi_1 _07297_ (.A1(net206),
    .A2(_02091_),
    .Y(_02201_),
    .B1(_02105_));
 sg13g2_nor2_1 _07298_ (.A(_00874_),
    .B(_02104_),
    .Y(_02202_));
 sg13g2_o21ai_1 _07299_ (.B1(_02202_),
    .Y(_02203_),
    .A1(_02177_),
    .A2(_02201_));
 sg13g2_buf_1 _07300_ (.A(_01286_),
    .X(_02204_));
 sg13g2_nand2_1 _07301_ (.Y(_02205_),
    .A(_02204_),
    .B(_01120_));
 sg13g2_a22oi_1 _07302_ (.Y(_02206_),
    .B1(_02205_),
    .B2(net261),
    .A2(_02195_),
    .A1(_02090_));
 sg13g2_nor4_1 _07303_ (.A(_02197_),
    .B(_02200_),
    .C(_02203_),
    .D(_02206_),
    .Y(_02207_));
 sg13g2_or3_1 _07304_ (.A(_02142_),
    .B(_02193_),
    .C(_02207_),
    .X(_02208_));
 sg13g2_o21ai_1 _07305_ (.B1(_02208_),
    .Y(_00295_),
    .A1(net297),
    .A2(net194));
 sg13g2_nand3_1 _07306_ (.B(net306),
    .C(net215),
    .A(net259),
    .Y(_02209_));
 sg13g2_o21ai_1 _07307_ (.B1(_02209_),
    .Y(_02210_),
    .A1(net215),
    .A2(net317));
 sg13g2_o21ai_1 _07308_ (.B1(net224),
    .Y(_02211_),
    .A1(_01126_),
    .A2(_02210_));
 sg13g2_nor2_1 _07309_ (.A(net284),
    .B(net182),
    .Y(_02212_));
 sg13g2_a221oi_1 _07310_ (.B2(net180),
    .C1(_02105_),
    .B1(_02212_),
    .A1(net206),
    .Y(_02213_),
    .A2(_00885_));
 sg13g2_a21oi_1 _07311_ (.A1(net259),
    .A2(net309),
    .Y(_02214_),
    .B1(net206));
 sg13g2_o21ai_1 _07312_ (.B1(_00981_),
    .Y(_02215_),
    .A1(net357),
    .A2(_01279_));
 sg13g2_nand2_1 _07313_ (.Y(_02216_),
    .A(net223),
    .B(_02128_));
 sg13g2_a21oi_1 _07314_ (.A1(_02090_),
    .A2(_01128_),
    .Y(_02217_),
    .B1(_02216_));
 sg13g2_a21oi_1 _07315_ (.A1(_02214_),
    .A2(_02215_),
    .Y(_02218_),
    .B1(_02217_));
 sg13g2_o21ai_1 _07316_ (.B1(_02218_),
    .Y(_02219_),
    .A1(net339),
    .A2(_02213_));
 sg13g2_nand2_1 _07317_ (.Y(_02220_),
    .A(net306),
    .B(net302));
 sg13g2_a21oi_1 _07318_ (.A1(net171),
    .A2(_02220_),
    .Y(_02221_),
    .B1(_02216_));
 sg13g2_and3_1 _07319_ (.X(_02222_),
    .A(net317),
    .B(net171),
    .C(_01105_));
 sg13g2_o21ai_1 _07320_ (.B1(net300),
    .Y(_02223_),
    .A1(_02221_),
    .A2(_02222_));
 sg13g2_a21oi_1 _07321_ (.A1(net223),
    .A2(_02190_),
    .Y(_02224_),
    .B1(_01421_));
 sg13g2_o21ai_1 _07322_ (.B1(_02224_),
    .Y(_02225_),
    .A1(_01788_),
    .A2(_02120_));
 sg13g2_a21oi_1 _07323_ (.A1(net223),
    .A2(_00950_),
    .Y(_02226_),
    .B1(_01285_));
 sg13g2_a21oi_1 _07324_ (.A1(_02120_),
    .A2(_02123_),
    .Y(_02227_),
    .B1(_02187_));
 sg13g2_nor3_1 _07325_ (.A(net200),
    .B(_02226_),
    .C(_02227_),
    .Y(_02228_));
 sg13g2_o21ai_1 _07326_ (.B1(net265),
    .Y(_02229_),
    .A1(_02225_),
    .A2(_02228_));
 sg13g2_nand3_1 _07327_ (.B(_02223_),
    .C(_02229_),
    .A(net266),
    .Y(_02230_));
 sg13g2_o21ai_1 _07328_ (.B1(_02230_),
    .Y(_02231_),
    .A1(_02211_),
    .A2(_02219_));
 sg13g2_nand2_1 _07329_ (.Y(_02232_),
    .A(net294),
    .B(net196));
 sg13g2_o21ai_1 _07330_ (.B1(_02232_),
    .Y(_00296_),
    .A1(_02142_),
    .A2(_02231_));
 sg13g2_nor3_1 _07331_ (.A(net201),
    .B(net351),
    .C(net353),
    .Y(_02233_));
 sg13g2_nand2_1 _07332_ (.Y(_02234_),
    .A(net171),
    .B(_02233_));
 sg13g2_o21ai_1 _07333_ (.B1(_02234_),
    .Y(_02235_),
    .A1(_02128_),
    .A2(net171));
 sg13g2_and2_1 _07334_ (.A(_02138_),
    .B(_02235_),
    .X(_02236_));
 sg13g2_nor2_1 _07335_ (.A(net300),
    .B(_00886_),
    .Y(_02237_));
 sg13g2_a21oi_1 _07336_ (.A1(_01278_),
    .A2(_02236_),
    .Y(_02238_),
    .B1(_02237_));
 sg13g2_nor3_1 _07337_ (.A(net260),
    .B(_02122_),
    .C(_02236_),
    .Y(_02239_));
 sg13g2_a21o_1 _07338_ (.A2(_02238_),
    .A1(net260),
    .B1(_02239_),
    .X(_02240_));
 sg13g2_buf_1 _07339_ (.A(_01453_),
    .X(_02241_));
 sg13g2_nand2_1 _07340_ (.Y(_02242_),
    .A(net333),
    .B(net196));
 sg13g2_o21ai_1 _07341_ (.B1(_02242_),
    .Y(_00297_),
    .A1(_02142_),
    .A2(_02240_));
 sg13g2_a21oi_1 _07342_ (.A1(net115),
    .A2(_01346_),
    .Y(_02243_),
    .B1(_01317_));
 sg13g2_buf_1 _07343_ (.A(_02243_),
    .X(_02244_));
 sg13g2_buf_1 _07344_ (.A(_02244_),
    .X(_02245_));
 sg13g2_buf_1 _07345_ (.A(net168),
    .X(_02246_));
 sg13g2_buf_1 _07346_ (.A(net168),
    .X(_02247_));
 sg13g2_nand2_2 _07347_ (.Y(_02248_),
    .A(net276),
    .B(_01354_));
 sg13g2_nor2_1 _07348_ (.A(_01166_),
    .B(_02248_),
    .Y(_02249_));
 sg13g2_inv_1 _07349_ (.Y(_02250_),
    .A(_02249_));
 sg13g2_inv_1 _07350_ (.Y(_02251_),
    .A(_01354_));
 sg13g2_o21ai_1 _07351_ (.B1(_00747_),
    .Y(_02252_),
    .A1(_00930_),
    .A2(net322));
 sg13g2_nand3_1 _07352_ (.B(_00811_),
    .C(_02252_),
    .A(net245),
    .Y(_02253_));
 sg13g2_buf_1 _07353_ (.A(_02253_),
    .X(_02254_));
 sg13g2_nor2_1 _07354_ (.A(_01349_),
    .B(_01357_),
    .Y(_02255_));
 sg13g2_nor3_1 _07355_ (.A(_00878_),
    .B(net210),
    .C(_01282_),
    .Y(_02256_));
 sg13g2_o21ai_1 _07356_ (.B1(_01281_),
    .Y(_02257_),
    .A1(_02255_),
    .A2(_02256_));
 sg13g2_o21ai_1 _07357_ (.B1(_02257_),
    .Y(_02258_),
    .A1(_02251_),
    .A2(_02254_));
 sg13g2_nor2_1 _07358_ (.A(_01352_),
    .B(_00979_),
    .Y(_02259_));
 sg13g2_nand3_1 _07359_ (.B(_01558_),
    .C(_02259_),
    .A(_00808_),
    .Y(_02260_));
 sg13g2_buf_1 _07360_ (.A(_02260_),
    .X(_02261_));
 sg13g2_nand2_1 _07361_ (.Y(_02262_),
    .A(_00877_),
    .B(_01329_));
 sg13g2_a21o_1 _07362_ (.A2(_02262_),
    .A1(_01062_),
    .B1(_00831_),
    .X(_02263_));
 sg13g2_o21ai_1 _07363_ (.B1(_01044_),
    .Y(_02264_),
    .A1(net245),
    .A2(_01077_));
 sg13g2_nand2_1 _07364_ (.Y(_02265_),
    .A(_02263_),
    .B(_02264_));
 sg13g2_or2_1 _07365_ (.X(_02266_),
    .B(_01075_),
    .A(_01047_));
 sg13g2_buf_1 _07366_ (.A(_02266_),
    .X(_02267_));
 sg13g2_nand2_2 _07367_ (.Y(_02268_),
    .A(net274),
    .B(_01151_));
 sg13g2_nand2b_1 _07368_ (.Y(_02269_),
    .B(_02268_),
    .A_N(_02267_));
 sg13g2_o21ai_1 _07369_ (.B1(_00720_),
    .Y(_02270_),
    .A1(_00883_),
    .A2(_00734_));
 sg13g2_or4_1 _07370_ (.A(_02261_),
    .B(_02265_),
    .C(_02269_),
    .D(_02270_),
    .X(_02271_));
 sg13g2_buf_1 _07371_ (.A(_02271_),
    .X(_02272_));
 sg13g2_a21o_1 _07372_ (.A2(net230),
    .A1(_01429_),
    .B1(_02111_),
    .X(_02273_));
 sg13g2_inv_1 _07373_ (.Y(_02274_),
    .A(_00675_));
 sg13g2_nor2_1 _07374_ (.A(net234),
    .B(_02161_),
    .Y(_02275_));
 sg13g2_buf_1 _07375_ (.A(_00026_),
    .X(_02276_));
 sg13g2_nor2_2 _07376_ (.A(net360),
    .B(_01281_),
    .Y(_02277_));
 sg13g2_nand2b_1 _07377_ (.Y(_02278_),
    .B(_02277_),
    .A_N(_00853_));
 sg13g2_nor4_1 _07378_ (.A(net324),
    .B(net394),
    .C(_02276_),
    .D(_02278_),
    .Y(_02279_));
 sg13g2_nand2b_1 _07379_ (.Y(_02280_),
    .B(_02279_),
    .A_N(_01138_));
 sg13g2_nor4_1 _07380_ (.A(_00771_),
    .B(_02255_),
    .C(_02275_),
    .D(_02280_),
    .Y(_02281_));
 sg13g2_nand4_1 _07381_ (.B(_02274_),
    .C(_02254_),
    .A(_00819_),
    .Y(_02282_),
    .D(_02281_));
 sg13g2_nor3_1 _07382_ (.A(_02272_),
    .B(_02273_),
    .C(_02282_),
    .Y(_02283_));
 sg13g2_o21ai_1 _07383_ (.B1(net359),
    .Y(_02284_),
    .A1(_02258_),
    .A2(_02283_));
 sg13g2_nand2_1 _07384_ (.Y(_02285_),
    .A(_02250_),
    .B(_02284_));
 sg13g2_buf_1 _07385_ (.A(_02285_),
    .X(_02286_));
 sg13g2_inv_1 _07386_ (.Y(_02287_),
    .A(_02286_));
 sg13g2_buf_1 _07387_ (.A(_02287_),
    .X(_02288_));
 sg13g2_and2_1 _07388_ (.A(_01137_),
    .B(_01179_),
    .X(_02289_));
 sg13g2_buf_1 _07389_ (.A(_02289_),
    .X(_02290_));
 sg13g2_buf_1 _07390_ (.A(_02290_),
    .X(_02291_));
 sg13g2_buf_1 _07391_ (.A(_01197_),
    .X(_02292_));
 sg13g2_buf_1 _07392_ (.A(net145),
    .X(_02293_));
 sg13g2_buf_1 _07393_ (.A(\z80.tv80s.i_tv80_core.SP[0] ),
    .X(_02294_));
 sg13g2_nand2_1 _07394_ (.Y(_02295_),
    .A(_02294_),
    .B(net138));
 sg13g2_o21ai_1 _07395_ (.B1(_02295_),
    .Y(_02296_),
    .A1(_01452_),
    .A2(net138));
 sg13g2_buf_2 _07396_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .X(_02297_));
 sg13g2_nand2_2 _07397_ (.Y(_02298_),
    .A(net359),
    .B(_01081_));
 sg13g2_nand3_1 _07398_ (.B(_01294_),
    .C(_01435_),
    .A(_01434_),
    .Y(_02299_));
 sg13g2_or3_1 _07399_ (.A(_00802_),
    .B(_02298_),
    .C(_02299_),
    .X(_02300_));
 sg13g2_o21ai_1 _07400_ (.B1(_01057_),
    .Y(_02301_),
    .A1(net279),
    .A2(net240));
 sg13g2_nor3_1 _07401_ (.A(net310),
    .B(net269),
    .C(_00878_),
    .Y(_02302_));
 sg13g2_or3_1 _07402_ (.A(_01578_),
    .B(_01584_),
    .C(_02302_),
    .X(_02303_));
 sg13g2_nor4_1 _07403_ (.A(_01420_),
    .B(_02300_),
    .C(_02301_),
    .D(_02303_),
    .Y(_02304_));
 sg13g2_o21ai_1 _07404_ (.B1(_01369_),
    .Y(_02305_),
    .A1(_01273_),
    .A2(_02304_));
 sg13g2_buf_1 _07405_ (.A(_02305_),
    .X(_02306_));
 sg13g2_buf_1 _07406_ (.A(_02306_),
    .X(_02307_));
 sg13g2_buf_1 _07407_ (.A(net137),
    .X(_02308_));
 sg13g2_xor2_1 _07408_ (.B(_02308_),
    .A(_02297_),
    .X(_02309_));
 sg13g2_nor2_1 _07409_ (.A(_01031_),
    .B(\z80.tv80s.i_tv80_core.XY_State[0] ),
    .Y(_02310_));
 sg13g2_buf_2 _07410_ (.A(_02310_),
    .X(_02311_));
 sg13g2_buf_1 _07411_ (.A(_02311_),
    .X(_02312_));
 sg13g2_buf_1 _07412_ (.A(net352),
    .X(_02313_));
 sg13g2_buf_1 _07413_ (.A(_01029_),
    .X(_02314_));
 sg13g2_buf_2 _07414_ (.A(\z80.tv80s.i_tv80_core.PC[0] ),
    .X(_02315_));
 sg13g2_nor2b_1 _07415_ (.A(_02314_),
    .B_N(_02315_),
    .Y(_02316_));
 sg13g2_a21oi_1 _07416_ (.A1(net293),
    .A2(_02297_),
    .Y(_02317_),
    .B1(_02316_));
 sg13g2_buf_2 _07417_ (.A(\z80.tv80s.i_tv80_core.RegAddrC[1] ),
    .X(_02318_));
 sg13g2_buf_2 _07418_ (.A(\z80.tv80s.i_tv80_core.RegAddrC[0] ),
    .X(_02319_));
 sg13g2_mux4_1 _07419_ (.S0(_02318_),
    .A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .S1(_02319_),
    .X(_02320_));
 sg13g2_mux4_1 _07420_ (.S0(_02318_),
    .A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .S1(_02319_),
    .X(_02321_));
 sg13g2_buf_2 _07421_ (.A(\z80.tv80s.i_tv80_core.RegAddrC[2] ),
    .X(_02322_));
 sg13g2_mux2_1 _07422_ (.A0(_02320_),
    .A1(_02321_),
    .S(_02322_),
    .X(_02323_));
 sg13g2_buf_1 _07423_ (.A(_02323_),
    .X(_02324_));
 sg13g2_nand2_1 _07424_ (.Y(_02325_),
    .A(net254),
    .B(net253));
 sg13g2_o21ai_1 _07425_ (.B1(_02325_),
    .Y(_02326_),
    .A1(net254),
    .A2(_02317_));
 sg13g2_nor2_1 _07426_ (.A(net147),
    .B(_02326_),
    .Y(_02327_));
 sg13g2_a21oi_1 _07427_ (.A1(net147),
    .A2(_02309_),
    .Y(_02328_),
    .B1(_02327_));
 sg13g2_and2_1 _07428_ (.A(_01134_),
    .B(_01179_),
    .X(_02329_));
 sg13g2_and3_1 _07429_ (.X(_02330_),
    .A(_01035_),
    .B(_01131_),
    .C(_02329_));
 sg13g2_buf_1 _07430_ (.A(_02330_),
    .X(_02331_));
 sg13g2_buf_1 _07431_ (.A(_02331_),
    .X(_02332_));
 sg13g2_nand2_1 _07432_ (.Y(_02333_),
    .A(_01134_),
    .B(_01197_));
 sg13g2_nor2_1 _07433_ (.A(_01179_),
    .B(_02333_),
    .Y(_02334_));
 sg13g2_buf_1 _07434_ (.A(_02334_),
    .X(_02335_));
 sg13g2_buf_1 _07435_ (.A(_02335_),
    .X(_02336_));
 sg13g2_nand2_1 _07436_ (.Y(_02337_),
    .A(_00825_),
    .B(\z80.tv80s.i_tv80_core.IStatus[1] ));
 sg13g2_nor2_1 _07437_ (.A(net309),
    .B(_02337_),
    .Y(_02338_));
 sg13g2_buf_1 _07438_ (.A(_02338_),
    .X(_02339_));
 sg13g2_a221oi_1 _07439_ (.B2(_02315_),
    .C1(_02339_),
    .B1(_02336_),
    .A1(net253),
    .Y(_02340_),
    .A2(net113));
 sg13g2_inv_1 _07440_ (.Y(_02341_),
    .A(_02340_));
 sg13g2_a221oi_1 _07441_ (.B2(_01199_),
    .C1(_02341_),
    .B1(_02328_),
    .A1(net114),
    .Y(_02342_),
    .A2(_02296_));
 sg13g2_nand3_1 _07442_ (.B(_00825_),
    .C(\z80.tv80s.i_tv80_core.IStatus[1] ),
    .A(net357),
    .Y(_02343_));
 sg13g2_buf_1 _07443_ (.A(_02343_),
    .X(_02344_));
 sg13g2_buf_1 _07444_ (.A(net252),
    .X(_02345_));
 sg13g2_nor3_1 _07445_ (.A(_01153_),
    .B(_01433_),
    .C(_01581_),
    .Y(_02346_));
 sg13g2_buf_1 _07446_ (.A(_02346_),
    .X(_02347_));
 sg13g2_nor3_1 _07447_ (.A(net258),
    .B(\z80.tv80s.i_tv80_core.mcycles[1] ),
    .C(\z80.tv80s.i_tv80_core.mcycles[2] ),
    .Y(_02348_));
 sg13g2_nor2_1 _07448_ (.A(\z80.tv80s.i_tv80_core.mcycles[4] ),
    .B(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .Y(_02349_));
 sg13g2_a22oi_1 _07449_ (.Y(_02350_),
    .B1(\z80.tv80s.i_tv80_core.mcycles[2] ),
    .B2(net270),
    .A2(\z80.tv80s.i_tv80_core.mcycles[1] ),
    .A1(_00850_));
 sg13g2_a22oi_1 _07450_ (.Y(_02351_),
    .B1(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .B2(net357),
    .A2(\z80.tv80s.i_tv80_core.mcycles[4] ),
    .A1(_00852_));
 sg13g2_nand2_1 _07451_ (.Y(_02352_),
    .A(_02350_),
    .B(_02351_));
 sg13g2_a21oi_1 _07452_ (.A1(_02348_),
    .A2(_02349_),
    .Y(_02353_),
    .B1(_02352_));
 sg13g2_nor2b_1 _07453_ (.A(_02353_),
    .B_N(net394),
    .Y(_02354_));
 sg13g2_buf_1 _07454_ (.A(_02354_),
    .X(_02355_));
 sg13g2_or2_1 _07455_ (.X(_02356_),
    .B(_01414_),
    .A(_01408_));
 sg13g2_buf_1 _07456_ (.A(_02356_),
    .X(_02357_));
 sg13g2_or2_1 _07457_ (.X(_02358_),
    .B(_01565_),
    .A(_01553_));
 sg13g2_nand3_1 _07458_ (.B(_00655_),
    .C(_00730_),
    .A(_00756_),
    .Y(_02359_));
 sg13g2_nand2b_1 _07459_ (.Y(_02360_),
    .B(_02359_),
    .A_N(net205));
 sg13g2_nor4_1 _07460_ (.A(_00802_),
    .B(_00807_),
    .C(net208),
    .D(_02360_),
    .Y(_02361_));
 sg13g2_buf_1 _07461_ (.A(_02361_),
    .X(_02362_));
 sg13g2_nand3_1 _07462_ (.B(_01571_),
    .C(_02362_),
    .A(_01549_),
    .Y(_02363_));
 sg13g2_nor4_1 _07463_ (.A(_02357_),
    .B(_01559_),
    .C(_02358_),
    .D(_02363_),
    .Y(_02364_));
 sg13g2_nand2b_1 _07464_ (.Y(_02365_),
    .B(_01292_),
    .A_N(_02255_));
 sg13g2_nor4_1 _07465_ (.A(_02278_),
    .B(_02298_),
    .C(_02301_),
    .D(_02365_),
    .Y(_02366_));
 sg13g2_nand2_1 _07466_ (.Y(_02367_),
    .A(_02364_),
    .B(_02366_));
 sg13g2_inv_1 _07467_ (.Y(_02368_),
    .A(_01581_));
 sg13g2_nand2_1 _07468_ (.Y(_02369_),
    .A(_00657_),
    .B(_01444_));
 sg13g2_nor2_1 _07469_ (.A(_02369_),
    .B(_02273_),
    .Y(_02370_));
 sg13g2_nand4_1 _07470_ (.B(_01354_),
    .C(_02368_),
    .A(net359),
    .Y(_02371_),
    .D(_02370_));
 sg13g2_nand2_1 _07471_ (.Y(_02372_),
    .A(_02367_),
    .B(_02371_));
 sg13g2_buf_2 _07472_ (.A(_02372_),
    .X(_02373_));
 sg13g2_or2_1 _07473_ (.X(_02374_),
    .B(_02373_),
    .A(_02355_));
 sg13g2_buf_1 _07474_ (.A(_02374_),
    .X(_02375_));
 sg13g2_nor2_1 _07475_ (.A(_02347_),
    .B(net85),
    .Y(_02376_));
 sg13g2_o21ai_1 _07476_ (.B1(_02376_),
    .Y(_02377_),
    .A1(_02297_),
    .A2(net213));
 sg13g2_buf_1 _07477_ (.A(_02347_),
    .X(_02378_));
 sg13g2_nand2_1 _07478_ (.Y(_02379_),
    .A(net253),
    .B(net127));
 sg13g2_o21ai_1 _07479_ (.B1(_02379_),
    .Y(_02380_),
    .A1(_02342_),
    .A2(_02377_));
 sg13g2_nand2_1 _07480_ (.Y(_02381_),
    .A(net99),
    .B(_02380_));
 sg13g2_or3_1 _07481_ (.A(_01153_),
    .B(_01433_),
    .C(_01581_),
    .X(_02382_));
 sg13g2_buf_1 _07482_ (.A(_02382_),
    .X(_02383_));
 sg13g2_a21o_1 _07483_ (.A2(_02373_),
    .A1(net136),
    .B1(_02286_),
    .X(_02384_));
 sg13g2_buf_2 _07484_ (.A(_02384_),
    .X(_02385_));
 sg13g2_nand2_1 _07485_ (.Y(_02386_),
    .A(_02297_),
    .B(_02385_));
 sg13g2_nand3_1 _07486_ (.B(_02381_),
    .C(_02386_),
    .A(net158),
    .Y(_02387_));
 sg13g2_o21ai_1 _07487_ (.B1(_02387_),
    .Y(_02388_),
    .A1(_01606_),
    .A2(net159));
 sg13g2_buf_1 _07488_ (.A(_02244_),
    .X(_02389_));
 sg13g2_nand2_1 _07489_ (.Y(_02390_),
    .A(\addr_bus[0] ),
    .B(_02389_));
 sg13g2_o21ai_1 _07490_ (.B1(_02390_),
    .Y(_00298_),
    .A1(net71),
    .A2(_02388_));
 sg13g2_nor2_1 _07491_ (.A(_01740_),
    .B(net168),
    .Y(_02391_));
 sg13g2_buf_1 _07492_ (.A(_02286_),
    .X(_02392_));
 sg13g2_buf_1 _07493_ (.A(net111),
    .X(_02393_));
 sg13g2_buf_1 _07494_ (.A(_02347_),
    .X(_02394_));
 sg13g2_buf_1 _07495_ (.A(_02322_),
    .X(_02395_));
 sg13g2_buf_1 _07496_ (.A(net331),
    .X(_02396_));
 sg13g2_buf_1 _07497_ (.A(_02318_),
    .X(_02397_));
 sg13g2_buf_2 _07498_ (.A(net330),
    .X(_02398_));
 sg13g2_buf_1 _07499_ (.A(_02319_),
    .X(_02399_));
 sg13g2_buf_1 _07500_ (.A(_02399_),
    .X(_02400_));
 sg13g2_mux4_1 _07501_ (.S0(net291),
    .A0(_00051_),
    .A1(_00053_),
    .A2(_00052_),
    .A3(_00054_),
    .S1(net290),
    .X(_02401_));
 sg13g2_mux4_1 _07502_ (.S0(net291),
    .A0(_00047_),
    .A1(_00049_),
    .A2(_00048_),
    .A3(_00050_),
    .S1(net290),
    .X(_02402_));
 sg13g2_nor2b_1 _07503_ (.A(net292),
    .B_N(_02402_),
    .Y(_02403_));
 sg13g2_a21oi_2 _07504_ (.B1(_02403_),
    .Y(_02404_),
    .A2(_02401_),
    .A1(net292));
 sg13g2_inv_1 _07505_ (.Y(_02405_),
    .A(_02404_));
 sg13g2_a21oi_1 _07506_ (.A1(net126),
    .A2(_02405_),
    .Y(_02406_),
    .B1(_02392_));
 sg13g2_buf_1 _07507_ (.A(_01201_),
    .X(_02407_));
 sg13g2_buf_1 _07508_ (.A(net304),
    .X(_02408_));
 sg13g2_nand2_1 _07509_ (.Y(_02409_),
    .A(net293),
    .B(_00144_));
 sg13g2_buf_1 _07510_ (.A(_00145_),
    .X(_02410_));
 sg13g2_nand2b_1 _07511_ (.Y(_02411_),
    .B(_02410_),
    .A_N(net293));
 sg13g2_nand3_1 _07512_ (.B(_02409_),
    .C(_02411_),
    .A(net251),
    .Y(_02412_));
 sg13g2_o21ai_1 _07513_ (.B1(_02412_),
    .Y(_02413_),
    .A1(net251),
    .A2(_02405_));
 sg13g2_mux2_1 _07514_ (.A0(_01736_),
    .A1(\z80.tv80s.i_tv80_core.SP[10] ),
    .S(_02293_),
    .X(_02414_));
 sg13g2_and2_1 _07515_ (.A(net147),
    .B(_01199_),
    .X(_02415_));
 sg13g2_buf_1 _07516_ (.A(_02415_),
    .X(_02416_));
 sg13g2_buf_1 _07517_ (.A(_02416_),
    .X(_02417_));
 sg13g2_inv_1 _07518_ (.Y(_02418_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sg13g2_buf_1 _07519_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .X(_02419_));
 sg13g2_buf_1 _07520_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .X(_02420_));
 sg13g2_buf_1 _07521_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .X(_02421_));
 sg13g2_buf_2 _07522_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .X(_02422_));
 sg13g2_and2_1 _07523_ (.A(_02421_),
    .B(_02422_),
    .X(_02423_));
 sg13g2_buf_1 _07524_ (.A(_02423_),
    .X(_02424_));
 sg13g2_nand4_1 _07525_ (.B(_02419_),
    .C(_02420_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .Y(_02425_),
    .D(_02424_));
 sg13g2_buf_2 _07526_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .X(_02426_));
 sg13g2_nand2_2 _07527_ (.Y(_02427_),
    .A(_02426_),
    .B(_02297_));
 sg13g2_nor3_2 _07528_ (.A(_02418_),
    .B(_02425_),
    .C(_02427_),
    .Y(_02428_));
 sg13g2_and3_1 _07529_ (.X(_02429_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .C(_02428_));
 sg13g2_buf_1 _07530_ (.A(_02429_),
    .X(_02430_));
 sg13g2_xnor2_1 _07531_ (.Y(_02431_),
    .A(_00144_),
    .B(_02430_));
 sg13g2_nor2_1 _07532_ (.A(_02307_),
    .B(_02431_),
    .Y(_02432_));
 sg13g2_a21oi_1 _07533_ (.A1(_00143_),
    .A2(net128),
    .Y(_02433_),
    .B1(_02432_));
 sg13g2_nand2_1 _07534_ (.Y(_02434_),
    .A(_02417_),
    .B(_02433_));
 sg13g2_buf_2 _07535_ (.A(\z80.tv80s.i_tv80_core.PC[10] ),
    .X(_02435_));
 sg13g2_buf_1 _07536_ (.A(_02335_),
    .X(_02436_));
 sg13g2_a221oi_1 _07537_ (.B2(net113),
    .C1(_02339_),
    .B1(_02404_),
    .A1(_02435_),
    .Y(_02437_),
    .A2(net110));
 sg13g2_nand2_1 _07538_ (.Y(_02438_),
    .A(_02434_),
    .B(_02437_));
 sg13g2_a221oi_1 _07539_ (.B2(_02291_),
    .C1(_02438_),
    .B1(_02414_),
    .A1(net97),
    .Y(_02439_),
    .A2(_02413_));
 sg13g2_nor2_1 _07540_ (.A(_02355_),
    .B(_02373_),
    .Y(_02440_));
 sg13g2_buf_1 _07541_ (.A(_02440_),
    .X(_02441_));
 sg13g2_o21ai_1 _07542_ (.B1(net84),
    .Y(_02442_),
    .A1(_01740_),
    .A2(net213));
 sg13g2_buf_1 _07543_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .X(_02443_));
 sg13g2_buf_1 _07544_ (.A(_02373_),
    .X(_02444_));
 sg13g2_a21oi_1 _07545_ (.A1(_02443_),
    .A2(net95),
    .Y(_02445_),
    .B1(_02347_));
 sg13g2_o21ai_1 _07546_ (.B1(_02445_),
    .Y(_02446_),
    .A1(_02439_),
    .A2(_02442_));
 sg13g2_a221oi_1 _07547_ (.B2(_02446_),
    .C1(net179),
    .B1(_02406_),
    .A1(net389),
    .Y(_02447_),
    .A2(_02393_));
 sg13g2_or2_1 _07548_ (.X(_02448_),
    .B(_02447_),
    .A(_02391_));
 sg13g2_nand2_1 _07549_ (.Y(_02449_),
    .A(\addr_bus[10] ),
    .B(net70));
 sg13g2_o21ai_1 _07550_ (.B1(_02449_),
    .Y(_00299_),
    .A1(net71),
    .A2(_02448_));
 sg13g2_buf_1 _07551_ (.A(net179),
    .X(_02450_));
 sg13g2_mux4_1 _07552_ (.S0(net291),
    .A0(_00059_),
    .A1(_00061_),
    .A2(_00060_),
    .A3(_00062_),
    .S1(net290),
    .X(_02451_));
 sg13g2_mux4_1 _07553_ (.S0(net291),
    .A0(_00055_),
    .A1(_00057_),
    .A2(_00056_),
    .A3(_00058_),
    .S1(net290),
    .X(_02452_));
 sg13g2_nor2b_1 _07554_ (.A(_02396_),
    .B_N(_02452_),
    .Y(_02453_));
 sg13g2_a21o_1 _07555_ (.A2(_02451_),
    .A1(net292),
    .B1(_02453_),
    .X(_02454_));
 sg13g2_a21oi_1 _07556_ (.A1(net127),
    .A2(_02454_),
    .Y(_02455_),
    .B1(net111));
 sg13g2_buf_1 _07557_ (.A(_02339_),
    .X(_02456_));
 sg13g2_and2_1 _07558_ (.A(_01807_),
    .B(net193),
    .X(_02457_));
 sg13g2_buf_2 _07559_ (.A(\z80.tv80s.i_tv80_core.PC[11] ),
    .X(_02458_));
 sg13g2_inv_1 _07560_ (.Y(_02459_),
    .A(_02458_));
 sg13g2_inv_1 _07561_ (.Y(_02460_),
    .A(_00148_));
 sg13g2_nand2_1 _07562_ (.Y(_02461_),
    .A(net332),
    .B(_00147_));
 sg13g2_o21ai_1 _07563_ (.B1(_02461_),
    .Y(_02462_),
    .A1(net332),
    .A2(_02460_));
 sg13g2_buf_1 _07564_ (.A(_02396_),
    .X(_02463_));
 sg13g2_a21oi_1 _07565_ (.A1(net250),
    .A2(_02451_),
    .Y(_02464_),
    .B1(_02453_));
 sg13g2_nand2_1 _07566_ (.Y(_02465_),
    .A(net254),
    .B(_02464_));
 sg13g2_o21ai_1 _07567_ (.B1(_02465_),
    .Y(_02466_),
    .A1(net254),
    .A2(_02462_));
 sg13g2_nand2_1 _07568_ (.Y(_02467_),
    .A(_02443_),
    .B(_02430_));
 sg13g2_xor2_1 _07569_ (.B(_02467_),
    .A(_00147_),
    .X(_02468_));
 sg13g2_nor2_1 _07570_ (.A(net137),
    .B(_02468_),
    .Y(_02469_));
 sg13g2_a21oi_1 _07571_ (.A1(_00146_),
    .A2(net128),
    .Y(_02470_),
    .B1(_02469_));
 sg13g2_a22oi_1 _07572_ (.Y(_02471_),
    .B1(_02470_),
    .B2(net96),
    .A2(_02466_),
    .A1(net97));
 sg13g2_buf_1 _07573_ (.A(\z80.tv80s.i_tv80_core.SP[11] ),
    .X(_02472_));
 sg13g2_mux2_1 _07574_ (.A0(net379),
    .A1(_02472_),
    .S(net138),
    .X(_02473_));
 sg13g2_a221oi_1 _07575_ (.B2(net114),
    .C1(net110),
    .B1(_02473_),
    .A1(net113),
    .Y(_02474_),
    .A2(_02464_));
 sg13g2_a221oi_1 _07576_ (.B2(_02474_),
    .C1(net193),
    .B1(_02471_),
    .A1(_02459_),
    .Y(_02475_),
    .A2(net112));
 sg13g2_o21ai_1 _07577_ (.B1(net84),
    .Y(_02476_),
    .A1(_02457_),
    .A2(_02475_));
 sg13g2_buf_1 _07578_ (.A(_02347_),
    .X(_02477_));
 sg13g2_a21oi_1 _07579_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .A2(net95),
    .Y(_02478_),
    .B1(net125));
 sg13g2_nand2_1 _07580_ (.Y(_02479_),
    .A(_02476_),
    .B(_02478_));
 sg13g2_a22oi_1 _07581_ (.Y(_02480_),
    .B1(_02455_),
    .B2(_02479_),
    .A2(net98),
    .A1(net388));
 sg13g2_nor2_1 _07582_ (.A(_02450_),
    .B(_02480_),
    .Y(_02481_));
 sg13g2_a21oi_1 _07583_ (.A1(_01807_),
    .A2(net165),
    .Y(_02482_),
    .B1(_02481_));
 sg13g2_nand2_1 _07584_ (.Y(_02483_),
    .A(\addr_bus[11] ),
    .B(net70));
 sg13g2_o21ai_1 _07585_ (.B1(_02483_),
    .Y(_00300_),
    .A1(net71),
    .A2(_02482_));
 sg13g2_buf_1 _07586_ (.A(_02286_),
    .X(_02484_));
 sg13g2_buf_1 _07587_ (.A(net291),
    .X(_02485_));
 sg13g2_buf_1 _07588_ (.A(net290),
    .X(_02486_));
 sg13g2_mux4_1 _07589_ (.S0(net249),
    .A0(_00067_),
    .A1(_00069_),
    .A2(_00068_),
    .A3(_00070_),
    .S1(net248),
    .X(_02487_));
 sg13g2_mux4_1 _07590_ (.S0(net249),
    .A0(_00063_),
    .A1(_00065_),
    .A2(_00064_),
    .A3(_00066_),
    .S1(net248),
    .X(_02488_));
 sg13g2_nor2b_1 _07591_ (.A(net292),
    .B_N(_02488_),
    .Y(_02489_));
 sg13g2_a21o_1 _07592_ (.A2(_02487_),
    .A1(net250),
    .B1(_02489_),
    .X(_02490_));
 sg13g2_a21oi_1 _07593_ (.A1(net127),
    .A2(_02490_),
    .Y(_02491_),
    .B1(net111));
 sg13g2_buf_1 _07594_ (.A(_02339_),
    .X(_02492_));
 sg13g2_and2_1 _07595_ (.A(_01868_),
    .B(net192),
    .X(_02493_));
 sg13g2_buf_2 _07596_ (.A(\z80.tv80s.i_tv80_core.PC[12] ),
    .X(_02494_));
 sg13g2_inv_1 _07597_ (.Y(_02495_),
    .A(_02494_));
 sg13g2_buf_1 _07598_ (.A(net304),
    .X(_02496_));
 sg13g2_nand2_1 _07599_ (.Y(_02497_),
    .A(net332),
    .B(_00150_));
 sg13g2_buf_1 _07600_ (.A(_00151_),
    .X(_02498_));
 sg13g2_nand2b_1 _07601_ (.Y(_02499_),
    .B(_02498_),
    .A_N(net352));
 sg13g2_nand3_1 _07602_ (.B(_02497_),
    .C(_02499_),
    .A(net247),
    .Y(_02500_));
 sg13g2_o21ai_1 _07603_ (.B1(_02500_),
    .Y(_02501_),
    .A1(net251),
    .A2(_02490_));
 sg13g2_buf_1 _07604_ (.A(_00149_),
    .X(_02502_));
 sg13g2_nand3_1 _07605_ (.B(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .C(_02430_),
    .A(_02443_),
    .Y(_02503_));
 sg13g2_xor2_1 _07606_ (.B(_02503_),
    .A(_00150_),
    .X(_02504_));
 sg13g2_nor2_1 _07607_ (.A(net137),
    .B(_02504_),
    .Y(_02505_));
 sg13g2_a21oi_1 _07608_ (.A1(_02502_),
    .A2(net128),
    .Y(_02506_),
    .B1(_02505_));
 sg13g2_a22oi_1 _07609_ (.Y(_02507_),
    .B1(_02506_),
    .B2(net96),
    .A2(_02501_),
    .A1(net97));
 sg13g2_a21oi_1 _07610_ (.A1(net250),
    .A2(_02487_),
    .Y(_02508_),
    .B1(_02489_));
 sg13g2_buf_1 _07611_ (.A(\z80.tv80s.i_tv80_core.SP[12] ),
    .X(_02509_));
 sg13g2_mux2_1 _07612_ (.A0(_01864_),
    .A1(_02509_),
    .S(net138),
    .X(_02510_));
 sg13g2_a221oi_1 _07613_ (.B2(net114),
    .C1(net110),
    .B1(_02510_),
    .A1(net113),
    .Y(_02511_),
    .A2(_02508_));
 sg13g2_a221oi_1 _07614_ (.B2(_02511_),
    .C1(net193),
    .B1(_02507_),
    .A1(_02495_),
    .Y(_02512_),
    .A2(net112));
 sg13g2_o21ai_1 _07615_ (.B1(net84),
    .Y(_02513_),
    .A1(_02493_),
    .A2(_02512_));
 sg13g2_a21oi_1 _07616_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .A2(net95),
    .Y(_02514_),
    .B1(net125));
 sg13g2_nand2_1 _07617_ (.Y(_02515_),
    .A(_02513_),
    .B(_02514_));
 sg13g2_a22oi_1 _07618_ (.Y(_02516_),
    .B1(_02491_),
    .B2(_02515_),
    .A2(net109),
    .A1(net387));
 sg13g2_nor2_1 _07619_ (.A(net165),
    .B(_02516_),
    .Y(_02517_));
 sg13g2_a21oi_1 _07620_ (.A1(_01868_),
    .A2(net165),
    .Y(_02518_),
    .B1(_02517_));
 sg13g2_nand2_1 _07621_ (.Y(_02519_),
    .A(\addr_bus[12] ),
    .B(net70));
 sg13g2_o21ai_1 _07622_ (.B1(_02519_),
    .Y(_00301_),
    .A1(net71),
    .A2(_02518_));
 sg13g2_mux4_1 _07623_ (.S0(net249),
    .A0(_00075_),
    .A1(_00077_),
    .A2(_00076_),
    .A3(_00078_),
    .S1(net248),
    .X(_02520_));
 sg13g2_mux4_1 _07624_ (.S0(net249),
    .A0(_00071_),
    .A1(_00073_),
    .A2(_00072_),
    .A3(_00074_),
    .S1(net248),
    .X(_02521_));
 sg13g2_nor2b_1 _07625_ (.A(net292),
    .B_N(_02521_),
    .Y(_02522_));
 sg13g2_a21oi_2 _07626_ (.B1(_02522_),
    .Y(_02523_),
    .A2(_02520_),
    .A1(net250));
 sg13g2_inv_1 _07627_ (.Y(_02524_),
    .A(_02523_));
 sg13g2_a21oi_1 _07628_ (.A1(net127),
    .A2(_02524_),
    .Y(_02525_),
    .B1(net111));
 sg13g2_and2_1 _07629_ (.A(_01953_),
    .B(net192),
    .X(_02526_));
 sg13g2_buf_2 _07630_ (.A(\z80.tv80s.i_tv80_core.PC[13] ),
    .X(_02527_));
 sg13g2_inv_1 _07631_ (.Y(_02528_),
    .A(_02527_));
 sg13g2_nand2_1 _07632_ (.Y(_02529_),
    .A(net332),
    .B(_00153_));
 sg13g2_buf_1 _07633_ (.A(_00154_),
    .X(_02530_));
 sg13g2_nand2b_1 _07634_ (.Y(_02531_),
    .B(_02530_),
    .A_N(net352));
 sg13g2_nand3_1 _07635_ (.B(_02529_),
    .C(_02531_),
    .A(net247),
    .Y(_02532_));
 sg13g2_o21ai_1 _07636_ (.B1(_02532_),
    .Y(_02533_),
    .A1(net251),
    .A2(_02524_));
 sg13g2_inv_1 _07637_ (.Y(_02534_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[12] ));
 sg13g2_nor2_1 _07638_ (.A(_02534_),
    .B(_02503_),
    .Y(_02535_));
 sg13g2_xnor2_1 _07639_ (.Y(_02536_),
    .A(_00153_),
    .B(_02535_));
 sg13g2_nor2_1 _07640_ (.A(net137),
    .B(_02536_),
    .Y(_02537_));
 sg13g2_a21oi_1 _07641_ (.A1(_00152_),
    .A2(net128),
    .Y(_02538_),
    .B1(_02537_));
 sg13g2_a22oi_1 _07642_ (.Y(_02539_),
    .B1(_02538_),
    .B2(net96),
    .A2(_02533_),
    .A1(net97));
 sg13g2_buf_1 _07643_ (.A(\z80.tv80s.i_tv80_core.SP[13] ),
    .X(_02540_));
 sg13g2_mux2_1 _07644_ (.A0(net375),
    .A1(_02540_),
    .S(net145),
    .X(_02541_));
 sg13g2_a221oi_1 _07645_ (.B2(net114),
    .C1(net110),
    .B1(_02541_),
    .A1(net113),
    .Y(_02542_),
    .A2(_02523_));
 sg13g2_a221oi_1 _07646_ (.B2(_02542_),
    .C1(net193),
    .B1(_02539_),
    .A1(_02528_),
    .Y(_02543_),
    .A2(net112));
 sg13g2_o21ai_1 _07647_ (.B1(net84),
    .Y(_02544_),
    .A1(_02526_),
    .A2(_02543_));
 sg13g2_buf_1 _07648_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .X(_02545_));
 sg13g2_a21oi_1 _07649_ (.A1(_02545_),
    .A2(net95),
    .Y(_02546_),
    .B1(net125));
 sg13g2_nand2_1 _07650_ (.Y(_02547_),
    .A(_02544_),
    .B(_02546_));
 sg13g2_a22oi_1 _07651_ (.Y(_02548_),
    .B1(_02525_),
    .B2(_02547_),
    .A2(net109),
    .A1(net386));
 sg13g2_nor2_1 _07652_ (.A(net165),
    .B(_02548_),
    .Y(_02549_));
 sg13g2_a21oi_1 _07653_ (.A1(_01953_),
    .A2(net165),
    .Y(_02550_),
    .B1(_02549_));
 sg13g2_buf_1 _07654_ (.A(_02244_),
    .X(_02551_));
 sg13g2_nand2_1 _07655_ (.Y(_02552_),
    .A(\addr_bus[13] ),
    .B(net69));
 sg13g2_o21ai_1 _07656_ (.B1(_02552_),
    .Y(_00302_),
    .A1(net71),
    .A2(_02550_));
 sg13g2_mux4_1 _07657_ (.S0(net249),
    .A0(_00083_),
    .A1(_00085_),
    .A2(_00084_),
    .A3(_00086_),
    .S1(net248),
    .X(_02553_));
 sg13g2_mux4_1 _07658_ (.S0(net249),
    .A0(_00079_),
    .A1(_00081_),
    .A2(_00080_),
    .A3(_00082_),
    .S1(net248),
    .X(_02554_));
 sg13g2_nor2b_1 _07659_ (.A(net250),
    .B_N(_02554_),
    .Y(_02555_));
 sg13g2_a21oi_2 _07660_ (.B1(_02555_),
    .Y(_02556_),
    .A2(_02553_),
    .A1(net250));
 sg13g2_inv_1 _07661_ (.Y(_02557_),
    .A(_02556_));
 sg13g2_a21oi_1 _07662_ (.A1(net127),
    .A2(_02557_),
    .Y(_02558_),
    .B1(net111));
 sg13g2_and2_1 _07663_ (.A(_02011_),
    .B(net192),
    .X(_02559_));
 sg13g2_buf_1 _07664_ (.A(\z80.tv80s.i_tv80_core.PC[14] ),
    .X(_02560_));
 sg13g2_inv_1 _07665_ (.Y(_02561_),
    .A(_02560_));
 sg13g2_nand2_1 _07666_ (.Y(_02562_),
    .A(net332),
    .B(_00156_));
 sg13g2_nand2b_1 _07667_ (.Y(_02563_),
    .B(_00157_),
    .A_N(net352));
 sg13g2_nand3_1 _07668_ (.B(_02562_),
    .C(_02563_),
    .A(net247),
    .Y(_02564_));
 sg13g2_o21ai_1 _07669_ (.B1(_02564_),
    .Y(_02565_),
    .A1(net251),
    .A2(_02557_));
 sg13g2_buf_1 _07670_ (.A(_00155_),
    .X(_02566_));
 sg13g2_nand2_1 _07671_ (.Y(_02567_),
    .A(_02545_),
    .B(_02535_));
 sg13g2_xor2_1 _07672_ (.B(_02567_),
    .A(_00156_),
    .X(_02568_));
 sg13g2_nor2_1 _07673_ (.A(net137),
    .B(_02568_),
    .Y(_02569_));
 sg13g2_a21oi_1 _07674_ (.A1(_02566_),
    .A2(net128),
    .Y(_02570_),
    .B1(_02569_));
 sg13g2_a22oi_1 _07675_ (.Y(_02571_),
    .B1(_02570_),
    .B2(net96),
    .A2(_02565_),
    .A1(net97));
 sg13g2_buf_1 _07676_ (.A(\z80.tv80s.i_tv80_core.SP[14] ),
    .X(_02572_));
 sg13g2_mux2_1 _07677_ (.A0(_02007_),
    .A1(_02572_),
    .S(net145),
    .X(_02573_));
 sg13g2_a221oi_1 _07678_ (.B2(_02290_),
    .C1(net110),
    .B1(_02573_),
    .A1(_02331_),
    .Y(_02574_),
    .A2(_02556_));
 sg13g2_a221oi_1 _07679_ (.B2(_02574_),
    .C1(net193),
    .B1(_02571_),
    .A1(_02561_),
    .Y(_02575_),
    .A2(net112));
 sg13g2_o21ai_1 _07680_ (.B1(net84),
    .Y(_02576_),
    .A1(_02559_),
    .A2(_02575_));
 sg13g2_a21oi_1 _07681_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .A2(net95),
    .Y(_02577_),
    .B1(net125));
 sg13g2_nand2_1 _07682_ (.Y(_02578_),
    .A(_02576_),
    .B(_02577_));
 sg13g2_a22oi_1 _07683_ (.Y(_02579_),
    .B1(_02558_),
    .B2(_02578_),
    .A2(net109),
    .A1(net385));
 sg13g2_nor2_1 _07684_ (.A(net165),
    .B(_02579_),
    .Y(_02580_));
 sg13g2_a21oi_1 _07685_ (.A1(_02011_),
    .A2(net165),
    .Y(_02581_),
    .B1(_02580_));
 sg13g2_nand2_1 _07686_ (.Y(_02582_),
    .A(\addr_bus[14] ),
    .B(net69));
 sg13g2_o21ai_1 _07687_ (.B1(_02582_),
    .Y(_00303_),
    .A1(net71),
    .A2(_02581_));
 sg13g2_nor2_1 _07688_ (.A(_02080_),
    .B(net158),
    .Y(_02583_));
 sg13g2_mux4_1 _07689_ (.S0(net249),
    .A0(_00091_),
    .A1(_00093_),
    .A2(_00092_),
    .A3(_00094_),
    .S1(net248),
    .X(_02584_));
 sg13g2_mux4_1 _07690_ (.S0(_02485_),
    .A0(_00087_),
    .A1(_00089_),
    .A2(_00088_),
    .A3(_00090_),
    .S1(net248),
    .X(_02585_));
 sg13g2_nor2b_1 _07691_ (.A(net292),
    .B_N(_02585_),
    .Y(_02586_));
 sg13g2_a21o_1 _07692_ (.A2(_02584_),
    .A1(net250),
    .B1(_02586_),
    .X(_02587_));
 sg13g2_buf_1 _07693_ (.A(_02587_),
    .X(_02588_));
 sg13g2_a21oi_1 _07694_ (.A1(net127),
    .A2(_02588_),
    .Y(_02589_),
    .B1(net111));
 sg13g2_buf_1 _07695_ (.A(net192),
    .X(_02590_));
 sg13g2_inv_1 _07696_ (.Y(_02591_),
    .A(\z80.tv80s.i_tv80_core.PC[15] ));
 sg13g2_a21oi_1 _07697_ (.A1(net250),
    .A2(_02584_),
    .Y(_02592_),
    .B1(_02586_));
 sg13g2_buf_1 _07698_ (.A(\z80.tv80s.i_tv80_core.SP[15] ),
    .X(_02593_));
 sg13g2_mux2_1 _07699_ (.A0(_02076_),
    .A1(_02593_),
    .S(net138),
    .X(_02594_));
 sg13g2_a221oi_1 _07700_ (.B2(net114),
    .C1(net112),
    .B1(_02594_),
    .A1(net113),
    .Y(_02595_),
    .A2(_02592_));
 sg13g2_nand2_1 _07701_ (.Y(_02596_),
    .A(net332),
    .B(_00159_));
 sg13g2_nand2b_1 _07702_ (.Y(_02597_),
    .B(_00160_),
    .A_N(net332));
 sg13g2_nand3_1 _07703_ (.B(_02596_),
    .C(_02597_),
    .A(net251),
    .Y(_02598_));
 sg13g2_o21ai_1 _07704_ (.B1(_02598_),
    .Y(_02599_),
    .A1(net251),
    .A2(_02588_));
 sg13g2_nand3_1 _07705_ (.B(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .C(_02535_),
    .A(_02545_),
    .Y(_02600_));
 sg13g2_xor2_1 _07706_ (.B(_02600_),
    .A(_00159_),
    .X(_02601_));
 sg13g2_nor2_1 _07707_ (.A(net137),
    .B(_02601_),
    .Y(_02602_));
 sg13g2_a21oi_1 _07708_ (.A1(_00158_),
    .A2(net128),
    .Y(_02603_),
    .B1(_02602_));
 sg13g2_a22oi_1 _07709_ (.Y(_02604_),
    .B1(_02603_),
    .B2(net96),
    .A2(_02599_),
    .A1(net97));
 sg13g2_a221oi_1 _07710_ (.B2(_02604_),
    .C1(net174),
    .B1(_02595_),
    .A1(_02591_),
    .Y(_02605_),
    .A2(net112));
 sg13g2_a21oi_1 _07711_ (.A1(_02080_),
    .A2(net174),
    .Y(_02606_),
    .B1(_02605_));
 sg13g2_a21oi_1 _07712_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .A2(_02373_),
    .Y(_02607_),
    .B1(_02347_));
 sg13g2_o21ai_1 _07713_ (.B1(_02607_),
    .Y(_02608_),
    .A1(net85),
    .A2(_02606_));
 sg13g2_buf_1 _07714_ (.A(net179),
    .X(_02609_));
 sg13g2_a221oi_1 _07715_ (.B2(_02608_),
    .C1(net164),
    .B1(_02589_),
    .A1(net349),
    .Y(_02610_),
    .A2(net98));
 sg13g2_nor3_1 _07716_ (.A(net69),
    .B(_02583_),
    .C(_02610_),
    .Y(_02611_));
 sg13g2_a21o_1 _07717_ (.A2(net70),
    .A1(\addr_bus[15] ),
    .B1(_02611_),
    .X(_00304_));
 sg13g2_nor2_1 _07718_ (.A(\z80.tv80s.i_tv80_core.R[1] ),
    .B(net158),
    .Y(_02612_));
 sg13g2_o21ai_1 _07719_ (.B1(net136),
    .Y(_02613_),
    .A1(net174),
    .A2(_02373_));
 sg13g2_nand2_1 _07720_ (.Y(_02614_),
    .A(net99),
    .B(_02613_));
 sg13g2_mux4_1 _07721_ (.S0(net329),
    .A0(_00161_),
    .A1(_00162_),
    .A2(_00163_),
    .A3(_00164_),
    .S1(net330),
    .X(_02615_));
 sg13g2_mux4_1 _07722_ (.S0(net329),
    .A0(_00165_),
    .A1(_00166_),
    .A2(_00167_),
    .A3(_00168_),
    .S1(_02318_),
    .X(_02616_));
 sg13g2_mux2_1 _07723_ (.A0(_02615_),
    .A1(_02616_),
    .S(_02322_),
    .X(_02617_));
 sg13g2_buf_2 _07724_ (.A(_02617_),
    .X(_02618_));
 sg13g2_buf_1 _07725_ (.A(\z80.tv80s.i_tv80_core.PC[1] ),
    .X(_02619_));
 sg13g2_inv_1 _07726_ (.Y(_02620_),
    .A(_02619_));
 sg13g2_nand2_1 _07727_ (.Y(_02621_),
    .A(net352),
    .B(_00169_));
 sg13g2_nand2b_1 _07728_ (.Y(_02622_),
    .B(_00170_),
    .A_N(net352));
 sg13g2_nand3_1 _07729_ (.B(_02621_),
    .C(_02622_),
    .A(net304),
    .Y(_02623_));
 sg13g2_o21ai_1 _07730_ (.B1(_02623_),
    .Y(_02624_),
    .A1(net247),
    .A2(_02618_));
 sg13g2_xor2_1 _07731_ (.B(_02297_),
    .A(_02426_),
    .X(_02625_));
 sg13g2_nor2_1 _07732_ (.A(_02306_),
    .B(_02625_),
    .Y(_02626_));
 sg13g2_a21oi_1 _07733_ (.A1(_00169_),
    .A2(net137),
    .Y(_02627_),
    .B1(_02626_));
 sg13g2_a22oi_1 _07734_ (.Y(_02628_),
    .B1(_02627_),
    .B2(_02416_),
    .A2(_02624_),
    .A1(_01201_));
 sg13g2_inv_1 _07735_ (.Y(_02629_),
    .A(_02618_));
 sg13g2_buf_2 _07736_ (.A(\z80.tv80s.i_tv80_core.SP[1] ),
    .X(_02630_));
 sg13g2_mux2_1 _07737_ (.A0(net390),
    .A1(_02630_),
    .S(net145),
    .X(_02631_));
 sg13g2_a221oi_1 _07738_ (.B2(_02290_),
    .C1(net110),
    .B1(_02631_),
    .A1(_02331_),
    .Y(_02632_),
    .A2(_02629_));
 sg13g2_a221oi_1 _07739_ (.B2(_02632_),
    .C1(net192),
    .B1(_02628_),
    .A1(_02620_),
    .Y(_02633_),
    .A2(net112));
 sg13g2_nor2_1 _07740_ (.A(_02355_),
    .B(_02633_),
    .Y(_02634_));
 sg13g2_or3_1 _07741_ (.A(net125),
    .B(net95),
    .C(_02634_),
    .X(_02635_));
 sg13g2_o21ai_1 _07742_ (.B1(_02635_),
    .Y(_02636_),
    .A1(net136),
    .A2(_02618_));
 sg13g2_a221oi_1 _07743_ (.B2(net99),
    .C1(net164),
    .B1(_02636_),
    .A1(_02426_),
    .Y(_02637_),
    .A2(_02614_));
 sg13g2_nor3_1 _07744_ (.A(net69),
    .B(_02612_),
    .C(_02637_),
    .Y(_02638_));
 sg13g2_a21o_1 _07745_ (.A2(net70),
    .A1(\addr_bus[1] ),
    .B1(_02638_),
    .X(_00305_));
 sg13g2_nand2_1 _07746_ (.Y(_02639_),
    .A(net213),
    .B(_02376_));
 sg13g2_buf_2 _07747_ (.A(\z80.tv80s.i_tv80_core.PC[2] ),
    .X(_02640_));
 sg13g2_inv_1 _07748_ (.Y(_02641_),
    .A(_01199_));
 sg13g2_nor2_1 _07749_ (.A(_02306_),
    .B(_02427_),
    .Y(_02642_));
 sg13g2_xnor2_1 _07750_ (.Y(_02643_),
    .A(_00179_),
    .B(_02642_));
 sg13g2_mux4_1 _07751_ (.S0(_02319_),
    .A0(_00175_),
    .A1(_00176_),
    .A2(_00177_),
    .A3(_00178_),
    .S1(_02318_),
    .X(_02644_));
 sg13g2_mux4_1 _07752_ (.S0(_02319_),
    .A0(_00171_),
    .A1(_00172_),
    .A2(_00173_),
    .A3(_00174_),
    .S1(_02318_),
    .X(_02645_));
 sg13g2_nor2b_1 _07753_ (.A(_02322_),
    .B_N(_02645_),
    .Y(_02646_));
 sg13g2_a21oi_2 _07754_ (.B1(_02646_),
    .Y(_02647_),
    .A2(_02644_),
    .A1(_02322_));
 sg13g2_mux2_1 _07755_ (.A0(_00180_),
    .A1(_00179_),
    .S(_01029_),
    .X(_02648_));
 sg13g2_nand2_1 _07756_ (.Y(_02649_),
    .A(net247),
    .B(_02648_));
 sg13g2_o21ai_1 _07757_ (.B1(_02649_),
    .Y(_02650_),
    .A1(net247),
    .A2(_02647_));
 sg13g2_nor2_1 _07758_ (.A(net147),
    .B(_02650_),
    .Y(_02651_));
 sg13g2_a21oi_1 _07759_ (.A1(net147),
    .A2(_02643_),
    .Y(_02652_),
    .B1(_02651_));
 sg13g2_buf_1 _07760_ (.A(\z80.tv80s.i_tv80_core.SP[2] ),
    .X(_02653_));
 sg13g2_mux2_1 _07761_ (.A0(net389),
    .A1(_02653_),
    .S(net138),
    .X(_02654_));
 sg13g2_a22oi_1 _07762_ (.Y(_02655_),
    .B1(_02654_),
    .B2(net114),
    .A2(_02647_),
    .A1(_02332_));
 sg13g2_o21ai_1 _07763_ (.B1(_02655_),
    .Y(_02656_),
    .A1(_02641_),
    .A2(_02652_));
 sg13g2_or2_1 _07764_ (.X(_02657_),
    .B(_02333_),
    .A(_01179_));
 sg13g2_mux2_1 _07765_ (.A0(_02640_),
    .A1(_02656_),
    .S(_02657_),
    .X(_02658_));
 sg13g2_nand2b_1 _07766_ (.Y(_02659_),
    .B(net125),
    .A_N(_02647_));
 sg13g2_o21ai_1 _07767_ (.B1(_02659_),
    .Y(_02660_),
    .A1(_02639_),
    .A2(_02658_));
 sg13g2_nor2_1 _07768_ (.A(net252),
    .B(_02355_),
    .Y(_02661_));
 sg13g2_o21ai_1 _07769_ (.B1(net136),
    .Y(_02662_),
    .A1(_02373_),
    .A2(_02661_));
 sg13g2_nand2_2 _07770_ (.Y(_02663_),
    .A(_02287_),
    .B(_02662_));
 sg13g2_inv_1 _07771_ (.Y(_02664_),
    .A(_02420_));
 sg13g2_a221oi_1 _07772_ (.B2(_02664_),
    .C1(net164),
    .B1(_02663_),
    .A1(net99),
    .Y(_02665_),
    .A2(_02660_));
 sg13g2_a21o_1 _07773_ (.A2(_02450_),
    .A1(_01741_),
    .B1(_02665_),
    .X(_02666_));
 sg13g2_mux2_1 _07774_ (.A0(_02666_),
    .A1(\addr_bus[2] ),
    .S(net70),
    .X(_00306_));
 sg13g2_mux4_1 _07775_ (.S0(net330),
    .A0(_00099_),
    .A1(_00101_),
    .A2(_00100_),
    .A3(_00102_),
    .S1(net329),
    .X(_02667_));
 sg13g2_mux4_1 _07776_ (.S0(_02397_),
    .A0(_00095_),
    .A1(_00097_),
    .A2(_00096_),
    .A3(_00098_),
    .S1(net329),
    .X(_02668_));
 sg13g2_nor2b_1 _07777_ (.A(net331),
    .B_N(_02668_),
    .Y(_02669_));
 sg13g2_a21oi_1 _07778_ (.A1(net331),
    .A2(_02667_),
    .Y(_02670_),
    .B1(_02669_));
 sg13g2_buf_2 _07779_ (.A(_02670_),
    .X(_02671_));
 sg13g2_nand2_1 _07780_ (.Y(_02672_),
    .A(net293),
    .B(net247));
 sg13g2_nor3_2 _07781_ (.A(_02664_),
    .B(_02306_),
    .C(_02427_),
    .Y(_02673_));
 sg13g2_mux2_1 _07782_ (.A0(_02672_),
    .A1(_02673_),
    .S(net147),
    .X(_02674_));
 sg13g2_nand3b_1 _07783_ (.B(_02671_),
    .C(_02312_),
    .Y(_02675_),
    .A_N(net147));
 sg13g2_nand3_1 _07784_ (.B(net147),
    .C(_02673_),
    .A(_00181_),
    .Y(_02676_));
 sg13g2_and2_1 _07785_ (.A(_02675_),
    .B(_02676_),
    .X(_02677_));
 sg13g2_o21ai_1 _07786_ (.B1(_02677_),
    .Y(_02678_),
    .A1(_00181_),
    .A2(_02674_));
 sg13g2_nor2_1 _07787_ (.A(_02314_),
    .B(_02311_),
    .Y(_02679_));
 sg13g2_a21oi_1 _07788_ (.A1(_02679_),
    .A2(_01201_),
    .Y(_02680_),
    .B1(_02335_));
 sg13g2_buf_1 _07789_ (.A(\z80.tv80s.i_tv80_core.SP[3] ),
    .X(_02681_));
 sg13g2_nand2_1 _07790_ (.Y(_02682_),
    .A(_02681_),
    .B(_02292_));
 sg13g2_o21ai_1 _07791_ (.B1(_02682_),
    .Y(_02683_),
    .A1(_01796_),
    .A2(_02292_));
 sg13g2_a221oi_1 _07792_ (.B2(_02331_),
    .C1(_02339_),
    .B1(_02671_),
    .A1(_02290_),
    .Y(_02684_),
    .A2(_02683_));
 sg13g2_o21ai_1 _07793_ (.B1(_02684_),
    .Y(_02685_),
    .A1(_00182_),
    .A2(_02680_));
 sg13g2_a21o_1 _07794_ (.A2(_02678_),
    .A1(_01199_),
    .B1(_02685_),
    .X(_02686_));
 sg13g2_nand2_2 _07795_ (.Y(_02687_),
    .A(net136),
    .B(_02440_));
 sg13g2_a21oi_1 _07796_ (.A1(_00181_),
    .A2(net174),
    .Y(_02688_),
    .B1(_02687_));
 sg13g2_a22oi_1 _07797_ (.Y(_02689_),
    .B1(_02686_),
    .B2(_02688_),
    .A2(_02671_),
    .A1(_02378_));
 sg13g2_nor2_1 _07798_ (.A(net111),
    .B(_02689_),
    .Y(_02690_));
 sg13g2_a21oi_1 _07799_ (.A1(_02422_),
    .A2(_02385_),
    .Y(_02691_),
    .B1(_02690_));
 sg13g2_nand2_1 _07800_ (.Y(_02692_),
    .A(net159),
    .B(_02691_));
 sg13g2_o21ai_1 _07801_ (.B1(_02692_),
    .Y(_02693_),
    .A1(\z80.tv80s.i_tv80_core.R[3] ),
    .A2(net159));
 sg13g2_nand2_1 _07802_ (.Y(_02694_),
    .A(\addr_bus[3] ),
    .B(net69));
 sg13g2_o21ai_1 _07803_ (.B1(_02694_),
    .Y(_00307_),
    .A1(net71),
    .A2(_02693_));
 sg13g2_mux4_1 _07804_ (.S0(net330),
    .A0(_00107_),
    .A1(_00109_),
    .A2(_00108_),
    .A3(_00110_),
    .S1(net329),
    .X(_02695_));
 sg13g2_mux4_1 _07805_ (.S0(net330),
    .A0(_00103_),
    .A1(_00105_),
    .A2(_00104_),
    .A3(_00106_),
    .S1(net329),
    .X(_02696_));
 sg13g2_nor2b_1 _07806_ (.A(net331),
    .B_N(_02696_),
    .Y(_02697_));
 sg13g2_a21o_1 _07807_ (.A2(_02695_),
    .A1(net331),
    .B1(_02697_),
    .X(_02698_));
 sg13g2_buf_1 _07808_ (.A(_02698_),
    .X(_02699_));
 sg13g2_nor2_1 _07809_ (.A(_02383_),
    .B(_02699_),
    .Y(_02700_));
 sg13g2_a21oi_1 _07810_ (.A1(_02463_),
    .A2(_02695_),
    .Y(_02701_),
    .B1(_02697_));
 sg13g2_nand2_1 _07811_ (.Y(_02702_),
    .A(_02422_),
    .B(_02673_));
 sg13g2_xor2_1 _07812_ (.B(_02702_),
    .A(_00183_),
    .X(_02703_));
 sg13g2_o21ai_1 _07813_ (.B1(_02344_),
    .Y(_02704_),
    .A1(_00184_),
    .A2(_02657_));
 sg13g2_a221oi_1 _07814_ (.B2(net96),
    .C1(_02704_),
    .B1(_02703_),
    .A1(net113),
    .Y(_02705_),
    .A2(_02701_));
 sg13g2_nand2_1 _07815_ (.Y(_02706_),
    .A(net293),
    .B(_00183_));
 sg13g2_nand2b_1 _07816_ (.Y(_02707_),
    .B(_00184_),
    .A_N(net293));
 sg13g2_nand3_1 _07817_ (.B(_02706_),
    .C(_02707_),
    .A(_02408_),
    .Y(_02708_));
 sg13g2_o21ai_1 _07818_ (.B1(_02708_),
    .Y(_02709_),
    .A1(_02408_),
    .A2(_02699_));
 sg13g2_buf_1 _07819_ (.A(\z80.tv80s.i_tv80_core.SP[4] ),
    .X(_02710_));
 sg13g2_mux2_1 _07820_ (.A0(net387),
    .A1(_02710_),
    .S(net138),
    .X(_02711_));
 sg13g2_a22oi_1 _07821_ (.Y(_02712_),
    .B1(_02711_),
    .B2(net114),
    .A2(_02709_),
    .A1(_02407_));
 sg13g2_a221oi_1 _07822_ (.B2(_02712_),
    .C1(_02687_),
    .B1(_02705_),
    .A1(_00183_),
    .Y(_02713_),
    .A2(_02590_));
 sg13g2_o21ai_1 _07823_ (.B1(_02288_),
    .Y(_02714_),
    .A1(_02700_),
    .A2(_02713_));
 sg13g2_nand2_1 _07824_ (.Y(_02715_),
    .A(_02421_),
    .B(_02385_));
 sg13g2_nand3_1 _07825_ (.B(_02714_),
    .C(_02715_),
    .A(net158),
    .Y(_02716_));
 sg13g2_o21ai_1 _07826_ (.B1(_02716_),
    .Y(_02717_),
    .A1(\z80.tv80s.i_tv80_core.R[4] ),
    .A2(net159));
 sg13g2_nand2_1 _07827_ (.Y(_02718_),
    .A(\addr_bus[4] ),
    .B(_02551_));
 sg13g2_o21ai_1 _07828_ (.B1(_02718_),
    .Y(_00308_),
    .A1(_02245_),
    .A2(_02717_));
 sg13g2_nor2_1 _07829_ (.A(_01954_),
    .B(_02247_),
    .Y(_02719_));
 sg13g2_mux4_1 _07830_ (.S0(_02398_),
    .A0(_00111_),
    .A1(_00113_),
    .A2(_00112_),
    .A3(_00114_),
    .S1(_02400_),
    .X(_02720_));
 sg13g2_mux4_1 _07831_ (.S0(_02398_),
    .A0(_00115_),
    .A1(_00117_),
    .A2(_00116_),
    .A3(_00118_),
    .S1(_02400_),
    .X(_02721_));
 sg13g2_mux2_1 _07832_ (.A0(_02720_),
    .A1(_02721_),
    .S(net331),
    .X(_02722_));
 sg13g2_buf_2 _07833_ (.A(_02722_),
    .X(_02723_));
 sg13g2_inv_1 _07834_ (.Y(_02724_),
    .A(\z80.tv80s.i_tv80_core.PC[5] ));
 sg13g2_inv_1 _07835_ (.Y(_02725_),
    .A(_02723_));
 sg13g2_buf_2 _07836_ (.A(\z80.tv80s.i_tv80_core.SP[5] ),
    .X(_02726_));
 sg13g2_nand2_1 _07837_ (.Y(_02727_),
    .A(_02726_),
    .B(net145));
 sg13g2_o21ai_1 _07838_ (.B1(_02727_),
    .Y(_02728_),
    .A1(_01944_),
    .A2(net145));
 sg13g2_a221oi_1 _07839_ (.B2(_02290_),
    .C1(net110),
    .B1(_02728_),
    .A1(_02331_),
    .Y(_02729_),
    .A2(_02725_));
 sg13g2_nand2_1 _07840_ (.Y(_02730_),
    .A(net352),
    .B(_00185_));
 sg13g2_nand2b_1 _07841_ (.Y(_02731_),
    .B(_00186_),
    .A_N(_01029_));
 sg13g2_nand3_1 _07842_ (.B(_02730_),
    .C(_02731_),
    .A(net304),
    .Y(_02732_));
 sg13g2_o21ai_1 _07843_ (.B1(_02732_),
    .Y(_02733_),
    .A1(_02496_),
    .A2(_02723_));
 sg13g2_nand2_1 _07844_ (.Y(_02734_),
    .A(_02424_),
    .B(_02673_));
 sg13g2_xor2_1 _07845_ (.B(_02734_),
    .A(_00185_),
    .X(_02735_));
 sg13g2_a22oi_1 _07846_ (.Y(_02736_),
    .B1(_02735_),
    .B2(_02416_),
    .A2(_02733_),
    .A1(_01201_));
 sg13g2_a221oi_1 _07847_ (.B2(_02736_),
    .C1(net192),
    .B1(_02729_),
    .A1(_02724_),
    .Y(_02737_),
    .A2(_02436_));
 sg13g2_nor2_1 _07848_ (.A(_02355_),
    .B(_02737_),
    .Y(_02738_));
 sg13g2_or3_1 _07849_ (.A(_02477_),
    .B(net95),
    .C(_02738_),
    .X(_02739_));
 sg13g2_o21ai_1 _07850_ (.B1(_02739_),
    .Y(_02740_),
    .A1(net136),
    .A2(_02723_));
 sg13g2_a221oi_1 _07851_ (.B2(net99),
    .C1(net164),
    .B1(_02740_),
    .A1(_02419_),
    .Y(_02741_),
    .A2(_02614_));
 sg13g2_nor3_1 _07852_ (.A(net69),
    .B(_02719_),
    .C(_02741_),
    .Y(_02742_));
 sg13g2_a21o_1 _07853_ (.A2(net70),
    .A1(\addr_bus[5] ),
    .B1(_02742_),
    .X(_00309_));
 sg13g2_nor2_1 _07854_ (.A(\z80.tv80s.i_tv80_core.R[6] ),
    .B(_02247_),
    .Y(_02743_));
 sg13g2_mux4_1 _07855_ (.S0(net249),
    .A0(_00119_),
    .A1(_00121_),
    .A2(_00120_),
    .A3(_00122_),
    .S1(_02486_),
    .X(_02744_));
 sg13g2_mux4_1 _07856_ (.S0(net291),
    .A0(_00123_),
    .A1(_00125_),
    .A2(_00124_),
    .A3(_00126_),
    .S1(_02486_),
    .X(_02745_));
 sg13g2_mux2_1 _07857_ (.A0(_02744_),
    .A1(_02745_),
    .S(net292),
    .X(_02746_));
 sg13g2_buf_2 _07858_ (.A(_02746_),
    .X(_02747_));
 sg13g2_inv_1 _07859_ (.Y(_02748_),
    .A(\z80.tv80s.i_tv80_core.PC[6] ));
 sg13g2_nand2_1 _07860_ (.Y(_02749_),
    .A(_01030_),
    .B(_00187_));
 sg13g2_nand2b_1 _07861_ (.Y(_02750_),
    .B(_00188_),
    .A_N(_01029_));
 sg13g2_nand3_1 _07862_ (.B(_02749_),
    .C(_02750_),
    .A(net304),
    .Y(_02751_));
 sg13g2_o21ai_1 _07863_ (.B1(_02751_),
    .Y(_02752_),
    .A1(_02496_),
    .A2(_02747_));
 sg13g2_and4_1 _07864_ (.A(_02419_),
    .B(_02420_),
    .C(_02424_),
    .D(_02642_),
    .X(_02753_));
 sg13g2_xnor2_1 _07865_ (.Y(_02754_),
    .A(_00187_),
    .B(_02753_));
 sg13g2_a22oi_1 _07866_ (.Y(_02755_),
    .B1(_02754_),
    .B2(_02416_),
    .A2(_02752_),
    .A1(_01201_));
 sg13g2_inv_1 _07867_ (.Y(_02756_),
    .A(_02747_));
 sg13g2_buf_2 _07868_ (.A(\z80.tv80s.i_tv80_core.SP[6] ),
    .X(_02757_));
 sg13g2_mux2_1 _07869_ (.A0(\z80.tv80s.di_reg[6] ),
    .A1(_02757_),
    .S(net145),
    .X(_02758_));
 sg13g2_a221oi_1 _07870_ (.B2(_02290_),
    .C1(_02335_),
    .B1(_02758_),
    .A1(_02331_),
    .Y(_02759_),
    .A2(_02756_));
 sg13g2_a221oi_1 _07871_ (.B2(_02759_),
    .C1(_02492_),
    .B1(_02755_),
    .A1(_02748_),
    .Y(_02760_),
    .A2(_02436_));
 sg13g2_nor2_1 _07872_ (.A(_02355_),
    .B(_02760_),
    .Y(_02761_));
 sg13g2_or3_1 _07873_ (.A(net125),
    .B(net95),
    .C(_02761_),
    .X(_02762_));
 sg13g2_o21ai_1 _07874_ (.B1(_02762_),
    .Y(_02763_),
    .A1(net136),
    .A2(_02747_));
 sg13g2_a221oi_1 _07875_ (.B2(net99),
    .C1(net164),
    .B1(_02763_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .Y(_02764_),
    .A2(_02614_));
 sg13g2_nor3_1 _07876_ (.A(net69),
    .B(_02743_),
    .C(_02764_),
    .Y(_02765_));
 sg13g2_a21o_1 _07877_ (.A2(net70),
    .A1(\addr_bus[6] ),
    .B1(_02765_),
    .X(_00310_));
 sg13g2_buf_1 _07878_ (.A(\z80.tv80s.i_tv80_core.SP[7] ),
    .X(_02766_));
 sg13g2_mux2_1 _07879_ (.A0(_01400_),
    .A1(_02766_),
    .S(net138),
    .X(_02767_));
 sg13g2_nand2b_1 _07880_ (.Y(_02768_),
    .B(_02313_),
    .A_N(_00189_));
 sg13g2_mux4_1 _07881_ (.S0(net330),
    .A0(_00131_),
    .A1(_00133_),
    .A2(_00132_),
    .A3(_00134_),
    .S1(net329),
    .X(_02769_));
 sg13g2_inv_1 _07882_ (.Y(_02770_),
    .A(_00128_));
 sg13g2_inv_1 _07883_ (.Y(_02771_),
    .A(_00127_));
 sg13g2_inv_1 _07884_ (.Y(_02772_),
    .A(_00130_));
 sg13g2_inv_1 _07885_ (.Y(_02773_),
    .A(_00129_));
 sg13g2_inv_1 _07886_ (.Y(_02774_),
    .A(_02399_));
 sg13g2_mux4_1 _07887_ (.S0(_02774_),
    .A0(_02770_),
    .A1(_02771_),
    .A2(_02772_),
    .A3(_02773_),
    .S1(_02397_),
    .X(_02775_));
 sg13g2_nor2_1 _07888_ (.A(_02395_),
    .B(_02775_),
    .Y(_02776_));
 sg13g2_a21oi_2 _07889_ (.B1(_02776_),
    .Y(_02777_),
    .A2(_02769_),
    .A1(_02395_));
 sg13g2_nand2_1 _07890_ (.Y(_02778_),
    .A(net254),
    .B(_02777_));
 sg13g2_o21ai_1 _07891_ (.B1(_02778_),
    .Y(_02779_),
    .A1(net254),
    .A2(_02768_));
 sg13g2_a22oi_1 _07892_ (.Y(_02780_),
    .B1(_02779_),
    .B2(_02407_),
    .A2(_02767_),
    .A1(net114));
 sg13g2_nor3_1 _07893_ (.A(_02307_),
    .B(_02425_),
    .C(_02427_),
    .Y(_02781_));
 sg13g2_xnor2_1 _07894_ (.Y(_02782_),
    .A(_00189_),
    .B(_02781_));
 sg13g2_a221oi_1 _07895_ (.B2(_02417_),
    .C1(_02492_),
    .B1(_02782_),
    .A1(_02332_),
    .Y(_02783_),
    .A2(_02777_));
 sg13g2_nand2_1 _07896_ (.Y(_02784_),
    .A(_02780_),
    .B(_02783_));
 sg13g2_buf_1 _07897_ (.A(_00190_),
    .X(_02785_));
 sg13g2_nor2_1 _07898_ (.A(_02785_),
    .B(_02680_),
    .Y(_02786_));
 sg13g2_a21oi_1 _07899_ (.A1(_00189_),
    .A2(_02590_),
    .Y(_02787_),
    .B1(_02687_));
 sg13g2_o21ai_1 _07900_ (.B1(_02787_),
    .Y(_02788_),
    .A1(_02784_),
    .A2(_02786_));
 sg13g2_nand2_1 _07901_ (.Y(_02789_),
    .A(net125),
    .B(_02777_));
 sg13g2_nand2_1 _07902_ (.Y(_02790_),
    .A(_02788_),
    .B(_02789_));
 sg13g2_a22oi_1 _07903_ (.Y(_02791_),
    .B1(_02790_),
    .B2(_02288_),
    .A2(_02385_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sg13g2_nand2_1 _07904_ (.Y(_02792_),
    .A(net159),
    .B(_02791_));
 sg13g2_o21ai_1 _07905_ (.B1(_02792_),
    .Y(_02793_),
    .A1(\z80.tv80s.i_tv80_core.R[7] ),
    .A2(net159));
 sg13g2_nand2_1 _07906_ (.Y(_02794_),
    .A(\addr_bus[7] ),
    .B(_02551_));
 sg13g2_o21ai_1 _07907_ (.B1(_02794_),
    .Y(_00311_),
    .A1(_02245_),
    .A2(_02793_));
 sg13g2_mux4_1 _07908_ (.S0(net291),
    .A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .S1(net290),
    .X(_02795_));
 sg13g2_mux4_1 _07909_ (.S0(net330),
    .A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .S1(net290),
    .X(_02796_));
 sg13g2_mux2_1 _07910_ (.A0(_02795_),
    .A1(_02796_),
    .S(net331),
    .X(_02797_));
 sg13g2_inv_1 _07911_ (.Y(_02798_),
    .A(_02797_));
 sg13g2_a21oi_1 _07912_ (.A1(net127),
    .A2(_02798_),
    .Y(_02799_),
    .B1(net111));
 sg13g2_a21oi_1 _07913_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .A2(_02373_),
    .Y(_02800_),
    .B1(_02347_));
 sg13g2_and2_1 _07914_ (.A(_01605_),
    .B(net192),
    .X(_02801_));
 sg13g2_buf_1 _07915_ (.A(\z80.tv80s.i_tv80_core.PC[8] ),
    .X(_02802_));
 sg13g2_inv_1 _07916_ (.Y(_02803_),
    .A(net373));
 sg13g2_nand2_1 _07917_ (.Y(_02804_),
    .A(net332),
    .B(_00138_));
 sg13g2_nand2b_1 _07918_ (.Y(_02805_),
    .B(_00139_),
    .A_N(net352));
 sg13g2_nand3_1 _07919_ (.B(_02804_),
    .C(_02805_),
    .A(net247),
    .Y(_02806_));
 sg13g2_o21ai_1 _07920_ (.B1(_02806_),
    .Y(_02807_),
    .A1(net251),
    .A2(_02798_));
 sg13g2_xnor2_1 _07921_ (.Y(_02808_),
    .A(_00138_),
    .B(_02428_));
 sg13g2_nor2_1 _07922_ (.A(net137),
    .B(_02808_),
    .Y(_02809_));
 sg13g2_a21oi_1 _07923_ (.A1(_00137_),
    .A2(net128),
    .Y(_02810_),
    .B1(_02809_));
 sg13g2_a22oi_1 _07924_ (.Y(_02811_),
    .B1(_02810_),
    .B2(net96),
    .A2(_02807_),
    .A1(net97));
 sg13g2_buf_1 _07925_ (.A(\z80.tv80s.i_tv80_core.SP[8] ),
    .X(_02812_));
 sg13g2_mux2_1 _07926_ (.A0(_01545_),
    .A1(_02812_),
    .S(net145),
    .X(_02813_));
 sg13g2_a221oi_1 _07927_ (.B2(_02290_),
    .C1(net110),
    .B1(_02813_),
    .A1(_02331_),
    .Y(_02814_),
    .A2(_02797_));
 sg13g2_a221oi_1 _07928_ (.B2(_02814_),
    .C1(net193),
    .B1(_02811_),
    .A1(_02803_),
    .Y(_02815_),
    .A2(net112));
 sg13g2_o21ai_1 _07929_ (.B1(net84),
    .Y(_02816_),
    .A1(_02801_),
    .A2(_02815_));
 sg13g2_nand2_1 _07930_ (.Y(_02817_),
    .A(_02800_),
    .B(_02816_));
 sg13g2_a22oi_1 _07931_ (.Y(_02818_),
    .B1(_02799_),
    .B2(_02817_),
    .A2(net109),
    .A1(net350));
 sg13g2_nor2_1 _07932_ (.A(net164),
    .B(_02818_),
    .Y(_02819_));
 sg13g2_a21oi_1 _07933_ (.A1(_01605_),
    .A2(net165),
    .Y(_02820_),
    .B1(_02819_));
 sg13g2_nand2_1 _07934_ (.Y(_02821_),
    .A(\addr_bus[8] ),
    .B(net69));
 sg13g2_o21ai_1 _07935_ (.B1(_02821_),
    .Y(_00312_),
    .A1(net71),
    .A2(_02820_));
 sg13g2_mux4_1 _07936_ (.S0(net291),
    .A0(_00043_),
    .A1(_00045_),
    .A2(_00044_),
    .A3(_00046_),
    .S1(net290),
    .X(_02822_));
 sg13g2_mux4_1 _07937_ (.S0(net330),
    .A0(_00039_),
    .A1(_00041_),
    .A2(_00040_),
    .A3(_00042_),
    .S1(net329),
    .X(_02823_));
 sg13g2_nor2b_1 _07938_ (.A(net331),
    .B_N(_02823_),
    .Y(_02824_));
 sg13g2_a21oi_1 _07939_ (.A1(net292),
    .A2(_02822_),
    .Y(_02825_),
    .B1(_02824_));
 sg13g2_buf_1 _07940_ (.A(_02825_),
    .X(_02826_));
 sg13g2_o21ai_1 _07941_ (.B1(_02287_),
    .Y(_02827_),
    .A1(net136),
    .A2(_02826_));
 sg13g2_buf_2 _07942_ (.A(_00140_),
    .X(_02828_));
 sg13g2_nand2_1 _07943_ (.Y(_02829_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .B(_02428_));
 sg13g2_xor2_1 _07944_ (.B(_02829_),
    .A(_00141_),
    .X(_02830_));
 sg13g2_nor2_1 _07945_ (.A(net128),
    .B(_02830_),
    .Y(_02831_));
 sg13g2_a21oi_1 _07946_ (.A1(_02828_),
    .A2(_02308_),
    .Y(_02832_),
    .B1(_02831_));
 sg13g2_inv_1 _07947_ (.Y(_02833_),
    .A(_00142_));
 sg13g2_nand2_1 _07948_ (.Y(_02834_),
    .A(net293),
    .B(_00141_));
 sg13g2_o21ai_1 _07949_ (.B1(_02834_),
    .Y(_02835_),
    .A1(net293),
    .A2(_02833_));
 sg13g2_nand2_1 _07950_ (.Y(_02836_),
    .A(net254),
    .B(_02826_));
 sg13g2_o21ai_1 _07951_ (.B1(_02836_),
    .Y(_02837_),
    .A1(net254),
    .A2(_02835_));
 sg13g2_a22oi_1 _07952_ (.Y(_02838_),
    .B1(_02837_),
    .B2(net97),
    .A2(_02832_),
    .A1(net96));
 sg13g2_buf_1 _07953_ (.A(\z80.tv80s.i_tv80_core.PC[9] ),
    .X(_02839_));
 sg13g2_a221oi_1 _07954_ (.B2(net113),
    .C1(net193),
    .B1(_02826_),
    .A1(net372),
    .Y(_02840_),
    .A2(_02336_));
 sg13g2_buf_1 _07955_ (.A(\z80.tv80s.i_tv80_core.SP[9] ),
    .X(_02841_));
 sg13g2_mux2_1 _07956_ (.A0(_01683_),
    .A1(_02841_),
    .S(_02293_),
    .X(_02842_));
 sg13g2_nand2_1 _07957_ (.Y(_02843_),
    .A(_02291_),
    .B(_02842_));
 sg13g2_nand3_1 _07958_ (.B(_02840_),
    .C(_02843_),
    .A(_02838_),
    .Y(_02844_));
 sg13g2_a21oi_1 _07959_ (.A1(_01687_),
    .A2(net174),
    .Y(_02845_),
    .B1(_02375_));
 sg13g2_a221oi_1 _07960_ (.B2(_02845_),
    .C1(net126),
    .B1(_02844_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .Y(_02846_),
    .A2(_02444_));
 sg13g2_nand2_1 _07961_ (.Y(_02847_),
    .A(net390),
    .B(_02392_));
 sg13g2_o21ai_1 _07962_ (.B1(_02847_),
    .Y(_02848_),
    .A1(_02827_),
    .A2(_02846_));
 sg13g2_mux2_1 _07963_ (.A0(\z80.tv80s.i_tv80_core.I[1] ),
    .A1(_02848_),
    .S(_02246_),
    .X(_02849_));
 sg13g2_mux2_1 _07964_ (.A0(_02849_),
    .A1(\addr_bus[9] ),
    .S(_02389_),
    .X(_00313_));
 sg13g2_buf_2 _07965_ (.A(_00020_),
    .X(_02850_));
 sg13g2_nand2_1 _07966_ (.Y(_02851_),
    .A(_01346_),
    .B(_01573_));
 sg13g2_nor4_1 _07967_ (.A(_00802_),
    .B(_01420_),
    .C(_02267_),
    .D(_02851_),
    .Y(_02852_));
 sg13g2_mux2_1 _07968_ (.A0(\z80.tv80s.i_tv80_core.Alternate ),
    .A1(_02850_),
    .S(_02852_),
    .X(_00314_));
 sg13g2_nand3_1 _07969_ (.B(_01548_),
    .C(_01573_),
    .A(_01346_),
    .Y(_02853_));
 sg13g2_buf_1 _07970_ (.A(_02853_),
    .X(_02854_));
 sg13g2_buf_1 _07971_ (.A(_02854_),
    .X(_02855_));
 sg13g2_buf_1 _07972_ (.A(_02854_),
    .X(_02856_));
 sg13g2_nand2_1 _07973_ (.Y(_02857_),
    .A(_00229_),
    .B(net123));
 sg13g2_o21ai_1 _07974_ (.B1(_02857_),
    .Y(_00315_),
    .A1(_01545_),
    .A2(net124));
 sg13g2_nand2_1 _07975_ (.Y(_02858_),
    .A(_00230_),
    .B(net123));
 sg13g2_o21ai_1 _07976_ (.B1(_02858_),
    .Y(_00316_),
    .A1(_01683_),
    .A2(net124));
 sg13g2_nand2_1 _07977_ (.Y(_02859_),
    .A(_00231_),
    .B(net123));
 sg13g2_o21ai_1 _07978_ (.B1(_02859_),
    .Y(_00317_),
    .A1(_01736_),
    .A2(net124));
 sg13g2_nand2_1 _07979_ (.Y(_02860_),
    .A(_00232_),
    .B(_02856_));
 sg13g2_o21ai_1 _07980_ (.B1(_02860_),
    .Y(_00318_),
    .A1(net379),
    .A2(net124));
 sg13g2_buf_1 _07981_ (.A(_02854_),
    .X(_02861_));
 sg13g2_nand2_1 _07982_ (.Y(_02862_),
    .A(_00233_),
    .B(net122));
 sg13g2_o21ai_1 _07983_ (.B1(_02862_),
    .Y(_00319_),
    .A1(_01864_),
    .A2(net124));
 sg13g2_nand2_1 _07984_ (.Y(_02863_),
    .A(_00234_),
    .B(net122));
 sg13g2_o21ai_1 _07985_ (.B1(_02863_),
    .Y(_00320_),
    .A1(net375),
    .A2(net124));
 sg13g2_nand2_1 _07986_ (.Y(_02864_),
    .A(_00235_),
    .B(_02861_));
 sg13g2_o21ai_1 _07987_ (.B1(_02864_),
    .Y(_00321_),
    .A1(_02007_),
    .A2(_02855_));
 sg13g2_nand2_1 _07988_ (.Y(_02865_),
    .A(_00236_),
    .B(_02861_));
 sg13g2_o21ai_1 _07989_ (.B1(_02865_),
    .Y(_00322_),
    .A1(_02076_),
    .A2(_02855_));
 sg13g2_nand2_1 _07990_ (.Y(_02866_),
    .A(net219),
    .B(_01431_));
 sg13g2_nor3_1 _07991_ (.A(net242),
    .B(_00735_),
    .C(_01421_),
    .Y(_02867_));
 sg13g2_nand3_1 _07992_ (.B(_01423_),
    .C(_01428_),
    .A(_02867_),
    .Y(_02868_));
 sg13g2_buf_1 _07993_ (.A(_02868_),
    .X(_02869_));
 sg13g2_nor2_1 _07994_ (.A(_02866_),
    .B(_02869_),
    .Y(_02870_));
 sg13g2_nand3_1 _07995_ (.B(_02364_),
    .C(_02870_),
    .A(_02115_),
    .Y(_02871_));
 sg13g2_buf_1 _07996_ (.A(\z80.tv80s.i_tv80_core.Arith16_r ),
    .X(_02872_));
 sg13g2_nand2_1 _07997_ (.Y(_02873_),
    .A(_02872_),
    .B(_01747_));
 sg13g2_o21ai_1 _07998_ (.B1(_02873_),
    .Y(_00323_),
    .A1(_01239_),
    .A2(_02871_));
 sg13g2_nand2_1 _07999_ (.Y(_02874_),
    .A(net201),
    .B(_00922_));
 sg13g2_nand2_1 _08000_ (.Y(_02875_),
    .A(net214),
    .B(_01354_));
 sg13g2_o21ai_1 _08001_ (.B1(_02875_),
    .Y(_02876_),
    .A1(net214),
    .A2(net228));
 sg13g2_nor2_1 _08002_ (.A(_00984_),
    .B(net228),
    .Y(_02877_));
 sg13g2_nor2_2 _08003_ (.A(net229),
    .B(_00986_),
    .Y(_02878_));
 sg13g2_a22oi_1 _08004_ (.Y(_02879_),
    .B1(_02877_),
    .B2(_02878_),
    .A2(_02876_),
    .A1(_01120_));
 sg13g2_nor3_1 _08005_ (.A(_00769_),
    .B(_02299_),
    .C(_02303_),
    .Y(_02880_));
 sg13g2_nor3_1 _08006_ (.A(_02357_),
    .B(_01416_),
    .C(_02301_),
    .Y(_02881_));
 sg13g2_nor2_1 _08007_ (.A(_00802_),
    .B(_00833_),
    .Y(_02882_));
 sg13g2_and4_1 _08008_ (.A(_01081_),
    .B(_02880_),
    .C(_02881_),
    .D(_02882_),
    .X(_02883_));
 sg13g2_nand4_1 _08009_ (.B(net241),
    .C(_00720_),
    .A(net301),
    .Y(_02884_),
    .D(_02883_));
 sg13g2_o21ai_1 _08010_ (.B1(_02884_),
    .Y(_02885_),
    .A1(net266),
    .A2(_02879_));
 sg13g2_buf_1 _08011_ (.A(_02885_),
    .X(_02886_));
 sg13g2_nand2b_1 _08012_ (.Y(_02887_),
    .B(_02886_),
    .A_N(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ));
 sg13g2_a21oi_1 _08013_ (.A1(_02874_),
    .A2(_02887_),
    .Y(_02888_),
    .B1(net100));
 sg13g2_buf_1 _08014_ (.A(net399),
    .X(_02889_));
 sg13g2_mux2_1 _08015_ (.A0(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ),
    .A1(_02888_),
    .S(net328),
    .X(_00324_));
 sg13g2_nor2_1 _08016_ (.A(_00209_),
    .B(net100),
    .Y(_02890_));
 sg13g2_mux2_1 _08017_ (.A0(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ),
    .A1(_02890_),
    .S(net328),
    .X(_00325_));
 sg13g2_buf_1 _08018_ (.A(\z80.tv80s.i_tv80_core.BTR_r ),
    .X(_02891_));
 sg13g2_nor4_1 _08019_ (.A(\z80.tv80s.i_tv80_core.No_BTR ),
    .B(net182),
    .C(_02142_),
    .D(_02248_),
    .Y(_02892_));
 sg13g2_a21o_1 _08020_ (.A2(_02142_),
    .A1(_02891_),
    .B1(_02892_),
    .X(_00326_));
 sg13g2_a21oi_1 _08021_ (.A1(_00851_),
    .A2(_00028_),
    .Y(_02893_),
    .B1(_01368_));
 sg13g2_nand3_1 _08022_ (.B(net204),
    .C(_02893_),
    .A(_01071_),
    .Y(_02894_));
 sg13g2_buf_1 _08023_ (.A(_02894_),
    .X(_02895_));
 sg13g2_nor2_1 _08024_ (.A(net230),
    .B(_02895_),
    .Y(_02896_));
 sg13g2_nor2_1 _08025_ (.A(_02104_),
    .B(_02896_),
    .Y(_02897_));
 sg13g2_and2_1 _08026_ (.A(_01077_),
    .B(_01554_),
    .X(_02898_));
 sg13g2_buf_1 _08027_ (.A(_02898_),
    .X(_02899_));
 sg13g2_a21oi_1 _08028_ (.A1(_01054_),
    .A2(_01185_),
    .Y(_02900_),
    .B1(_02899_));
 sg13g2_nor2_1 _08029_ (.A(net230),
    .B(_01151_),
    .Y(_02901_));
 sg13g2_nand2_1 _08030_ (.Y(_02902_),
    .A(_01558_),
    .B(_02259_));
 sg13g2_nand3_1 _08031_ (.B(_01362_),
    .C(_01444_),
    .A(_01434_),
    .Y(_02903_));
 sg13g2_a21oi_1 _08032_ (.A1(net240),
    .A2(_01550_),
    .Y(_02904_),
    .B1(net234));
 sg13g2_nor3_1 _08033_ (.A(_02902_),
    .B(_02903_),
    .C(_02904_),
    .Y(_02905_));
 sg13g2_nand4_1 _08034_ (.B(_02900_),
    .C(_02901_),
    .A(_02870_),
    .Y(_02906_),
    .D(_02905_));
 sg13g2_nor4_1 _08035_ (.A(_00802_),
    .B(_01420_),
    .C(_01547_),
    .D(_02906_),
    .Y(_02907_));
 sg13g2_nor2_1 _08036_ (.A(net285),
    .B(_00796_),
    .Y(_02908_));
 sg13g2_nand2_1 _08037_ (.Y(_02909_),
    .A(net245),
    .B(_02908_));
 sg13g2_nor4_1 _08038_ (.A(_00961_),
    .B(net351),
    .C(_02909_),
    .D(net230),
    .Y(_02910_));
 sg13g2_o21ai_1 _08039_ (.B1(net301),
    .Y(_02911_),
    .A1(_02907_),
    .A2(_02910_));
 sg13g2_o21ai_1 _08040_ (.B1(_02911_),
    .Y(_02912_),
    .A1(_01229_),
    .A2(_02897_));
 sg13g2_buf_1 _08041_ (.A(_02912_),
    .X(_02913_));
 sg13g2_a21oi_1 _08042_ (.A1(_00951_),
    .A2(_01371_),
    .Y(_02914_),
    .B1(_00933_));
 sg13g2_nor2_1 _08043_ (.A(_01289_),
    .B(_02914_),
    .Y(_02915_));
 sg13g2_nor2_1 _08044_ (.A(_01062_),
    .B(_00831_),
    .Y(_02916_));
 sg13g2_nor2b_1 _08045_ (.A(_02277_),
    .B_N(_02916_),
    .Y(_02917_));
 sg13g2_a22oi_1 _08046_ (.Y(_02918_),
    .B1(_02917_),
    .B2(_00977_),
    .A2(_02915_),
    .A1(_00721_));
 sg13g2_nor2_1 _08047_ (.A(net351),
    .B(net267),
    .Y(_02919_));
 sg13g2_a221oi_1 _08048_ (.B2(net203),
    .C1(_02122_),
    .B1(_02919_),
    .A1(net209),
    .Y(_02920_),
    .A2(net219));
 sg13g2_nor2_1 _08049_ (.A(_01388_),
    .B(_01005_),
    .Y(_02921_));
 sg13g2_nand2_1 _08050_ (.Y(_02922_),
    .A(net175),
    .B(net228));
 sg13g2_nand2_1 _08051_ (.Y(_02923_),
    .A(_00821_),
    .B(_00850_));
 sg13g2_a21oi_1 _08052_ (.A1(_00923_),
    .A2(_02923_),
    .Y(_02924_),
    .B1(_00639_));
 sg13g2_and2_1 _08053_ (.A(net205),
    .B(_02924_),
    .X(_02925_));
 sg13g2_buf_1 _08054_ (.A(_02925_),
    .X(_02926_));
 sg13g2_a221oi_1 _08055_ (.B2(_01117_),
    .C1(_02926_),
    .B1(_02922_),
    .A1(_02899_),
    .Y(_02927_),
    .A2(_02921_));
 sg13g2_or3_1 _08056_ (.A(_01052_),
    .B(_01061_),
    .C(_01082_),
    .X(_02928_));
 sg13g2_buf_1 _08057_ (.A(_02928_),
    .X(_02929_));
 sg13g2_a21oi_1 _08058_ (.A1(net306),
    .A2(_02133_),
    .Y(_02930_),
    .B1(_02929_));
 sg13g2_nand2_1 _08059_ (.Y(_02931_),
    .A(net258),
    .B(_00797_));
 sg13g2_buf_1 _08060_ (.A(_02931_),
    .X(_02932_));
 sg13g2_nand2_1 _08061_ (.Y(_02933_),
    .A(_01352_),
    .B(net200));
 sg13g2_o21ai_1 _08062_ (.B1(_02933_),
    .Y(_02934_),
    .A1(net257),
    .A2(_02932_));
 sg13g2_nor3_1 _08063_ (.A(net270),
    .B(_00971_),
    .C(_02932_),
    .Y(_02935_));
 sg13g2_a221oi_1 _08064_ (.B2(net235),
    .C1(_02935_),
    .B1(_02934_),
    .A1(_00933_),
    .Y(_02936_),
    .A2(_02930_));
 sg13g2_nand2b_1 _08065_ (.Y(_02937_),
    .B(net223),
    .A_N(_02936_));
 sg13g2_nand4_1 _08066_ (.B(_02920_),
    .C(_02927_),
    .A(_02918_),
    .Y(_02938_),
    .D(_02937_));
 sg13g2_or2_1 _08067_ (.X(_02939_),
    .B(_01248_),
    .A(_00871_));
 sg13g2_a21oi_1 _08068_ (.A1(net301),
    .A2(_02938_),
    .Y(_02940_),
    .B1(_02939_));
 sg13g2_nor2_1 _08069_ (.A(net272),
    .B(net351),
    .Y(_02941_));
 sg13g2_nand3_1 _08070_ (.B(_00815_),
    .C(_02941_),
    .A(_01111_),
    .Y(_02942_));
 sg13g2_inv_1 _08071_ (.Y(_02943_),
    .A(_02942_));
 sg13g2_nand2_1 _08072_ (.Y(_02944_),
    .A(_00933_),
    .B(_02943_));
 sg13g2_o21ai_1 _08073_ (.B1(_02944_),
    .Y(_02945_),
    .A1(net257),
    .A2(_02895_));
 sg13g2_a221oi_1 _08074_ (.B2(_01191_),
    .C1(net266),
    .B1(_01371_),
    .A1(net241),
    .Y(_02946_),
    .A2(_00885_));
 sg13g2_inv_1 _08075_ (.Y(_02947_),
    .A(_02946_));
 sg13g2_a221oi_1 _08076_ (.B2(_01259_),
    .C1(_02947_),
    .B1(_02945_),
    .A1(net170),
    .Y(_02948_),
    .A2(net219));
 sg13g2_or2_1 _08077_ (.X(_02949_),
    .B(_02948_),
    .A(_02940_));
 sg13g2_buf_1 _08078_ (.A(_02949_),
    .X(_02950_));
 sg13g2_nor2_1 _08079_ (.A(net217),
    .B(_01084_),
    .Y(_02951_));
 sg13g2_nor3_1 _08080_ (.A(net267),
    .B(_02929_),
    .C(_02951_),
    .Y(_02952_));
 sg13g2_o21ai_1 _08081_ (.B1(net270),
    .Y(_02953_),
    .A1(_01241_),
    .A2(_02952_));
 sg13g2_o21ai_1 _08082_ (.B1(_02953_),
    .Y(_02954_),
    .A1(net184),
    .A2(_01380_));
 sg13g2_nor2_1 _08083_ (.A(_02277_),
    .B(_02932_),
    .Y(_02955_));
 sg13g2_o21ai_1 _08084_ (.B1(_01331_),
    .Y(_02956_),
    .A1(_02954_),
    .A2(_02955_));
 sg13g2_mux2_1 _08085_ (.A0(_02919_),
    .A1(_02922_),
    .S(_00978_),
    .X(_02957_));
 sg13g2_a21oi_1 _08086_ (.A1(net310),
    .A2(_02957_),
    .Y(_02958_),
    .B1(_02122_));
 sg13g2_nand2_1 _08087_ (.Y(_02959_),
    .A(_01410_),
    .B(_02917_));
 sg13g2_nand2_1 _08088_ (.Y(_02960_),
    .A(_00935_),
    .B(_01172_));
 sg13g2_nand2_1 _08089_ (.Y(_02961_),
    .A(_02177_),
    .B(_01290_));
 sg13g2_nand3_1 _08090_ (.B(_02960_),
    .C(_02961_),
    .A(net208),
    .Y(_02962_));
 sg13g2_nand4_1 _08091_ (.B(_02958_),
    .C(_02959_),
    .A(_02956_),
    .Y(_02963_),
    .D(_02962_));
 sg13g2_a21o_1 _08092_ (.A2(net358),
    .A1(_00984_),
    .B1(_00871_),
    .X(_02964_));
 sg13g2_a21oi_1 _08093_ (.A1(net301),
    .A2(_02963_),
    .Y(_02965_),
    .B1(_02964_));
 sg13g2_nor2_1 _08094_ (.A(net184),
    .B(_02942_),
    .Y(_02966_));
 sg13g2_nor2_1 _08095_ (.A(_01259_),
    .B(_02895_),
    .Y(_02967_));
 sg13g2_o21ai_1 _08096_ (.B1(_01331_),
    .Y(_02968_),
    .A1(_02966_),
    .A2(_02967_));
 sg13g2_nand3b_1 _08097_ (.B(_02946_),
    .C(_02968_),
    .Y(_02969_),
    .A_N(_02104_));
 sg13g2_nand2b_1 _08098_ (.Y(_02970_),
    .B(_02969_),
    .A_N(_02965_));
 sg13g2_buf_1 _08099_ (.A(_02970_),
    .X(_02971_));
 sg13g2_nand2_1 _08100_ (.Y(_02972_),
    .A(_02950_),
    .B(_02971_));
 sg13g2_a21o_1 _08101_ (.A2(_02972_),
    .A1(_02913_),
    .B1(_01266_),
    .X(_02973_));
 sg13g2_buf_2 _08102_ (.A(_02973_),
    .X(_02974_));
 sg13g2_nor3_1 _08103_ (.A(_02913_),
    .B(_02950_),
    .C(_02971_),
    .Y(_02975_));
 sg13g2_buf_2 _08104_ (.A(_02975_),
    .X(_02976_));
 sg13g2_xnor2_1 _08105_ (.Y(_02977_),
    .A(_00850_),
    .B(net199));
 sg13g2_a22oi_1 _08106_ (.Y(_02978_),
    .B1(_02943_),
    .B2(net176),
    .A2(net170),
    .A1(net235));
 sg13g2_o21ai_1 _08107_ (.B1(_02978_),
    .Y(_02979_),
    .A1(_02895_),
    .A2(_02977_));
 sg13g2_nand2_1 _08108_ (.Y(_02980_),
    .A(_00845_),
    .B(_02932_));
 sg13g2_nand2_1 _08109_ (.Y(_02981_),
    .A(_01077_),
    .B(_01554_));
 sg13g2_nand3_1 _08110_ (.B(net199),
    .C(_02916_),
    .A(net357),
    .Y(_02982_));
 sg13g2_o21ai_1 _08111_ (.B1(_02982_),
    .Y(_02983_),
    .A1(_02981_),
    .A2(_02923_));
 sg13g2_a22oi_1 _08112_ (.Y(_02984_),
    .B1(net230),
    .B2(_02916_),
    .A2(_01352_),
    .A1(net195));
 sg13g2_nand2_1 _08113_ (.Y(_02985_),
    .A(_00970_),
    .B(_02984_));
 sg13g2_o21ai_1 _08114_ (.B1(_02985_),
    .Y(_02986_),
    .A1(net235),
    .A2(_02983_));
 sg13g2_nand2_1 _08115_ (.Y(_02987_),
    .A(_00891_),
    .B(net199));
 sg13g2_inv_1 _08116_ (.Y(_02988_),
    .A(_02092_));
 sg13g2_nand3_1 _08117_ (.B(_00719_),
    .C(net200),
    .A(_02988_),
    .Y(_02989_));
 sg13g2_o21ai_1 _08118_ (.B1(_02989_),
    .Y(_02990_),
    .A1(_02932_),
    .A2(_02987_));
 sg13g2_a21oi_1 _08119_ (.A1(net205),
    .A2(_01371_),
    .Y(_02991_),
    .B1(_02990_));
 sg13g2_nand3_1 _08120_ (.B(_02986_),
    .C(_02991_),
    .A(_02958_),
    .Y(_02992_));
 sg13g2_a221oi_1 _08121_ (.B2(_01296_),
    .C1(_02992_),
    .B1(_02980_),
    .A1(net176),
    .Y(_02993_),
    .A2(_02930_));
 sg13g2_a21oi_1 _08122_ (.A1(net214),
    .A2(_00863_),
    .Y(_02994_),
    .B1(net276));
 sg13g2_o21ai_1 _08123_ (.B1(_02994_),
    .Y(_02995_),
    .A1(net305),
    .A2(_02993_));
 sg13g2_o21ai_1 _08124_ (.B1(_02995_),
    .Y(_02996_),
    .A1(_02947_),
    .A2(_02979_));
 sg13g2_buf_1 _08125_ (.A(_02996_),
    .X(_02997_));
 sg13g2_buf_1 _08126_ (.A(_02997_),
    .X(_02998_));
 sg13g2_mux2_1 _08127_ (.A0(_01545_),
    .A1(net350),
    .S(net108),
    .X(_02999_));
 sg13g2_inv_1 _08128_ (.Y(_03000_),
    .A(_02913_));
 sg13g2_nor2_1 _08129_ (.A(_03000_),
    .B(_02972_),
    .Y(_03001_));
 sg13g2_buf_2 _08130_ (.A(_03001_),
    .X(_03002_));
 sg13g2_mux2_1 _08131_ (.A0(_02812_),
    .A1(_02294_),
    .S(net108),
    .X(_03003_));
 sg13g2_o21ai_1 _08132_ (.B1(_03000_),
    .Y(_03004_),
    .A1(_02950_),
    .A2(_02971_));
 sg13g2_buf_2 _08133_ (.A(_03004_),
    .X(_03005_));
 sg13g2_buf_1 _08134_ (.A(_02997_),
    .X(_03006_));
 sg13g2_buf_1 _08135_ (.A(_03006_),
    .X(_03007_));
 sg13g2_nand2_1 _08136_ (.Y(_03008_),
    .A(_00870_),
    .B(_01377_));
 sg13g2_a21oi_2 _08137_ (.B1(_03008_),
    .Y(_03009_),
    .A2(_01128_),
    .A1(_01166_));
 sg13g2_nor2b_1 _08138_ (.A(_01360_),
    .B_N(_00849_),
    .Y(_03010_));
 sg13g2_buf_1 _08139_ (.A(_03010_),
    .X(_03011_));
 sg13g2_nor2b_1 _08140_ (.A(net394),
    .B_N(_02276_),
    .Y(_03012_));
 sg13g2_nor2_1 _08141_ (.A(_01115_),
    .B(_03012_),
    .Y(_03013_));
 sg13g2_a22oi_1 _08142_ (.Y(_03014_),
    .B1(_03013_),
    .B2(_00833_),
    .A2(_01376_),
    .A1(_01156_));
 sg13g2_nor2_1 _08143_ (.A(_00023_),
    .B(net395),
    .Y(_03015_));
 sg13g2_a22oi_1 _08144_ (.Y(_03016_),
    .B1(_01283_),
    .B2(_03015_),
    .A2(_01184_),
    .A1(_00847_));
 sg13g2_nand2_2 _08145_ (.Y(_03017_),
    .A(_03014_),
    .B(_03016_));
 sg13g2_inv_1 _08146_ (.Y(_03018_),
    .A(_01377_));
 sg13g2_a21oi_1 _08147_ (.A1(_02909_),
    .A2(_02254_),
    .Y(_03019_),
    .B1(_03018_));
 sg13g2_nor2_1 _08148_ (.A(_02177_),
    .B(_01585_),
    .Y(_03020_));
 sg13g2_nor4_1 _08149_ (.A(_00928_),
    .B(_03017_),
    .C(_03019_),
    .D(_03020_),
    .Y(_03021_));
 sg13g2_a221oi_1 _08150_ (.B2(_00913_),
    .C1(net355),
    .B1(_03021_),
    .A1(_00940_),
    .Y(_03022_),
    .A2(_03011_));
 sg13g2_nor2_2 _08151_ (.A(_03009_),
    .B(_03022_),
    .Y(_03023_));
 sg13g2_nor4_1 _08152_ (.A(_00732_),
    .B(_00928_),
    .C(_03017_),
    .D(_03019_),
    .Y(_03024_));
 sg13g2_a221oi_1 _08153_ (.B2(_00940_),
    .C1(net355),
    .B1(_03011_),
    .A1(_00913_),
    .Y(_03025_),
    .A2(_03024_));
 sg13g2_buf_2 _08154_ (.A(_03025_),
    .X(_03026_));
 sg13g2_a22oi_1 _08155_ (.Y(_03027_),
    .B1(_01171_),
    .B2(net283),
    .A2(_00877_),
    .A1(net360));
 sg13g2_a21oi_1 _08156_ (.A1(net207),
    .A2(_03027_),
    .Y(_03028_),
    .B1(_01121_));
 sg13g2_nor2_1 _08157_ (.A(_03008_),
    .B(_03028_),
    .Y(_03029_));
 sg13g2_buf_2 _08158_ (.A(_03029_),
    .X(_03030_));
 sg13g2_a21o_1 _08159_ (.A2(_03026_),
    .A1(net317),
    .B1(_03030_),
    .X(_03031_));
 sg13g2_buf_8 _08160_ (.A(_03031_),
    .X(_03032_));
 sg13g2_inv_1 _08161_ (.Y(_03033_),
    .A(_01307_));
 sg13g2_and4_1 _08162_ (.A(_03033_),
    .B(_01418_),
    .C(_01571_),
    .D(_02362_),
    .X(_03034_));
 sg13g2_buf_1 _08163_ (.A(_03034_),
    .X(_03035_));
 sg13g2_and2_1 _08164_ (.A(_01566_),
    .B(_03035_),
    .X(_03036_));
 sg13g2_buf_1 _08165_ (.A(_03036_),
    .X(_03037_));
 sg13g2_buf_8 _08166_ (.A(_03037_),
    .X(_03038_));
 sg13g2_and4_1 _08167_ (.A(net393),
    .B(_01418_),
    .C(_01571_),
    .D(_02362_),
    .X(_03039_));
 sg13g2_buf_1 _08168_ (.A(_03039_),
    .X(_03040_));
 sg13g2_buf_1 _08169_ (.A(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ),
    .X(_03041_));
 sg13g2_a21oi_1 _08170_ (.A1(_01566_),
    .A2(_03040_),
    .Y(_03042_),
    .B1(_03041_));
 sg13g2_o21ai_1 _08171_ (.B1(net304),
    .Y(_03043_),
    .A1(net144),
    .A2(_03042_));
 sg13g2_a21o_1 _08172_ (.A2(_03032_),
    .A1(_03023_),
    .B1(_03043_),
    .X(_03044_));
 sg13g2_buf_8 _08173_ (.A(_03044_),
    .X(_03045_));
 sg13g2_inv_1 _08174_ (.Y(_03046_),
    .A(\z80.tv80s.i_tv80_core.ts[3] ));
 sg13g2_nor2_1 _08175_ (.A(_00881_),
    .B(_03046_),
    .Y(_03047_));
 sg13g2_nand2_1 _08176_ (.Y(_03048_),
    .A(_00859_),
    .B(_03047_));
 sg13g2_a221oi_1 _08177_ (.B2(_00940_),
    .C1(_03048_),
    .B1(_03011_),
    .A1(_00913_),
    .Y(_03049_),
    .A2(_03024_));
 sg13g2_buf_2 _08178_ (.A(_03049_),
    .X(_03050_));
 sg13g2_nand2_1 _08179_ (.Y(_03051_),
    .A(net243),
    .B(net395));
 sg13g2_a21oi_1 _08180_ (.A1(_01115_),
    .A2(_03051_),
    .Y(_03052_),
    .B1(net281));
 sg13g2_nor2_1 _08181_ (.A(net243),
    .B(_01171_),
    .Y(_03053_));
 sg13g2_o21ai_1 _08182_ (.B1(net207),
    .Y(_03054_),
    .A1(_03052_),
    .A2(_03053_));
 sg13g2_nand2_1 _08183_ (.Y(_03055_),
    .A(_00870_),
    .B(_03047_));
 sg13g2_o21ai_1 _08184_ (.B1(_00032_),
    .Y(_03056_),
    .A1(_03054_),
    .A2(_03055_));
 sg13g2_buf_1 _08185_ (.A(_03056_),
    .X(_03057_));
 sg13g2_and2_1 _08186_ (.A(_02311_),
    .B(_03057_),
    .X(_03058_));
 sg13g2_a21o_1 _08187_ (.A2(_03050_),
    .A1(_02311_),
    .B1(_03058_),
    .X(_03059_));
 sg13g2_buf_8 _08188_ (.A(_03059_),
    .X(_03060_));
 sg13g2_or2_1 _08189_ (.X(_03061_),
    .B(_03042_),
    .A(_03037_));
 sg13g2_nor2_1 _08190_ (.A(_03057_),
    .B(_03050_),
    .Y(_03062_));
 sg13g2_a22oi_1 _08191_ (.Y(_03063_),
    .B1(_03061_),
    .B2(_03062_),
    .A2(_03023_),
    .A1(_03060_));
 sg13g2_buf_8 _08192_ (.A(_03063_),
    .X(_03064_));
 sg13g2_nand2_2 _08193_ (.Y(_03065_),
    .A(_03045_),
    .B(_03064_));
 sg13g2_buf_16 _08194_ (.X(_03066_),
    .A(_03065_));
 sg13g2_buf_8 _08195_ (.A(_03066_),
    .X(_03067_));
 sg13g2_buf_8 _08196_ (.A(net68),
    .X(_03068_));
 sg13g2_nor3_1 _08197_ (.A(_00928_),
    .B(_03017_),
    .C(_03019_),
    .Y(_03069_));
 sg13g2_nor2_1 _08198_ (.A(_03009_),
    .B(_03020_),
    .Y(_03070_));
 sg13g2_and3_1 _08199_ (.X(_03071_),
    .A(_00913_),
    .B(_03069_),
    .C(_03070_));
 sg13g2_buf_1 _08200_ (.A(_03071_),
    .X(_03072_));
 sg13g2_nor2_1 _08201_ (.A(_00859_),
    .B(_03009_),
    .Y(_03073_));
 sg13g2_a21o_1 _08202_ (.A2(_03011_),
    .A1(_00940_),
    .B1(_03073_),
    .X(_03074_));
 sg13g2_buf_1 _08203_ (.A(_03074_),
    .X(_03075_));
 sg13g2_nor2_2 _08204_ (.A(_03072_),
    .B(_03075_),
    .Y(_03076_));
 sg13g2_a21oi_2 _08205_ (.B1(_03030_),
    .Y(_03077_),
    .A2(_03026_),
    .A1(net317));
 sg13g2_inv_1 _08206_ (.Y(_03078_),
    .A(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ));
 sg13g2_a21oi_2 _08207_ (.B1(_03078_),
    .Y(_03079_),
    .A2(_03040_),
    .A1(net151));
 sg13g2_nor3_1 _08208_ (.A(_02311_),
    .B(_03079_),
    .C(net144),
    .Y(_03080_));
 sg13g2_o21ai_1 _08209_ (.B1(_03080_),
    .Y(_03081_),
    .A1(_03076_),
    .A2(_03077_));
 sg13g2_buf_1 _08210_ (.A(_03081_),
    .X(_03082_));
 sg13g2_nor2_1 _08211_ (.A(net396),
    .B(_01585_),
    .Y(_03083_));
 sg13g2_nor4_1 _08212_ (.A(_00928_),
    .B(_03017_),
    .C(_03019_),
    .D(_03083_),
    .Y(_03084_));
 sg13g2_a221oi_1 _08213_ (.B2(_00913_),
    .C1(net355),
    .B1(_03084_),
    .A1(_00940_),
    .Y(_03085_),
    .A2(_03011_));
 sg13g2_nor2_1 _08214_ (.A(_03030_),
    .B(_03085_),
    .Y(_03086_));
 sg13g2_nor2_1 _08215_ (.A(_03079_),
    .B(_03038_),
    .Y(_03087_));
 sg13g2_a22oi_1 _08216_ (.Y(_03088_),
    .B1(_03087_),
    .B2(_03062_),
    .A2(_03086_),
    .A1(_03060_));
 sg13g2_buf_1 _08217_ (.A(_03088_),
    .X(_03089_));
 sg13g2_and2_1 _08218_ (.A(_03082_),
    .B(_03089_),
    .X(_03090_));
 sg13g2_buf_2 _08219_ (.A(_03090_),
    .X(_03091_));
 sg13g2_buf_8 _08220_ (.A(_03091_),
    .X(_03092_));
 sg13g2_mux4_1 _08221_ (.S0(_03068_),
    .A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .S1(net67),
    .X(_03093_));
 sg13g2_mux4_1 _08222_ (.S0(net60),
    .A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .S1(_03091_),
    .X(_03094_));
 sg13g2_inv_1 _08223_ (.Y(_03095_),
    .A(_00037_));
 sg13g2_o21ai_1 _08224_ (.B1(net304),
    .Y(_03096_),
    .A1(_03057_),
    .A2(_03050_));
 sg13g2_or4_1 _08225_ (.A(_03095_),
    .B(_03076_),
    .C(_03077_),
    .D(_03096_),
    .X(_03097_));
 sg13g2_nand2b_1 _08226_ (.Y(_03098_),
    .B(_01307_),
    .A_N(net393));
 sg13g2_and4_1 _08227_ (.A(_01418_),
    .B(_01571_),
    .C(_02362_),
    .D(_03098_),
    .X(_03099_));
 sg13g2_nand3_1 _08228_ (.B(net151),
    .C(_03099_),
    .A(_02850_),
    .Y(_03100_));
 sg13g2_or4_1 _08229_ (.A(_01433_),
    .B(_01553_),
    .C(_01559_),
    .D(_01565_),
    .X(_03101_));
 sg13g2_buf_1 _08230_ (.A(_03101_),
    .X(_03102_));
 sg13g2_nand4_1 _08231_ (.B(_01571_),
    .C(_02362_),
    .A(_01418_),
    .Y(_03103_),
    .D(_03098_));
 sg13g2_buf_1 _08232_ (.A(_03103_),
    .X(_03104_));
 sg13g2_o21ai_1 _08233_ (.B1(_00038_),
    .Y(_03105_),
    .A1(_03102_),
    .A2(_03104_));
 sg13g2_a21oi_1 _08234_ (.A1(_03100_),
    .A2(_03105_),
    .Y(_03106_),
    .B1(_02311_));
 sg13g2_o21ai_1 _08235_ (.B1(_03106_),
    .Y(_03107_),
    .A1(_03076_),
    .A2(_03077_));
 sg13g2_a221oi_1 _08236_ (.B2(_03105_),
    .C1(_03057_),
    .B1(_03100_),
    .A1(_03047_),
    .Y(_03108_),
    .A2(_03026_));
 sg13g2_a21oi_1 _08237_ (.A1(_02850_),
    .A2(_03060_),
    .Y(_03109_),
    .B1(_03108_));
 sg13g2_and3_1 _08238_ (.X(_03110_),
    .A(_03097_),
    .B(_03107_),
    .C(_03109_));
 sg13g2_buf_8 _08239_ (.A(_03110_),
    .X(_03111_));
 sg13g2_buf_8 _08240_ (.A(_03111_),
    .X(_03112_));
 sg13g2_buf_8 _08241_ (.A(_03112_),
    .X(_03113_));
 sg13g2_mux2_1 _08242_ (.A0(_03093_),
    .A1(_03094_),
    .S(net66),
    .X(_03114_));
 sg13g2_buf_2 _08243_ (.A(_03114_),
    .X(_03115_));
 sg13g2_nand3_1 _08244_ (.B(net83),
    .C(net68),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .Y(_03116_));
 sg13g2_nand3_1 _08245_ (.B(_03107_),
    .C(_03109_),
    .A(_03097_),
    .Y(_03117_));
 sg13g2_buf_2 _08246_ (.A(_03117_),
    .X(_03118_));
 sg13g2_and2_1 _08247_ (.A(_03045_),
    .B(_03064_),
    .X(_03119_));
 sg13g2_buf_8 _08248_ (.A(_03119_),
    .X(_03120_));
 sg13g2_nand3_1 _08249_ (.B(_03118_),
    .C(_03120_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .Y(_03121_));
 sg13g2_nand2_1 _08250_ (.Y(_03122_),
    .A(_03082_),
    .B(_03089_));
 sg13g2_buf_2 _08251_ (.A(_03122_),
    .X(_03123_));
 sg13g2_buf_8 _08252_ (.A(_03123_),
    .X(_03124_));
 sg13g2_a21oi_1 _08253_ (.A1(_03116_),
    .A2(_03121_),
    .Y(_03125_),
    .B1(net65));
 sg13g2_nand3_1 _08254_ (.B(_03091_),
    .C(net68),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .Y(_03126_));
 sg13g2_nor2_1 _08255_ (.A(_03041_),
    .B(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ),
    .Y(_03127_));
 sg13g2_o21ai_1 _08256_ (.B1(_03127_),
    .Y(_03128_),
    .A1(_03102_),
    .A2(_03104_));
 sg13g2_nand2b_1 _08257_ (.Y(_03129_),
    .B(_01033_),
    .A_N(_03128_));
 sg13g2_a21oi_2 _08258_ (.B1(_03129_),
    .Y(_03130_),
    .A2(_03032_),
    .A1(_03023_));
 sg13g2_o21ai_1 _08259_ (.B1(_02311_),
    .Y(_03131_),
    .A1(_03057_),
    .A2(_03050_));
 sg13g2_or4_1 _08260_ (.A(_03009_),
    .B(_03030_),
    .C(_03085_),
    .D(_03022_),
    .X(_03132_));
 sg13g2_or3_1 _08261_ (.A(_03057_),
    .B(_03050_),
    .C(_03128_),
    .X(_03133_));
 sg13g2_o21ai_1 _08262_ (.B1(_03133_),
    .Y(_03134_),
    .A1(_03131_),
    .A2(_03132_));
 sg13g2_buf_2 _08263_ (.A(_03134_),
    .X(_03135_));
 sg13g2_or2_1 _08264_ (.X(_03136_),
    .B(_03135_),
    .A(_03130_));
 sg13g2_buf_2 _08265_ (.A(_03136_),
    .X(_03137_));
 sg13g2_nand2_1 _08266_ (.Y(_03138_),
    .A(_03041_),
    .B(_03078_));
 sg13g2_nand2_1 _08267_ (.Y(_03139_),
    .A(net151),
    .B(_03040_));
 sg13g2_buf_1 _08268_ (.A(_03139_),
    .X(_03140_));
 sg13g2_nand2_1 _08269_ (.Y(_03141_),
    .A(net151),
    .B(_03035_));
 sg13g2_buf_1 _08270_ (.A(_03141_),
    .X(_03142_));
 sg13g2_nand2_1 _08271_ (.Y(_03143_),
    .A(_01033_),
    .B(_03142_));
 sg13g2_a221oi_1 _08272_ (.B2(_03140_),
    .C1(_03143_),
    .B1(_03138_),
    .A1(_03023_),
    .Y(_03144_),
    .A2(_03032_));
 sg13g2_buf_2 _08273_ (.A(_03144_),
    .X(_03145_));
 sg13g2_nor4_1 _08274_ (.A(_03030_),
    .B(_03085_),
    .C(_03072_),
    .D(_03075_),
    .Y(_03146_));
 sg13g2_a22oi_1 _08275_ (.Y(_03147_),
    .B1(net151),
    .B2(_03040_),
    .A2(_03078_),
    .A1(_03041_));
 sg13g2_nor4_1 _08276_ (.A(_03057_),
    .B(_03050_),
    .C(net144),
    .D(_03147_),
    .Y(_03148_));
 sg13g2_a21o_1 _08277_ (.A2(_03146_),
    .A1(_03060_),
    .B1(_03148_),
    .X(_03149_));
 sg13g2_buf_2 _08278_ (.A(_03149_),
    .X(_03150_));
 sg13g2_or2_1 _08279_ (.X(_03151_),
    .B(_03150_),
    .A(_03145_));
 sg13g2_buf_2 _08280_ (.A(_03151_),
    .X(_03152_));
 sg13g2_buf_8 _08281_ (.A(_03111_),
    .X(_03153_));
 sg13g2_a221oi_1 _08282_ (.B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ),
    .C1(net82),
    .B1(_03152_),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ),
    .Y(_03154_),
    .A2(_03137_));
 sg13g2_o21ai_1 _08283_ (.B1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .Y(_03155_),
    .A1(_03130_),
    .A2(_03135_));
 sg13g2_o21ai_1 _08284_ (.B1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .Y(_03156_),
    .A1(_03145_),
    .A2(_03150_));
 sg13g2_inv_1 _08285_ (.Y(_03157_),
    .A(_03041_));
 sg13g2_a21oi_1 _08286_ (.A1(net151),
    .A2(_03035_),
    .Y(_03158_),
    .B1(_03157_));
 sg13g2_a21oi_1 _08287_ (.A1(_03079_),
    .A2(_03158_),
    .Y(_03159_),
    .B1(_02311_));
 sg13g2_o21ai_1 _08288_ (.B1(_03159_),
    .Y(_03160_),
    .A1(_03076_),
    .A2(_03077_));
 sg13g2_buf_2 _08289_ (.A(_03160_),
    .X(_03161_));
 sg13g2_nor2_1 _08290_ (.A(_03030_),
    .B(_03083_),
    .Y(_03162_));
 sg13g2_and3_1 _08291_ (.X(_03163_),
    .A(_00913_),
    .B(_03069_),
    .C(_03162_));
 sg13g2_nor2_1 _08292_ (.A(_00859_),
    .B(_03030_),
    .Y(_03164_));
 sg13g2_a21o_1 _08293_ (.A2(_03011_),
    .A1(_00940_),
    .B1(_03164_),
    .X(_03165_));
 sg13g2_or4_1 _08294_ (.A(_03163_),
    .B(_03165_),
    .C(_03072_),
    .D(_03075_),
    .X(_03166_));
 sg13g2_buf_1 _08295_ (.A(_03166_),
    .X(_03167_));
 sg13g2_nand2_1 _08296_ (.Y(_03168_),
    .A(_03079_),
    .B(_03158_));
 sg13g2_a22oi_1 _08297_ (.Y(_03169_),
    .B1(_03168_),
    .B2(_03062_),
    .A2(_03167_),
    .A1(_03060_));
 sg13g2_buf_2 _08298_ (.A(_03169_),
    .X(_03170_));
 sg13g2_nand3_1 _08299_ (.B(_03161_),
    .C(_03170_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .Y(_03171_));
 sg13g2_and4_1 _08300_ (.A(net82),
    .B(_03155_),
    .C(_03156_),
    .D(_03171_),
    .X(_03172_));
 sg13g2_a21oi_1 _08301_ (.A1(_03126_),
    .A2(_03154_),
    .Y(_03173_),
    .B1(_03172_));
 sg13g2_nor2_1 _08302_ (.A(_03125_),
    .B(_03173_),
    .Y(_03174_));
 sg13g2_buf_2 _08303_ (.A(_03174_),
    .X(_03175_));
 sg13g2_nor2_1 _08304_ (.A(net107),
    .B(_03175_),
    .Y(_03176_));
 sg13g2_a21oi_1 _08305_ (.A1(_03007_),
    .A2(_03115_),
    .Y(_03177_),
    .B1(_03176_));
 sg13g2_nor2_1 _08306_ (.A(_03005_),
    .B(_03177_),
    .Y(_03178_));
 sg13g2_a221oi_1 _08307_ (.B2(_03003_),
    .C1(_03178_),
    .B1(_03002_),
    .A1(_02976_),
    .Y(_03179_),
    .A2(_02999_));
 sg13g2_nand2_1 _08308_ (.Y(_03180_),
    .A(_01468_),
    .B(_01747_));
 sg13g2_o21ai_1 _08309_ (.B1(_03180_),
    .Y(_00327_),
    .A1(_02974_),
    .A2(_03179_));
 sg13g2_mux2_1 _08310_ (.A0(_01683_),
    .A1(net390),
    .S(net108),
    .X(_03181_));
 sg13g2_mux2_1 _08311_ (.A0(_02841_),
    .A1(_02630_),
    .S(net94),
    .X(_03182_));
 sg13g2_nor2_2 _08312_ (.A(_03123_),
    .B(_03118_),
    .Y(_03183_));
 sg13g2_mux2_1 _08313_ (.A0(_00039_),
    .A1(_00041_),
    .S(_03091_),
    .X(_03184_));
 sg13g2_buf_8 _08314_ (.A(_03118_),
    .X(_03185_));
 sg13g2_buf_1 _08315_ (.A(net81),
    .X(_03186_));
 sg13g2_a22oi_1 _08316_ (.Y(_03187_),
    .B1(_03184_),
    .B2(net64),
    .A2(_03183_),
    .A1(_00045_));
 sg13g2_inv_1 _08317_ (.Y(_03188_),
    .A(_00043_));
 sg13g2_nor2_2 _08318_ (.A(_03130_),
    .B(_03135_),
    .Y(_03189_));
 sg13g2_nand3_1 _08319_ (.B(_03161_),
    .C(_03170_),
    .A(_00046_),
    .Y(_03190_));
 sg13g2_o21ai_1 _08320_ (.B1(_03190_),
    .Y(_03191_),
    .A1(_03188_),
    .A2(_03189_));
 sg13g2_mux2_1 _08321_ (.A0(_00040_),
    .A1(_00044_),
    .S(net83),
    .X(_03192_));
 sg13g2_and2_1 _08322_ (.A(_03161_),
    .B(_03170_),
    .X(_03193_));
 sg13g2_buf_1 _08323_ (.A(_03193_),
    .X(_03194_));
 sg13g2_and3_1 _08324_ (.X(_03195_),
    .A(_00042_),
    .B(net81),
    .C(net80));
 sg13g2_a221oi_1 _08325_ (.B2(_03152_),
    .C1(_03195_),
    .B1(_03192_),
    .A1(_03113_),
    .Y(_03196_),
    .A2(_03191_));
 sg13g2_o21ai_1 _08326_ (.B1(_03196_),
    .Y(_03197_),
    .A1(_03120_),
    .A2(_03187_));
 sg13g2_buf_1 _08327_ (.A(_03197_),
    .X(_03198_));
 sg13g2_buf_1 _08328_ (.A(_03198_),
    .X(_03199_));
 sg13g2_inv_1 _08329_ (.Y(_03200_),
    .A(net52));
 sg13g2_inv_1 _08330_ (.Y(_03201_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ));
 sg13g2_inv_1 _08331_ (.Y(_03202_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ));
 sg13g2_inv_1 _08332_ (.Y(_03203_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ));
 sg13g2_inv_1 _08333_ (.Y(_03204_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ));
 sg13g2_mux4_1 _08334_ (.S0(_03066_),
    .A0(_03201_),
    .A1(_03202_),
    .A2(_03203_),
    .A3(_03204_),
    .S1(net82),
    .X(_03205_));
 sg13g2_inv_1 _08335_ (.Y(_03206_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ));
 sg13g2_inv_1 _08336_ (.Y(_03207_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ));
 sg13g2_inv_1 _08337_ (.Y(_03208_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ));
 sg13g2_inv_1 _08338_ (.Y(_03209_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ));
 sg13g2_mux4_1 _08339_ (.S0(_03066_),
    .A0(_03206_),
    .A1(_03207_),
    .A2(_03208_),
    .A3(_03209_),
    .S1(net82),
    .X(_03210_));
 sg13g2_mux2_1 _08340_ (.A0(_03205_),
    .A1(_03210_),
    .S(net65),
    .X(_03211_));
 sg13g2_buf_2 _08341_ (.A(_03211_),
    .X(_03212_));
 sg13g2_nor2_1 _08342_ (.A(net107),
    .B(_03212_),
    .Y(_03213_));
 sg13g2_a21oi_1 _08343_ (.A1(net94),
    .A2(_03200_),
    .Y(_03214_),
    .B1(_03213_));
 sg13g2_nor2_1 _08344_ (.A(_03005_),
    .B(_03214_),
    .Y(_03215_));
 sg13g2_a221oi_1 _08345_ (.B2(_03002_),
    .C1(_03215_),
    .B1(_03182_),
    .A1(_02976_),
    .Y(_03216_),
    .A2(_03181_));
 sg13g2_buf_1 _08346_ (.A(net216),
    .X(_03217_));
 sg13g2_nand2_1 _08347_ (.Y(_03218_),
    .A(net342),
    .B(net191));
 sg13g2_o21ai_1 _08348_ (.B1(_03218_),
    .Y(_00328_),
    .A1(_02974_),
    .A2(_03216_));
 sg13g2_mux2_1 _08349_ (.A0(_01736_),
    .A1(net389),
    .S(net108),
    .X(_03219_));
 sg13g2_inv_1 _08350_ (.Y(_03220_),
    .A(\z80.tv80s.i_tv80_core.SP[10] ));
 sg13g2_nand2_1 _08351_ (.Y(_03221_),
    .A(_02653_),
    .B(net108));
 sg13g2_o21ai_1 _08352_ (.B1(_03221_),
    .Y(_03222_),
    .A1(_03220_),
    .A2(net94));
 sg13g2_nand3_1 _08353_ (.B(_03091_),
    .C(net68),
    .A(_00173_),
    .Y(_03223_));
 sg13g2_nand2_1 _08354_ (.Y(_03224_),
    .A(_00172_),
    .B(_03152_));
 sg13g2_and3_1 _08355_ (.X(_03225_),
    .A(net81),
    .B(_03223_),
    .C(_03224_));
 sg13g2_buf_8 _08356_ (.A(_03112_),
    .X(_03226_));
 sg13g2_nand2_1 _08357_ (.Y(_03227_),
    .A(_00178_),
    .B(net80));
 sg13g2_nand2_1 _08358_ (.Y(_03228_),
    .A(_00175_),
    .B(_03137_));
 sg13g2_and3_1 _08359_ (.X(_03229_),
    .A(net63),
    .B(_03227_),
    .C(_03228_));
 sg13g2_and3_1 _08360_ (.X(_03230_),
    .A(_00174_),
    .B(_03082_),
    .C(_03089_));
 sg13g2_inv_1 _08361_ (.Y(_03231_),
    .A(_00176_));
 sg13g2_a21oi_1 _08362_ (.A1(_03082_),
    .A2(_03089_),
    .Y(_03232_),
    .B1(_03231_));
 sg13g2_mux2_1 _08363_ (.A0(_03230_),
    .A1(_03232_),
    .S(_03153_),
    .X(_03233_));
 sg13g2_and2_1 _08364_ (.A(_00177_),
    .B(net68),
    .X(_03234_));
 sg13g2_and4_1 _08365_ (.A(_00171_),
    .B(_03123_),
    .C(net81),
    .D(net68),
    .X(_03235_));
 sg13g2_a221oi_1 _08366_ (.B2(_03183_),
    .C1(_03235_),
    .B1(_03234_),
    .A1(_03120_),
    .Y(_03236_),
    .A2(_03233_));
 sg13g2_o21ai_1 _08367_ (.B1(_03236_),
    .Y(_03237_),
    .A1(_03225_),
    .A2(_03229_));
 sg13g2_buf_2 _08368_ (.A(_03237_),
    .X(_03238_));
 sg13g2_nor2_2 _08369_ (.A(_03123_),
    .B(_03120_),
    .Y(_03239_));
 sg13g2_a21o_1 _08370_ (.A2(_03137_),
    .A1(_00047_),
    .B1(net63),
    .X(_03240_));
 sg13g2_a221oi_1 _08371_ (.B2(_00048_),
    .C1(_03240_),
    .B1(_03152_),
    .A1(_00049_),
    .Y(_03241_),
    .A2(_03239_));
 sg13g2_a21o_1 _08372_ (.A2(_03137_),
    .A1(_00051_),
    .B1(net81),
    .X(_03242_));
 sg13g2_a221oi_1 _08373_ (.B2(_00054_),
    .C1(_03242_),
    .B1(net80),
    .A1(_00052_),
    .Y(_03243_),
    .A2(_03152_));
 sg13g2_nand3_1 _08374_ (.B(net63),
    .C(net60),
    .A(_00053_),
    .Y(_03244_));
 sg13g2_nand3_1 _08375_ (.B(net81),
    .C(_03120_),
    .A(_00050_),
    .Y(_03245_));
 sg13g2_a21o_1 _08376_ (.A2(_03245_),
    .A1(_03244_),
    .B1(net65),
    .X(_03246_));
 sg13g2_o21ai_1 _08377_ (.B1(_03246_),
    .Y(_03247_),
    .A1(_03241_),
    .A2(_03243_));
 sg13g2_buf_1 _08378_ (.A(_03247_),
    .X(_03248_));
 sg13g2_mux2_1 _08379_ (.A0(_03238_),
    .A1(net42),
    .S(_03006_),
    .X(_03249_));
 sg13g2_nor2_1 _08380_ (.A(_03005_),
    .B(_03249_),
    .Y(_03250_));
 sg13g2_a221oi_1 _08381_ (.B2(_03002_),
    .C1(_03250_),
    .B1(_03222_),
    .A1(_02976_),
    .Y(_03251_),
    .A2(_03219_));
 sg13g2_nand2_1 _08382_ (.Y(_03252_),
    .A(net341),
    .B(net191));
 sg13g2_o21ai_1 _08383_ (.B1(_03252_),
    .Y(_00329_),
    .A1(_02974_),
    .A2(_03251_));
 sg13g2_mux2_1 _08384_ (.A0(net379),
    .A1(net388),
    .S(net108),
    .X(_03253_));
 sg13g2_mux2_1 _08385_ (.A0(_02472_),
    .A1(_02681_),
    .S(_03007_),
    .X(_03254_));
 sg13g2_inv_1 _08386_ (.Y(_03255_),
    .A(_00101_));
 sg13g2_a21oi_1 _08387_ (.A1(_03045_),
    .A2(_03064_),
    .Y(_03256_),
    .B1(_03255_));
 sg13g2_a21oi_1 _08388_ (.A1(_00102_),
    .A2(_03120_),
    .Y(_03257_),
    .B1(_03256_));
 sg13g2_nand3_1 _08389_ (.B(_03091_),
    .C(_03066_),
    .A(_00097_),
    .Y(_03258_));
 sg13g2_nand3_1 _08390_ (.B(_03161_),
    .C(_03170_),
    .A(_00098_),
    .Y(_03259_));
 sg13g2_o21ai_1 _08391_ (.B1(_00095_),
    .Y(_03260_),
    .A1(_03130_),
    .A2(_03135_));
 sg13g2_o21ai_1 _08392_ (.B1(_00096_),
    .Y(_03261_),
    .A1(_03145_),
    .A2(_03150_));
 sg13g2_and4_1 _08393_ (.A(_03118_),
    .B(_03259_),
    .C(_03260_),
    .D(_03261_),
    .X(_03262_));
 sg13g2_buf_1 _08394_ (.A(_03262_),
    .X(_03263_));
 sg13g2_nand3_1 _08395_ (.B(_03045_),
    .C(_03064_),
    .A(_00100_),
    .Y(_03264_));
 sg13g2_inv_1 _08396_ (.Y(_03265_),
    .A(_00099_));
 sg13g2_a21o_1 _08397_ (.A2(_03064_),
    .A1(_03045_),
    .B1(_03265_),
    .X(_03266_));
 sg13g2_and4_1 _08398_ (.A(_03123_),
    .B(net82),
    .C(_03264_),
    .D(_03266_),
    .X(_03267_));
 sg13g2_a221oi_1 _08399_ (.B2(_03263_),
    .C1(_03267_),
    .B1(_03258_),
    .A1(_03183_),
    .Y(_03268_),
    .A2(_03257_));
 sg13g2_buf_1 _08400_ (.A(_03268_),
    .X(_03269_));
 sg13g2_buf_8 _08401_ (.A(_03269_),
    .X(_03270_));
 sg13g2_buf_1 _08402_ (.A(_03137_),
    .X(_03271_));
 sg13g2_mux2_1 _08403_ (.A0(_00055_),
    .A1(_00059_),
    .S(net66),
    .X(_03272_));
 sg13g2_mux2_1 _08404_ (.A0(_00058_),
    .A1(_00062_),
    .S(net66),
    .X(_03273_));
 sg13g2_a22oi_1 _08405_ (.Y(_03274_),
    .B1(_03273_),
    .B2(net80),
    .A2(_03272_),
    .A1(_03271_));
 sg13g2_mux2_1 _08406_ (.A0(_00057_),
    .A1(_00061_),
    .S(net63),
    .X(_03275_));
 sg13g2_mux2_1 _08407_ (.A0(_00056_),
    .A1(_00060_),
    .S(net66),
    .X(_03276_));
 sg13g2_buf_1 _08408_ (.A(_03152_),
    .X(_03277_));
 sg13g2_a22oi_1 _08409_ (.Y(_03278_),
    .B1(_03276_),
    .B2(_03277_),
    .A2(_03275_),
    .A1(_03239_));
 sg13g2_nand2_1 _08410_ (.Y(_03279_),
    .A(_03274_),
    .B(_03278_));
 sg13g2_buf_2 _08411_ (.A(_03279_),
    .X(_03280_));
 sg13g2_mux2_1 _08412_ (.A0(net55),
    .A1(_03280_),
    .S(net107),
    .X(_03281_));
 sg13g2_nor2_1 _08413_ (.A(_03005_),
    .B(_03281_),
    .Y(_03282_));
 sg13g2_a221oi_1 _08414_ (.B2(_03002_),
    .C1(_03282_),
    .B1(_03254_),
    .A1(_02976_),
    .Y(_03283_),
    .A2(_03253_));
 sg13g2_nand2_1 _08415_ (.Y(_03284_),
    .A(net340),
    .B(net191));
 sg13g2_o21ai_1 _08416_ (.B1(_03284_),
    .Y(_00330_),
    .A1(_02974_),
    .A2(_03283_));
 sg13g2_mux2_1 _08417_ (.A0(_01864_),
    .A1(net387),
    .S(net108),
    .X(_03285_));
 sg13g2_mux2_1 _08418_ (.A0(_02509_),
    .A1(_02710_),
    .S(net94),
    .X(_03286_));
 sg13g2_mux4_1 _08419_ (.S0(net60),
    .A0(_00104_),
    .A1(_00103_),
    .A2(_00108_),
    .A3(_00107_),
    .S1(net63),
    .X(_03287_));
 sg13g2_nand2_1 _08420_ (.Y(_03288_),
    .A(net65),
    .B(_03287_));
 sg13g2_mux2_1 _08421_ (.A0(_00105_),
    .A1(_00109_),
    .S(net83),
    .X(_03289_));
 sg13g2_mux2_1 _08422_ (.A0(_00106_),
    .A1(_00110_),
    .S(net83),
    .X(_03290_));
 sg13g2_a22oi_1 _08423_ (.Y(_03291_),
    .B1(_03290_),
    .B2(_03194_),
    .A2(_03289_),
    .A1(_03239_));
 sg13g2_buf_1 _08424_ (.A(_03291_),
    .X(_03292_));
 sg13g2_nand2_1 _08425_ (.Y(_03293_),
    .A(_03288_),
    .B(_03292_));
 sg13g2_buf_2 _08426_ (.A(_03293_),
    .X(_03294_));
 sg13g2_a22oi_1 _08427_ (.Y(_03295_),
    .B1(net80),
    .B2(_00070_),
    .A2(net79),
    .A1(_00067_));
 sg13g2_nand3_1 _08428_ (.B(_03091_),
    .C(net60),
    .A(_00069_),
    .Y(_03296_));
 sg13g2_and3_1 _08429_ (.X(_03297_),
    .A(net66),
    .B(_03295_),
    .C(_03296_));
 sg13g2_mux2_1 _08430_ (.A0(_00066_),
    .A1(_00065_),
    .S(net60),
    .X(_03298_));
 sg13g2_a221oi_1 _08431_ (.B2(net67),
    .C1(net66),
    .B1(_03298_),
    .A1(_00063_),
    .Y(_03299_),
    .A2(_03271_));
 sg13g2_mux2_1 _08432_ (.A0(_00064_),
    .A1(_00068_),
    .S(net63),
    .X(_03300_));
 sg13g2_nand2_1 _08433_ (.Y(_03301_),
    .A(_03277_),
    .B(_03300_));
 sg13g2_o21ai_1 _08434_ (.B1(_03301_),
    .Y(_03302_),
    .A1(_03297_),
    .A2(_03299_));
 sg13g2_buf_2 _08435_ (.A(_03302_),
    .X(_03303_));
 sg13g2_mux2_1 _08436_ (.A0(_03294_),
    .A1(_03303_),
    .S(net107),
    .X(_03304_));
 sg13g2_nor2_1 _08437_ (.A(_03005_),
    .B(_03304_),
    .Y(_03305_));
 sg13g2_a221oi_1 _08438_ (.B2(_03002_),
    .C1(_03305_),
    .B1(_03286_),
    .A1(_02976_),
    .Y(_03306_),
    .A2(_03285_));
 sg13g2_nand2_1 _08439_ (.Y(_03307_),
    .A(net338),
    .B(net191));
 sg13g2_o21ai_1 _08440_ (.B1(_03307_),
    .Y(_00331_),
    .A1(_02974_),
    .A2(_03306_));
 sg13g2_mux2_1 _08441_ (.A0(net375),
    .A1(net386),
    .S(_02998_),
    .X(_03308_));
 sg13g2_mux2_1 _08442_ (.A0(_02540_),
    .A1(_02726_),
    .S(net94),
    .X(_03309_));
 sg13g2_nand3_1 _08443_ (.B(_03161_),
    .C(_03170_),
    .A(_00114_),
    .Y(_03310_));
 sg13g2_o21ai_1 _08444_ (.B1(_00112_),
    .Y(_03311_),
    .A1(_03145_),
    .A2(_03150_));
 sg13g2_nand3_1 _08445_ (.B(_03310_),
    .C(_03311_),
    .A(net81),
    .Y(_03312_));
 sg13g2_o21ai_1 _08446_ (.B1(_00116_),
    .Y(_03313_),
    .A1(_03145_),
    .A2(_03150_));
 sg13g2_o21ai_1 _08447_ (.B1(_00115_),
    .Y(_03314_),
    .A1(_03130_),
    .A2(_03135_));
 sg13g2_nand3_1 _08448_ (.B(_03313_),
    .C(_03314_),
    .A(net63),
    .Y(_03315_));
 sg13g2_and3_1 _08449_ (.X(_03316_),
    .A(_00118_),
    .B(_03045_),
    .C(_03064_));
 sg13g2_inv_1 _08450_ (.Y(_03317_),
    .A(_00113_));
 sg13g2_a21oi_1 _08451_ (.A1(_03045_),
    .A2(_03064_),
    .Y(_03318_),
    .B1(_03317_));
 sg13g2_mux2_1 _08452_ (.A0(_03316_),
    .A1(_03318_),
    .S(net81),
    .X(_03319_));
 sg13g2_a22oi_1 _08453_ (.Y(_03320_),
    .B1(_03319_),
    .B2(net67),
    .A2(_03315_),
    .A1(_03312_));
 sg13g2_buf_2 _08454_ (.A(_03320_),
    .X(_03321_));
 sg13g2_nand3_1 _08455_ (.B(_03091_),
    .C(net63),
    .A(_00117_),
    .Y(_03322_));
 sg13g2_nand3_1 _08456_ (.B(net65),
    .C(_03185_),
    .A(_00111_),
    .Y(_03323_));
 sg13g2_a21o_1 _08457_ (.A2(_03323_),
    .A1(_03322_),
    .B1(_03120_),
    .X(_03324_));
 sg13g2_buf_2 _08458_ (.A(_03324_),
    .X(_03325_));
 sg13g2_nand2_2 _08459_ (.Y(_03326_),
    .A(_03321_),
    .B(_03325_));
 sg13g2_buf_1 _08460_ (.A(net66),
    .X(_03327_));
 sg13g2_a221oi_1 _08461_ (.B2(_00072_),
    .C1(net59),
    .B1(net62),
    .A1(_00071_),
    .Y(_03328_),
    .A2(net79));
 sg13g2_a221oi_1 _08462_ (.B2(_00076_),
    .C1(net64),
    .B1(net62),
    .A1(_00075_),
    .Y(_03329_),
    .A2(net79));
 sg13g2_mux4_1 _08463_ (.S0(net60),
    .A0(_00074_),
    .A1(_00073_),
    .A2(_00078_),
    .A3(_00077_),
    .S1(net59),
    .X(_03330_));
 sg13g2_nand2_1 _08464_ (.Y(_03331_),
    .A(net67),
    .B(_03330_));
 sg13g2_o21ai_1 _08465_ (.B1(_03331_),
    .Y(_03332_),
    .A1(_03328_),
    .A2(_03329_));
 sg13g2_buf_1 _08466_ (.A(_03332_),
    .X(_03333_));
 sg13g2_mux2_1 _08467_ (.A0(_03326_),
    .A1(_03333_),
    .S(net107),
    .X(_03334_));
 sg13g2_nor2_1 _08468_ (.A(_03005_),
    .B(_03334_),
    .Y(_03335_));
 sg13g2_a221oi_1 _08469_ (.B2(_03002_),
    .C1(_03335_),
    .B1(_03309_),
    .A1(_02976_),
    .Y(_03336_),
    .A2(_03308_));
 sg13g2_nand2_1 _08470_ (.Y(_03337_),
    .A(_01889_),
    .B(net191));
 sg13g2_o21ai_1 _08471_ (.B1(_03337_),
    .Y(_00332_),
    .A1(_02974_),
    .A2(_03336_));
 sg13g2_mux2_1 _08472_ (.A0(_02007_),
    .A1(_01399_),
    .S(_02998_),
    .X(_03338_));
 sg13g2_mux2_1 _08473_ (.A0(_02572_),
    .A1(_02757_),
    .S(net94),
    .X(_03339_));
 sg13g2_mux4_1 _08474_ (.S0(net67),
    .A0(_00119_),
    .A1(_00121_),
    .A2(_00123_),
    .A3(_00125_),
    .S1(net66),
    .X(_03340_));
 sg13g2_nand2_2 _08475_ (.Y(_03341_),
    .A(_03068_),
    .B(_03340_));
 sg13g2_mux2_1 _08476_ (.A0(_00122_),
    .A1(_00126_),
    .S(net83),
    .X(_03342_));
 sg13g2_mux2_1 _08477_ (.A0(_00120_),
    .A1(_00124_),
    .S(net83),
    .X(_03343_));
 sg13g2_a22oi_1 _08478_ (.Y(_03344_),
    .B1(_03343_),
    .B2(net62),
    .A2(_03342_),
    .A1(net80));
 sg13g2_buf_1 _08479_ (.A(_03344_),
    .X(_03345_));
 sg13g2_nand2_2 _08480_ (.Y(_03346_),
    .A(_03341_),
    .B(_03345_));
 sg13g2_a221oi_1 _08481_ (.B2(_00080_),
    .C1(net59),
    .B1(net62),
    .A1(_00079_),
    .Y(_03347_),
    .A2(net79));
 sg13g2_a221oi_1 _08482_ (.B2(_00084_),
    .C1(net64),
    .B1(net62),
    .A1(_00083_),
    .Y(_03348_),
    .A2(net79));
 sg13g2_mux4_1 _08483_ (.S0(net60),
    .A0(_00082_),
    .A1(_00081_),
    .A2(_00086_),
    .A3(_00085_),
    .S1(net59),
    .X(_03349_));
 sg13g2_nand2_1 _08484_ (.Y(_03350_),
    .A(net67),
    .B(_03349_));
 sg13g2_o21ai_1 _08485_ (.B1(_03350_),
    .Y(_03351_),
    .A1(_03347_),
    .A2(_03348_));
 sg13g2_buf_2 _08486_ (.A(_03351_),
    .X(_03352_));
 sg13g2_mux2_1 _08487_ (.A0(_03346_),
    .A1(_03352_),
    .S(net107),
    .X(_03353_));
 sg13g2_nor2_1 _08488_ (.A(_03005_),
    .B(_03353_),
    .Y(_03354_));
 sg13g2_a221oi_1 _08489_ (.B2(_03002_),
    .C1(_03354_),
    .B1(_03339_),
    .A1(_02976_),
    .Y(_03355_),
    .A2(_03338_));
 sg13g2_nand2_1 _08490_ (.Y(_03356_),
    .A(net335),
    .B(_03217_));
 sg13g2_o21ai_1 _08491_ (.B1(_03356_),
    .Y(_00333_),
    .A1(_02974_),
    .A2(_03355_));
 sg13g2_mux2_1 _08492_ (.A0(_02076_),
    .A1(net349),
    .S(net107),
    .X(_03357_));
 sg13g2_inv_1 _08493_ (.Y(_03358_),
    .A(_02593_));
 sg13g2_nand2_1 _08494_ (.Y(_03359_),
    .A(_02766_),
    .B(net108));
 sg13g2_o21ai_1 _08495_ (.B1(_03359_),
    .Y(_03360_),
    .A1(_03358_),
    .A2(net94));
 sg13g2_inv_1 _08496_ (.Y(_03361_),
    .A(_00132_));
 sg13g2_inv_1 _08497_ (.Y(_03362_),
    .A(_00131_));
 sg13g2_mux4_1 _08498_ (.S0(net68),
    .A0(_02770_),
    .A1(_02771_),
    .A2(_03361_),
    .A3(_03362_),
    .S1(net83),
    .X(_03363_));
 sg13g2_inv_1 _08499_ (.Y(_03364_),
    .A(_00134_));
 sg13g2_inv_1 _08500_ (.Y(_03365_),
    .A(_00133_));
 sg13g2_mux4_1 _08501_ (.S0(net68),
    .A0(_02772_),
    .A1(_02773_),
    .A2(_03364_),
    .A3(_03365_),
    .S1(net83),
    .X(_03366_));
 sg13g2_nand2b_1 _08502_ (.Y(_03367_),
    .B(net67),
    .A_N(_03366_));
 sg13g2_o21ai_1 _08503_ (.B1(_03367_),
    .Y(_03368_),
    .A1(_03092_),
    .A2(_03363_));
 sg13g2_mux2_1 _08504_ (.A0(_00090_),
    .A1(_00094_),
    .S(net59),
    .X(_03369_));
 sg13g2_mux2_1 _08505_ (.A0(_00088_),
    .A1(_00092_),
    .S(net59),
    .X(_03370_));
 sg13g2_a22oi_1 _08506_ (.Y(_03371_),
    .B1(_03370_),
    .B2(net62),
    .A2(_03369_),
    .A1(net80));
 sg13g2_mux2_1 _08507_ (.A0(_00087_),
    .A1(_00091_),
    .S(net59),
    .X(_03372_));
 sg13g2_mux2_1 _08508_ (.A0(_00089_),
    .A1(_00093_),
    .S(net59),
    .X(_03373_));
 sg13g2_a22oi_1 _08509_ (.Y(_03374_),
    .B1(_03373_),
    .B2(_03239_),
    .A2(_03372_),
    .A1(net79));
 sg13g2_nand2_2 _08510_ (.Y(_03375_),
    .A(_03371_),
    .B(_03374_));
 sg13g2_mux2_1 _08511_ (.A0(_03368_),
    .A1(_03375_),
    .S(net107),
    .X(_03376_));
 sg13g2_nor2_1 _08512_ (.A(_03005_),
    .B(_03376_),
    .Y(_03377_));
 sg13g2_a221oi_1 _08513_ (.B2(_03002_),
    .C1(_03377_),
    .B1(_03360_),
    .A1(_02976_),
    .Y(_03378_),
    .A2(_03357_));
 sg13g2_nand2_1 _08514_ (.Y(_03379_),
    .A(net376),
    .B(_03217_));
 sg13g2_o21ai_1 _08515_ (.B1(_03379_),
    .Y(_00334_),
    .A1(_02974_),
    .A2(_03378_));
 sg13g2_inv_1 _08516_ (.Y(_03380_),
    .A(_00031_));
 sg13g2_a22oi_1 _08517_ (.Y(_03381_),
    .B1(_01000_),
    .B2(_03380_),
    .A2(_01011_),
    .A1(_00998_));
 sg13g2_inv_1 _08518_ (.Y(_00335_),
    .A(_03381_));
 sg13g2_o21ai_1 _08519_ (.B1(net204),
    .Y(_03382_),
    .A1(_01092_),
    .A2(_01383_));
 sg13g2_a21oi_1 _08520_ (.A1(_02105_),
    .A2(_03382_),
    .Y(_03383_),
    .B1(_01229_));
 sg13g2_nand3_1 _08521_ (.B(_01064_),
    .C(_02878_),
    .A(net272),
    .Y(_03384_));
 sg13g2_or4_1 _08522_ (.A(_00854_),
    .B(net236),
    .C(_01357_),
    .D(_01162_),
    .X(_03385_));
 sg13g2_buf_1 _08523_ (.A(_03385_),
    .X(_03386_));
 sg13g2_o21ai_1 _08524_ (.B1(_03386_),
    .Y(_03387_),
    .A1(_00971_),
    .A2(_01279_));
 sg13g2_nand2_1 _08525_ (.Y(_03388_),
    .A(_01295_),
    .B(_03387_));
 sg13g2_a21o_1 _08526_ (.A2(_03388_),
    .A1(_03384_),
    .B1(_01253_),
    .X(_03389_));
 sg13g2_a22oi_1 _08527_ (.Y(_03390_),
    .B1(_01191_),
    .B2(net258),
    .A2(_00880_),
    .A1(_01410_));
 sg13g2_nand2b_1 _08528_ (.Y(_03391_),
    .B(net270),
    .A_N(_03390_));
 sg13g2_a21oi_1 _08529_ (.A1(_01156_),
    .A2(_01120_),
    .Y(_03392_),
    .B1(_02104_));
 sg13g2_nand4_1 _08530_ (.B(_03389_),
    .C(_03391_),
    .A(_00886_),
    .Y(_03393_),
    .D(_03392_));
 sg13g2_inv_1 _08531_ (.Y(_03394_),
    .A(_00027_));
 sg13g2_nor3_1 _08532_ (.A(_00739_),
    .B(_01309_),
    .C(net244),
    .Y(_03395_));
 sg13g2_a21oi_1 _08533_ (.A1(_03394_),
    .A2(_01290_),
    .Y(_03396_),
    .B1(_03395_));
 sg13g2_a22oi_1 _08534_ (.Y(_03397_),
    .B1(_00935_),
    .B2(_01352_),
    .A2(net175),
    .A1(_01141_));
 sg13g2_nand2_1 _08535_ (.Y(_03398_),
    .A(_00877_),
    .B(_00740_));
 sg13g2_a21oi_1 _08536_ (.A1(_01329_),
    .A2(_00823_),
    .Y(_03399_),
    .B1(_01088_));
 sg13g2_nor3_1 _08537_ (.A(net268),
    .B(_03398_),
    .C(_03399_),
    .Y(_03400_));
 sg13g2_nand3_1 _08538_ (.B(_01359_),
    .C(_01092_),
    .A(_00854_),
    .Y(_03401_));
 sg13g2_nor2b_1 _08539_ (.A(_03400_),
    .B_N(_03401_),
    .Y(_03402_));
 sg13g2_o21ai_1 _08540_ (.B1(_03402_),
    .Y(_03403_),
    .A1(_00703_),
    .A2(_03397_));
 sg13g2_nor2_1 _08541_ (.A(net267),
    .B(_01172_),
    .Y(_03404_));
 sg13g2_a21oi_1 _08542_ (.A1(_03394_),
    .A2(_01101_),
    .Y(_03405_),
    .B1(_03404_));
 sg13g2_a22oi_1 _08543_ (.Y(_03406_),
    .B1(_02960_),
    .B2(net208),
    .A2(_00959_),
    .A1(net272));
 sg13g2_buf_1 _08544_ (.A(_03406_),
    .X(_03407_));
 sg13g2_o21ai_1 _08545_ (.B1(_03407_),
    .Y(_03408_),
    .A1(_00894_),
    .A2(_03405_));
 sg13g2_and2_1 _08546_ (.A(_01123_),
    .B(_01151_),
    .X(_03409_));
 sg13g2_buf_1 _08547_ (.A(_03409_),
    .X(_03410_));
 sg13g2_nand2b_1 _08548_ (.Y(_03411_),
    .B(_00712_),
    .A_N(_02277_));
 sg13g2_nor2_1 _08549_ (.A(_00951_),
    .B(_03411_),
    .Y(_03412_));
 sg13g2_a21oi_1 _08550_ (.A1(_01147_),
    .A2(_03410_),
    .Y(_03413_),
    .B1(_03412_));
 sg13g2_nor2_1 _08551_ (.A(_01253_),
    .B(_03413_),
    .Y(_03414_));
 sg13g2_nor3_1 _08552_ (.A(_03403_),
    .B(_03408_),
    .C(_03414_),
    .Y(_03415_));
 sg13g2_o21ai_1 _08553_ (.B1(_03415_),
    .Y(_03416_),
    .A1(_01380_),
    .A2(_03396_));
 sg13g2_a22oi_1 _08554_ (.Y(_03417_),
    .B1(_03416_),
    .B2(_00860_),
    .A2(_03393_),
    .A1(_03383_));
 sg13g2_o21ai_1 _08555_ (.B1(net237),
    .Y(_03418_),
    .A1(net358),
    .A2(_00866_));
 sg13g2_o21ai_1 _08556_ (.B1(_03418_),
    .Y(_03419_),
    .A1(net353),
    .A2(_03417_));
 sg13g2_buf_1 _08557_ (.A(_03419_),
    .X(_03420_));
 sg13g2_nand2_1 _08558_ (.Y(_03421_),
    .A(net282),
    .B(_00640_));
 sg13g2_nor2_1 _08559_ (.A(_00752_),
    .B(_03421_),
    .Y(_03422_));
 sg13g2_nor3_1 _08560_ (.A(net307),
    .B(net233),
    .C(_02277_),
    .Y(_03423_));
 sg13g2_o21ai_1 _08561_ (.B1(_02878_),
    .Y(_03424_),
    .A1(_03422_),
    .A2(_03423_));
 sg13g2_o21ai_1 _08562_ (.B1(_03424_),
    .Y(_03425_),
    .A1(net307),
    .A2(_03386_));
 sg13g2_nand2_1 _08563_ (.Y(_03426_),
    .A(_00886_),
    .B(_02202_));
 sg13g2_a221oi_1 _08564_ (.B2(net271),
    .C1(_03426_),
    .B1(_03425_),
    .A1(net183),
    .Y(_03427_),
    .A2(_01371_));
 sg13g2_inv_1 _08565_ (.Y(_03428_),
    .A(_00025_));
 sg13g2_nor3_1 _08566_ (.A(net275),
    .B(_01309_),
    .C(net244),
    .Y(_03429_));
 sg13g2_a21oi_1 _08567_ (.A1(_03428_),
    .A2(net244),
    .Y(_03430_),
    .B1(_03429_));
 sg13g2_a21oi_1 _08568_ (.A1(_03428_),
    .A2(_01101_),
    .Y(_03431_),
    .B1(_03404_));
 sg13g2_nand2_1 _08569_ (.Y(_03432_),
    .A(_00897_),
    .B(_01363_));
 sg13g2_o21ai_1 _08570_ (.B1(_03432_),
    .Y(_03433_),
    .A1(_00894_),
    .A2(_03431_));
 sg13g2_o21ai_1 _08571_ (.B1(_03411_),
    .Y(_03434_),
    .A1(_01161_),
    .A2(_02268_));
 sg13g2_a22oi_1 _08572_ (.Y(_03435_),
    .B1(_03434_),
    .B2(_00760_),
    .A2(_03410_),
    .A1(_00640_));
 sg13g2_o21ai_1 _08573_ (.B1(_01582_),
    .Y(_03436_),
    .A1(net185),
    .A2(_03012_));
 sg13g2_a22oi_1 _08574_ (.Y(_03437_),
    .B1(_03436_),
    .B2(_01156_),
    .A2(_01283_),
    .A1(_01163_));
 sg13g2_o21ai_1 _08575_ (.B1(_03437_),
    .Y(_03438_),
    .A1(_01295_),
    .A2(_03435_));
 sg13g2_nor4_1 _08576_ (.A(_02926_),
    .B(_03403_),
    .C(_03433_),
    .D(_03438_),
    .Y(_03439_));
 sg13g2_o21ai_1 _08577_ (.B1(_03439_),
    .Y(_03440_),
    .A1(_01380_),
    .A2(_03430_));
 sg13g2_a21oi_1 _08578_ (.A1(_00860_),
    .A2(_03440_),
    .Y(_03441_),
    .B1(_02939_));
 sg13g2_nor3_2 _08579_ (.A(_00866_),
    .B(_03427_),
    .C(_03441_),
    .Y(_03442_));
 sg13g2_nor2_1 _08580_ (.A(_00845_),
    .B(net277),
    .Y(_03443_));
 sg13g2_a22oi_1 _08581_ (.Y(_03444_),
    .B1(_03443_),
    .B2(_01329_),
    .A2(_00897_),
    .A1(_00847_));
 sg13g2_nor4_1 _08582_ (.A(net324),
    .B(_00923_),
    .C(_00802_),
    .D(net230),
    .Y(_03445_));
 sg13g2_nand3_1 _08583_ (.B(_01413_),
    .C(_03445_),
    .A(_00955_),
    .Y(_03446_));
 sg13g2_nand3_1 _08584_ (.B(_00655_),
    .C(_00918_),
    .A(_01410_),
    .Y(_03447_));
 sg13g2_and2_1 _08585_ (.A(_02263_),
    .B(_02981_),
    .X(_03448_));
 sg13g2_nand4_1 _08586_ (.B(_03447_),
    .C(_01435_),
    .A(_02909_),
    .Y(_03449_),
    .D(_03448_));
 sg13g2_nor4_1 _08587_ (.A(_00848_),
    .B(_02365_),
    .C(_03446_),
    .D(_03449_),
    .Y(_03450_));
 sg13g2_nand3b_1 _08588_ (.B(_02905_),
    .C(_03450_),
    .Y(_03451_),
    .A_N(_02273_));
 sg13g2_nand4_1 _08589_ (.B(_03437_),
    .C(_03444_),
    .A(_03407_),
    .Y(_03452_),
    .D(_03451_));
 sg13g2_a21oi_1 _08590_ (.A1(net214),
    .A2(_02878_),
    .Y(_03453_),
    .B1(net237));
 sg13g2_nand2_1 _08591_ (.Y(_03454_),
    .A(net273),
    .B(_00728_));
 sg13g2_a21oi_1 _08592_ (.A1(_02878_),
    .A2(_03454_),
    .Y(_03455_),
    .B1(net183));
 sg13g2_nand2_1 _08593_ (.Y(_03456_),
    .A(_01064_),
    .B(_02878_));
 sg13g2_o21ai_1 _08594_ (.B1(_02090_),
    .Y(_03457_),
    .A1(net244),
    .A2(_03456_));
 sg13g2_o21ai_1 _08595_ (.B1(_03386_),
    .Y(_03458_),
    .A1(_01279_),
    .A2(net277));
 sg13g2_a22oi_1 _08596_ (.Y(_03459_),
    .B1(_03458_),
    .B2(_01329_),
    .A2(_03457_),
    .A1(_00942_));
 sg13g2_nor4_1 _08597_ (.A(_00863_),
    .B(_03453_),
    .C(_03455_),
    .D(_03459_),
    .Y(_03460_));
 sg13g2_mux2_1 _08598_ (.A0(_03452_),
    .A1(_03460_),
    .S(_00967_),
    .X(_03461_));
 sg13g2_and2_1 _08599_ (.A(net302),
    .B(_03461_),
    .X(_03462_));
 sg13g2_buf_1 _08600_ (.A(_03462_),
    .X(_03463_));
 sg13g2_nand2b_1 _08601_ (.Y(_03464_),
    .B(_03463_),
    .A_N(_03442_));
 sg13g2_nor2_1 _08602_ (.A(_03420_),
    .B(_03464_),
    .Y(_03465_));
 sg13g2_buf_1 _08603_ (.A(_03465_),
    .X(_03466_));
 sg13g2_inv_2 _08604_ (.Y(_03467_),
    .A(_02294_));
 sg13g2_or2_1 _08605_ (.X(_03468_),
    .B(_03384_),
    .A(_01252_));
 sg13g2_nand3_1 _08606_ (.B(net230),
    .C(net170),
    .A(_01016_),
    .Y(_03469_));
 sg13g2_nand3_1 _08607_ (.B(_03468_),
    .C(_03469_),
    .A(_02202_),
    .Y(_03470_));
 sg13g2_nand2_1 _08608_ (.Y(_03471_),
    .A(_01044_),
    .B(_01330_));
 sg13g2_o21ai_1 _08609_ (.B1(_03471_),
    .Y(_03472_),
    .A1(net199),
    .A2(_01357_));
 sg13g2_and2_1 _08610_ (.A(net199),
    .B(_03015_),
    .X(_03473_));
 sg13g2_a22oi_1 _08611_ (.Y(_03474_),
    .B1(_03473_),
    .B2(_01092_),
    .A2(_03472_),
    .A1(_00891_));
 sg13g2_nor3_1 _08612_ (.A(_01016_),
    .B(net236),
    .C(_03474_),
    .Y(_03475_));
 sg13g2_or2_1 _08613_ (.X(_03476_),
    .B(_03421_),
    .A(net244));
 sg13g2_nor2_1 _08614_ (.A(_00215_),
    .B(_02133_),
    .Y(_03477_));
 sg13g2_nand2_1 _08615_ (.Y(_03478_),
    .A(_00723_),
    .B(_03477_));
 sg13g2_a21oi_1 _08616_ (.A1(_03476_),
    .A2(_03478_),
    .Y(_03479_),
    .B1(_02929_));
 sg13g2_a22oi_1 _08617_ (.Y(_03480_),
    .B1(_03477_),
    .B2(_01117_),
    .A2(_01371_),
    .A1(net205));
 sg13g2_nand3_1 _08618_ (.B(net209),
    .C(_01084_),
    .A(_00970_),
    .Y(_03481_));
 sg13g2_a21oi_1 _08619_ (.A1(_00942_),
    .A2(_01329_),
    .Y(_03482_),
    .B1(_02941_));
 sg13g2_nand2b_1 _08620_ (.Y(_03483_),
    .B(_03410_),
    .A_N(_03482_));
 sg13g2_nand4_1 _08621_ (.B(_03480_),
    .C(_03481_),
    .A(_03402_),
    .Y(_03484_),
    .D(_03483_));
 sg13g2_a21oi_1 _08622_ (.A1(net209),
    .A2(net199),
    .Y(_03485_),
    .B1(_01363_));
 sg13g2_nor2_1 _08623_ (.A(net234),
    .B(net240),
    .Y(_03486_));
 sg13g2_o21ai_1 _08624_ (.B1(_00961_),
    .Y(_03487_),
    .A1(_00962_),
    .A2(_03486_));
 sg13g2_o21ai_1 _08625_ (.B1(_03487_),
    .Y(_03488_),
    .A1(_00705_),
    .A2(_03485_));
 sg13g2_nor4_1 _08626_ (.A(net270),
    .B(_00971_),
    .C(_00657_),
    .D(net210),
    .Y(_03489_));
 sg13g2_nor4_1 _08627_ (.A(_03479_),
    .B(_03484_),
    .C(_03488_),
    .D(_03489_),
    .Y(_03490_));
 sg13g2_o21ai_1 _08628_ (.B1(_02994_),
    .Y(_03491_),
    .A1(net305),
    .A2(_03490_));
 sg13g2_o21ai_1 _08629_ (.B1(_03491_),
    .Y(_03492_),
    .A1(_03470_),
    .A2(_03475_));
 sg13g2_and2_1 _08630_ (.A(net353),
    .B(_00215_),
    .X(_03493_));
 sg13g2_a21oi_1 _08631_ (.A1(net302),
    .A2(_03492_),
    .Y(_03494_),
    .B1(_03493_));
 sg13g2_buf_2 _08632_ (.A(_03494_),
    .X(_03495_));
 sg13g2_buf_1 _08633_ (.A(_03495_),
    .X(_03496_));
 sg13g2_nand2_1 _08634_ (.Y(_03497_),
    .A(_02812_),
    .B(net92));
 sg13g2_o21ai_1 _08635_ (.B1(_03497_),
    .Y(_03498_),
    .A1(_03467_),
    .A2(net92));
 sg13g2_buf_1 _08636_ (.A(_03420_),
    .X(_03499_));
 sg13g2_and2_1 _08637_ (.A(_03461_),
    .B(_03442_),
    .X(_03500_));
 sg13g2_nor2b_1 _08638_ (.A(_03499_),
    .B_N(_03500_),
    .Y(_03501_));
 sg13g2_buf_1 _08639_ (.A(_03501_),
    .X(_03502_));
 sg13g2_mux2_1 _08640_ (.A0(_02315_),
    .A1(_02802_),
    .S(net92),
    .X(_03503_));
 sg13g2_a22oi_1 _08641_ (.Y(_03504_),
    .B1(_03502_),
    .B2(_03503_),
    .A2(_03498_),
    .A1(_03466_));
 sg13g2_a21oi_2 _08642_ (.B1(_03442_),
    .Y(_03505_),
    .A2(_00866_),
    .A1(_03428_));
 sg13g2_nor2_1 _08643_ (.A(_03463_),
    .B(_03505_),
    .Y(_03506_));
 sg13g2_inv_1 _08644_ (.Y(_03507_),
    .A(_03464_));
 sg13g2_a21oi_1 _08645_ (.A1(net350),
    .A2(_03506_),
    .Y(_03508_),
    .B1(_03507_));
 sg13g2_and2_1 _08646_ (.A(_01545_),
    .B(_03495_),
    .X(_03509_));
 sg13g2_a22oi_1 _08647_ (.Y(_03510_),
    .B1(_03506_),
    .B2(_03509_),
    .A2(_03507_),
    .A1(net391));
 sg13g2_o21ai_1 _08648_ (.B1(_03510_),
    .Y(_03511_),
    .A1(net92),
    .A2(_03508_));
 sg13g2_inv_1 _08649_ (.Y(_03512_),
    .A(_03505_));
 sg13g2_a21oi_1 _08650_ (.A1(net106),
    .A2(_03512_),
    .Y(_03513_),
    .B1(_03463_));
 sg13g2_buf_2 _08651_ (.A(_03513_),
    .X(_03514_));
 sg13g2_buf_1 _08652_ (.A(_03142_),
    .X(_03515_));
 sg13g2_buf_1 _08653_ (.A(net143),
    .X(_03516_));
 sg13g2_nand2b_1 _08654_ (.Y(_03517_),
    .B(net135),
    .A_N(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ));
 sg13g2_nand2b_1 _08655_ (.Y(_03518_),
    .B(net135),
    .A_N(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ));
 sg13g2_mux2_1 _08656_ (.A0(_02850_),
    .A1(_00213_),
    .S(_03142_),
    .X(_03519_));
 sg13g2_buf_2 _08657_ (.A(_03519_),
    .X(_03520_));
 sg13g2_buf_1 _08658_ (.A(_03520_),
    .X(_03521_));
 sg13g2_buf_1 _08659_ (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .X(_03522_));
 sg13g2_buf_1 _08660_ (.A(_03522_),
    .X(_03523_));
 sg13g2_buf_1 _08661_ (.A(net327),
    .X(_03524_));
 sg13g2_mux4_1 _08662_ (.S0(net121),
    .A0(_03517_),
    .A1(_03518_),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .S1(net289),
    .X(_03525_));
 sg13g2_buf_2 _08663_ (.A(_03520_),
    .X(_03526_));
 sg13g2_nor2_1 _08664_ (.A(_03522_),
    .B(net144),
    .Y(_03527_));
 sg13g2_buf_2 _08665_ (.A(_03527_),
    .X(_03528_));
 sg13g2_mux4_1 _08666_ (.S0(net120),
    .A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ),
    .S1(_03528_),
    .X(_03529_));
 sg13g2_buf_1 _08667_ (.A(net143),
    .X(_03530_));
 sg13g2_nand2b_1 _08668_ (.Y(_03531_),
    .B(net134),
    .A_N(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ));
 sg13g2_nand2b_1 _08669_ (.Y(_03532_),
    .B(net134),
    .A_N(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ));
 sg13g2_mux4_1 _08670_ (.S0(net121),
    .A0(_03531_),
    .A1(_03532_),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .S1(net289),
    .X(_03533_));
 sg13g2_buf_2 _08671_ (.A(_03520_),
    .X(_03534_));
 sg13g2_buf_1 _08672_ (.A(_03528_),
    .X(_03535_));
 sg13g2_mux4_1 _08673_ (.S0(net119),
    .A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ),
    .S1(net105),
    .X(_03536_));
 sg13g2_nand2_1 _08674_ (.Y(_03537_),
    .A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .B(_03515_));
 sg13g2_buf_4 _08675_ (.X(_03538_),
    .A(_03537_));
 sg13g2_mux4_1 _08676_ (.S0(_03538_),
    .A0(_03525_),
    .A1(_03529_),
    .A2(_03533_),
    .A3(_03536_),
    .S1(net92),
    .X(_03539_));
 sg13g2_a22oi_1 _08677_ (.Y(_03540_),
    .B1(_03514_),
    .B2(_03539_),
    .A2(_03511_),
    .A1(net106));
 sg13g2_a21o_1 _08678_ (.A2(_03500_),
    .A1(net106),
    .B1(net263),
    .X(_03541_));
 sg13g2_buf_2 _08679_ (.A(_03541_),
    .X(_03542_));
 sg13g2_a21oi_1 _08680_ (.A1(_03504_),
    .A2(_03540_),
    .Y(_03543_),
    .B1(_03542_));
 sg13g2_a21o_1 _08681_ (.A2(net197),
    .A1(net348),
    .B1(_03543_),
    .X(_00336_));
 sg13g2_nand2b_1 _08682_ (.Y(_03544_),
    .B(net134),
    .A_N(_00045_));
 sg13g2_nand2b_1 _08683_ (.Y(_03545_),
    .B(net134),
    .A_N(_00041_));
 sg13g2_mux4_1 _08684_ (.S0(net121),
    .A0(_03544_),
    .A1(_03545_),
    .A2(_00046_),
    .A3(_00042_),
    .S1(net289),
    .X(_03546_));
 sg13g2_mux4_1 _08685_ (.S0(net119),
    .A0(_00044_),
    .A1(_00040_),
    .A2(_00043_),
    .A3(_00039_),
    .S1(net105),
    .X(_03547_));
 sg13g2_buf_1 _08686_ (.A(_03142_),
    .X(_03548_));
 sg13g2_nand2b_1 _08687_ (.Y(_03549_),
    .B(net142),
    .A_N(_00167_));
 sg13g2_nand2b_1 _08688_ (.Y(_03550_),
    .B(_03530_),
    .A_N(_00163_));
 sg13g2_mux4_1 _08689_ (.S0(net121),
    .A0(_03549_),
    .A1(_03550_),
    .A2(_00168_),
    .A3(_00164_),
    .S1(net289),
    .X(_03551_));
 sg13g2_inv_1 _08690_ (.Y(_03552_),
    .A(_03520_));
 sg13g2_mux4_1 _08691_ (.S0(_03552_),
    .A0(_00162_),
    .A1(_00166_),
    .A2(_00161_),
    .A3(_00165_),
    .S1(net105),
    .X(_03553_));
 sg13g2_mux4_1 _08692_ (.S0(_03538_),
    .A0(_03546_),
    .A1(_03547_),
    .A2(_03551_),
    .A3(_03553_),
    .S1(net92),
    .X(_03554_));
 sg13g2_inv_1 _08693_ (.Y(_03555_),
    .A(_03554_));
 sg13g2_and2_1 _08694_ (.A(_03420_),
    .B(_03506_),
    .X(_03556_));
 sg13g2_buf_1 _08695_ (.A(_03556_),
    .X(_03557_));
 sg13g2_nor2b_1 _08696_ (.A(_03495_),
    .B_N(net91),
    .Y(_03558_));
 sg13g2_buf_1 _08697_ (.A(_03558_),
    .X(_03559_));
 sg13g2_buf_1 _08698_ (.A(_03495_),
    .X(_03560_));
 sg13g2_nor2_1 _08699_ (.A(_02619_),
    .B(net90),
    .Y(_03561_));
 sg13g2_a21oi_1 _08700_ (.A1(_00142_),
    .A2(net90),
    .Y(_03562_),
    .B1(_03561_));
 sg13g2_nand2_1 _08701_ (.Y(_03563_),
    .A(net78),
    .B(_03562_));
 sg13g2_nor3_1 _08702_ (.A(net106),
    .B(_03464_),
    .C(_03495_),
    .Y(_03564_));
 sg13g2_and3_1 _08703_ (.X(_03565_),
    .A(net106),
    .B(_03507_),
    .C(_03495_));
 sg13g2_buf_1 _08704_ (.A(_03565_),
    .X(_03566_));
 sg13g2_a22oi_1 _08705_ (.Y(_03567_),
    .B1(_03566_),
    .B2(net337),
    .A2(_03564_),
    .A1(_02630_));
 sg13g2_a22oi_1 _08706_ (.Y(_03568_),
    .B1(net91),
    .B2(_01683_),
    .A2(net93),
    .A1(_02841_));
 sg13g2_buf_1 _08707_ (.A(net90),
    .X(_03569_));
 sg13g2_nand2b_1 _08708_ (.Y(_03570_),
    .B(net77),
    .A_N(_03568_));
 sg13g2_nand3_1 _08709_ (.B(_03567_),
    .C(_03570_),
    .A(_03563_),
    .Y(_03571_));
 sg13g2_a221oi_1 _08710_ (.B2(net390),
    .C1(_03571_),
    .B1(_03559_),
    .A1(_03514_),
    .Y(_03572_),
    .A2(_03555_));
 sg13g2_nand2_1 _08711_ (.Y(_03573_),
    .A(_01636_),
    .B(net191));
 sg13g2_o21ai_1 _08712_ (.B1(_03573_),
    .Y(_00337_),
    .A1(_03542_),
    .A2(_03572_));
 sg13g2_nand2b_1 _08713_ (.Y(_03574_),
    .B(net134),
    .A_N(_00053_));
 sg13g2_nand2b_1 _08714_ (.Y(_03575_),
    .B(net134),
    .A_N(_00049_));
 sg13g2_mux4_1 _08715_ (.S0(net121),
    .A0(_03574_),
    .A1(_03575_),
    .A2(_00054_),
    .A3(_00050_),
    .S1(net289),
    .X(_03576_));
 sg13g2_mux4_1 _08716_ (.S0(net119),
    .A0(_00052_),
    .A1(_00048_),
    .A2(_00051_),
    .A3(_00047_),
    .S1(net105),
    .X(_03577_));
 sg13g2_nand2b_1 _08717_ (.Y(_03578_),
    .B(net142),
    .A_N(_00177_));
 sg13g2_nand2b_1 _08718_ (.Y(_03579_),
    .B(net142),
    .A_N(_00173_));
 sg13g2_mux4_1 _08719_ (.S0(net119),
    .A0(_03578_),
    .A1(_03579_),
    .A2(_00178_),
    .A3(_00174_),
    .S1(_03524_),
    .X(_03580_));
 sg13g2_mux4_1 _08720_ (.S0(_03552_),
    .A0(_00172_),
    .A1(_00176_),
    .A2(_00171_),
    .A3(_00175_),
    .S1(net105),
    .X(_03581_));
 sg13g2_mux4_1 _08721_ (.S0(_03538_),
    .A0(_03576_),
    .A1(_03577_),
    .A2(_03580_),
    .A3(_03581_),
    .S1(net92),
    .X(_03582_));
 sg13g2_nor2b_1 _08722_ (.A(_03582_),
    .B_N(_03514_),
    .Y(_03583_));
 sg13g2_and2_1 _08723_ (.A(net389),
    .B(_03559_),
    .X(_03584_));
 sg13g2_nand2_1 _08724_ (.Y(_03585_),
    .A(net90),
    .B(_03501_));
 sg13g2_nand2_1 _08725_ (.Y(_03586_),
    .A(_00685_),
    .B(_03566_));
 sg13g2_o21ai_1 _08726_ (.B1(_03586_),
    .Y(_03587_),
    .A1(_02410_),
    .A2(_03585_));
 sg13g2_a22oi_1 _08727_ (.Y(_03588_),
    .B1(net91),
    .B2(_01736_),
    .A2(net93),
    .A1(\z80.tv80s.i_tv80_core.SP[10] ));
 sg13g2_a221oi_1 _08728_ (.B2(_02640_),
    .C1(net77),
    .B1(net78),
    .A1(_02653_),
    .Y(_03589_),
    .A2(net93));
 sg13g2_a21oi_1 _08729_ (.A1(net77),
    .A2(_03588_),
    .Y(_03590_),
    .B1(_03589_));
 sg13g2_nor4_1 _08730_ (.A(_03583_),
    .B(_03584_),
    .C(_03587_),
    .D(_03590_),
    .Y(_03591_));
 sg13g2_nand2_1 _08731_ (.Y(_03592_),
    .A(net380),
    .B(net191));
 sg13g2_o21ai_1 _08732_ (.B1(_03592_),
    .Y(_00338_),
    .A1(_03542_),
    .A2(_03591_));
 sg13g2_a22oi_1 _08733_ (.Y(_03593_),
    .B1(net91),
    .B2(net379),
    .A2(net78),
    .A1(_02460_));
 sg13g2_buf_1 _08734_ (.A(\z80.tv80s.i_tv80_core.PC[3] ),
    .X(_03594_));
 sg13g2_a221oi_1 _08735_ (.B2(net388),
    .C1(_03496_),
    .B1(net91),
    .A1(_03594_),
    .Y(_03595_),
    .A2(net78));
 sg13g2_a21o_1 _08736_ (.A2(_03593_),
    .A1(net77),
    .B1(_03595_),
    .X(_03596_));
 sg13g2_mux2_1 _08737_ (.A0(_02681_),
    .A1(_02472_),
    .S(_03495_),
    .X(_03597_));
 sg13g2_nand2b_1 _08738_ (.Y(_03598_),
    .B(_03597_),
    .A_N(_03499_));
 sg13g2_buf_1 _08739_ (.A(\z80.tv80s.i_tv80_core.F[3] ),
    .X(_03599_));
 sg13g2_nand3_1 _08740_ (.B(net106),
    .C(net90),
    .A(_03599_),
    .Y(_03600_));
 sg13g2_nand2_1 _08741_ (.Y(_03601_),
    .A(_03598_),
    .B(_03600_));
 sg13g2_nand2b_1 _08742_ (.Y(_03602_),
    .B(net143),
    .A_N(_00061_));
 sg13g2_nand2b_1 _08743_ (.Y(_03603_),
    .B(net143),
    .A_N(_00057_));
 sg13g2_mux4_1 _08744_ (.S0(net120),
    .A0(_03602_),
    .A1(_03603_),
    .A2(_00062_),
    .A3(_00058_),
    .S1(net327),
    .X(_03604_));
 sg13g2_mux4_1 _08745_ (.S0(net120),
    .A0(_00060_),
    .A1(_00056_),
    .A2(_00059_),
    .A3(_00055_),
    .S1(_03528_),
    .X(_03605_));
 sg13g2_nand2_1 _08746_ (.Y(_03606_),
    .A(_03255_),
    .B(net143));
 sg13g2_nand2b_1 _08747_ (.Y(_03607_),
    .B(_03515_),
    .A_N(_00097_));
 sg13g2_mux4_1 _08748_ (.S0(_03526_),
    .A0(_03606_),
    .A1(_03607_),
    .A2(_00102_),
    .A3(_00098_),
    .S1(net327),
    .X(_03608_));
 sg13g2_mux4_1 _08749_ (.S0(_03520_),
    .A0(_00100_),
    .A1(_00096_),
    .A2(_00099_),
    .A3(_00095_),
    .S1(_03528_),
    .X(_03609_));
 sg13g2_mux4_1 _08750_ (.S0(_03538_),
    .A0(_03604_),
    .A1(_03605_),
    .A2(_03608_),
    .A3(_03609_),
    .S1(net90),
    .X(_03610_));
 sg13g2_nor2b_1 _08751_ (.A(_03610_),
    .B_N(_03514_),
    .Y(_03611_));
 sg13g2_a21oi_1 _08752_ (.A1(_03507_),
    .A2(_03601_),
    .Y(_03612_),
    .B1(_03611_));
 sg13g2_a21oi_1 _08753_ (.A1(_03596_),
    .A2(_03612_),
    .Y(_03613_),
    .B1(_03542_));
 sg13g2_a21o_1 _08754_ (.A2(net197),
    .A1(_01757_),
    .B1(_03613_),
    .X(_00339_));
 sg13g2_nand2b_1 _08755_ (.Y(_03614_),
    .B(net142),
    .A_N(_00069_));
 sg13g2_nand2b_1 _08756_ (.Y(_03615_),
    .B(net142),
    .A_N(_00065_));
 sg13g2_mux4_1 _08757_ (.S0(net119),
    .A0(_03614_),
    .A1(_03615_),
    .A2(_00070_),
    .A3(_00066_),
    .S1(net327),
    .X(_03616_));
 sg13g2_mux4_1 _08758_ (.S0(net119),
    .A0(_00068_),
    .A1(_00064_),
    .A2(_00067_),
    .A3(_00063_),
    .S1(net105),
    .X(_03617_));
 sg13g2_nand2b_1 _08759_ (.Y(_03618_),
    .B(net143),
    .A_N(_00109_));
 sg13g2_nand2b_1 _08760_ (.Y(_03619_),
    .B(net142),
    .A_N(_00105_));
 sg13g2_mux4_1 _08761_ (.S0(_03526_),
    .A0(_03618_),
    .A1(_03619_),
    .A2(_00110_),
    .A3(_00106_),
    .S1(net327),
    .X(_03620_));
 sg13g2_mux4_1 _08762_ (.S0(net120),
    .A0(_00108_),
    .A1(_00104_),
    .A2(_00107_),
    .A3(_00103_),
    .S1(_03528_),
    .X(_03621_));
 sg13g2_mux4_1 _08763_ (.S0(_03538_),
    .A0(_03616_),
    .A1(_03617_),
    .A2(_03620_),
    .A3(_03621_),
    .S1(net90),
    .X(_03622_));
 sg13g2_nand2b_1 _08764_ (.Y(_03623_),
    .B(_03514_),
    .A_N(_03622_));
 sg13g2_nor2_1 _08765_ (.A(_02498_),
    .B(_03585_),
    .Y(_03624_));
 sg13g2_a221oi_1 _08766_ (.B2(_01653_),
    .C1(_03624_),
    .B1(_03566_),
    .A1(net387),
    .Y(_03625_),
    .A2(_03559_));
 sg13g2_a22oi_1 _08767_ (.Y(_03626_),
    .B1(net91),
    .B2(_01864_),
    .A2(net93),
    .A1(_02509_));
 sg13g2_buf_2 _08768_ (.A(\z80.tv80s.i_tv80_core.PC[4] ),
    .X(_03627_));
 sg13g2_a221oi_1 _08769_ (.B2(_03627_),
    .C1(_03560_),
    .B1(net78),
    .A1(_02710_),
    .Y(_03628_),
    .A2(net93));
 sg13g2_a21o_1 _08770_ (.A2(_03626_),
    .A1(net77),
    .B1(_03628_),
    .X(_03629_));
 sg13g2_nand3_1 _08771_ (.B(_03625_),
    .C(_03629_),
    .A(_03623_),
    .Y(_03630_));
 sg13g2_nand2b_1 _08772_ (.Y(_03631_),
    .B(_03630_),
    .A_N(_03542_));
 sg13g2_o21ai_1 _08773_ (.B1(_03631_),
    .Y(_00340_),
    .A1(_01830_),
    .A2(net194));
 sg13g2_nand2b_1 _08774_ (.Y(_03632_),
    .B(net134),
    .A_N(_00077_));
 sg13g2_nand2b_1 _08775_ (.Y(_03633_),
    .B(net134),
    .A_N(_00073_));
 sg13g2_mux4_1 _08776_ (.S0(net121),
    .A0(_03632_),
    .A1(_03633_),
    .A2(_00078_),
    .A3(_00074_),
    .S1(net289),
    .X(_03634_));
 sg13g2_mux4_1 _08777_ (.S0(net119),
    .A0(_00076_),
    .A1(_00072_),
    .A2(_00075_),
    .A3(_00071_),
    .S1(net105),
    .X(_03635_));
 sg13g2_nand2b_1 _08778_ (.Y(_03636_),
    .B(_03548_),
    .A_N(_00117_));
 sg13g2_nand2_1 _08779_ (.Y(_03637_),
    .A(_03317_),
    .B(_03548_));
 sg13g2_mux4_1 _08780_ (.S0(net119),
    .A0(_03636_),
    .A1(_03637_),
    .A2(_00118_),
    .A3(_00114_),
    .S1(net289),
    .X(_03638_));
 sg13g2_mux4_1 _08781_ (.S0(_03534_),
    .A0(_00116_),
    .A1(_00112_),
    .A2(_00115_),
    .A3(_00111_),
    .S1(_03535_),
    .X(_03639_));
 sg13g2_mux4_1 _08782_ (.S0(_03538_),
    .A0(_03634_),
    .A1(_03635_),
    .A2(_03638_),
    .A3(_03639_),
    .S1(net92),
    .X(_03640_));
 sg13g2_nor2b_1 _08783_ (.A(_03640_),
    .B_N(_03514_),
    .Y(_03641_));
 sg13g2_and2_1 _08784_ (.A(net386),
    .B(_03559_),
    .X(_03642_));
 sg13g2_buf_1 _08785_ (.A(\z80.tv80s.i_tv80_core.F[5] ),
    .X(_03643_));
 sg13g2_nand2_1 _08786_ (.Y(_03644_),
    .A(_03643_),
    .B(_03566_));
 sg13g2_o21ai_1 _08787_ (.B1(_03644_),
    .Y(_03645_),
    .A1(_02530_),
    .A2(_03585_));
 sg13g2_a22oi_1 _08788_ (.Y(_03646_),
    .B1(net91),
    .B2(_01948_),
    .A2(net93),
    .A1(_02540_));
 sg13g2_a221oi_1 _08789_ (.B2(\z80.tv80s.i_tv80_core.PC[5] ),
    .C1(net77),
    .B1(net78),
    .A1(_02726_),
    .Y(_03647_),
    .A2(net93));
 sg13g2_a21oi_1 _08790_ (.A1(net77),
    .A2(_03646_),
    .Y(_03648_),
    .B1(_03647_));
 sg13g2_nor4_1 _08791_ (.A(_03641_),
    .B(_03642_),
    .C(_03645_),
    .D(_03648_),
    .Y(_03649_));
 sg13g2_nand2_1 _08792_ (.Y(_03650_),
    .A(_01876_),
    .B(net191));
 sg13g2_o21ai_1 _08793_ (.B1(_03650_),
    .Y(_00341_),
    .A1(_03542_),
    .A2(_03649_));
 sg13g2_nand2b_1 _08794_ (.Y(_03651_),
    .B(net142),
    .A_N(_00085_));
 sg13g2_nand2b_1 _08795_ (.Y(_03652_),
    .B(net142),
    .A_N(_00081_));
 sg13g2_mux4_1 _08796_ (.S0(net120),
    .A0(_03651_),
    .A1(_03652_),
    .A2(_00086_),
    .A3(_00082_),
    .S1(net327),
    .X(_03653_));
 sg13g2_mux4_1 _08797_ (.S0(net120),
    .A0(_00084_),
    .A1(_00080_),
    .A2(_00083_),
    .A3(_00079_),
    .S1(_03528_),
    .X(_03654_));
 sg13g2_nand2b_1 _08798_ (.Y(_03655_),
    .B(net143),
    .A_N(_00125_));
 sg13g2_nand2b_1 _08799_ (.Y(_03656_),
    .B(net143),
    .A_N(_00121_));
 sg13g2_mux4_1 _08800_ (.S0(net120),
    .A0(_03655_),
    .A1(_03656_),
    .A2(_00126_),
    .A3(_00122_),
    .S1(net327),
    .X(_03657_));
 sg13g2_mux4_1 _08801_ (.S0(net120),
    .A0(_00124_),
    .A1(_00120_),
    .A2(_00123_),
    .A3(_00119_),
    .S1(_03528_),
    .X(_03658_));
 sg13g2_mux4_1 _08802_ (.S0(_03538_),
    .A0(_03653_),
    .A1(_03654_),
    .A2(_03657_),
    .A3(_03658_),
    .S1(net90),
    .X(_03659_));
 sg13g2_nand2b_1 _08803_ (.Y(_03660_),
    .B(_03514_),
    .A_N(_03659_));
 sg13g2_nor2_1 _08804_ (.A(_00157_),
    .B(_03585_),
    .Y(_03661_));
 sg13g2_a221oi_1 _08805_ (.B2(net397),
    .C1(_03661_),
    .B1(_03566_),
    .A1(net385),
    .Y(_03662_),
    .A2(_03559_));
 sg13g2_a22oi_1 _08806_ (.Y(_03663_),
    .B1(net91),
    .B2(_02007_),
    .A2(_03466_),
    .A1(_02572_));
 sg13g2_a221oi_1 _08807_ (.B2(\z80.tv80s.i_tv80_core.PC[6] ),
    .C1(_03560_),
    .B1(_03502_),
    .A1(_02757_),
    .Y(_03664_),
    .A2(_03465_));
 sg13g2_a21o_1 _08808_ (.A2(_03663_),
    .A1(_03569_),
    .B1(_03664_),
    .X(_03665_));
 sg13g2_nand3_1 _08809_ (.B(_03662_),
    .C(_03665_),
    .A(_03660_),
    .Y(_03666_));
 sg13g2_nand2b_1 _08810_ (.Y(_03667_),
    .B(_03666_),
    .A_N(_03542_));
 sg13g2_o21ai_1 _08811_ (.B1(_03667_),
    .Y(_00342_),
    .A1(_01962_),
    .A2(net194));
 sg13g2_nand2b_1 _08812_ (.Y(_03668_),
    .B(net135),
    .A_N(_00093_));
 sg13g2_nand2b_1 _08813_ (.Y(_03669_),
    .B(net135),
    .A_N(_00089_));
 sg13g2_mux4_1 _08814_ (.S0(net121),
    .A0(_03668_),
    .A1(_03669_),
    .A2(_00094_),
    .A3(_00090_),
    .S1(net289),
    .X(_03670_));
 sg13g2_mux4_1 _08815_ (.S0(net121),
    .A0(_00092_),
    .A1(_00088_),
    .A2(_00091_),
    .A3(_00087_),
    .S1(net105),
    .X(_03671_));
 sg13g2_a21oi_1 _08816_ (.A1(_03365_),
    .A2(_03530_),
    .Y(_03672_),
    .B1(net327));
 sg13g2_a21oi_1 _08817_ (.A1(_00134_),
    .A2(_03523_),
    .Y(_03673_),
    .B1(_03672_));
 sg13g2_nor2_1 _08818_ (.A(_00129_),
    .B(_03522_),
    .Y(_03674_));
 sg13g2_a22oi_1 _08819_ (.Y(_03675_),
    .B1(net135),
    .B2(_03674_),
    .A2(_03523_),
    .A1(_02772_));
 sg13g2_nand2_1 _08820_ (.Y(_03676_),
    .A(_03521_),
    .B(_03675_));
 sg13g2_o21ai_1 _08821_ (.B1(_03676_),
    .Y(_03677_),
    .A1(_03521_),
    .A2(_03673_));
 sg13g2_mux4_1 _08822_ (.S0(_03534_),
    .A0(_00132_),
    .A1(_00128_),
    .A2(_00131_),
    .A3(_00127_),
    .S1(_03535_),
    .X(_03678_));
 sg13g2_mux4_1 _08823_ (.S0(_03538_),
    .A0(_03670_),
    .A1(_03671_),
    .A2(_03677_),
    .A3(_03678_),
    .S1(_03569_),
    .X(_03679_));
 sg13g2_inv_1 _08824_ (.Y(_03680_),
    .A(_03679_));
 sg13g2_inv_1 _08825_ (.Y(_03681_),
    .A(_00160_));
 sg13g2_a22oi_1 _08826_ (.Y(_03682_),
    .B1(net78),
    .B2(_03681_),
    .A2(net93),
    .A1(_02593_));
 sg13g2_nand2b_1 _08827_ (.Y(_03683_),
    .B(net77),
    .A_N(_03682_));
 sg13g2_mux2_1 _08828_ (.A0(net349),
    .A1(_02076_),
    .S(_03495_),
    .X(_03684_));
 sg13g2_buf_1 _08829_ (.A(\z80.tv80s.i_tv80_core.PC[7] ),
    .X(_03685_));
 sg13g2_inv_2 _08830_ (.Y(_03686_),
    .A(_03685_));
 sg13g2_nor2_1 _08831_ (.A(_03686_),
    .B(_03496_),
    .Y(_03687_));
 sg13g2_a22oi_1 _08832_ (.Y(_03688_),
    .B1(_03687_),
    .B2(net78),
    .A2(_03684_),
    .A1(_03557_));
 sg13g2_a22oi_1 _08833_ (.Y(_03689_),
    .B1(_03566_),
    .B2(_00697_),
    .A2(_03564_),
    .A1(_02766_));
 sg13g2_nand3_1 _08834_ (.B(_03688_),
    .C(_03689_),
    .A(_03683_),
    .Y(_03690_));
 sg13g2_a21oi_1 _08835_ (.A1(_03514_),
    .A2(_03680_),
    .Y(_03691_),
    .B1(_03690_));
 sg13g2_buf_1 _08836_ (.A(net216),
    .X(_03692_));
 sg13g2_nand2_1 _08837_ (.Y(_03693_),
    .A(net334),
    .B(net190));
 sg13g2_o21ai_1 _08838_ (.B1(_03693_),
    .Y(_00343_),
    .A1(_03542_),
    .A2(_03691_));
 sg13g2_buf_1 _08839_ (.A(net399),
    .X(_03694_));
 sg13g2_nor2_1 _08840_ (.A(_03694_),
    .B(\z80.tv80s.i_tv80_core.BusReq_s ),
    .Y(_03695_));
 sg13g2_a21oi_1 _08841_ (.A1(net328),
    .A2(net5),
    .Y(_00344_),
    .B1(_03695_));
 sg13g2_inv_1 _08842_ (.Y(_03696_),
    .A(_01528_));
 sg13g2_nand2_2 _08843_ (.Y(_03697_),
    .A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .B(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ));
 sg13g2_inv_1 _08844_ (.Y(_03698_),
    .A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ));
 sg13g2_nand2_1 _08845_ (.Y(_03699_),
    .A(_03698_),
    .B(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ));
 sg13g2_or3_1 _08846_ (.A(_01534_),
    .B(_03697_),
    .C(_03699_),
    .X(_03700_));
 sg13g2_buf_2 _08847_ (.A(_03700_),
    .X(_03701_));
 sg13g2_nand2_1 _08848_ (.Y(_03702_),
    .A(net176),
    .B(net382));
 sg13g2_o21ai_1 _08849_ (.B1(_03702_),
    .Y(_03703_),
    .A1(_02101_),
    .A2(_01494_));
 sg13g2_nor4_1 _08850_ (.A(_01749_),
    .B(net296),
    .C(_01879_),
    .D(_03703_),
    .Y(_03704_));
 sg13g2_nor2_1 _08851_ (.A(_01255_),
    .B(_01486_),
    .Y(_03705_));
 sg13g2_o21ai_1 _08852_ (.B1(net333),
    .Y(_03706_),
    .A1(_03704_),
    .A2(_03705_));
 sg13g2_or2_1 _08853_ (.X(_03707_),
    .B(net334),
    .A(net381));
 sg13g2_nand3_1 _08854_ (.B(net374),
    .C(_03707_),
    .A(net255),
    .Y(_03708_));
 sg13g2_or3_1 _08855_ (.A(net255),
    .B(net374),
    .C(_02061_),
    .X(_03709_));
 sg13g2_a22oi_1 _08856_ (.Y(_03710_),
    .B1(_03708_),
    .B2(_03709_),
    .A2(net149),
    .A1(net335));
 sg13g2_xnor2_1 _08857_ (.Y(_03711_),
    .A(net255),
    .B(_02018_));
 sg13g2_nor2_1 _08858_ (.A(net335),
    .B(net149),
    .Y(_03712_));
 sg13g2_a21oi_1 _08859_ (.A1(net381),
    .A2(_03711_),
    .Y(_03713_),
    .B1(_03712_));
 sg13g2_nor2_1 _08860_ (.A(net381),
    .B(_03711_),
    .Y(_03714_));
 sg13g2_nor2_1 _08861_ (.A(_03713_),
    .B(_03714_),
    .Y(_03715_));
 sg13g2_a21oi_1 _08862_ (.A1(net294),
    .A2(net299),
    .Y(_03716_),
    .B1(net297));
 sg13g2_buf_1 _08863_ (.A(_03716_),
    .X(_03717_));
 sg13g2_o21ai_1 _08864_ (.B1(_03717_),
    .Y(_03718_),
    .A1(_03710_),
    .A2(_03715_));
 sg13g2_or4_1 _08865_ (.A(net294),
    .B(net255),
    .C(_03710_),
    .D(_03715_),
    .X(_03719_));
 sg13g2_a21o_1 _08866_ (.A2(_03719_),
    .A1(_03718_),
    .B1(net333),
    .X(_03720_));
 sg13g2_nand2_1 _08867_ (.Y(_03721_),
    .A(net376),
    .B(_01907_));
 sg13g2_nand2_1 _08868_ (.Y(_03722_),
    .A(_01915_),
    .B(_01907_));
 sg13g2_xnor2_1 _08869_ (.Y(_03723_),
    .A(_01494_),
    .B(_03722_));
 sg13g2_nand2_1 _08870_ (.Y(_03724_),
    .A(_01921_),
    .B(_03723_));
 sg13g2_o21ai_1 _08871_ (.B1(_03724_),
    .Y(_03725_),
    .A1(_01921_),
    .A2(_03721_));
 sg13g2_nor2b_1 _08872_ (.A(_02021_),
    .B_N(_02025_),
    .Y(_03726_));
 sg13g2_o21ai_1 _08873_ (.B1(net337),
    .Y(_03727_),
    .A1(_01927_),
    .A2(_03726_));
 sg13g2_o21ai_1 _08874_ (.B1(_03727_),
    .Y(_03728_),
    .A1(net337),
    .A2(_03725_));
 sg13g2_a21o_1 _08875_ (.A2(_03728_),
    .A1(_01255_),
    .B1(_01511_),
    .X(_03729_));
 sg13g2_nand2_1 _08876_ (.Y(_03730_),
    .A(_00845_),
    .B(_01156_));
 sg13g2_nor4_2 _08877_ (.A(_03102_),
    .B(_02116_),
    .C(_02363_),
    .Y(_03731_),
    .D(_03730_));
 sg13g2_nor2_1 _08878_ (.A(_00191_),
    .B(_03731_),
    .Y(_03732_));
 sg13g2_nor2_1 _08879_ (.A(_01712_),
    .B(_03732_),
    .Y(_03733_));
 sg13g2_buf_1 _08880_ (.A(_03733_),
    .X(_03734_));
 sg13g2_nor2_1 _08881_ (.A(\z80.tv80s.i_tv80_core.PreserveC_r ),
    .B(_03734_),
    .Y(_03735_));
 sg13g2_and4_1 _08882_ (.A(_03706_),
    .B(_03720_),
    .C(_03729_),
    .D(_03735_),
    .X(_03736_));
 sg13g2_nor3_1 _08883_ (.A(_00780_),
    .B(net268),
    .C(_01059_),
    .Y(_03737_));
 sg13g2_nand2b_1 _08884_ (.Y(_03738_),
    .B(_01422_),
    .A_N(_03737_));
 sg13g2_inv_1 _08885_ (.Y(_03739_),
    .A(_01588_));
 sg13g2_nor2_1 _08886_ (.A(_03739_),
    .B(_02298_),
    .Y(_03740_));
 sg13g2_nand2_1 _08887_ (.Y(_03741_),
    .A(_00995_),
    .B(_03740_));
 sg13g2_a21oi_1 _08888_ (.A1(net391),
    .A2(_03738_),
    .Y(_03742_),
    .B1(_03741_));
 sg13g2_mux2_1 _08889_ (.A0(_03742_),
    .A1(\z80.tv80s.i_tv80_core.Fp[0] ),
    .S(net129),
    .X(_03743_));
 sg13g2_nand3_1 _08890_ (.B(_00888_),
    .C(_01054_),
    .A(net262),
    .Y(_03744_));
 sg13g2_nand3_1 _08891_ (.B(_03744_),
    .C(_03740_),
    .A(_00995_),
    .Y(_03745_));
 sg13g2_nand2b_1 _08892_ (.Y(_03746_),
    .B(_03745_),
    .A_N(net129));
 sg13g2_nand2_1 _08893_ (.Y(_03747_),
    .A(net178),
    .B(_03746_));
 sg13g2_a221oi_1 _08894_ (.B2(net391),
    .C1(_03735_),
    .B1(_03747_),
    .A1(_01603_),
    .Y(_03748_),
    .A2(_03743_));
 sg13g2_o21ai_1 _08895_ (.B1(_03701_),
    .Y(_03749_),
    .A1(_03736_),
    .A2(_03748_));
 sg13g2_o21ai_1 _08896_ (.B1(_03749_),
    .Y(_03750_),
    .A1(_03696_),
    .A2(_03701_));
 sg13g2_mux2_1 _08897_ (.A0(_00237_),
    .A1(_03750_),
    .S(net227),
    .X(_00345_));
 sg13g2_nor3_2 _08898_ (.A(_01534_),
    .B(_03697_),
    .C(_03699_),
    .Y(_03751_));
 sg13g2_inv_1 _08899_ (.Y(_03752_),
    .A(_00995_));
 sg13g2_nor4_1 _08900_ (.A(_02159_),
    .B(net104),
    .C(net228),
    .D(_01335_),
    .Y(_03753_));
 sg13g2_buf_2 _08901_ (.A(_03753_),
    .X(_03754_));
 sg13g2_buf_1 _08902_ (.A(_00135_),
    .X(_03755_));
 sg13g2_nor4_2 _08903_ (.A(_03755_),
    .B(net284),
    .C(net182),
    .Y(_03756_),
    .D(_02248_));
 sg13g2_nor3_1 _08904_ (.A(_03751_),
    .B(_03754_),
    .C(_03756_),
    .Y(_03757_));
 sg13g2_buf_1 _08905_ (.A(_03734_),
    .X(_03758_));
 sg13g2_or2_1 _08906_ (.X(_03759_),
    .B(_03717_),
    .A(_01662_));
 sg13g2_a22oi_1 _08907_ (.Y(_03760_),
    .B1(_03759_),
    .B2(_01843_),
    .A2(_03717_),
    .A1(_01487_));
 sg13g2_a21oi_1 _08908_ (.A1(\z80.tv80s.i_tv80_core.Fp[1] ),
    .A2(net130),
    .Y(_03761_),
    .B1(_01592_));
 sg13g2_o21ai_1 _08909_ (.B1(_01834_),
    .Y(_03762_),
    .A1(net198),
    .A2(_03761_));
 sg13g2_nand2b_1 _08910_ (.Y(_03763_),
    .B(net130),
    .A_N(\z80.tv80s.i_tv80_core.Fp[1] ));
 sg13g2_o21ai_1 _08911_ (.B1(_03763_),
    .Y(_03764_),
    .A1(net129),
    .A2(_03741_));
 sg13g2_nand2_1 _08912_ (.Y(_03765_),
    .A(net178),
    .B(_03764_));
 sg13g2_nand4_1 _08913_ (.B(net118),
    .C(_03762_),
    .A(_01543_),
    .Y(_03766_),
    .D(_03765_));
 sg13g2_o21ai_1 _08914_ (.B1(_03766_),
    .Y(_03767_),
    .A1(net118),
    .A2(_03760_));
 sg13g2_a221oi_1 _08915_ (.B2(_03767_),
    .C1(_01267_),
    .B1(_03757_),
    .A1(_01681_),
    .Y(_03768_),
    .A2(_03751_));
 sg13g2_a21o_1 _08916_ (.A2(net197),
    .A1(_00238_),
    .B1(_03768_),
    .X(_00346_));
 sg13g2_nand2_2 _08917_ (.Y(_03769_),
    .A(net333),
    .B(_03717_));
 sg13g2_xnor2_1 _08918_ (.Y(_03770_),
    .A(_01468_),
    .B(_01661_));
 sg13g2_xnor2_1 _08919_ (.Y(_03771_),
    .A(_01720_),
    .B(_03770_));
 sg13g2_xnor2_1 _08920_ (.Y(_03772_),
    .A(_01777_),
    .B(_03771_));
 sg13g2_xnor2_1 _08921_ (.Y(_03773_),
    .A(_01846_),
    .B(_03772_));
 sg13g2_xnor2_1 _08922_ (.Y(_03774_),
    .A(_03728_),
    .B(_03773_));
 sg13g2_xnor2_1 _08923_ (.Y(_03775_),
    .A(_02034_),
    .B(_03774_));
 sg13g2_xnor2_1 _08924_ (.Y(_03776_),
    .A(_01934_),
    .B(_01991_));
 sg13g2_xnor2_1 _08925_ (.Y(_03777_),
    .A(_03775_),
    .B(_03776_));
 sg13g2_xor2_1 _08926_ (.B(_01650_),
    .A(_01499_),
    .X(_03778_));
 sg13g2_xnor2_1 _08927_ (.Y(_03779_),
    .A(_01519_),
    .B(_01648_));
 sg13g2_nor2_1 _08928_ (.A(_01514_),
    .B(_03779_),
    .Y(_03780_));
 sg13g2_a21oi_1 _08929_ (.A1(net296),
    .A2(_03778_),
    .Y(_03781_),
    .B1(_03780_));
 sg13g2_xnor2_1 _08930_ (.Y(_03782_),
    .A(_01722_),
    .B(_01780_));
 sg13g2_xnor2_1 _08931_ (.Y(_03783_),
    .A(net336),
    .B(_01914_));
 sg13g2_xnor2_1 _08932_ (.Y(_03784_),
    .A(_01994_),
    .B(net338));
 sg13g2_xnor2_1 _08933_ (.Y(_03785_),
    .A(_03783_),
    .B(_03784_));
 sg13g2_xnor2_1 _08934_ (.Y(_03786_),
    .A(_03782_),
    .B(_03785_));
 sg13g2_xnor2_1 _08935_ (.Y(_03787_),
    .A(_03781_),
    .B(_03786_));
 sg13g2_xnor2_1 _08936_ (.Y(_03788_),
    .A(net382),
    .B(_01496_));
 sg13g2_xor2_1 _08937_ (.B(_01911_),
    .A(net381),
    .X(_03789_));
 sg13g2_nand2_1 _08938_ (.Y(_03790_),
    .A(net195),
    .B(_03789_));
 sg13g2_o21ai_1 _08939_ (.B1(_03790_),
    .Y(_03791_),
    .A1(_01896_),
    .A2(_03788_));
 sg13g2_xnor2_1 _08940_ (.Y(_03792_),
    .A(_01850_),
    .B(_03791_));
 sg13g2_xnor2_1 _08941_ (.Y(_03793_),
    .A(_01723_),
    .B(_01782_));
 sg13g2_xnor2_1 _08942_ (.Y(_03794_),
    .A(_01492_),
    .B(_01670_));
 sg13g2_xnor2_1 _08943_ (.Y(_03795_),
    .A(_03793_),
    .B(_03794_));
 sg13g2_xnor2_1 _08944_ (.Y(_03796_),
    .A(_02044_),
    .B(_03795_));
 sg13g2_xnor2_1 _08945_ (.Y(_03797_),
    .A(_03792_),
    .B(_03796_));
 sg13g2_nand2_1 _08946_ (.Y(_03798_),
    .A(_01230_),
    .B(_00685_));
 sg13g2_o21ai_1 _08947_ (.B1(_03798_),
    .Y(_03799_),
    .A1(_01230_),
    .A2(_03797_));
 sg13g2_nor2_1 _08948_ (.A(_01648_),
    .B(_01666_),
    .Y(_03800_));
 sg13g2_o21ai_1 _08949_ (.B1(_01712_),
    .Y(_03801_),
    .A1(_01519_),
    .A2(_01073_));
 sg13g2_inv_1 _08950_ (.Y(_03802_),
    .A(_01499_));
 sg13g2_and2_1 _08951_ (.A(net339),
    .B(_00202_),
    .X(_03803_));
 sg13g2_a21oi_1 _08952_ (.A1(net317),
    .A2(_00206_),
    .Y(_03804_),
    .B1(_03803_));
 sg13g2_a22oi_1 _08953_ (.Y(_03805_),
    .B1(_03804_),
    .B2(_00694_),
    .A2(_01847_),
    .A1(_03802_));
 sg13g2_o21ai_1 _08954_ (.B1(_03805_),
    .Y(_03806_),
    .A1(_01778_),
    .A2(_01789_));
 sg13g2_nor2_1 _08955_ (.A(_01650_),
    .B(_01897_),
    .Y(_03807_));
 sg13g2_or4_1 _08956_ (.A(_03800_),
    .B(_03801_),
    .C(_03806_),
    .D(_03807_),
    .X(_03808_));
 sg13g2_o21ai_1 _08957_ (.B1(_03769_),
    .Y(_03809_),
    .A1(_02037_),
    .A2(_03808_));
 sg13g2_a221oi_1 _08958_ (.B2(_01490_),
    .C1(_03809_),
    .B1(_03799_),
    .A1(_01507_),
    .Y(_03810_),
    .A2(_03787_));
 sg13g2_o21ai_1 _08959_ (.B1(_03810_),
    .Y(_03811_),
    .A1(_01511_),
    .A2(_03777_));
 sg13g2_nand2_1 _08960_ (.Y(_03812_),
    .A(_01487_),
    .B(_02872_));
 sg13g2_nand2b_1 _08961_ (.Y(_03813_),
    .B(_03812_),
    .A_N(_03811_));
 sg13g2_a22oi_1 _08962_ (.Y(_03814_),
    .B1(_03813_),
    .B2(_00685_),
    .A2(_03811_),
    .A1(_03769_));
 sg13g2_xor2_1 _08963_ (.B(_02070_),
    .A(_01894_),
    .X(_03815_));
 sg13g2_xnor2_1 _08964_ (.Y(_03816_),
    .A(_01483_),
    .B(_03815_));
 sg13g2_xnor2_1 _08965_ (.Y(_03817_),
    .A(_01647_),
    .B(_03816_));
 sg13g2_xnor2_1 _08966_ (.Y(_03818_),
    .A(_01710_),
    .B(_03817_));
 sg13g2_xnor2_1 _08967_ (.Y(_03819_),
    .A(_01766_),
    .B(_03818_));
 sg13g2_xnor2_1 _08968_ (.Y(_03820_),
    .A(_01833_),
    .B(_03819_));
 sg13g2_xnor2_1 _08969_ (.Y(_03821_),
    .A(_01981_),
    .B(_03820_));
 sg13g2_nand2_1 _08970_ (.Y(_03822_),
    .A(net381),
    .B(_02018_));
 sg13g2_nand2_1 _08971_ (.Y(_03823_),
    .A(_01962_),
    .B(net149));
 sg13g2_o21ai_1 _08972_ (.B1(net335),
    .Y(_03824_),
    .A1(_01962_),
    .A2(net149));
 sg13g2_nand2_1 _08973_ (.Y(_03825_),
    .A(_03823_),
    .B(_03824_));
 sg13g2_mux2_1 _08974_ (.A0(_03707_),
    .A1(_03822_),
    .S(_03825_),
    .X(_03826_));
 sg13g2_a21o_1 _08975_ (.A2(net149),
    .A1(_01961_),
    .B1(net335),
    .X(_03827_));
 sg13g2_o21ai_1 _08976_ (.B1(_03827_),
    .Y(_03828_),
    .A1(_01961_),
    .A2(net149));
 sg13g2_mux2_1 _08977_ (.A0(_02062_),
    .A1(_02061_),
    .S(_03828_),
    .X(_03829_));
 sg13g2_nor2_1 _08978_ (.A(net255),
    .B(_03829_),
    .Y(_03830_));
 sg13g2_a221oi_1 _08979_ (.B2(net255),
    .C1(_03830_),
    .B1(_03826_),
    .A1(net294),
    .Y(_03831_),
    .A2(_01619_));
 sg13g2_a21oi_1 _08980_ (.A1(_01621_),
    .A2(_03821_),
    .Y(_03832_),
    .B1(_03831_));
 sg13g2_or3_1 _08981_ (.A(net333),
    .B(_02872_),
    .C(_03832_),
    .X(_03833_));
 sg13g2_a21o_1 _08982_ (.A2(_03833_),
    .A1(_03814_),
    .B1(_03758_),
    .X(_03834_));
 sg13g2_nor2_1 _08983_ (.A(net266),
    .B(_02251_),
    .Y(_03835_));
 sg13g2_nand2_2 _08984_ (.Y(_03836_),
    .A(_01594_),
    .B(_01575_));
 sg13g2_mux2_1 _08985_ (.A0(\z80.tv80s.i_tv80_core.Fp[2] ),
    .A1(_00685_),
    .S(_03836_),
    .X(_03837_));
 sg13g2_mux2_1 _08986_ (.A0(\z80.tv80s.i_tv80_core.IntE_FF2 ),
    .A1(_03837_),
    .S(_01542_),
    .X(_03838_));
 sg13g2_a221oi_1 _08987_ (.B2(_03838_),
    .C1(_03754_),
    .B1(net118),
    .A1(_01191_),
    .Y(_03839_),
    .A2(_03835_));
 sg13g2_xor2_1 _08988_ (.B(net388),
    .A(_01395_),
    .X(_03840_));
 sg13g2_xnor2_1 _08989_ (.Y(_03841_),
    .A(net350),
    .B(_01394_));
 sg13g2_xnor2_1 _08990_ (.Y(_03842_),
    .A(_03840_),
    .B(_03841_));
 sg13g2_xnor2_1 _08991_ (.Y(_03843_),
    .A(_01399_),
    .B(_01401_));
 sg13g2_xnor2_1 _08992_ (.Y(_03844_),
    .A(net387),
    .B(_01398_));
 sg13g2_xnor2_1 _08993_ (.Y(_03845_),
    .A(_03843_),
    .B(_03844_));
 sg13g2_xnor2_1 _08994_ (.Y(_03846_),
    .A(_03842_),
    .B(_03845_));
 sg13g2_nor4_1 _08995_ (.A(net237),
    .B(\z80.tv80s.i_tv80_core.IncDecZ ),
    .C(net182),
    .D(_02248_),
    .Y(_03847_));
 sg13g2_a221oi_1 _08996_ (.B2(_03754_),
    .C1(_03847_),
    .B1(_03846_),
    .A1(_03834_),
    .Y(_03848_),
    .A2(_03839_));
 sg13g2_nand2_1 _08997_ (.Y(_03849_),
    .A(net264),
    .B(_03701_));
 sg13g2_buf_1 _08998_ (.A(net225),
    .X(_03850_));
 sg13g2_nor2_1 _08999_ (.A(_01266_),
    .B(_03701_),
    .Y(_03851_));
 sg13g2_a22oi_1 _09000_ (.Y(_03852_),
    .B1(_01735_),
    .B2(_03851_),
    .A2(net189),
    .A1(_00239_));
 sg13g2_o21ai_1 _09001_ (.B1(_03852_),
    .Y(_00347_),
    .A1(_03848_),
    .A2(_03849_));
 sg13g2_nor3_1 _09002_ (.A(_01340_),
    .B(_01712_),
    .C(_03732_),
    .Y(_03853_));
 sg13g2_nor2_1 _09003_ (.A(_03599_),
    .B(net115),
    .Y(_03854_));
 sg13g2_nand2b_1 _09004_ (.Y(_03855_),
    .B(_00995_),
    .A_N(_01591_));
 sg13g2_o21ai_1 _09005_ (.B1(_01803_),
    .Y(_03856_),
    .A1(_03739_),
    .A2(_02298_));
 sg13g2_a21oi_1 _09006_ (.A1(_03599_),
    .A2(_03855_),
    .Y(_03857_),
    .B1(_03856_));
 sg13g2_nand2b_1 _09007_ (.Y(_03858_),
    .B(_01591_),
    .A_N(_03599_));
 sg13g2_a21oi_1 _09008_ (.A1(_03741_),
    .A2(_03858_),
    .Y(_03859_),
    .B1(_01803_));
 sg13g2_nor4_1 _09009_ (.A(net129),
    .B(_03854_),
    .C(_03857_),
    .D(_03859_),
    .Y(_03860_));
 sg13g2_a21oi_1 _09010_ (.A1(\z80.tv80s.i_tv80_core.Fp[3] ),
    .A2(net129),
    .Y(_03861_),
    .B1(_03860_));
 sg13g2_nor2_1 _09011_ (.A(_03734_),
    .B(_03769_),
    .Y(_03862_));
 sg13g2_a21oi_1 _09012_ (.A1(net198),
    .A2(_03734_),
    .Y(_03863_),
    .B1(_03862_));
 sg13g2_or2_1 _09013_ (.X(_03864_),
    .B(_01619_),
    .A(_00208_));
 sg13g2_buf_1 _09014_ (.A(_03864_),
    .X(_03865_));
 sg13g2_mux2_1 _09015_ (.A0(_01778_),
    .A1(_01766_),
    .S(_03865_),
    .X(_03866_));
 sg13g2_and2_1 _09016_ (.A(_02241_),
    .B(_03717_),
    .X(_03867_));
 sg13g2_buf_1 _09017_ (.A(_03867_),
    .X(_03868_));
 sg13g2_nor3_1 _09018_ (.A(_01778_),
    .B(net175),
    .C(_01665_),
    .Y(_03869_));
 sg13g2_nor4_1 _09019_ (.A(_01787_),
    .B(_03734_),
    .C(_03868_),
    .D(_03869_),
    .Y(_03870_));
 sg13g2_o21ai_1 _09020_ (.B1(_03870_),
    .Y(_03871_),
    .A1(net333),
    .A2(_03866_));
 sg13g2_o21ai_1 _09021_ (.B1(_03871_),
    .Y(_03872_),
    .A1(_03599_),
    .A2(_03863_));
 sg13g2_a21oi_1 _09022_ (.A1(_03853_),
    .A2(_03861_),
    .Y(_03873_),
    .B1(_03872_));
 sg13g2_inv_1 _09023_ (.Y(_03874_),
    .A(_03756_));
 sg13g2_mux2_1 _09024_ (.A0(_01795_),
    .A1(_03873_),
    .S(_03874_),
    .X(_03875_));
 sg13g2_a22oi_1 _09025_ (.Y(_03876_),
    .B1(_01802_),
    .B2(_03851_),
    .A2(net189),
    .A1(_00240_));
 sg13g2_o21ai_1 _09026_ (.B1(_03876_),
    .Y(_00348_),
    .A1(_03849_),
    .A2(_03875_));
 sg13g2_inv_1 _09027_ (.Y(_03877_),
    .A(_01863_));
 sg13g2_nand2_1 _09028_ (.Y(_03878_),
    .A(_01654_),
    .B(net179));
 sg13g2_nand2_1 _09029_ (.Y(_03879_),
    .A(\z80.tv80s.i_tv80_core.Fp[4] ),
    .B(_01600_));
 sg13g2_and3_1 _09030_ (.X(_03880_),
    .A(_01654_),
    .B(_03855_),
    .C(_03745_));
 sg13g2_or3_1 _09031_ (.A(net130),
    .B(_03742_),
    .C(_03880_),
    .X(_03881_));
 sg13g2_nand3_1 _09032_ (.B(_03879_),
    .C(_03881_),
    .A(net178),
    .Y(_03882_));
 sg13g2_nand3_1 _09033_ (.B(_03878_),
    .C(_03882_),
    .A(_01543_),
    .Y(_03883_));
 sg13g2_or2_1 _09034_ (.X(_03884_),
    .B(_00208_),
    .A(net296));
 sg13g2_o21ai_1 _09035_ (.B1(_03884_),
    .Y(_03885_),
    .A1(net294),
    .A2(_01819_));
 sg13g2_a22oi_1 _09036_ (.Y(_03886_),
    .B1(_03885_),
    .B2(net297),
    .A2(_03717_),
    .A1(_01819_));
 sg13g2_nand2b_1 _09037_ (.Y(_03887_),
    .B(_01696_),
    .A_N(_01492_));
 sg13g2_nand3_1 _09038_ (.B(_01653_),
    .C(_03887_),
    .A(_01843_),
    .Y(_03888_));
 sg13g2_nand3_1 _09039_ (.B(_01834_),
    .C(_01769_),
    .A(_01760_),
    .Y(_03889_));
 sg13g2_o21ai_1 _09040_ (.B1(_03889_),
    .Y(_03890_),
    .A1(_01760_),
    .A2(_03888_));
 sg13g2_a221oi_1 _09041_ (.B2(_01662_),
    .C1(_01712_),
    .B1(_03890_),
    .A1(_01653_),
    .Y(_03891_),
    .A2(_03868_));
 sg13g2_o21ai_1 _09042_ (.B1(_03891_),
    .Y(_03892_),
    .A1(net333),
    .A2(_03886_));
 sg13g2_nor2_1 _09043_ (.A(_03758_),
    .B(_03892_),
    .Y(_03893_));
 sg13g2_a21oi_1 _09044_ (.A1(net118),
    .A2(_03883_),
    .Y(_03894_),
    .B1(_03893_));
 sg13g2_a221oi_1 _09045_ (.B2(_03894_),
    .C1(net202),
    .B1(_03757_),
    .A1(_03877_),
    .Y(_03895_),
    .A2(_03751_));
 sg13g2_a21o_1 _09046_ (.A2(net197),
    .A1(_00241_),
    .B1(_03895_),
    .X(_00349_));
 sg13g2_nor2_1 _09047_ (.A(_03643_),
    .B(net115),
    .Y(_03896_));
 sg13g2_o21ai_1 _09048_ (.B1(_01948_),
    .Y(_03897_),
    .A1(_03739_),
    .A2(_02298_));
 sg13g2_a21oi_1 _09049_ (.A1(_03643_),
    .A2(_03855_),
    .Y(_03898_),
    .B1(_03897_));
 sg13g2_nand2b_1 _09050_ (.Y(_03899_),
    .B(_01591_),
    .A_N(_03643_));
 sg13g2_a21oi_1 _09051_ (.A1(_03741_),
    .A2(_03899_),
    .Y(_03900_),
    .B1(net375));
 sg13g2_nor4_1 _09052_ (.A(net130),
    .B(_03896_),
    .C(_03898_),
    .D(_03900_),
    .Y(_03901_));
 sg13g2_a21oi_1 _09053_ (.A1(\z80.tv80s.i_tv80_core.Fp[5] ),
    .A2(_01600_),
    .Y(_03902_),
    .B1(_03901_));
 sg13g2_and2_1 _09054_ (.A(_03853_),
    .B(_03902_),
    .X(_03903_));
 sg13g2_nor2_1 _09055_ (.A(_01650_),
    .B(_03865_),
    .Y(_03904_));
 sg13g2_a21oi_1 _09056_ (.A1(_01895_),
    .A2(_03865_),
    .Y(_03905_),
    .B1(_03904_));
 sg13g2_nor3_1 _09057_ (.A(_01650_),
    .B(net175),
    .C(_01665_),
    .Y(_03906_));
 sg13g2_nor3_1 _09058_ (.A(_03734_),
    .B(_03868_),
    .C(_03906_),
    .Y(_03907_));
 sg13g2_and2_1 _09059_ (.A(_01939_),
    .B(_03907_),
    .X(_03908_));
 sg13g2_o21ai_1 _09060_ (.B1(_03908_),
    .Y(_03909_),
    .A1(_02241_),
    .A2(_03905_));
 sg13g2_o21ai_1 _09061_ (.B1(_03909_),
    .Y(_03910_),
    .A1(_03643_),
    .A2(_03863_));
 sg13g2_nor3_1 _09062_ (.A(_03756_),
    .B(_03903_),
    .C(_03910_),
    .Y(_03911_));
 sg13g2_o21ai_1 _09063_ (.B1(_03701_),
    .Y(_03912_),
    .A1(_01677_),
    .A2(_03874_));
 sg13g2_nand3_1 _09064_ (.B(_01946_),
    .C(_03751_),
    .A(_01943_),
    .Y(_03913_));
 sg13g2_o21ai_1 _09065_ (.B1(_03913_),
    .Y(_03914_),
    .A1(_03911_),
    .A2(_03912_));
 sg13g2_mux2_1 _09066_ (.A0(_00242_),
    .A1(_03914_),
    .S(net227),
    .X(_00350_));
 sg13g2_inv_1 _09067_ (.Y(_03915_),
    .A(_01661_));
 sg13g2_nand4_1 _09068_ (.B(_01662_),
    .C(_03915_),
    .A(net382),
    .Y(_03916_),
    .D(_01720_));
 sg13g2_nor2b_1 _09069_ (.A(_03916_),
    .B_N(_01777_),
    .Y(_03917_));
 sg13g2_nand4_1 _09070_ (.B(_01991_),
    .C(_02034_),
    .A(_01846_),
    .Y(_03918_),
    .D(_03917_));
 sg13g2_a22oi_1 _09071_ (.Y(_03919_),
    .B1(_01995_),
    .B2(_01911_),
    .A2(_01724_),
    .A1(_01464_));
 sg13g2_nand4_1 _09072_ (.B(_01723_),
    .C(_01782_),
    .A(_01670_),
    .Y(_03920_),
    .D(net377));
 sg13g2_nor4_1 _09073_ (.A(net359),
    .B(_01497_),
    .C(_03919_),
    .D(_03920_),
    .Y(_03921_));
 sg13g2_a22oi_1 _09074_ (.Y(_03922_),
    .B1(_02044_),
    .B2(_03921_),
    .A2(net397),
    .A1(net301));
 sg13g2_nor2_1 _09075_ (.A(_01935_),
    .B(_03922_),
    .Y(_03923_));
 sg13g2_a22oi_1 _09076_ (.Y(_03924_),
    .B1(_01651_),
    .B2(_00206_),
    .A2(_01649_),
    .A1(_00202_));
 sg13g2_mux2_1 _09077_ (.A0(_01519_),
    .A1(_01499_),
    .S(net296),
    .X(_03925_));
 sg13g2_nor2_1 _09078_ (.A(_01825_),
    .B(_01914_),
    .Y(_03926_));
 sg13g2_nand4_1 _09079_ (.B(_01925_),
    .C(_03925_),
    .A(_01780_),
    .Y(_03927_),
    .D(_03926_));
 sg13g2_nor3_1 _09080_ (.A(_01508_),
    .B(_03924_),
    .C(_03927_),
    .Y(_03928_));
 sg13g2_nor3_1 _09081_ (.A(_03809_),
    .B(_03923_),
    .C(_03928_),
    .Y(_03929_));
 sg13g2_o21ai_1 _09082_ (.B1(_03929_),
    .Y(_03930_),
    .A1(_01934_),
    .A2(_03918_));
 sg13g2_a21oi_1 _09083_ (.A1(_03769_),
    .A2(_03930_),
    .Y(_03931_),
    .B1(_00684_));
 sg13g2_nor2b_1 _09084_ (.A(_03930_),
    .B_N(_03812_),
    .Y(_03932_));
 sg13g2_nor2_1 _09085_ (.A(\z80.tv80s.i_tv80_core.Z16_r ),
    .B(_02872_),
    .Y(_03933_));
 sg13g2_o21ai_1 _09086_ (.B1(_01487_),
    .Y(_03934_),
    .A1(_00684_),
    .A2(_03933_));
 sg13g2_nor3_1 _09087_ (.A(_01484_),
    .B(_01647_),
    .C(_03934_),
    .Y(_03935_));
 sg13g2_nand3_1 _09088_ (.B(_01766_),
    .C(_03935_),
    .A(_01710_),
    .Y(_03936_));
 sg13g2_nor4_1 _09089_ (.A(_01833_),
    .B(_01981_),
    .C(_02071_),
    .D(_03936_),
    .Y(_03937_));
 sg13g2_nand2b_1 _09090_ (.Y(_03938_),
    .B(_03937_),
    .A_N(_01895_));
 sg13g2_o21ai_1 _09091_ (.B1(_03938_),
    .Y(_03939_),
    .A1(_03931_),
    .A2(_03932_));
 sg13g2_nor4_1 _09092_ (.A(_01868_),
    .B(_01953_),
    .C(_02011_),
    .D(_02080_),
    .Y(_03940_));
 sg13g2_nor4_1 _09093_ (.A(_01605_),
    .B(\z80.tv80s.i_tv80_core.I[1] ),
    .C(_01740_),
    .D(_01807_),
    .Y(_03941_));
 sg13g2_a21oi_1 _09094_ (.A1(_03940_),
    .A2(_03941_),
    .Y(_03942_),
    .B1(_01542_));
 sg13g2_mux2_1 _09095_ (.A0(\z80.tv80s.i_tv80_core.Fp[6] ),
    .A1(net397),
    .S(_03836_),
    .X(_03943_));
 sg13g2_nor2b_1 _09096_ (.A(_03943_),
    .B_N(_01542_),
    .Y(_03944_));
 sg13g2_o21ai_1 _09097_ (.B1(net118),
    .Y(_03945_),
    .A1(_03942_),
    .A2(_03944_));
 sg13g2_o21ai_1 _09098_ (.B1(_03945_),
    .Y(_03946_),
    .A1(net118),
    .A2(_03939_));
 sg13g2_nor4_1 _09099_ (.A(_01397_),
    .B(_01398_),
    .C(net385),
    .D(net349),
    .Y(_03947_));
 sg13g2_nor4_1 _09100_ (.A(_01393_),
    .B(_01394_),
    .C(net389),
    .D(_01396_),
    .Y(_03948_));
 sg13g2_nand3_1 _09101_ (.B(_03947_),
    .C(_03948_),
    .A(_03754_),
    .Y(_03949_));
 sg13g2_o21ai_1 _09102_ (.B1(_03949_),
    .Y(_03950_),
    .A1(_03754_),
    .A2(_03946_));
 sg13g2_mux2_1 _09103_ (.A0(_02006_),
    .A1(_03950_),
    .S(_03701_),
    .X(_03951_));
 sg13g2_nand2_1 _09104_ (.Y(_03952_),
    .A(_00243_),
    .B(_03692_));
 sg13g2_o21ai_1 _09105_ (.B1(_03952_),
    .Y(_00351_),
    .A1(net177),
    .A2(_03951_));
 sg13g2_nand2b_1 _09106_ (.Y(_03953_),
    .B(_02872_),
    .A_N(_00697_));
 sg13g2_o21ai_1 _09107_ (.B1(_03953_),
    .Y(_03954_),
    .A1(_02872_),
    .A2(_02071_));
 sg13g2_o21ai_1 _09108_ (.B1(_03769_),
    .Y(_03955_),
    .A1(net305),
    .A2(_01935_));
 sg13g2_a221oi_1 _09109_ (.B2(_00697_),
    .C1(_02039_),
    .B1(_03955_),
    .A1(net260),
    .Y(_03956_),
    .A2(_02045_));
 sg13g2_o21ai_1 _09110_ (.B1(_03956_),
    .Y(_03957_),
    .A1(net333),
    .A2(_03954_));
 sg13g2_nor2_1 _09111_ (.A(_02080_),
    .B(net155),
    .Y(_03958_));
 sg13g2_mux2_1 _09112_ (.A0(\z80.tv80s.i_tv80_core.Fp[7] ),
    .A1(_00697_),
    .S(_03836_),
    .X(_03959_));
 sg13g2_nor2b_1 _09113_ (.A(_03959_),
    .B_N(_01542_),
    .Y(_03960_));
 sg13g2_o21ai_1 _09114_ (.B1(net118),
    .Y(_03961_),
    .A1(_03958_),
    .A2(_03960_));
 sg13g2_o21ai_1 _09115_ (.B1(_03961_),
    .Y(_03962_),
    .A1(net118),
    .A2(_03957_));
 sg13g2_nand2_1 _09116_ (.Y(_03963_),
    .A(_01401_),
    .B(_03754_));
 sg13g2_o21ai_1 _09117_ (.B1(_03963_),
    .Y(_03964_),
    .A1(_03754_),
    .A2(_03962_));
 sg13g2_a22oi_1 _09118_ (.Y(_03965_),
    .B1(_02075_),
    .B2(_03851_),
    .A2(net189),
    .A1(_00244_));
 sg13g2_o21ai_1 _09119_ (.B1(_03965_),
    .Y(_00352_),
    .A1(_03849_),
    .A2(_03964_));
 sg13g2_nand2_1 _09120_ (.Y(_03966_),
    .A(_00245_),
    .B(net122));
 sg13g2_o21ai_1 _09121_ (.B1(_03966_),
    .Y(_00353_),
    .A1(net391),
    .A2(net124));
 sg13g2_nand2_1 _09122_ (.Y(_03967_),
    .A(_00246_),
    .B(net122));
 sg13g2_o21ai_1 _09123_ (.B1(_03967_),
    .Y(_00354_),
    .A1(net337),
    .A2(net124));
 sg13g2_nand2_1 _09124_ (.Y(_03968_),
    .A(_00247_),
    .B(net122));
 sg13g2_o21ai_1 _09125_ (.B1(_03968_),
    .Y(_00355_),
    .A1(_00685_),
    .A2(net123));
 sg13g2_nand2_1 _09126_ (.Y(_03969_),
    .A(_00248_),
    .B(net122));
 sg13g2_o21ai_1 _09127_ (.B1(_03969_),
    .Y(_00356_),
    .A1(_03599_),
    .A2(net123));
 sg13g2_nand2_1 _09128_ (.Y(_03970_),
    .A(_00249_),
    .B(net122));
 sg13g2_o21ai_1 _09129_ (.B1(_03970_),
    .Y(_00357_),
    .A1(_01653_),
    .A2(net123));
 sg13g2_nand2_1 _09130_ (.Y(_03971_),
    .A(_00250_),
    .B(net122));
 sg13g2_o21ai_1 _09131_ (.B1(_03971_),
    .Y(_00358_),
    .A1(_03643_),
    .A2(net123));
 sg13g2_nand2_1 _09132_ (.Y(_03972_),
    .A(_00251_),
    .B(_02854_));
 sg13g2_o21ai_1 _09133_ (.B1(_03972_),
    .Y(_00359_),
    .A1(net397),
    .A2(net123));
 sg13g2_nand2_1 _09134_ (.Y(_03973_),
    .A(_00252_),
    .B(_02854_));
 sg13g2_o21ai_1 _09135_ (.B1(_03973_),
    .Y(_00360_),
    .A1(_00697_),
    .A2(_02856_));
 sg13g2_inv_1 _09136_ (.Y(_03974_),
    .A(_00035_));
 sg13g2_and2_1 _09137_ (.A(net115),
    .B(_00997_),
    .X(_03975_));
 sg13g2_nand2_1 _09138_ (.Y(_03976_),
    .A(_01085_),
    .B(_01447_));
 sg13g2_nor2b_1 _09139_ (.A(_03976_),
    .B_N(_00999_),
    .Y(_03977_));
 sg13g2_a22oi_1 _09140_ (.Y(_03978_),
    .B1(_03975_),
    .B2(_03977_),
    .A2(_00827_),
    .A1(_03974_));
 sg13g2_nor2_1 _09141_ (.A(net326),
    .B(\z80.tv80s.i_tv80_core.Halt_FF ),
    .Y(_03979_));
 sg13g2_a21oi_1 _09142_ (.A1(net328),
    .A2(_03978_),
    .Y(_00361_),
    .B1(_03979_));
 sg13g2_nor2_1 _09143_ (.A(net326),
    .B(\z80.tv80s.i_tv80_core.INT_s ),
    .Y(_03980_));
 sg13g2_a21oi_1 _09144_ (.A1(_02889_),
    .A2(net3),
    .Y(_00362_),
    .B1(_03980_));
 sg13g2_and2_1 _09145_ (.A(net300),
    .B(net353),
    .X(_03981_));
 sg13g2_o21ai_1 _09146_ (.B1(_01315_),
    .Y(_03982_),
    .A1(net198),
    .A2(_03981_));
 sg13g2_buf_1 _09147_ (.A(_03982_),
    .X(_03983_));
 sg13g2_and2_1 _09148_ (.A(_00825_),
    .B(\z80.tv80s.i_tv80_core.IStatus[2] ),
    .X(_03984_));
 sg13g2_a21oi_1 _09149_ (.A1(_02609_),
    .A2(_03984_),
    .Y(_03985_),
    .B1(net163));
 sg13g2_buf_2 _09150_ (.A(_03985_),
    .X(_03986_));
 sg13g2_nand3b_1 _09151_ (.B(_00016_),
    .C(_02337_),
    .Y(_03987_),
    .A_N(\z80.tv80s.i_tv80_core.Halt_FF ));
 sg13g2_nand2_1 _09152_ (.Y(_03988_),
    .A(_01341_),
    .B(_03987_));
 sg13g2_buf_2 _09153_ (.A(_03988_),
    .X(_03989_));
 sg13g2_nand2_1 _09154_ (.Y(_03990_),
    .A(net6),
    .B(_03989_));
 sg13g2_a22oi_1 _09155_ (.Y(_00363_),
    .B1(_03986_),
    .B2(_03990_),
    .A2(net163),
    .A1(net243));
 sg13g2_nand2_1 _09156_ (.Y(_03991_),
    .A(net7),
    .B(_03989_));
 sg13g2_a22oi_1 _09157_ (.Y(_00364_),
    .B1(_03986_),
    .B2(_03991_),
    .A2(net163),
    .A1(net283));
 sg13g2_nand2_1 _09158_ (.Y(_03992_),
    .A(net8),
    .B(_03989_));
 sg13g2_a22oi_1 _09159_ (.Y(_00365_),
    .B1(_03986_),
    .B2(_03992_),
    .A2(net163),
    .A1(net275));
 sg13g2_nand2_1 _09160_ (.Y(_03993_),
    .A(net9),
    .B(_03989_));
 sg13g2_a22oi_1 _09161_ (.Y(_00366_),
    .B1(_03986_),
    .B2(_03993_),
    .A2(net163),
    .A1(net262));
 sg13g2_nand2_1 _09162_ (.Y(_03994_),
    .A(net10),
    .B(_03989_));
 sg13g2_a22oi_1 _09163_ (.Y(_00367_),
    .B1(_03986_),
    .B2(_03994_),
    .A2(net163),
    .A1(net261));
 sg13g2_nand2_1 _09164_ (.Y(_03995_),
    .A(net11),
    .B(_03989_));
 sg13g2_a22oi_1 _09165_ (.Y(_00368_),
    .B1(_03986_),
    .B2(_03995_),
    .A2(net163),
    .A1(net259));
 sg13g2_nand2_1 _09166_ (.Y(_03996_),
    .A(net12),
    .B(_03989_));
 sg13g2_a22oi_1 _09167_ (.Y(_00369_),
    .B1(_03986_),
    .B2(_03996_),
    .A2(net163),
    .A1(_00978_));
 sg13g2_nand2_1 _09168_ (.Y(_03997_),
    .A(net13),
    .B(_03989_));
 sg13g2_a22oi_1 _09169_ (.Y(_00370_),
    .B1(_03986_),
    .B2(_03997_),
    .A2(_03983_),
    .A1(_00800_));
 sg13g2_nor3_1 _09170_ (.A(net220),
    .B(net266),
    .C(_00890_),
    .Y(_03998_));
 sg13g2_nor3_1 _09171_ (.A(_01307_),
    .B(net263),
    .C(_01608_),
    .Y(_03999_));
 sg13g2_nand2_1 _09172_ (.Y(_04000_),
    .A(_03998_),
    .B(_03999_));
 sg13g2_buf_4 _09173_ (.X(_04001_),
    .A(_04000_));
 sg13g2_mux2_1 _09174_ (.A0(_01545_),
    .A1(_01605_),
    .S(_04001_),
    .X(_00371_));
 sg13g2_mux2_1 _09175_ (.A0(_01683_),
    .A1(\z80.tv80s.i_tv80_core.I[1] ),
    .S(_04001_),
    .X(_00372_));
 sg13g2_mux2_1 _09176_ (.A0(_01736_),
    .A1(_01740_),
    .S(_04001_),
    .X(_00373_));
 sg13g2_mux2_1 _09177_ (.A0(net379),
    .A1(_01807_),
    .S(_04001_),
    .X(_00374_));
 sg13g2_mux2_1 _09178_ (.A0(_01864_),
    .A1(_01868_),
    .S(_04001_),
    .X(_00375_));
 sg13g2_mux2_1 _09179_ (.A0(net375),
    .A1(_01953_),
    .S(_04001_),
    .X(_00376_));
 sg13g2_mux2_1 _09180_ (.A0(_02007_),
    .A1(_02011_),
    .S(_04001_),
    .X(_00377_));
 sg13g2_mux2_1 _09181_ (.A0(_02076_),
    .A1(_02080_),
    .S(_04001_),
    .X(_00378_));
 sg13g2_mux4_1 _09182_ (.S0(_03066_),
    .A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ),
    .S1(net82),
    .X(_04002_));
 sg13g2_mux4_1 _09183_ (.S0(_03066_),
    .A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ),
    .S1(net82),
    .X(_04003_));
 sg13g2_mux2_1 _09184_ (.A0(_04002_),
    .A1(_04003_),
    .S(_03123_),
    .X(_04004_));
 sg13g2_buf_2 _09185_ (.A(_04004_),
    .X(_04005_));
 sg13g2_o21ai_1 _09186_ (.B1(_04005_),
    .Y(_04006_),
    .A1(_03125_),
    .A2(_03173_));
 sg13g2_buf_2 _09187_ (.A(_04006_),
    .X(_04007_));
 sg13g2_a22oi_1 _09188_ (.Y(_04008_),
    .B1(_02098_),
    .B2(_00704_),
    .A2(_02988_),
    .A1(_00820_));
 sg13g2_o21ai_1 _09189_ (.B1(_00882_),
    .Y(_04009_),
    .A1(net282),
    .A2(_04008_));
 sg13g2_nand3_1 _09190_ (.B(_00877_),
    .C(_00823_),
    .A(_00881_),
    .Y(_04010_));
 sg13g2_o21ai_1 _09191_ (.B1(_04010_),
    .Y(_04011_),
    .A1(_00703_),
    .A2(net232));
 sg13g2_nor3_1 _09192_ (.A(_00638_),
    .B(net303),
    .C(_04008_),
    .Y(_04012_));
 sg13g2_a221oi_1 _09193_ (.B2(net273),
    .C1(_04012_),
    .B1(_04011_),
    .A1(_00739_),
    .Y(_04013_),
    .A2(_04009_));
 sg13g2_nand3b_1 _09194_ (.B(net207),
    .C(_00870_),
    .Y(_04014_),
    .A_N(_04013_));
 sg13g2_buf_1 _09195_ (.A(_04014_),
    .X(_04015_));
 sg13g2_nor2_1 _09196_ (.A(net268),
    .B(_01348_),
    .Y(_04016_));
 sg13g2_nor3_1 _09197_ (.A(_00928_),
    .B(_03017_),
    .C(_04016_),
    .Y(_04017_));
 sg13g2_nor2_1 _09198_ (.A(_00638_),
    .B(_02278_),
    .Y(_04018_));
 sg13g2_nand4_1 _09199_ (.B(_00839_),
    .C(_00849_),
    .A(_00837_),
    .Y(_04019_),
    .D(_04018_));
 sg13g2_a21o_1 _09200_ (.A2(_04019_),
    .A1(_04017_),
    .B1(net355),
    .X(_04020_));
 sg13g2_buf_1 _09201_ (.A(_04020_),
    .X(_04021_));
 sg13g2_and2_1 _09202_ (.A(_04015_),
    .B(_04021_),
    .X(_04022_));
 sg13g2_buf_1 _09203_ (.A(_04022_),
    .X(_04023_));
 sg13g2_buf_1 _09204_ (.A(_04023_),
    .X(_04024_));
 sg13g2_mux4_1 _09205_ (.S0(_03067_),
    .A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .S1(_03226_),
    .X(_04025_));
 sg13g2_mux4_1 _09206_ (.S0(_03067_),
    .A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .S1(_03226_),
    .X(_04026_));
 sg13g2_mux2_1 _09207_ (.A0(_04025_),
    .A1(_04026_),
    .S(net65),
    .X(_04027_));
 sg13g2_buf_1 _09208_ (.A(_04027_),
    .X(_04028_));
 sg13g2_nand3b_1 _09209_ (.B(net133),
    .C(_04028_),
    .Y(_04029_),
    .A_N(net55));
 sg13g2_nor2_1 _09210_ (.A(_04007_),
    .B(_04029_),
    .Y(_04030_));
 sg13g2_nand3_1 _09211_ (.B(_03223_),
    .C(_03224_),
    .A(_03185_),
    .Y(_04031_));
 sg13g2_nand3_1 _09212_ (.B(_03227_),
    .C(_03228_),
    .A(_03113_),
    .Y(_04032_));
 sg13g2_a21o_1 _09213_ (.A2(_03234_),
    .A1(_03183_),
    .B1(_03235_),
    .X(_04033_));
 sg13g2_a221oi_1 _09214_ (.B2(_03120_),
    .C1(_04033_),
    .B1(_03233_),
    .A1(_04031_),
    .Y(_04034_),
    .A2(_04032_));
 sg13g2_a21o_1 _09215_ (.A2(_03121_),
    .A1(_03116_),
    .B1(net65),
    .X(_04035_));
 sg13g2_buf_1 _09216_ (.A(_04035_),
    .X(_04036_));
 sg13g2_a21o_1 _09217_ (.A2(_03154_),
    .A1(_03126_),
    .B1(_03172_),
    .X(_04037_));
 sg13g2_buf_1 _09218_ (.A(_04037_),
    .X(_04038_));
 sg13g2_a21oi_1 _09219_ (.A1(_04036_),
    .A2(_04038_),
    .Y(_04039_),
    .B1(_04028_));
 sg13g2_nand2_1 _09220_ (.Y(_04040_),
    .A(_04015_),
    .B(_04021_));
 sg13g2_buf_1 _09221_ (.A(_04040_),
    .X(_04041_));
 sg13g2_nand2_1 _09222_ (.Y(_04042_),
    .A(net55),
    .B(net141));
 sg13g2_nor4_2 _09223_ (.A(_04005_),
    .B(_04034_),
    .C(_04039_),
    .Y(_04043_),
    .D(_04042_));
 sg13g2_mux2_1 _09224_ (.A0(_04030_),
    .A1(_04043_),
    .S(_03294_),
    .X(_04044_));
 sg13g2_xnor2_1 _09225_ (.Y(_04045_),
    .A(_03326_),
    .B(_04044_));
 sg13g2_mux2_1 _09226_ (.A0(_03366_),
    .A1(_03363_),
    .S(net65),
    .X(_04046_));
 sg13g2_buf_1 _09227_ (.A(_04046_),
    .X(_04047_));
 sg13g2_a21oi_1 _09228_ (.A1(_03341_),
    .A2(_03345_),
    .Y(_04048_),
    .B1(_04047_));
 sg13g2_a221oi_1 _09229_ (.B2(_03325_),
    .C1(_03115_),
    .B1(_03321_),
    .A1(_03288_),
    .Y(_04049_),
    .A2(_03292_));
 sg13g2_and4_1 _09230_ (.A(net52),
    .B(net42),
    .C(_04048_),
    .D(_04049_),
    .X(_04050_));
 sg13g2_buf_1 _09231_ (.A(_04050_),
    .X(_04051_));
 sg13g2_nor4_1 _09232_ (.A(net52),
    .B(net42),
    .C(_04007_),
    .D(_04029_),
    .Y(_04052_));
 sg13g2_inv_1 _09233_ (.Y(_04053_),
    .A(_03115_));
 sg13g2_nand4_1 _09234_ (.B(_03292_),
    .C(_03321_),
    .A(_03288_),
    .Y(_04054_),
    .D(_03325_));
 sg13g2_buf_2 _09235_ (.A(_04054_),
    .X(_04055_));
 sg13g2_nand3_1 _09236_ (.B(_03345_),
    .C(_04047_),
    .A(_03341_),
    .Y(_04056_));
 sg13g2_buf_2 _09237_ (.A(_04056_),
    .X(_04057_));
 sg13g2_nor3_1 _09238_ (.A(_04053_),
    .B(_04055_),
    .C(_04057_),
    .Y(_04058_));
 sg13g2_a22oi_1 _09239_ (.Y(_04059_),
    .B1(_04052_),
    .B2(_04058_),
    .A2(_04051_),
    .A1(_04043_));
 sg13g2_xnor2_1 _09240_ (.Y(_04060_),
    .A(_03280_),
    .B(_04059_));
 sg13g2_nor2b_1 _09241_ (.A(_04045_),
    .B_N(_04060_),
    .Y(_04061_));
 sg13g2_and4_1 _09242_ (.A(_03280_),
    .B(_03303_),
    .C(net41),
    .D(_03352_),
    .X(_04062_));
 sg13g2_nand3_1 _09243_ (.B(_04051_),
    .C(_04062_),
    .A(_04043_),
    .Y(_04063_));
 sg13g2_or3_1 _09244_ (.A(_04053_),
    .B(_04055_),
    .C(_04057_),
    .X(_04064_));
 sg13g2_nand3_1 _09245_ (.B(_03278_),
    .C(net133),
    .A(_03274_),
    .Y(_04065_));
 sg13g2_or4_1 _09246_ (.A(_03198_),
    .B(net42),
    .C(_03303_),
    .D(_04065_),
    .X(_04066_));
 sg13g2_buf_1 _09247_ (.A(_04066_),
    .X(_04067_));
 sg13g2_or3_1 _09248_ (.A(_03352_),
    .B(_04007_),
    .C(_04029_),
    .X(_04068_));
 sg13g2_or4_1 _09249_ (.A(net41),
    .B(_04064_),
    .C(_04067_),
    .D(_04068_),
    .X(_04069_));
 sg13g2_nand3_1 _09250_ (.B(_04063_),
    .C(_04069_),
    .A(_03375_),
    .Y(_04070_));
 sg13g2_a21o_1 _09251_ (.A2(_04069_),
    .A1(_04063_),
    .B1(_03375_),
    .X(_04071_));
 sg13g2_inv_1 _09252_ (.Y(_04072_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ));
 sg13g2_inv_1 _09253_ (.Y(_04073_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ));
 sg13g2_inv_1 _09254_ (.Y(_04074_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ));
 sg13g2_inv_1 _09255_ (.Y(_04075_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ));
 sg13g2_mux4_1 _09256_ (.S0(_03066_),
    .A0(_04072_),
    .A1(_04073_),
    .A2(_04074_),
    .A3(_04075_),
    .S1(_03153_),
    .X(_04076_));
 sg13g2_inv_1 _09257_ (.Y(_04077_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ));
 sg13g2_inv_1 _09258_ (.Y(_04078_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ));
 sg13g2_inv_1 _09259_ (.Y(_04079_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ));
 sg13g2_inv_1 _09260_ (.Y(_04080_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ));
 sg13g2_mux4_1 _09261_ (.S0(_03066_),
    .A0(_04077_),
    .A1(_04078_),
    .A2(_04079_),
    .A3(_04080_),
    .S1(net82),
    .X(_04081_));
 sg13g2_mux2_1 _09262_ (.A0(_04076_),
    .A1(_04081_),
    .S(_03124_),
    .X(_04082_));
 sg13g2_buf_2 _09263_ (.A(_04082_),
    .X(_04083_));
 sg13g2_nand2_1 _09264_ (.Y(_04084_),
    .A(net141),
    .B(_04083_));
 sg13g2_nand2_1 _09265_ (.Y(_04085_),
    .A(_04005_),
    .B(_04028_));
 sg13g2_a21o_1 _09266_ (.A2(_04085_),
    .A1(_04084_),
    .B1(_03175_),
    .X(_04086_));
 sg13g2_o21ai_1 _09267_ (.B1(net141),
    .Y(_04087_),
    .A1(_04005_),
    .A2(_04034_));
 sg13g2_a22oi_1 _09268_ (.Y(_04088_),
    .B1(_03321_),
    .B2(_03325_),
    .A2(_03292_),
    .A1(_03288_));
 sg13g2_buf_1 _09269_ (.A(_04088_),
    .X(_04089_));
 sg13g2_nor2_1 _09270_ (.A(_03115_),
    .B(net133),
    .Y(_04090_));
 sg13g2_and3_1 _09271_ (.X(_04091_),
    .A(_04089_),
    .B(_04048_),
    .C(_04090_));
 sg13g2_buf_8 _09272_ (.A(_04091_),
    .X(_04092_));
 sg13g2_nand4_1 _09273_ (.B(_04086_),
    .C(_04087_),
    .A(_03270_),
    .Y(_04093_),
    .D(_04092_));
 sg13g2_a21o_1 _09274_ (.A2(_03257_),
    .A1(_03183_),
    .B1(_03267_),
    .X(_04094_));
 sg13g2_a21o_1 _09275_ (.A2(_03263_),
    .A1(_03258_),
    .B1(_04094_),
    .X(_04095_));
 sg13g2_nand3_1 _09276_ (.B(net133),
    .C(_04028_),
    .A(_03115_),
    .Y(_04096_));
 sg13g2_nor4_1 _09277_ (.A(_04007_),
    .B(_04055_),
    .C(_04057_),
    .D(_04096_),
    .Y(_04097_));
 sg13g2_a21oi_1 _09278_ (.A1(_04095_),
    .A2(_04097_),
    .Y(_04098_),
    .B1(_03200_));
 sg13g2_nand3_1 _09279_ (.B(_04048_),
    .C(_04090_),
    .A(_04089_),
    .Y(_04099_));
 sg13g2_nor3_1 _09280_ (.A(net52),
    .B(_04095_),
    .C(_04099_),
    .Y(_04100_));
 sg13g2_and2_1 _09281_ (.A(_04086_),
    .B(_04087_),
    .X(_04101_));
 sg13g2_buf_1 _09282_ (.A(_04101_),
    .X(_04102_));
 sg13g2_or4_1 _09283_ (.A(_04007_),
    .B(_04055_),
    .C(_04057_),
    .D(_04096_),
    .X(_04103_));
 sg13g2_nor3_1 _09284_ (.A(net52),
    .B(net55),
    .C(_04103_),
    .Y(_04104_));
 sg13g2_a221oi_1 _09285_ (.B2(_04102_),
    .C1(_04104_),
    .B1(_04100_),
    .A1(_04093_),
    .Y(_04105_),
    .A2(_04098_));
 sg13g2_a21oi_1 _09286_ (.A1(_04070_),
    .A2(_04071_),
    .Y(_04106_),
    .B1(_04105_));
 sg13g2_nor3_1 _09287_ (.A(net41),
    .B(_04064_),
    .C(_04067_),
    .Y(_04107_));
 sg13g2_nand2_1 _09288_ (.Y(_04108_),
    .A(net52),
    .B(net42));
 sg13g2_nand3_1 _09289_ (.B(_03303_),
    .C(net41),
    .A(_03280_),
    .Y(_04109_));
 sg13g2_nor3_1 _09290_ (.A(_04108_),
    .B(_04109_),
    .C(_04099_),
    .Y(_04110_));
 sg13g2_or3_1 _09291_ (.A(_03212_),
    .B(_03269_),
    .C(_04083_),
    .X(_04111_));
 sg13g2_a21o_1 _09292_ (.A2(_04111_),
    .A1(_04084_),
    .B1(_03175_),
    .X(_04112_));
 sg13g2_buf_2 _09293_ (.A(_04112_),
    .X(_04113_));
 sg13g2_a221oi_1 _09294_ (.B2(_04005_),
    .C1(_04094_),
    .B1(_04083_),
    .A1(_03258_),
    .Y(_04114_),
    .A2(_03263_));
 sg13g2_a21o_1 _09295_ (.A2(_04114_),
    .A1(_03238_),
    .B1(net133),
    .X(_04115_));
 sg13g2_buf_8 _09296_ (.A(_04115_),
    .X(_04116_));
 sg13g2_and2_1 _09297_ (.A(_04113_),
    .B(_04116_),
    .X(_04117_));
 sg13g2_buf_1 _09298_ (.A(_04117_),
    .X(_04118_));
 sg13g2_mux2_1 _09299_ (.A0(_04107_),
    .A1(_04110_),
    .S(_04118_),
    .X(_04119_));
 sg13g2_xor2_1 _09300_ (.B(_04119_),
    .A(_03352_),
    .X(_04120_));
 sg13g2_and2_1 _09301_ (.A(_04089_),
    .B(_04048_),
    .X(_04121_));
 sg13g2_nand4_1 _09302_ (.B(_04113_),
    .C(_04121_),
    .A(net141),
    .Y(_04122_),
    .D(_04116_));
 sg13g2_a21oi_2 _09303_ (.B1(_03175_),
    .Y(_04123_),
    .A2(_04111_),
    .A1(_04084_));
 sg13g2_nor3_1 _09304_ (.A(net141),
    .B(_04055_),
    .C(_04057_),
    .Y(_04124_));
 sg13g2_a21oi_1 _09305_ (.A1(_04123_),
    .A2(_04124_),
    .Y(_04125_),
    .B1(_04053_));
 sg13g2_and3_1 _09306_ (.X(_04126_),
    .A(_04053_),
    .B(_04123_),
    .C(_04124_));
 sg13g2_a221oi_1 _09307_ (.B2(_04125_),
    .C1(_04126_),
    .B1(_04122_),
    .A1(_04092_),
    .Y(_04127_),
    .A2(_04118_));
 sg13g2_and4_1 _09308_ (.A(_04061_),
    .B(_04106_),
    .C(_04120_),
    .D(_04127_),
    .X(_04128_));
 sg13g2_nand4_1 _09309_ (.B(_03346_),
    .C(_03368_),
    .A(_03326_),
    .Y(_04129_),
    .D(_04090_));
 sg13g2_nand2_1 _09310_ (.Y(_04130_),
    .A(_04129_),
    .B(_04103_));
 sg13g2_a21oi_1 _09311_ (.A1(net55),
    .A2(_04129_),
    .Y(_04131_),
    .B1(_04067_));
 sg13g2_nand2_1 _09312_ (.Y(_04132_),
    .A(_03280_),
    .B(_03303_));
 sg13g2_nand2_1 _09313_ (.Y(_04133_),
    .A(net55),
    .B(_03294_));
 sg13g2_nor4_1 _09314_ (.A(_04108_),
    .B(_04132_),
    .C(_04129_),
    .D(_04133_),
    .Y(_04134_));
 sg13g2_a22oi_1 _09315_ (.Y(_04135_),
    .B1(_04134_),
    .B2(_04102_),
    .A2(_04131_),
    .A1(_04130_));
 sg13g2_xor2_1 _09316_ (.B(_04135_),
    .A(net41),
    .X(_04136_));
 sg13g2_nand2_1 _09317_ (.Y(_04137_),
    .A(_04113_),
    .B(_04116_));
 sg13g2_nand3_1 _09318_ (.B(net141),
    .C(_04051_),
    .A(_03280_),
    .Y(_04138_));
 sg13g2_nor2_1 _09319_ (.A(_04055_),
    .B(_04057_),
    .Y(_04139_));
 sg13g2_nor4_1 _09320_ (.A(_04053_),
    .B(net52),
    .C(net42),
    .D(_04065_),
    .Y(_04140_));
 sg13g2_nand3_1 _09321_ (.B(_04139_),
    .C(_04140_),
    .A(_04123_),
    .Y(_04141_));
 sg13g2_o21ai_1 _09322_ (.B1(_04141_),
    .Y(_04142_),
    .A1(_04137_),
    .A2(_04138_));
 sg13g2_xnor2_1 _09323_ (.Y(_04143_),
    .A(_03303_),
    .B(_04142_));
 sg13g2_and2_1 _09324_ (.A(_03341_),
    .B(_03345_),
    .X(_04144_));
 sg13g2_nor2_1 _09325_ (.A(_03294_),
    .B(_03326_),
    .Y(_04145_));
 sg13g2_and4_1 _09326_ (.A(_03238_),
    .B(_04041_),
    .C(_04089_),
    .D(_04114_),
    .X(_04146_));
 sg13g2_a22oi_1 _09327_ (.Y(_04147_),
    .B1(_04146_),
    .B2(_04113_),
    .A2(_04145_),
    .A1(_04030_));
 sg13g2_xnor2_1 _09328_ (.Y(_04148_),
    .A(_04144_),
    .B(_04147_));
 sg13g2_nand4_1 _09329_ (.B(_04113_),
    .C(_04092_),
    .A(_03199_),
    .Y(_04149_),
    .D(_04116_));
 sg13g2_nand2_1 _09330_ (.Y(_04150_),
    .A(_03115_),
    .B(net133));
 sg13g2_nor4_1 _09331_ (.A(_03199_),
    .B(_04055_),
    .C(_04057_),
    .D(_04150_),
    .Y(_04151_));
 sg13g2_inv_1 _09332_ (.Y(_04152_),
    .A(net42));
 sg13g2_a21oi_1 _09333_ (.A1(_04123_),
    .A2(_04151_),
    .Y(_04153_),
    .B1(_04152_));
 sg13g2_nor3_1 _09334_ (.A(_03200_),
    .B(_03248_),
    .C(_04099_),
    .Y(_04154_));
 sg13g2_and3_1 _09335_ (.X(_04155_),
    .A(_04152_),
    .B(_04123_),
    .C(_04151_));
 sg13g2_a221oi_1 _09336_ (.B2(_04118_),
    .C1(_04155_),
    .B1(_04154_),
    .A1(_04149_),
    .Y(_04156_),
    .A2(_04153_));
 sg13g2_buf_1 _09337_ (.A(net133),
    .X(_04157_));
 sg13g2_o21ai_1 _09338_ (.B1(_04157_),
    .Y(_04158_),
    .A1(_03212_),
    .A2(_03238_));
 sg13g2_nor2_1 _09339_ (.A(_03175_),
    .B(_04083_),
    .Y(_04159_));
 sg13g2_nand2b_1 _09340_ (.Y(_04160_),
    .B(net133),
    .A_N(_03270_));
 sg13g2_nand2_1 _09341_ (.Y(_04161_),
    .A(_04036_),
    .B(_04038_));
 sg13g2_a21oi_1 _09342_ (.A1(_04160_),
    .A2(_04042_),
    .Y(_04162_),
    .B1(_04161_));
 sg13g2_a21oi_1 _09343_ (.A1(net55),
    .A2(_04159_),
    .Y(_04163_),
    .B1(_04162_));
 sg13g2_nand2_1 _09344_ (.Y(_04164_),
    .A(_04095_),
    .B(_04039_));
 sg13g2_nand4_1 _09345_ (.B(_04158_),
    .C(_04163_),
    .A(_04087_),
    .Y(_04165_),
    .D(_04164_));
 sg13g2_nor2_1 _09346_ (.A(_03346_),
    .B(_04055_),
    .Y(_04166_));
 sg13g2_nor4_1 _09347_ (.A(_04005_),
    .B(_04034_),
    .C(_04144_),
    .D(_04042_),
    .Y(_04167_));
 sg13g2_nor2b_1 _09348_ (.A(_04039_),
    .B_N(_04089_),
    .Y(_04168_));
 sg13g2_a22oi_1 _09349_ (.Y(_04169_),
    .B1(_04167_),
    .B2(_04168_),
    .A2(_04166_),
    .A1(_04030_));
 sg13g2_xnor2_1 _09350_ (.Y(_04170_),
    .A(_04047_),
    .B(_04169_));
 sg13g2_xnor2_1 _09351_ (.Y(_04171_),
    .A(_03294_),
    .B(_04157_));
 sg13g2_a21oi_1 _09352_ (.A1(_04113_),
    .A2(_04116_),
    .Y(_04172_),
    .B1(_04171_));
 sg13g2_and3_1 _09353_ (.X(_04173_),
    .A(_04113_),
    .B(_04116_),
    .C(_04171_));
 sg13g2_nor3_1 _09354_ (.A(net270),
    .B(net233),
    .C(net182),
    .Y(_04174_));
 sg13g2_o21ai_1 _09355_ (.B1(_01377_),
    .Y(_04175_),
    .A1(_01121_),
    .A2(_04174_));
 sg13g2_a21oi_1 _09356_ (.A1(_03054_),
    .A2(_04175_),
    .Y(_04176_),
    .B1(_00874_));
 sg13g2_or2_1 _09357_ (.X(_04177_),
    .B(_04176_),
    .A(_03026_));
 sg13g2_buf_1 _09358_ (.A(_04177_),
    .X(_04178_));
 sg13g2_buf_1 _09359_ (.A(_03046_),
    .X(_04179_));
 sg13g2_buf_1 _09360_ (.A(net325),
    .X(_04180_));
 sg13g2_o21ai_1 _09361_ (.B1(_00032_),
    .Y(_04181_),
    .A1(net215),
    .A2(_04180_));
 sg13g2_nand4_1 _09362_ (.B(_03023_),
    .C(_04178_),
    .A(_03086_),
    .Y(_04182_),
    .D(_04181_));
 sg13g2_a221oi_1 _09363_ (.B2(_04038_),
    .C1(_04182_),
    .B1(_04036_),
    .A1(\z80.tv80s.i_tv80_core.IncDecZ ),
    .Y(_04183_),
    .A2(net263));
 sg13g2_o21ai_1 _09364_ (.B1(_04183_),
    .Y(_04184_),
    .A1(_04172_),
    .A2(_04173_));
 sg13g2_or4_1 _09365_ (.A(_04156_),
    .B(_04165_),
    .C(_04170_),
    .D(_04184_),
    .X(_04185_));
 sg13g2_nor4_1 _09366_ (.A(_04136_),
    .B(_04143_),
    .C(_04148_),
    .D(_04185_),
    .Y(_04186_));
 sg13g2_nand2_1 _09367_ (.Y(_04187_),
    .A(net343),
    .B(_03731_));
 sg13g2_a21oi_1 _09368_ (.A1(_04187_),
    .A2(_04182_),
    .Y(_04188_),
    .B1(net225));
 sg13g2_or3_1 _09369_ (.A(_01246_),
    .B(_03939_),
    .C(_04187_),
    .X(_04189_));
 sg13g2_o21ai_1 _09370_ (.B1(_04189_),
    .Y(_04190_),
    .A1(\z80.tv80s.i_tv80_core.IncDecZ ),
    .A2(_04188_));
 sg13g2_a21oi_1 _09371_ (.A1(_04128_),
    .A2(_04186_),
    .Y(_00379_),
    .B1(_04190_));
 sg13g2_or4_1 _09372_ (.A(_03738_),
    .B(_01581_),
    .C(_01584_),
    .D(_01586_),
    .X(_04191_));
 sg13g2_or3_1 _09373_ (.A(_01426_),
    .B(_01427_),
    .C(_04191_),
    .X(_04192_));
 sg13g2_buf_1 _09374_ (.A(_04192_),
    .X(_04193_));
 sg13g2_nand3_1 _09375_ (.B(\z80.tv80s.i_tv80_core.INT_s ),
    .C(_04193_),
    .A(\z80.tv80s.i_tv80_core.IntE ),
    .Y(_04194_));
 sg13g2_a21oi_1 _09376_ (.A1(_01071_),
    .A2(net239),
    .Y(_04195_),
    .B1(_01063_));
 sg13g2_nor3_2 _09377_ (.A(_01260_),
    .B(net234),
    .C(_04195_),
    .Y(_04196_));
 sg13g2_nor3_1 _09378_ (.A(\z80.tv80s.i_tv80_core.NMI_s ),
    .B(_04194_),
    .C(_04196_),
    .Y(_04197_));
 sg13g2_nand3_1 _09379_ (.B(\z80.tv80s.i_tv80_core.IncDecZ ),
    .C(_03731_),
    .A(_01296_),
    .Y(_04198_));
 sg13g2_nand3b_1 _09380_ (.B(_02353_),
    .C(_04198_),
    .Y(_04199_),
    .A_N(\z80.tv80s.i_tv80_core.No_BTR ));
 sg13g2_buf_1 _09381_ (.A(_04199_),
    .X(_04200_));
 sg13g2_nand2_1 _09382_ (.Y(_04201_),
    .A(net302),
    .B(_04200_));
 sg13g2_nor2_1 _09383_ (.A(net72),
    .B(_04201_),
    .Y(_04202_));
 sg13g2_nand2_1 _09384_ (.Y(_04203_),
    .A(_01002_),
    .B(_04202_));
 sg13g2_mux2_1 _09385_ (.A0(_04197_),
    .A1(_00825_),
    .S(_04203_),
    .X(_00380_));
 sg13g2_nor2b_1 _09386_ (.A(\z80.tv80s.i_tv80_core.IntE_FF2 ),
    .B_N(net398),
    .Y(_04204_));
 sg13g2_nor3_1 _09387_ (.A(\z80.tv80s.i_tv80_core.BusReq_s ),
    .B(net72),
    .C(_04201_),
    .Y(_04205_));
 sg13g2_and2_1 _09388_ (.A(_03975_),
    .B(_04205_),
    .X(_04206_));
 sg13g2_buf_1 _09389_ (.A(_04206_),
    .X(_04207_));
 sg13g2_inv_1 _09390_ (.Y(_04208_),
    .A(\z80.tv80s.i_tv80_core.NMI_s ));
 sg13g2_a21oi_1 _09391_ (.A1(_04208_),
    .A2(_04194_),
    .Y(_04209_),
    .B1(_04196_));
 sg13g2_or3_1 _09392_ (.A(_04180_),
    .B(_01425_),
    .C(_01426_),
    .X(_04210_));
 sg13g2_o21ai_1 _09393_ (.B1(net399),
    .Y(_04211_),
    .A1(_04191_),
    .A2(_04210_));
 sg13g2_a221oi_1 _09394_ (.B2(_04209_),
    .C1(_04211_),
    .B1(_04207_),
    .A1(_02249_),
    .Y(_04212_),
    .A2(_04204_));
 sg13g2_inv_1 _09395_ (.Y(_04213_),
    .A(_04212_));
 sg13g2_o21ai_1 _09396_ (.B1(_02250_),
    .Y(_04214_),
    .A1(net394),
    .A2(_04193_));
 sg13g2_nand3_1 _09397_ (.B(_04212_),
    .C(_04214_),
    .A(net398),
    .Y(_04215_));
 sg13g2_inv_1 _09398_ (.Y(_04216_),
    .A(\z80.tv80s.i_tv80_core.IntE ));
 sg13g2_a22oi_1 _09399_ (.Y(_00381_),
    .B1(_04215_),
    .B2(_04216_),
    .A2(_04213_),
    .A1(net328));
 sg13g2_inv_1 _09400_ (.Y(_04217_),
    .A(_04193_));
 sg13g2_nand2_1 _09401_ (.Y(_04218_),
    .A(_00637_),
    .B(_04217_));
 sg13g2_a221oi_1 _09402_ (.B2(_00136_),
    .C1(_04211_),
    .B1(_04218_),
    .A1(_04197_),
    .Y(_04219_),
    .A2(_04207_));
 sg13g2_nand2b_1 _09403_ (.Y(_04220_),
    .B(\z80.tv80s.i_tv80_core.IntE_FF2 ),
    .A_N(_00636_));
 sg13g2_nand2b_1 _09404_ (.Y(_00382_),
    .B(_04220_),
    .A_N(_04219_));
 sg13g2_nor3_1 _09405_ (.A(_04208_),
    .B(_04196_),
    .C(_04203_),
    .Y(_04221_));
 sg13g2_a21o_1 _09406_ (.A2(_04203_),
    .A1(net394),
    .B1(_04221_),
    .X(_00383_));
 sg13g2_inv_1 _09407_ (.Y(_04222_),
    .A(_00016_));
 sg13g2_nand3b_1 _09408_ (.B(\z80.tv80s.i_tv80_core.Oldnmi_n ),
    .C(net399),
    .Y(_04223_),
    .A_N(net4));
 sg13g2_a22oi_1 _09409_ (.Y(_00384_),
    .B1(_04208_),
    .B2(_04223_),
    .A2(_04222_),
    .A1(_02889_));
 sg13g2_o21ai_1 _09410_ (.B1(net220),
    .Y(_04224_),
    .A1(net237),
    .A2(_00685_));
 sg13g2_a21oi_1 _09411_ (.A1(net397),
    .A2(net284),
    .Y(_04225_),
    .B1(_04224_));
 sg13g2_nor3_1 _09412_ (.A(net182),
    .B(_02248_),
    .C(_04225_),
    .Y(_04226_));
 sg13g2_mux2_1 _09413_ (.A0(\z80.tv80s.i_tv80_core.No_BTR ),
    .A1(_04226_),
    .S(_03694_),
    .X(_00385_));
 sg13g2_mux2_1 _09414_ (.A0(\z80.tv80s.i_tv80_core.Oldnmi_n ),
    .A1(net4),
    .S(net326),
    .X(_00386_));
 sg13g2_nor2b_1 _09415_ (.A(\z80.tv80s.i_tv80_core.Halt_FF ),
    .B_N(_03012_),
    .Y(_04227_));
 sg13g2_nand4_1 _09416_ (.B(_02367_),
    .C(_03976_),
    .A(_01315_),
    .Y(_04228_),
    .D(_04227_));
 sg13g2_nor2_1 _09417_ (.A(_02286_),
    .B(_04228_),
    .Y(_04229_));
 sg13g2_nor2_1 _09418_ (.A(_01346_),
    .B(_04229_),
    .Y(_04230_));
 sg13g2_buf_2 _09419_ (.A(_04230_),
    .X(_04231_));
 sg13g2_buf_1 _09420_ (.A(_04231_),
    .X(_04232_));
 sg13g2_nor2_1 _09421_ (.A(net174),
    .B(_02687_),
    .Y(_04233_));
 sg13g2_a22oi_1 _09422_ (.Y(_04234_),
    .B1(_04233_),
    .B2(_02315_),
    .A2(net126),
    .A1(net253));
 sg13g2_nand2_1 _09423_ (.Y(_04235_),
    .A(_02297_),
    .B(_02663_));
 sg13g2_o21ai_1 _09424_ (.B1(_04235_),
    .Y(_04236_),
    .A1(net98),
    .A2(_04234_));
 sg13g2_nand3_1 _09425_ (.B(_00955_),
    .C(_01068_),
    .A(_00786_),
    .Y(_04237_));
 sg13g2_and2_1 _09426_ (.A(_01054_),
    .B(_01554_),
    .X(_04238_));
 sg13g2_buf_1 _09427_ (.A(_04238_),
    .X(_04239_));
 sg13g2_or4_1 _09428_ (.A(_00680_),
    .B(_01298_),
    .C(_01363_),
    .D(_04239_),
    .X(_04240_));
 sg13g2_buf_1 _09429_ (.A(_04240_),
    .X(_04241_));
 sg13g2_inv_1 _09430_ (.Y(_04242_),
    .A(_04241_));
 sg13g2_a21oi_1 _09431_ (.A1(_03448_),
    .A2(_04242_),
    .Y(_04243_),
    .B1(net277));
 sg13g2_a221oi_1 _09432_ (.B2(_01296_),
    .C1(_04243_),
    .B1(_04237_),
    .A1(_00959_),
    .Y(_04244_),
    .A2(_01371_));
 sg13g2_a21o_1 _09433_ (.A2(_00734_),
    .A1(_00773_),
    .B1(_00883_),
    .X(_04245_));
 sg13g2_nand3_1 _09434_ (.B(_01444_),
    .C(_04245_),
    .A(_01081_),
    .Y(_04246_));
 sg13g2_nor3_1 _09435_ (.A(_01156_),
    .B(_02129_),
    .C(_02923_),
    .Y(_04247_));
 sg13g2_nand4_1 _09436_ (.B(_01434_),
    .C(_02172_),
    .A(_00720_),
    .Y(_04248_),
    .D(_04247_));
 sg13g2_nor4_1 _09437_ (.A(_02162_),
    .B(_04237_),
    .C(_04246_),
    .D(_04248_),
    .Y(_04249_));
 sg13g2_nor2_1 _09438_ (.A(_00878_),
    .B(net279),
    .Y(_04250_));
 sg13g2_or4_1 _09439_ (.A(_00826_),
    .B(_02276_),
    .C(_04241_),
    .D(_04250_),
    .X(_04251_));
 sg13g2_nor2_1 _09440_ (.A(_03449_),
    .B(_04251_),
    .Y(_04252_));
 sg13g2_nand4_1 _09441_ (.B(_02268_),
    .C(_04249_),
    .A(_01057_),
    .Y(_04253_),
    .D(_04252_));
 sg13g2_a21oi_1 _09442_ (.A1(_04244_),
    .A2(_04253_),
    .Y(_04254_),
    .B1(_00968_));
 sg13g2_nand2_1 _09443_ (.Y(_04255_),
    .A(net219),
    .B(_01273_));
 sg13g2_o21ai_1 _09444_ (.B1(_01014_),
    .Y(_04256_),
    .A1(_02138_),
    .A2(_01028_));
 sg13g2_nor4_2 _09445_ (.A(_02261_),
    .B(_02265_),
    .C(_02269_),
    .Y(_04257_),
    .D(_02270_));
 sg13g2_a21oi_1 _09446_ (.A1(net307),
    .A2(_00881_),
    .Y(_04258_),
    .B1(net271));
 sg13g2_nand3_1 _09447_ (.B(_00918_),
    .C(_04258_),
    .A(_00655_),
    .Y(_04259_));
 sg13g2_a21oi_1 _09448_ (.A1(_01079_),
    .A2(_00665_),
    .Y(_04260_),
    .B1(_03737_));
 sg13g2_nand4_1 _09449_ (.B(_00823_),
    .C(_04259_),
    .A(_00859_),
    .Y(_04261_),
    .D(_04260_));
 sg13g2_nand2_1 _09450_ (.Y(_04262_),
    .A(_01053_),
    .B(_02115_));
 sg13g2_nor4_2 _09451_ (.A(_02162_),
    .B(_02869_),
    .C(_04261_),
    .Y(_04263_),
    .D(_04262_));
 sg13g2_a21oi_1 _09452_ (.A1(_04257_),
    .A2(_04263_),
    .Y(_04264_),
    .B1(_02891_));
 sg13g2_nand4_1 _09453_ (.B(_04255_),
    .C(_04256_),
    .A(_00214_),
    .Y(_04265_),
    .D(_04264_));
 sg13g2_o21ai_1 _09454_ (.B1(_01312_),
    .Y(_04266_),
    .A1(_04254_),
    .A2(_04265_));
 sg13g2_nand2_1 _09455_ (.Y(_04267_),
    .A(_01594_),
    .B(_04266_));
 sg13g2_buf_1 _09456_ (.A(_04267_),
    .X(_04268_));
 sg13g2_nor2_1 _09457_ (.A(net104),
    .B(_04268_),
    .Y(_04269_));
 sg13g2_buf_1 _09458_ (.A(_04269_),
    .X(_04270_));
 sg13g2_nand2_1 _09459_ (.Y(_04271_),
    .A(_04257_),
    .B(_04263_));
 sg13g2_buf_2 _09460_ (.A(_04271_),
    .X(_04272_));
 sg13g2_mux2_1 _09461_ (.A0(_00137_),
    .A1(_02891_),
    .S(_04272_),
    .X(_04273_));
 sg13g2_nor2_1 _09462_ (.A(_02315_),
    .B(_04273_),
    .Y(_04274_));
 sg13g2_buf_1 _09463_ (.A(_04268_),
    .X(_04275_));
 sg13g2_a22oi_1 _09464_ (.Y(_04276_),
    .B1(_04274_),
    .B2(net89),
    .A2(net76),
    .A1(_04236_));
 sg13g2_inv_2 _09465_ (.Y(_04277_),
    .A(_04231_));
 sg13g2_o21ai_1 _09466_ (.B1(_04277_),
    .Y(_04278_),
    .A1(_02088_),
    .A2(_04268_));
 sg13g2_buf_1 _09467_ (.A(_04278_),
    .X(_04279_));
 sg13g2_and2_1 _09468_ (.A(_04268_),
    .B(_04273_),
    .X(_04280_));
 sg13g2_o21ai_1 _09469_ (.B1(_02315_),
    .Y(_04281_),
    .A1(_04279_),
    .A2(_04280_));
 sg13g2_o21ai_1 _09470_ (.B1(_04281_),
    .Y(_00387_),
    .A1(net61),
    .A2(_04276_));
 sg13g2_inv_1 _09471_ (.Y(_04282_),
    .A(_02435_));
 sg13g2_buf_1 _09472_ (.A(_04279_),
    .X(_04283_));
 sg13g2_inv_1 _09473_ (.Y(_04284_),
    .A(_04268_));
 sg13g2_inv_1 _09474_ (.Y(_04285_),
    .A(_02566_));
 sg13g2_or4_1 _09475_ (.A(_02162_),
    .B(_02869_),
    .C(_04261_),
    .D(_04262_),
    .X(_04286_));
 sg13g2_buf_1 _09476_ (.A(_04286_),
    .X(_04287_));
 sg13g2_o21ai_1 _09477_ (.B1(_00211_),
    .Y(_04288_),
    .A1(_02272_),
    .A2(_04287_));
 sg13g2_buf_1 _09478_ (.A(_04288_),
    .X(_04289_));
 sg13g2_o21ai_1 _09479_ (.B1(_04289_),
    .Y(_04290_),
    .A1(_04285_),
    .A2(_04272_));
 sg13g2_or2_1 _09480_ (.X(_04291_),
    .B(_04290_),
    .A(_00188_));
 sg13g2_buf_1 _09481_ (.A(_04291_),
    .X(_04292_));
 sg13g2_xnor2_1 _09482_ (.Y(_04293_),
    .A(_02748_),
    .B(_04290_));
 sg13g2_nand2_1 _09483_ (.Y(_04294_),
    .A(_04292_),
    .B(_04293_));
 sg13g2_xnor2_1 _09484_ (.Y(_04295_),
    .A(_02828_),
    .B(_02619_));
 sg13g2_nand2b_1 _09485_ (.Y(_04296_),
    .B(_04295_),
    .A_N(_00137_));
 sg13g2_nor3_1 _09486_ (.A(_02272_),
    .B(_04287_),
    .C(_04296_),
    .Y(_04297_));
 sg13g2_xor2_1 _09487_ (.B(_00211_),
    .A(_02619_),
    .X(_04298_));
 sg13g2_or2_1 _09488_ (.X(_04299_),
    .B(_04298_),
    .A(_02891_));
 sg13g2_a21oi_1 _09489_ (.A1(_04257_),
    .A2(_04263_),
    .Y(_04300_),
    .B1(_04299_));
 sg13g2_o21ai_1 _09490_ (.B1(_02315_),
    .Y(_04301_),
    .A1(_04297_),
    .A2(_04300_));
 sg13g2_nand3_1 _09491_ (.B(_04257_),
    .C(_04263_),
    .A(_02828_),
    .Y(_04302_));
 sg13g2_nand3b_1 _09492_ (.B(_04289_),
    .C(_04302_),
    .Y(_04303_),
    .A_N(_00170_));
 sg13g2_inv_1 _09493_ (.Y(_04304_),
    .A(_00211_));
 sg13g2_a21oi_1 _09494_ (.A1(_04257_),
    .A2(_04263_),
    .Y(_04305_),
    .B1(_04304_));
 sg13g2_buf_1 _09495_ (.A(_04305_),
    .X(_04306_));
 sg13g2_inv_1 _09496_ (.Y(_04307_),
    .A(_00143_));
 sg13g2_nor3_1 _09497_ (.A(_04307_),
    .B(_02272_),
    .C(_04287_),
    .Y(_04308_));
 sg13g2_o21ai_1 _09498_ (.B1(_02640_),
    .Y(_04309_),
    .A1(_04306_),
    .A2(_04308_));
 sg13g2_or3_1 _09499_ (.A(_02640_),
    .B(_04306_),
    .C(_04308_),
    .X(_04310_));
 sg13g2_a22oi_1 _09500_ (.Y(_04311_),
    .B1(_04309_),
    .B2(_04310_),
    .A2(_04303_),
    .A1(_04301_));
 sg13g2_or2_1 _09501_ (.X(_04312_),
    .B(_04308_),
    .A(_04306_));
 sg13g2_nor2_1 _09502_ (.A(_00180_),
    .B(_04312_),
    .Y(_04313_));
 sg13g2_inv_1 _09503_ (.Y(_04314_),
    .A(_00146_));
 sg13g2_nor3_1 _09504_ (.A(_04314_),
    .B(_02272_),
    .C(_04287_),
    .Y(_04315_));
 sg13g2_o21ai_1 _09505_ (.B1(_03594_),
    .Y(_04316_),
    .A1(_04306_),
    .A2(_04315_));
 sg13g2_or3_1 _09506_ (.A(_03594_),
    .B(_04306_),
    .C(_04315_),
    .X(_04317_));
 sg13g2_a21oi_1 _09507_ (.A1(_04316_),
    .A2(_04317_),
    .Y(_04318_),
    .B1(_03627_));
 sg13g2_o21ai_1 _09508_ (.B1(_04318_),
    .Y(_04319_),
    .A1(_04311_),
    .A2(_04313_));
 sg13g2_or2_1 _09509_ (.X(_04320_),
    .B(_04315_),
    .A(_04306_));
 sg13g2_nor3_1 _09510_ (.A(_00182_),
    .B(_03627_),
    .C(_04320_),
    .Y(_04321_));
 sg13g2_nor2b_1 _09511_ (.A(_04321_),
    .B_N(_00184_),
    .Y(_04322_));
 sg13g2_inv_1 _09512_ (.Y(_04323_),
    .A(_00152_));
 sg13g2_o21ai_1 _09513_ (.B1(_04289_),
    .Y(_04324_),
    .A1(_04323_),
    .A2(_04272_));
 sg13g2_xnor2_1 _09514_ (.Y(_04325_),
    .A(_02724_),
    .B(_04324_));
 sg13g2_inv_1 _09515_ (.Y(_04326_),
    .A(_02502_));
 sg13g2_o21ai_1 _09516_ (.B1(_04289_),
    .Y(_04327_),
    .A1(_04326_),
    .A2(_04272_));
 sg13g2_inv_1 _09517_ (.Y(_04328_),
    .A(_04327_));
 sg13g2_nand2b_1 _09518_ (.Y(_04329_),
    .B(_04328_),
    .A_N(_04325_));
 sg13g2_a21o_1 _09519_ (.A2(_04322_),
    .A1(_04319_),
    .B1(_04329_),
    .X(_04330_));
 sg13g2_buf_1 _09520_ (.A(_04330_),
    .X(_04331_));
 sg13g2_nand2_1 _09521_ (.Y(_04332_),
    .A(_04316_),
    .B(_04317_));
 sg13g2_o21ai_1 _09522_ (.B1(_04332_),
    .Y(_04333_),
    .A1(_04311_),
    .A2(_04313_));
 sg13g2_or2_1 _09523_ (.X(_04334_),
    .B(_04320_),
    .A(_00182_));
 sg13g2_and2_1 _09524_ (.A(_03627_),
    .B(_04327_),
    .X(_04335_));
 sg13g2_nand2b_1 _09525_ (.Y(_04336_),
    .B(_04335_),
    .A_N(_04325_));
 sg13g2_a21o_1 _09526_ (.A2(_04334_),
    .A1(_04333_),
    .B1(_04336_),
    .X(_04337_));
 sg13g2_buf_1 _09527_ (.A(_04337_),
    .X(_04338_));
 sg13g2_or2_1 _09528_ (.X(_04339_),
    .B(_04324_),
    .A(_00186_));
 sg13g2_buf_1 _09529_ (.A(_04339_),
    .X(_04340_));
 sg13g2_and2_1 _09530_ (.A(_04292_),
    .B(_04340_),
    .X(_04341_));
 sg13g2_nand3_1 _09531_ (.B(_04338_),
    .C(_04341_),
    .A(_04331_),
    .Y(_04342_));
 sg13g2_and3_1 _09532_ (.X(_04343_),
    .A(_03686_),
    .B(_04294_),
    .C(_04342_));
 sg13g2_inv_1 _09533_ (.Y(_04344_),
    .A(_00158_));
 sg13g2_o21ai_1 _09534_ (.B1(_04289_),
    .Y(_04345_),
    .A1(_04344_),
    .A2(_04272_));
 sg13g2_buf_1 _09535_ (.A(_04345_),
    .X(_04346_));
 sg13g2_nor3_1 _09536_ (.A(net373),
    .B(net372),
    .C(_04346_),
    .Y(_04347_));
 sg13g2_nor2_1 _09537_ (.A(_04344_),
    .B(_04272_),
    .Y(_04348_));
 sg13g2_nor2_1 _09538_ (.A(_04306_),
    .B(_04348_),
    .Y(_04349_));
 sg13g2_buf_2 _09539_ (.A(_04349_),
    .X(_04350_));
 sg13g2_nor3_1 _09540_ (.A(_02803_),
    .B(_03686_),
    .C(_04350_),
    .Y(_04351_));
 sg13g2_and3_1 _09541_ (.X(_04352_),
    .A(_04294_),
    .B(_04342_),
    .C(_04351_));
 sg13g2_o21ai_1 _09542_ (.B1(_00139_),
    .Y(_04353_),
    .A1(net373),
    .A2(_02785_));
 sg13g2_nand2b_1 _09543_ (.Y(_04354_),
    .B(_04353_),
    .A_N(net372));
 sg13g2_a21oi_1 _09544_ (.A1(_00142_),
    .A2(_04354_),
    .Y(_04355_),
    .B1(_04346_));
 sg13g2_a221oi_1 _09545_ (.B2(net372),
    .C1(_04355_),
    .B1(_04352_),
    .A1(_04343_),
    .Y(_04356_),
    .A2(_04347_));
 sg13g2_buf_1 _09546_ (.A(_04346_),
    .X(_04357_));
 sg13g2_xnor2_1 _09547_ (.Y(_04358_),
    .A(_02435_),
    .B(net103));
 sg13g2_xnor2_1 _09548_ (.Y(_04359_),
    .A(_04356_),
    .B(_04358_));
 sg13g2_nor2_1 _09549_ (.A(_04282_),
    .B(net174),
    .Y(_04360_));
 sg13g2_a21oi_1 _09550_ (.A1(_01740_),
    .A2(net174),
    .Y(_04361_),
    .B1(_04360_));
 sg13g2_o21ai_1 _09551_ (.B1(_02445_),
    .Y(_04362_),
    .A1(net85),
    .A2(_04361_));
 sg13g2_a22oi_1 _09552_ (.Y(_04363_),
    .B1(_02406_),
    .B2(_04362_),
    .A2(net98),
    .A1(net389));
 sg13g2_nand2_1 _09553_ (.Y(_04364_),
    .A(net76),
    .B(_04363_));
 sg13g2_o21ai_1 _09554_ (.B1(_04364_),
    .Y(_04365_),
    .A1(net88),
    .A2(_04359_));
 sg13g2_a22oi_1 _09555_ (.Y(_00388_),
    .B1(_04365_),
    .B2(_04277_),
    .A2(net54),
    .A1(_04282_));
 sg13g2_nand2_1 _09556_ (.Y(_04366_),
    .A(_02833_),
    .B(_04282_));
 sg13g2_a21oi_1 _09557_ (.A1(_02410_),
    .A2(_04366_),
    .Y(_04367_),
    .B1(net103));
 sg13g2_nand4_1 _09558_ (.B(_04331_),
    .C(_04338_),
    .A(_02785_),
    .Y(_04368_),
    .D(_04341_));
 sg13g2_and3_1 _09559_ (.X(_04369_),
    .A(_02785_),
    .B(_04292_),
    .C(_04293_));
 sg13g2_a21oi_1 _09560_ (.A1(_02785_),
    .A2(_03685_),
    .Y(_04370_),
    .B1(_04369_));
 sg13g2_nand4_1 _09561_ (.B(_04350_),
    .C(_04368_),
    .A(_02803_),
    .Y(_04371_),
    .D(_04370_));
 sg13g2_nand3_1 _09562_ (.B(_03685_),
    .C(_04346_),
    .A(net373),
    .Y(_04372_));
 sg13g2_or2_1 _09563_ (.X(_04373_),
    .B(_04372_),
    .A(_04293_));
 sg13g2_a21oi_1 _09564_ (.A1(_04331_),
    .A2(_04338_),
    .Y(_04374_),
    .B1(_04373_));
 sg13g2_nor2_1 _09565_ (.A(_04292_),
    .B(_04372_),
    .Y(_04375_));
 sg13g2_nor3_1 _09566_ (.A(_04293_),
    .B(_04340_),
    .C(_04372_),
    .Y(_04376_));
 sg13g2_nor2_1 _09567_ (.A(_00139_),
    .B(_04346_),
    .Y(_04377_));
 sg13g2_nor4_1 _09568_ (.A(_04374_),
    .B(_04375_),
    .C(_04376_),
    .D(_04377_),
    .Y(_04378_));
 sg13g2_nand3_1 _09569_ (.B(_02435_),
    .C(_04346_),
    .A(net372),
    .Y(_04379_));
 sg13g2_or3_1 _09570_ (.A(net372),
    .B(_02435_),
    .C(_04346_),
    .X(_04380_));
 sg13g2_a22oi_1 _09571_ (.Y(_04381_),
    .B1(_04379_),
    .B2(_04380_),
    .A2(_04378_),
    .A1(_04371_));
 sg13g2_nor2_2 _09572_ (.A(_04367_),
    .B(_04381_),
    .Y(_04382_));
 sg13g2_xnor2_1 _09573_ (.Y(_04383_),
    .A(_02458_),
    .B(net103));
 sg13g2_xnor2_1 _09574_ (.Y(_04384_),
    .A(_04382_),
    .B(_04383_));
 sg13g2_a21oi_1 _09575_ (.A1(_02458_),
    .A2(net213),
    .Y(_04385_),
    .B1(_02457_));
 sg13g2_o21ai_1 _09576_ (.B1(_02478_),
    .Y(_04386_),
    .A1(_02375_),
    .A2(_04385_));
 sg13g2_a22oi_1 _09577_ (.Y(_04387_),
    .B1(_02455_),
    .B2(_04386_),
    .A2(_02393_),
    .A1(net388));
 sg13g2_nand2_1 _09578_ (.Y(_04388_),
    .A(net76),
    .B(_04387_));
 sg13g2_o21ai_1 _09579_ (.B1(_04388_),
    .Y(_04389_),
    .A1(net88),
    .A2(_04384_));
 sg13g2_a22oi_1 _09580_ (.Y(_00389_),
    .B1(_04389_),
    .B2(_04277_),
    .A2(net54),
    .A1(_02459_));
 sg13g2_inv_1 _09581_ (.Y(_04390_),
    .A(_04269_));
 sg13g2_a21oi_1 _09582_ (.A1(_02494_),
    .A2(net213),
    .Y(_04391_),
    .B1(_02493_));
 sg13g2_o21ai_1 _09583_ (.B1(_02514_),
    .Y(_04392_),
    .A1(net85),
    .A2(_04391_));
 sg13g2_a22oi_1 _09584_ (.Y(_04393_),
    .B1(_02491_),
    .B2(_04392_),
    .A2(net98),
    .A1(net387));
 sg13g2_nor3_1 _09585_ (.A(net61),
    .B(_04390_),
    .C(_04393_),
    .Y(_04394_));
 sg13g2_nor2_2 _09586_ (.A(_04231_),
    .B(net88),
    .Y(_04395_));
 sg13g2_nor2_1 _09587_ (.A(_02410_),
    .B(_02458_),
    .Y(_04396_));
 sg13g2_o21ai_1 _09588_ (.B1(_04350_),
    .Y(_04397_),
    .A1(_02460_),
    .A2(_04396_));
 sg13g2_nand3_1 _09589_ (.B(_02459_),
    .C(_04350_),
    .A(_04282_),
    .Y(_04398_));
 sg13g2_nand3_1 _09590_ (.B(_02458_),
    .C(net103),
    .A(_02435_),
    .Y(_04399_));
 sg13g2_a21o_1 _09591_ (.A2(_04399_),
    .A1(_04398_),
    .B1(_04356_),
    .X(_04400_));
 sg13g2_nand2_1 _09592_ (.Y(_04401_),
    .A(_04397_),
    .B(_04400_));
 sg13g2_xnor2_1 _09593_ (.Y(_04402_),
    .A(_02495_),
    .B(net103));
 sg13g2_xnor2_1 _09594_ (.Y(_04403_),
    .A(_04401_),
    .B(_04402_));
 sg13g2_a22oi_1 _09595_ (.Y(_04404_),
    .B1(_04395_),
    .B2(_04403_),
    .A2(net54),
    .A1(_02494_));
 sg13g2_nand2b_1 _09596_ (.Y(_00390_),
    .B(_04404_),
    .A_N(_04394_));
 sg13g2_nor2_1 _09597_ (.A(_02460_),
    .B(_02459_),
    .Y(_04405_));
 sg13g2_and2_1 _09598_ (.A(_02498_),
    .B(_04350_),
    .X(_04406_));
 sg13g2_buf_1 _09599_ (.A(_04406_),
    .X(_04407_));
 sg13g2_o21ai_1 _09600_ (.B1(_04407_),
    .Y(_04408_),
    .A1(_02494_),
    .A2(_04405_));
 sg13g2_nand3_1 _09601_ (.B(_02494_),
    .C(net103),
    .A(_02458_),
    .Y(_04409_));
 sg13g2_nand2_1 _09602_ (.Y(_04410_),
    .A(_00148_),
    .B(_04407_));
 sg13g2_mux2_1 _09603_ (.A0(_04409_),
    .A1(_04410_),
    .S(_04382_),
    .X(_04411_));
 sg13g2_nand2_1 _09604_ (.Y(_04412_),
    .A(_02528_),
    .B(_04395_));
 sg13g2_a21oi_1 _09605_ (.A1(_04408_),
    .A2(_04411_),
    .Y(_04413_),
    .B1(_04412_));
 sg13g2_nand4_1 _09606_ (.B(net89),
    .C(_04408_),
    .A(_02527_),
    .Y(_04414_),
    .D(_04411_));
 sg13g2_a21oi_1 _09607_ (.A1(_02527_),
    .A2(net213),
    .Y(_04415_),
    .B1(_02526_));
 sg13g2_o21ai_1 _09608_ (.B1(_02546_),
    .Y(_04416_),
    .A1(net85),
    .A2(_04415_));
 sg13g2_a22oi_1 _09609_ (.Y(_04417_),
    .B1(_02525_),
    .B2(_04416_),
    .A2(net109),
    .A1(net386));
 sg13g2_nor2_1 _09610_ (.A(_04390_),
    .B(_04417_),
    .Y(_04418_));
 sg13g2_a22oi_1 _09611_ (.Y(_04419_),
    .B1(_04418_),
    .B2(_04277_),
    .A2(_04279_),
    .A1(_02527_));
 sg13g2_nand3b_1 _09612_ (.B(_04414_),
    .C(_04419_),
    .Y(_00391_),
    .A_N(_04413_));
 sg13g2_a21oi_1 _09613_ (.A1(_02560_),
    .A2(net213),
    .Y(_04420_),
    .B1(_02559_));
 sg13g2_o21ai_1 _09614_ (.B1(_02577_),
    .Y(_04421_),
    .A1(net85),
    .A2(_04420_));
 sg13g2_a22oi_1 _09615_ (.Y(_04422_),
    .B1(_02558_),
    .B2(_04421_),
    .A2(net98),
    .A1(net385));
 sg13g2_nor3_1 _09616_ (.A(_04231_),
    .B(_04390_),
    .C(_04422_),
    .Y(_04423_));
 sg13g2_a21oi_1 _09617_ (.A1(_02560_),
    .A2(net54),
    .Y(_04424_),
    .B1(_04423_));
 sg13g2_nand2_1 _09618_ (.Y(_04425_),
    .A(_02560_),
    .B(_04268_));
 sg13g2_nand2_1 _09619_ (.Y(_04426_),
    .A(_02561_),
    .B(_04395_));
 sg13g2_nor4_1 _09620_ (.A(_02495_),
    .B(_02528_),
    .C(_04350_),
    .D(_04400_),
    .Y(_04427_));
 sg13g2_and2_1 _09621_ (.A(_02530_),
    .B(_04350_),
    .X(_04428_));
 sg13g2_nand4_1 _09622_ (.B(_04397_),
    .C(_04400_),
    .A(_02498_),
    .Y(_04429_),
    .D(_04428_));
 sg13g2_and2_1 _09623_ (.A(_02498_),
    .B(_02494_),
    .X(_04430_));
 sg13g2_o21ai_1 _09624_ (.B1(_04428_),
    .Y(_04431_),
    .A1(_02527_),
    .A2(_04430_));
 sg13g2_nand3b_1 _09625_ (.B(_04429_),
    .C(_04431_),
    .Y(_04432_),
    .A_N(_04427_));
 sg13g2_mux2_1 _09626_ (.A0(_04425_),
    .A1(_04426_),
    .S(_04432_),
    .X(_04433_));
 sg13g2_nand2_1 _09627_ (.Y(_00392_),
    .A(_04424_),
    .B(_04433_));
 sg13g2_nand4_1 _09628_ (.B(_02494_),
    .C(_02527_),
    .A(_02458_),
    .Y(_04434_),
    .D(_02560_));
 sg13g2_nand2b_1 _09629_ (.Y(_04435_),
    .B(net103),
    .A_N(_04434_));
 sg13g2_a21o_1 _09630_ (.A2(_02527_),
    .A1(_02530_),
    .B1(_02560_),
    .X(_04436_));
 sg13g2_nand3_1 _09631_ (.B(_04350_),
    .C(_04436_),
    .A(_00157_),
    .Y(_04437_));
 sg13g2_o21ai_1 _09632_ (.B1(_04437_),
    .Y(_04438_),
    .A1(_04382_),
    .A2(_04435_));
 sg13g2_o21ai_1 _09633_ (.B1(_02459_),
    .Y(_04439_),
    .A1(_04367_),
    .A2(_04381_));
 sg13g2_nand2_1 _09634_ (.Y(_04440_),
    .A(_02460_),
    .B(_02495_));
 sg13g2_and4_1 _09635_ (.A(_02530_),
    .B(_00157_),
    .C(_04407_),
    .D(_04440_),
    .X(_04441_));
 sg13g2_o21ai_1 _09636_ (.B1(_04441_),
    .Y(_04442_),
    .A1(_02494_),
    .A2(_04439_));
 sg13g2_nand2b_1 _09637_ (.Y(_04443_),
    .B(_04442_),
    .A_N(_04438_));
 sg13g2_nor3_1 _09638_ (.A(_02591_),
    .B(net61),
    .C(net88),
    .Y(_04444_));
 sg13g2_o21ai_1 _09639_ (.B1(_04277_),
    .Y(_04445_),
    .A1(net88),
    .A2(_04443_));
 sg13g2_nor2_1 _09640_ (.A(_02591_),
    .B(net192),
    .Y(_04446_));
 sg13g2_a21oi_1 _09641_ (.A1(_02080_),
    .A2(net193),
    .Y(_04447_),
    .B1(_04446_));
 sg13g2_o21ai_1 _09642_ (.B1(_02607_),
    .Y(_04448_),
    .A1(net85),
    .A2(_04447_));
 sg13g2_a221oi_1 _09643_ (.B2(_04448_),
    .C1(_04231_),
    .B1(_02589_),
    .A1(net349),
    .Y(_04449_),
    .A2(net109));
 sg13g2_nand2_1 _09644_ (.Y(_04450_),
    .A(\z80.tv80s.i_tv80_core.PC[15] ),
    .B(net104));
 sg13g2_o21ai_1 _09645_ (.B1(_04450_),
    .Y(_04451_),
    .A1(net104),
    .A2(_04449_));
 sg13g2_nor2_1 _09646_ (.A(net89),
    .B(_04451_),
    .Y(_04452_));
 sg13g2_a221oi_1 _09647_ (.B2(_02591_),
    .C1(_04452_),
    .B1(_04445_),
    .A1(_04443_),
    .Y(_00393_),
    .A2(_04444_));
 sg13g2_nor2_1 _09648_ (.A(_02426_),
    .B(net252),
    .Y(_04453_));
 sg13g2_a21oi_1 _09649_ (.A1(_02620_),
    .A2(net252),
    .Y(_04454_),
    .B1(_04453_));
 sg13g2_nor2_1 _09650_ (.A(_02378_),
    .B(_04454_),
    .Y(_04455_));
 sg13g2_a22oi_1 _09651_ (.Y(_04456_),
    .B1(_04455_),
    .B2(_02441_),
    .A2(_02618_),
    .A1(net126));
 sg13g2_nand2b_1 _09652_ (.Y(_04457_),
    .B(_02385_),
    .A_N(_02426_));
 sg13g2_o21ai_1 _09653_ (.B1(_04457_),
    .Y(_04458_),
    .A1(_02484_),
    .A2(_04456_));
 sg13g2_and2_1 _09654_ (.A(_04272_),
    .B(_04298_),
    .X(_04459_));
 sg13g2_nor2_1 _09655_ (.A(_04272_),
    .B(_04295_),
    .Y(_04460_));
 sg13g2_nor2_1 _09656_ (.A(_04459_),
    .B(_04460_),
    .Y(_04461_));
 sg13g2_nor2_1 _09657_ (.A(_02315_),
    .B(_04461_),
    .Y(_04462_));
 sg13g2_a221oi_1 _09658_ (.B2(_00137_),
    .C1(_04462_),
    .B1(_04460_),
    .A1(_02891_),
    .Y(_04463_),
    .A2(_04459_));
 sg13g2_nand2_1 _09659_ (.Y(_04464_),
    .A(_04301_),
    .B(_04463_));
 sg13g2_a22oi_1 _09660_ (.Y(_04465_),
    .B1(_04464_),
    .B2(net89),
    .A2(_04458_),
    .A1(net76));
 sg13g2_nor2_1 _09661_ (.A(_04232_),
    .B(_04465_),
    .Y(_04466_));
 sg13g2_a21oi_1 _09662_ (.A1(_02620_),
    .A2(net54),
    .Y(_00394_),
    .B1(_04466_));
 sg13g2_nand2_1 _09663_ (.Y(_04467_),
    .A(_02640_),
    .B(_02345_));
 sg13g2_o21ai_1 _09664_ (.B1(_04467_),
    .Y(_04468_),
    .A1(_02664_),
    .A2(_02345_));
 sg13g2_o21ai_1 _09665_ (.B1(_02659_),
    .Y(_04469_),
    .A1(_02687_),
    .A2(_04468_));
 sg13g2_a22oi_1 _09666_ (.Y(_04470_),
    .B1(_04469_),
    .B2(net99),
    .A2(_02385_),
    .A1(_02664_));
 sg13g2_nand2_1 _09667_ (.Y(_04471_),
    .A(_04301_),
    .B(_04303_));
 sg13g2_xnor2_1 _09668_ (.Y(_04472_),
    .A(_04471_),
    .B(_04312_));
 sg13g2_nor2b_1 _09669_ (.A(_02640_),
    .B_N(_04472_),
    .Y(_04473_));
 sg13g2_a22oi_1 _09670_ (.Y(_04474_),
    .B1(_04473_),
    .B2(_04275_),
    .A2(_04470_),
    .A1(_04270_));
 sg13g2_nor2_1 _09671_ (.A(net88),
    .B(_04472_),
    .Y(_04475_));
 sg13g2_o21ai_1 _09672_ (.B1(_02640_),
    .Y(_04476_),
    .A1(_04279_),
    .A2(_04475_));
 sg13g2_o21ai_1 _09673_ (.B1(_04476_),
    .Y(_00395_),
    .A1(net61),
    .A2(_04474_));
 sg13g2_a22oi_1 _09674_ (.Y(_04477_),
    .B1(_02671_),
    .B2(net126),
    .A2(_04233_),
    .A1(_03594_));
 sg13g2_nand2_1 _09675_ (.Y(_04478_),
    .A(_02422_),
    .B(_02663_));
 sg13g2_o21ai_1 _09676_ (.B1(_04478_),
    .Y(_04479_),
    .A1(net98),
    .A2(_04477_));
 sg13g2_nor2_1 _09677_ (.A(_04311_),
    .B(_04313_),
    .Y(_04480_));
 sg13g2_xnor2_1 _09678_ (.Y(_04481_),
    .A(_04480_),
    .B(_04332_));
 sg13g2_a22oi_1 _09679_ (.Y(_04482_),
    .B1(_04481_),
    .B2(net89),
    .A2(_04479_),
    .A1(net76));
 sg13g2_nand2_1 _09680_ (.Y(_04483_),
    .A(_03594_),
    .B(_04283_));
 sg13g2_o21ai_1 _09681_ (.B1(_04483_),
    .Y(_00396_),
    .A1(net61),
    .A2(_04482_));
 sg13g2_a21oi_1 _09682_ (.A1(_03627_),
    .A2(_04233_),
    .Y(_04484_),
    .B1(_02700_));
 sg13g2_nand2_1 _09683_ (.Y(_04485_),
    .A(_02421_),
    .B(_02663_));
 sg13g2_o21ai_1 _09684_ (.B1(_04485_),
    .Y(_04486_),
    .A1(net98),
    .A2(_04484_));
 sg13g2_nand2_1 _09685_ (.Y(_04487_),
    .A(_04333_),
    .B(_04334_));
 sg13g2_xor2_1 _09686_ (.B(_04327_),
    .A(_03627_),
    .X(_04488_));
 sg13g2_xnor2_1 _09687_ (.Y(_04489_),
    .A(_04487_),
    .B(_04488_));
 sg13g2_a22oi_1 _09688_ (.Y(_04490_),
    .B1(_04489_),
    .B2(net89),
    .A2(_04486_),
    .A1(net76));
 sg13g2_nand2_1 _09689_ (.Y(_04491_),
    .A(_03627_),
    .B(net54));
 sg13g2_o21ai_1 _09690_ (.B1(_04491_),
    .Y(_00397_),
    .A1(net61),
    .A2(_04490_));
 sg13g2_inv_1 _09691_ (.Y(_04492_),
    .A(_02419_));
 sg13g2_nand2_1 _09692_ (.Y(_04493_),
    .A(_04492_),
    .B(_02456_));
 sg13g2_nand2_1 _09693_ (.Y(_04494_),
    .A(_02724_),
    .B(net252));
 sg13g2_a21oi_1 _09694_ (.A1(_04493_),
    .A2(_04494_),
    .Y(_04495_),
    .B1(net127));
 sg13g2_a22oi_1 _09695_ (.Y(_04496_),
    .B1(_04495_),
    .B2(_02441_),
    .A2(_02723_),
    .A1(net126));
 sg13g2_nor2_1 _09696_ (.A(net109),
    .B(_04496_),
    .Y(_04497_));
 sg13g2_a21oi_1 _09697_ (.A1(_04492_),
    .A2(_02385_),
    .Y(_04498_),
    .B1(_04497_));
 sg13g2_nand2_1 _09698_ (.Y(_04499_),
    .A(_04319_),
    .B(_04322_));
 sg13g2_a22oi_1 _09699_ (.Y(_04500_),
    .B1(_04499_),
    .B2(_04328_),
    .A2(_04335_),
    .A1(_04487_));
 sg13g2_xor2_1 _09700_ (.B(_04500_),
    .A(_04325_),
    .X(_04501_));
 sg13g2_a22oi_1 _09701_ (.Y(_04502_),
    .B1(_04501_),
    .B2(_04275_),
    .A2(_04498_),
    .A1(net76));
 sg13g2_nand2_1 _09702_ (.Y(_04503_),
    .A(\z80.tv80s.i_tv80_core.PC[5] ),
    .B(net54));
 sg13g2_o21ai_1 _09703_ (.B1(_04503_),
    .Y(_00398_),
    .A1(net61),
    .A2(_04502_));
 sg13g2_inv_1 _09704_ (.Y(_04504_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sg13g2_nand2_1 _09705_ (.Y(_04505_),
    .A(_04504_),
    .B(_02456_));
 sg13g2_nand2_1 _09706_ (.Y(_04506_),
    .A(_02748_),
    .B(net252));
 sg13g2_a21oi_1 _09707_ (.A1(_04505_),
    .A2(_04506_),
    .Y(_04507_),
    .B1(_02477_));
 sg13g2_a22oi_1 _09708_ (.Y(_04508_),
    .B1(_04507_),
    .B2(net84),
    .A2(_02747_),
    .A1(net126));
 sg13g2_nor2_1 _09709_ (.A(_02484_),
    .B(_04508_),
    .Y(_04509_));
 sg13g2_a21oi_1 _09710_ (.A1(_04504_),
    .A2(_02385_),
    .Y(_04510_),
    .B1(_04509_));
 sg13g2_nand3_1 _09711_ (.B(_04338_),
    .C(_04340_),
    .A(_04331_),
    .Y(_04511_));
 sg13g2_xnor2_1 _09712_ (.Y(_04512_),
    .A(_04293_),
    .B(_04511_));
 sg13g2_a22oi_1 _09713_ (.Y(_04513_),
    .B1(_04512_),
    .B2(net89),
    .A2(_04510_),
    .A1(_04270_));
 sg13g2_nand2_1 _09714_ (.Y(_04514_),
    .A(\z80.tv80s.i_tv80_core.PC[6] ),
    .B(net54));
 sg13g2_o21ai_1 _09715_ (.B1(_04514_),
    .Y(_00399_),
    .A1(net61),
    .A2(_04513_));
 sg13g2_o21ai_1 _09716_ (.B1(_02789_),
    .Y(_04515_),
    .A1(_03686_),
    .A2(_02639_));
 sg13g2_a22oi_1 _09717_ (.Y(_04516_),
    .B1(_04515_),
    .B2(net99),
    .A2(_02663_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sg13g2_and2_1 _09718_ (.A(_04294_),
    .B(_04342_),
    .X(_04517_));
 sg13g2_buf_1 _09719_ (.A(_04517_),
    .X(_04518_));
 sg13g2_xnor2_1 _09720_ (.Y(_04519_),
    .A(_03685_),
    .B(_04357_));
 sg13g2_xnor2_1 _09721_ (.Y(_04520_),
    .A(_04518_),
    .B(_04519_));
 sg13g2_a22oi_1 _09722_ (.Y(_04521_),
    .B1(_04520_),
    .B2(net89),
    .A2(_04516_),
    .A1(net76));
 sg13g2_nor2_1 _09723_ (.A(_04232_),
    .B(_04521_),
    .Y(_04522_));
 sg13g2_a21oi_1 _09724_ (.A1(_03686_),
    .A2(_04283_),
    .Y(_00400_),
    .B1(_04522_));
 sg13g2_a21oi_1 _09725_ (.A1(net373),
    .A2(net213),
    .Y(_04523_),
    .B1(_02801_));
 sg13g2_o21ai_1 _09726_ (.B1(_02800_),
    .Y(_04524_),
    .A1(net85),
    .A2(_04523_));
 sg13g2_a221oi_1 _09727_ (.B2(_04524_),
    .C1(_04231_),
    .B1(_02799_),
    .A1(net350),
    .Y(_04525_),
    .A2(net109));
 sg13g2_nor2_1 _09728_ (.A(net104),
    .B(_04525_),
    .Y(_04526_));
 sg13g2_a21oi_1 _09729_ (.A1(net373),
    .A2(net104),
    .Y(_04527_),
    .B1(_04526_));
 sg13g2_nand2_1 _09730_ (.Y(_04528_),
    .A(_03686_),
    .B(_04518_));
 sg13g2_mux2_1 _09731_ (.A0(_02785_),
    .A1(_04518_),
    .S(net103),
    .X(_04529_));
 sg13g2_nand3_1 _09732_ (.B(_04395_),
    .C(_04529_),
    .A(_04528_),
    .Y(_04530_));
 sg13g2_a21oi_1 _09733_ (.A1(_04528_),
    .A2(_04529_),
    .Y(_04531_),
    .B1(_04284_));
 sg13g2_nor3_1 _09734_ (.A(net373),
    .B(_04231_),
    .C(_04531_),
    .Y(_04532_));
 sg13g2_a21oi_1 _09735_ (.A1(net373),
    .A2(_04530_),
    .Y(_04533_),
    .B1(_04532_));
 sg13g2_a21oi_1 _09736_ (.A1(net88),
    .A2(_04527_),
    .Y(_00401_),
    .B1(_04533_));
 sg13g2_nand2_1 _09737_ (.Y(_04534_),
    .A(_04371_),
    .B(_04378_));
 sg13g2_xnor2_1 _09738_ (.Y(_04535_),
    .A(net372),
    .B(_04357_));
 sg13g2_xnor2_1 _09739_ (.Y(_04536_),
    .A(_04534_),
    .B(_04535_));
 sg13g2_nand2_1 _09740_ (.Y(_04537_),
    .A(_02839_),
    .B(net252));
 sg13g2_o21ai_1 _09741_ (.B1(_04537_),
    .Y(_04538_),
    .A1(_01687_),
    .A2(net252));
 sg13g2_a221oi_1 _09742_ (.B2(_04538_),
    .C1(net126),
    .B1(net84),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .Y(_04539_),
    .A2(_02444_));
 sg13g2_o21ai_1 _09743_ (.B1(_02847_),
    .Y(_04540_),
    .A1(_02827_),
    .A2(_04539_));
 sg13g2_nand2_1 _09744_ (.Y(_04541_),
    .A(_04269_),
    .B(_04540_));
 sg13g2_o21ai_1 _09745_ (.B1(_04541_),
    .Y(_04542_),
    .A1(net88),
    .A2(_04536_));
 sg13g2_and2_1 _09746_ (.A(net372),
    .B(_04279_),
    .X(_04543_));
 sg13g2_a21o_1 _09747_ (.A2(_04542_),
    .A1(_04277_),
    .B1(_04543_),
    .X(_00402_));
 sg13g2_nand4_1 _09748_ (.B(_01292_),
    .C(_02883_),
    .A(_01261_),
    .Y(_04544_),
    .D(_02960_));
 sg13g2_nor4_1 _09749_ (.A(net266),
    .B(_01126_),
    .C(net228),
    .D(_01246_),
    .Y(_04545_));
 sg13g2_a21oi_1 _09750_ (.A1(\z80.tv80s.i_tv80_core.PreserveC_r ),
    .A2(net189),
    .Y(_04546_),
    .B1(_04545_));
 sg13g2_nand2_1 _09751_ (.Y(_00403_),
    .A(_04544_),
    .B(_04546_));
 sg13g2_nor2_1 _09752_ (.A(_01606_),
    .B(_01317_),
    .Y(_04547_));
 sg13g2_buf_1 _09753_ (.A(net295),
    .X(_04548_));
 sg13g2_buf_1 _09754_ (.A(net246),
    .X(_04549_));
 sg13g2_nand3_1 _09755_ (.B(_01607_),
    .C(_03998_),
    .A(net212),
    .Y(_04550_));
 sg13g2_buf_1 _09756_ (.A(_04550_),
    .X(_04551_));
 sg13g2_nand2_1 _09757_ (.Y(_04552_),
    .A(_01606_),
    .B(_01320_));
 sg13g2_a21oi_1 _09758_ (.A1(net154),
    .A2(_04552_),
    .Y(_04553_),
    .B1(net225));
 sg13g2_nor2_1 _09759_ (.A(net225),
    .B(_04551_),
    .Y(_04554_));
 sg13g2_nand2_1 _09760_ (.Y(_04555_),
    .A(_01545_),
    .B(_04554_));
 sg13g2_o21ai_1 _09761_ (.B1(_04555_),
    .Y(_00404_),
    .A1(_04547_),
    .A2(_04553_));
 sg13g2_buf_1 _09762_ (.A(net226),
    .X(_04556_));
 sg13g2_buf_1 _09763_ (.A(net154),
    .X(_04557_));
 sg13g2_and3_1 _09764_ (.X(_04558_),
    .A(_01606_),
    .B(\z80.tv80s.i_tv80_core.R[1] ),
    .C(_01320_));
 sg13g2_buf_1 _09765_ (.A(_04558_),
    .X(_04559_));
 sg13g2_nand2_1 _09766_ (.Y(_04560_),
    .A(net150),
    .B(_04559_));
 sg13g2_o21ai_1 _09767_ (.B1(_04560_),
    .Y(_04561_),
    .A1(_01683_),
    .A2(_04557_));
 sg13g2_nor2_1 _09768_ (.A(\z80.tv80s.i_tv80_core.R[1] ),
    .B(_04553_),
    .Y(_04562_));
 sg13g2_a21oi_1 _09769_ (.A1(_04556_),
    .A2(_04561_),
    .Y(_00405_),
    .B1(_04562_));
 sg13g2_nand3_1 _09770_ (.B(net154),
    .C(_04559_),
    .A(_01741_),
    .Y(_04563_));
 sg13g2_o21ai_1 _09771_ (.B1(_04563_),
    .Y(_04564_),
    .A1(_01736_),
    .A2(net150));
 sg13g2_inv_1 _09772_ (.Y(_04565_),
    .A(_04559_));
 sg13g2_a21oi_1 _09773_ (.A1(net150),
    .A2(_04565_),
    .Y(_04566_),
    .B1(_01614_));
 sg13g2_nor2_1 _09774_ (.A(_01741_),
    .B(_04566_),
    .Y(_04567_));
 sg13g2_a21oi_1 _09775_ (.A1(net188),
    .A2(_04564_),
    .Y(_00406_),
    .B1(_04567_));
 sg13g2_nand3_1 _09776_ (.B(\z80.tv80s.i_tv80_core.R[3] ),
    .C(_04559_),
    .A(_01741_),
    .Y(_04568_));
 sg13g2_buf_1 _09777_ (.A(_04568_),
    .X(_04569_));
 sg13g2_nand2b_1 _09778_ (.Y(_04570_),
    .B(net154),
    .A_N(_04569_));
 sg13g2_o21ai_1 _09779_ (.B1(_04570_),
    .Y(_04571_),
    .A1(net379),
    .A2(net150));
 sg13g2_nand2_1 _09780_ (.Y(_04572_),
    .A(_01741_),
    .B(_04559_));
 sg13g2_a21oi_1 _09781_ (.A1(net150),
    .A2(_04572_),
    .Y(_04573_),
    .B1(_01614_));
 sg13g2_nor2_1 _09782_ (.A(\z80.tv80s.i_tv80_core.R[3] ),
    .B(_04573_),
    .Y(_04574_));
 sg13g2_a21oi_1 _09783_ (.A1(net188),
    .A2(_04571_),
    .Y(_00407_),
    .B1(_04574_));
 sg13g2_inv_1 _09784_ (.Y(_04575_),
    .A(\z80.tv80s.i_tv80_core.R[4] ));
 sg13g2_or2_1 _09785_ (.X(_04576_),
    .B(net154),
    .A(_01864_));
 sg13g2_o21ai_1 _09786_ (.B1(_04576_),
    .Y(_04577_),
    .A1(_04575_),
    .A2(_04570_));
 sg13g2_a21o_1 _09787_ (.A2(_04569_),
    .A1(_04557_),
    .B1(net189),
    .X(_04578_));
 sg13g2_a22oi_1 _09788_ (.Y(_00408_),
    .B1(_04578_),
    .B2(_04575_),
    .A2(_04577_),
    .A1(net194));
 sg13g2_nor2_1 _09789_ (.A(_04575_),
    .B(_04569_),
    .Y(_04579_));
 sg13g2_nand3_1 _09790_ (.B(net154),
    .C(_04579_),
    .A(_01954_),
    .Y(_04580_));
 sg13g2_o21ai_1 _09791_ (.B1(_04580_),
    .Y(_04581_),
    .A1(net375),
    .A2(net150));
 sg13g2_o21ai_1 _09792_ (.B1(net154),
    .Y(_04582_),
    .A1(_04575_),
    .A2(_04569_));
 sg13g2_a21oi_1 _09793_ (.A1(net226),
    .A2(_04582_),
    .Y(_04583_),
    .B1(_01954_));
 sg13g2_a21oi_1 _09794_ (.A1(net194),
    .A2(_04581_),
    .Y(_00409_),
    .B1(_04583_));
 sg13g2_nand4_1 _09795_ (.B(\z80.tv80s.i_tv80_core.R[6] ),
    .C(net154),
    .A(_01954_),
    .Y(_04584_),
    .D(_04579_));
 sg13g2_o21ai_1 _09796_ (.B1(_04584_),
    .Y(_04585_),
    .A1(_02007_),
    .A2(net150));
 sg13g2_nand2_1 _09797_ (.Y(_04586_),
    .A(_01954_),
    .B(_04579_));
 sg13g2_a21oi_1 _09798_ (.A1(net150),
    .A2(_04586_),
    .Y(_04587_),
    .B1(net216));
 sg13g2_nor2_1 _09799_ (.A(\z80.tv80s.i_tv80_core.R[6] ),
    .B(_04587_),
    .Y(_04588_));
 sg13g2_a21oi_1 _09800_ (.A1(net194),
    .A2(_04585_),
    .Y(_00410_),
    .B1(_04588_));
 sg13g2_mux2_1 _09801_ (.A0(\z80.tv80s.i_tv80_core.R[7] ),
    .A1(_02076_),
    .S(_04554_),
    .X(_00411_));
 sg13g2_inv_1 _09802_ (.Y(_04589_),
    .A(_01530_));
 sg13g2_buf_1 _09803_ (.A(_01236_),
    .X(_04590_));
 sg13g2_nand2b_1 _09804_ (.Y(_04591_),
    .B(_04239_),
    .A_N(_00023_));
 sg13g2_nand3_1 _09805_ (.B(_01359_),
    .C(_00824_),
    .A(_01071_),
    .Y(_04592_));
 sg13g2_or4_1 _09806_ (.A(net351),
    .B(_01563_),
    .C(_01556_),
    .D(_04239_),
    .X(_04593_));
 sg13g2_nor4_1 _09807_ (.A(_01578_),
    .B(_03486_),
    .C(_02363_),
    .D(_04593_),
    .Y(_04594_));
 sg13g2_nand3_1 _09808_ (.B(_02370_),
    .C(_04594_),
    .A(_01418_),
    .Y(_04595_));
 sg13g2_nand3_1 _09809_ (.B(_04592_),
    .C(_04595_),
    .A(_04591_),
    .Y(_04596_));
 sg13g2_a22oi_1 _09810_ (.Y(_04597_),
    .B1(_04596_),
    .B2(net265),
    .A2(_02104_),
    .A1(net224));
 sg13g2_buf_1 _09811_ (.A(_04597_),
    .X(_04598_));
 sg13g2_nand2_1 _09812_ (.Y(_04599_),
    .A(net94),
    .B(_04598_));
 sg13g2_nand3_1 _09813_ (.B(net211),
    .C(_04599_),
    .A(net100),
    .Y(_04600_));
 sg13g2_o21ai_1 _09814_ (.B1(_04600_),
    .Y(_00412_),
    .A1(_04589_),
    .A2(net194));
 sg13g2_a21oi_1 _09815_ (.A1(_02971_),
    .A2(_04598_),
    .Y(_04601_),
    .B1(_03752_));
 sg13g2_nand2_1 _09816_ (.Y(_04602_),
    .A(net211),
    .B(_04601_));
 sg13g2_o21ai_1 _09817_ (.B1(_04602_),
    .Y(_00413_),
    .A1(_01529_),
    .A2(_02087_));
 sg13g2_a21oi_1 _09818_ (.A1(_02950_),
    .A2(_04598_),
    .Y(_04603_),
    .B1(_03752_));
 sg13g2_mux2_1 _09819_ (.A0(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ),
    .A1(_04603_),
    .S(net227),
    .X(_00414_));
 sg13g2_nand4_1 _09820_ (.B(_01238_),
    .C(_02913_),
    .A(net100),
    .Y(_04604_),
    .D(_04598_));
 sg13g2_o21ai_1 _09821_ (.B1(_04604_),
    .Y(_00415_),
    .A1(_01535_),
    .A2(_02087_));
 sg13g2_inv_1 _09822_ (.Y(_04605_),
    .A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ));
 sg13g2_inv_1 _09823_ (.Y(_04606_),
    .A(_02171_));
 sg13g2_o21ai_1 _09824_ (.B1(net283),
    .Y(_04607_),
    .A1(net214),
    .A2(net239));
 sg13g2_a21oi_1 _09825_ (.A1(_02262_),
    .A2(_04607_),
    .Y(_04608_),
    .B1(_00831_));
 sg13g2_nor3_1 _09826_ (.A(_02267_),
    .B(_04246_),
    .C(_04608_),
    .Y(_04609_));
 sg13g2_nor2_1 _09827_ (.A(_00741_),
    .B(_01330_),
    .Y(_04610_));
 sg13g2_a21oi_1 _09828_ (.A1(net275),
    .A2(_00914_),
    .Y(_04611_),
    .B1(net237));
 sg13g2_o21ai_1 _09829_ (.B1(_00842_),
    .Y(_04612_),
    .A1(_02144_),
    .A2(_04611_));
 sg13g2_nor3_1 _09830_ (.A(_02908_),
    .B(_04610_),
    .C(_04612_),
    .Y(_04613_));
 sg13g2_nor3_1 _09831_ (.A(_00769_),
    .B(_00807_),
    .C(_04613_),
    .Y(_04614_));
 sg13g2_nand4_1 _09832_ (.B(_04606_),
    .C(_04609_),
    .A(_01558_),
    .Y(_04615_),
    .D(_04614_));
 sg13g2_a22oi_1 _09833_ (.Y(_04616_),
    .B1(_04615_),
    .B2(net166),
    .A2(_02233_),
    .A1(_01103_));
 sg13g2_nand2b_1 _09834_ (.Y(_04617_),
    .B(_01278_),
    .A_N(_04616_));
 sg13g2_nor2_1 _09835_ (.A(_02159_),
    .B(net228),
    .Y(_04618_));
 sg13g2_a22oi_1 _09836_ (.Y(_04619_),
    .B1(_04618_),
    .B2(net200),
    .A2(_01364_),
    .A1(_01071_));
 sg13g2_o21ai_1 _09837_ (.B1(_01279_),
    .Y(_04620_),
    .A1(net235),
    .A2(_00981_));
 sg13g2_a22oi_1 _09838_ (.Y(_04621_),
    .B1(_04620_),
    .B2(net219),
    .A2(_01120_),
    .A1(net180));
 sg13g2_o21ai_1 _09839_ (.B1(_04621_),
    .Y(_04622_),
    .A1(net236),
    .A2(_04619_));
 sg13g2_o21ai_1 _09840_ (.B1(_01111_),
    .Y(_04623_),
    .A1(_01412_),
    .A2(_01071_));
 sg13g2_nand3_1 _09841_ (.B(_02090_),
    .C(_04623_),
    .A(_00981_),
    .Y(_04624_));
 sg13g2_nand3_1 _09842_ (.B(_04622_),
    .C(_04624_),
    .A(net224),
    .Y(_04625_));
 sg13g2_nand2_1 _09843_ (.Y(_04626_),
    .A(net231),
    .B(_00730_));
 sg13g2_nand2_1 _09844_ (.Y(_04627_),
    .A(_04626_),
    .B(_02932_));
 sg13g2_a221oi_1 _09845_ (.B2(_01388_),
    .C1(_02926_),
    .B1(_04627_),
    .A1(_01364_),
    .Y(_04628_),
    .A2(_02899_));
 sg13g2_nand3_1 _09846_ (.B(_03407_),
    .C(_04628_),
    .A(_02958_),
    .Y(_04629_));
 sg13g2_o21ai_1 _09847_ (.B1(_01231_),
    .Y(_04630_),
    .A1(_02954_),
    .A2(_04629_));
 sg13g2_nand4_1 _09848_ (.B(_04617_),
    .C(_04625_),
    .A(_04598_),
    .Y(_04631_),
    .D(_04630_));
 sg13g2_nand3_1 _09849_ (.B(_01238_),
    .C(_04631_),
    .A(net100),
    .Y(_04632_));
 sg13g2_o21ai_1 _09850_ (.B1(_04632_),
    .Y(_00416_),
    .A1(_04605_),
    .A2(_01237_));
 sg13g2_nor2_1 _09851_ (.A(_01034_),
    .B(_02950_),
    .Y(_04633_));
 sg13g2_nor2_1 _09852_ (.A(_03850_),
    .B(_04633_),
    .Y(_04634_));
 sg13g2_a22oi_1 _09853_ (.Y(_00417_),
    .B1(_02971_),
    .B2(_04634_),
    .A2(net181),
    .A1(_03157_));
 sg13g2_nand2_1 _09854_ (.Y(_04635_),
    .A(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ),
    .B(_03692_));
 sg13g2_o21ai_1 _09855_ (.B1(_04635_),
    .Y(_00418_),
    .A1(_01960_),
    .A2(_02950_));
 sg13g2_nand2_1 _09856_ (.Y(_04636_),
    .A(_02971_),
    .B(_04633_));
 sg13g2_mux2_1 _09857_ (.A0(_01031_),
    .A1(\z80.tv80s.i_tv80_core.Alternate ),
    .S(_04636_),
    .X(_04637_));
 sg13g2_mux2_1 _09858_ (.A0(\z80.tv80s.i_tv80_core.RegAddrA_r[2] ),
    .A1(_04637_),
    .S(_01237_),
    .X(_00419_));
 sg13g2_a21oi_1 _09859_ (.A1(_02679_),
    .A2(_03512_),
    .Y(_04638_),
    .B1(net106));
 sg13g2_nand2_1 _09860_ (.Y(_04639_),
    .A(_03524_),
    .B(net190));
 sg13g2_o21ai_1 _09861_ (.B1(_04639_),
    .Y(_00420_),
    .A1(net177),
    .A2(_04638_));
 sg13g2_nand2_1 _09862_ (.Y(_04640_),
    .A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .B(net190));
 sg13g2_o21ai_1 _09863_ (.B1(_04640_),
    .Y(_00421_),
    .A1(net177),
    .A2(_03505_));
 sg13g2_nor3_1 _09864_ (.A(_01034_),
    .B(net106),
    .C(_03505_),
    .Y(_04641_));
 sg13g2_mux2_1 _09865_ (.A0(\z80.tv80s.i_tv80_core.Alternate ),
    .A1(_01031_),
    .S(_04641_),
    .X(_04642_));
 sg13g2_mux2_1 _09866_ (.A0(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ),
    .A1(_04642_),
    .S(net211),
    .X(_00422_));
 sg13g2_nor4_1 _09867_ (.A(net305),
    .B(net242),
    .C(_00781_),
    .D(_03739_),
    .Y(_04643_));
 sg13g2_buf_1 _09868_ (.A(_04643_),
    .X(_04644_));
 sg13g2_nor2_1 _09869_ (.A(_02394_),
    .B(net102),
    .Y(_04645_));
 sg13g2_mux2_1 _09870_ (.A0(_02312_),
    .A1(_02333_),
    .S(_04645_),
    .X(_04646_));
 sg13g2_nor2_1 _09871_ (.A(net354),
    .B(_01267_),
    .Y(_04647_));
 sg13g2_a22oi_1 _09872_ (.Y(_00423_),
    .B1(_04646_),
    .B2(_04647_),
    .A2(net181),
    .A1(_02774_));
 sg13g2_inv_1 _09873_ (.Y(_04648_),
    .A(_02485_));
 sg13g2_a22oi_1 _09874_ (.Y(_00424_),
    .B1(_02329_),
    .B2(_04647_),
    .A2(_01277_),
    .A1(_04648_));
 sg13g2_nand2b_1 _09875_ (.Y(_04649_),
    .B(_04645_),
    .A_N(net354));
 sg13g2_nor2b_1 _09876_ (.A(net354),
    .B_N(\z80.tv80s.i_tv80_core.Alternate ),
    .Y(_04650_));
 sg13g2_o21ai_1 _09877_ (.B1(\z80.tv80s.i_tv80_core.XY_State[0] ),
    .Y(_04651_),
    .A1(_02394_),
    .A2(_04644_));
 sg13g2_a22oi_1 _09878_ (.Y(_04652_),
    .B1(_04650_),
    .B2(_04651_),
    .A2(_04649_),
    .A1(_01031_));
 sg13g2_nand2_1 _09879_ (.Y(_04653_),
    .A(_02463_),
    .B(net190));
 sg13g2_o21ai_1 _09880_ (.B1(_04653_),
    .Y(_00425_),
    .A1(net177),
    .A2(_04652_));
 sg13g2_nand2_1 _09881_ (.Y(_04654_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[0] ),
    .B(net190));
 sg13g2_o21ai_1 _09882_ (.B1(_04654_),
    .Y(_00426_),
    .A1(_01960_),
    .A2(_03175_));
 sg13g2_nand2_1 _09883_ (.Y(_04655_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[10] ),
    .B(net190));
 sg13g2_o21ai_1 _09884_ (.B1(_04655_),
    .Y(_00427_),
    .A1(net177),
    .A2(net42));
 sg13g2_nand2_1 _09885_ (.Y(_04656_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[11] ),
    .B(net190));
 sg13g2_o21ai_1 _09886_ (.B1(_04656_),
    .Y(_00428_),
    .A1(net177),
    .A2(_03280_));
 sg13g2_buf_1 _09887_ (.A(net202),
    .X(_04657_));
 sg13g2_nand2_1 _09888_ (.Y(_04658_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[12] ),
    .B(net190));
 sg13g2_o21ai_1 _09889_ (.B1(_04658_),
    .Y(_00429_),
    .A1(net173),
    .A2(_03303_));
 sg13g2_buf_1 _09890_ (.A(net216),
    .X(_04659_));
 sg13g2_nand2_1 _09891_ (.Y(_04660_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[13] ),
    .B(net187));
 sg13g2_o21ai_1 _09892_ (.B1(_04660_),
    .Y(_00430_),
    .A1(net173),
    .A2(net41));
 sg13g2_nand2_1 _09893_ (.Y(_04661_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[14] ),
    .B(net187));
 sg13g2_o21ai_1 _09894_ (.B1(_04661_),
    .Y(_00431_),
    .A1(net173),
    .A2(_03352_));
 sg13g2_nand2_1 _09895_ (.Y(_04662_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[15] ),
    .B(net187));
 sg13g2_o21ai_1 _09896_ (.B1(_04662_),
    .Y(_00432_),
    .A1(net173),
    .A2(_03375_));
 sg13g2_nand2_1 _09897_ (.Y(_04663_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[1] ),
    .B(net187));
 sg13g2_o21ai_1 _09898_ (.B1(_04663_),
    .Y(_00433_),
    .A1(net173),
    .A2(_03212_));
 sg13g2_nand2_1 _09899_ (.Y(_04664_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[2] ),
    .B(net187));
 sg13g2_o21ai_1 _09900_ (.B1(_04664_),
    .Y(_00434_),
    .A1(net173),
    .A2(_04083_));
 sg13g2_nand2_1 _09901_ (.Y(_04665_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[3] ),
    .B(_04659_));
 sg13g2_o21ai_1 _09902_ (.B1(_04665_),
    .Y(_00435_),
    .A1(_04657_),
    .A2(net55));
 sg13g2_nand2_1 _09903_ (.Y(_04666_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[4] ),
    .B(net187));
 sg13g2_o21ai_1 _09904_ (.B1(_04666_),
    .Y(_00436_),
    .A1(net173),
    .A2(_03294_));
 sg13g2_nand2_1 _09905_ (.Y(_04667_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[5] ),
    .B(_04659_));
 sg13g2_o21ai_1 _09906_ (.B1(_04667_),
    .Y(_00437_),
    .A1(_04657_),
    .A2(_03326_));
 sg13g2_nand2_1 _09907_ (.Y(_04668_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[6] ),
    .B(net187));
 sg13g2_o21ai_1 _09908_ (.B1(_04668_),
    .Y(_00438_),
    .A1(net173),
    .A2(_03346_));
 sg13g2_buf_1 _09909_ (.A(net202),
    .X(_04669_));
 sg13g2_nand2_1 _09910_ (.Y(_04670_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[7] ),
    .B(net187));
 sg13g2_o21ai_1 _09911_ (.B1(_04670_),
    .Y(_00439_),
    .A1(_04669_),
    .A2(_03368_));
 sg13g2_buf_1 _09912_ (.A(net216),
    .X(_04671_));
 sg13g2_nand2_1 _09913_ (.Y(_04672_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[8] ),
    .B(net186));
 sg13g2_o21ai_1 _09914_ (.B1(_04672_),
    .Y(_00440_),
    .A1(net172),
    .A2(_04053_));
 sg13g2_nand2_1 _09915_ (.Y(_04673_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[9] ),
    .B(net186));
 sg13g2_o21ai_1 _09916_ (.B1(_04673_),
    .Y(_00441_),
    .A1(net172),
    .A2(net52));
 sg13g2_nand2_1 _09917_ (.Y(_04674_),
    .A(_01529_),
    .B(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ));
 sg13g2_nor2_1 _09918_ (.A(_03699_),
    .B(_04674_),
    .Y(_04675_));
 sg13g2_nand3_1 _09919_ (.B(_01533_),
    .C(_04675_),
    .A(_04589_),
    .Y(_04676_));
 sg13g2_buf_1 _09920_ (.A(_04676_),
    .X(_04677_));
 sg13g2_buf_1 _09921_ (.A(_04677_),
    .X(_04678_));
 sg13g2_nand2_1 _09922_ (.Y(_04679_),
    .A(net238),
    .B(net393));
 sg13g2_a21oi_1 _09923_ (.A1(_01319_),
    .A2(_04679_),
    .Y(_04680_),
    .B1(_03167_));
 sg13g2_o21ai_1 _09924_ (.B1(_01595_),
    .Y(_04681_),
    .A1(_04643_),
    .A2(_04680_));
 sg13g2_buf_1 _09925_ (.A(_04681_),
    .X(_04682_));
 sg13g2_buf_1 _09926_ (.A(_04682_),
    .X(_04683_));
 sg13g2_or4_1 _09927_ (.A(net305),
    .B(net242),
    .C(_00781_),
    .D(_03739_),
    .X(_04684_));
 sg13g2_buf_2 _09928_ (.A(_04684_),
    .X(_04685_));
 sg13g2_nand3_1 _09929_ (.B(net253),
    .C(_04685_),
    .A(_01392_),
    .Y(_04686_));
 sg13g2_o21ai_1 _09930_ (.B1(_04686_),
    .Y(_04687_),
    .A1(_01393_),
    .A2(net253));
 sg13g2_nor2_1 _09931_ (.A(net392),
    .B(_03467_),
    .Y(_04688_));
 sg13g2_a22oi_1 _09932_ (.Y(_04689_),
    .B1(_04688_),
    .B2(_04685_),
    .A2(_04687_),
    .A1(net212));
 sg13g2_buf_1 _09933_ (.A(_04680_),
    .X(_04690_));
 sg13g2_nand2b_1 _09934_ (.Y(_04691_),
    .B(_04690_),
    .A_N(_04689_));
 sg13g2_o21ai_1 _09935_ (.B1(_04691_),
    .Y(_04692_),
    .A1(net253),
    .A2(_04685_));
 sg13g2_a22oi_1 _09936_ (.Y(_04693_),
    .B1(_04692_),
    .B2(_01951_),
    .A2(net75),
    .A1(_03467_));
 sg13g2_nand2_1 _09937_ (.Y(_04694_),
    .A(net162),
    .B(_04693_));
 sg13g2_o21ai_1 _09938_ (.B1(_04694_),
    .Y(_04695_),
    .A1(_01528_),
    .A2(net162));
 sg13g2_nand2_1 _09939_ (.Y(_04696_),
    .A(_00253_),
    .B(net186));
 sg13g2_o21ai_1 _09940_ (.B1(_04696_),
    .Y(_00442_),
    .A1(net172),
    .A2(_04695_));
 sg13g2_inv_1 _09941_ (.Y(_04697_),
    .A(_04682_));
 sg13g2_nor2_1 _09942_ (.A(net198),
    .B(_04685_),
    .Y(_04698_));
 sg13g2_buf_2 _09943_ (.A(_04698_),
    .X(_04699_));
 sg13g2_nand3_1 _09944_ (.B(_01533_),
    .C(_04675_),
    .A(_01530_),
    .Y(_04700_));
 sg13g2_buf_1 _09945_ (.A(_04700_),
    .X(_04701_));
 sg13g2_nand2_1 _09946_ (.Y(_04702_),
    .A(net264),
    .B(_04701_));
 sg13g2_buf_2 _09947_ (.A(_04702_),
    .X(_04703_));
 sg13g2_a21oi_1 _09948_ (.A1(_02404_),
    .A2(_04699_),
    .Y(_04704_),
    .B1(_04703_));
 sg13g2_o21ai_1 _09949_ (.B1(_04704_),
    .Y(_04705_),
    .A1(_03220_),
    .A2(_04697_));
 sg13g2_nor2b_1 _09950_ (.A(net356),
    .B_N(\z80.tv80s.i_tv80_core.SP[10] ),
    .Y(_04706_));
 sg13g2_a21oi_2 _09951_ (.B1(_04706_),
    .Y(_04707_),
    .A2(_02404_),
    .A1(net356));
 sg13g2_nor2b_1 _09952_ (.A(net356),
    .B_N(_02841_),
    .Y(_04708_));
 sg13g2_a21oi_1 _09953_ (.A1(net356),
    .A2(_02826_),
    .Y(_04709_),
    .B1(_04708_));
 sg13g2_nor2_1 _09954_ (.A(net356),
    .B(_02812_),
    .Y(_04710_));
 sg13g2_a21oi_2 _09955_ (.B1(_04710_),
    .Y(_04711_),
    .A2(_02798_),
    .A1(net356));
 sg13g2_nor2_1 _09956_ (.A(net392),
    .B(_04041_),
    .Y(_04712_));
 sg13g2_a21oi_1 _09957_ (.A1(net356),
    .A2(_00158_),
    .Y(_04713_),
    .B1(_04712_));
 sg13g2_buf_2 _09958_ (.A(_04713_),
    .X(_04714_));
 sg13g2_and2_1 _09959_ (.A(net356),
    .B(_02777_),
    .X(_04715_));
 sg13g2_a21oi_2 _09960_ (.B1(_04715_),
    .Y(_04716_),
    .A2(_02766_),
    .A1(net325));
 sg13g2_nor2_1 _09961_ (.A(_04714_),
    .B(_04716_),
    .Y(_04717_));
 sg13g2_nand3b_1 _09962_ (.B(_04711_),
    .C(_04717_),
    .Y(_04718_),
    .A_N(_04709_));
 sg13g2_nand2_1 _09963_ (.Y(_04719_),
    .A(_04707_),
    .B(_04718_));
 sg13g2_or2_1 _09964_ (.X(_04720_),
    .B(_04718_),
    .A(_04707_));
 sg13g2_buf_1 _09965_ (.A(_04720_),
    .X(_04721_));
 sg13g2_o21ai_1 _09966_ (.B1(net325),
    .Y(_04722_),
    .A1(_02710_),
    .A2(_02726_));
 sg13g2_nor2_1 _09967_ (.A(_00152_),
    .B(_02723_),
    .Y(_04723_));
 sg13g2_nor2_1 _09968_ (.A(_02502_),
    .B(_02699_),
    .Y(_04724_));
 sg13g2_o21ai_1 _09969_ (.B1(net295),
    .Y(_04725_),
    .A1(_04723_),
    .A2(_04724_));
 sg13g2_o21ai_1 _09970_ (.B1(_04725_),
    .Y(_04726_),
    .A1(_04023_),
    .A2(_04722_));
 sg13g2_nand2_1 _09971_ (.Y(_04727_),
    .A(net325),
    .B(_02710_));
 sg13g2_o21ai_1 _09972_ (.B1(_04727_),
    .Y(_04728_),
    .A1(net325),
    .A2(_02699_));
 sg13g2_nand3_1 _09973_ (.B(_04015_),
    .C(_04021_),
    .A(_03046_),
    .Y(_04729_));
 sg13g2_o21ai_1 _09974_ (.B1(_04729_),
    .Y(_04730_),
    .A1(net325),
    .A2(_04326_));
 sg13g2_xnor2_1 _09975_ (.Y(_04731_),
    .A(_04728_),
    .B(_04730_));
 sg13g2_o21ai_1 _09976_ (.B1(_04729_),
    .Y(_04732_),
    .A1(net325),
    .A2(_04314_));
 sg13g2_nor2_1 _09977_ (.A(_03046_),
    .B(_01452_),
    .Y(_04733_));
 sg13g2_a21oi_2 _09978_ (.B1(_04688_),
    .Y(_04734_),
    .A2(_04733_),
    .A1(net253));
 sg13g2_a21o_1 _09979_ (.A2(_04734_),
    .A1(_02618_),
    .B1(_02828_),
    .X(_04735_));
 sg13g2_o21ai_1 _09980_ (.B1(_04735_),
    .Y(_04736_),
    .A1(_02618_),
    .A2(_04734_));
 sg13g2_nand2_1 _09981_ (.Y(_04737_),
    .A(_00908_),
    .B(_04736_));
 sg13g2_nand3_1 _09982_ (.B(_04015_),
    .C(_04021_),
    .A(_03467_),
    .Y(_04738_));
 sg13g2_nand3_1 _09983_ (.B(_02630_),
    .C(_04738_),
    .A(_04179_),
    .Y(_04739_));
 sg13g2_a221oi_1 _09984_ (.B2(_04739_),
    .C1(_04712_),
    .B1(_04737_),
    .A1(net392),
    .Y(_04740_),
    .A2(_00143_));
 sg13g2_mux2_1 _09985_ (.A0(_02653_),
    .A1(_02647_),
    .S(net392),
    .X(_04741_));
 sg13g2_buf_1 _09986_ (.A(_04741_),
    .X(_04742_));
 sg13g2_nand2_1 _09987_ (.Y(_04743_),
    .A(_02630_),
    .B(_04742_));
 sg13g2_a22oi_1 _09988_ (.Y(_04744_),
    .B1(_04743_),
    .B2(_03467_),
    .A2(_04021_),
    .A1(_04015_));
 sg13g2_nor2_1 _09989_ (.A(_03467_),
    .B(_04743_),
    .Y(_04745_));
 sg13g2_o21ai_1 _09990_ (.B1(_04179_),
    .Y(_04746_),
    .A1(_04744_),
    .A2(_04745_));
 sg13g2_nand3_1 _09991_ (.B(_04736_),
    .C(_04742_),
    .A(net392),
    .Y(_04747_));
 sg13g2_nand2_1 _09992_ (.Y(_04748_),
    .A(net392),
    .B(_00143_));
 sg13g2_nand3_1 _09993_ (.B(_04748_),
    .C(_04742_),
    .A(_04729_),
    .Y(_04749_));
 sg13g2_nand3_1 _09994_ (.B(_04747_),
    .C(_04749_),
    .A(_04746_),
    .Y(_04750_));
 sg13g2_nor2b_1 _09995_ (.A(net392),
    .B_N(_02681_),
    .Y(_04751_));
 sg13g2_a21oi_1 _09996_ (.A1(net392),
    .A2(_02671_),
    .Y(_04752_),
    .B1(_04751_));
 sg13g2_inv_1 _09997_ (.Y(_04753_),
    .A(_04752_));
 sg13g2_nor3_1 _09998_ (.A(_04740_),
    .B(_04750_),
    .C(_04753_),
    .Y(_04754_));
 sg13g2_o21ai_1 _09999_ (.B1(_04753_),
    .Y(_04755_),
    .A1(_04740_),
    .A2(_04750_));
 sg13g2_o21ai_1 _10000_ (.B1(_04755_),
    .Y(_04756_),
    .A1(_04732_),
    .A2(_04754_));
 sg13g2_and2_1 _10001_ (.A(_04731_),
    .B(_04756_),
    .X(_04757_));
 sg13g2_nor2_1 _10002_ (.A(_04323_),
    .B(_02725_),
    .Y(_04758_));
 sg13g2_nor2_1 _10003_ (.A(net295),
    .B(_02726_),
    .Y(_04759_));
 sg13g2_a22oi_1 _10004_ (.Y(_04760_),
    .B1(_04759_),
    .B2(_04024_),
    .A2(_04758_),
    .A1(net295));
 sg13g2_o21ai_1 _10005_ (.B1(_04760_),
    .Y(_04761_),
    .A1(_04726_),
    .A2(_04757_));
 sg13g2_buf_2 _10006_ (.A(_04761_),
    .X(_04762_));
 sg13g2_inv_1 _10007_ (.Y(_04763_),
    .A(_02757_));
 sg13g2_o21ai_1 _10008_ (.B1(_04763_),
    .Y(_04764_),
    .A1(net117),
    .A2(_04762_));
 sg13g2_a21oi_1 _10009_ (.A1(net117),
    .A2(_04762_),
    .Y(_04765_),
    .B1(net246));
 sg13g2_o21ai_1 _10010_ (.B1(_02566_),
    .Y(_04766_),
    .A1(_02747_),
    .A2(_04762_));
 sg13g2_a21oi_1 _10011_ (.A1(_02747_),
    .A2(_04762_),
    .Y(_04767_),
    .B1(net288));
 sg13g2_a22oi_1 _10012_ (.Y(_04768_),
    .B1(_04766_),
    .B2(_04767_),
    .A2(_04765_),
    .A1(_04764_));
 sg13g2_buf_1 _10013_ (.A(_04768_),
    .X(_04769_));
 sg13g2_buf_1 _10014_ (.A(_04769_),
    .X(_04770_));
 sg13g2_a21o_1 _10015_ (.A2(_04721_),
    .A1(_04719_),
    .B1(net40),
    .X(_04771_));
 sg13g2_nor2b_1 _10016_ (.A(_04711_),
    .B_N(_04716_),
    .Y(_04772_));
 sg13g2_and3_1 _10017_ (.X(_04773_),
    .A(_04709_),
    .B(_04714_),
    .C(_04772_));
 sg13g2_buf_1 _10018_ (.A(_04773_),
    .X(_04774_));
 sg13g2_nand3b_1 _10019_ (.B(net40),
    .C(_04707_),
    .Y(_04775_),
    .A_N(_04774_));
 sg13g2_nand3b_1 _10020_ (.B(net40),
    .C(_04774_),
    .Y(_04776_),
    .A_N(_04707_));
 sg13g2_nand3_1 _10021_ (.B(_04685_),
    .C(net101),
    .A(net169),
    .Y(_04777_));
 sg13g2_inv_1 _10022_ (.Y(_04778_),
    .A(_04777_));
 sg13g2_and4_1 _10023_ (.A(_04771_),
    .B(_04775_),
    .C(_04776_),
    .D(_04778_),
    .X(_04779_));
 sg13g2_nor2_1 _10024_ (.A(_01244_),
    .B(_04701_),
    .Y(_04780_));
 sg13g2_buf_2 _10025_ (.A(_04780_),
    .X(_04781_));
 sg13g2_a22oi_1 _10026_ (.Y(_04782_),
    .B1(_01735_),
    .B2(_04781_),
    .A2(net189),
    .A1(_00254_));
 sg13g2_o21ai_1 _10027_ (.B1(_04782_),
    .Y(_00443_),
    .A1(_04705_),
    .A2(_04779_));
 sg13g2_a22oi_1 _10028_ (.Y(_04783_),
    .B1(_01802_),
    .B2(_04781_),
    .A2(net222),
    .A1(_00255_));
 sg13g2_a221oi_1 _10029_ (.B2(_02464_),
    .C1(_04703_),
    .B1(_04699_),
    .A1(_02472_),
    .Y(_04784_),
    .A2(net75));
 sg13g2_inv_1 _10030_ (.Y(_04785_),
    .A(_04784_));
 sg13g2_nor2_1 _10031_ (.A(net325),
    .B(_02454_),
    .Y(_04786_));
 sg13g2_a21oi_2 _10032_ (.B1(_04786_),
    .Y(_04787_),
    .A2(_02472_),
    .A1(net288));
 sg13g2_nand2_1 _10033_ (.Y(_04788_),
    .A(_04707_),
    .B(_04774_));
 sg13g2_mux2_1 _10034_ (.A0(_04721_),
    .A1(_04788_),
    .S(_04769_),
    .X(_04789_));
 sg13g2_xor2_1 _10035_ (.B(_04789_),
    .A(_04787_),
    .X(_04790_));
 sg13g2_and2_1 _10036_ (.A(_04778_),
    .B(_04783_),
    .X(_04791_));
 sg13g2_a22oi_1 _10037_ (.Y(_00444_),
    .B1(_04790_),
    .B2(_04791_),
    .A2(_04785_),
    .A1(_04783_));
 sg13g2_a22oi_1 _10038_ (.Y(_04792_),
    .B1(_01863_),
    .B2(_04781_),
    .A2(net222),
    .A1(_00256_));
 sg13g2_a221oi_1 _10039_ (.B2(_02508_),
    .C1(_04703_),
    .B1(_04699_),
    .A1(_02509_),
    .Y(_04793_),
    .A2(net75));
 sg13g2_inv_1 _10040_ (.Y(_04794_),
    .A(_04793_));
 sg13g2_nor2_1 _10041_ (.A(net288),
    .B(_02490_),
    .Y(_04795_));
 sg13g2_a21oi_2 _10042_ (.B1(_04795_),
    .Y(_04796_),
    .A2(_02509_),
    .A1(net288));
 sg13g2_inv_1 _10043_ (.Y(_04797_),
    .A(_04796_));
 sg13g2_or2_1 _10044_ (.X(_04798_),
    .B(_04787_),
    .A(_04721_));
 sg13g2_buf_1 _10045_ (.A(_04798_),
    .X(_04799_));
 sg13g2_nand3_1 _10046_ (.B(_04774_),
    .C(_04787_),
    .A(_04707_),
    .Y(_04800_));
 sg13g2_mux2_1 _10047_ (.A0(_04799_),
    .A1(_04800_),
    .S(net40),
    .X(_04801_));
 sg13g2_xnor2_1 _10048_ (.Y(_04802_),
    .A(_04797_),
    .B(_04801_));
 sg13g2_and2_1 _10049_ (.A(_04778_),
    .B(_04792_),
    .X(_04803_));
 sg13g2_a22oi_1 _10050_ (.Y(_00445_),
    .B1(_04802_),
    .B2(_04803_),
    .A2(_04794_),
    .A1(_04792_));
 sg13g2_nor2b_1 _10051_ (.A(net295),
    .B_N(_02540_),
    .Y(_04804_));
 sg13g2_a21oi_1 _10052_ (.A1(net246),
    .A2(_02523_),
    .Y(_04805_),
    .B1(_04804_));
 sg13g2_buf_1 _10053_ (.A(_04805_),
    .X(_04806_));
 sg13g2_o21ai_1 _10054_ (.B1(_04806_),
    .Y(_04807_),
    .A1(_04799_),
    .A2(_04796_));
 sg13g2_nor2_1 _10055_ (.A(_04799_),
    .B(_04796_),
    .Y(_04808_));
 sg13g2_nand2b_1 _10056_ (.Y(_04809_),
    .B(_04808_),
    .A_N(_04806_));
 sg13g2_a21o_1 _10057_ (.A2(_04809_),
    .A1(_04807_),
    .B1(net40),
    .X(_04810_));
 sg13g2_nor2_1 _10058_ (.A(_04797_),
    .B(_04800_),
    .Y(_04811_));
 sg13g2_nor2b_1 _10059_ (.A(_04811_),
    .B_N(_04806_),
    .Y(_04812_));
 sg13g2_nor3_1 _10060_ (.A(_04797_),
    .B(_04800_),
    .C(_04806_),
    .Y(_04813_));
 sg13g2_o21ai_1 _10061_ (.B1(net40),
    .Y(_04814_),
    .A1(_04812_),
    .A2(_04813_));
 sg13g2_a21oi_1 _10062_ (.A1(_02523_),
    .A2(_04699_),
    .Y(_04815_),
    .B1(_04703_));
 sg13g2_nand3_1 _10063_ (.B(net101),
    .C(_04815_),
    .A(net159),
    .Y(_04816_));
 sg13g2_a21oi_1 _10064_ (.A1(_04810_),
    .A2(_04814_),
    .Y(_04817_),
    .B1(_04816_));
 sg13g2_nand2_1 _10065_ (.Y(_04818_),
    .A(_02540_),
    .B(net179));
 sg13g2_nand2_1 _10066_ (.Y(_04819_),
    .A(net169),
    .B(_02523_));
 sg13g2_nand4_1 _10067_ (.B(_04701_),
    .C(_04818_),
    .A(net102),
    .Y(_04820_),
    .D(_04819_));
 sg13g2_o21ai_1 _10068_ (.B1(_04820_),
    .Y(_04821_),
    .A1(_01947_),
    .A2(_04701_));
 sg13g2_a21oi_1 _10069_ (.A1(net168),
    .A2(net101),
    .Y(_04822_),
    .B1(_02540_));
 sg13g2_and2_1 _10070_ (.A(_00257_),
    .B(net225),
    .X(_04823_));
 sg13g2_a221oi_1 _10071_ (.B2(_04822_),
    .C1(_04823_),
    .B1(_04815_),
    .A1(net226),
    .Y(_04824_),
    .A2(_04821_));
 sg13g2_nand2b_1 _10072_ (.Y(_00446_),
    .B(_04824_),
    .A_N(_04817_));
 sg13g2_a21oi_1 _10073_ (.A1(net168),
    .A2(net101),
    .Y(_04825_),
    .B1(_02572_));
 sg13g2_nor2_1 _10074_ (.A(net102),
    .B(_04703_),
    .Y(_04826_));
 sg13g2_inv_1 _10075_ (.Y(_04827_),
    .A(_04826_));
 sg13g2_inv_1 _10076_ (.Y(_04828_),
    .A(_00258_));
 sg13g2_nand2_1 _10077_ (.Y(_04829_),
    .A(_02572_),
    .B(net198));
 sg13g2_nand3_1 _10078_ (.B(_02556_),
    .C(net102),
    .A(net178),
    .Y(_04830_));
 sg13g2_a21oi_1 _10079_ (.A1(_04829_),
    .A2(_04830_),
    .Y(_04831_),
    .B1(_04703_));
 sg13g2_a221oi_1 _10080_ (.B2(_04781_),
    .C1(_04831_),
    .B1(_02006_),
    .A1(_04828_),
    .Y(_04832_),
    .A2(net263));
 sg13g2_o21ai_1 _10081_ (.B1(_04832_),
    .Y(_04833_),
    .A1(_04825_),
    .A2(_04827_));
 sg13g2_nand2_1 _10082_ (.Y(_04834_),
    .A(_04806_),
    .B(_04811_));
 sg13g2_mux2_1 _10083_ (.A0(_04809_),
    .A1(_04834_),
    .S(_04769_),
    .X(_04835_));
 sg13g2_nor2b_1 _10084_ (.A(net246),
    .B_N(_02572_),
    .Y(_04836_));
 sg13g2_a21oi_2 _10085_ (.B1(_04836_),
    .Y(_04837_),
    .A2(_02556_),
    .A1(net212));
 sg13g2_nand3b_1 _10086_ (.B(net101),
    .C(_04832_),
    .Y(_04838_),
    .A_N(_04837_));
 sg13g2_or2_1 _10087_ (.X(_04839_),
    .B(_04838_),
    .A(_04835_));
 sg13g2_nand4_1 _10088_ (.B(_04832_),
    .C(_04835_),
    .A(net101),
    .Y(_04840_),
    .D(_04837_));
 sg13g2_nand3_1 _10089_ (.B(_04839_),
    .C(_04840_),
    .A(_04833_),
    .Y(_00447_));
 sg13g2_a22oi_1 _10090_ (.Y(_04841_),
    .B1(_04699_),
    .B2(_02588_),
    .A2(_04682_),
    .A1(_03358_));
 sg13g2_nand2_1 _10091_ (.Y(_04842_),
    .A(_04701_),
    .B(_04841_));
 sg13g2_o21ai_1 _10092_ (.B1(_04842_),
    .Y(_04843_),
    .A1(_02075_),
    .A2(_04701_));
 sg13g2_nand2_1 _10093_ (.Y(_04844_),
    .A(net226),
    .B(_04843_));
 sg13g2_o21ai_1 _10094_ (.B1(_04844_),
    .Y(_04845_),
    .A1(_00259_),
    .A2(net211));
 sg13g2_nor2_1 _10095_ (.A(net288),
    .B(_02588_),
    .Y(_04846_));
 sg13g2_a21o_1 _10096_ (.A2(_02593_),
    .A1(net288),
    .B1(_04846_),
    .X(_04847_));
 sg13g2_nand2_1 _10097_ (.Y(_04848_),
    .A(_02593_),
    .B(net179));
 sg13g2_nand4_1 _10098_ (.B(_04826_),
    .C(_04847_),
    .A(net101),
    .Y(_04849_),
    .D(_04848_));
 sg13g2_a21oi_1 _10099_ (.A1(net288),
    .A2(_02593_),
    .Y(_04850_),
    .B1(_04846_));
 sg13g2_nand4_1 _10100_ (.B(_04826_),
    .C(_04850_),
    .A(net101),
    .Y(_04851_),
    .D(_04848_));
 sg13g2_nor3_1 _10101_ (.A(_04714_),
    .B(_04806_),
    .C(_04837_),
    .Y(_04852_));
 sg13g2_nand2_1 _10102_ (.Y(_04853_),
    .A(_04808_),
    .B(_04852_));
 sg13g2_nand3_1 _10103_ (.B(_04811_),
    .C(_04837_),
    .A(_04806_),
    .Y(_04854_));
 sg13g2_mux2_1 _10104_ (.A0(_04853_),
    .A1(_04854_),
    .S(net40),
    .X(_04855_));
 sg13g2_mux2_1 _10105_ (.A0(_04849_),
    .A1(_04851_),
    .S(_04855_),
    .X(_04856_));
 sg13g2_nand2_1 _10106_ (.Y(_00448_),
    .A(_04845_),
    .B(_04856_));
 sg13g2_and2_1 _10107_ (.A(_04685_),
    .B(_04690_),
    .X(_04857_));
 sg13g2_buf_2 _10108_ (.A(_04857_),
    .X(_04858_));
 sg13g2_xnor2_1 _10109_ (.Y(_04859_),
    .A(_02630_),
    .B(net117));
 sg13g2_xnor2_1 _10110_ (.Y(_04860_),
    .A(_02828_),
    .B(_02618_));
 sg13g2_nand2_1 _10111_ (.Y(_04861_),
    .A(_04548_),
    .B(_04860_));
 sg13g2_o21ai_1 _10112_ (.B1(_04861_),
    .Y(_04862_),
    .A1(net212),
    .A2(_04859_));
 sg13g2_xor2_1 _10113_ (.B(_04862_),
    .A(_04734_),
    .X(_04863_));
 sg13g2_nand2_1 _10114_ (.Y(_04864_),
    .A(_04858_),
    .B(_04863_));
 sg13g2_o21ai_1 _10115_ (.B1(_04864_),
    .Y(_04865_),
    .A1(_02618_),
    .A2(_04685_));
 sg13g2_a22oi_1 _10116_ (.Y(_04866_),
    .B1(_04865_),
    .B2(net158),
    .A2(net75),
    .A1(_02630_));
 sg13g2_nor2_1 _10117_ (.A(_01681_),
    .B(net162),
    .Y(_04867_));
 sg13g2_a21oi_1 _10118_ (.A1(_04678_),
    .A2(_04866_),
    .Y(_04868_),
    .B1(_04867_));
 sg13g2_nand2_1 _10119_ (.Y(_04869_),
    .A(_00260_),
    .B(net186));
 sg13g2_o21ai_1 _10120_ (.B1(_04869_),
    .Y(_00449_),
    .A1(net172),
    .A2(_04868_));
 sg13g2_nand2_1 _10121_ (.Y(_04870_),
    .A(_04737_),
    .B(_04739_));
 sg13g2_nor3_1 _10122_ (.A(_02294_),
    .B(net117),
    .C(_04870_),
    .Y(_04871_));
 sg13g2_a21oi_1 _10123_ (.A1(net117),
    .A2(_04870_),
    .Y(_04872_),
    .B1(_04871_));
 sg13g2_xnor2_1 _10124_ (.Y(_04873_),
    .A(_04307_),
    .B(_04870_));
 sg13g2_mux2_1 _10125_ (.A0(_04872_),
    .A1(_04873_),
    .S(net246),
    .X(_04874_));
 sg13g2_xnor2_1 _10126_ (.Y(_04875_),
    .A(_04742_),
    .B(_04874_));
 sg13g2_a22oi_1 _10127_ (.Y(_04876_),
    .B1(_04858_),
    .B2(_04875_),
    .A2(_04644_),
    .A1(_02647_));
 sg13g2_inv_1 _10128_ (.Y(_04877_),
    .A(_04876_));
 sg13g2_a22oi_1 _10129_ (.Y(_04878_),
    .B1(_04877_),
    .B2(net158),
    .A2(net75),
    .A1(_02653_));
 sg13g2_nor2_1 _10130_ (.A(_01734_),
    .B(_04678_),
    .Y(_04879_));
 sg13g2_a21oi_1 _10131_ (.A1(net162),
    .A2(_04878_),
    .Y(_04880_),
    .B1(_04879_));
 sg13g2_nand2_1 _10132_ (.Y(_04881_),
    .A(_00261_),
    .B(_04671_));
 sg13g2_o21ai_1 _10133_ (.B1(_04881_),
    .Y(_00450_),
    .A1(net172),
    .A2(_04880_));
 sg13g2_nor2_1 _10134_ (.A(_04740_),
    .B(_04750_),
    .Y(_04882_));
 sg13g2_xnor2_1 _10135_ (.Y(_04883_),
    .A(_04753_),
    .B(_04732_));
 sg13g2_xnor2_1 _10136_ (.Y(_04884_),
    .A(_04882_),
    .B(_04883_));
 sg13g2_a22oi_1 _10137_ (.Y(_04885_),
    .B1(_04858_),
    .B2(_04884_),
    .A2(net102),
    .A1(_02671_));
 sg13g2_inv_1 _10138_ (.Y(_04886_),
    .A(_04885_));
 sg13g2_a22oi_1 _10139_ (.Y(_04887_),
    .B1(_04886_),
    .B2(net158),
    .A2(_04683_),
    .A1(_02681_));
 sg13g2_nor2_1 _10140_ (.A(_01801_),
    .B(_04677_),
    .Y(_04888_));
 sg13g2_a21oi_1 _10141_ (.A1(net162),
    .A2(_04887_),
    .Y(_04889_),
    .B1(_04888_));
 sg13g2_nand2_1 _10142_ (.Y(_04890_),
    .A(_00262_),
    .B(net186));
 sg13g2_o21ai_1 _10143_ (.B1(_04890_),
    .Y(_00451_),
    .A1(_04669_),
    .A2(_04889_));
 sg13g2_xnor2_1 _10144_ (.Y(_04891_),
    .A(_04731_),
    .B(_04756_));
 sg13g2_nand2b_1 _10145_ (.Y(_04892_),
    .B(_04858_),
    .A_N(_04891_));
 sg13g2_o21ai_1 _10146_ (.B1(_04892_),
    .Y(_04893_),
    .A1(_02699_),
    .A2(_04685_));
 sg13g2_a22oi_1 _10147_ (.Y(_04894_),
    .B1(_04893_),
    .B2(net158),
    .A2(_04683_),
    .A1(_02710_));
 sg13g2_nor2_1 _10148_ (.A(_03877_),
    .B(_04677_),
    .Y(_04895_));
 sg13g2_a21oi_1 _10149_ (.A1(net162),
    .A2(_04894_),
    .Y(_04896_),
    .B1(_04895_));
 sg13g2_nand2_1 _10150_ (.Y(_04897_),
    .A(_00263_),
    .B(net186));
 sg13g2_o21ai_1 _10151_ (.B1(_04897_),
    .Y(_00452_),
    .A1(net172),
    .A2(_04896_));
 sg13g2_o21ai_1 _10152_ (.B1(_02502_),
    .Y(_04898_),
    .A1(_00146_),
    .A2(_04754_));
 sg13g2_o21ai_1 _10153_ (.B1(_04755_),
    .Y(_04899_),
    .A1(net295),
    .A2(_04024_));
 sg13g2_a21o_1 _10154_ (.A2(_04898_),
    .A1(net295),
    .B1(_04899_),
    .X(_04900_));
 sg13g2_a21oi_1 _10155_ (.A1(_00146_),
    .A2(_04755_),
    .Y(_04901_),
    .B1(_02502_));
 sg13g2_nand2b_1 _10156_ (.Y(_04902_),
    .B(net246),
    .A_N(_04901_));
 sg13g2_nor2_1 _10157_ (.A(_04712_),
    .B(_04754_),
    .Y(_04903_));
 sg13g2_a22oi_1 _10158_ (.Y(_04904_),
    .B1(_04902_),
    .B2(_04903_),
    .A2(_04900_),
    .A1(_04728_));
 sg13g2_xnor2_1 _10159_ (.Y(_04905_),
    .A(_02726_),
    .B(net117));
 sg13g2_o21ai_1 _10160_ (.B1(_04548_),
    .Y(_04906_),
    .A1(_04758_),
    .A2(_04723_));
 sg13g2_o21ai_1 _10161_ (.B1(_04906_),
    .Y(_04907_),
    .A1(net212),
    .A2(_04905_));
 sg13g2_xnor2_1 _10162_ (.Y(_04908_),
    .A(_04904_),
    .B(_04907_));
 sg13g2_a22oi_1 _10163_ (.Y(_04909_),
    .B1(_04858_),
    .B2(_04908_),
    .A2(net102),
    .A1(_02723_));
 sg13g2_nor2_1 _10164_ (.A(net164),
    .B(_04909_),
    .Y(_04910_));
 sg13g2_o21ai_1 _10165_ (.B1(_04677_),
    .Y(_04911_),
    .A1(_02726_),
    .A2(_04697_));
 sg13g2_nand2b_1 _10166_ (.Y(_04912_),
    .B(_01947_),
    .A_N(_04677_));
 sg13g2_o21ai_1 _10167_ (.B1(_04912_),
    .Y(_04913_),
    .A1(_04910_),
    .A2(_04911_));
 sg13g2_nand2_1 _10168_ (.Y(_04914_),
    .A(_00264_),
    .B(net186));
 sg13g2_o21ai_1 _10169_ (.B1(_04914_),
    .Y(_00453_),
    .A1(net172),
    .A2(_04913_));
 sg13g2_xnor2_1 _10170_ (.Y(_04915_),
    .A(_02757_),
    .B(net117));
 sg13g2_xnor2_1 _10171_ (.Y(_04916_),
    .A(_02566_),
    .B(_02747_));
 sg13g2_nand2_1 _10172_ (.Y(_04917_),
    .A(net246),
    .B(_04916_));
 sg13g2_o21ai_1 _10173_ (.B1(_04917_),
    .Y(_04918_),
    .A1(net212),
    .A2(_04915_));
 sg13g2_xor2_1 _10174_ (.B(_04918_),
    .A(_04762_),
    .X(_04919_));
 sg13g2_a22oi_1 _10175_ (.Y(_04920_),
    .B1(_04858_),
    .B2(_04919_),
    .A2(net102),
    .A1(_02756_));
 sg13g2_nand2_1 _10176_ (.Y(_04921_),
    .A(_02757_),
    .B(net75));
 sg13g2_o21ai_1 _10177_ (.B1(_04921_),
    .Y(_04922_),
    .A1(net179),
    .A2(_04920_));
 sg13g2_mux2_1 _10178_ (.A0(_02006_),
    .A1(_04922_),
    .S(net162),
    .X(_04923_));
 sg13g2_nand2_1 _10179_ (.Y(_04924_),
    .A(_00265_),
    .B(net186));
 sg13g2_o21ai_1 _10180_ (.B1(_04924_),
    .Y(_00454_),
    .A1(net172),
    .A2(_04923_));
 sg13g2_xnor2_1 _10181_ (.Y(_04925_),
    .A(_04714_),
    .B(_04716_));
 sg13g2_xnor2_1 _10182_ (.Y(_04926_),
    .A(_04770_),
    .B(_04925_));
 sg13g2_nand2_1 _10183_ (.Y(_04927_),
    .A(_02766_),
    .B(_04682_));
 sg13g2_nand3_1 _10184_ (.B(_04677_),
    .C(_04927_),
    .A(net264),
    .Y(_04928_));
 sg13g2_a221oi_1 _10185_ (.B2(_04926_),
    .C1(_04928_),
    .B1(_04858_),
    .A1(_02777_),
    .Y(_04929_),
    .A2(net102));
 sg13g2_nor2_1 _10186_ (.A(net216),
    .B(net162),
    .Y(_04930_));
 sg13g2_a22oi_1 _10187_ (.Y(_04931_),
    .B1(_02075_),
    .B2(_04930_),
    .A2(net189),
    .A1(_00266_));
 sg13g2_or2_1 _10188_ (.X(_04932_),
    .B(_04928_),
    .A(net159));
 sg13g2_nand3b_1 _10189_ (.B(_04931_),
    .C(_04932_),
    .Y(_00455_),
    .A_N(_04929_));
 sg13g2_a22oi_1 _10190_ (.Y(_04933_),
    .B1(_01528_),
    .B2(_04781_),
    .A2(net222),
    .A1(_00267_));
 sg13g2_a221oi_1 _10191_ (.B2(_02797_),
    .C1(_04703_),
    .B1(_04699_),
    .A1(_02812_),
    .Y(_04934_),
    .A2(net75));
 sg13g2_inv_1 _10192_ (.Y(_04935_),
    .A(_04934_));
 sg13g2_or2_1 _10193_ (.X(_04936_),
    .B(_04716_),
    .A(_04714_));
 sg13g2_nand2_1 _10194_ (.Y(_04937_),
    .A(_04714_),
    .B(_04716_));
 sg13g2_mux2_1 _10195_ (.A0(_04936_),
    .A1(_04937_),
    .S(_04769_),
    .X(_04938_));
 sg13g2_xnor2_1 _10196_ (.Y(_04939_),
    .A(_04711_),
    .B(_04938_));
 sg13g2_and2_1 _10197_ (.A(_04778_),
    .B(_04933_),
    .X(_04940_));
 sg13g2_a22oi_1 _10198_ (.Y(_00456_),
    .B1(_04939_),
    .B2(_04940_),
    .A2(_04935_),
    .A1(_04933_));
 sg13g2_a221oi_1 _10199_ (.B2(_02826_),
    .C1(_04703_),
    .B1(_04699_),
    .A1(_02841_),
    .Y(_04941_),
    .A2(net75));
 sg13g2_a22oi_1 _10200_ (.Y(_04942_),
    .B1(_01682_),
    .B2(_04781_),
    .A2(net222),
    .A1(_00268_));
 sg13g2_nand2b_1 _10201_ (.Y(_04943_),
    .B(_04942_),
    .A_N(_04941_));
 sg13g2_a221oi_1 _10202_ (.B2(_04772_),
    .C1(_04708_),
    .B1(_04714_),
    .A1(net212),
    .Y(_04944_),
    .A2(_02826_));
 sg13g2_nor3_1 _10203_ (.A(_04709_),
    .B(_04711_),
    .C(_04937_),
    .Y(_04945_));
 sg13g2_o21ai_1 _10204_ (.B1(_04770_),
    .Y(_04946_),
    .A1(_04944_),
    .A2(_04945_));
 sg13g2_nand2_1 _10205_ (.Y(_04947_),
    .A(_04711_),
    .B(_04717_));
 sg13g2_nand2_1 _10206_ (.Y(_04948_),
    .A(_04709_),
    .B(_04947_));
 sg13g2_a21o_1 _10207_ (.A2(_04948_),
    .A1(_04718_),
    .B1(net40),
    .X(_04949_));
 sg13g2_nand4_1 _10208_ (.B(_04942_),
    .C(_04946_),
    .A(_04778_),
    .Y(_04950_),
    .D(_04949_));
 sg13g2_and2_1 _10209_ (.A(_04943_),
    .B(_04950_),
    .X(_00457_));
 sg13g2_nand2_1 _10210_ (.Y(_04951_),
    .A(_02920_),
    .B(_03407_));
 sg13g2_nor2_1 _10211_ (.A(_00959_),
    .B(_02122_),
    .Y(_04952_));
 sg13g2_nand2_1 _10212_ (.Y(_04953_),
    .A(_01141_),
    .B(net175));
 sg13g2_nand4_1 _10213_ (.B(_04952_),
    .C(_02880_),
    .A(_00720_),
    .Y(_04954_),
    .D(_04953_));
 sg13g2_or2_1 _10214_ (.X(_04955_),
    .B(_04954_),
    .A(_02119_));
 sg13g2_mux2_1 _10215_ (.A0(_02922_),
    .A1(_04951_),
    .S(_04955_),
    .X(_04956_));
 sg13g2_a21oi_1 _10216_ (.A1(_01231_),
    .A2(_04956_),
    .Y(_04957_),
    .B1(net224));
 sg13g2_o21ai_1 _10217_ (.B1(_02202_),
    .Y(_04958_),
    .A1(_01126_),
    .A2(net228));
 sg13g2_inv_1 _10218_ (.Y(_04959_),
    .A(_04958_));
 sg13g2_a221oi_1 _10219_ (.B2(_04621_),
    .C1(_02142_),
    .B1(_04959_),
    .A1(_04617_),
    .Y(_04960_),
    .A2(_04957_));
 sg13g2_a21o_1 _10220_ (.A2(_01615_),
    .A1(net343),
    .B1(_04960_),
    .X(_00458_));
 sg13g2_o21ai_1 _10221_ (.B1(_02900_),
    .Y(_04961_),
    .A1(net201),
    .A2(_02254_));
 sg13g2_o21ai_1 _10222_ (.B1(net301),
    .Y(_04962_),
    .A1(_04241_),
    .A2(_04961_));
 sg13g2_o21ai_1 _10223_ (.B1(net224),
    .Y(_04963_),
    .A1(_01124_),
    .A2(_01167_));
 sg13g2_nand2_1 _10224_ (.Y(_04964_),
    .A(_04962_),
    .B(_04963_));
 sg13g2_nor2_1 _10225_ (.A(net201),
    .B(_01369_),
    .Y(_04965_));
 sg13g2_nand4_1 _10226_ (.B(_01292_),
    .C(_02254_),
    .A(_01289_),
    .Y(_04966_),
    .D(_02900_));
 sg13g2_nor4_1 _10227_ (.A(_01578_),
    .B(_03486_),
    .C(_04965_),
    .D(_04966_),
    .Y(_04967_));
 sg13g2_nor3_1 _10228_ (.A(_01061_),
    .B(_02300_),
    .C(_04251_),
    .Y(_04968_));
 sg13g2_a22oi_1 _10229_ (.Y(_04969_),
    .B1(_04967_),
    .B2(_04968_),
    .A2(_04964_),
    .A1(net206));
 sg13g2_nor2_2 _10230_ (.A(net288),
    .B(_04969_),
    .Y(_04970_));
 sg13g2_buf_1 _10231_ (.A(_04970_),
    .X(_04971_));
 sg13g2_nor2_1 _10232_ (.A(_01319_),
    .B(_03984_),
    .Y(_04972_));
 sg13g2_and2_1 _10233_ (.A(_03987_),
    .B(_04972_),
    .X(_04973_));
 sg13g2_buf_2 _10234_ (.A(_04973_),
    .X(_04974_));
 sg13g2_nand2_1 _10235_ (.Y(_04975_),
    .A(_01003_),
    .B(net295));
 sg13g2_buf_1 _10236_ (.A(_04975_),
    .X(_04976_));
 sg13g2_or2_1 _10237_ (.X(_04977_),
    .B(_02371_),
    .A(_01319_));
 sg13g2_buf_2 _10238_ (.A(_04977_),
    .X(_04978_));
 sg13g2_and2_1 _10239_ (.A(_04976_),
    .B(_04978_),
    .X(_04979_));
 sg13g2_buf_1 _10240_ (.A(_04979_),
    .X(_04980_));
 sg13g2_nand2_1 _10241_ (.Y(_04981_),
    .A(_01594_),
    .B(_04980_));
 sg13g2_o21ai_1 _10242_ (.B1(_04981_),
    .Y(_04982_),
    .A1(net178),
    .A2(_04974_));
 sg13g2_buf_1 _10243_ (.A(_04982_),
    .X(_04983_));
 sg13g2_inv_1 _10244_ (.Y(_04984_),
    .A(_04983_));
 sg13g2_o21ai_1 _10245_ (.B1(net226),
    .Y(_04985_),
    .A1(net132),
    .A2(_04984_));
 sg13g2_and2_1 _10246_ (.A(net198),
    .B(_04974_),
    .X(_04986_));
 sg13g2_buf_1 _10247_ (.A(_04986_),
    .X(_04987_));
 sg13g2_and2_1 _10248_ (.A(_01003_),
    .B(net246),
    .X(_04988_));
 sg13g2_buf_1 _10249_ (.A(_04988_),
    .X(_04989_));
 sg13g2_nand2_1 _10250_ (.Y(_04990_),
    .A(net178),
    .B(_04989_));
 sg13g2_nor2_1 _10251_ (.A(net350),
    .B(_04990_),
    .Y(_04991_));
 sg13g2_a22oi_1 _10252_ (.Y(_04992_),
    .B1(_04991_),
    .B2(_02324_),
    .A2(_04987_),
    .A1(net6));
 sg13g2_nor2_1 _10253_ (.A(_02324_),
    .B(_04990_),
    .Y(_04993_));
 sg13g2_o21ai_1 _10254_ (.B1(net350),
    .Y(_04994_),
    .A1(_04970_),
    .A2(_04993_));
 sg13g2_o21ai_1 _10255_ (.B1(_04994_),
    .Y(_04995_),
    .A1(net132),
    .A2(_04992_));
 sg13g2_a22oi_1 _10256_ (.Y(_04996_),
    .B1(_04995_),
    .B2(net227),
    .A2(_04985_),
    .A1(_02297_));
 sg13g2_inv_1 _10257_ (.Y(_00459_),
    .A(_04996_));
 sg13g2_nand3_1 _10258_ (.B(_01289_),
    .C(net241),
    .A(net301),
    .Y(_04997_));
 sg13g2_nor4_1 _10259_ (.A(_02357_),
    .B(_02275_),
    .C(_02365_),
    .D(_04997_),
    .Y(_04998_));
 sg13g2_nand4_1 _10260_ (.B(_02268_),
    .C(_04609_),
    .A(_01057_),
    .Y(_04999_),
    .D(_04998_));
 sg13g2_nand2_1 _10261_ (.Y(_05000_),
    .A(net241),
    .B(_01273_));
 sg13g2_o21ai_1 _10262_ (.B1(_05000_),
    .Y(_05001_),
    .A1(_02261_),
    .A2(_04999_));
 sg13g2_nand2_1 _10263_ (.Y(_05002_),
    .A(net212),
    .B(_05001_));
 sg13g2_buf_2 _10264_ (.A(_05002_),
    .X(_05003_));
 sg13g2_nand2_1 _10265_ (.Y(_05004_),
    .A(_01346_),
    .B(_05003_));
 sg13g2_a21oi_1 _10266_ (.A1(_02443_),
    .A2(_04980_),
    .Y(_05005_),
    .B1(_05004_));
 sg13g2_nand4_1 _10267_ (.B(_04775_),
    .C(_04776_),
    .A(_04771_),
    .Y(_05006_),
    .D(_04989_));
 sg13g2_a21oi_1 _10268_ (.A1(net164),
    .A2(_05003_),
    .Y(_05007_),
    .B1(net225));
 sg13g2_nor2_2 _10269_ (.A(net263),
    .B(_05003_),
    .Y(_05008_));
 sg13g2_nand2b_1 _10270_ (.Y(_05009_),
    .B(_05008_),
    .A_N(net389));
 sg13g2_o21ai_1 _10271_ (.B1(_05009_),
    .Y(_05010_),
    .A1(_02443_),
    .A2(_05007_));
 sg13g2_a21oi_1 _10272_ (.A1(_05005_),
    .A2(_05006_),
    .Y(_00460_),
    .B1(_05010_));
 sg13g2_xnor2_1 _10273_ (.Y(_05011_),
    .A(_04787_),
    .B(_04789_));
 sg13g2_nor2_1 _10274_ (.A(net198),
    .B(_04976_),
    .Y(_05012_));
 sg13g2_nand3_1 _10275_ (.B(_05012_),
    .C(_05003_),
    .A(net264),
    .Y(_05013_));
 sg13g2_buf_1 _10276_ (.A(_05013_),
    .X(_05014_));
 sg13g2_inv_1 _10277_ (.Y(_05015_),
    .A(_05014_));
 sg13g2_nand2_1 _10278_ (.Y(_05016_),
    .A(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .B(_04978_));
 sg13g2_nand4_1 _10279_ (.B(_04976_),
    .C(_05003_),
    .A(net168),
    .Y(_05017_),
    .D(_05016_));
 sg13g2_o21ai_1 _10280_ (.B1(_05017_),
    .Y(_05018_),
    .A1(net388),
    .A2(_05003_));
 sg13g2_nor2_1 _10281_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .B(_05007_),
    .Y(_05019_));
 sg13g2_a221oi_1 _10282_ (.B2(net227),
    .C1(_05019_),
    .B1(_05018_),
    .A1(_05011_),
    .Y(_00461_),
    .A2(_05015_));
 sg13g2_xnor2_1 _10283_ (.Y(_05020_),
    .A(_04796_),
    .B(_04801_));
 sg13g2_o21ai_1 _10284_ (.B1(_05003_),
    .Y(_05021_),
    .A1(net198),
    .A2(_04980_));
 sg13g2_nand2_1 _10285_ (.Y(_05022_),
    .A(net264),
    .B(_05021_));
 sg13g2_buf_2 _10286_ (.A(_05022_),
    .X(_05023_));
 sg13g2_a22oi_1 _10287_ (.Y(_05024_),
    .B1(_05023_),
    .B2(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .A2(_05008_),
    .A1(net387));
 sg13g2_o21ai_1 _10288_ (.B1(_05024_),
    .Y(_00462_),
    .A1(_05020_),
    .A2(_05014_));
 sg13g2_nand3_1 _10289_ (.B(_04814_),
    .C(_05015_),
    .A(_04810_),
    .Y(_05025_));
 sg13g2_a22oi_1 _10290_ (.Y(_05026_),
    .B1(_05023_),
    .B2(_02545_),
    .A2(_05008_),
    .A1(net386));
 sg13g2_nand2_1 _10291_ (.Y(_00463_),
    .A(_05025_),
    .B(_05026_));
 sg13g2_xnor2_1 _10292_ (.Y(_05027_),
    .A(_04835_),
    .B(_04837_));
 sg13g2_a22oi_1 _10293_ (.Y(_05028_),
    .B1(_05023_),
    .B2(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .A2(_05008_),
    .A1(net385));
 sg13g2_o21ai_1 _10294_ (.B1(_05028_),
    .Y(_00464_),
    .A1(_05027_),
    .A2(_05014_));
 sg13g2_nand3b_1 _10295_ (.B(_05015_),
    .C(_04850_),
    .Y(_05029_),
    .A_N(_04855_));
 sg13g2_nand3_1 _10296_ (.B(_04855_),
    .C(_05015_),
    .A(_04847_),
    .Y(_05030_));
 sg13g2_a22oi_1 _10297_ (.Y(_05031_),
    .B1(_05023_),
    .B2(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .A2(_05008_),
    .A1(net349));
 sg13g2_nand3_1 _10298_ (.B(_05030_),
    .C(_05031_),
    .A(_05029_),
    .Y(_00465_));
 sg13g2_nand2_1 _10299_ (.Y(_05032_),
    .A(_04863_),
    .B(_05012_));
 sg13g2_a22oi_1 _10300_ (.Y(_05033_),
    .B1(_04987_),
    .B2(net7),
    .A2(_04983_),
    .A1(_02426_));
 sg13g2_nand2_1 _10301_ (.Y(_05034_),
    .A(_05032_),
    .B(_05033_));
 sg13g2_mux2_1 _10302_ (.A0(_05034_),
    .A1(net390),
    .S(net132),
    .X(_05035_));
 sg13g2_mux2_1 _10303_ (.A0(_02426_),
    .A1(_05035_),
    .S(net211),
    .X(_00466_));
 sg13g2_nand2_1 _10304_ (.Y(_05036_),
    .A(_04875_),
    .B(_05012_));
 sg13g2_a22oi_1 _10305_ (.Y(_05037_),
    .B1(_04987_),
    .B2(net8),
    .A2(_04983_),
    .A1(_02420_));
 sg13g2_nand2_1 _10306_ (.Y(_05038_),
    .A(_05036_),
    .B(_05037_));
 sg13g2_mux2_1 _10307_ (.A0(_05038_),
    .A1(net389),
    .S(net132),
    .X(_05039_));
 sg13g2_nand2_1 _10308_ (.Y(_05040_),
    .A(net211),
    .B(_05039_));
 sg13g2_o21ai_1 _10309_ (.B1(_05040_),
    .Y(_00467_),
    .A1(_02664_),
    .A2(net227));
 sg13g2_nand2_1 _10310_ (.Y(_05041_),
    .A(_02422_),
    .B(_04978_));
 sg13g2_o21ai_1 _10311_ (.B1(_05041_),
    .Y(_05042_),
    .A1(net262),
    .A2(_04978_));
 sg13g2_and2_1 _10312_ (.A(_04976_),
    .B(_05042_),
    .X(_05043_));
 sg13g2_a221oi_1 _10313_ (.B2(_04989_),
    .C1(_05043_),
    .B1(_04884_),
    .A1(net166),
    .Y(_05044_),
    .A2(_01593_));
 sg13g2_mux2_1 _10314_ (.A0(_02422_),
    .A1(net9),
    .S(_04974_),
    .X(_05045_));
 sg13g2_nor2_1 _10315_ (.A(_01951_),
    .B(_05045_),
    .Y(_05046_));
 sg13g2_nor3_1 _10316_ (.A(_04971_),
    .B(_05044_),
    .C(_05046_),
    .Y(_05047_));
 sg13g2_a21oi_1 _10317_ (.A1(net388),
    .A2(_04971_),
    .Y(_05048_),
    .B1(_05047_));
 sg13g2_nand2_1 _10318_ (.Y(_05049_),
    .A(_02422_),
    .B(_04671_));
 sg13g2_o21ai_1 _10319_ (.B1(_05049_),
    .Y(_00468_),
    .A1(net197),
    .A2(_05048_));
 sg13g2_mux2_1 _10320_ (.A0(_02421_),
    .A1(net10),
    .S(_04974_),
    .X(_05050_));
 sg13g2_nor2_1 _10321_ (.A(net261),
    .B(_04978_),
    .Y(_05051_));
 sg13g2_a221oi_1 _10322_ (.B2(_04978_),
    .C1(_05051_),
    .B1(_02421_),
    .A1(_01008_),
    .Y(_05052_),
    .A2(_04549_));
 sg13g2_a221oi_1 _10323_ (.B2(_04989_),
    .C1(_05052_),
    .B1(_04891_),
    .A1(net166),
    .Y(_05053_),
    .A2(_01593_));
 sg13g2_a21oi_1 _10324_ (.A1(_02609_),
    .A2(_05050_),
    .Y(_05054_),
    .B1(_05053_));
 sg13g2_nand2_1 _10325_ (.Y(_05055_),
    .A(net387),
    .B(net132));
 sg13g2_o21ai_1 _10326_ (.B1(_05055_),
    .Y(_05056_),
    .A1(net132),
    .A2(_05054_));
 sg13g2_mux2_1 _10327_ (.A0(_02421_),
    .A1(_05056_),
    .S(_04590_),
    .X(_00469_));
 sg13g2_nand2_1 _10328_ (.Y(_05057_),
    .A(_02419_),
    .B(_04978_));
 sg13g2_o21ai_1 _10329_ (.B1(_05057_),
    .Y(_05058_),
    .A1(net259),
    .A2(_04978_));
 sg13g2_nand2_1 _10330_ (.Y(_05059_),
    .A(_04976_),
    .B(_05058_));
 sg13g2_o21ai_1 _10331_ (.B1(_05059_),
    .Y(_05060_),
    .A1(_04908_),
    .A2(_04976_));
 sg13g2_nand2_1 _10332_ (.Y(_05061_),
    .A(net11),
    .B(_04974_));
 sg13g2_o21ai_1 _10333_ (.B1(_05061_),
    .Y(_05062_),
    .A1(_04492_),
    .A2(_04974_));
 sg13g2_mux2_1 _10334_ (.A0(_05060_),
    .A1(_05062_),
    .S(_01341_),
    .X(_05063_));
 sg13g2_mux2_1 _10335_ (.A0(_05063_),
    .A1(net386),
    .S(net132),
    .X(_05064_));
 sg13g2_mux2_1 _10336_ (.A0(_02419_),
    .A1(_05064_),
    .S(_04590_),
    .X(_00470_));
 sg13g2_xnor2_1 _10337_ (.Y(_05065_),
    .A(_04762_),
    .B(_04918_));
 sg13g2_a22oi_1 _10338_ (.Y(_05066_),
    .B1(_04987_),
    .B2(net12),
    .A2(_04983_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sg13g2_o21ai_1 _10339_ (.B1(_05066_),
    .Y(_05067_),
    .A1(_05065_),
    .A2(_04990_));
 sg13g2_mux2_1 _10340_ (.A0(_05067_),
    .A1(net385),
    .S(_04970_),
    .X(_05068_));
 sg13g2_nand2_1 _10341_ (.Y(_05069_),
    .A(net211),
    .B(_05068_));
 sg13g2_o21ai_1 _10342_ (.B1(_05069_),
    .Y(_00471_),
    .A1(_04504_),
    .A2(net227));
 sg13g2_nor2_1 _10343_ (.A(net349),
    .B(net202),
    .Y(_05070_));
 sg13g2_a221oi_1 _10344_ (.B2(net13),
    .C1(_04970_),
    .B1(_04987_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .Y(_05071_),
    .A2(_04983_));
 sg13g2_nand2_1 _10345_ (.Y(_05072_),
    .A(net264),
    .B(_05071_));
 sg13g2_a21oi_1 _10346_ (.A1(_04926_),
    .A2(_05012_),
    .Y(_05073_),
    .B1(_05072_));
 sg13g2_a221oi_1 _10347_ (.B2(_05070_),
    .C1(_05073_),
    .B1(net132),
    .A1(_02418_),
    .Y(_00472_),
    .A2(net197));
 sg13g2_nor3_1 _10348_ (.A(_01452_),
    .B(net222),
    .C(_05003_),
    .Y(_05074_));
 sg13g2_a21o_1 _10349_ (.A2(_05023_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .B1(_05074_),
    .X(_05075_));
 sg13g2_a21o_1 _10350_ (.A2(_05015_),
    .A1(_04939_),
    .B1(_05075_),
    .X(_00473_));
 sg13g2_nand3_1 _10351_ (.B(_04949_),
    .C(_05015_),
    .A(_04946_),
    .Y(_05076_));
 sg13g2_a22oi_1 _10352_ (.Y(_05077_),
    .B1(_05023_),
    .B2(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .A2(_05008_),
    .A1(net390));
 sg13g2_nand2_1 _10353_ (.Y(_00474_),
    .A(_05076_),
    .B(_05077_));
 sg13g2_nand4_1 _10354_ (.B(net265),
    .C(net203),
    .A(net220),
    .Y(_05078_),
    .D(_00672_));
 sg13g2_inv_1 _10355_ (.Y(_05079_),
    .A(_05078_));
 sg13g2_a221oi_1 _10356_ (.B2(_05079_),
    .C1(net263),
    .B1(_01320_),
    .A1(_00214_),
    .Y(_05080_),
    .A2(net169));
 sg13g2_nand3_1 _10357_ (.B(_01344_),
    .C(_05080_),
    .A(_01312_),
    .Y(_05081_));
 sg13g2_a22oi_1 _10358_ (.Y(_05082_),
    .B1(_05081_),
    .B2(_02313_),
    .A2(_05080_),
    .A1(_02246_));
 sg13g2_inv_1 _10359_ (.Y(_00475_),
    .A(_05082_));
 sg13g2_nor2_1 _10360_ (.A(_01342_),
    .B(_05078_),
    .Y(_05083_));
 sg13g2_nand2_1 _10361_ (.Y(_05084_),
    .A(_01317_),
    .B(_01344_));
 sg13g2_a22oi_1 _10362_ (.Y(_05085_),
    .B1(_05084_),
    .B2(\z80.tv80s.i_tv80_core.XY_State[0] ),
    .A2(_05083_),
    .A1(net339));
 sg13g2_inv_1 _10363_ (.Y(_00476_),
    .A(_05085_));
 sg13g2_a22oi_1 _10364_ (.Y(_05086_),
    .B1(_05084_),
    .B2(_01031_),
    .A2(_05083_),
    .A1(net223));
 sg13g2_inv_1 _10365_ (.Y(_00477_),
    .A(_05086_));
 sg13g2_nand4_1 _10366_ (.B(\z80.tv80s.i_tv80_core.ISet[1] ),
    .C(_02140_),
    .A(net357),
    .Y(_05087_),
    .D(_02231_));
 sg13g2_nand2_1 _10367_ (.Y(_05088_),
    .A(\z80.tv80s.i_tv80_core.Z16_r ),
    .B(_03850_));
 sg13g2_o21ai_1 _10368_ (.B1(_05088_),
    .Y(_00478_),
    .A1(_01615_),
    .A2(_05087_));
 sg13g2_inv_1 _10369_ (.Y(_05089_),
    .A(net22));
 sg13g2_nand2_1 _10370_ (.Y(_05090_),
    .A(_04589_),
    .B(_01533_));
 sg13g2_nor3_1 _10371_ (.A(_01536_),
    .B(_03697_),
    .C(_05090_),
    .Y(_05091_));
 sg13g2_inv_1 _10372_ (.Y(_05092_),
    .A(\z80.tv80s.i_tv80_core.ts[1] ));
 sg13g2_nor2_1 _10373_ (.A(_05092_),
    .B(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ),
    .Y(_05093_));
 sg13g2_buf_1 _10374_ (.A(_05093_),
    .X(_05094_));
 sg13g2_o21ai_1 _10375_ (.B1(_01236_),
    .Y(_05095_),
    .A1(_05091_),
    .A2(_05094_));
 sg13g2_buf_2 _10376_ (.A(_05095_),
    .X(_05096_));
 sg13g2_or3_1 _10377_ (.A(_01536_),
    .B(_03697_),
    .C(_05090_),
    .X(_05097_));
 sg13g2_buf_1 _10378_ (.A(_05097_),
    .X(_05098_));
 sg13g2_buf_1 _10379_ (.A(_05098_),
    .X(_05099_));
 sg13g2_buf_1 _10380_ (.A(_01390_),
    .X(_05100_));
 sg13g2_buf_1 _10381_ (.A(net167),
    .X(_05101_));
 sg13g2_nand2b_1 _10382_ (.Y(_05102_),
    .B(net156),
    .A_N(_01468_));
 sg13g2_o21ai_1 _10383_ (.B1(_05102_),
    .Y(_05103_),
    .A1(net156),
    .A2(net378));
 sg13g2_nand2_1 _10384_ (.Y(_05104_),
    .A(_05100_),
    .B(_05103_));
 sg13g2_o21ai_1 _10385_ (.B1(_05104_),
    .Y(_05105_),
    .A1(net348),
    .A2(net153));
 sg13g2_nand3_1 _10386_ (.B(net287),
    .C(_05105_),
    .A(_05099_),
    .Y(_05106_));
 sg13g2_o21ai_1 _10387_ (.B1(_05106_),
    .Y(_05107_),
    .A1(_03696_),
    .A2(_05099_));
 sg13g2_a22oi_1 _10388_ (.Y(_00479_),
    .B1(_05107_),
    .B2(_04556_),
    .A2(_05096_),
    .A1(_05089_));
 sg13g2_inv_1 _10389_ (.Y(_05108_),
    .A(net23));
 sg13g2_nand2b_1 _10390_ (.Y(_05109_),
    .B(net156),
    .A_N(net342));
 sg13g2_o21ai_1 _10391_ (.B1(_05109_),
    .Y(_05110_),
    .A1(net156),
    .A2(_01876_));
 sg13g2_nand2_1 _10392_ (.Y(_05111_),
    .A(net153),
    .B(_05110_));
 sg13g2_o21ai_1 _10393_ (.B1(_05111_),
    .Y(_05112_),
    .A1(_01636_),
    .A2(net153));
 sg13g2_nand3_1 _10394_ (.B(net287),
    .C(_05112_),
    .A(net157),
    .Y(_05113_));
 sg13g2_o21ai_1 _10395_ (.B1(_05113_),
    .Y(_05114_),
    .A1(_01681_),
    .A2(net157));
 sg13g2_a22oi_1 _10396_ (.Y(_00480_),
    .B1(_05114_),
    .B2(net188),
    .A2(_05096_),
    .A1(_05108_));
 sg13g2_inv_1 _10397_ (.Y(_05115_),
    .A(net24));
 sg13g2_nand2b_1 _10398_ (.Y(_05116_),
    .B(net167),
    .A_N(net341));
 sg13g2_o21ai_1 _10399_ (.B1(_05116_),
    .Y(_05117_),
    .A1(_05101_),
    .A2(net374));
 sg13g2_nand2_1 _10400_ (.Y(_05118_),
    .A(_01390_),
    .B(_05117_));
 sg13g2_o21ai_1 _10401_ (.B1(_05118_),
    .Y(_05119_),
    .A1(net380),
    .A2(net153));
 sg13g2_nand3_1 _10402_ (.B(net287),
    .C(_05119_),
    .A(net157),
    .Y(_05120_));
 sg13g2_o21ai_1 _10403_ (.B1(_05120_),
    .Y(_05121_),
    .A1(_01734_),
    .A2(net157));
 sg13g2_a22oi_1 _10404_ (.Y(_00481_),
    .B1(_05121_),
    .B2(net188),
    .A2(_05096_),
    .A1(_05115_));
 sg13g2_inv_1 _10405_ (.Y(_05122_),
    .A(net25));
 sg13g2_nand2b_1 _10406_ (.Y(_05123_),
    .B(net167),
    .A_N(net340));
 sg13g2_o21ai_1 _10407_ (.B1(_05123_),
    .Y(_05124_),
    .A1(net156),
    .A2(net334));
 sg13g2_nand2_1 _10408_ (.Y(_05125_),
    .A(_01390_),
    .B(_05124_));
 sg13g2_o21ai_1 _10409_ (.B1(_05125_),
    .Y(_05126_),
    .A1(_01757_),
    .A2(net153));
 sg13g2_nand3_1 _10410_ (.B(net287),
    .C(_05126_),
    .A(_05098_),
    .Y(_05127_));
 sg13g2_o21ai_1 _10411_ (.B1(_05127_),
    .Y(_05128_),
    .A1(_01801_),
    .A2(net157));
 sg13g2_a22oi_1 _10412_ (.Y(_00482_),
    .B1(_05128_),
    .B2(net188),
    .A2(_05096_),
    .A1(_05122_));
 sg13g2_inv_1 _10413_ (.Y(_05129_),
    .A(net26));
 sg13g2_nand2b_1 _10414_ (.Y(_05130_),
    .B(net167),
    .A_N(net348));
 sg13g2_o21ai_1 _10415_ (.B1(_05130_),
    .Y(_05131_),
    .A1(net156),
    .A2(_01468_));
 sg13g2_nand2_1 _10416_ (.Y(_05132_),
    .A(_01390_),
    .B(_05131_));
 sg13g2_o21ai_1 _10417_ (.B1(_05132_),
    .Y(_05133_),
    .A1(net378),
    .A2(net153));
 sg13g2_nand3_1 _10418_ (.B(net287),
    .C(_05133_),
    .A(_05098_),
    .Y(_05134_));
 sg13g2_o21ai_1 _10419_ (.B1(_05134_),
    .Y(_05135_),
    .A1(_03877_),
    .A2(net157));
 sg13g2_a22oi_1 _10420_ (.Y(_00483_),
    .B1(_05135_),
    .B2(net188),
    .A2(_05096_),
    .A1(_05129_));
 sg13g2_inv_1 _10421_ (.Y(_05136_),
    .A(net27));
 sg13g2_nand2b_1 _10422_ (.Y(_05137_),
    .B(net167),
    .A_N(_01636_));
 sg13g2_o21ai_1 _10423_ (.B1(_05137_),
    .Y(_05138_),
    .A1(net156),
    .A2(net342));
 sg13g2_nand2_1 _10424_ (.Y(_05139_),
    .A(_01390_),
    .B(_05138_));
 sg13g2_o21ai_1 _10425_ (.B1(_05139_),
    .Y(_05140_),
    .A1(_01876_),
    .A2(net153));
 sg13g2_nand3_1 _10426_ (.B(net287),
    .C(_05140_),
    .A(_05098_),
    .Y(_05141_));
 sg13g2_o21ai_1 _10427_ (.B1(_05141_),
    .Y(_05142_),
    .A1(_01947_),
    .A2(net157));
 sg13g2_a22oi_1 _10428_ (.Y(_00484_),
    .B1(_05142_),
    .B2(net188),
    .A2(_05096_),
    .A1(_05136_));
 sg13g2_inv_1 _10429_ (.Y(_05143_),
    .A(net28));
 sg13g2_nand2b_1 _10430_ (.Y(_05144_),
    .B(net167),
    .A_N(net380));
 sg13g2_o21ai_1 _10431_ (.B1(_05144_),
    .Y(_05145_),
    .A1(_05101_),
    .A2(net341));
 sg13g2_nand2_1 _10432_ (.Y(_05146_),
    .A(_01390_),
    .B(_05145_));
 sg13g2_o21ai_1 _10433_ (.B1(_05146_),
    .Y(_05147_),
    .A1(net374),
    .A2(_05100_));
 sg13g2_nand3_1 _10434_ (.B(net287),
    .C(_05147_),
    .A(_05098_),
    .Y(_05148_));
 sg13g2_o21ai_1 _10435_ (.B1(_05148_),
    .Y(_05149_),
    .A1(_02006_),
    .A2(net157));
 sg13g2_a22oi_1 _10436_ (.Y(_00485_),
    .B1(_05149_),
    .B2(net188),
    .A2(_05096_),
    .A1(_05143_));
 sg13g2_inv_1 _10437_ (.Y(_05150_),
    .A(net29));
 sg13g2_nand2_1 _10438_ (.Y(_05151_),
    .A(_02075_),
    .B(_05091_));
 sg13g2_nand2b_1 _10439_ (.Y(_05152_),
    .B(net167),
    .A_N(_01757_));
 sg13g2_o21ai_1 _10440_ (.B1(_05152_),
    .Y(_05153_),
    .A1(net156),
    .A2(net340));
 sg13g2_nand2_1 _10441_ (.Y(_05154_),
    .A(_01390_),
    .B(_05153_));
 sg13g2_o21ai_1 _10442_ (.B1(_05154_),
    .Y(_05155_),
    .A1(net334),
    .A2(net153));
 sg13g2_nand3_1 _10443_ (.B(net287),
    .C(_05155_),
    .A(_05098_),
    .Y(_05156_));
 sg13g2_a21oi_1 _10444_ (.A1(_05151_),
    .A2(_05156_),
    .Y(_05157_),
    .B1(net189));
 sg13g2_a21oi_1 _10445_ (.A1(_05150_),
    .A2(_05096_),
    .Y(_00486_),
    .B1(_05157_));
 sg13g2_nor2_1 _10446_ (.A(net238),
    .B(_01319_),
    .Y(_05158_));
 sg13g2_a21oi_1 _10447_ (.A1(net238),
    .A2(_03033_),
    .Y(_05159_),
    .B1(_05158_));
 sg13g2_nand2_1 _10448_ (.Y(_05160_),
    .A(_03167_),
    .B(_04178_));
 sg13g2_and4_1 _10449_ (.A(_01418_),
    .B(_01567_),
    .C(_01571_),
    .D(_02362_),
    .X(_05161_));
 sg13g2_buf_1 _10450_ (.A(_05161_),
    .X(_05162_));
 sg13g2_o21ai_1 _10451_ (.B1(_05162_),
    .Y(_05163_),
    .A1(net393),
    .A2(_01540_));
 sg13g2_o21ai_1 _10452_ (.B1(_05163_),
    .Y(_05164_),
    .A1(_05159_),
    .A2(_05160_));
 sg13g2_or3_1 _10453_ (.A(_01530_),
    .B(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .C(_00210_),
    .X(_05165_));
 sg13g2_a21oi_1 _10454_ (.A1(_03697_),
    .A2(_05165_),
    .Y(_05166_),
    .B1(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ));
 sg13g2_a21oi_1 _10455_ (.A1(_04589_),
    .A2(_03698_),
    .Y(_05167_),
    .B1(_04674_));
 sg13g2_o21ai_1 _10456_ (.B1(_01535_),
    .Y(_05168_),
    .A1(_05166_),
    .A2(_05167_));
 sg13g2_nor2_1 _10457_ (.A(_05090_),
    .B(_05168_),
    .Y(_05169_));
 sg13g2_o21ai_1 _10458_ (.B1(_01235_),
    .Y(_05170_),
    .A1(_05164_),
    .A2(_05169_));
 sg13g2_buf_1 _10459_ (.A(_05170_),
    .X(_05171_));
 sg13g2_nor2_1 _10460_ (.A(_03327_),
    .B(_05171_),
    .Y(_05172_));
 sg13g2_nand2_1 _10461_ (.Y(_05173_),
    .A(net79),
    .B(_05172_));
 sg13g2_buf_2 _10462_ (.A(_05173_),
    .X(_05174_));
 sg13g2_nor2_1 _10463_ (.A(_03516_),
    .B(_03529_),
    .Y(_05175_));
 sg13g2_nor2_1 _10464_ (.A(net258),
    .B(_03033_),
    .Y(_05176_));
 sg13g2_a21oi_1 _10465_ (.A1(net258),
    .A2(_00032_),
    .Y(_05177_),
    .B1(_05176_));
 sg13g2_and2_1 _10466_ (.A(_04178_),
    .B(_05177_),
    .X(_05178_));
 sg13g2_buf_1 _10467_ (.A(_05178_),
    .X(_05179_));
 sg13g2_buf_1 _10468_ (.A(_05179_),
    .X(_05180_));
 sg13g2_buf_1 _10469_ (.A(net87),
    .X(_05181_));
 sg13g2_nor2_2 _10470_ (.A(_03140_),
    .B(net144),
    .Y(_05182_));
 sg13g2_nand2b_1 _10471_ (.Y(_05183_),
    .B(_05182_),
    .A_N(\z80.tv80s.i_tv80_core.RegBusA_r[8] ));
 sg13g2_nand2_1 _10472_ (.Y(_05184_),
    .A(net74),
    .B(_05183_));
 sg13g2_nor3_1 _10473_ (.A(_04127_),
    .B(_05175_),
    .C(_05184_),
    .Y(_05185_));
 sg13g2_inv_1 _10474_ (.Y(_05186_),
    .A(_05179_));
 sg13g2_nand3_1 _10475_ (.B(net86),
    .C(_05183_),
    .A(_03696_),
    .Y(_05187_));
 sg13g2_nor2_2 _10476_ (.A(_03102_),
    .B(_03104_),
    .Y(_05188_));
 sg13g2_nand2_1 _10477_ (.Y(_05189_),
    .A(_05188_),
    .B(_05183_));
 sg13g2_a21oi_1 _10478_ (.A1(_05187_),
    .A2(_05189_),
    .Y(_05190_),
    .B1(_05175_));
 sg13g2_nor2_1 _10479_ (.A(_05185_),
    .B(_05190_),
    .Y(_05191_));
 sg13g2_buf_2 _10480_ (.A(_05191_),
    .X(_05192_));
 sg13g2_nand2_1 _10481_ (.Y(_05193_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ),
    .B(_05174_));
 sg13g2_o21ai_1 _10482_ (.B1(_05193_),
    .Y(_00487_),
    .A1(_05174_),
    .A2(_05192_));
 sg13g2_nor3_1 _10483_ (.A(_03327_),
    .B(_03189_),
    .C(_05171_),
    .Y(_05194_));
 sg13g2_buf_2 _10484_ (.A(_05194_),
    .X(_05195_));
 sg13g2_nand2_1 _10485_ (.Y(_05196_),
    .A(_01681_),
    .B(net86));
 sg13g2_inv_1 _10486_ (.Y(_05197_),
    .A(_05196_));
 sg13g2_a221oi_1 _10487_ (.B2(net74),
    .C1(_05197_),
    .B1(_04105_),
    .A1(_05162_),
    .Y(_05198_),
    .A2(_03098_));
 sg13g2_buf_1 _10488_ (.A(net144),
    .X(_05199_));
 sg13g2_buf_1 _10489_ (.A(_03140_),
    .X(_05200_));
 sg13g2_nor3_1 _10490_ (.A(\z80.tv80s.i_tv80_core.RegBusA_r[9] ),
    .B(net140),
    .C(net144),
    .Y(_05201_));
 sg13g2_a21oi_1 _10491_ (.A1(net131),
    .A2(_03547_),
    .Y(_05202_),
    .B1(_05201_));
 sg13g2_nand2b_1 _10492_ (.Y(_05203_),
    .B(_05202_),
    .A_N(_05198_));
 sg13g2_buf_2 _10493_ (.A(_05203_),
    .X(_05204_));
 sg13g2_nor2_1 _10494_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ),
    .B(_05195_),
    .Y(_05205_));
 sg13g2_a21oi_1 _10495_ (.A1(_05195_),
    .A2(_05204_),
    .Y(_00488_),
    .B1(_05205_));
 sg13g2_inv_1 _10496_ (.Y(_05206_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[10] ));
 sg13g2_nand2_1 _10497_ (.Y(_05207_),
    .A(net151),
    .B(_03099_));
 sg13g2_nand2_1 _10498_ (.Y(_05208_),
    .A(_01734_),
    .B(_05186_));
 sg13g2_nand2_1 _10499_ (.Y(_05209_),
    .A(_05207_),
    .B(_05208_));
 sg13g2_a21oi_1 _10500_ (.A1(_04156_),
    .A2(net74),
    .Y(_05210_),
    .B1(_05209_));
 sg13g2_a221oi_1 _10501_ (.B2(_05206_),
    .C1(_05210_),
    .B1(_05182_),
    .A1(net131),
    .Y(_05211_),
    .A2(_03577_));
 sg13g2_buf_2 _10502_ (.A(_05211_),
    .X(_05212_));
 sg13g2_mux2_1 _10503_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ),
    .A1(_05212_),
    .S(_05195_),
    .X(_00489_));
 sg13g2_mux2_1 _10504_ (.A0(_00060_),
    .A1(_00056_),
    .S(_02850_),
    .X(_05213_));
 sg13g2_nor2_1 _10505_ (.A(_01801_),
    .B(_05180_),
    .Y(_05214_));
 sg13g2_a21o_1 _10506_ (.A2(_05181_),
    .A1(_04060_),
    .B1(_05214_),
    .X(_05215_));
 sg13g2_nor3_1 _10507_ (.A(\z80.tv80s.i_tv80_core.RegBusA_r[11] ),
    .B(net140),
    .C(net131),
    .Y(_05216_));
 sg13g2_a221oi_1 _10508_ (.B2(_05207_),
    .C1(_05216_),
    .B1(_05215_),
    .A1(net131),
    .Y(_05217_),
    .A2(_05213_));
 sg13g2_buf_2 _10509_ (.A(_05217_),
    .X(_05218_));
 sg13g2_mux2_1 _10510_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ),
    .A1(_05218_),
    .S(_05195_),
    .X(_00490_));
 sg13g2_nand2b_1 _10511_ (.Y(_05219_),
    .B(net86),
    .A_N(_01863_));
 sg13g2_nand2_1 _10512_ (.Y(_05220_),
    .A(_05207_),
    .B(_05219_));
 sg13g2_inv_1 _10513_ (.Y(_05221_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[12] ));
 sg13g2_mux2_1 _10514_ (.A0(_00068_),
    .A1(_00064_),
    .S(_02850_),
    .X(_05222_));
 sg13g2_a22oi_1 _10515_ (.Y(_05223_),
    .B1(_05222_),
    .B2(net144),
    .A2(_05182_),
    .A1(_05221_));
 sg13g2_and2_1 _10516_ (.A(net74),
    .B(_05223_),
    .X(_05224_));
 sg13g2_a22oi_1 _10517_ (.Y(_05225_),
    .B1(_05224_),
    .B2(_04143_),
    .A2(_05223_),
    .A1(_05220_));
 sg13g2_buf_2 _10518_ (.A(_05225_),
    .X(_05226_));
 sg13g2_nand2_1 _10519_ (.Y(_05227_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ),
    .B(_05174_));
 sg13g2_o21ai_1 _10520_ (.B1(_05227_),
    .Y(_00491_),
    .A1(_05174_),
    .A2(_05226_));
 sg13g2_inv_1 _10521_ (.Y(_05228_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ));
 sg13g2_nand2_1 _10522_ (.Y(_05229_),
    .A(_03140_),
    .B(net87));
 sg13g2_nand2b_1 _10523_ (.Y(_05230_),
    .B(net41),
    .A_N(_05229_));
 sg13g2_a21oi_1 _10524_ (.A1(_01943_),
    .A2(_01946_),
    .Y(_05231_),
    .B1(_05180_));
 sg13g2_nand2_1 _10525_ (.Y(_05232_),
    .A(net140),
    .B(_05231_));
 sg13g2_o21ai_1 _10526_ (.B1(_05232_),
    .Y(_05233_),
    .A1(_04135_),
    .A2(_05230_));
 sg13g2_nor2_1 _10527_ (.A(net41),
    .B(_05229_),
    .Y(_05234_));
 sg13g2_and2_1 _10528_ (.A(net151),
    .B(_03040_),
    .X(_05235_));
 sg13g2_buf_1 _10529_ (.A(_05235_),
    .X(_05236_));
 sg13g2_and2_1 _10530_ (.A(\z80.tv80s.i_tv80_core.RegBusA_r[13] ),
    .B(net148),
    .X(_05237_));
 sg13g2_a21o_1 _10531_ (.A2(_05234_),
    .A1(_04135_),
    .B1(_05237_),
    .X(_05238_));
 sg13g2_buf_1 _10532_ (.A(net135),
    .X(_05239_));
 sg13g2_o21ai_1 _10533_ (.B1(net116),
    .Y(_05240_),
    .A1(_05233_),
    .A2(_05238_));
 sg13g2_buf_2 _10534_ (.A(_05240_),
    .X(_05241_));
 sg13g2_nor2_2 _10535_ (.A(net116),
    .B(_03635_),
    .Y(_05242_));
 sg13g2_nor2_1 _10536_ (.A(_05174_),
    .B(_05242_),
    .Y(_05243_));
 sg13g2_a22oi_1 _10537_ (.Y(_00492_),
    .B1(_05241_),
    .B2(_05243_),
    .A2(_05174_),
    .A1(_05228_));
 sg13g2_inv_1 _10538_ (.Y(_05244_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ));
 sg13g2_or2_1 _10539_ (.X(_05245_),
    .B(_05229_),
    .A(_03352_));
 sg13g2_nand2b_1 _10540_ (.Y(_05246_),
    .B(_03352_),
    .A_N(_05229_));
 sg13g2_mux2_1 _10541_ (.A0(_05245_),
    .A1(_05246_),
    .S(_04119_),
    .X(_05247_));
 sg13g2_nor2_1 _10542_ (.A(net148),
    .B(net74),
    .Y(_05248_));
 sg13g2_a22oi_1 _10543_ (.Y(_05249_),
    .B1(_05248_),
    .B2(_02006_),
    .A2(net148),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[14] ));
 sg13g2_a21o_1 _10544_ (.A2(_05249_),
    .A1(_05247_),
    .B1(net131),
    .X(_05250_));
 sg13g2_buf_2 _10545_ (.A(_05250_),
    .X(_05251_));
 sg13g2_nor2_2 _10546_ (.A(net116),
    .B(_03654_),
    .Y(_05252_));
 sg13g2_nor2_1 _10547_ (.A(_05174_),
    .B(_05252_),
    .Y(_05253_));
 sg13g2_a22oi_1 _10548_ (.Y(_00493_),
    .B1(_05251_),
    .B2(_05253_),
    .A2(_05174_),
    .A1(_05244_));
 sg13g2_inv_1 _10549_ (.Y(_05254_),
    .A(_03671_));
 sg13g2_and2_1 _10550_ (.A(_04070_),
    .B(_04071_),
    .X(_05255_));
 sg13g2_nor2_1 _10551_ (.A(_05188_),
    .B(net86),
    .Y(_05256_));
 sg13g2_nor3_1 _10552_ (.A(_02075_),
    .B(_05188_),
    .C(net87),
    .Y(_05257_));
 sg13g2_a21o_1 _10553_ (.A2(_05182_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[15] ),
    .B1(_05257_),
    .X(_05258_));
 sg13g2_a221oi_1 _10554_ (.B2(_05256_),
    .C1(_05258_),
    .B1(_05255_),
    .A1(net131),
    .Y(_05259_),
    .A2(_05254_));
 sg13g2_buf_2 _10555_ (.A(_05259_),
    .X(_05260_));
 sg13g2_nor2_1 _10556_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ),
    .B(_05195_),
    .Y(_05261_));
 sg13g2_a21oi_1 _10557_ (.A1(_05195_),
    .A2(_05260_),
    .Y(_00494_),
    .B1(_05261_));
 sg13g2_nor2_1 _10558_ (.A(_03696_),
    .B(net87),
    .Y(_05262_));
 sg13g2_a21oi_1 _10559_ (.A1(_04127_),
    .A2(net74),
    .Y(_05263_),
    .B1(_05262_));
 sg13g2_o21ai_1 _10560_ (.B1(_05183_),
    .Y(_05264_),
    .A1(_05188_),
    .A2(_05263_));
 sg13g2_nand2_1 _10561_ (.Y(_05265_),
    .A(net62),
    .B(_05172_));
 sg13g2_buf_1 _10562_ (.A(_05265_),
    .X(_05266_));
 sg13g2_nand2_1 _10563_ (.Y(_05267_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ),
    .B(net51));
 sg13g2_o21ai_1 _10564_ (.B1(_05267_),
    .Y(_00495_),
    .A1(_05264_),
    .A2(_05266_));
 sg13g2_a21oi_1 _10565_ (.A1(_04105_),
    .A2(_05181_),
    .Y(_05268_),
    .B1(_05197_));
 sg13g2_nor2_1 _10566_ (.A(\z80.tv80s.i_tv80_core.RegBusA_r[9] ),
    .B(net140),
    .Y(_05269_));
 sg13g2_a221oi_1 _10567_ (.B2(_05268_),
    .C1(_05269_),
    .B1(net140),
    .A1(_03033_),
    .Y(_05270_),
    .A2(_05162_));
 sg13g2_mux2_1 _10568_ (.A0(_05270_),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ),
    .S(_05266_),
    .X(_00496_));
 sg13g2_mux2_1 _10569_ (.A0(_05212_),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ),
    .S(net51),
    .X(_00497_));
 sg13g2_mux2_1 _10570_ (.A0(_05218_),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ),
    .S(net51),
    .X(_00498_));
 sg13g2_nand2_1 _10571_ (.Y(_05271_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ),
    .B(net51));
 sg13g2_o21ai_1 _10572_ (.B1(_05271_),
    .Y(_00499_),
    .A1(_05226_),
    .A2(net51));
 sg13g2_nand2_1 _10573_ (.Y(_05272_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ),
    .B(_05265_));
 sg13g2_o21ai_1 _10574_ (.B1(_05272_),
    .Y(_00500_),
    .A1(_05241_),
    .A2(net51));
 sg13g2_nand2_1 _10575_ (.Y(_05273_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ),
    .B(_05265_));
 sg13g2_o21ai_1 _10576_ (.B1(_05273_),
    .Y(_00501_),
    .A1(_05251_),
    .A2(net51));
 sg13g2_a21oi_1 _10577_ (.A1(_05255_),
    .A2(_05256_),
    .Y(_05274_),
    .B1(_05258_));
 sg13g2_nand2_1 _10578_ (.Y(_05275_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ),
    .B(_05265_));
 sg13g2_o21ai_1 _10579_ (.B1(_05275_),
    .Y(_00502_),
    .A1(_05274_),
    .A2(net51));
 sg13g2_nand2_1 _10580_ (.Y(_05276_),
    .A(_03239_),
    .B(_05172_));
 sg13g2_buf_1 _10581_ (.A(_05276_),
    .X(_05277_));
 sg13g2_buf_1 _10582_ (.A(_05277_),
    .X(_05278_));
 sg13g2_nand2_1 _10583_ (.Y(_05279_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .B(net39));
 sg13g2_o21ai_1 _10584_ (.B1(_05279_),
    .Y(_00503_),
    .A1(_05192_),
    .A2(net39));
 sg13g2_nand2_1 _10585_ (.Y(_05280_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .B(net39));
 sg13g2_o21ai_1 _10586_ (.B1(_05280_),
    .Y(_00504_),
    .A1(_05204_),
    .A2(net39));
 sg13g2_mux2_1 _10587_ (.A0(_05212_),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .S(_05278_),
    .X(_00505_));
 sg13g2_mux2_1 _10588_ (.A0(_05218_),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .S(_05278_),
    .X(_00506_));
 sg13g2_nand2_1 _10589_ (.Y(_05281_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .B(_05277_));
 sg13g2_o21ai_1 _10590_ (.B1(_05281_),
    .Y(_00507_),
    .A1(_05226_),
    .A2(net39));
 sg13g2_inv_1 _10591_ (.Y(_05282_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ));
 sg13g2_nor2_1 _10592_ (.A(_05242_),
    .B(_05277_),
    .Y(_05283_));
 sg13g2_a22oi_1 _10593_ (.Y(_00508_),
    .B1(_05283_),
    .B2(_05241_),
    .A2(net39),
    .A1(_05282_));
 sg13g2_inv_1 _10594_ (.Y(_05284_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ));
 sg13g2_nor2_1 _10595_ (.A(_05252_),
    .B(_05277_),
    .Y(_05285_));
 sg13g2_a22oi_1 _10596_ (.Y(_00509_),
    .B1(_05285_),
    .B2(_05251_),
    .A2(net39),
    .A1(_05284_));
 sg13g2_nand2_1 _10597_ (.Y(_05286_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ),
    .B(_05277_));
 sg13g2_o21ai_1 _10598_ (.B1(_05286_),
    .Y(_00510_),
    .A1(_05260_),
    .A2(net39));
 sg13g2_nand2_1 _10599_ (.Y(_05287_),
    .A(net80),
    .B(_05172_));
 sg13g2_buf_1 _10600_ (.A(_05287_),
    .X(_05288_));
 sg13g2_buf_1 _10601_ (.A(_05288_),
    .X(_05289_));
 sg13g2_nand2_1 _10602_ (.Y(_05290_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .B(net38));
 sg13g2_o21ai_1 _10603_ (.B1(_05290_),
    .Y(_00511_),
    .A1(_05192_),
    .A2(net38));
 sg13g2_nand2_1 _10604_ (.Y(_05291_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .B(net38));
 sg13g2_o21ai_1 _10605_ (.B1(_05291_),
    .Y(_00512_),
    .A1(_05204_),
    .A2(_05289_));
 sg13g2_mux2_1 _10606_ (.A0(_05212_),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .S(_05289_),
    .X(_00513_));
 sg13g2_mux2_1 _10607_ (.A0(_05218_),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .S(net38),
    .X(_00514_));
 sg13g2_nand2_1 _10608_ (.Y(_05292_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ),
    .B(_05288_));
 sg13g2_o21ai_1 _10609_ (.B1(_05292_),
    .Y(_00515_),
    .A1(_05226_),
    .A2(net38));
 sg13g2_inv_1 _10610_ (.Y(_05293_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ));
 sg13g2_nor2_1 _10611_ (.A(_05242_),
    .B(_05288_),
    .Y(_05294_));
 sg13g2_a22oi_1 _10612_ (.Y(_00516_),
    .B1(_05294_),
    .B2(_05241_),
    .A2(net38),
    .A1(_05293_));
 sg13g2_inv_1 _10613_ (.Y(_05295_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ));
 sg13g2_nor2_1 _10614_ (.A(_05252_),
    .B(_05288_),
    .Y(_05296_));
 sg13g2_a22oi_1 _10615_ (.Y(_00517_),
    .B1(_05296_),
    .B2(_05251_),
    .A2(net38),
    .A1(_05295_));
 sg13g2_nand2_1 _10616_ (.Y(_05297_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ),
    .B(_05288_));
 sg13g2_o21ai_1 _10617_ (.B1(_05297_),
    .Y(_00518_),
    .A1(_05260_),
    .A2(net38));
 sg13g2_nor2_1 _10618_ (.A(net64),
    .B(_05171_),
    .Y(_05298_));
 sg13g2_nand2_1 _10619_ (.Y(_05299_),
    .A(net79),
    .B(_05298_));
 sg13g2_buf_1 _10620_ (.A(_05299_),
    .X(_05300_));
 sg13g2_buf_1 _10621_ (.A(_05300_),
    .X(_05301_));
 sg13g2_nand2_1 _10622_ (.Y(_05302_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ),
    .B(net50));
 sg13g2_o21ai_1 _10623_ (.B1(_05302_),
    .Y(_00519_),
    .A1(_05192_),
    .A2(net50));
 sg13g2_nand2_1 _10624_ (.Y(_05303_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ),
    .B(net50));
 sg13g2_o21ai_1 _10625_ (.B1(_05303_),
    .Y(_00520_),
    .A1(_05204_),
    .A2(_05301_));
 sg13g2_mux2_1 _10626_ (.A0(_05212_),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ),
    .S(net50),
    .X(_00521_));
 sg13g2_mux2_1 _10627_ (.A0(_05218_),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ),
    .S(_05301_),
    .X(_00522_));
 sg13g2_nand2_1 _10628_ (.Y(_05304_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ),
    .B(_05300_));
 sg13g2_o21ai_1 _10629_ (.B1(_05304_),
    .Y(_00523_),
    .A1(_05226_),
    .A2(net50));
 sg13g2_inv_1 _10630_ (.Y(_05305_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ));
 sg13g2_nor2_1 _10631_ (.A(_05242_),
    .B(_05300_),
    .Y(_05306_));
 sg13g2_a22oi_1 _10632_ (.Y(_00524_),
    .B1(_05306_),
    .B2(_05241_),
    .A2(net50),
    .A1(_05305_));
 sg13g2_inv_1 _10633_ (.Y(_05307_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ));
 sg13g2_nor2_1 _10634_ (.A(_05252_),
    .B(_05300_),
    .Y(_05308_));
 sg13g2_a22oi_1 _10635_ (.Y(_00525_),
    .B1(_05308_),
    .B2(_05251_),
    .A2(net50),
    .A1(_05307_));
 sg13g2_nand2_1 _10636_ (.Y(_05309_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ),
    .B(_05300_));
 sg13g2_o21ai_1 _10637_ (.B1(_05309_),
    .Y(_00526_),
    .A1(_05260_),
    .A2(net50));
 sg13g2_nand2_1 _10638_ (.Y(_05310_),
    .A(net62),
    .B(_05298_));
 sg13g2_buf_1 _10639_ (.A(_05310_),
    .X(_05311_));
 sg13g2_nand2_1 _10640_ (.Y(_05312_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ),
    .B(net53));
 sg13g2_o21ai_1 _10641_ (.B1(_05312_),
    .Y(_00527_),
    .A1(_05264_),
    .A2(net53));
 sg13g2_mux2_1 _10642_ (.A0(_05270_),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ),
    .S(net53),
    .X(_00528_));
 sg13g2_mux2_1 _10643_ (.A0(_05212_),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ),
    .S(net53),
    .X(_00529_));
 sg13g2_mux2_1 _10644_ (.A0(_05218_),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ),
    .S(net53),
    .X(_00530_));
 sg13g2_nand2_1 _10645_ (.Y(_05313_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ),
    .B(net53));
 sg13g2_o21ai_1 _10646_ (.B1(_05313_),
    .Y(_00531_),
    .A1(_05226_),
    .A2(_05311_));
 sg13g2_nand2_1 _10647_ (.Y(_05314_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ),
    .B(_05310_));
 sg13g2_o21ai_1 _10648_ (.B1(_05314_),
    .Y(_00532_),
    .A1(_05241_),
    .A2(net53));
 sg13g2_nand2_1 _10649_ (.Y(_05315_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ),
    .B(_05310_));
 sg13g2_o21ai_1 _10650_ (.B1(_05315_),
    .Y(_00533_),
    .A1(_05251_),
    .A2(net53));
 sg13g2_nand2_1 _10651_ (.Y(_05316_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ),
    .B(_05310_));
 sg13g2_o21ai_1 _10652_ (.B1(_05316_),
    .Y(_00534_),
    .A1(_05274_),
    .A2(_05311_));
 sg13g2_nand2_1 _10653_ (.Y(_05317_),
    .A(_03239_),
    .B(_05298_));
 sg13g2_buf_2 _10654_ (.A(_05317_),
    .X(_05318_));
 sg13g2_nand2_1 _10655_ (.Y(_05319_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .B(_05318_));
 sg13g2_o21ai_1 _10656_ (.B1(_05319_),
    .Y(_00535_),
    .A1(_05192_),
    .A2(_05318_));
 sg13g2_nand2_1 _10657_ (.Y(_05320_),
    .A(net67),
    .B(net60));
 sg13g2_nor3_1 _10658_ (.A(net64),
    .B(_05320_),
    .C(_05171_),
    .Y(_05321_));
 sg13g2_buf_2 _10659_ (.A(_05321_),
    .X(_05322_));
 sg13g2_nor2_1 _10660_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .B(_05322_),
    .Y(_05323_));
 sg13g2_a21oi_1 _10661_ (.A1(_05204_),
    .A2(_05322_),
    .Y(_00536_),
    .B1(_05323_));
 sg13g2_mux2_1 _10662_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .A1(_05212_),
    .S(_05322_),
    .X(_00537_));
 sg13g2_mux2_1 _10663_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .A1(_05218_),
    .S(_05322_),
    .X(_00538_));
 sg13g2_nand2_1 _10664_ (.Y(_05324_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .B(_05318_));
 sg13g2_o21ai_1 _10665_ (.B1(_05324_),
    .Y(_00539_),
    .A1(_05226_),
    .A2(_05318_));
 sg13g2_inv_1 _10666_ (.Y(_05325_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ));
 sg13g2_nor2_1 _10667_ (.A(_05242_),
    .B(_05318_),
    .Y(_05326_));
 sg13g2_a22oi_1 _10668_ (.Y(_00540_),
    .B1(_05326_),
    .B2(_05241_),
    .A2(_05318_),
    .A1(_05325_));
 sg13g2_inv_1 _10669_ (.Y(_05327_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ));
 sg13g2_nor2_1 _10670_ (.A(_05252_),
    .B(_05318_),
    .Y(_05328_));
 sg13g2_a22oi_1 _10671_ (.Y(_00541_),
    .B1(_05328_),
    .B2(_05251_),
    .A2(_05318_),
    .A1(_05327_));
 sg13g2_nor2_1 _10672_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ),
    .B(_05322_),
    .Y(_05329_));
 sg13g2_a21oi_1 _10673_ (.A1(_05260_),
    .A2(_05322_),
    .Y(_00542_),
    .B1(_05329_));
 sg13g2_nand2_1 _10674_ (.Y(_05330_),
    .A(_03161_),
    .B(_03170_));
 sg13g2_or3_1 _10675_ (.A(net64),
    .B(_05330_),
    .C(_05171_),
    .X(_05331_));
 sg13g2_buf_2 _10676_ (.A(_05331_),
    .X(_05332_));
 sg13g2_nand2_1 _10677_ (.Y(_05333_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .B(_05332_));
 sg13g2_o21ai_1 _10678_ (.B1(_05333_),
    .Y(_00543_),
    .A1(_05192_),
    .A2(_05332_));
 sg13g2_nor3_1 _10679_ (.A(net64),
    .B(_05330_),
    .C(_05171_),
    .Y(_05334_));
 sg13g2_buf_2 _10680_ (.A(_05334_),
    .X(_05335_));
 sg13g2_nor2_1 _10681_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .B(_05335_),
    .Y(_05336_));
 sg13g2_a21oi_1 _10682_ (.A1(_05204_),
    .A2(_05335_),
    .Y(_00544_),
    .B1(_05336_));
 sg13g2_mux2_1 _10683_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .A1(_05212_),
    .S(_05335_),
    .X(_00545_));
 sg13g2_mux2_1 _10684_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ),
    .A1(_05218_),
    .S(_05335_),
    .X(_00546_));
 sg13g2_nand2_1 _10685_ (.Y(_05337_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ),
    .B(_05332_));
 sg13g2_o21ai_1 _10686_ (.B1(_05337_),
    .Y(_00547_),
    .A1(_05226_),
    .A2(_05332_));
 sg13g2_inv_1 _10687_ (.Y(_05338_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ));
 sg13g2_nor2_1 _10688_ (.A(_05242_),
    .B(_05332_),
    .Y(_05339_));
 sg13g2_a22oi_1 _10689_ (.Y(_00548_),
    .B1(_05339_),
    .B2(_05241_),
    .A2(_05332_),
    .A1(_05338_));
 sg13g2_inv_1 _10690_ (.Y(_05340_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ));
 sg13g2_nor2_1 _10691_ (.A(_05252_),
    .B(_05332_),
    .Y(_05341_));
 sg13g2_a22oi_1 _10692_ (.Y(_00549_),
    .B1(_05341_),
    .B2(_05251_),
    .A2(_05332_),
    .A1(_05340_));
 sg13g2_nor2_1 _10693_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ),
    .B(_05335_),
    .Y(_05342_));
 sg13g2_a21oi_1 _10694_ (.A1(_05260_),
    .A2(_05335_),
    .Y(_00550_),
    .B1(_05342_));
 sg13g2_a21oi_1 _10695_ (.A1(_04161_),
    .A2(net87),
    .Y(_05343_),
    .B1(_05262_));
 sg13g2_or2_1 _10696_ (.X(_05344_),
    .B(_05343_),
    .A(net148));
 sg13g2_o21ai_1 _10697_ (.B1(_05344_),
    .Y(_05345_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[0] ),
    .A2(_05200_));
 sg13g2_nand2_1 _10698_ (.Y(_05346_),
    .A(net131),
    .B(_03536_));
 sg13g2_o21ai_1 _10699_ (.B1(_05346_),
    .Y(_05347_),
    .A1(net131),
    .A2(_05345_));
 sg13g2_buf_2 _10700_ (.A(_05347_),
    .X(_05348_));
 sg13g2_nor2_1 _10701_ (.A(_01534_),
    .B(_05168_),
    .Y(_05349_));
 sg13g2_o21ai_1 _10702_ (.B1(_01235_),
    .Y(_05350_),
    .A1(_05164_),
    .A2(_05349_));
 sg13g2_nand2b_1 _10703_ (.Y(_05351_),
    .B(net64),
    .A_N(_05350_));
 sg13g2_buf_1 _10704_ (.A(_05351_),
    .X(_05352_));
 sg13g2_nor2_1 _10705_ (.A(_03189_),
    .B(_05352_),
    .Y(_05353_));
 sg13g2_buf_1 _10706_ (.A(_05353_),
    .X(_05354_));
 sg13g2_mux2_1 _10707_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ),
    .A1(_05348_),
    .S(net49),
    .X(_00551_));
 sg13g2_xnor2_1 _10708_ (.Y(_05355_),
    .A(_03212_),
    .B(net117));
 sg13g2_xnor2_1 _10709_ (.Y(_05356_),
    .A(_04161_),
    .B(_05355_));
 sg13g2_a21oi_1 _10710_ (.A1(net87),
    .A2(_05356_),
    .Y(_05357_),
    .B1(_05197_));
 sg13g2_nand2_1 _10711_ (.Y(_05358_),
    .A(\z80.tv80s.i_tv80_core.RegBusA_r[1] ),
    .B(net148));
 sg13g2_o21ai_1 _10712_ (.B1(_05358_),
    .Y(_05359_),
    .A1(net148),
    .A2(_05357_));
 sg13g2_nand2_1 _10713_ (.Y(_05360_),
    .A(net116),
    .B(_05359_));
 sg13g2_o21ai_1 _10714_ (.B1(_05360_),
    .Y(_05361_),
    .A1(net116),
    .A2(_03553_));
 sg13g2_buf_2 _10715_ (.A(_05361_),
    .X(_05362_));
 sg13g2_mux2_1 _10716_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ),
    .A1(_05362_),
    .S(net49),
    .X(_00552_));
 sg13g2_nor3_1 _10717_ (.A(_03125_),
    .B(_03173_),
    .C(_04005_),
    .Y(_05363_));
 sg13g2_nand2_1 _10718_ (.Y(_05364_),
    .A(_03092_),
    .B(_04002_));
 sg13g2_nand2_1 _10719_ (.Y(_05365_),
    .A(_03124_),
    .B(_04003_));
 sg13g2_a221oi_1 _10720_ (.B2(_05365_),
    .C1(net141),
    .B1(_05364_),
    .A1(_04036_),
    .Y(_05366_),
    .A2(_04038_));
 sg13g2_a21oi_1 _10721_ (.A1(net141),
    .A2(_05363_),
    .Y(_05367_),
    .B1(_05366_));
 sg13g2_xnor2_1 _10722_ (.Y(_05368_),
    .A(_03238_),
    .B(_05367_));
 sg13g2_o21ai_1 _10723_ (.B1(_05208_),
    .Y(_05369_),
    .A1(net86),
    .A2(_05368_));
 sg13g2_mux2_1 _10724_ (.A0(\z80.tv80s.i_tv80_core.RegBusA_r[2] ),
    .A1(_05369_),
    .S(_05200_),
    .X(_05370_));
 sg13g2_nor2_1 _10725_ (.A(net116),
    .B(_03581_),
    .Y(_05371_));
 sg13g2_a21o_1 _10726_ (.A2(_05370_),
    .A1(net116),
    .B1(_05371_),
    .X(_05372_));
 sg13g2_buf_2 _10727_ (.A(_05372_),
    .X(_05373_));
 sg13g2_mux2_1 _10728_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .A1(_05373_),
    .S(_05354_),
    .X(_00553_));
 sg13g2_inv_1 _10729_ (.Y(_05374_),
    .A(_05354_));
 sg13g2_nand2_1 _10730_ (.Y(_05375_),
    .A(_04160_),
    .B(_04042_));
 sg13g2_xor2_1 _10731_ (.B(_05375_),
    .A(_04102_),
    .X(_05376_));
 sg13g2_a221oi_1 _10732_ (.B2(_05376_),
    .C1(_05214_),
    .B1(net87),
    .A1(net393),
    .Y(_05377_),
    .A2(_05162_));
 sg13g2_buf_1 _10733_ (.A(_05377_),
    .X(_05378_));
 sg13g2_a21o_1 _10734_ (.A2(_05236_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[3] ),
    .B1(_03038_),
    .X(_05379_));
 sg13g2_buf_1 _10735_ (.A(_05379_),
    .X(_05380_));
 sg13g2_nand2_1 _10736_ (.Y(_05381_),
    .A(_05199_),
    .B(_03609_));
 sg13g2_o21ai_1 _10737_ (.B1(_05381_),
    .Y(_05382_),
    .A1(_05378_),
    .A2(_05380_));
 sg13g2_buf_2 _10738_ (.A(_05382_),
    .X(_05383_));
 sg13g2_nand2_1 _10739_ (.Y(_05384_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ),
    .B(_05374_));
 sg13g2_o21ai_1 _10740_ (.B1(_05384_),
    .Y(_00554_),
    .A1(_05374_),
    .A2(_05383_));
 sg13g2_inv_1 _10741_ (.Y(_05385_),
    .A(_05219_));
 sg13g2_nor3_1 _10742_ (.A(_04172_),
    .B(_04173_),
    .C(net86),
    .Y(_05386_));
 sg13g2_or3_1 _10743_ (.A(net148),
    .B(_05385_),
    .C(_05386_),
    .X(_05387_));
 sg13g2_o21ai_1 _10744_ (.B1(net135),
    .Y(_05388_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[4] ),
    .A2(net140));
 sg13g2_inv_1 _10745_ (.Y(_05389_),
    .A(_05388_));
 sg13g2_nor2_1 _10746_ (.A(_05239_),
    .B(_03621_),
    .Y(_05390_));
 sg13g2_a21oi_1 _10747_ (.A1(_05387_),
    .A2(_05389_),
    .Y(_05391_),
    .B1(_05390_));
 sg13g2_buf_2 _10748_ (.A(_05391_),
    .X(_05392_));
 sg13g2_nor2_1 _10749_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ),
    .B(net49),
    .Y(_05393_));
 sg13g2_a21oi_1 _10750_ (.A1(net49),
    .A2(_05392_),
    .Y(_00555_),
    .B1(_05393_));
 sg13g2_a221oi_1 _10751_ (.B2(net87),
    .C1(_05231_),
    .B1(_04045_),
    .A1(net393),
    .Y(_05394_),
    .A2(_05162_));
 sg13g2_o21ai_1 _10752_ (.B1(_05239_),
    .Y(_05395_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[5] ),
    .A2(net140));
 sg13g2_nand2b_1 _10753_ (.Y(_05396_),
    .B(_05199_),
    .A_N(_03639_));
 sg13g2_o21ai_1 _10754_ (.B1(_05396_),
    .Y(_05397_),
    .A1(_05394_),
    .A2(_05395_));
 sg13g2_buf_2 _10755_ (.A(_05397_),
    .X(_05398_));
 sg13g2_mux2_1 _10756_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ),
    .A1(_05398_),
    .S(net49),
    .X(_00556_));
 sg13g2_xnor2_1 _10757_ (.Y(_05399_),
    .A(_03346_),
    .B(_04147_));
 sg13g2_a21oi_1 _10758_ (.A1(_02006_),
    .A2(net86),
    .Y(_05400_),
    .B1(net148));
 sg13g2_o21ai_1 _10759_ (.B1(_05400_),
    .Y(_05401_),
    .A1(_05399_),
    .A2(net86));
 sg13g2_o21ai_1 _10760_ (.B1(_03516_),
    .Y(_05402_),
    .A1(\z80.tv80s.i_tv80_core.RegBusA_r[6] ),
    .A2(net140));
 sg13g2_inv_1 _10761_ (.Y(_05403_),
    .A(_05402_));
 sg13g2_nor2_1 _10762_ (.A(net116),
    .B(_03658_),
    .Y(_05404_));
 sg13g2_a21oi_1 _10763_ (.A1(_05401_),
    .A2(_05403_),
    .Y(_05405_),
    .B1(_05404_));
 sg13g2_buf_2 _10764_ (.A(_05405_),
    .X(_05406_));
 sg13g2_nor2_1 _10765_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ),
    .B(net49),
    .Y(_05407_));
 sg13g2_a21oi_1 _10766_ (.A1(net49),
    .A2(_05406_),
    .Y(_00557_),
    .B1(_05407_));
 sg13g2_nor2_1 _10767_ (.A(_02075_),
    .B(net74),
    .Y(_05408_));
 sg13g2_a21oi_1 _10768_ (.A1(_04170_),
    .A2(net74),
    .Y(_05409_),
    .B1(_05408_));
 sg13g2_nor2_1 _10769_ (.A(net135),
    .B(_03678_),
    .Y(_05410_));
 sg13g2_a21oi_1 _10770_ (.A1(\z80.tv80s.i_tv80_core.RegBusA_r[7] ),
    .A2(_05182_),
    .Y(_05411_),
    .B1(_05410_));
 sg13g2_o21ai_1 _10771_ (.B1(_05411_),
    .Y(_05412_),
    .A1(_05188_),
    .A2(_05409_));
 sg13g2_buf_2 _10772_ (.A(_05412_),
    .X(_05413_));
 sg13g2_mux2_1 _10773_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ),
    .A1(_05413_),
    .S(net49),
    .X(_00558_));
 sg13g2_nor2_1 _10774_ (.A(_03145_),
    .B(_03150_),
    .Y(_05414_));
 sg13g2_nor2_1 _10775_ (.A(_05414_),
    .B(_05352_),
    .Y(_05415_));
 sg13g2_buf_1 _10776_ (.A(_05415_),
    .X(_05416_));
 sg13g2_mux2_1 _10777_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ),
    .A1(_05348_),
    .S(net48),
    .X(_00559_));
 sg13g2_mux2_1 _10778_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ),
    .A1(_05362_),
    .S(net48),
    .X(_00560_));
 sg13g2_mux2_1 _10779_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .A1(_05373_),
    .S(_05416_),
    .X(_00561_));
 sg13g2_inv_1 _10780_ (.Y(_05417_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ));
 sg13g2_o21ai_1 _10781_ (.B1(_05415_),
    .Y(_05418_),
    .A1(_05378_),
    .A2(_05380_));
 sg13g2_o21ai_1 _10782_ (.B1(_05418_),
    .Y(_00562_),
    .A1(_05417_),
    .A2(_05416_));
 sg13g2_nor2_1 _10783_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ),
    .B(net48),
    .Y(_05419_));
 sg13g2_a21oi_1 _10784_ (.A1(_05392_),
    .A2(net48),
    .Y(_00563_),
    .B1(_05419_));
 sg13g2_nor2_1 _10785_ (.A(_05394_),
    .B(_05395_),
    .Y(_05420_));
 sg13g2_mux2_1 _10786_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ),
    .A1(_05420_),
    .S(net48),
    .X(_00564_));
 sg13g2_nor2_1 _10787_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ),
    .B(net48),
    .Y(_05421_));
 sg13g2_a21oi_1 _10788_ (.A1(_05406_),
    .A2(net48),
    .Y(_00565_),
    .B1(_05421_));
 sg13g2_mux2_1 _10789_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ),
    .A1(_05413_),
    .S(net48),
    .X(_00566_));
 sg13g2_nor2_1 _10790_ (.A(_05320_),
    .B(_05352_),
    .Y(_05422_));
 sg13g2_buf_1 _10791_ (.A(_05422_),
    .X(_05423_));
 sg13g2_mux2_1 _10792_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .A1(_05348_),
    .S(net47),
    .X(_00567_));
 sg13g2_mux2_1 _10793_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ),
    .A1(_05362_),
    .S(net47),
    .X(_00568_));
 sg13g2_mux2_1 _10794_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .A1(_05373_),
    .S(_05423_),
    .X(_00569_));
 sg13g2_inv_1 _10795_ (.Y(_05424_),
    .A(_05423_));
 sg13g2_nand2_1 _10796_ (.Y(_05425_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .B(_05424_));
 sg13g2_o21ai_1 _10797_ (.B1(_05425_),
    .Y(_00570_),
    .A1(_05383_),
    .A2(_05424_));
 sg13g2_nor2_1 _10798_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .B(net47),
    .Y(_05426_));
 sg13g2_a21oi_1 _10799_ (.A1(_05392_),
    .A2(net47),
    .Y(_00571_),
    .B1(_05426_));
 sg13g2_mux2_1 _10800_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ),
    .A1(_05398_),
    .S(net47),
    .X(_00572_));
 sg13g2_nor2_1 _10801_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .B(net47),
    .Y(_05427_));
 sg13g2_a21oi_1 _10802_ (.A1(_05406_),
    .A2(net47),
    .Y(_00573_),
    .B1(_05427_));
 sg13g2_mux2_1 _10803_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .A1(_05413_),
    .S(net47),
    .X(_00574_));
 sg13g2_nor2_1 _10804_ (.A(_05330_),
    .B(_05352_),
    .Y(_05428_));
 sg13g2_buf_1 _10805_ (.A(_05428_),
    .X(_05429_));
 sg13g2_mux2_1 _10806_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .A1(_05348_),
    .S(net46),
    .X(_00575_));
 sg13g2_mux2_1 _10807_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .A1(_05362_),
    .S(net46),
    .X(_00576_));
 sg13g2_mux2_1 _10808_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .A1(_05373_),
    .S(_05429_),
    .X(_00577_));
 sg13g2_inv_1 _10809_ (.Y(_05430_),
    .A(net46));
 sg13g2_nand2_1 _10810_ (.Y(_05431_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .B(_05430_));
 sg13g2_o21ai_1 _10811_ (.B1(_05431_),
    .Y(_00578_),
    .A1(_05383_),
    .A2(_05430_));
 sg13g2_nor2_1 _10812_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .B(net46),
    .Y(_05432_));
 sg13g2_a21oi_1 _10813_ (.A1(_05392_),
    .A2(net46),
    .Y(_00579_),
    .B1(_05432_));
 sg13g2_mux2_1 _10814_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .A1(_05398_),
    .S(_05429_),
    .X(_00580_));
 sg13g2_nor2_1 _10815_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .B(net46),
    .Y(_05433_));
 sg13g2_a21oi_1 _10816_ (.A1(_05406_),
    .A2(net46),
    .Y(_00581_),
    .B1(_05433_));
 sg13g2_mux2_1 _10817_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ),
    .A1(_05413_),
    .S(net46),
    .X(_00582_));
 sg13g2_or2_1 _10818_ (.X(_05434_),
    .B(_05350_),
    .A(_03186_));
 sg13g2_buf_1 _10819_ (.A(_05434_),
    .X(_05435_));
 sg13g2_nor2_1 _10820_ (.A(_03189_),
    .B(_05435_),
    .Y(_05436_));
 sg13g2_buf_1 _10821_ (.A(_05436_),
    .X(_05437_));
 sg13g2_mux2_1 _10822_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .A1(_05348_),
    .S(net45),
    .X(_00583_));
 sg13g2_mux2_1 _10823_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ),
    .A1(_05362_),
    .S(net45),
    .X(_00584_));
 sg13g2_mux2_1 _10824_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .A1(_05373_),
    .S(_05437_),
    .X(_00585_));
 sg13g2_inv_1 _10825_ (.Y(_05438_),
    .A(_05437_));
 sg13g2_nand2_1 _10826_ (.Y(_05439_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ),
    .B(_05438_));
 sg13g2_o21ai_1 _10827_ (.B1(_05439_),
    .Y(_00586_),
    .A1(_05383_),
    .A2(_05438_));
 sg13g2_nor2_1 _10828_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ),
    .B(net45),
    .Y(_05440_));
 sg13g2_a21oi_1 _10829_ (.A1(_05392_),
    .A2(net45),
    .Y(_00587_),
    .B1(_05440_));
 sg13g2_mux2_1 _10830_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ),
    .A1(_05398_),
    .S(net45),
    .X(_00588_));
 sg13g2_nor2_1 _10831_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ),
    .B(net45),
    .Y(_05441_));
 sg13g2_a21oi_1 _10832_ (.A1(_05406_),
    .A2(net45),
    .Y(_00589_),
    .B1(_05441_));
 sg13g2_mux2_1 _10833_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ),
    .A1(_05413_),
    .S(net45),
    .X(_00590_));
 sg13g2_nor2_1 _10834_ (.A(_05414_),
    .B(_05435_),
    .Y(_05442_));
 sg13g2_buf_1 _10835_ (.A(_05442_),
    .X(_05443_));
 sg13g2_mux2_1 _10836_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .A1(_05348_),
    .S(_05443_),
    .X(_00591_));
 sg13g2_mux2_1 _10837_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .A1(_05362_),
    .S(net44),
    .X(_00592_));
 sg13g2_mux2_1 _10838_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .A1(_05373_),
    .S(_05443_),
    .X(_00593_));
 sg13g2_inv_1 _10839_ (.Y(_05444_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ));
 sg13g2_o21ai_1 _10840_ (.B1(_05442_),
    .Y(_05445_),
    .A1(_05378_),
    .A2(_05380_));
 sg13g2_o21ai_1 _10841_ (.B1(_05445_),
    .Y(_00594_),
    .A1(_05444_),
    .A2(net44));
 sg13g2_nor2_1 _10842_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ),
    .B(net44),
    .Y(_05446_));
 sg13g2_a21oi_1 _10843_ (.A1(_05392_),
    .A2(net44),
    .Y(_00595_),
    .B1(_05446_));
 sg13g2_mux2_1 _10844_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ),
    .A1(_05420_),
    .S(net44),
    .X(_00596_));
 sg13g2_nor2_1 _10845_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ),
    .B(net44),
    .Y(_05447_));
 sg13g2_a21oi_1 _10846_ (.A1(_05406_),
    .A2(net44),
    .Y(_00597_),
    .B1(_05447_));
 sg13g2_mux2_1 _10847_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ),
    .A1(_05413_),
    .S(net44),
    .X(_00598_));
 sg13g2_nor2_1 _10848_ (.A(_05320_),
    .B(_05435_),
    .Y(_05448_));
 sg13g2_buf_1 _10849_ (.A(_05448_),
    .X(_05449_));
 sg13g2_mux2_1 _10850_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .A1(_05348_),
    .S(net43),
    .X(_00599_));
 sg13g2_mux2_1 _10851_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ),
    .A1(_05362_),
    .S(net43),
    .X(_00600_));
 sg13g2_mux2_1 _10852_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .A1(_05373_),
    .S(_05449_),
    .X(_00601_));
 sg13g2_inv_1 _10853_ (.Y(_05450_),
    .A(_05449_));
 sg13g2_nand2_1 _10854_ (.Y(_05451_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .B(_05450_));
 sg13g2_o21ai_1 _10855_ (.B1(_05451_),
    .Y(_00602_),
    .A1(_05383_),
    .A2(_05450_));
 sg13g2_nor2_1 _10856_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .B(net43),
    .Y(_05452_));
 sg13g2_a21oi_1 _10857_ (.A1(_05392_),
    .A2(net43),
    .Y(_00603_),
    .B1(_05452_));
 sg13g2_mux2_1 _10858_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .A1(_05398_),
    .S(net43),
    .X(_00604_));
 sg13g2_nor2_1 _10859_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ),
    .B(net43),
    .Y(_05453_));
 sg13g2_a21oi_1 _10860_ (.A1(_05406_),
    .A2(net43),
    .Y(_00605_),
    .B1(_05453_));
 sg13g2_mux2_1 _10861_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ),
    .A1(_05413_),
    .S(net43),
    .X(_00606_));
 sg13g2_nor3_1 _10862_ (.A(_03186_),
    .B(_05330_),
    .C(_05350_),
    .Y(_05454_));
 sg13g2_buf_1 _10863_ (.A(_05454_),
    .X(_05455_));
 sg13g2_mux2_1 _10864_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .A1(_05348_),
    .S(net57),
    .X(_00607_));
 sg13g2_mux2_1 _10865_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ),
    .A1(_05362_),
    .S(net57),
    .X(_00608_));
 sg13g2_mux2_1 _10866_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ),
    .A1(_05373_),
    .S(_05455_),
    .X(_00609_));
 sg13g2_inv_1 _10867_ (.Y(_05456_),
    .A(_05455_));
 sg13g2_nand2_1 _10868_ (.Y(_05457_),
    .A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ),
    .B(_05456_));
 sg13g2_o21ai_1 _10869_ (.B1(_05457_),
    .Y(_00610_),
    .A1(_05383_),
    .A2(_05456_));
 sg13g2_nor2_1 _10870_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .B(net57),
    .Y(_05458_));
 sg13g2_a21oi_1 _10871_ (.A1(_05392_),
    .A2(net57),
    .Y(_00611_),
    .B1(_05458_));
 sg13g2_mux2_1 _10872_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .A1(_05398_),
    .S(net57),
    .X(_00612_));
 sg13g2_nor2_1 _10873_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .B(net57),
    .Y(_05459_));
 sg13g2_a21oi_1 _10874_ (.A1(_05406_),
    .A2(net57),
    .Y(_00613_),
    .B1(_05459_));
 sg13g2_mux2_1 _10875_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ),
    .A1(_05413_),
    .S(net57),
    .X(_00614_));
 sg13g2_nor2_1 _10876_ (.A(\z80.m1_n ),
    .B(_01320_),
    .Y(_05460_));
 sg13g2_nor3_1 _10877_ (.A(\z80.tv80s.i_tv80_core.ts[0] ),
    .B(_04207_),
    .C(_05460_),
    .Y(_05461_));
 sg13g2_nor2_1 _10878_ (.A(net326),
    .B(_00269_),
    .Y(_05462_));
 sg13g2_a21oi_1 _10879_ (.A1(net328),
    .A2(_05461_),
    .Y(_00615_),
    .B1(_05462_));
 sg13g2_buf_1 _10880_ (.A(_01013_),
    .X(_05463_));
 sg13g2_buf_1 _10881_ (.A(_00218_),
    .X(_05464_));
 sg13g2_buf_1 _10882_ (.A(_00219_),
    .X(_05465_));
 sg13g2_and3_1 _10883_ (.X(_05466_),
    .A(_05464_),
    .B(_05465_),
    .C(_00220_));
 sg13g2_nor3_1 _10884_ (.A(_05464_),
    .B(_05465_),
    .C(_00220_),
    .Y(_05467_));
 sg13g2_o21ai_1 _10885_ (.B1(net353),
    .Y(_05468_),
    .A1(_05466_),
    .A2(_05467_));
 sg13g2_a21oi_1 _10886_ (.A1(_04201_),
    .A2(_05468_),
    .Y(_05469_),
    .B1(net72));
 sg13g2_nand2_1 _10887_ (.Y(_05470_),
    .A(_00270_),
    .B(net73));
 sg13g2_o21ai_1 _10888_ (.B1(_05470_),
    .Y(_00616_),
    .A1(net73),
    .A2(_05469_));
 sg13g2_nor2b_1 _10889_ (.A(_05465_),
    .B_N(_05464_),
    .Y(_05471_));
 sg13g2_nor2_1 _10890_ (.A(net302),
    .B(_00220_),
    .Y(_05472_));
 sg13g2_a22oi_1 _10891_ (.Y(_05473_),
    .B1(_05471_),
    .B2(_05472_),
    .A2(net302),
    .A1(_02204_));
 sg13g2_nor2b_1 _10892_ (.A(net72),
    .B_N(_04201_),
    .Y(_05474_));
 sg13g2_nand2b_1 _10893_ (.Y(_05475_),
    .B(_05474_),
    .A_N(_05473_));
 sg13g2_nand2_1 _10894_ (.Y(_05476_),
    .A(_01017_),
    .B(net73));
 sg13g2_o21ai_1 _10895_ (.B1(_05476_),
    .Y(_00617_),
    .A1(_05463_),
    .A2(_05475_));
 sg13g2_inv_1 _10896_ (.Y(_05477_),
    .A(_04200_));
 sg13g2_nor2b_1 _10897_ (.A(_05464_),
    .B_N(_05465_),
    .Y(_05478_));
 sg13g2_a22oi_1 _10898_ (.Y(_05479_),
    .B1(_05472_),
    .B2(_05478_),
    .A2(_05477_),
    .A1(_00867_));
 sg13g2_or3_1 _10899_ (.A(_05463_),
    .B(net72),
    .C(_05479_),
    .X(_05480_));
 sg13g2_o21ai_1 _10900_ (.B1(_05480_),
    .Y(_00618_),
    .A1(_00924_),
    .A2(_01211_));
 sg13g2_nand3_1 _10901_ (.B(_05465_),
    .C(_05472_),
    .A(_05464_),
    .Y(_05481_));
 sg13g2_o21ai_1 _10902_ (.B1(_05481_),
    .Y(_05482_),
    .A1(_00924_),
    .A2(net353));
 sg13g2_nand3_1 _10903_ (.B(_05474_),
    .C(_05482_),
    .A(_01211_),
    .Y(_05483_));
 sg13g2_o21ai_1 _10904_ (.B1(_05483_),
    .Y(_00619_),
    .A1(_00851_),
    .A2(_01211_));
 sg13g2_nor2_1 _10905_ (.A(_05464_),
    .B(_05465_),
    .Y(_05484_));
 sg13g2_and2_1 _10906_ (.A(net353),
    .B(_00220_),
    .X(_05485_));
 sg13g2_buf_1 _10907_ (.A(_05485_),
    .X(_05486_));
 sg13g2_a22oi_1 _10908_ (.Y(_05487_),
    .B1(_05484_),
    .B2(_05486_),
    .A2(net302),
    .A1(_00850_));
 sg13g2_nand2b_1 _10909_ (.Y(_05488_),
    .B(_05474_),
    .A_N(_05487_));
 sg13g2_nand2_1 _10910_ (.Y(_05489_),
    .A(_00852_),
    .B(net73));
 sg13g2_o21ai_1 _10911_ (.B1(_05489_),
    .Y(_00620_),
    .A1(net73),
    .A2(_05488_));
 sg13g2_nor2_1 _10912_ (.A(_00028_),
    .B(_04200_),
    .Y(_05490_));
 sg13g2_a221oi_1 _10913_ (.B2(_01216_),
    .C1(net72),
    .B1(_05490_),
    .A1(_05471_),
    .Y(_05491_),
    .A2(_05486_));
 sg13g2_nand2_1 _10914_ (.Y(_05492_),
    .A(_01008_),
    .B(net73));
 sg13g2_o21ai_1 _10915_ (.B1(_05492_),
    .Y(_00621_),
    .A1(net73),
    .A2(_05491_));
 sg13g2_nand2_1 _10916_ (.Y(_05493_),
    .A(_05478_),
    .B(_05486_));
 sg13g2_a21oi_1 _10917_ (.A1(_01217_),
    .A2(_05493_),
    .Y(_05494_),
    .B1(_01206_));
 sg13g2_o21ai_1 _10918_ (.B1(_01216_),
    .Y(_05495_),
    .A1(_01013_),
    .A2(_04200_));
 sg13g2_o21ai_1 _10919_ (.B1(_05495_),
    .Y(_05496_),
    .A1(net73),
    .A2(_05494_));
 sg13g2_inv_1 _10920_ (.Y(_00622_),
    .A(_05496_));
 sg13g2_a21oi_1 _10921_ (.A1(_01307_),
    .A2(_01319_),
    .Y(_05497_),
    .B1(net215));
 sg13g2_mux2_1 _10922_ (.A0(_00271_),
    .A1(_05497_),
    .S(net326),
    .X(_00623_));
 sg13g2_inv_1 _10923_ (.Y(_05498_),
    .A(_00272_));
 sg13g2_nand2b_1 _10924_ (.Y(_05499_),
    .B(_02886_),
    .A_N(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ));
 sg13g2_o21ai_1 _10925_ (.B1(_05499_),
    .Y(_05500_),
    .A1(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ),
    .A2(_02874_));
 sg13g2_nand2_1 _10926_ (.Y(_05501_),
    .A(_00031_),
    .B(net115));
 sg13g2_o21ai_1 _10927_ (.B1(_05501_),
    .Y(_05502_),
    .A1(net115),
    .A2(_05500_));
 sg13g2_nand4_1 _10928_ (.B(_00997_),
    .C(_00999_),
    .A(net399),
    .Y(_05503_),
    .D(_05502_));
 sg13g2_buf_1 _10929_ (.A(_05503_),
    .X(_05504_));
 sg13g2_buf_1 _10930_ (.A(_05504_),
    .X(_05505_));
 sg13g2_nor3_1 _10931_ (.A(_00030_),
    .B(net100),
    .C(_05505_),
    .Y(_05506_));
 sg13g2_a21oi_1 _10932_ (.A1(_05498_),
    .A2(net56),
    .Y(_00624_),
    .B1(_05506_));
 sg13g2_nor3_1 _10933_ (.A(\z80.tv80s.i_tv80_core.ts[0] ),
    .B(net100),
    .C(_05504_),
    .Y(_05507_));
 sg13g2_a21oi_1 _10934_ (.A1(_05092_),
    .A2(net56),
    .Y(_00625_),
    .B1(_05507_));
 sg13g2_nor3_1 _10935_ (.A(_03755_),
    .B(_02089_),
    .C(_05504_),
    .Y(_05508_));
 sg13g2_a21o_1 _10936_ (.A2(_05505_),
    .A1(net398),
    .B1(_05508_),
    .X(_00626_));
 sg13g2_nor3_1 _10937_ (.A(_00032_),
    .B(_02089_),
    .C(_05504_),
    .Y(_05509_));
 sg13g2_a21o_1 _10938_ (.A2(net56),
    .A1(_04549_),
    .B1(_05509_),
    .X(_00627_));
 sg13g2_nor3_1 _10939_ (.A(_01307_),
    .B(net115),
    .C(_05504_),
    .Y(_05510_));
 sg13g2_a21o_1 _10940_ (.A2(net56),
    .A1(net393),
    .B1(_05510_),
    .X(_00628_));
 sg13g2_nand2_1 _10941_ (.Y(_05511_),
    .A(_00905_),
    .B(net104));
 sg13g2_nand2_1 _10942_ (.Y(_05512_),
    .A(\z80.tv80s.i_tv80_core.ts[5] ),
    .B(net56));
 sg13g2_o21ai_1 _10943_ (.B1(_05512_),
    .Y(_00629_),
    .A1(net56),
    .A2(_05511_));
 sg13g2_nand2_1 _10944_ (.Y(_05513_),
    .A(\z80.tv80s.i_tv80_core.ts[5] ),
    .B(net104));
 sg13g2_nand2_1 _10945_ (.Y(_05514_),
    .A(\z80.tv80s.i_tv80_core.ts[6] ),
    .B(net56));
 sg13g2_o21ai_1 _10946_ (.B1(_05514_),
    .Y(_00630_),
    .A1(net56),
    .A2(_05513_));
 sg13g2_a21oi_1 _10947_ (.A1(_03755_),
    .A2(_00997_),
    .Y(_05515_),
    .B1(_02276_));
 sg13g2_nand2_1 _10948_ (.Y(_05516_),
    .A(_03755_),
    .B(_00997_));
 sg13g2_nand2_1 _10949_ (.Y(_05517_),
    .A(doe),
    .B(_05516_));
 sg13g2_o21ai_1 _10950_ (.B1(_00955_),
    .Y(_05518_),
    .A1(net201),
    .A2(_03447_));
 sg13g2_nand2_1 _10951_ (.Y(_05519_),
    .A(net241),
    .B(_05518_));
 sg13g2_a21o_1 _10952_ (.A2(_05519_),
    .A1(_02871_),
    .B1(net305),
    .X(_05520_));
 sg13g2_nor2_1 _10953_ (.A(net232),
    .B(_01146_),
    .Y(_05521_));
 sg13g2_a21oi_1 _10954_ (.A1(net232),
    .A2(_01369_),
    .Y(_05522_),
    .B1(_05521_));
 sg13g2_nor3_1 _10955_ (.A(net201),
    .B(_01119_),
    .C(_05522_),
    .Y(_05523_));
 sg13g2_a221oi_1 _10956_ (.B2(_01296_),
    .C1(_05523_),
    .B1(_02091_),
    .A1(net170),
    .Y(_05524_),
    .A2(net219));
 sg13g2_nand2b_1 _10957_ (.Y(_05525_),
    .B(net224),
    .A_N(_05524_));
 sg13g2_nand3b_1 _10958_ (.B(_00034_),
    .C(_01014_),
    .Y(_05526_),
    .A_N(_01028_));
 sg13g2_nand4_1 _10959_ (.B(_05520_),
    .C(_05525_),
    .A(_05516_),
    .Y(_05527_),
    .D(_05526_));
 sg13g2_nand2_1 _10960_ (.Y(_05528_),
    .A(_05517_),
    .B(_05527_));
 sg13g2_and2_1 _10961_ (.A(net215),
    .B(_02886_),
    .X(_05529_));
 sg13g2_a22oi_1 _10962_ (.Y(_05530_),
    .B1(_05528_),
    .B2(_05529_),
    .A2(_05515_),
    .A1(net166));
 sg13g2_nor2_1 _10963_ (.A(net326),
    .B(_00273_),
    .Y(_05531_));
 sg13g2_a21oi_1 _10964_ (.A1(net328),
    .A2(_05530_),
    .Y(_00631_),
    .B1(_05531_));
 sg13g2_nand2_1 _10965_ (.Y(_05532_),
    .A(_02276_),
    .B(_05516_));
 sg13g2_nand2b_1 _10966_ (.Y(_05533_),
    .B(_05528_),
    .A_N(_02886_));
 sg13g2_a22oi_1 _10967_ (.Y(_05534_),
    .B1(_05533_),
    .B2(net215),
    .A2(_05532_),
    .A1(_05176_));
 sg13g2_mux2_1 _10968_ (.A0(_00274_),
    .A1(_05534_),
    .S(net326),
    .X(_00632_));
 sg13g2_and2_1 _10969_ (.A(_02276_),
    .B(_05516_),
    .X(_05535_));
 sg13g2_nor3_1 _10970_ (.A(net166),
    .B(doe),
    .C(_05527_),
    .Y(_05536_));
 sg13g2_a21oi_1 _10971_ (.A1(net166),
    .A2(_05535_),
    .Y(_05537_),
    .B1(_05536_));
 sg13g2_nor2_1 _10972_ (.A(net399),
    .B(_00275_),
    .Y(_05538_));
 sg13g2_a21oi_1 _10973_ (.A1(net328),
    .A2(_05537_),
    .Y(_00633_),
    .B1(_05538_));
 sg13g2_nor2_1 _10974_ (.A(net166),
    .B(_05517_),
    .Y(_05539_));
 sg13g2_mux2_1 _10975_ (.A0(_00276_),
    .A1(_05539_),
    .S(net326),
    .X(_00634_));
 sg13g2_nor3_1 _10976_ (.A(net300),
    .B(_01132_),
    .C(_01421_),
    .Y(_05540_));
 sg13g2_nand4_1 _10977_ (.B(_04196_),
    .C(_05078_),
    .A(_02259_),
    .Y(_05541_),
    .D(_05540_));
 sg13g2_a221oi_1 _10978_ (.B2(net354),
    .C1(_00214_),
    .B1(_01344_),
    .A1(net166),
    .Y(_05542_),
    .A2(_01593_));
 sg13g2_o21ai_1 _10979_ (.B1(net211),
    .Y(_05543_),
    .A1(_01320_),
    .A2(_05542_));
 sg13g2_a22oi_1 _10980_ (.Y(_00277_),
    .B1(_05543_),
    .B2(net265),
    .A2(_05541_),
    .A1(_01317_));
 sg13g2_buf_1 _10981_ (.A(ui_in[7]),
    .X(_05544_));
 sg13g2_buf_1 _10982_ (.A(_05544_),
    .X(_05545_));
 sg13g2_buf_1 _10983_ (.A(ui_in[6]),
    .X(_05546_));
 sg13g2_buf_1 _10984_ (.A(_05546_),
    .X(_05547_));
 sg13g2_nor2b_1 _10985_ (.A(_05547_),
    .B_N(\addr_bus[0] ),
    .Y(_05548_));
 sg13g2_a21oi_1 _10986_ (.A1(\addr_bus[8] ),
    .A2(net370),
    .Y(_05549_),
    .B1(_05548_));
 sg13g2_nand2_1 _10987_ (.Y(_05550_),
    .A(\z80.m1_n ),
    .B(_05544_));
 sg13g2_o21ai_1 _10988_ (.B1(_05550_),
    .Y(net30),
    .A1(net371),
    .A2(_05549_));
 sg13g2_nor2b_1 _10989_ (.A(net370),
    .B_N(\addr_bus[1] ),
    .Y(_05551_));
 sg13g2_a21oi_1 _10990_ (.A1(net370),
    .A2(\addr_bus[9] ),
    .Y(_05552_),
    .B1(_05551_));
 sg13g2_nand2_1 _10991_ (.Y(_05553_),
    .A(_05545_),
    .B(\z80.mreq_n ));
 sg13g2_o21ai_1 _10992_ (.B1(_05553_),
    .Y(net31),
    .A1(_05545_),
    .A2(_05552_));
 sg13g2_nor2b_1 _10993_ (.A(net370),
    .B_N(\addr_bus[2] ),
    .Y(_05554_));
 sg13g2_a21oi_1 _10994_ (.A1(_05547_),
    .A2(\addr_bus[10] ),
    .Y(_05555_),
    .B1(_05554_));
 sg13g2_nand2_1 _10995_ (.Y(_05556_),
    .A(net371),
    .B(\z80.iorq_n ));
 sg13g2_o21ai_1 _10996_ (.B1(_05556_),
    .Y(net32),
    .A1(net371),
    .A2(_05555_));
 sg13g2_nor2b_1 _10997_ (.A(_05546_),
    .B_N(\addr_bus[3] ),
    .Y(_05557_));
 sg13g2_a21oi_1 _10998_ (.A1(net370),
    .A2(\addr_bus[11] ),
    .Y(_05558_),
    .B1(_05557_));
 sg13g2_nand2_1 _10999_ (.Y(_05559_),
    .A(_05544_),
    .B(\z80.rd_n ));
 sg13g2_o21ai_1 _11000_ (.B1(_05559_),
    .Y(net33),
    .A1(net371),
    .A2(_05558_));
 sg13g2_nor2b_1 _11001_ (.A(_05546_),
    .B_N(\addr_bus[4] ),
    .Y(_05560_));
 sg13g2_a21oi_1 _11002_ (.A1(net370),
    .A2(\addr_bus[12] ),
    .Y(_05561_),
    .B1(_05560_));
 sg13g2_nand2_1 _11003_ (.Y(_05562_),
    .A(_05544_),
    .B(\z80.tv80s.wr_n ));
 sg13g2_o21ai_1 _11004_ (.B1(_05562_),
    .Y(net34),
    .A1(net371),
    .A2(_05561_));
 sg13g2_nor2b_1 _11005_ (.A(_05546_),
    .B_N(\addr_bus[5] ),
    .Y(_05563_));
 sg13g2_a21oi_1 _11006_ (.A1(net370),
    .A2(\addr_bus[13] ),
    .Y(_05564_),
    .B1(_05563_));
 sg13g2_nand2_1 _11007_ (.Y(_05565_),
    .A(_05544_),
    .B(\z80.rfsh_n ));
 sg13g2_o21ai_1 _11008_ (.B1(_05565_),
    .Y(net35),
    .A1(net371),
    .A2(_05564_));
 sg13g2_mux2_1 _11009_ (.A0(\addr_bus[6] ),
    .A1(\addr_bus[14] ),
    .S(_05546_),
    .X(_05566_));
 sg13g2_nor2_1 _11010_ (.A(_05544_),
    .B(_05566_),
    .Y(_05567_));
 sg13g2_a21oi_1 _11011_ (.A1(_03974_),
    .A2(net371),
    .Y(net36),
    .B1(_05567_));
 sg13g2_nor2b_1 _11012_ (.A(_05546_),
    .B_N(\addr_bus[7] ),
    .Y(_05568_));
 sg13g2_a21oi_1 _11013_ (.A1(net370),
    .A2(\addr_bus[15] ),
    .Y(_05569_),
    .B1(_05568_));
 sg13g2_nand2_1 _11014_ (.Y(_05570_),
    .A(_05544_),
    .B(_00036_));
 sg13g2_o21ai_1 _11015_ (.B1(_05570_),
    .Y(net37),
    .A1(net371),
    .A2(_05569_));
 sg13g2_dfrbp_1 _11016_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net430),
    .D(_00017_),
    .Q_N(_05678_),
    .Q(_00218_));
 sg13g2_dfrbp_1 _11017_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net430),
    .D(_00018_),
    .Q_N(_05679_),
    .Q(_00219_));
 sg13g2_dfrbp_1 _11018_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net430),
    .D(_00019_),
    .Q_N(_05677_),
    .Q(_00220_));
 sg13g2_buf_4 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_1 _11020_ (.A(net146),
    .X(net14));
 sg13g2_buf_1 _11021_ (.A(net146),
    .X(net15));
 sg13g2_buf_1 _11022_ (.A(net146),
    .X(net16));
 sg13g2_buf_1 _11023_ (.A(net146),
    .X(net17));
 sg13g2_buf_1 _11024_ (.A(net146),
    .X(net18));
 sg13g2_buf_1 _11025_ (.A(net146),
    .X(net19));
 sg13g2_buf_1 _11026_ (.A(net146),
    .X(net20));
 sg13g2_buf_1 _11027_ (.A(net146),
    .X(net21));
 sg13g2_dfrbp_1 \z80.tv80s.di_reg[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net418),
    .D(_00278_),
    .Q_N(_00137_),
    .Q(\z80.tv80s.di_reg[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.di_reg[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net416),
    .D(_00279_),
    .Q_N(_00140_),
    .Q(\z80.tv80s.di_reg[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.di_reg[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net413),
    .D(_00280_),
    .Q_N(_00143_),
    .Q(\z80.tv80s.di_reg[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.di_reg[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net413),
    .D(_00281_),
    .Q_N(_00146_),
    .Q(\z80.tv80s.di_reg[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.di_reg[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net413),
    .D(_00282_),
    .Q_N(_00149_),
    .Q(\z80.tv80s.di_reg[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.di_reg[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net413),
    .D(_00283_),
    .Q_N(_00152_),
    .Q(\z80.tv80s.di_reg[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.di_reg[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net415),
    .D(_00284_),
    .Q_N(_00155_),
    .Q(\z80.tv80s.di_reg[6] ));
 sg13g2_dfrbp_1 \z80.tv80s.di_reg[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net413),
    .D(_00285_),
    .Q_N(_00158_),
    .Q(\z80.tv80s.di_reg[7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ACC[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net412),
    .D(_00286_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[0] ),
    .Q(_00221_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ACC[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net412),
    .D(_00287_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[1] ),
    .Q(_00222_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ACC[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net414),
    .D(_00288_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[2] ),
    .Q(_00223_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ACC[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net412),
    .D(_00289_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[3] ),
    .Q(_00224_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ACC[4]$_DFFE_PN1P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net414),
    .D(_00290_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[4] ),
    .Q(_00225_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ACC[5]$_DFFE_PN1P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net414),
    .D(_00291_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[5] ),
    .Q(_00226_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ACC[6]$_DFFE_PN1P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net414),
    .D(_00292_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[6] ),
    .Q(_00227_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ACC[7]$_DFFE_PN1P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net414),
    .D(_00293_),
    .Q_N(\z80.tv80s.i_tv80_core.ACC[7] ),
    .Q(_00228_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ALU_Op_r[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net433),
    .D(_00294_),
    .Q_N(_05676_),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ALU_Op_r[1]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net433),
    .D(_00295_),
    .Q_N(_05675_),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ALU_Op_r[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net433),
    .D(_00296_),
    .Q_N(_00208_),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ALU_Op_r[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net433),
    .D(_00297_),
    .Q_N(_05674_),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net416),
    .D(_00298_),
    .Q_N(_05673_),
    .Q(\addr_bus[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net409),
    .D(_00299_),
    .Q_N(_05672_),
    .Q(\addr_bus[10] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net406),
    .D(_00300_),
    .Q_N(_05671_),
    .Q(\addr_bus[11] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net406),
    .D(_00301_),
    .Q_N(_05670_),
    .Q(\addr_bus[12] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net404),
    .D(_00302_),
    .Q_N(_05669_),
    .Q(\addr_bus[13] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net404),
    .D(_00303_),
    .Q_N(_05668_),
    .Q(\addr_bus[14] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net406),
    .D(_00304_),
    .Q_N(_05667_),
    .Q(\addr_bus[15] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net417),
    .D(_00305_),
    .Q_N(_05666_),
    .Q(\addr_bus[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net406),
    .D(_00306_),
    .Q_N(_05665_),
    .Q(\addr_bus[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net417),
    .D(_00307_),
    .Q_N(_05664_),
    .Q(\addr_bus[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net417),
    .D(_00308_),
    .Q_N(_05663_),
    .Q(\addr_bus[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net409),
    .D(_00309_),
    .Q_N(_05662_),
    .Q(\addr_bus[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net410),
    .D(_00310_),
    .Q_N(_05661_),
    .Q(\addr_bus[6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net416),
    .D(_00311_),
    .Q_N(_05660_),
    .Q(\addr_bus[7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net404),
    .D(_00312_),
    .Q_N(_05659_),
    .Q(\addr_bus[8] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.A[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net416),
    .D(_00313_),
    .Q_N(_05658_),
    .Q(\addr_bus[9] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Alternate$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net426),
    .D(_00314_),
    .Q_N(_00020_),
    .Q(\z80.tv80s.i_tv80_core.Alternate ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Ap[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net419),
    .D(_00315_),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[0] ),
    .Q(_00229_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Ap[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net419),
    .D(_00316_),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[1] ),
    .Q(_00230_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Ap[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net419),
    .D(_00317_),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[2] ),
    .Q(_00231_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Ap[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net419),
    .D(_00318_),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[3] ),
    .Q(_00232_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Ap[4]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net419),
    .D(_00319_),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[4] ),
    .Q(_00233_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Ap[5]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net420),
    .D(_00320_),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[5] ),
    .Q(_00234_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Ap[6]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net419),
    .D(_00321_),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[6] ),
    .Q(_00235_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Ap[7]$_DFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net419),
    .D(_00322_),
    .Q_N(\z80.tv80s.i_tv80_core.Ap[7] ),
    .Q(_00236_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Arith16_r$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net424),
    .D(_00323_),
    .Q_N(_05657_),
    .Q(\z80.tv80s.i_tv80_core.Arith16_r ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Auto_Wait_t1$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net421),
    .D(_00324_),
    .Q_N(_00209_),
    .Q(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Auto_Wait_t2$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net421),
    .D(_00325_),
    .Q_N(_05656_),
    .Q(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BTR_r$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net410),
    .D(_00326_),
    .Q_N(_00211_),
    .Q(\z80.tv80s.i_tv80_core.BTR_r ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusA[0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net436),
    .D(_00327_),
    .Q_N(_00194_),
    .Q(\z80.tv80s.i_tv80_core.BusA[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusA[1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net437),
    .D(_00328_),
    .Q_N(_00192_),
    .Q(\z80.tv80s.i_tv80_core.BusA[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusA[2]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net438),
    .D(_00329_),
    .Q_N(_00195_),
    .Q(\z80.tv80s.i_tv80_core.BusA[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusA[3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net439),
    .D(_00330_),
    .Q_N(_00196_),
    .Q(\z80.tv80s.i_tv80_core.BusA[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusA[4]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net440),
    .D(_00331_),
    .Q_N(_00197_),
    .Q(\z80.tv80s.i_tv80_core.BusA[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusA[5]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net441),
    .D(_00332_),
    .Q_N(_00198_),
    .Q(\z80.tv80s.i_tv80_core.BusA[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusA[6]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net442),
    .D(_00333_),
    .Q_N(_00199_),
    .Q(\z80.tv80s.i_tv80_core.BusA[6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusA[7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net443),
    .D(_00334_),
    .Q_N(_00193_),
    .Q(\z80.tv80s.i_tv80_core.BusA[7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusAck$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net421),
    .D(_00335_),
    .Q_N(_00036_),
    .Q(\z80.tv80s.i_tv80_core.BusAck ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusB[0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net444),
    .D(_00336_),
    .Q_N(_00200_),
    .Q(\z80.tv80s.i_tv80_core.BusB[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusB[1]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net445),
    .D(_00337_),
    .Q_N(_00201_),
    .Q(\z80.tv80s.i_tv80_core.BusB[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusB[2]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net446),
    .D(_00338_),
    .Q_N(_00202_),
    .Q(\z80.tv80s.i_tv80_core.BusB[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusB[3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net447),
    .D(_00339_),
    .Q_N(_00203_),
    .Q(\z80.tv80s.i_tv80_core.BusB[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusB[4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net448),
    .D(_00340_),
    .Q_N(_00204_),
    .Q(\z80.tv80s.i_tv80_core.BusB[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusB[5]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net449),
    .D(_00341_),
    .Q_N(_00205_),
    .Q(\z80.tv80s.i_tv80_core.BusB[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusB[6]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net450),
    .D(_00342_),
    .Q_N(_00206_),
    .Q(\z80.tv80s.i_tv80_core.BusB[6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusB[7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net451),
    .D(_00343_),
    .Q_N(_00207_),
    .Q(\z80.tv80s.i_tv80_core.BusB[7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.BusReq_s$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net422),
    .D(_00344_),
    .Q_N(_00031_),
    .Q(\z80.tv80s.i_tv80_core.BusReq_s ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.F[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net424),
    .D(_00345_),
    .Q_N(\z80.tv80s.i_tv80_core.F[0] ),
    .Q(_00237_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.F[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net425),
    .D(_00346_),
    .Q_N(\z80.tv80s.i_tv80_core.F[1] ),
    .Q(_00238_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.F[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net424),
    .D(_00347_),
    .Q_N(\z80.tv80s.i_tv80_core.F[2] ),
    .Q(_00239_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.F[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net425),
    .D(_00348_),
    .Q_N(\z80.tv80s.i_tv80_core.F[3] ),
    .Q(_00240_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.F[4]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net425),
    .D(_00349_),
    .Q_N(\z80.tv80s.i_tv80_core.F[4] ),
    .Q(_00241_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.F[5]$_DFFE_PN1P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net424),
    .D(_00350_),
    .Q_N(\z80.tv80s.i_tv80_core.F[5] ),
    .Q(_00242_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.F[6]$_DFFE_PN1P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net425),
    .D(_00351_),
    .Q_N(\z80.tv80s.i_tv80_core.F[6] ),
    .Q(_00243_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.F[7]$_DFFE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net413),
    .D(_00352_),
    .Q_N(\z80.tv80s.i_tv80_core.F[7] ),
    .Q(_00244_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Fp[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net413),
    .D(_00353_),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[0] ),
    .Q(_00245_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Fp[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net424),
    .D(_00354_),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[1] ),
    .Q(_00246_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Fp[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net420),
    .D(_00355_),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[2] ),
    .Q(_00247_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Fp[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net413),
    .D(_00356_),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[3] ),
    .Q(_00248_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Fp[4]$_DFFE_PN1P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net424),
    .D(_00357_),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[4] ),
    .Q(_00249_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Fp[5]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net415),
    .D(_00358_),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[5] ),
    .Q(_00250_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Fp[6]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net420),
    .D(_00359_),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[6] ),
    .Q(_00251_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Fp[7]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net420),
    .D(_00360_),
    .Q_N(\z80.tv80s.i_tv80_core.Fp[7] ),
    .Q(_00252_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Halt_FF$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net422),
    .D(_00361_),
    .Q_N(_00035_),
    .Q(\z80.tv80s.i_tv80_core.Halt_FF ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.INT_s$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net422),
    .D(_00362_),
    .Q_N(_05655_),
    .Q(\z80.tv80s.i_tv80_core.INT_s ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IR[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net432),
    .D(_00363_),
    .Q_N(_00215_),
    .Q(\z80.tv80s.i_tv80_core.IR[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IR[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net432),
    .D(_00364_),
    .Q_N(_00027_),
    .Q(\z80.tv80s.i_tv80_core.IR[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IR[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net432),
    .D(_00365_),
    .Q_N(_00025_),
    .Q(\z80.tv80s.i_tv80_core.IR[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IR[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net432),
    .D(_00366_),
    .Q_N(_00033_),
    .Q(\z80.tv80s.i_tv80_core.IR[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IR[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net432),
    .D(_00367_),
    .Q_N(_00029_),
    .Q(\z80.tv80s.i_tv80_core.IR[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IR[5]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net432),
    .D(_00368_),
    .Q_N(_00021_),
    .Q(\z80.tv80s.i_tv80_core.IR[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IR[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net432),
    .D(_00369_),
    .Q_N(_05654_),
    .Q(\z80.tv80s.i_tv80_core.IR[6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IR[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net433),
    .D(_00370_),
    .Q_N(_00216_),
    .Q(\z80.tv80s.i_tv80_core.IR[7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ISet[0]$_DFF_PN1_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net429),
    .D(_00277_),
    .Q_N(\z80.tv80s.i_tv80_core.ISet[0] ),
    .Q(_05692_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ISet[1]$_DFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net429),
    .D(_00000_),
    .Q_N(_05680_),
    .Q(\z80.tv80s.i_tv80_core.ISet[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ISet[2]$_DFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net429),
    .D(_00001_),
    .Q_N(_00034_),
    .Q(\z80.tv80s.i_tv80_core.ISet[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.ISet[3]$_DFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net429),
    .D(_00002_),
    .Q_N(_05681_),
    .Q(\z80.tv80s.i_tv80_core.ISet[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IStatus[1]$_DFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net427),
    .D(_00003_),
    .Q_N(_05682_),
    .Q(\z80.tv80s.i_tv80_core.IStatus[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IStatus[2]$_DFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net427),
    .D(_00004_),
    .Q_N(_05653_),
    .Q(\z80.tv80s.i_tv80_core.IStatus[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.I[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net404),
    .D(_00371_),
    .Q_N(_05652_),
    .Q(\z80.tv80s.i_tv80_core.I[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.I[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net417),
    .D(_00372_),
    .Q_N(_05651_),
    .Q(\z80.tv80s.i_tv80_core.I[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.I[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net406),
    .D(_00373_),
    .Q_N(_05650_),
    .Q(\z80.tv80s.i_tv80_core.I[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.I[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net405),
    .D(_00374_),
    .Q_N(_05649_),
    .Q(\z80.tv80s.i_tv80_core.I[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.I[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net404),
    .D(_00375_),
    .Q_N(_05648_),
    .Q(\z80.tv80s.i_tv80_core.I[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.I[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net405),
    .D(_00376_),
    .Q_N(_05647_),
    .Q(\z80.tv80s.i_tv80_core.I[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.I[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net405),
    .D(_00377_),
    .Q_N(_05646_),
    .Q(\z80.tv80s.i_tv80_core.I[6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.I[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net404),
    .D(_00378_),
    .Q_N(_05645_),
    .Q(\z80.tv80s.i_tv80_core.I[7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IncDecZ$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net452),
    .D(_00379_),
    .Q_N(_05644_),
    .Q(\z80.tv80s.i_tv80_core.IncDecZ ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IntCycle$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net428),
    .D(_00380_),
    .Q_N(_00026_),
    .Q(\z80.tv80s.i_tv80_core.IntCycle ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IntE_FF1$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net427),
    .D(_00381_),
    .Q_N(_05643_),
    .Q(\z80.tv80s.i_tv80_core.IntE ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.IntE_FF2$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net427),
    .D(_00382_),
    .Q_N(_00136_),
    .Q(\z80.tv80s.i_tv80_core.IntE_FF2 ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.NMICycle$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net427),
    .D(_00383_),
    .Q_N(_00016_),
    .Q(\z80.tv80s.i_tv80_core.NMICycle ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.NMI_s$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net427),
    .D(_00384_),
    .Q_N(_05642_),
    .Q(\z80.tv80s.i_tv80_core.NMI_s ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.No_BTR$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net429),
    .D(_00385_),
    .Q_N(_05641_),
    .Q(\z80.tv80s.i_tv80_core.No_BTR ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Oldnmi_n$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net421),
    .D(_00386_),
    .Q_N(_05640_),
    .Q(\z80.tv80s.i_tv80_core.Oldnmi_n ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net406),
    .D(_00387_),
    .Q_N(_05639_),
    .Q(\z80.tv80s.i_tv80_core.PC[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net400),
    .D(_00388_),
    .Q_N(_00145_),
    .Q(\z80.tv80s.i_tv80_core.PC[10] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net400),
    .D(_00389_),
    .Q_N(_00148_),
    .Q(\z80.tv80s.i_tv80_core.PC[11] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net400),
    .D(_00390_),
    .Q_N(_00151_),
    .Q(\z80.tv80s.i_tv80_core.PC[12] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net400),
    .D(_00391_),
    .Q_N(_00154_),
    .Q(\z80.tv80s.i_tv80_core.PC[13] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net400),
    .D(_00392_),
    .Q_N(_00157_),
    .Q(\z80.tv80s.i_tv80_core.PC[14] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net400),
    .D(_00393_),
    .Q_N(_00160_),
    .Q(\z80.tv80s.i_tv80_core.PC[15] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net408),
    .D(_00394_),
    .Q_N(_00170_),
    .Q(\z80.tv80s.i_tv80_core.PC[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net406),
    .D(_00395_),
    .Q_N(_00180_),
    .Q(\z80.tv80s.i_tv80_core.PC[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net404),
    .D(_00396_),
    .Q_N(_00182_),
    .Q(\z80.tv80s.i_tv80_core.PC[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net404),
    .D(_00397_),
    .Q_N(_00184_),
    .Q(\z80.tv80s.i_tv80_core.PC[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net408),
    .D(_00398_),
    .Q_N(_00186_),
    .Q(\z80.tv80s.i_tv80_core.PC[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net408),
    .D(_00399_),
    .Q_N(_00188_),
    .Q(\z80.tv80s.i_tv80_core.PC[6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net408),
    .D(_00400_),
    .Q_N(_00190_),
    .Q(\z80.tv80s.i_tv80_core.PC[7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net408),
    .D(_00401_),
    .Q_N(_00139_),
    .Q(\z80.tv80s.i_tv80_core.PC[8] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PC[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net408),
    .D(_00402_),
    .Q_N(_00142_),
    .Q(\z80.tv80s.i_tv80_core.PC[9] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Pre_XY_F_M[1]$_DFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net430),
    .D(_00005_),
    .Q_N(_05683_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Pre_XY_F_M[2]$_DFF_PN0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net428),
    .D(_00006_),
    .Q_N(_05684_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Pre_XY_F_M[3]$_DFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net430),
    .D(_00007_),
    .Q_N(_05685_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Pre_XY_F_M[4]$_DFF_PN0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net428),
    .D(_00008_),
    .Q_N(_05686_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Pre_XY_F_M[5]$_DFF_PN0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net428),
    .D(_00009_),
    .Q_N(_05687_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Pre_XY_F_M[6]$_DFF_PN0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net427),
    .D(_00010_),
    .Q_N(_05688_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Pre_XY_F_M[7]$_DFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net430),
    .D(_00011_),
    .Q_N(_05638_),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.PreserveC_r$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net426),
    .D(_00403_),
    .Q_N(_05637_),
    .Q(\z80.tv80s.i_tv80_core.PreserveC_r ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.R[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net416),
    .D(_00404_),
    .Q_N(_05636_),
    .Q(\z80.tv80s.i_tv80_core.R[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.R[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net417),
    .D(_00405_),
    .Q_N(_05635_),
    .Q(\z80.tv80s.i_tv80_core.R[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.R[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net407),
    .D(_00406_),
    .Q_N(_05634_),
    .Q(\z80.tv80s.i_tv80_core.R[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.R[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net410),
    .D(_00407_),
    .Q_N(_05633_),
    .Q(\z80.tv80s.i_tv80_core.R[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.R[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net410),
    .D(_00408_),
    .Q_N(_05632_),
    .Q(\z80.tv80s.i_tv80_core.R[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.R[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net409),
    .D(_00409_),
    .Q_N(_05631_),
    .Q(\z80.tv80s.i_tv80_core.R[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.R[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net409),
    .D(_00410_),
    .Q_N(_05630_),
    .Q(\z80.tv80s.i_tv80_core.R[6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.R[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net416),
    .D(_00411_),
    .Q_N(_05629_),
    .Q(\z80.tv80s.i_tv80_core.R[7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Read_To_Reg_r[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net414),
    .D(_00412_),
    .Q_N(_05628_),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Read_To_Reg_r[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net425),
    .D(_00413_),
    .Q_N(_05627_),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Read_To_Reg_r[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net425),
    .D(_00414_),
    .Q_N(_05626_),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Read_To_Reg_r[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net414),
    .D(_00415_),
    .Q_N(_05625_),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Read_To_Reg_r[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net425),
    .D(_00416_),
    .Q_N(_00210_),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegAddrA_r[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net453),
    .D(_00417_),
    .Q_N(_05624_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegAddrA_r[1]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net454),
    .D(_00418_),
    .Q_N(_05623_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegAddrA_r[2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net455),
    .D(_00419_),
    .Q_N(_00038_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegAddrB_r[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net456),
    .D(_00420_),
    .Q_N(_05622_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegAddrB_r[1]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net457),
    .D(_00421_),
    .Q_N(_05621_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegAddrB_r[2]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net458),
    .D(_00422_),
    .Q_N(_00213_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegAddrC[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net459),
    .D(_00423_),
    .Q_N(_05620_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegAddrC[1]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net460),
    .D(_00424_),
    .Q_N(_05619_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegAddrC[2]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net461),
    .D(_00425_),
    .Q_N(_05618_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[0]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net462),
    .D(_00426_),
    .Q_N(_05617_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[10]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net463),
    .D(_00427_),
    .Q_N(_05616_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[10] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[11]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net464),
    .D(_00428_),
    .Q_N(_05615_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[11] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[12]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net465),
    .D(_00429_),
    .Q_N(_05614_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[12] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[13]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net466),
    .D(_00430_),
    .Q_N(_05613_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[13] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[14]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net467),
    .D(_00431_),
    .Q_N(_05612_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[14] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[15]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net468),
    .D(_00432_),
    .Q_N(_05611_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[15] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[1]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net469),
    .D(_00433_),
    .Q_N(_05610_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net470),
    .D(_00434_),
    .Q_N(_05609_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[3]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net471),
    .D(_00435_),
    .Q_N(_05608_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[4]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net472),
    .D(_00436_),
    .Q_N(_05607_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net473),
    .D(_00437_),
    .Q_N(_05606_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[6]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net474),
    .D(_00438_),
    .Q_N(_05605_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[7]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net475),
    .D(_00439_),
    .Q_N(_05604_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[8]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net476),
    .D(_00440_),
    .Q_N(_05603_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[8] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.RegBusA_r[9]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net477),
    .D(_00441_),
    .Q_N(_05602_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[9] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net402),
    .D(_00442_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[0] ),
    .Q(_00253_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[10]$_DFFE_PN1P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net412),
    .D(_00443_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[10] ),
    .Q(_00254_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[11]$_DFFE_PN1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net402),
    .D(_00444_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[11] ),
    .Q(_00255_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[12]$_DFFE_PN1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net402),
    .D(_00445_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[12] ),
    .Q(_00256_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[13]$_DFFE_PN1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net401),
    .D(_00446_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[13] ),
    .Q(_00257_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[14]$_DFFE_PN1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net402),
    .D(_00447_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[14] ),
    .Q(_00258_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[15]$_DFFE_PN1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net401),
    .D(_00448_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[15] ),
    .Q(_00259_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net402),
    .D(_00449_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[1] ),
    .Q(_00260_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net402),
    .D(_00450_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[2] ),
    .Q(_00261_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net412),
    .D(_00451_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[3] ),
    .Q(_00262_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[4]$_DFFE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net412),
    .D(_00452_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[4] ),
    .Q(_00263_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[5]$_DFFE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net412),
    .D(_00453_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[5] ),
    .Q(_00264_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[6]$_DFFE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net412),
    .D(_00454_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[6] ),
    .Q(_00265_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[7]$_DFFE_PN1P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net402),
    .D(_00455_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[7] ),
    .Q(_00266_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[8]$_DFFE_PN1P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net402),
    .D(_00456_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[8] ),
    .Q(_00267_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.SP[9]$_DFFE_PN1P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net403),
    .D(_00457_),
    .Q_N(\z80.tv80s.i_tv80_core.SP[9] ),
    .Q(_00268_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Save_ALU_r$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net426),
    .D(_00458_),
    .Q_N(_00191_),
    .Q(\z80.tv80s.i_tv80_core.Save_ALU_r ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net418),
    .D(_00459_),
    .Q_N(_05601_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net403),
    .D(_00460_),
    .Q_N(_00144_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[10] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net403),
    .D(_00461_),
    .Q_N(_00147_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[11] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net400),
    .D(_00462_),
    .Q_N(_00150_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[12] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net401),
    .D(_00463_),
    .Q_N(_00153_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[13] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net400),
    .D(_00464_),
    .Q_N(_00156_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[14] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net401),
    .D(_00465_),
    .Q_N(_00159_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[15] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net418),
    .D(_00466_),
    .Q_N(_00169_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net418),
    .D(_00467_),
    .Q_N(_00179_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net418),
    .D(_00468_),
    .Q_N(_00181_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net419),
    .D(_00469_),
    .Q_N(_00183_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net418),
    .D(_00470_),
    .Q_N(_00185_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net418),
    .D(_00471_),
    .Q_N(_00187_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net418),
    .D(_00472_),
    .Q_N(_00189_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net403),
    .D(_00473_),
    .Q_N(_00138_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[8] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.TmpAddr[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net403),
    .D(_00474_),
    .Q_N(_00141_),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[9] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.XY_Ind$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net406),
    .D(_00475_),
    .Q_N(_05600_),
    .Q(\z80.tv80s.i_tv80_core.XY_Ind ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.XY_State[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net424),
    .D(_00476_),
    .Q_N(_05599_),
    .Q(\z80.tv80s.i_tv80_core.XY_State[0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.XY_State[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net425),
    .D(_00477_),
    .Q_N(_00037_),
    .Q(\z80.tv80s.i_tv80_core.XY_State[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.Z16_r$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net426),
    .D(_00478_),
    .Q_N(_05598_),
    .Q(\z80.tv80s.i_tv80_core.Z16_r ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.dout[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net410),
    .D(_00479_),
    .Q_N(_05597_),
    .Q(net22));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.dout[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net410),
    .D(_00480_),
    .Q_N(_05596_),
    .Q(net23));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.dout[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net410),
    .D(_00481_),
    .Q_N(_05595_),
    .Q(net24));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.dout[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net409),
    .D(_00482_),
    .Q_N(_05594_),
    .Q(net25));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.dout[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net409),
    .D(_00483_),
    .Q_N(_05593_),
    .Q(net26));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.dout[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net409),
    .D(_00484_),
    .Q_N(_05592_),
    .Q(net27));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.dout[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net409),
    .D(_00485_),
    .Q_N(_05591_),
    .Q(net28));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.dout[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net405),
    .D(_00486_),
    .Q_N(_05590_),
    .Q(net29));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net478),
    .D(_00487_),
    .Q_N(_05589_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net479),
    .D(_00488_),
    .Q_N(_00039_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net480),
    .D(_00489_),
    .Q_N(_00047_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net481),
    .D(_00490_),
    .Q_N(_00055_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net482),
    .D(_00491_),
    .Q_N(_00063_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net483),
    .D(_00492_),
    .Q_N(_00071_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net484),
    .D(_00493_),
    .Q_N(_00079_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net485),
    .D(_00494_),
    .Q_N(_00087_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net486),
    .D(_00495_),
    .Q_N(_05588_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net487),
    .D(_00496_),
    .Q_N(_00040_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net488),
    .D(_00497_),
    .Q_N(_00048_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net489),
    .D(_00498_),
    .Q_N(_00056_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net490),
    .D(_00499_),
    .Q_N(_00064_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net491),
    .D(_00500_),
    .Q_N(_00072_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net492),
    .D(_00501_),
    .Q_N(_00080_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net493),
    .D(_00502_),
    .Q_N(_00088_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net494),
    .D(_00503_),
    .Q_N(_05587_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net495),
    .D(_00504_),
    .Q_N(_00041_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net496),
    .D(_00505_),
    .Q_N(_00049_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net497),
    .D(_00506_),
    .Q_N(_00057_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net498),
    .D(_00507_),
    .Q_N(_00065_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net499),
    .D(_00508_),
    .Q_N(_00073_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net500),
    .D(_00509_),
    .Q_N(_00081_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net501),
    .D(_00510_),
    .Q_N(_00089_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net502),
    .D(_00511_),
    .Q_N(_05586_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net503),
    .D(_00512_),
    .Q_N(_00042_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net504),
    .D(_00513_),
    .Q_N(_00050_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net505),
    .D(_00514_),
    .Q_N(_00058_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net506),
    .D(_00515_),
    .Q_N(_00066_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net507),
    .D(_00516_),
    .Q_N(_00074_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net508),
    .D(_00517_),
    .Q_N(_00082_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net509),
    .D(_00518_),
    .Q_N(_00090_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net510),
    .D(_00519_),
    .Q_N(_05585_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net511),
    .D(_00520_),
    .Q_N(_00043_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net512),
    .D(_00521_),
    .Q_N(_00051_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net513),
    .D(_00522_),
    .Q_N(_00059_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net514),
    .D(_00523_),
    .Q_N(_00067_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net515),
    .D(_00524_),
    .Q_N(_00075_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net516),
    .D(_00525_),
    .Q_N(_00083_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net517),
    .D(_00526_),
    .Q_N(_00091_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net518),
    .D(_00527_),
    .Q_N(_05584_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net519),
    .D(_00528_),
    .Q_N(_00044_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net520),
    .D(_00529_),
    .Q_N(_00052_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net521),
    .D(_00530_),
    .Q_N(_00060_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net522),
    .D(_00531_),
    .Q_N(_00068_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net523),
    .D(_00532_),
    .Q_N(_00076_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net524),
    .D(_00533_),
    .Q_N(_00084_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net525),
    .D(_00534_),
    .Q_N(_00092_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net526),
    .D(_00535_),
    .Q_N(_05583_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net527),
    .D(_00536_),
    .Q_N(_00045_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net528),
    .D(_00537_),
    .Q_N(_00053_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net529),
    .D(_00538_),
    .Q_N(_00061_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net530),
    .D(_00539_),
    .Q_N(_00069_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net531),
    .D(_00540_),
    .Q_N(_00077_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net532),
    .D(_00541_),
    .Q_N(_00085_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net533),
    .D(_00542_),
    .Q_N(_00093_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net534),
    .D(_00543_),
    .Q_N(_05582_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net535),
    .D(_00544_),
    .Q_N(_00046_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net536),
    .D(_00545_),
    .Q_N(_00054_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net537),
    .D(_00546_),
    .Q_N(_00062_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net538),
    .D(_00547_),
    .Q_N(_00070_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net539),
    .D(_00548_),
    .Q_N(_00078_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net540),
    .D(_00549_),
    .Q_N(_00086_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsH[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net541),
    .D(_00550_),
    .Q_N(_00094_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net542),
    .D(_00551_),
    .Q_N(_05581_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net543),
    .D(_00552_),
    .Q_N(_00161_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net544),
    .D(_00553_),
    .Q_N(_00171_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net545),
    .D(_00554_),
    .Q_N(_00095_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net546),
    .D(_00555_),
    .Q_N(_00103_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net547),
    .D(_00556_),
    .Q_N(_00111_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net548),
    .D(_00557_),
    .Q_N(_00119_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net549),
    .D(_00558_),
    .Q_N(_00127_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net550),
    .D(_00559_),
    .Q_N(_05580_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net551),
    .D(_00560_),
    .Q_N(_00162_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net552),
    .D(_00561_),
    .Q_N(_00172_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net553),
    .D(_00562_),
    .Q_N(_00096_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net554),
    .D(_00563_),
    .Q_N(_00104_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net555),
    .D(_00564_),
    .Q_N(_00112_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net556),
    .D(_00565_),
    .Q_N(_00120_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net557),
    .D(_00566_),
    .Q_N(_00128_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net558),
    .D(_00567_),
    .Q_N(_05579_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net559),
    .D(_00568_),
    .Q_N(_00163_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net560),
    .D(_00569_),
    .Q_N(_00173_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net561),
    .D(_00570_),
    .Q_N(_00097_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net562),
    .D(_00571_),
    .Q_N(_00105_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net563),
    .D(_00572_),
    .Q_N(_00113_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net564),
    .D(_00573_),
    .Q_N(_00121_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net565),
    .D(_00574_),
    .Q_N(_00129_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net566),
    .D(_00575_),
    .Q_N(_05578_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net567),
    .D(_00576_),
    .Q_N(_00164_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[3][2]$_DFFE_PP_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net568),
    .D(_00577_),
    .Q_N(_00174_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net569),
    .D(_00578_),
    .Q_N(_00098_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net570),
    .D(_00579_),
    .Q_N(_00106_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net571),
    .D(_00580_),
    .Q_N(_00114_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net572),
    .D(_00581_),
    .Q_N(_00122_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net573),
    .D(_00582_),
    .Q_N(_00130_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net574),
    .D(_00583_),
    .Q_N(_05577_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net575),
    .D(_00584_),
    .Q_N(_00165_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net576),
    .D(_00585_),
    .Q_N(_00175_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net577),
    .D(_00586_),
    .Q_N(_00099_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net578),
    .D(_00587_),
    .Q_N(_00107_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net579),
    .D(_00588_),
    .Q_N(_00115_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net580),
    .D(_00589_),
    .Q_N(_00123_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net581),
    .D(_00590_),
    .Q_N(_00131_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net582),
    .D(_00591_),
    .Q_N(_05576_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net583),
    .D(_00592_),
    .Q_N(_00166_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net584),
    .D(_00593_),
    .Q_N(_00176_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net585),
    .D(_00594_),
    .Q_N(_00100_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net586),
    .D(_00595_),
    .Q_N(_00108_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net587),
    .D(_00596_),
    .Q_N(_00116_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net588),
    .D(_00597_),
    .Q_N(_00124_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net589),
    .D(_00598_),
    .Q_N(_00132_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net590),
    .D(_00599_),
    .Q_N(_05575_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net591),
    .D(_00600_),
    .Q_N(_00167_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net592),
    .D(_00601_),
    .Q_N(_00177_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net593),
    .D(_00602_),
    .Q_N(_00101_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net594),
    .D(_00603_),
    .Q_N(_00109_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net595),
    .D(_00604_),
    .Q_N(_00117_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net596),
    .D(_00605_),
    .Q_N(_00125_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net597),
    .D(_00606_),
    .Q_N(_00133_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net598),
    .D(_00607_),
    .Q_N(_05574_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net599),
    .D(_00608_),
    .Q_N(_00168_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net600),
    .D(_00609_),
    .Q_N(_00178_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net601),
    .D(_00610_),
    .Q_N(_00102_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net602),
    .D(_00611_),
    .Q_N(_00110_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net603),
    .D(_00612_),
    .Q_N(_00118_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net604),
    .D(_00613_),
    .Q_N(_00126_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.i_reg.RegsL[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net605),
    .D(_00614_),
    .Q_N(_00134_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.m1_n$_DFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net422),
    .D(_00615_),
    .Q_N(\z80.m1_n ),
    .Q(_00269_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.mcycle[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net431),
    .D(_00616_),
    .Q_N(\z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ),
    .Q(_00270_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.mcycle[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net432),
    .D(_00617_),
    .Q_N(_00217_),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.mcycle[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net431),
    .D(_00618_),
    .Q_N(_00022_),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.mcycle[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net431),
    .D(_00619_),
    .Q_N(_00023_),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.mcycle[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net430),
    .D(_00620_),
    .Q_N(_00028_),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.mcycle[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net428),
    .D(_00621_),
    .Q_N(_00214_),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.mcycle[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net430),
    .D(_00622_),
    .Q_N(_00212_),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.mcycles[1]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net424),
    .D(_00012_),
    .Q_N(_05689_),
    .Q(\z80.tv80s.i_tv80_core.mcycles[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.mcycles[2]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net426),
    .D(_00013_),
    .Q_N(_05690_),
    .Q(\z80.tv80s.i_tv80_core.mcycles[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.mcycles[4]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net429),
    .D(_00014_),
    .Q_N(_05691_),
    .Q(\z80.tv80s.i_tv80_core.mcycles[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.mcycles[5]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net426),
    .D(_00015_),
    .Q_N(_05573_),
    .Q(\z80.tv80s.i_tv80_core.mcycles[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.rfsh_n$_DFFE_PN1P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net416),
    .D(_00623_),
    .Q_N(\z80.rfsh_n ),
    .Q(_00271_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.tstate[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net421),
    .D(_00624_),
    .Q_N(\z80.tv80s.i_tv80_core.ts[0] ),
    .Q(_00272_));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.tstate[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net422),
    .D(_00625_),
    .Q_N(_00135_),
    .Q(\z80.tv80s.i_tv80_core.ts[1] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.tstate[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net427),
    .D(_00626_),
    .Q_N(_00032_),
    .Q(\z80.tv80s.i_tv80_core.ts[2] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.tstate[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net421),
    .D(_00627_),
    .Q_N(_00024_),
    .Q(\z80.tv80s.i_tv80_core.ts[3] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.tstate[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net416),
    .D(_00628_),
    .Q_N(_05572_),
    .Q(\z80.tv80s.i_tv80_core.ts[4] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.tstate[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net421),
    .D(_00629_),
    .Q_N(_05571_),
    .Q(\z80.tv80s.i_tv80_core.ts[5] ));
 sg13g2_dfrbp_1 \z80.tv80s.i_tv80_core.tstate[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net421),
    .D(_00630_),
    .Q_N(_00030_),
    .Q(\z80.tv80s.i_tv80_core.ts[6] ));
 sg13g2_dfrbp_1 \z80.tv80s.iorq_n$_DFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net422),
    .D(_00631_),
    .Q_N(\z80.iorq_n ),
    .Q(_00273_));
 sg13g2_dfrbp_1 \z80.tv80s.mreq_n$_DFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net417),
    .D(_00632_),
    .Q_N(\z80.mreq_n ),
    .Q(_00274_));
 sg13g2_dfrbp_1 \z80.tv80s.rd_n$_DFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net422),
    .D(_00633_),
    .Q_N(\z80.rd_n ),
    .Q(_00275_));
 sg13g2_dfrbp_1 \z80.tv80s.wr_n$_DFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net417),
    .D(_00634_),
    .Q_N(\z80.tv80s.wr_n ),
    .Q(_00276_));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[5]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[6]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_oe[0]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[1]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_oe[2]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_oe[3]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_oe[4]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_oe[5]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_oe[6]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_oe[7]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[0]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[1]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[2]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uio_out[3]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uio_out[4]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uio_out[5]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uio_out[6]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uio_out[7]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[0]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[1]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uo_out[2]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(uo_out[3]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(uo_out[4]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(uo_out[5]));
 sg13g2_buf_1 output36 (.A(net36),
    .X(uo_out[6]));
 sg13g2_buf_1 output37 (.A(net37),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout38 (.A(_05289_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_05278_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_04770_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_03333_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_03248_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_05449_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_05443_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_05437_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_05429_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_05423_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_05416_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_05354_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_05301_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_05266_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_03199_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_05311_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_04283_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_03270_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_05505_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_05455_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_01208_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_03327_),
    .X(net59));
 sg13g2_buf_4 fanout60 (.X(net60),
    .A(_03068_));
 sg13g2_buf_2 fanout61 (.A(_04232_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_03277_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_03226_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_03186_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_03124_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_03113_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_03092_),
    .X(net67));
 sg13g2_buf_4 fanout68 (.X(net68),
    .A(_03067_));
 sg13g2_buf_2 fanout69 (.A(_02551_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_02389_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_02245_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_01206_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_05463_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_05181_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_04683_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_04270_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_03569_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_03502_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_03271_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_03194_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_03185_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_03153_),
    .X(net82));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(_03112_));
 sg13g2_buf_2 fanout84 (.A(_02441_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_02375_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_05186_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_05180_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_04284_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_04275_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_03560_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_03557_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_03496_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_03466_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_03007_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_02444_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_02417_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_02407_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_02393_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_02288_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_02089_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_04690_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_04644_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_04357_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_03752_),
    .X(net104));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(_03535_));
 sg13g2_buf_2 fanout106 (.A(_03499_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_03006_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_02998_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_02484_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_02436_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_02392_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_02336_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_02332_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_02291_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_02088_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_05239_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_04157_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_03758_),
    .X(net118));
 sg13g2_buf_8 fanout119 (.A(_03534_),
    .X(net119));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(_03526_));
 sg13g2_buf_8 fanout121 (.A(_03521_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_02861_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_02856_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_02855_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_02477_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_02394_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_02378_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_02308_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_01600_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_01576_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_05199_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_04971_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_04024_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_03530_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_03516_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_02383_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_02307_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_02293_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_01695_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_05200_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_04041_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_03548_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_03515_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_03038_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_02292_),
    .X(net145));
 sg13g2_buf_1 fanout146 (.A(doe),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_01137_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_05236_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_01973_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_04557_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_01567_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_01544_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_05100_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_04551_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_01543_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_05101_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_05099_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_02247_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_02246_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_01608_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_01539_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_04678_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_03983_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_02609_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_02450_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_02204_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_02101_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_01951_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_01603_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_00880_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_00865_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_04669_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_04657_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_02590_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_02133_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_02048_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_01960_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_01595_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_01341_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_01286_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_01277_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_01119_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_00973_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_00935_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_00920_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_04671_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_04659_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_04556_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_03850_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_03692_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_03217_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_02492_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_02456_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_02087_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_01896_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_01747_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_01615_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_01340_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_01330_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_01290_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_01285_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_01267_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_01141_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_01111_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_01047_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_01017_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_00896_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_00719_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_00712_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_00701_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_04590_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_04549_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_02345_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_02144_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_02128_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_01614_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_01491_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_01461_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_01388_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_01332_),
    .X(net220));
 sg13g2_buf_4 fanout221 (.X(net221),
    .A(_01314_));
 sg13g2_buf_2 fanout222 (.A(_01266_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_01259_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_01247_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_01246_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_01238_),
    .X(net226));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(_01237_));
 sg13g2_buf_2 fanout228 (.A(_01172_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_01123_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_01084_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_01064_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_01062_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_01042_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_01038_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_01016_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_00986_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_00984_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_00961_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_00914_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_00883_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_00824_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_00779_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_00749_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_00723_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_00649_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_04548_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_02496_),
    .X(net247));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(_02486_));
 sg13g2_buf_4 fanout249 (.X(net249),
    .A(_02485_));
 sg13g2_buf_2 fanout250 (.A(_02463_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_02408_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_02344_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_02324_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_02312_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_01879_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_01467_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_01331_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_01309_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_01295_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_01260_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_01253_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_01252_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_01245_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_01236_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_01231_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_01229_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_01101_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_01024_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_00977_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_00970_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_00951_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_00942_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_00916_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_00915_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_00875_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_00871_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_00829_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_00788_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_00773_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_00754_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_00752_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_00751_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_00739_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_00678_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_00668_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_00660_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_05094_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_04180_),
    .X(net288));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(_03524_));
 sg13g2_buf_2 fanout290 (.A(_02400_),
    .X(net290));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(_02398_));
 sg13g2_buf_2 fanout292 (.A(_02396_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_02313_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_01749_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_01540_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_01514_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_01502_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_01478_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_01476_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_01278_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_01230_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_01216_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_01045_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_01033_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_00968_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_00950_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_00931_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_00930_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_00924_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_00917_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_00882_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_00854_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_00747_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_00743_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_00742_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_00738_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_00721_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_00713_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_00710_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_00708_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_00669_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_00664_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_00643_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_00640_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_04179_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_03694_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_03523_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_02889_),
    .X(net328));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(_02399_));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(_02397_));
 sg13g2_buf_2 fanout331 (.A(_02395_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_02314_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_02241_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_02018_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_01994_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_01889_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_01843_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_01825_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_01788_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_01760_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_01696_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_01642_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_01512_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_01462_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_01458_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_01455_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_01451_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_01403_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_01401_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_01393_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_01161_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_01030_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_01014_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_01008_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_00967_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_00909_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_00891_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_00863_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_00860_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_00820_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_00715_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_00692_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_00686_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_00681_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_00653_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_00651_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_00645_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_00642_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_00639_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_05547_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_05545_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_02839_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_02802_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_01961_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_01948_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_01914_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_01850_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_01820_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_01803_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_01697_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_01493_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_01464_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_01457_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_01456_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_01399_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_01398_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_01397_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_01396_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_01395_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_01394_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_01254_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_00908_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_00905_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_00826_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_00704_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_00688_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_00684_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_00637_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_00636_),
    .X(net399));
 sg13g2_buf_4 fanout400 (.X(net400),
    .A(net401));
 sg13g2_buf_2 fanout401 (.A(net411),
    .X(net401));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(net403));
 sg13g2_buf_2 fanout403 (.A(net411),
    .X(net403));
 sg13g2_buf_4 fanout404 (.X(net404),
    .A(net407));
 sg13g2_buf_2 fanout405 (.A(net407),
    .X(net405));
 sg13g2_buf_4 fanout406 (.X(net406),
    .A(net407));
 sg13g2_buf_1 fanout407 (.A(net408),
    .X(net407));
 sg13g2_buf_4 fanout408 (.X(net408),
    .A(net411));
 sg13g2_buf_4 fanout409 (.X(net409),
    .A(net411));
 sg13g2_buf_4 fanout410 (.X(net410),
    .A(net411));
 sg13g2_buf_1 fanout411 (.A(net435),
    .X(net411));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(net415));
 sg13g2_buf_4 fanout413 (.X(net413),
    .A(net414));
 sg13g2_buf_4 fanout414 (.X(net414),
    .A(net415));
 sg13g2_buf_2 fanout415 (.A(net435),
    .X(net415));
 sg13g2_buf_4 fanout416 (.X(net416),
    .A(net417));
 sg13g2_buf_4 fanout417 (.X(net417),
    .A(net423));
 sg13g2_buf_4 fanout418 (.X(net418),
    .A(net423));
 sg13g2_buf_4 fanout419 (.X(net419),
    .A(net423));
 sg13g2_buf_2 fanout420 (.A(net423),
    .X(net420));
 sg13g2_buf_4 fanout421 (.X(net421),
    .A(net422));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(net423));
 sg13g2_buf_1 fanout423 (.A(net435),
    .X(net423));
 sg13g2_buf_4 fanout424 (.X(net424),
    .A(net426));
 sg13g2_buf_4 fanout425 (.X(net425),
    .A(net426));
 sg13g2_buf_4 fanout426 (.X(net426),
    .A(net434));
 sg13g2_buf_4 fanout427 (.X(net427),
    .A(net429));
 sg13g2_buf_2 fanout428 (.A(net429),
    .X(net428));
 sg13g2_buf_4 fanout429 (.X(net429),
    .A(net434));
 sg13g2_buf_4 fanout430 (.X(net430),
    .A(net431));
 sg13g2_buf_2 fanout431 (.A(net434),
    .X(net431));
 sg13g2_buf_4 fanout432 (.X(net432),
    .A(net433));
 sg13g2_buf_2 fanout433 (.A(net434),
    .X(net433));
 sg13g2_buf_1 fanout434 (.A(net435),
    .X(net434));
 sg13g2_buf_1 fanout435 (.A(net1),
    .X(net435));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusA[0]$_DFFE_PP__436  (.L_HI(net436));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusA[1]$_DFFE_PP__437  (.L_HI(net437));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusA[2]$_DFFE_PP__438  (.L_HI(net438));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusA[3]$_DFFE_PP__439  (.L_HI(net439));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusA[4]$_DFFE_PP__440  (.L_HI(net440));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusA[5]$_DFFE_PP__441  (.L_HI(net441));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusA[6]$_DFFE_PP__442  (.L_HI(net442));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusA[7]$_DFFE_PP__443  (.L_HI(net443));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusB[0]$_DFFE_PP__444  (.L_HI(net444));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusB[1]$_DFFE_PP__445  (.L_HI(net445));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusB[2]$_DFFE_PP__446  (.L_HI(net446));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusB[3]$_DFFE_PP__447  (.L_HI(net447));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusB[4]$_DFFE_PP__448  (.L_HI(net448));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusB[5]$_DFFE_PP__449  (.L_HI(net449));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusB[6]$_DFFE_PP__450  (.L_HI(net450));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.BusB[7]$_DFFE_PP__451  (.L_HI(net451));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.IncDecZ$_DFFE_PP__452  (.L_HI(net452));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegAddrA_r[0]$_SDFFCE_PP1P__453  (.L_HI(net453));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegAddrA_r[1]$_SDFFCE_PP1P__454  (.L_HI(net454));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegAddrA_r[2]$_DFFE_PP__455  (.L_HI(net455));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegAddrB_r[0]$_SDFFCE_PP1P__456  (.L_HI(net456));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegAddrB_r[1]$_SDFFCE_PP1P__457  (.L_HI(net457));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegAddrB_r[2]$_DFFE_PP__458  (.L_HI(net458));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegAddrC[0]$_SDFFCE_PP1P__459  (.L_HI(net459));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegAddrC[1]$_SDFFCE_PP1P__460  (.L_HI(net460));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegAddrC[2]$_DFFE_PP__461  (.L_HI(net461));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[0]$_DFFE_PP__462  (.L_HI(net462));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[10]$_DFFE_PP__463  (.L_HI(net463));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[11]$_DFFE_PP__464  (.L_HI(net464));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[12]$_DFFE_PP__465  (.L_HI(net465));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[13]$_DFFE_PP__466  (.L_HI(net466));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[14]$_DFFE_PP__467  (.L_HI(net467));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[15]$_DFFE_PP__468  (.L_HI(net468));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[1]$_DFFE_PP__469  (.L_HI(net469));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[2]$_DFFE_PP__470  (.L_HI(net470));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[3]$_DFFE_PP__471  (.L_HI(net471));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[4]$_DFFE_PP__472  (.L_HI(net472));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[5]$_DFFE_PP__473  (.L_HI(net473));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[6]$_DFFE_PP__474  (.L_HI(net474));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[7]$_DFFE_PP__475  (.L_HI(net475));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[8]$_DFFE_PP__476  (.L_HI(net476));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.RegBusA_r[9]$_DFFE_PP__477  (.L_HI(net477));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[0][0]$_DFFE_PP__478  (.L_HI(net478));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[0][1]$_DFFE_PP__479  (.L_HI(net479));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[0][2]$_DFFE_PP__480  (.L_HI(net480));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[0][3]$_DFFE_PP__481  (.L_HI(net481));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[0][4]$_DFFE_PP__482  (.L_HI(net482));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[0][5]$_DFFE_PP__483  (.L_HI(net483));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[0][6]$_DFFE_PP__484  (.L_HI(net484));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[0][7]$_DFFE_PP__485  (.L_HI(net485));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[1][0]$_DFFE_PP__486  (.L_HI(net486));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[1][1]$_DFFE_PP__487  (.L_HI(net487));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[1][2]$_DFFE_PP__488  (.L_HI(net488));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[1][3]$_DFFE_PP__489  (.L_HI(net489));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[1][4]$_DFFE_PP__490  (.L_HI(net490));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[1][5]$_DFFE_PP__491  (.L_HI(net491));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[1][6]$_DFFE_PP__492  (.L_HI(net492));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[1][7]$_DFFE_PP__493  (.L_HI(net493));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[2][0]$_DFFE_PP__494  (.L_HI(net494));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[2][1]$_DFFE_PP__495  (.L_HI(net495));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[2][2]$_DFFE_PP__496  (.L_HI(net496));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[2][3]$_DFFE_PP__497  (.L_HI(net497));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[2][4]$_DFFE_PP__498  (.L_HI(net498));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[2][5]$_DFFE_PP__499  (.L_HI(net499));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[2][6]$_DFFE_PP__500  (.L_HI(net500));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[2][7]$_DFFE_PP__501  (.L_HI(net501));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[3][0]$_DFFE_PP__502  (.L_HI(net502));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[3][1]$_DFFE_PP__503  (.L_HI(net503));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[3][2]$_DFFE_PP__504  (.L_HI(net504));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[3][3]$_DFFE_PP__505  (.L_HI(net505));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[3][4]$_DFFE_PP__506  (.L_HI(net506));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[3][5]$_DFFE_PP__507  (.L_HI(net507));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[3][6]$_DFFE_PP__508  (.L_HI(net508));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[3][7]$_DFFE_PP__509  (.L_HI(net509));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[4][0]$_DFFE_PP__510  (.L_HI(net510));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[4][1]$_DFFE_PP__511  (.L_HI(net511));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[4][2]$_DFFE_PP__512  (.L_HI(net512));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[4][3]$_DFFE_PP__513  (.L_HI(net513));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[4][4]$_DFFE_PP__514  (.L_HI(net514));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[4][5]$_DFFE_PP__515  (.L_HI(net515));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[4][6]$_DFFE_PP__516  (.L_HI(net516));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[4][7]$_DFFE_PP__517  (.L_HI(net517));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[5][0]$_DFFE_PP__518  (.L_HI(net518));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[5][1]$_DFFE_PP__519  (.L_HI(net519));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[5][2]$_DFFE_PP__520  (.L_HI(net520));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[5][3]$_DFFE_PP__521  (.L_HI(net521));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[5][4]$_DFFE_PP__522  (.L_HI(net522));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[5][5]$_DFFE_PP__523  (.L_HI(net523));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[5][6]$_DFFE_PP__524  (.L_HI(net524));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[5][7]$_DFFE_PP__525  (.L_HI(net525));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[6][0]$_DFFE_PP__526  (.L_HI(net526));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[6][1]$_DFFE_PP__527  (.L_HI(net527));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[6][2]$_DFFE_PP__528  (.L_HI(net528));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[6][3]$_DFFE_PP__529  (.L_HI(net529));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[6][4]$_DFFE_PP__530  (.L_HI(net530));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[6][5]$_DFFE_PP__531  (.L_HI(net531));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[6][6]$_DFFE_PP__532  (.L_HI(net532));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[6][7]$_DFFE_PP__533  (.L_HI(net533));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[7][0]$_DFFE_PP__534  (.L_HI(net534));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[7][1]$_DFFE_PP__535  (.L_HI(net535));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[7][2]$_DFFE_PP__536  (.L_HI(net536));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[7][3]$_DFFE_PP__537  (.L_HI(net537));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[7][4]$_DFFE_PP__538  (.L_HI(net538));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[7][5]$_DFFE_PP__539  (.L_HI(net539));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[7][6]$_DFFE_PP__540  (.L_HI(net540));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsH[7][7]$_DFFE_PP__541  (.L_HI(net541));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[0][0]$_DFFE_PP__542  (.L_HI(net542));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[0][1]$_DFFE_PP__543  (.L_HI(net543));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[0][2]$_DFFE_PP__544  (.L_HI(net544));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[0][3]$_DFFE_PP__545  (.L_HI(net545));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[0][4]$_DFFE_PP__546  (.L_HI(net546));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[0][5]$_DFFE_PP__547  (.L_HI(net547));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[0][6]$_DFFE_PP__548  (.L_HI(net548));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[0][7]$_DFFE_PP__549  (.L_HI(net549));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[1][0]$_DFFE_PP__550  (.L_HI(net550));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[1][1]$_DFFE_PP__551  (.L_HI(net551));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[1][2]$_DFFE_PP__552  (.L_HI(net552));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[1][3]$_DFFE_PP__553  (.L_HI(net553));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[1][4]$_DFFE_PP__554  (.L_HI(net554));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[1][5]$_DFFE_PP__555  (.L_HI(net555));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[1][6]$_DFFE_PP__556  (.L_HI(net556));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[1][7]$_DFFE_PP__557  (.L_HI(net557));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[2][0]$_DFFE_PP__558  (.L_HI(net558));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[2][1]$_DFFE_PP__559  (.L_HI(net559));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[2][2]$_DFFE_PP__560  (.L_HI(net560));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[2][3]$_DFFE_PP__561  (.L_HI(net561));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[2][4]$_DFFE_PP__562  (.L_HI(net562));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[2][5]$_DFFE_PP__563  (.L_HI(net563));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[2][6]$_DFFE_PP__564  (.L_HI(net564));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[2][7]$_DFFE_PP__565  (.L_HI(net565));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[3][0]$_DFFE_PP__566  (.L_HI(net566));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[3][1]$_DFFE_PP__567  (.L_HI(net567));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[3][2]$_DFFE_PP__568  (.L_HI(net568));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[3][3]$_DFFE_PP__569  (.L_HI(net569));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[3][4]$_DFFE_PP__570  (.L_HI(net570));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[3][5]$_DFFE_PP__571  (.L_HI(net571));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[3][6]$_DFFE_PP__572  (.L_HI(net572));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[3][7]$_DFFE_PP__573  (.L_HI(net573));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[4][0]$_DFFE_PP__574  (.L_HI(net574));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[4][1]$_DFFE_PP__575  (.L_HI(net575));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[4][2]$_DFFE_PP__576  (.L_HI(net576));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[4][3]$_DFFE_PP__577  (.L_HI(net577));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[4][4]$_DFFE_PP__578  (.L_HI(net578));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[4][5]$_DFFE_PP__579  (.L_HI(net579));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[4][6]$_DFFE_PP__580  (.L_HI(net580));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[4][7]$_DFFE_PP__581  (.L_HI(net581));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[5][0]$_DFFE_PP__582  (.L_HI(net582));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[5][1]$_DFFE_PP__583  (.L_HI(net583));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[5][2]$_DFFE_PP__584  (.L_HI(net584));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[5][3]$_DFFE_PP__585  (.L_HI(net585));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[5][4]$_DFFE_PP__586  (.L_HI(net586));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[5][5]$_DFFE_PP__587  (.L_HI(net587));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[5][6]$_DFFE_PP__588  (.L_HI(net588));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[5][7]$_DFFE_PP__589  (.L_HI(net589));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[6][0]$_DFFE_PP__590  (.L_HI(net590));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[6][1]$_DFFE_PP__591  (.L_HI(net591));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[6][2]$_DFFE_PP__592  (.L_HI(net592));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[6][3]$_DFFE_PP__593  (.L_HI(net593));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[6][4]$_DFFE_PP__594  (.L_HI(net594));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[6][5]$_DFFE_PP__595  (.L_HI(net595));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[6][6]$_DFFE_PP__596  (.L_HI(net596));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[6][7]$_DFFE_PP__597  (.L_HI(net597));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[7][0]$_DFFE_PP__598  (.L_HI(net598));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[7][1]$_DFFE_PP__599  (.L_HI(net599));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[7][2]$_DFFE_PP__600  (.L_HI(net600));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[7][3]$_DFFE_PP__601  (.L_HI(net601));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[7][4]$_DFFE_PP__602  (.L_HI(net602));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[7][5]$_DFFE_PP__603  (.L_HI(net603));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[7][6]$_DFFE_PP__604  (.L_HI(net604));
 sg13g2_tiehi \z80.tv80s.i_tv80_core.i_reg.RegsL[7][7]$_DFFE_PP__605  (.L_HI(net605));
 sg13g2_buf_4 clkbuf_leaf_1_clk (.X(clknet_leaf_1_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_3_clk (.X(clknet_leaf_3_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_5_clk (.X(clknet_leaf_5_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_9_clk (.X(clknet_leaf_9_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_10_clk (.X(clknet_leaf_10_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_11_clk (.X(clknet_leaf_11_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_15_clk (.X(clknet_leaf_15_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_19_clk (.X(clknet_leaf_19_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_22_clk (.X(clknet_leaf_22_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_24_clk (.X(clknet_leaf_24_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_25_clk (.X(clknet_leaf_25_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_26_clk (.X(clknet_leaf_26_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_27_clk (.X(clknet_leaf_27_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_28_clk (.X(clknet_leaf_28_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_29_clk (.X(clknet_leaf_29_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_30_clk (.X(clknet_leaf_30_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_31_clk (.X(clknet_leaf_31_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_32_clk (.X(clknet_leaf_32_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_33_clk (.X(clknet_leaf_33_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_34_clk (.X(clknet_leaf_34_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_35_clk (.X(clknet_leaf_35_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_37_clk (.X(clknet_leaf_37_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_38_clk (.X(clknet_leaf_38_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_39_clk (.X(clknet_leaf_39_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_40_clk (.X(clknet_leaf_40_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_41_clk (.X(clknet_leaf_41_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_42_clk (.X(clknet_leaf_42_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_44_clk (.X(clknet_leaf_44_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_45_clk (.X(clknet_leaf_45_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_47_clk (.X(clknet_leaf_47_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_48_clk (.X(clknet_leaf_48_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_49_clk (.X(clknet_leaf_49_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_50_clk (.X(clknet_leaf_50_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_51_clk (.X(clknet_leaf_51_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_52_clk (.X(clknet_leaf_52_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_53_clk (.X(clknet_leaf_53_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_54_clk (.X(clknet_leaf_54_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_55_clk (.X(clknet_leaf_55_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_56_clk (.X(clknet_leaf_56_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_57_clk (.X(clknet_leaf_57_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_58_clk (.X(clknet_leaf_58_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkbuf_leaf_59_clk (.X(clknet_leaf_59_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_60_clk (.X(clknet_leaf_60_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkbuf_leaf_61_clk (.X(clknet_leaf_61_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_0_0_clk (.X(clknet_4_0_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_1_0_clk (.X(clknet_4_1_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_2_0_clk (.X(clknet_4_2_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_3_0_clk (.X(clknet_4_3_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_4_0_clk (.X(clknet_4_4_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_5_0_clk (.X(clknet_4_5_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_6_0_clk (.X(clknet_4_6_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_7_0_clk (.X(clknet_4_7_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_8_0_clk (.X(clknet_4_8_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_9_0_clk (.X(clknet_4_9_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_10_0_clk (.X(clknet_4_10_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_11_0_clk (.X(clknet_4_11_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_12_0_clk (.X(clknet_4_12_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_13_0_clk (.X(clknet_4_13_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_14_0_clk (.X(clknet_4_14_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_15_0_clk (.X(clknet_4_15_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_4_8_0_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_4_11_0_clk));
 sg13g2_inv_2 clkload3 (.A(clknet_4_15_0_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_58_clk));
 sg13g2_buf_16 clkload5 (.A(clknet_leaf_60_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_leaf_1_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_3_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_57_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_59_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_8_clk));
 sg13g2_buf_16 clkload11 (.A(clknet_leaf_52_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_5_clk));
 sg13g2_buf_16 clkload13 (.A(clknet_leaf_14_clk));
 sg13g2_buf_16 clkload14 (.A(clknet_leaf_11_clk));
 sg13g2_buf_8 clkload15 (.A(clknet_leaf_12_clk));
 sg13g2_buf_16 clkload16 (.A(clknet_leaf_47_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_48_clk));
 sg13g2_buf_16 clkload18 (.A(clknet_leaf_39_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_51_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_40_clk));
 sg13g2_buf_16 clkload21 (.A(clknet_leaf_44_clk));
 sg13g2_buf_8 clkload22 (.A(clknet_leaf_49_clk));
 sg13g2_buf_16 clkload23 (.A(clknet_leaf_37_clk));
 sg13g2_buf_16 clkload24 (.A(clknet_leaf_42_clk));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_27_clk));
 sg13g2_buf_16 clkload26 (.A(clknet_leaf_28_clk));
 sg13g2_buf_8 clkload27 (.A(clknet_leaf_29_clk));
 sg13g2_inv_1 clkload28 (.A(clknet_leaf_23_clk));
 sg13g2_buf_8 clkload29 (.A(clknet_leaf_25_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_30_clk));
 sg13g2_inv_1 clkload31 (.A(clknet_leaf_33_clk));
 sg13g2_buf_8 clkload32 (.A(clknet_leaf_35_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00296_));
 sg13g2_antennanp ANTENNA_2 (.A(_00296_));
 sg13g2_antennanp ANTENNA_3 (.A(_00368_));
 sg13g2_antennanp ANTENNA_4 (.A(_00368_));
 sg13g2_antennanp ANTENNA_5 (.A(_05157_));
 sg13g2_antennanp ANTENNA_6 (.A(doe));
 sg13g2_antennanp ANTENNA_7 (.A(doe));
 sg13g2_antennanp ANTENNA_8 (.A(doe));
 sg13g2_antennanp ANTENNA_9 (.A(_00368_));
 sg13g2_antennanp ANTENNA_10 (.A(_00368_));
 sg13g2_antennanp ANTENNA_11 (.A(_05157_));
 sg13g2_antennanp ANTENNA_12 (.A(_00368_));
 sg13g2_antennanp ANTENNA_13 (.A(_00368_));
 sg13g2_antennanp ANTENNA_14 (.A(_00368_));
 sg13g2_antennanp ANTENNA_15 (.A(_00368_));
 sg13g2_antennanp ANTENNA_16 (.A(_00368_));
 sg13g2_antennanp ANTENNA_17 (.A(_00368_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_fill_2 FILLER_0_875 ();
 sg13g2_fill_1 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_fill_2 FILLER_1_875 ();
 sg13g2_fill_1 FILLER_1_877 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_2_868 ();
 sg13g2_fill_2 FILLER_2_875 ();
 sg13g2_fill_1 FILLER_2_877 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_decap_8 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_3_868 ();
 sg13g2_fill_2 FILLER_3_875 ();
 sg13g2_fill_1 FILLER_3_877 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_decap_8 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_4_868 ();
 sg13g2_fill_2 FILLER_4_875 ();
 sg13g2_fill_1 FILLER_4_877 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_decap_8 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_5_868 ();
 sg13g2_fill_2 FILLER_5_875 ();
 sg13g2_fill_1 FILLER_5_877 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_229 ();
 sg13g2_decap_4 FILLER_6_236 ();
 sg13g2_fill_1 FILLER_6_270 ();
 sg13g2_fill_1 FILLER_6_275 ();
 sg13g2_decap_4 FILLER_6_306 ();
 sg13g2_fill_2 FILLER_6_310 ();
 sg13g2_fill_2 FILLER_6_322 ();
 sg13g2_fill_1 FILLER_6_324 ();
 sg13g2_decap_4 FILLER_6_329 ();
 sg13g2_fill_2 FILLER_6_333 ();
 sg13g2_fill_2 FILLER_6_339 ();
 sg13g2_fill_1 FILLER_6_341 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_fill_1 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_403 ();
 sg13g2_decap_8 FILLER_6_410 ();
 sg13g2_decap_8 FILLER_6_417 ();
 sg13g2_decap_8 FILLER_6_424 ();
 sg13g2_decap_8 FILLER_6_431 ();
 sg13g2_decap_8 FILLER_6_438 ();
 sg13g2_decap_8 FILLER_6_445 ();
 sg13g2_decap_8 FILLER_6_452 ();
 sg13g2_decap_8 FILLER_6_459 ();
 sg13g2_decap_8 FILLER_6_466 ();
 sg13g2_decap_8 FILLER_6_473 ();
 sg13g2_decap_8 FILLER_6_480 ();
 sg13g2_decap_8 FILLER_6_487 ();
 sg13g2_decap_8 FILLER_6_494 ();
 sg13g2_decap_8 FILLER_6_501 ();
 sg13g2_decap_8 FILLER_6_508 ();
 sg13g2_decap_8 FILLER_6_515 ();
 sg13g2_decap_8 FILLER_6_522 ();
 sg13g2_decap_8 FILLER_6_529 ();
 sg13g2_decap_8 FILLER_6_536 ();
 sg13g2_decap_8 FILLER_6_543 ();
 sg13g2_decap_8 FILLER_6_550 ();
 sg13g2_decap_8 FILLER_6_557 ();
 sg13g2_decap_8 FILLER_6_564 ();
 sg13g2_decap_8 FILLER_6_571 ();
 sg13g2_decap_8 FILLER_6_578 ();
 sg13g2_decap_8 FILLER_6_585 ();
 sg13g2_decap_8 FILLER_6_592 ();
 sg13g2_decap_8 FILLER_6_599 ();
 sg13g2_decap_8 FILLER_6_606 ();
 sg13g2_decap_8 FILLER_6_613 ();
 sg13g2_decap_8 FILLER_6_620 ();
 sg13g2_decap_8 FILLER_6_627 ();
 sg13g2_decap_8 FILLER_6_634 ();
 sg13g2_decap_8 FILLER_6_641 ();
 sg13g2_decap_8 FILLER_6_648 ();
 sg13g2_decap_8 FILLER_6_655 ();
 sg13g2_decap_8 FILLER_6_662 ();
 sg13g2_decap_8 FILLER_6_669 ();
 sg13g2_decap_8 FILLER_6_676 ();
 sg13g2_decap_8 FILLER_6_683 ();
 sg13g2_decap_8 FILLER_6_690 ();
 sg13g2_decap_8 FILLER_6_697 ();
 sg13g2_decap_8 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_711 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_decap_8 FILLER_6_725 ();
 sg13g2_decap_8 FILLER_6_732 ();
 sg13g2_decap_8 FILLER_6_739 ();
 sg13g2_decap_8 FILLER_6_746 ();
 sg13g2_decap_8 FILLER_6_753 ();
 sg13g2_decap_8 FILLER_6_760 ();
 sg13g2_decap_8 FILLER_6_767 ();
 sg13g2_decap_8 FILLER_6_774 ();
 sg13g2_decap_8 FILLER_6_781 ();
 sg13g2_decap_8 FILLER_6_788 ();
 sg13g2_decap_8 FILLER_6_795 ();
 sg13g2_decap_8 FILLER_6_802 ();
 sg13g2_decap_8 FILLER_6_809 ();
 sg13g2_decap_8 FILLER_6_816 ();
 sg13g2_decap_8 FILLER_6_823 ();
 sg13g2_decap_8 FILLER_6_830 ();
 sg13g2_decap_8 FILLER_6_837 ();
 sg13g2_decap_8 FILLER_6_844 ();
 sg13g2_decap_8 FILLER_6_851 ();
 sg13g2_decap_8 FILLER_6_858 ();
 sg13g2_decap_8 FILLER_6_865 ();
 sg13g2_decap_4 FILLER_6_872 ();
 sg13g2_fill_2 FILLER_6_876 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_4 FILLER_7_203 ();
 sg13g2_fill_2 FILLER_7_207 ();
 sg13g2_decap_4 FILLER_7_213 ();
 sg13g2_fill_2 FILLER_7_347 ();
 sg13g2_fill_1 FILLER_7_349 ();
 sg13g2_decap_8 FILLER_7_425 ();
 sg13g2_decap_8 FILLER_7_432 ();
 sg13g2_decap_8 FILLER_7_439 ();
 sg13g2_decap_8 FILLER_7_446 ();
 sg13g2_decap_8 FILLER_7_453 ();
 sg13g2_decap_8 FILLER_7_460 ();
 sg13g2_decap_8 FILLER_7_467 ();
 sg13g2_decap_8 FILLER_7_474 ();
 sg13g2_decap_8 FILLER_7_481 ();
 sg13g2_decap_8 FILLER_7_488 ();
 sg13g2_decap_8 FILLER_7_495 ();
 sg13g2_decap_8 FILLER_7_502 ();
 sg13g2_decap_8 FILLER_7_509 ();
 sg13g2_decap_8 FILLER_7_516 ();
 sg13g2_decap_8 FILLER_7_523 ();
 sg13g2_decap_8 FILLER_7_530 ();
 sg13g2_decap_8 FILLER_7_537 ();
 sg13g2_decap_8 FILLER_7_544 ();
 sg13g2_decap_8 FILLER_7_551 ();
 sg13g2_decap_8 FILLER_7_558 ();
 sg13g2_decap_8 FILLER_7_565 ();
 sg13g2_decap_8 FILLER_7_572 ();
 sg13g2_decap_8 FILLER_7_579 ();
 sg13g2_decap_8 FILLER_7_586 ();
 sg13g2_decap_8 FILLER_7_593 ();
 sg13g2_decap_8 FILLER_7_600 ();
 sg13g2_decap_8 FILLER_7_607 ();
 sg13g2_decap_8 FILLER_7_614 ();
 sg13g2_decap_8 FILLER_7_621 ();
 sg13g2_decap_8 FILLER_7_628 ();
 sg13g2_decap_8 FILLER_7_635 ();
 sg13g2_decap_8 FILLER_7_642 ();
 sg13g2_decap_8 FILLER_7_649 ();
 sg13g2_decap_8 FILLER_7_656 ();
 sg13g2_decap_8 FILLER_7_663 ();
 sg13g2_decap_8 FILLER_7_670 ();
 sg13g2_decap_8 FILLER_7_677 ();
 sg13g2_decap_8 FILLER_7_684 ();
 sg13g2_decap_8 FILLER_7_691 ();
 sg13g2_decap_8 FILLER_7_698 ();
 sg13g2_decap_8 FILLER_7_705 ();
 sg13g2_decap_8 FILLER_7_712 ();
 sg13g2_decap_8 FILLER_7_719 ();
 sg13g2_decap_8 FILLER_7_726 ();
 sg13g2_decap_8 FILLER_7_733 ();
 sg13g2_decap_8 FILLER_7_740 ();
 sg13g2_decap_8 FILLER_7_747 ();
 sg13g2_decap_8 FILLER_7_754 ();
 sg13g2_decap_8 FILLER_7_761 ();
 sg13g2_decap_8 FILLER_7_768 ();
 sg13g2_decap_8 FILLER_7_775 ();
 sg13g2_decap_8 FILLER_7_782 ();
 sg13g2_decap_8 FILLER_7_789 ();
 sg13g2_decap_8 FILLER_7_796 ();
 sg13g2_decap_8 FILLER_7_803 ();
 sg13g2_decap_8 FILLER_7_810 ();
 sg13g2_decap_8 FILLER_7_817 ();
 sg13g2_decap_8 FILLER_7_824 ();
 sg13g2_decap_8 FILLER_7_831 ();
 sg13g2_decap_8 FILLER_7_838 ();
 sg13g2_decap_8 FILLER_7_845 ();
 sg13g2_decap_8 FILLER_7_852 ();
 sg13g2_decap_8 FILLER_7_859 ();
 sg13g2_decap_8 FILLER_7_866 ();
 sg13g2_decap_4 FILLER_7_873 ();
 sg13g2_fill_1 FILLER_7_877 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_fill_2 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_171 ();
 sg13g2_decap_8 FILLER_8_178 ();
 sg13g2_decap_8 FILLER_8_185 ();
 sg13g2_decap_8 FILLER_8_192 ();
 sg13g2_decap_8 FILLER_8_199 ();
 sg13g2_fill_2 FILLER_8_206 ();
 sg13g2_decap_4 FILLER_8_212 ();
 sg13g2_fill_2 FILLER_8_220 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_fill_2 FILLER_8_243 ();
 sg13g2_fill_2 FILLER_8_262 ();
 sg13g2_fill_1 FILLER_8_276 ();
 sg13g2_decap_4 FILLER_8_301 ();
 sg13g2_fill_1 FILLER_8_305 ();
 sg13g2_fill_1 FILLER_8_332 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_fill_2 FILLER_8_350 ();
 sg13g2_fill_1 FILLER_8_352 ();
 sg13g2_decap_4 FILLER_8_357 ();
 sg13g2_fill_1 FILLER_8_361 ();
 sg13g2_fill_2 FILLER_8_372 ();
 sg13g2_fill_1 FILLER_8_374 ();
 sg13g2_decap_4 FILLER_8_379 ();
 sg13g2_fill_1 FILLER_8_383 ();
 sg13g2_decap_4 FILLER_8_389 ();
 sg13g2_fill_1 FILLER_8_393 ();
 sg13g2_fill_1 FILLER_8_411 ();
 sg13g2_fill_1 FILLER_8_438 ();
 sg13g2_decap_8 FILLER_8_465 ();
 sg13g2_decap_8 FILLER_8_472 ();
 sg13g2_decap_8 FILLER_8_479 ();
 sg13g2_fill_2 FILLER_8_486 ();
 sg13g2_fill_1 FILLER_8_488 ();
 sg13g2_decap_8 FILLER_8_499 ();
 sg13g2_decap_8 FILLER_8_506 ();
 sg13g2_decap_8 FILLER_8_513 ();
 sg13g2_decap_8 FILLER_8_520 ();
 sg13g2_decap_8 FILLER_8_527 ();
 sg13g2_decap_8 FILLER_8_534 ();
 sg13g2_decap_8 FILLER_8_541 ();
 sg13g2_decap_8 FILLER_8_548 ();
 sg13g2_decap_8 FILLER_8_555 ();
 sg13g2_decap_8 FILLER_8_562 ();
 sg13g2_decap_8 FILLER_8_569 ();
 sg13g2_decap_8 FILLER_8_576 ();
 sg13g2_decap_8 FILLER_8_583 ();
 sg13g2_decap_8 FILLER_8_590 ();
 sg13g2_decap_8 FILLER_8_597 ();
 sg13g2_decap_8 FILLER_8_604 ();
 sg13g2_decap_8 FILLER_8_611 ();
 sg13g2_decap_8 FILLER_8_618 ();
 sg13g2_decap_8 FILLER_8_625 ();
 sg13g2_decap_8 FILLER_8_632 ();
 sg13g2_decap_8 FILLER_8_639 ();
 sg13g2_decap_8 FILLER_8_646 ();
 sg13g2_decap_8 FILLER_8_653 ();
 sg13g2_decap_8 FILLER_8_660 ();
 sg13g2_decap_8 FILLER_8_667 ();
 sg13g2_decap_8 FILLER_8_674 ();
 sg13g2_decap_8 FILLER_8_681 ();
 sg13g2_decap_8 FILLER_8_688 ();
 sg13g2_decap_8 FILLER_8_695 ();
 sg13g2_decap_8 FILLER_8_702 ();
 sg13g2_decap_8 FILLER_8_709 ();
 sg13g2_decap_8 FILLER_8_716 ();
 sg13g2_decap_8 FILLER_8_723 ();
 sg13g2_decap_8 FILLER_8_730 ();
 sg13g2_decap_8 FILLER_8_737 ();
 sg13g2_decap_8 FILLER_8_744 ();
 sg13g2_decap_8 FILLER_8_751 ();
 sg13g2_decap_8 FILLER_8_758 ();
 sg13g2_decap_8 FILLER_8_765 ();
 sg13g2_decap_8 FILLER_8_772 ();
 sg13g2_decap_8 FILLER_8_779 ();
 sg13g2_decap_8 FILLER_8_786 ();
 sg13g2_decap_8 FILLER_8_793 ();
 sg13g2_decap_8 FILLER_8_800 ();
 sg13g2_decap_8 FILLER_8_807 ();
 sg13g2_decap_8 FILLER_8_814 ();
 sg13g2_decap_8 FILLER_8_821 ();
 sg13g2_decap_8 FILLER_8_828 ();
 sg13g2_decap_8 FILLER_8_835 ();
 sg13g2_decap_8 FILLER_8_842 ();
 sg13g2_decap_8 FILLER_8_849 ();
 sg13g2_decap_8 FILLER_8_856 ();
 sg13g2_decap_8 FILLER_8_863 ();
 sg13g2_decap_8 FILLER_8_870 ();
 sg13g2_fill_1 FILLER_8_877 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_fill_2 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_188 ();
 sg13g2_decap_8 FILLER_9_195 ();
 sg13g2_fill_1 FILLER_9_232 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_fill_2 FILLER_9_245 ();
 sg13g2_fill_1 FILLER_9_247 ();
 sg13g2_decap_4 FILLER_9_274 ();
 sg13g2_fill_1 FILLER_9_283 ();
 sg13g2_fill_1 FILLER_9_288 ();
 sg13g2_fill_2 FILLER_9_319 ();
 sg13g2_fill_1 FILLER_9_321 ();
 sg13g2_decap_4 FILLER_9_342 ();
 sg13g2_fill_1 FILLER_9_372 ();
 sg13g2_decap_4 FILLER_9_377 ();
 sg13g2_fill_2 FILLER_9_415 ();
 sg13g2_fill_1 FILLER_9_417 ();
 sg13g2_fill_1 FILLER_9_421 ();
 sg13g2_fill_2 FILLER_9_426 ();
 sg13g2_fill_1 FILLER_9_428 ();
 sg13g2_decap_4 FILLER_9_475 ();
 sg13g2_fill_2 FILLER_9_479 ();
 sg13g2_fill_2 FILLER_9_491 ();
 sg13g2_fill_1 FILLER_9_493 ();
 sg13g2_decap_8 FILLER_9_520 ();
 sg13g2_decap_8 FILLER_9_527 ();
 sg13g2_decap_8 FILLER_9_534 ();
 sg13g2_decap_8 FILLER_9_541 ();
 sg13g2_decap_8 FILLER_9_548 ();
 sg13g2_decap_8 FILLER_9_555 ();
 sg13g2_decap_8 FILLER_9_562 ();
 sg13g2_decap_8 FILLER_9_569 ();
 sg13g2_decap_8 FILLER_9_576 ();
 sg13g2_decap_8 FILLER_9_583 ();
 sg13g2_decap_8 FILLER_9_590 ();
 sg13g2_decap_8 FILLER_9_597 ();
 sg13g2_decap_8 FILLER_9_604 ();
 sg13g2_decap_8 FILLER_9_611 ();
 sg13g2_decap_8 FILLER_9_618 ();
 sg13g2_decap_8 FILLER_9_625 ();
 sg13g2_decap_8 FILLER_9_632 ();
 sg13g2_decap_8 FILLER_9_639 ();
 sg13g2_decap_8 FILLER_9_646 ();
 sg13g2_decap_8 FILLER_9_653 ();
 sg13g2_decap_8 FILLER_9_660 ();
 sg13g2_decap_8 FILLER_9_667 ();
 sg13g2_decap_8 FILLER_9_674 ();
 sg13g2_decap_8 FILLER_9_681 ();
 sg13g2_decap_8 FILLER_9_688 ();
 sg13g2_decap_8 FILLER_9_695 ();
 sg13g2_decap_8 FILLER_9_702 ();
 sg13g2_decap_8 FILLER_9_709 ();
 sg13g2_decap_8 FILLER_9_716 ();
 sg13g2_decap_8 FILLER_9_723 ();
 sg13g2_decap_8 FILLER_9_730 ();
 sg13g2_decap_8 FILLER_9_737 ();
 sg13g2_decap_8 FILLER_9_744 ();
 sg13g2_decap_8 FILLER_9_751 ();
 sg13g2_decap_8 FILLER_9_758 ();
 sg13g2_decap_8 FILLER_9_765 ();
 sg13g2_decap_8 FILLER_9_772 ();
 sg13g2_decap_8 FILLER_9_779 ();
 sg13g2_decap_8 FILLER_9_786 ();
 sg13g2_decap_8 FILLER_9_793 ();
 sg13g2_decap_8 FILLER_9_800 ();
 sg13g2_decap_8 FILLER_9_807 ();
 sg13g2_decap_8 FILLER_9_814 ();
 sg13g2_decap_8 FILLER_9_821 ();
 sg13g2_decap_8 FILLER_9_828 ();
 sg13g2_decap_8 FILLER_9_835 ();
 sg13g2_decap_8 FILLER_9_842 ();
 sg13g2_decap_8 FILLER_9_849 ();
 sg13g2_decap_8 FILLER_9_856 ();
 sg13g2_decap_8 FILLER_9_863 ();
 sg13g2_decap_8 FILLER_9_870 ();
 sg13g2_fill_1 FILLER_9_877 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_fill_2 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_128 ();
 sg13g2_decap_8 FILLER_10_155 ();
 sg13g2_decap_8 FILLER_10_162 ();
 sg13g2_decap_8 FILLER_10_169 ();
 sg13g2_decap_4 FILLER_10_176 ();
 sg13g2_fill_2 FILLER_10_184 ();
 sg13g2_fill_1 FILLER_10_186 ();
 sg13g2_fill_1 FILLER_10_257 ();
 sg13g2_fill_1 FILLER_10_262 ();
 sg13g2_fill_1 FILLER_10_267 ();
 sg13g2_decap_4 FILLER_10_294 ();
 sg13g2_fill_1 FILLER_10_298 ();
 sg13g2_fill_2 FILLER_10_304 ();
 sg13g2_fill_1 FILLER_10_310 ();
 sg13g2_fill_2 FILLER_10_349 ();
 sg13g2_fill_1 FILLER_10_351 ();
 sg13g2_fill_1 FILLER_10_356 ();
 sg13g2_decap_4 FILLER_10_406 ();
 sg13g2_fill_2 FILLER_10_410 ();
 sg13g2_fill_1 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_425 ();
 sg13g2_decap_8 FILLER_10_432 ();
 sg13g2_decap_8 FILLER_10_439 ();
 sg13g2_decap_8 FILLER_10_450 ();
 sg13g2_fill_2 FILLER_10_461 ();
 sg13g2_fill_1 FILLER_10_466 ();
 sg13g2_fill_2 FILLER_10_470 ();
 sg13g2_fill_1 FILLER_10_472 ();
 sg13g2_decap_8 FILLER_10_507 ();
 sg13g2_decap_8 FILLER_10_514 ();
 sg13g2_decap_8 FILLER_10_521 ();
 sg13g2_decap_8 FILLER_10_528 ();
 sg13g2_decap_8 FILLER_10_535 ();
 sg13g2_decap_8 FILLER_10_542 ();
 sg13g2_decap_8 FILLER_10_549 ();
 sg13g2_decap_8 FILLER_10_556 ();
 sg13g2_decap_8 FILLER_10_563 ();
 sg13g2_decap_8 FILLER_10_570 ();
 sg13g2_decap_8 FILLER_10_577 ();
 sg13g2_decap_8 FILLER_10_584 ();
 sg13g2_decap_8 FILLER_10_591 ();
 sg13g2_decap_8 FILLER_10_598 ();
 sg13g2_decap_8 FILLER_10_605 ();
 sg13g2_decap_8 FILLER_10_612 ();
 sg13g2_decap_8 FILLER_10_619 ();
 sg13g2_decap_8 FILLER_10_626 ();
 sg13g2_decap_8 FILLER_10_633 ();
 sg13g2_decap_8 FILLER_10_640 ();
 sg13g2_decap_8 FILLER_10_647 ();
 sg13g2_decap_8 FILLER_10_654 ();
 sg13g2_decap_8 FILLER_10_661 ();
 sg13g2_decap_8 FILLER_10_668 ();
 sg13g2_decap_8 FILLER_10_675 ();
 sg13g2_decap_8 FILLER_10_682 ();
 sg13g2_decap_8 FILLER_10_689 ();
 sg13g2_decap_8 FILLER_10_696 ();
 sg13g2_decap_8 FILLER_10_703 ();
 sg13g2_decap_8 FILLER_10_710 ();
 sg13g2_decap_8 FILLER_10_717 ();
 sg13g2_decap_8 FILLER_10_724 ();
 sg13g2_decap_8 FILLER_10_731 ();
 sg13g2_decap_8 FILLER_10_738 ();
 sg13g2_decap_8 FILLER_10_745 ();
 sg13g2_decap_8 FILLER_10_752 ();
 sg13g2_decap_8 FILLER_10_759 ();
 sg13g2_decap_8 FILLER_10_766 ();
 sg13g2_decap_8 FILLER_10_773 ();
 sg13g2_decap_8 FILLER_10_780 ();
 sg13g2_decap_8 FILLER_10_787 ();
 sg13g2_decap_8 FILLER_10_794 ();
 sg13g2_decap_8 FILLER_10_801 ();
 sg13g2_decap_8 FILLER_10_808 ();
 sg13g2_decap_8 FILLER_10_815 ();
 sg13g2_decap_8 FILLER_10_822 ();
 sg13g2_decap_8 FILLER_10_829 ();
 sg13g2_decap_8 FILLER_10_836 ();
 sg13g2_decap_8 FILLER_10_843 ();
 sg13g2_decap_8 FILLER_10_850 ();
 sg13g2_decap_8 FILLER_10_857 ();
 sg13g2_decap_8 FILLER_10_864 ();
 sg13g2_decap_8 FILLER_10_871 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_fill_2 FILLER_11_120 ();
 sg13g2_fill_1 FILLER_11_122 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_fill_2 FILLER_11_133 ();
 sg13g2_fill_1 FILLER_11_135 ();
 sg13g2_fill_2 FILLER_11_140 ();
 sg13g2_fill_1 FILLER_11_142 ();
 sg13g2_fill_2 FILLER_11_195 ();
 sg13g2_fill_1 FILLER_11_197 ();
 sg13g2_fill_1 FILLER_11_237 ();
 sg13g2_fill_1 FILLER_11_242 ();
 sg13g2_fill_2 FILLER_11_248 ();
 sg13g2_fill_2 FILLER_11_254 ();
 sg13g2_fill_2 FILLER_11_265 ();
 sg13g2_fill_1 FILLER_11_284 ();
 sg13g2_fill_2 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_fill_2 FILLER_11_395 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_fill_1 FILLER_11_451 ();
 sg13g2_fill_2 FILLER_11_455 ();
 sg13g2_fill_1 FILLER_11_486 ();
 sg13g2_decap_8 FILLER_11_508 ();
 sg13g2_fill_2 FILLER_11_518 ();
 sg13g2_fill_2 FILLER_11_526 ();
 sg13g2_decap_8 FILLER_11_531 ();
 sg13g2_decap_8 FILLER_11_538 ();
 sg13g2_decap_8 FILLER_11_545 ();
 sg13g2_decap_8 FILLER_11_552 ();
 sg13g2_decap_8 FILLER_11_559 ();
 sg13g2_decap_8 FILLER_11_566 ();
 sg13g2_decap_8 FILLER_11_573 ();
 sg13g2_decap_8 FILLER_11_580 ();
 sg13g2_decap_8 FILLER_11_587 ();
 sg13g2_decap_8 FILLER_11_594 ();
 sg13g2_decap_8 FILLER_11_601 ();
 sg13g2_decap_8 FILLER_11_608 ();
 sg13g2_decap_8 FILLER_11_615 ();
 sg13g2_decap_8 FILLER_11_622 ();
 sg13g2_decap_8 FILLER_11_629 ();
 sg13g2_decap_8 FILLER_11_636 ();
 sg13g2_decap_8 FILLER_11_643 ();
 sg13g2_decap_8 FILLER_11_650 ();
 sg13g2_decap_8 FILLER_11_657 ();
 sg13g2_decap_8 FILLER_11_664 ();
 sg13g2_decap_8 FILLER_11_671 ();
 sg13g2_decap_8 FILLER_11_678 ();
 sg13g2_decap_8 FILLER_11_685 ();
 sg13g2_decap_8 FILLER_11_692 ();
 sg13g2_decap_8 FILLER_11_699 ();
 sg13g2_decap_8 FILLER_11_706 ();
 sg13g2_decap_8 FILLER_11_713 ();
 sg13g2_decap_8 FILLER_11_720 ();
 sg13g2_decap_8 FILLER_11_727 ();
 sg13g2_decap_8 FILLER_11_734 ();
 sg13g2_decap_8 FILLER_11_741 ();
 sg13g2_decap_8 FILLER_11_748 ();
 sg13g2_decap_8 FILLER_11_755 ();
 sg13g2_decap_8 FILLER_11_762 ();
 sg13g2_decap_8 FILLER_11_769 ();
 sg13g2_decap_8 FILLER_11_776 ();
 sg13g2_decap_8 FILLER_11_783 ();
 sg13g2_decap_8 FILLER_11_790 ();
 sg13g2_decap_8 FILLER_11_797 ();
 sg13g2_decap_8 FILLER_11_804 ();
 sg13g2_decap_8 FILLER_11_811 ();
 sg13g2_decap_8 FILLER_11_818 ();
 sg13g2_decap_8 FILLER_11_825 ();
 sg13g2_decap_8 FILLER_11_832 ();
 sg13g2_decap_8 FILLER_11_839 ();
 sg13g2_decap_8 FILLER_11_846 ();
 sg13g2_decap_8 FILLER_11_853 ();
 sg13g2_decap_8 FILLER_11_860 ();
 sg13g2_decap_8 FILLER_11_867 ();
 sg13g2_decap_4 FILLER_11_874 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_4 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_60 ();
 sg13g2_decap_4 FILLER_12_68 ();
 sg13g2_fill_2 FILLER_12_72 ();
 sg13g2_decap_4 FILLER_12_78 ();
 sg13g2_fill_2 FILLER_12_99 ();
 sg13g2_fill_1 FILLER_12_127 ();
 sg13g2_decap_4 FILLER_12_137 ();
 sg13g2_fill_1 FILLER_12_146 ();
 sg13g2_decap_4 FILLER_12_155 ();
 sg13g2_fill_2 FILLER_12_180 ();
 sg13g2_fill_1 FILLER_12_182 ();
 sg13g2_fill_1 FILLER_12_203 ();
 sg13g2_fill_1 FILLER_12_208 ();
 sg13g2_fill_1 FILLER_12_213 ();
 sg13g2_fill_1 FILLER_12_240 ();
 sg13g2_fill_1 FILLER_12_267 ();
 sg13g2_fill_1 FILLER_12_320 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_fill_1 FILLER_12_354 ();
 sg13g2_fill_1 FILLER_12_374 ();
 sg13g2_fill_1 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_409 ();
 sg13g2_fill_1 FILLER_12_415 ();
 sg13g2_decap_4 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_463 ();
 sg13g2_fill_2 FILLER_12_470 ();
 sg13g2_fill_2 FILLER_12_482 ();
 sg13g2_decap_8 FILLER_12_541 ();
 sg13g2_decap_8 FILLER_12_548 ();
 sg13g2_decap_8 FILLER_12_555 ();
 sg13g2_decap_8 FILLER_12_562 ();
 sg13g2_decap_8 FILLER_12_569 ();
 sg13g2_decap_8 FILLER_12_576 ();
 sg13g2_decap_8 FILLER_12_583 ();
 sg13g2_decap_8 FILLER_12_590 ();
 sg13g2_decap_8 FILLER_12_597 ();
 sg13g2_decap_8 FILLER_12_604 ();
 sg13g2_decap_8 FILLER_12_611 ();
 sg13g2_decap_8 FILLER_12_618 ();
 sg13g2_decap_8 FILLER_12_625 ();
 sg13g2_decap_8 FILLER_12_632 ();
 sg13g2_decap_8 FILLER_12_639 ();
 sg13g2_decap_8 FILLER_12_646 ();
 sg13g2_decap_8 FILLER_12_653 ();
 sg13g2_decap_8 FILLER_12_660 ();
 sg13g2_decap_8 FILLER_12_667 ();
 sg13g2_decap_8 FILLER_12_674 ();
 sg13g2_decap_8 FILLER_12_681 ();
 sg13g2_decap_8 FILLER_12_688 ();
 sg13g2_decap_8 FILLER_12_695 ();
 sg13g2_decap_8 FILLER_12_702 ();
 sg13g2_decap_8 FILLER_12_709 ();
 sg13g2_decap_8 FILLER_12_716 ();
 sg13g2_decap_8 FILLER_12_723 ();
 sg13g2_decap_8 FILLER_12_730 ();
 sg13g2_decap_8 FILLER_12_737 ();
 sg13g2_decap_8 FILLER_12_744 ();
 sg13g2_decap_8 FILLER_12_751 ();
 sg13g2_decap_8 FILLER_12_758 ();
 sg13g2_decap_8 FILLER_12_765 ();
 sg13g2_decap_8 FILLER_12_772 ();
 sg13g2_decap_8 FILLER_12_779 ();
 sg13g2_decap_8 FILLER_12_786 ();
 sg13g2_decap_8 FILLER_12_793 ();
 sg13g2_decap_8 FILLER_12_800 ();
 sg13g2_decap_8 FILLER_12_807 ();
 sg13g2_decap_8 FILLER_12_814 ();
 sg13g2_decap_8 FILLER_12_821 ();
 sg13g2_decap_8 FILLER_12_828 ();
 sg13g2_decap_8 FILLER_12_835 ();
 sg13g2_decap_8 FILLER_12_842 ();
 sg13g2_decap_8 FILLER_12_849 ();
 sg13g2_decap_8 FILLER_12_856 ();
 sg13g2_decap_8 FILLER_12_863 ();
 sg13g2_decap_8 FILLER_12_870 ();
 sg13g2_fill_1 FILLER_12_877 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_35 ();
 sg13g2_fill_1 FILLER_13_37 ();
 sg13g2_decap_4 FILLER_13_48 ();
 sg13g2_fill_2 FILLER_13_62 ();
 sg13g2_decap_4 FILLER_13_94 ();
 sg13g2_fill_2 FILLER_13_101 ();
 sg13g2_fill_1 FILLER_13_103 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_152 ();
 sg13g2_decap_8 FILLER_13_159 ();
 sg13g2_decap_4 FILLER_13_166 ();
 sg13g2_fill_2 FILLER_13_170 ();
 sg13g2_fill_2 FILLER_13_198 ();
 sg13g2_fill_2 FILLER_13_230 ();
 sg13g2_decap_4 FILLER_13_286 ();
 sg13g2_fill_2 FILLER_13_314 ();
 sg13g2_decap_4 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_4 FILLER_13_437 ();
 sg13g2_decap_8 FILLER_13_449 ();
 sg13g2_decap_8 FILLER_13_456 ();
 sg13g2_decap_4 FILLER_13_463 ();
 sg13g2_fill_2 FILLER_13_467 ();
 sg13g2_decap_4 FILLER_13_490 ();
 sg13g2_fill_1 FILLER_13_494 ();
 sg13g2_decap_8 FILLER_13_513 ();
 sg13g2_decap_8 FILLER_13_520 ();
 sg13g2_decap_8 FILLER_13_527 ();
 sg13g2_decap_8 FILLER_13_534 ();
 sg13g2_decap_8 FILLER_13_541 ();
 sg13g2_decap_8 FILLER_13_548 ();
 sg13g2_decap_8 FILLER_13_555 ();
 sg13g2_decap_8 FILLER_13_562 ();
 sg13g2_decap_8 FILLER_13_569 ();
 sg13g2_decap_8 FILLER_13_576 ();
 sg13g2_decap_8 FILLER_13_583 ();
 sg13g2_decap_8 FILLER_13_590 ();
 sg13g2_decap_8 FILLER_13_597 ();
 sg13g2_decap_8 FILLER_13_604 ();
 sg13g2_decap_8 FILLER_13_611 ();
 sg13g2_decap_8 FILLER_13_618 ();
 sg13g2_decap_8 FILLER_13_625 ();
 sg13g2_decap_8 FILLER_13_632 ();
 sg13g2_decap_8 FILLER_13_639 ();
 sg13g2_decap_8 FILLER_13_646 ();
 sg13g2_decap_8 FILLER_13_653 ();
 sg13g2_decap_8 FILLER_13_660 ();
 sg13g2_decap_8 FILLER_13_667 ();
 sg13g2_decap_8 FILLER_13_674 ();
 sg13g2_decap_8 FILLER_13_681 ();
 sg13g2_decap_8 FILLER_13_688 ();
 sg13g2_decap_8 FILLER_13_695 ();
 sg13g2_decap_8 FILLER_13_702 ();
 sg13g2_decap_8 FILLER_13_709 ();
 sg13g2_decap_8 FILLER_13_716 ();
 sg13g2_decap_8 FILLER_13_723 ();
 sg13g2_decap_8 FILLER_13_730 ();
 sg13g2_decap_8 FILLER_13_737 ();
 sg13g2_decap_8 FILLER_13_744 ();
 sg13g2_decap_8 FILLER_13_751 ();
 sg13g2_decap_8 FILLER_13_758 ();
 sg13g2_decap_8 FILLER_13_765 ();
 sg13g2_decap_8 FILLER_13_772 ();
 sg13g2_decap_8 FILLER_13_779 ();
 sg13g2_decap_8 FILLER_13_786 ();
 sg13g2_decap_8 FILLER_13_793 ();
 sg13g2_decap_8 FILLER_13_800 ();
 sg13g2_decap_8 FILLER_13_807 ();
 sg13g2_decap_8 FILLER_13_814 ();
 sg13g2_decap_8 FILLER_13_821 ();
 sg13g2_decap_8 FILLER_13_828 ();
 sg13g2_decap_8 FILLER_13_835 ();
 sg13g2_decap_8 FILLER_13_842 ();
 sg13g2_decap_8 FILLER_13_849 ();
 sg13g2_decap_8 FILLER_13_856 ();
 sg13g2_decap_8 FILLER_13_863 ();
 sg13g2_decap_8 FILLER_13_870 ();
 sg13g2_fill_1 FILLER_13_877 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_65 ();
 sg13g2_fill_1 FILLER_14_67 ();
 sg13g2_fill_2 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_128 ();
 sg13g2_fill_1 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_160 ();
 sg13g2_fill_2 FILLER_14_167 ();
 sg13g2_fill_1 FILLER_14_169 ();
 sg13g2_decap_8 FILLER_14_204 ();
 sg13g2_fill_2 FILLER_14_236 ();
 sg13g2_fill_1 FILLER_14_238 ();
 sg13g2_fill_1 FILLER_14_243 ();
 sg13g2_fill_1 FILLER_14_270 ();
 sg13g2_fill_1 FILLER_14_301 ();
 sg13g2_fill_1 FILLER_14_323 ();
 sg13g2_fill_1 FILLER_14_345 ();
 sg13g2_fill_2 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_426 ();
 sg13g2_fill_1 FILLER_14_433 ();
 sg13g2_fill_2 FILLER_14_499 ();
 sg13g2_fill_1 FILLER_14_501 ();
 sg13g2_decap_4 FILLER_14_528 ();
 sg13g2_decap_8 FILLER_14_545 ();
 sg13g2_decap_8 FILLER_14_552 ();
 sg13g2_decap_8 FILLER_14_559 ();
 sg13g2_decap_8 FILLER_14_566 ();
 sg13g2_decap_8 FILLER_14_573 ();
 sg13g2_decap_8 FILLER_14_580 ();
 sg13g2_decap_8 FILLER_14_587 ();
 sg13g2_decap_8 FILLER_14_594 ();
 sg13g2_decap_8 FILLER_14_601 ();
 sg13g2_decap_8 FILLER_14_608 ();
 sg13g2_decap_8 FILLER_14_615 ();
 sg13g2_decap_8 FILLER_14_622 ();
 sg13g2_decap_8 FILLER_14_629 ();
 sg13g2_decap_8 FILLER_14_636 ();
 sg13g2_decap_8 FILLER_14_643 ();
 sg13g2_decap_8 FILLER_14_650 ();
 sg13g2_decap_8 FILLER_14_657 ();
 sg13g2_decap_8 FILLER_14_664 ();
 sg13g2_decap_8 FILLER_14_671 ();
 sg13g2_decap_8 FILLER_14_678 ();
 sg13g2_decap_8 FILLER_14_685 ();
 sg13g2_decap_8 FILLER_14_692 ();
 sg13g2_decap_8 FILLER_14_699 ();
 sg13g2_decap_8 FILLER_14_706 ();
 sg13g2_decap_8 FILLER_14_713 ();
 sg13g2_decap_8 FILLER_14_720 ();
 sg13g2_decap_8 FILLER_14_727 ();
 sg13g2_decap_8 FILLER_14_734 ();
 sg13g2_decap_8 FILLER_14_741 ();
 sg13g2_decap_8 FILLER_14_748 ();
 sg13g2_decap_8 FILLER_14_755 ();
 sg13g2_decap_8 FILLER_14_762 ();
 sg13g2_decap_8 FILLER_14_769 ();
 sg13g2_decap_8 FILLER_14_776 ();
 sg13g2_decap_8 FILLER_14_783 ();
 sg13g2_decap_8 FILLER_14_790 ();
 sg13g2_decap_8 FILLER_14_797 ();
 sg13g2_decap_8 FILLER_14_804 ();
 sg13g2_decap_8 FILLER_14_811 ();
 sg13g2_decap_8 FILLER_14_818 ();
 sg13g2_decap_8 FILLER_14_825 ();
 sg13g2_decap_8 FILLER_14_832 ();
 sg13g2_decap_8 FILLER_14_839 ();
 sg13g2_decap_8 FILLER_14_846 ();
 sg13g2_decap_8 FILLER_14_853 ();
 sg13g2_decap_8 FILLER_14_860 ();
 sg13g2_decap_8 FILLER_14_867 ();
 sg13g2_decap_4 FILLER_14_874 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_12 ();
 sg13g2_decap_4 FILLER_15_19 ();
 sg13g2_fill_1 FILLER_15_23 ();
 sg13g2_fill_2 FILLER_15_27 ();
 sg13g2_decap_4 FILLER_15_55 ();
 sg13g2_fill_1 FILLER_15_66 ();
 sg13g2_fill_2 FILLER_15_110 ();
 sg13g2_fill_1 FILLER_15_143 ();
 sg13g2_fill_1 FILLER_15_204 ();
 sg13g2_fill_2 FILLER_15_244 ();
 sg13g2_fill_1 FILLER_15_246 ();
 sg13g2_fill_1 FILLER_15_252 ();
 sg13g2_fill_2 FILLER_15_282 ();
 sg13g2_fill_1 FILLER_15_284 ();
 sg13g2_fill_1 FILLER_15_306 ();
 sg13g2_fill_1 FILLER_15_310 ();
 sg13g2_fill_1 FILLER_15_332 ();
 sg13g2_fill_2 FILLER_15_336 ();
 sg13g2_fill_2 FILLER_15_341 ();
 sg13g2_decap_4 FILLER_15_351 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_fill_1 FILLER_15_410 ();
 sg13g2_fill_2 FILLER_15_420 ();
 sg13g2_decap_4 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_436 ();
 sg13g2_decap_8 FILLER_15_447 ();
 sg13g2_fill_2 FILLER_15_496 ();
 sg13g2_fill_2 FILLER_15_502 ();
 sg13g2_fill_2 FILLER_15_514 ();
 sg13g2_fill_1 FILLER_15_516 ();
 sg13g2_decap_8 FILLER_15_521 ();
 sg13g2_decap_8 FILLER_15_565 ();
 sg13g2_decap_8 FILLER_15_572 ();
 sg13g2_decap_8 FILLER_15_579 ();
 sg13g2_decap_8 FILLER_15_586 ();
 sg13g2_decap_8 FILLER_15_593 ();
 sg13g2_decap_8 FILLER_15_600 ();
 sg13g2_decap_8 FILLER_15_607 ();
 sg13g2_decap_8 FILLER_15_614 ();
 sg13g2_decap_8 FILLER_15_621 ();
 sg13g2_decap_8 FILLER_15_628 ();
 sg13g2_decap_8 FILLER_15_635 ();
 sg13g2_decap_8 FILLER_15_642 ();
 sg13g2_decap_8 FILLER_15_649 ();
 sg13g2_decap_8 FILLER_15_656 ();
 sg13g2_decap_8 FILLER_15_663 ();
 sg13g2_decap_8 FILLER_15_670 ();
 sg13g2_decap_8 FILLER_15_677 ();
 sg13g2_decap_8 FILLER_15_684 ();
 sg13g2_decap_8 FILLER_15_691 ();
 sg13g2_decap_8 FILLER_15_698 ();
 sg13g2_decap_8 FILLER_15_705 ();
 sg13g2_decap_8 FILLER_15_712 ();
 sg13g2_decap_8 FILLER_15_719 ();
 sg13g2_decap_8 FILLER_15_726 ();
 sg13g2_decap_8 FILLER_15_733 ();
 sg13g2_decap_8 FILLER_15_740 ();
 sg13g2_decap_8 FILLER_15_747 ();
 sg13g2_decap_8 FILLER_15_754 ();
 sg13g2_decap_8 FILLER_15_761 ();
 sg13g2_decap_8 FILLER_15_768 ();
 sg13g2_decap_8 FILLER_15_775 ();
 sg13g2_decap_8 FILLER_15_782 ();
 sg13g2_decap_8 FILLER_15_789 ();
 sg13g2_decap_8 FILLER_15_796 ();
 sg13g2_decap_8 FILLER_15_803 ();
 sg13g2_decap_8 FILLER_15_810 ();
 sg13g2_decap_8 FILLER_15_817 ();
 sg13g2_decap_8 FILLER_15_824 ();
 sg13g2_decap_8 FILLER_15_831 ();
 sg13g2_decap_8 FILLER_15_838 ();
 sg13g2_decap_8 FILLER_15_845 ();
 sg13g2_decap_8 FILLER_15_852 ();
 sg13g2_decap_8 FILLER_15_859 ();
 sg13g2_decap_8 FILLER_15_866 ();
 sg13g2_decap_4 FILLER_15_873 ();
 sg13g2_fill_1 FILLER_15_877 ();
 sg13g2_fill_1 FILLER_16_36 ();
 sg13g2_decap_4 FILLER_16_41 ();
 sg13g2_fill_1 FILLER_16_74 ();
 sg13g2_fill_2 FILLER_16_79 ();
 sg13g2_decap_8 FILLER_16_102 ();
 sg13g2_fill_2 FILLER_16_109 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_fill_1 FILLER_16_147 ();
 sg13g2_fill_2 FILLER_16_174 ();
 sg13g2_fill_1 FILLER_16_212 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_250 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_269 ();
 sg13g2_fill_1 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_289 ();
 sg13g2_fill_1 FILLER_16_296 ();
 sg13g2_fill_2 FILLER_16_310 ();
 sg13g2_fill_1 FILLER_16_312 ();
 sg13g2_fill_1 FILLER_16_316 ();
 sg13g2_fill_2 FILLER_16_320 ();
 sg13g2_fill_2 FILLER_16_327 ();
 sg13g2_fill_1 FILLER_16_354 ();
 sg13g2_fill_2 FILLER_16_387 ();
 sg13g2_fill_2 FILLER_16_400 ();
 sg13g2_fill_1 FILLER_16_402 ();
 sg13g2_fill_2 FILLER_16_431 ();
 sg13g2_fill_1 FILLER_16_433 ();
 sg13g2_decap_4 FILLER_16_447 ();
 sg13g2_fill_2 FILLER_16_504 ();
 sg13g2_decap_4 FILLER_16_532 ();
 sg13g2_fill_1 FILLER_16_536 ();
 sg13g2_fill_2 FILLER_16_564 ();
 sg13g2_fill_1 FILLER_16_566 ();
 sg13g2_decap_8 FILLER_16_593 ();
 sg13g2_decap_8 FILLER_16_600 ();
 sg13g2_decap_8 FILLER_16_607 ();
 sg13g2_decap_8 FILLER_16_614 ();
 sg13g2_decap_8 FILLER_16_621 ();
 sg13g2_decap_8 FILLER_16_628 ();
 sg13g2_decap_8 FILLER_16_635 ();
 sg13g2_decap_8 FILLER_16_642 ();
 sg13g2_decap_8 FILLER_16_649 ();
 sg13g2_decap_8 FILLER_16_656 ();
 sg13g2_decap_8 FILLER_16_663 ();
 sg13g2_decap_8 FILLER_16_670 ();
 sg13g2_decap_8 FILLER_16_677 ();
 sg13g2_decap_8 FILLER_16_684 ();
 sg13g2_decap_8 FILLER_16_691 ();
 sg13g2_decap_8 FILLER_16_698 ();
 sg13g2_decap_8 FILLER_16_705 ();
 sg13g2_decap_8 FILLER_16_712 ();
 sg13g2_decap_8 FILLER_16_719 ();
 sg13g2_decap_8 FILLER_16_726 ();
 sg13g2_decap_8 FILLER_16_733 ();
 sg13g2_decap_8 FILLER_16_740 ();
 sg13g2_decap_8 FILLER_16_747 ();
 sg13g2_decap_8 FILLER_16_754 ();
 sg13g2_decap_8 FILLER_16_761 ();
 sg13g2_decap_8 FILLER_16_768 ();
 sg13g2_decap_8 FILLER_16_775 ();
 sg13g2_decap_8 FILLER_16_782 ();
 sg13g2_decap_8 FILLER_16_789 ();
 sg13g2_decap_8 FILLER_16_796 ();
 sg13g2_decap_8 FILLER_16_803 ();
 sg13g2_decap_8 FILLER_16_810 ();
 sg13g2_decap_8 FILLER_16_817 ();
 sg13g2_decap_8 FILLER_16_824 ();
 sg13g2_decap_8 FILLER_16_831 ();
 sg13g2_decap_8 FILLER_16_838 ();
 sg13g2_decap_8 FILLER_16_845 ();
 sg13g2_decap_8 FILLER_16_852 ();
 sg13g2_decap_8 FILLER_16_859 ();
 sg13g2_decap_8 FILLER_16_866 ();
 sg13g2_decap_4 FILLER_16_873 ();
 sg13g2_fill_1 FILLER_16_877 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_11 ();
 sg13g2_decap_4 FILLER_17_18 ();
 sg13g2_fill_1 FILLER_17_31 ();
 sg13g2_fill_1 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_61 ();
 sg13g2_fill_1 FILLER_17_68 ();
 sg13g2_fill_2 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_137 ();
 sg13g2_fill_1 FILLER_17_144 ();
 sg13g2_decap_8 FILLER_17_179 ();
 sg13g2_decap_4 FILLER_17_186 ();
 sg13g2_decap_8 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_209 ();
 sg13g2_fill_2 FILLER_17_216 ();
 sg13g2_fill_1 FILLER_17_218 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_259 ();
 sg13g2_decap_4 FILLER_17_286 ();
 sg13g2_fill_1 FILLER_17_290 ();
 sg13g2_fill_1 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_decap_4 FILLER_17_339 ();
 sg13g2_fill_1 FILLER_17_343 ();
 sg13g2_fill_1 FILLER_17_359 ();
 sg13g2_fill_2 FILLER_17_391 ();
 sg13g2_fill_2 FILLER_17_400 ();
 sg13g2_fill_1 FILLER_17_402 ();
 sg13g2_fill_1 FILLER_17_434 ();
 sg13g2_decap_4 FILLER_17_481 ();
 sg13g2_fill_1 FILLER_17_485 ();
 sg13g2_fill_1 FILLER_17_516 ();
 sg13g2_decap_4 FILLER_17_543 ();
 sg13g2_decap_8 FILLER_17_568 ();
 sg13g2_fill_1 FILLER_17_575 ();
 sg13g2_decap_8 FILLER_17_580 ();
 sg13g2_decap_8 FILLER_17_587 ();
 sg13g2_decap_8 FILLER_17_594 ();
 sg13g2_decap_8 FILLER_17_601 ();
 sg13g2_decap_8 FILLER_17_608 ();
 sg13g2_decap_8 FILLER_17_615 ();
 sg13g2_decap_8 FILLER_17_622 ();
 sg13g2_decap_8 FILLER_17_629 ();
 sg13g2_decap_8 FILLER_17_636 ();
 sg13g2_decap_8 FILLER_17_643 ();
 sg13g2_decap_8 FILLER_17_650 ();
 sg13g2_decap_8 FILLER_17_657 ();
 sg13g2_decap_8 FILLER_17_664 ();
 sg13g2_decap_8 FILLER_17_671 ();
 sg13g2_decap_8 FILLER_17_678 ();
 sg13g2_decap_8 FILLER_17_685 ();
 sg13g2_decap_8 FILLER_17_692 ();
 sg13g2_decap_8 FILLER_17_699 ();
 sg13g2_decap_8 FILLER_17_706 ();
 sg13g2_decap_8 FILLER_17_713 ();
 sg13g2_decap_8 FILLER_17_720 ();
 sg13g2_decap_8 FILLER_17_727 ();
 sg13g2_decap_8 FILLER_17_734 ();
 sg13g2_decap_8 FILLER_17_741 ();
 sg13g2_decap_8 FILLER_17_748 ();
 sg13g2_decap_8 FILLER_17_755 ();
 sg13g2_decap_8 FILLER_17_762 ();
 sg13g2_decap_8 FILLER_17_769 ();
 sg13g2_decap_8 FILLER_17_776 ();
 sg13g2_decap_8 FILLER_17_783 ();
 sg13g2_decap_8 FILLER_17_790 ();
 sg13g2_decap_8 FILLER_17_797 ();
 sg13g2_decap_8 FILLER_17_804 ();
 sg13g2_decap_8 FILLER_17_811 ();
 sg13g2_decap_8 FILLER_17_818 ();
 sg13g2_decap_8 FILLER_17_825 ();
 sg13g2_decap_8 FILLER_17_832 ();
 sg13g2_decap_8 FILLER_17_839 ();
 sg13g2_decap_8 FILLER_17_846 ();
 sg13g2_decap_8 FILLER_17_853 ();
 sg13g2_decap_8 FILLER_17_860 ();
 sg13g2_decap_8 FILLER_17_867 ();
 sg13g2_decap_4 FILLER_17_874 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_30 ();
 sg13g2_fill_1 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_65 ();
 sg13g2_fill_2 FILLER_18_72 ();
 sg13g2_fill_2 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_102 ();
 sg13g2_fill_2 FILLER_18_109 ();
 sg13g2_fill_2 FILLER_18_137 ();
 sg13g2_fill_1 FILLER_18_139 ();
 sg13g2_fill_1 FILLER_18_184 ();
 sg13g2_fill_2 FILLER_18_203 ();
 sg13g2_fill_1 FILLER_18_210 ();
 sg13g2_fill_2 FILLER_18_215 ();
 sg13g2_fill_1 FILLER_18_227 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_4 FILLER_18_276 ();
 sg13g2_fill_1 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_286 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_fill_1 FILLER_18_312 ();
 sg13g2_fill_1 FILLER_18_321 ();
 sg13g2_decap_8 FILLER_18_327 ();
 sg13g2_fill_1 FILLER_18_334 ();
 sg13g2_fill_1 FILLER_18_357 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_2 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_436 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_4 FILLER_18_455 ();
 sg13g2_fill_2 FILLER_18_459 ();
 sg13g2_fill_1 FILLER_18_519 ();
 sg13g2_fill_2 FILLER_18_534 ();
 sg13g2_fill_2 FILLER_18_569 ();
 sg13g2_decap_4 FILLER_18_585 ();
 sg13g2_fill_1 FILLER_18_589 ();
 sg13g2_decap_8 FILLER_18_598 ();
 sg13g2_decap_8 FILLER_18_605 ();
 sg13g2_decap_8 FILLER_18_612 ();
 sg13g2_decap_8 FILLER_18_619 ();
 sg13g2_decap_8 FILLER_18_626 ();
 sg13g2_decap_8 FILLER_18_633 ();
 sg13g2_decap_8 FILLER_18_640 ();
 sg13g2_decap_8 FILLER_18_647 ();
 sg13g2_decap_8 FILLER_18_654 ();
 sg13g2_decap_8 FILLER_18_661 ();
 sg13g2_decap_8 FILLER_18_668 ();
 sg13g2_decap_8 FILLER_18_675 ();
 sg13g2_decap_8 FILLER_18_682 ();
 sg13g2_decap_8 FILLER_18_689 ();
 sg13g2_decap_8 FILLER_18_696 ();
 sg13g2_decap_8 FILLER_18_703 ();
 sg13g2_decap_8 FILLER_18_710 ();
 sg13g2_decap_8 FILLER_18_717 ();
 sg13g2_decap_8 FILLER_18_724 ();
 sg13g2_decap_8 FILLER_18_731 ();
 sg13g2_decap_8 FILLER_18_738 ();
 sg13g2_decap_8 FILLER_18_745 ();
 sg13g2_decap_8 FILLER_18_752 ();
 sg13g2_decap_8 FILLER_18_759 ();
 sg13g2_decap_8 FILLER_18_766 ();
 sg13g2_decap_8 FILLER_18_773 ();
 sg13g2_decap_8 FILLER_18_780 ();
 sg13g2_decap_8 FILLER_18_787 ();
 sg13g2_decap_8 FILLER_18_794 ();
 sg13g2_decap_8 FILLER_18_801 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_8 FILLER_18_815 ();
 sg13g2_decap_8 FILLER_18_822 ();
 sg13g2_decap_8 FILLER_18_829 ();
 sg13g2_decap_8 FILLER_18_836 ();
 sg13g2_decap_8 FILLER_18_843 ();
 sg13g2_decap_8 FILLER_18_850 ();
 sg13g2_decap_8 FILLER_18_857 ();
 sg13g2_decap_8 FILLER_18_864 ();
 sg13g2_decap_8 FILLER_18_871 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_53 ();
 sg13g2_decap_4 FILLER_19_69 ();
 sg13g2_fill_2 FILLER_19_73 ();
 sg13g2_fill_2 FILLER_19_96 ();
 sg13g2_fill_1 FILLER_19_118 ();
 sg13g2_fill_1 FILLER_19_127 ();
 sg13g2_decap_8 FILLER_19_136 ();
 sg13g2_fill_1 FILLER_19_153 ();
 sg13g2_fill_2 FILLER_19_158 ();
 sg13g2_decap_4 FILLER_19_226 ();
 sg13g2_decap_8 FILLER_19_236 ();
 sg13g2_decap_4 FILLER_19_243 ();
 sg13g2_fill_2 FILLER_19_272 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_fill_2 FILLER_19_288 ();
 sg13g2_decap_4 FILLER_19_319 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_4 FILLER_19_336 ();
 sg13g2_fill_1 FILLER_19_340 ();
 sg13g2_fill_2 FILLER_19_345 ();
 sg13g2_fill_1 FILLER_19_347 ();
 sg13g2_decap_4 FILLER_19_353 ();
 sg13g2_fill_1 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_363 ();
 sg13g2_fill_1 FILLER_19_370 ();
 sg13g2_fill_1 FILLER_19_380 ();
 sg13g2_fill_1 FILLER_19_420 ();
 sg13g2_fill_1 FILLER_19_426 ();
 sg13g2_decap_8 FILLER_19_436 ();
 sg13g2_fill_2 FILLER_19_443 ();
 sg13g2_fill_2 FILLER_19_471 ();
 sg13g2_fill_1 FILLER_19_569 ();
 sg13g2_decap_8 FILLER_19_621 ();
 sg13g2_decap_8 FILLER_19_628 ();
 sg13g2_decap_8 FILLER_19_635 ();
 sg13g2_decap_8 FILLER_19_642 ();
 sg13g2_decap_8 FILLER_19_649 ();
 sg13g2_decap_8 FILLER_19_656 ();
 sg13g2_decap_8 FILLER_19_663 ();
 sg13g2_decap_8 FILLER_19_670 ();
 sg13g2_decap_8 FILLER_19_677 ();
 sg13g2_decap_8 FILLER_19_684 ();
 sg13g2_decap_8 FILLER_19_691 ();
 sg13g2_decap_8 FILLER_19_698 ();
 sg13g2_decap_8 FILLER_19_705 ();
 sg13g2_decap_8 FILLER_19_712 ();
 sg13g2_decap_8 FILLER_19_719 ();
 sg13g2_decap_8 FILLER_19_726 ();
 sg13g2_decap_8 FILLER_19_733 ();
 sg13g2_decap_8 FILLER_19_740 ();
 sg13g2_decap_8 FILLER_19_747 ();
 sg13g2_decap_8 FILLER_19_754 ();
 sg13g2_decap_8 FILLER_19_761 ();
 sg13g2_decap_8 FILLER_19_768 ();
 sg13g2_decap_8 FILLER_19_775 ();
 sg13g2_decap_8 FILLER_19_782 ();
 sg13g2_decap_8 FILLER_19_789 ();
 sg13g2_decap_8 FILLER_19_796 ();
 sg13g2_decap_8 FILLER_19_803 ();
 sg13g2_decap_8 FILLER_19_810 ();
 sg13g2_decap_8 FILLER_19_817 ();
 sg13g2_decap_8 FILLER_19_824 ();
 sg13g2_decap_8 FILLER_19_831 ();
 sg13g2_decap_8 FILLER_19_838 ();
 sg13g2_decap_8 FILLER_19_845 ();
 sg13g2_decap_8 FILLER_19_852 ();
 sg13g2_decap_8 FILLER_19_859 ();
 sg13g2_decap_8 FILLER_19_866 ();
 sg13g2_decap_4 FILLER_19_873 ();
 sg13g2_fill_1 FILLER_19_877 ();
 sg13g2_fill_1 FILLER_20_26 ();
 sg13g2_fill_2 FILLER_20_37 ();
 sg13g2_fill_1 FILLER_20_39 ();
 sg13g2_decap_4 FILLER_20_78 ();
 sg13g2_fill_1 FILLER_20_82 ();
 sg13g2_fill_2 FILLER_20_108 ();
 sg13g2_fill_2 FILLER_20_136 ();
 sg13g2_fill_2 FILLER_20_143 ();
 sg13g2_fill_2 FILLER_20_171 ();
 sg13g2_fill_2 FILLER_20_199 ();
 sg13g2_fill_1 FILLER_20_247 ();
 sg13g2_fill_2 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_271 ();
 sg13g2_fill_1 FILLER_20_288 ();
 sg13g2_fill_1 FILLER_20_321 ();
 sg13g2_fill_2 FILLER_20_326 ();
 sg13g2_fill_1 FILLER_20_328 ();
 sg13g2_fill_2 FILLER_20_343 ();
 sg13g2_fill_1 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_351 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_fill_1 FILLER_20_394 ();
 sg13g2_fill_1 FILLER_20_400 ();
 sg13g2_fill_1 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_428 ();
 sg13g2_fill_1 FILLER_20_434 ();
 sg13g2_decap_4 FILLER_20_439 ();
 sg13g2_fill_2 FILLER_20_443 ();
 sg13g2_decap_4 FILLER_20_450 ();
 sg13g2_fill_2 FILLER_20_454 ();
 sg13g2_fill_1 FILLER_20_466 ();
 sg13g2_fill_1 FILLER_20_496 ();
 sg13g2_fill_1 FILLER_20_509 ();
 sg13g2_fill_2 FILLER_20_528 ();
 sg13g2_fill_1 FILLER_20_530 ();
 sg13g2_fill_1 FILLER_20_541 ();
 sg13g2_fill_2 FILLER_20_568 ();
 sg13g2_decap_8 FILLER_20_596 ();
 sg13g2_decap_8 FILLER_20_603 ();
 sg13g2_decap_8 FILLER_20_610 ();
 sg13g2_decap_8 FILLER_20_617 ();
 sg13g2_decap_8 FILLER_20_624 ();
 sg13g2_decap_8 FILLER_20_631 ();
 sg13g2_decap_8 FILLER_20_638 ();
 sg13g2_decap_8 FILLER_20_645 ();
 sg13g2_decap_8 FILLER_20_652 ();
 sg13g2_decap_8 FILLER_20_659 ();
 sg13g2_decap_8 FILLER_20_666 ();
 sg13g2_decap_8 FILLER_20_673 ();
 sg13g2_decap_8 FILLER_20_680 ();
 sg13g2_decap_8 FILLER_20_687 ();
 sg13g2_decap_8 FILLER_20_694 ();
 sg13g2_decap_8 FILLER_20_701 ();
 sg13g2_decap_8 FILLER_20_708 ();
 sg13g2_decap_8 FILLER_20_715 ();
 sg13g2_decap_8 FILLER_20_722 ();
 sg13g2_decap_8 FILLER_20_729 ();
 sg13g2_decap_8 FILLER_20_736 ();
 sg13g2_decap_8 FILLER_20_743 ();
 sg13g2_decap_8 FILLER_20_750 ();
 sg13g2_decap_8 FILLER_20_757 ();
 sg13g2_decap_8 FILLER_20_764 ();
 sg13g2_decap_8 FILLER_20_771 ();
 sg13g2_decap_8 FILLER_20_778 ();
 sg13g2_decap_8 FILLER_20_785 ();
 sg13g2_decap_8 FILLER_20_792 ();
 sg13g2_decap_8 FILLER_20_799 ();
 sg13g2_decap_8 FILLER_20_806 ();
 sg13g2_decap_8 FILLER_20_813 ();
 sg13g2_decap_8 FILLER_20_820 ();
 sg13g2_decap_8 FILLER_20_827 ();
 sg13g2_decap_8 FILLER_20_834 ();
 sg13g2_decap_8 FILLER_20_841 ();
 sg13g2_decap_8 FILLER_20_848 ();
 sg13g2_decap_8 FILLER_20_855 ();
 sg13g2_decap_8 FILLER_20_862 ();
 sg13g2_decap_8 FILLER_20_869 ();
 sg13g2_fill_2 FILLER_20_876 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_11 ();
 sg13g2_fill_2 FILLER_21_81 ();
 sg13g2_decap_4 FILLER_21_108 ();
 sg13g2_fill_1 FILLER_21_124 ();
 sg13g2_fill_1 FILLER_21_134 ();
 sg13g2_fill_1 FILLER_21_149 ();
 sg13g2_decap_8 FILLER_21_202 ();
 sg13g2_decap_8 FILLER_21_209 ();
 sg13g2_fill_2 FILLER_21_216 ();
 sg13g2_fill_1 FILLER_21_218 ();
 sg13g2_fill_1 FILLER_21_224 ();
 sg13g2_fill_2 FILLER_21_246 ();
 sg13g2_fill_2 FILLER_21_258 ();
 sg13g2_decap_4 FILLER_21_265 ();
 sg13g2_fill_1 FILLER_21_289 ();
 sg13g2_fill_2 FILLER_21_314 ();
 sg13g2_fill_1 FILLER_21_316 ();
 sg13g2_fill_2 FILLER_21_348 ();
 sg13g2_fill_1 FILLER_21_350 ();
 sg13g2_decap_4 FILLER_21_356 ();
 sg13g2_fill_1 FILLER_21_374 ();
 sg13g2_fill_1 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_415 ();
 sg13g2_fill_1 FILLER_21_423 ();
 sg13g2_fill_2 FILLER_21_432 ();
 sg13g2_fill_2 FILLER_21_441 ();
 sg13g2_fill_1 FILLER_21_443 ();
 sg13g2_fill_2 FILLER_21_449 ();
 sg13g2_fill_1 FILLER_21_451 ();
 sg13g2_fill_1 FILLER_21_465 ();
 sg13g2_fill_2 FILLER_21_501 ();
 sg13g2_fill_1 FILLER_21_513 ();
 sg13g2_fill_2 FILLER_21_527 ();
 sg13g2_decap_4 FILLER_21_575 ();
 sg13g2_decap_8 FILLER_21_583 ();
 sg13g2_decap_8 FILLER_21_590 ();
 sg13g2_decap_8 FILLER_21_597 ();
 sg13g2_decap_8 FILLER_21_604 ();
 sg13g2_decap_8 FILLER_21_611 ();
 sg13g2_decap_8 FILLER_21_618 ();
 sg13g2_decap_8 FILLER_21_625 ();
 sg13g2_decap_8 FILLER_21_632 ();
 sg13g2_decap_8 FILLER_21_639 ();
 sg13g2_decap_8 FILLER_21_646 ();
 sg13g2_decap_8 FILLER_21_653 ();
 sg13g2_decap_8 FILLER_21_660 ();
 sg13g2_decap_8 FILLER_21_667 ();
 sg13g2_decap_8 FILLER_21_674 ();
 sg13g2_decap_8 FILLER_21_681 ();
 sg13g2_decap_8 FILLER_21_688 ();
 sg13g2_decap_8 FILLER_21_695 ();
 sg13g2_decap_8 FILLER_21_702 ();
 sg13g2_decap_8 FILLER_21_709 ();
 sg13g2_decap_8 FILLER_21_716 ();
 sg13g2_decap_8 FILLER_21_723 ();
 sg13g2_decap_8 FILLER_21_730 ();
 sg13g2_decap_8 FILLER_21_737 ();
 sg13g2_decap_8 FILLER_21_744 ();
 sg13g2_decap_8 FILLER_21_751 ();
 sg13g2_decap_8 FILLER_21_758 ();
 sg13g2_decap_8 FILLER_21_765 ();
 sg13g2_decap_8 FILLER_21_772 ();
 sg13g2_decap_8 FILLER_21_779 ();
 sg13g2_decap_8 FILLER_21_786 ();
 sg13g2_decap_8 FILLER_21_793 ();
 sg13g2_decap_8 FILLER_21_800 ();
 sg13g2_decap_8 FILLER_21_807 ();
 sg13g2_decap_8 FILLER_21_814 ();
 sg13g2_decap_8 FILLER_21_821 ();
 sg13g2_decap_8 FILLER_21_828 ();
 sg13g2_decap_8 FILLER_21_835 ();
 sg13g2_decap_8 FILLER_21_842 ();
 sg13g2_decap_8 FILLER_21_849 ();
 sg13g2_decap_8 FILLER_21_856 ();
 sg13g2_decap_8 FILLER_21_863 ();
 sg13g2_decap_8 FILLER_21_870 ();
 sg13g2_fill_1 FILLER_21_877 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_14 ();
 sg13g2_fill_1 FILLER_22_25 ();
 sg13g2_fill_1 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_45 ();
 sg13g2_fill_1 FILLER_22_58 ();
 sg13g2_fill_2 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_78 ();
 sg13g2_fill_2 FILLER_22_83 ();
 sg13g2_fill_2 FILLER_22_93 ();
 sg13g2_fill_1 FILLER_22_95 ();
 sg13g2_fill_2 FILLER_22_122 ();
 sg13g2_fill_1 FILLER_22_124 ();
 sg13g2_decap_4 FILLER_22_151 ();
 sg13g2_decap_4 FILLER_22_173 ();
 sg13g2_fill_1 FILLER_22_177 ();
 sg13g2_decap_4 FILLER_22_182 ();
 sg13g2_fill_2 FILLER_22_190 ();
 sg13g2_fill_1 FILLER_22_192 ();
 sg13g2_fill_1 FILLER_22_243 ();
 sg13g2_fill_2 FILLER_22_249 ();
 sg13g2_decap_4 FILLER_22_262 ();
 sg13g2_fill_1 FILLER_22_266 ();
 sg13g2_fill_2 FILLER_22_306 ();
 sg13g2_fill_2 FILLER_22_339 ();
 sg13g2_fill_1 FILLER_22_367 ();
 sg13g2_fill_2 FILLER_22_373 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_423 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_4 FILLER_22_441 ();
 sg13g2_fill_2 FILLER_22_479 ();
 sg13g2_fill_1 FILLER_22_496 ();
 sg13g2_fill_2 FILLER_22_515 ();
 sg13g2_fill_2 FILLER_22_527 ();
 sg13g2_fill_1 FILLER_22_529 ();
 sg13g2_fill_1 FILLER_22_539 ();
 sg13g2_fill_2 FILLER_22_558 ();
 sg13g2_fill_1 FILLER_22_560 ();
 sg13g2_fill_2 FILLER_22_571 ();
 sg13g2_fill_1 FILLER_22_573 ();
 sg13g2_decap_8 FILLER_22_600 ();
 sg13g2_decap_8 FILLER_22_607 ();
 sg13g2_decap_8 FILLER_22_614 ();
 sg13g2_decap_8 FILLER_22_621 ();
 sg13g2_decap_8 FILLER_22_628 ();
 sg13g2_decap_8 FILLER_22_635 ();
 sg13g2_decap_8 FILLER_22_642 ();
 sg13g2_decap_8 FILLER_22_649 ();
 sg13g2_decap_8 FILLER_22_656 ();
 sg13g2_decap_8 FILLER_22_663 ();
 sg13g2_decap_8 FILLER_22_670 ();
 sg13g2_decap_8 FILLER_22_677 ();
 sg13g2_decap_8 FILLER_22_684 ();
 sg13g2_decap_8 FILLER_22_691 ();
 sg13g2_decap_8 FILLER_22_698 ();
 sg13g2_decap_8 FILLER_22_705 ();
 sg13g2_decap_8 FILLER_22_712 ();
 sg13g2_decap_8 FILLER_22_719 ();
 sg13g2_decap_8 FILLER_22_726 ();
 sg13g2_decap_8 FILLER_22_733 ();
 sg13g2_decap_8 FILLER_22_740 ();
 sg13g2_decap_8 FILLER_22_747 ();
 sg13g2_decap_8 FILLER_22_754 ();
 sg13g2_decap_8 FILLER_22_761 ();
 sg13g2_decap_8 FILLER_22_768 ();
 sg13g2_decap_8 FILLER_22_775 ();
 sg13g2_decap_8 FILLER_22_782 ();
 sg13g2_decap_8 FILLER_22_789 ();
 sg13g2_decap_8 FILLER_22_796 ();
 sg13g2_decap_8 FILLER_22_803 ();
 sg13g2_decap_8 FILLER_22_810 ();
 sg13g2_decap_8 FILLER_22_817 ();
 sg13g2_decap_8 FILLER_22_824 ();
 sg13g2_decap_8 FILLER_22_831 ();
 sg13g2_decap_8 FILLER_22_838 ();
 sg13g2_decap_8 FILLER_22_845 ();
 sg13g2_decap_8 FILLER_22_852 ();
 sg13g2_decap_8 FILLER_22_859 ();
 sg13g2_decap_8 FILLER_22_866 ();
 sg13g2_decap_4 FILLER_22_873 ();
 sg13g2_fill_1 FILLER_22_877 ();
 sg13g2_fill_2 FILLER_23_26 ();
 sg13g2_fill_2 FILLER_23_67 ();
 sg13g2_fill_1 FILLER_23_69 ();
 sg13g2_fill_1 FILLER_23_75 ();
 sg13g2_fill_2 FILLER_23_89 ();
 sg13g2_fill_1 FILLER_23_91 ();
 sg13g2_decap_4 FILLER_23_96 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_4 FILLER_23_133 ();
 sg13g2_fill_1 FILLER_23_137 ();
 sg13g2_fill_1 FILLER_23_153 ();
 sg13g2_fill_1 FILLER_23_159 ();
 sg13g2_fill_1 FILLER_23_170 ();
 sg13g2_fill_1 FILLER_23_197 ();
 sg13g2_fill_1 FILLER_23_224 ();
 sg13g2_fill_2 FILLER_23_230 ();
 sg13g2_fill_1 FILLER_23_240 ();
 sg13g2_fill_2 FILLER_23_251 ();
 sg13g2_fill_1 FILLER_23_253 ();
 sg13g2_fill_2 FILLER_23_271 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_decap_4 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_4 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_368 ();
 sg13g2_fill_1 FILLER_23_387 ();
 sg13g2_fill_1 FILLER_23_397 ();
 sg13g2_fill_2 FILLER_23_467 ();
 sg13g2_fill_2 FILLER_23_514 ();
 sg13g2_fill_2 FILLER_23_526 ();
 sg13g2_fill_2 FILLER_23_554 ();
 sg13g2_fill_2 FILLER_23_582 ();
 sg13g2_fill_1 FILLER_23_584 ();
 sg13g2_decap_8 FILLER_23_589 ();
 sg13g2_decap_8 FILLER_23_596 ();
 sg13g2_decap_8 FILLER_23_603 ();
 sg13g2_decap_8 FILLER_23_610 ();
 sg13g2_decap_8 FILLER_23_617 ();
 sg13g2_decap_8 FILLER_23_624 ();
 sg13g2_decap_8 FILLER_23_631 ();
 sg13g2_decap_8 FILLER_23_638 ();
 sg13g2_decap_8 FILLER_23_645 ();
 sg13g2_decap_8 FILLER_23_652 ();
 sg13g2_decap_8 FILLER_23_659 ();
 sg13g2_decap_8 FILLER_23_666 ();
 sg13g2_decap_8 FILLER_23_673 ();
 sg13g2_decap_8 FILLER_23_680 ();
 sg13g2_decap_8 FILLER_23_687 ();
 sg13g2_decap_8 FILLER_23_694 ();
 sg13g2_decap_8 FILLER_23_701 ();
 sg13g2_decap_8 FILLER_23_708 ();
 sg13g2_decap_8 FILLER_23_715 ();
 sg13g2_decap_8 FILLER_23_722 ();
 sg13g2_decap_8 FILLER_23_729 ();
 sg13g2_decap_8 FILLER_23_736 ();
 sg13g2_decap_8 FILLER_23_743 ();
 sg13g2_decap_8 FILLER_23_750 ();
 sg13g2_decap_8 FILLER_23_757 ();
 sg13g2_decap_8 FILLER_23_764 ();
 sg13g2_decap_8 FILLER_23_771 ();
 sg13g2_decap_8 FILLER_23_778 ();
 sg13g2_decap_8 FILLER_23_785 ();
 sg13g2_decap_8 FILLER_23_792 ();
 sg13g2_decap_8 FILLER_23_799 ();
 sg13g2_decap_8 FILLER_23_806 ();
 sg13g2_decap_8 FILLER_23_813 ();
 sg13g2_decap_8 FILLER_23_820 ();
 sg13g2_decap_8 FILLER_23_827 ();
 sg13g2_decap_8 FILLER_23_834 ();
 sg13g2_decap_8 FILLER_23_841 ();
 sg13g2_decap_8 FILLER_23_848 ();
 sg13g2_decap_8 FILLER_23_855 ();
 sg13g2_decap_8 FILLER_23_862 ();
 sg13g2_decap_8 FILLER_23_869 ();
 sg13g2_fill_2 FILLER_23_876 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_fill_2 FILLER_24_18 ();
 sg13g2_fill_1 FILLER_24_20 ();
 sg13g2_decap_4 FILLER_24_25 ();
 sg13g2_fill_1 FILLER_24_29 ();
 sg13g2_fill_1 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_88 ();
 sg13g2_decap_4 FILLER_24_95 ();
 sg13g2_fill_2 FILLER_24_99 ();
 sg13g2_fill_1 FILLER_24_132 ();
 sg13g2_fill_1 FILLER_24_139 ();
 sg13g2_fill_2 FILLER_24_155 ();
 sg13g2_fill_2 FILLER_24_177 ();
 sg13g2_fill_1 FILLER_24_179 ();
 sg13g2_decap_8 FILLER_24_198 ();
 sg13g2_fill_2 FILLER_24_240 ();
 sg13g2_fill_2 FILLER_24_260 ();
 sg13g2_fill_1 FILLER_24_271 ();
 sg13g2_fill_2 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_320 ();
 sg13g2_fill_2 FILLER_24_327 ();
 sg13g2_fill_1 FILLER_24_333 ();
 sg13g2_fill_1 FILLER_24_344 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_fill_1 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_fill_1 FILLER_24_393 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_2 FILLER_24_439 ();
 sg13g2_fill_1 FILLER_24_455 ();
 sg13g2_fill_1 FILLER_24_498 ();
 sg13g2_decap_4 FILLER_24_529 ();
 sg13g2_fill_1 FILLER_24_533 ();
 sg13g2_fill_1 FILLER_24_542 ();
 sg13g2_decap_4 FILLER_24_557 ();
 sg13g2_fill_2 FILLER_24_561 ();
 sg13g2_decap_8 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_574 ();
 sg13g2_decap_8 FILLER_24_581 ();
 sg13g2_decap_8 FILLER_24_588 ();
 sg13g2_decap_8 FILLER_24_595 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_decap_8 FILLER_24_609 ();
 sg13g2_decap_8 FILLER_24_616 ();
 sg13g2_decap_8 FILLER_24_623 ();
 sg13g2_decap_8 FILLER_24_630 ();
 sg13g2_decap_8 FILLER_24_637 ();
 sg13g2_decap_8 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_651 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_672 ();
 sg13g2_decap_8 FILLER_24_679 ();
 sg13g2_decap_8 FILLER_24_686 ();
 sg13g2_decap_8 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_decap_8 FILLER_24_707 ();
 sg13g2_decap_8 FILLER_24_714 ();
 sg13g2_decap_8 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_728 ();
 sg13g2_decap_8 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_749 ();
 sg13g2_decap_8 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_763 ();
 sg13g2_decap_8 FILLER_24_770 ();
 sg13g2_decap_8 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_8 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_847 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_decap_8 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_24_868 ();
 sg13g2_fill_2 FILLER_24_875 ();
 sg13g2_fill_1 FILLER_24_877 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_64 ();
 sg13g2_fill_1 FILLER_25_70 ();
 sg13g2_fill_1 FILLER_25_96 ();
 sg13g2_fill_1 FILLER_25_118 ();
 sg13g2_fill_1 FILLER_25_140 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_fill_2 FILLER_25_162 ();
 sg13g2_fill_1 FILLER_25_195 ();
 sg13g2_fill_2 FILLER_25_222 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_fill_1 FILLER_25_265 ();
 sg13g2_fill_1 FILLER_25_270 ();
 sg13g2_fill_1 FILLER_25_275 ();
 sg13g2_decap_8 FILLER_25_281 ();
 sg13g2_fill_1 FILLER_25_288 ();
 sg13g2_fill_2 FILLER_25_297 ();
 sg13g2_decap_4 FILLER_25_348 ();
 sg13g2_fill_1 FILLER_25_352 ();
 sg13g2_fill_2 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_fill_1 FILLER_25_397 ();
 sg13g2_fill_2 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_412 ();
 sg13g2_fill_2 FILLER_25_419 ();
 sg13g2_fill_1 FILLER_25_421 ();
 sg13g2_fill_2 FILLER_25_426 ();
 sg13g2_fill_1 FILLER_25_432 ();
 sg13g2_fill_1 FILLER_25_449 ();
 sg13g2_fill_2 FILLER_25_508 ();
 sg13g2_fill_2 FILLER_25_520 ();
 sg13g2_fill_2 FILLER_25_526 ();
 sg13g2_fill_1 FILLER_25_528 ();
 sg13g2_fill_2 FILLER_25_555 ();
 sg13g2_fill_1 FILLER_25_557 ();
 sg13g2_fill_2 FILLER_25_568 ();
 sg13g2_fill_1 FILLER_25_570 ();
 sg13g2_decap_8 FILLER_25_597 ();
 sg13g2_decap_8 FILLER_25_604 ();
 sg13g2_decap_8 FILLER_25_611 ();
 sg13g2_decap_8 FILLER_25_618 ();
 sg13g2_decap_8 FILLER_25_625 ();
 sg13g2_decap_8 FILLER_25_632 ();
 sg13g2_decap_8 FILLER_25_639 ();
 sg13g2_decap_8 FILLER_25_646 ();
 sg13g2_decap_8 FILLER_25_653 ();
 sg13g2_decap_8 FILLER_25_660 ();
 sg13g2_decap_8 FILLER_25_667 ();
 sg13g2_decap_8 FILLER_25_674 ();
 sg13g2_decap_8 FILLER_25_681 ();
 sg13g2_decap_8 FILLER_25_688 ();
 sg13g2_decap_8 FILLER_25_695 ();
 sg13g2_decap_8 FILLER_25_702 ();
 sg13g2_decap_8 FILLER_25_709 ();
 sg13g2_decap_8 FILLER_25_716 ();
 sg13g2_decap_8 FILLER_25_723 ();
 sg13g2_decap_8 FILLER_25_730 ();
 sg13g2_decap_8 FILLER_25_737 ();
 sg13g2_decap_8 FILLER_25_744 ();
 sg13g2_decap_8 FILLER_25_751 ();
 sg13g2_decap_8 FILLER_25_758 ();
 sg13g2_decap_8 FILLER_25_765 ();
 sg13g2_decap_8 FILLER_25_772 ();
 sg13g2_decap_8 FILLER_25_779 ();
 sg13g2_decap_8 FILLER_25_786 ();
 sg13g2_decap_8 FILLER_25_793 ();
 sg13g2_decap_8 FILLER_25_800 ();
 sg13g2_decap_8 FILLER_25_807 ();
 sg13g2_decap_8 FILLER_25_814 ();
 sg13g2_decap_8 FILLER_25_821 ();
 sg13g2_decap_8 FILLER_25_828 ();
 sg13g2_decap_8 FILLER_25_835 ();
 sg13g2_decap_8 FILLER_25_842 ();
 sg13g2_decap_8 FILLER_25_849 ();
 sg13g2_decap_8 FILLER_25_856 ();
 sg13g2_decap_8 FILLER_25_863 ();
 sg13g2_decap_8 FILLER_25_870 ();
 sg13g2_fill_1 FILLER_25_877 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_19 ();
 sg13g2_fill_2 FILLER_26_26 ();
 sg13g2_fill_1 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_33 ();
 sg13g2_decap_4 FILLER_26_39 ();
 sg13g2_fill_1 FILLER_26_43 ();
 sg13g2_decap_4 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_53 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_4 FILLER_26_101 ();
 sg13g2_decap_8 FILLER_26_110 ();
 sg13g2_fill_2 FILLER_26_117 ();
 sg13g2_fill_1 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_156 ();
 sg13g2_fill_2 FILLER_26_162 ();
 sg13g2_fill_2 FILLER_26_169 ();
 sg13g2_fill_1 FILLER_26_171 ();
 sg13g2_fill_2 FILLER_26_193 ();
 sg13g2_decap_4 FILLER_26_199 ();
 sg13g2_decap_4 FILLER_26_207 ();
 sg13g2_fill_2 FILLER_26_216 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_decap_4 FILLER_26_246 ();
 sg13g2_fill_2 FILLER_26_250 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_4 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_decap_4 FILLER_26_283 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_fill_1 FILLER_26_324 ();
 sg13g2_fill_2 FILLER_26_329 ();
 sg13g2_fill_1 FILLER_26_331 ();
 sg13g2_fill_1 FILLER_26_346 ();
 sg13g2_fill_1 FILLER_26_353 ();
 sg13g2_fill_1 FILLER_26_364 ();
 sg13g2_fill_2 FILLER_26_371 ();
 sg13g2_fill_2 FILLER_26_378 ();
 sg13g2_fill_1 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_26_409 ();
 sg13g2_fill_2 FILLER_26_416 ();
 sg13g2_fill_1 FILLER_26_418 ();
 sg13g2_fill_2 FILLER_26_428 ();
 sg13g2_fill_1 FILLER_26_430 ();
 sg13g2_fill_1 FILLER_26_439 ();
 sg13g2_fill_1 FILLER_26_445 ();
 sg13g2_fill_1 FILLER_26_465 ();
 sg13g2_fill_1 FILLER_26_491 ();
 sg13g2_fill_1 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_537 ();
 sg13g2_decap_4 FILLER_26_544 ();
 sg13g2_fill_2 FILLER_26_548 ();
 sg13g2_decap_8 FILLER_26_593 ();
 sg13g2_decap_8 FILLER_26_600 ();
 sg13g2_decap_8 FILLER_26_607 ();
 sg13g2_decap_8 FILLER_26_614 ();
 sg13g2_decap_8 FILLER_26_621 ();
 sg13g2_decap_8 FILLER_26_628 ();
 sg13g2_decap_8 FILLER_26_635 ();
 sg13g2_decap_8 FILLER_26_642 ();
 sg13g2_decap_8 FILLER_26_649 ();
 sg13g2_decap_8 FILLER_26_656 ();
 sg13g2_decap_8 FILLER_26_663 ();
 sg13g2_decap_8 FILLER_26_670 ();
 sg13g2_decap_8 FILLER_26_677 ();
 sg13g2_decap_8 FILLER_26_684 ();
 sg13g2_decap_8 FILLER_26_691 ();
 sg13g2_decap_8 FILLER_26_698 ();
 sg13g2_decap_8 FILLER_26_705 ();
 sg13g2_decap_8 FILLER_26_712 ();
 sg13g2_decap_8 FILLER_26_719 ();
 sg13g2_decap_8 FILLER_26_726 ();
 sg13g2_decap_8 FILLER_26_733 ();
 sg13g2_decap_8 FILLER_26_740 ();
 sg13g2_decap_8 FILLER_26_747 ();
 sg13g2_decap_8 FILLER_26_754 ();
 sg13g2_decap_8 FILLER_26_761 ();
 sg13g2_decap_8 FILLER_26_768 ();
 sg13g2_decap_8 FILLER_26_775 ();
 sg13g2_decap_8 FILLER_26_782 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_796 ();
 sg13g2_decap_8 FILLER_26_803 ();
 sg13g2_decap_8 FILLER_26_810 ();
 sg13g2_decap_8 FILLER_26_817 ();
 sg13g2_decap_8 FILLER_26_824 ();
 sg13g2_decap_8 FILLER_26_831 ();
 sg13g2_decap_8 FILLER_26_838 ();
 sg13g2_decap_8 FILLER_26_845 ();
 sg13g2_decap_8 FILLER_26_852 ();
 sg13g2_decap_8 FILLER_26_859 ();
 sg13g2_decap_8 FILLER_26_866 ();
 sg13g2_decap_4 FILLER_26_873 ();
 sg13g2_fill_1 FILLER_26_877 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_27 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_decap_4 FILLER_27_60 ();
 sg13g2_fill_2 FILLER_27_72 ();
 sg13g2_fill_1 FILLER_27_74 ();
 sg13g2_fill_1 FILLER_27_85 ();
 sg13g2_fill_1 FILLER_27_100 ();
 sg13g2_fill_1 FILLER_27_158 ();
 sg13g2_fill_2 FILLER_27_169 ();
 sg13g2_fill_2 FILLER_27_187 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_2 FILLER_27_249 ();
 sg13g2_fill_1 FILLER_27_288 ();
 sg13g2_decap_8 FILLER_27_293 ();
 sg13g2_decap_4 FILLER_27_300 ();
 sg13g2_fill_1 FILLER_27_312 ();
 sg13g2_fill_1 FILLER_27_330 ();
 sg13g2_fill_1 FILLER_27_338 ();
 sg13g2_fill_1 FILLER_27_345 ();
 sg13g2_fill_2 FILLER_27_350 ();
 sg13g2_fill_2 FILLER_27_394 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_fill_2 FILLER_27_420 ();
 sg13g2_decap_4 FILLER_27_427 ();
 sg13g2_fill_2 FILLER_27_431 ();
 sg13g2_fill_2 FILLER_27_442 ();
 sg13g2_fill_1 FILLER_27_444 ();
 sg13g2_fill_1 FILLER_27_450 ();
 sg13g2_fill_2 FILLER_27_460 ();
 sg13g2_fill_1 FILLER_27_462 ();
 sg13g2_fill_2 FILLER_27_472 ();
 sg13g2_fill_1 FILLER_27_474 ();
 sg13g2_fill_1 FILLER_27_480 ();
 sg13g2_fill_1 FILLER_27_489 ();
 sg13g2_fill_1 FILLER_27_495 ();
 sg13g2_fill_2 FILLER_27_501 ();
 sg13g2_fill_2 FILLER_27_552 ();
 sg13g2_fill_1 FILLER_27_554 ();
 sg13g2_decap_8 FILLER_27_572 ();
 sg13g2_decap_8 FILLER_27_579 ();
 sg13g2_decap_8 FILLER_27_586 ();
 sg13g2_decap_8 FILLER_27_593 ();
 sg13g2_decap_8 FILLER_27_600 ();
 sg13g2_decap_8 FILLER_27_607 ();
 sg13g2_decap_8 FILLER_27_614 ();
 sg13g2_decap_8 FILLER_27_621 ();
 sg13g2_decap_8 FILLER_27_628 ();
 sg13g2_decap_8 FILLER_27_635 ();
 sg13g2_decap_8 FILLER_27_642 ();
 sg13g2_decap_8 FILLER_27_649 ();
 sg13g2_decap_8 FILLER_27_656 ();
 sg13g2_decap_8 FILLER_27_663 ();
 sg13g2_decap_8 FILLER_27_670 ();
 sg13g2_decap_8 FILLER_27_677 ();
 sg13g2_decap_8 FILLER_27_684 ();
 sg13g2_decap_8 FILLER_27_691 ();
 sg13g2_decap_8 FILLER_27_698 ();
 sg13g2_decap_8 FILLER_27_705 ();
 sg13g2_decap_8 FILLER_27_712 ();
 sg13g2_decap_8 FILLER_27_719 ();
 sg13g2_decap_8 FILLER_27_726 ();
 sg13g2_decap_8 FILLER_27_733 ();
 sg13g2_decap_8 FILLER_27_740 ();
 sg13g2_decap_8 FILLER_27_747 ();
 sg13g2_decap_8 FILLER_27_754 ();
 sg13g2_decap_8 FILLER_27_761 ();
 sg13g2_decap_8 FILLER_27_768 ();
 sg13g2_decap_8 FILLER_27_775 ();
 sg13g2_decap_8 FILLER_27_782 ();
 sg13g2_decap_8 FILLER_27_789 ();
 sg13g2_decap_8 FILLER_27_796 ();
 sg13g2_decap_8 FILLER_27_803 ();
 sg13g2_decap_8 FILLER_27_810 ();
 sg13g2_decap_8 FILLER_27_817 ();
 sg13g2_decap_8 FILLER_27_824 ();
 sg13g2_decap_8 FILLER_27_831 ();
 sg13g2_decap_8 FILLER_27_838 ();
 sg13g2_decap_8 FILLER_27_845 ();
 sg13g2_decap_8 FILLER_27_852 ();
 sg13g2_decap_8 FILLER_27_859 ();
 sg13g2_decap_8 FILLER_27_866 ();
 sg13g2_decap_4 FILLER_27_873 ();
 sg13g2_fill_1 FILLER_27_877 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_14 ();
 sg13g2_fill_1 FILLER_28_16 ();
 sg13g2_decap_8 FILLER_28_47 ();
 sg13g2_decap_4 FILLER_28_54 ();
 sg13g2_fill_2 FILLER_28_58 ();
 sg13g2_fill_2 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_81 ();
 sg13g2_fill_2 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_121 ();
 sg13g2_decap_8 FILLER_28_128 ();
 sg13g2_fill_1 FILLER_28_135 ();
 sg13g2_fill_1 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_175 ();
 sg13g2_fill_2 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_194 ();
 sg13g2_decap_8 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_211 ();
 sg13g2_decap_8 FILLER_28_218 ();
 sg13g2_fill_2 FILLER_28_225 ();
 sg13g2_decap_4 FILLER_28_232 ();
 sg13g2_fill_2 FILLER_28_250 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_294 ();
 sg13g2_fill_1 FILLER_28_299 ();
 sg13g2_fill_2 FILLER_28_318 ();
 sg13g2_fill_2 FILLER_28_325 ();
 sg13g2_fill_1 FILLER_28_327 ();
 sg13g2_fill_1 FILLER_28_335 ();
 sg13g2_fill_2 FILLER_28_344 ();
 sg13g2_fill_1 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_391 ();
 sg13g2_fill_1 FILLER_28_398 ();
 sg13g2_fill_1 FILLER_28_410 ();
 sg13g2_fill_2 FILLER_28_435 ();
 sg13g2_fill_1 FILLER_28_437 ();
 sg13g2_decap_4 FILLER_28_443 ();
 sg13g2_fill_1 FILLER_28_447 ();
 sg13g2_fill_1 FILLER_28_453 ();
 sg13g2_decap_8 FILLER_28_459 ();
 sg13g2_decap_4 FILLER_28_466 ();
 sg13g2_fill_2 FILLER_28_501 ();
 sg13g2_fill_2 FILLER_28_508 ();
 sg13g2_fill_1 FILLER_28_510 ();
 sg13g2_decap_8 FILLER_28_515 ();
 sg13g2_decap_8 FILLER_28_522 ();
 sg13g2_fill_2 FILLER_28_529 ();
 sg13g2_fill_1 FILLER_28_531 ();
 sg13g2_decap_8 FILLER_28_545 ();
 sg13g2_fill_2 FILLER_28_552 ();
 sg13g2_fill_1 FILLER_28_554 ();
 sg13g2_decap_8 FILLER_28_563 ();
 sg13g2_decap_8 FILLER_28_570 ();
 sg13g2_decap_8 FILLER_28_577 ();
 sg13g2_decap_8 FILLER_28_584 ();
 sg13g2_decap_8 FILLER_28_591 ();
 sg13g2_decap_8 FILLER_28_598 ();
 sg13g2_decap_8 FILLER_28_605 ();
 sg13g2_decap_8 FILLER_28_612 ();
 sg13g2_decap_8 FILLER_28_619 ();
 sg13g2_decap_8 FILLER_28_626 ();
 sg13g2_decap_8 FILLER_28_633 ();
 sg13g2_decap_8 FILLER_28_640 ();
 sg13g2_decap_8 FILLER_28_647 ();
 sg13g2_decap_8 FILLER_28_654 ();
 sg13g2_decap_8 FILLER_28_661 ();
 sg13g2_decap_8 FILLER_28_668 ();
 sg13g2_decap_8 FILLER_28_675 ();
 sg13g2_decap_8 FILLER_28_682 ();
 sg13g2_decap_8 FILLER_28_689 ();
 sg13g2_decap_8 FILLER_28_696 ();
 sg13g2_decap_8 FILLER_28_703 ();
 sg13g2_decap_8 FILLER_28_710 ();
 sg13g2_decap_8 FILLER_28_717 ();
 sg13g2_decap_8 FILLER_28_724 ();
 sg13g2_decap_8 FILLER_28_731 ();
 sg13g2_decap_8 FILLER_28_738 ();
 sg13g2_decap_8 FILLER_28_745 ();
 sg13g2_decap_8 FILLER_28_752 ();
 sg13g2_decap_8 FILLER_28_759 ();
 sg13g2_decap_8 FILLER_28_766 ();
 sg13g2_decap_8 FILLER_28_773 ();
 sg13g2_decap_8 FILLER_28_780 ();
 sg13g2_decap_8 FILLER_28_787 ();
 sg13g2_decap_8 FILLER_28_794 ();
 sg13g2_decap_8 FILLER_28_801 ();
 sg13g2_decap_8 FILLER_28_808 ();
 sg13g2_decap_8 FILLER_28_815 ();
 sg13g2_decap_8 FILLER_28_822 ();
 sg13g2_decap_8 FILLER_28_829 ();
 sg13g2_decap_8 FILLER_28_836 ();
 sg13g2_decap_8 FILLER_28_843 ();
 sg13g2_decap_8 FILLER_28_850 ();
 sg13g2_decap_8 FILLER_28_857 ();
 sg13g2_decap_8 FILLER_28_864 ();
 sg13g2_decap_8 FILLER_28_871 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_4 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_25 ();
 sg13g2_decap_4 FILLER_29_71 ();
 sg13g2_fill_2 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_167 ();
 sg13g2_decap_4 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_193 ();
 sg13g2_decap_8 FILLER_29_198 ();
 sg13g2_decap_4 FILLER_29_205 ();
 sg13g2_fill_1 FILLER_29_209 ();
 sg13g2_decap_4 FILLER_29_231 ();
 sg13g2_fill_2 FILLER_29_235 ();
 sg13g2_decap_4 FILLER_29_242 ();
 sg13g2_fill_2 FILLER_29_251 ();
 sg13g2_fill_1 FILLER_29_253 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_269 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_282 ();
 sg13g2_fill_1 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_333 ();
 sg13g2_fill_2 FILLER_29_340 ();
 sg13g2_decap_4 FILLER_29_346 ();
 sg13g2_decap_8 FILLER_29_354 ();
 sg13g2_decap_4 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_458 ();
 sg13g2_decap_8 FILLER_29_465 ();
 sg13g2_fill_1 FILLER_29_472 ();
 sg13g2_fill_1 FILLER_29_477 ();
 sg13g2_decap_4 FILLER_29_491 ();
 sg13g2_fill_1 FILLER_29_495 ();
 sg13g2_fill_2 FILLER_29_501 ();
 sg13g2_fill_1 FILLER_29_503 ();
 sg13g2_decap_8 FILLER_29_539 ();
 sg13g2_decap_8 FILLER_29_546 ();
 sg13g2_decap_8 FILLER_29_553 ();
 sg13g2_decap_8 FILLER_29_560 ();
 sg13g2_decap_8 FILLER_29_567 ();
 sg13g2_decap_8 FILLER_29_574 ();
 sg13g2_decap_8 FILLER_29_581 ();
 sg13g2_decap_8 FILLER_29_588 ();
 sg13g2_decap_8 FILLER_29_595 ();
 sg13g2_decap_8 FILLER_29_602 ();
 sg13g2_decap_8 FILLER_29_609 ();
 sg13g2_decap_8 FILLER_29_616 ();
 sg13g2_decap_8 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_630 ();
 sg13g2_decap_8 FILLER_29_637 ();
 sg13g2_decap_8 FILLER_29_644 ();
 sg13g2_decap_8 FILLER_29_651 ();
 sg13g2_decap_8 FILLER_29_658 ();
 sg13g2_decap_8 FILLER_29_665 ();
 sg13g2_decap_8 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_679 ();
 sg13g2_decap_8 FILLER_29_686 ();
 sg13g2_decap_8 FILLER_29_693 ();
 sg13g2_decap_8 FILLER_29_700 ();
 sg13g2_decap_8 FILLER_29_707 ();
 sg13g2_decap_8 FILLER_29_714 ();
 sg13g2_decap_8 FILLER_29_721 ();
 sg13g2_decap_8 FILLER_29_728 ();
 sg13g2_decap_8 FILLER_29_735 ();
 sg13g2_decap_8 FILLER_29_742 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_8 FILLER_29_756 ();
 sg13g2_decap_8 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_770 ();
 sg13g2_decap_8 FILLER_29_777 ();
 sg13g2_decap_8 FILLER_29_784 ();
 sg13g2_decap_8 FILLER_29_791 ();
 sg13g2_decap_8 FILLER_29_798 ();
 sg13g2_decap_8 FILLER_29_805 ();
 sg13g2_decap_8 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_819 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_decap_8 FILLER_29_847 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_decap_8 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_29_868 ();
 sg13g2_fill_2 FILLER_29_875 ();
 sg13g2_fill_1 FILLER_29_877 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_23 ();
 sg13g2_fill_2 FILLER_30_50 ();
 sg13g2_decap_4 FILLER_30_86 ();
 sg13g2_decap_8 FILLER_30_115 ();
 sg13g2_fill_1 FILLER_30_122 ();
 sg13g2_decap_8 FILLER_30_146 ();
 sg13g2_fill_2 FILLER_30_153 ();
 sg13g2_fill_2 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_178 ();
 sg13g2_decap_4 FILLER_30_214 ();
 sg13g2_fill_2 FILLER_30_218 ();
 sg13g2_fill_2 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_277 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_305 ();
 sg13g2_fill_1 FILLER_30_315 ();
 sg13g2_fill_2 FILLER_30_355 ();
 sg13g2_fill_2 FILLER_30_362 ();
 sg13g2_fill_1 FILLER_30_364 ();
 sg13g2_fill_1 FILLER_30_368 ();
 sg13g2_fill_1 FILLER_30_377 ();
 sg13g2_fill_1 FILLER_30_390 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_417 ();
 sg13g2_decap_4 FILLER_30_429 ();
 sg13g2_fill_2 FILLER_30_433 ();
 sg13g2_fill_1 FILLER_30_447 ();
 sg13g2_decap_8 FILLER_30_484 ();
 sg13g2_fill_2 FILLER_30_498 ();
 sg13g2_decap_8 FILLER_30_521 ();
 sg13g2_decap_8 FILLER_30_528 ();
 sg13g2_decap_4 FILLER_30_535 ();
 sg13g2_fill_1 FILLER_30_539 ();
 sg13g2_decap_8 FILLER_30_553 ();
 sg13g2_decap_8 FILLER_30_560 ();
 sg13g2_decap_8 FILLER_30_567 ();
 sg13g2_decap_8 FILLER_30_574 ();
 sg13g2_decap_8 FILLER_30_581 ();
 sg13g2_decap_8 FILLER_30_588 ();
 sg13g2_decap_8 FILLER_30_595 ();
 sg13g2_decap_8 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_8 FILLER_30_616 ();
 sg13g2_decap_8 FILLER_30_623 ();
 sg13g2_decap_8 FILLER_30_630 ();
 sg13g2_decap_8 FILLER_30_637 ();
 sg13g2_decap_8 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_8 FILLER_30_658 ();
 sg13g2_decap_8 FILLER_30_665 ();
 sg13g2_decap_8 FILLER_30_672 ();
 sg13g2_decap_8 FILLER_30_679 ();
 sg13g2_decap_8 FILLER_30_686 ();
 sg13g2_decap_8 FILLER_30_693 ();
 sg13g2_decap_8 FILLER_30_700 ();
 sg13g2_decap_8 FILLER_30_707 ();
 sg13g2_decap_8 FILLER_30_714 ();
 sg13g2_decap_8 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_742 ();
 sg13g2_decap_8 FILLER_30_749 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_decap_8 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_30_868 ();
 sg13g2_fill_2 FILLER_30_875 ();
 sg13g2_fill_1 FILLER_30_877 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_4 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_36 ();
 sg13g2_decap_8 FILLER_31_43 ();
 sg13g2_decap_8 FILLER_31_50 ();
 sg13g2_decap_4 FILLER_31_57 ();
 sg13g2_fill_1 FILLER_31_61 ();
 sg13g2_fill_1 FILLER_31_66 ();
 sg13g2_decap_4 FILLER_31_71 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_fill_2 FILLER_31_90 ();
 sg13g2_fill_1 FILLER_31_92 ();
 sg13g2_fill_2 FILLER_31_105 ();
 sg13g2_fill_1 FILLER_31_107 ();
 sg13g2_decap_8 FILLER_31_117 ();
 sg13g2_fill_2 FILLER_31_124 ();
 sg13g2_decap_4 FILLER_31_152 ();
 sg13g2_decap_8 FILLER_31_160 ();
 sg13g2_decap_8 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_174 ();
 sg13g2_fill_1 FILLER_31_176 ();
 sg13g2_decap_8 FILLER_31_186 ();
 sg13g2_decap_4 FILLER_31_193 ();
 sg13g2_fill_2 FILLER_31_197 ();
 sg13g2_fill_1 FILLER_31_225 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_312 ();
 sg13g2_fill_1 FILLER_31_314 ();
 sg13g2_decap_4 FILLER_31_341 ();
 sg13g2_fill_1 FILLER_31_345 ();
 sg13g2_fill_1 FILLER_31_361 ();
 sg13g2_fill_2 FILLER_31_389 ();
 sg13g2_fill_2 FILLER_31_403 ();
 sg13g2_fill_1 FILLER_31_410 ();
 sg13g2_fill_1 FILLER_31_469 ();
 sg13g2_fill_1 FILLER_31_484 ();
 sg13g2_fill_2 FILLER_31_517 ();
 sg13g2_decap_8 FILLER_31_524 ();
 sg13g2_fill_1 FILLER_31_531 ();
 sg13g2_decap_8 FILLER_31_544 ();
 sg13g2_decap_8 FILLER_31_551 ();
 sg13g2_decap_8 FILLER_31_558 ();
 sg13g2_decap_8 FILLER_31_565 ();
 sg13g2_decap_8 FILLER_31_572 ();
 sg13g2_decap_8 FILLER_31_579 ();
 sg13g2_decap_8 FILLER_31_586 ();
 sg13g2_decap_8 FILLER_31_593 ();
 sg13g2_decap_8 FILLER_31_600 ();
 sg13g2_decap_8 FILLER_31_607 ();
 sg13g2_decap_8 FILLER_31_614 ();
 sg13g2_decap_8 FILLER_31_621 ();
 sg13g2_decap_8 FILLER_31_628 ();
 sg13g2_decap_8 FILLER_31_635 ();
 sg13g2_decap_8 FILLER_31_642 ();
 sg13g2_decap_8 FILLER_31_649 ();
 sg13g2_decap_8 FILLER_31_656 ();
 sg13g2_fill_1 FILLER_31_663 ();
 sg13g2_decap_8 FILLER_31_701 ();
 sg13g2_decap_8 FILLER_31_725 ();
 sg13g2_decap_8 FILLER_31_732 ();
 sg13g2_decap_8 FILLER_31_739 ();
 sg13g2_decap_8 FILLER_31_746 ();
 sg13g2_decap_8 FILLER_31_753 ();
 sg13g2_decap_8 FILLER_31_760 ();
 sg13g2_decap_8 FILLER_31_767 ();
 sg13g2_decap_8 FILLER_31_774 ();
 sg13g2_decap_8 FILLER_31_781 ();
 sg13g2_decap_8 FILLER_31_788 ();
 sg13g2_decap_8 FILLER_31_795 ();
 sg13g2_decap_8 FILLER_31_802 ();
 sg13g2_decap_8 FILLER_31_809 ();
 sg13g2_decap_8 FILLER_31_816 ();
 sg13g2_decap_8 FILLER_31_823 ();
 sg13g2_decap_8 FILLER_31_830 ();
 sg13g2_decap_8 FILLER_31_837 ();
 sg13g2_decap_8 FILLER_31_844 ();
 sg13g2_decap_8 FILLER_31_851 ();
 sg13g2_decap_8 FILLER_31_858 ();
 sg13g2_decap_8 FILLER_31_865 ();
 sg13g2_decap_4 FILLER_31_872 ();
 sg13g2_fill_2 FILLER_31_876 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_4 FILLER_32_56 ();
 sg13g2_fill_2 FILLER_32_86 ();
 sg13g2_fill_2 FILLER_32_114 ();
 sg13g2_fill_1 FILLER_32_116 ();
 sg13g2_fill_1 FILLER_32_147 ();
 sg13g2_fill_1 FILLER_32_174 ();
 sg13g2_fill_1 FILLER_32_206 ();
 sg13g2_fill_2 FILLER_32_257 ();
 sg13g2_fill_1 FILLER_32_259 ();
 sg13g2_fill_2 FILLER_32_274 ();
 sg13g2_fill_1 FILLER_32_276 ();
 sg13g2_fill_1 FILLER_32_281 ();
 sg13g2_fill_1 FILLER_32_287 ();
 sg13g2_fill_2 FILLER_32_303 ();
 sg13g2_decap_4 FILLER_32_312 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_fill_2 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_373 ();
 sg13g2_decap_8 FILLER_32_380 ();
 sg13g2_fill_2 FILLER_32_387 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_fill_1 FILLER_32_400 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_fill_2 FILLER_32_414 ();
 sg13g2_fill_2 FILLER_32_448 ();
 sg13g2_fill_1 FILLER_32_450 ();
 sg13g2_fill_2 FILLER_32_471 ();
 sg13g2_fill_2 FILLER_32_490 ();
 sg13g2_fill_1 FILLER_32_497 ();
 sg13g2_decap_4 FILLER_32_526 ();
 sg13g2_fill_1 FILLER_32_535 ();
 sg13g2_decap_8 FILLER_32_549 ();
 sg13g2_decap_8 FILLER_32_556 ();
 sg13g2_decap_8 FILLER_32_563 ();
 sg13g2_decap_8 FILLER_32_570 ();
 sg13g2_decap_8 FILLER_32_577 ();
 sg13g2_decap_8 FILLER_32_584 ();
 sg13g2_decap_8 FILLER_32_595 ();
 sg13g2_fill_1 FILLER_32_602 ();
 sg13g2_decap_8 FILLER_32_608 ();
 sg13g2_fill_1 FILLER_32_615 ();
 sg13g2_fill_1 FILLER_32_620 ();
 sg13g2_decap_8 FILLER_32_651 ();
 sg13g2_decap_8 FILLER_32_658 ();
 sg13g2_fill_1 FILLER_32_665 ();
 sg13g2_decap_4 FILLER_32_669 ();
 sg13g2_fill_2 FILLER_32_682 ();
 sg13g2_fill_1 FILLER_32_684 ();
 sg13g2_fill_1 FILLER_32_690 ();
 sg13g2_decap_8 FILLER_32_695 ();
 sg13g2_fill_1 FILLER_32_702 ();
 sg13g2_fill_2 FILLER_32_727 ();
 sg13g2_decap_4 FILLER_32_733 ();
 sg13g2_fill_2 FILLER_32_746 ();
 sg13g2_fill_1 FILLER_32_748 ();
 sg13g2_fill_2 FILLER_32_761 ();
 sg13g2_fill_1 FILLER_32_763 ();
 sg13g2_decap_8 FILLER_32_768 ();
 sg13g2_decap_8 FILLER_32_775 ();
 sg13g2_decap_8 FILLER_32_782 ();
 sg13g2_decap_8 FILLER_32_789 ();
 sg13g2_decap_8 FILLER_32_796 ();
 sg13g2_decap_8 FILLER_32_803 ();
 sg13g2_decap_8 FILLER_32_810 ();
 sg13g2_decap_8 FILLER_32_817 ();
 sg13g2_decap_8 FILLER_32_824 ();
 sg13g2_decap_8 FILLER_32_831 ();
 sg13g2_decap_8 FILLER_32_838 ();
 sg13g2_decap_8 FILLER_32_845 ();
 sg13g2_decap_8 FILLER_32_852 ();
 sg13g2_decap_8 FILLER_32_859 ();
 sg13g2_decap_8 FILLER_32_866 ();
 sg13g2_decap_4 FILLER_32_873 ();
 sg13g2_fill_1 FILLER_32_877 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_4 FILLER_33_49 ();
 sg13g2_decap_4 FILLER_33_88 ();
 sg13g2_decap_8 FILLER_33_96 ();
 sg13g2_fill_2 FILLER_33_113 ();
 sg13g2_fill_2 FILLER_33_120 ();
 sg13g2_fill_1 FILLER_33_122 ();
 sg13g2_fill_2 FILLER_33_127 ();
 sg13g2_fill_1 FILLER_33_129 ();
 sg13g2_fill_2 FILLER_33_140 ();
 sg13g2_fill_1 FILLER_33_142 ();
 sg13g2_fill_1 FILLER_33_185 ();
 sg13g2_decap_4 FILLER_33_190 ();
 sg13g2_fill_1 FILLER_33_194 ();
 sg13g2_fill_2 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_decap_8 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_268 ();
 sg13g2_fill_2 FILLER_33_275 ();
 sg13g2_fill_2 FILLER_33_286 ();
 sg13g2_fill_1 FILLER_33_308 ();
 sg13g2_fill_2 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_328 ();
 sg13g2_fill_2 FILLER_33_334 ();
 sg13g2_fill_1 FILLER_33_336 ();
 sg13g2_fill_2 FILLER_33_376 ();
 sg13g2_fill_1 FILLER_33_378 ();
 sg13g2_decap_4 FILLER_33_383 ();
 sg13g2_fill_1 FILLER_33_416 ();
 sg13g2_fill_2 FILLER_33_430 ();
 sg13g2_fill_1 FILLER_33_432 ();
 sg13g2_decap_8 FILLER_33_464 ();
 sg13g2_fill_2 FILLER_33_471 ();
 sg13g2_decap_8 FILLER_33_477 ();
 sg13g2_fill_1 FILLER_33_484 ();
 sg13g2_fill_2 FILLER_33_490 ();
 sg13g2_fill_1 FILLER_33_513 ();
 sg13g2_fill_1 FILLER_33_529 ();
 sg13g2_decap_4 FILLER_33_547 ();
 sg13g2_fill_1 FILLER_33_564 ();
 sg13g2_fill_1 FILLER_33_569 ();
 sg13g2_decap_4 FILLER_33_578 ();
 sg13g2_fill_2 FILLER_33_582 ();
 sg13g2_fill_2 FILLER_33_615 ();
 sg13g2_fill_1 FILLER_33_617 ();
 sg13g2_fill_1 FILLER_33_622 ();
 sg13g2_decap_4 FILLER_33_627 ();
 sg13g2_fill_1 FILLER_33_631 ();
 sg13g2_decap_4 FILLER_33_636 ();
 sg13g2_fill_2 FILLER_33_645 ();
 sg13g2_fill_1 FILLER_33_651 ();
 sg13g2_fill_2 FILLER_33_660 ();
 sg13g2_fill_1 FILLER_33_667 ();
 sg13g2_fill_1 FILLER_33_681 ();
 sg13g2_decap_8 FILLER_33_698 ();
 sg13g2_fill_2 FILLER_33_710 ();
 sg13g2_fill_2 FILLER_33_739 ();
 sg13g2_fill_1 FILLER_33_741 ();
 sg13g2_decap_8 FILLER_33_789 ();
 sg13g2_decap_8 FILLER_33_796 ();
 sg13g2_decap_8 FILLER_33_803 ();
 sg13g2_decap_8 FILLER_33_810 ();
 sg13g2_decap_8 FILLER_33_817 ();
 sg13g2_decap_8 FILLER_33_824 ();
 sg13g2_decap_8 FILLER_33_831 ();
 sg13g2_decap_8 FILLER_33_838 ();
 sg13g2_decap_8 FILLER_33_845 ();
 sg13g2_decap_8 FILLER_33_852 ();
 sg13g2_decap_8 FILLER_33_859 ();
 sg13g2_decap_8 FILLER_33_866 ();
 sg13g2_decap_4 FILLER_33_873 ();
 sg13g2_fill_1 FILLER_33_877 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_fill_2 FILLER_34_63 ();
 sg13g2_decap_4 FILLER_34_69 ();
 sg13g2_fill_1 FILLER_34_73 ();
 sg13g2_fill_2 FILLER_34_83 ();
 sg13g2_fill_2 FILLER_34_111 ();
 sg13g2_fill_2 FILLER_34_118 ();
 sg13g2_fill_1 FILLER_34_120 ();
 sg13g2_fill_2 FILLER_34_157 ();
 sg13g2_decap_4 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_218 ();
 sg13g2_fill_2 FILLER_34_224 ();
 sg13g2_fill_1 FILLER_34_252 ();
 sg13g2_fill_2 FILLER_34_258 ();
 sg13g2_fill_2 FILLER_34_286 ();
 sg13g2_fill_1 FILLER_34_288 ();
 sg13g2_fill_1 FILLER_34_299 ();
 sg13g2_fill_1 FILLER_34_337 ();
 sg13g2_decap_8 FILLER_34_342 ();
 sg13g2_decap_4 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_fill_2 FILLER_34_384 ();
 sg13g2_fill_1 FILLER_34_386 ();
 sg13g2_fill_2 FILLER_34_391 ();
 sg13g2_fill_1 FILLER_34_415 ();
 sg13g2_fill_2 FILLER_34_420 ();
 sg13g2_fill_1 FILLER_34_448 ();
 sg13g2_decap_8 FILLER_34_453 ();
 sg13g2_decap_4 FILLER_34_460 ();
 sg13g2_fill_1 FILLER_34_464 ();
 sg13g2_fill_1 FILLER_34_481 ();
 sg13g2_decap_8 FILLER_34_504 ();
 sg13g2_decap_4 FILLER_34_511 ();
 sg13g2_decap_8 FILLER_34_543 ();
 sg13g2_decap_8 FILLER_34_550 ();
 sg13g2_fill_1 FILLER_34_557 ();
 sg13g2_fill_2 FILLER_34_613 ();
 sg13g2_fill_1 FILLER_34_615 ();
 sg13g2_fill_2 FILLER_34_660 ();
 sg13g2_fill_1 FILLER_34_662 ();
 sg13g2_fill_2 FILLER_34_687 ();
 sg13g2_fill_1 FILLER_34_693 ();
 sg13g2_fill_2 FILLER_34_705 ();
 sg13g2_fill_2 FILLER_34_712 ();
 sg13g2_fill_1 FILLER_34_714 ();
 sg13g2_fill_1 FILLER_34_723 ();
 sg13g2_fill_2 FILLER_34_732 ();
 sg13g2_fill_1 FILLER_34_734 ();
 sg13g2_fill_1 FILLER_34_748 ();
 sg13g2_fill_2 FILLER_34_759 ();
 sg13g2_fill_1 FILLER_34_765 ();
 sg13g2_decap_8 FILLER_34_794 ();
 sg13g2_decap_8 FILLER_34_801 ();
 sg13g2_decap_8 FILLER_34_808 ();
 sg13g2_decap_8 FILLER_34_815 ();
 sg13g2_decap_8 FILLER_34_822 ();
 sg13g2_decap_8 FILLER_34_829 ();
 sg13g2_decap_8 FILLER_34_836 ();
 sg13g2_decap_8 FILLER_34_843 ();
 sg13g2_decap_8 FILLER_34_850 ();
 sg13g2_decap_8 FILLER_34_857 ();
 sg13g2_decap_8 FILLER_34_864 ();
 sg13g2_decap_8 FILLER_34_871 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_fill_1 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_120 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_fill_1 FILLER_35_137 ();
 sg13g2_fill_1 FILLER_35_142 ();
 sg13g2_fill_1 FILLER_35_153 ();
 sg13g2_fill_2 FILLER_35_161 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_fill_2 FILLER_35_200 ();
 sg13g2_fill_1 FILLER_35_228 ();
 sg13g2_fill_2 FILLER_35_233 ();
 sg13g2_fill_1 FILLER_35_265 ();
 sg13g2_fill_2 FILLER_35_274 ();
 sg13g2_fill_1 FILLER_35_281 ();
 sg13g2_fill_2 FILLER_35_286 ();
 sg13g2_fill_1 FILLER_35_296 ();
 sg13g2_fill_2 FILLER_35_323 ();
 sg13g2_fill_2 FILLER_35_334 ();
 sg13g2_fill_2 FILLER_35_346 ();
 sg13g2_fill_1 FILLER_35_348 ();
 sg13g2_fill_2 FILLER_35_364 ();
 sg13g2_fill_1 FILLER_35_366 ();
 sg13g2_fill_1 FILLER_35_387 ();
 sg13g2_decap_4 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_fill_1 FILLER_35_413 ();
 sg13g2_fill_1 FILLER_35_418 ();
 sg13g2_fill_1 FILLER_35_423 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_fill_1 FILLER_35_438 ();
 sg13g2_fill_2 FILLER_35_452 ();
 sg13g2_decap_8 FILLER_35_458 ();
 sg13g2_fill_2 FILLER_35_514 ();
 sg13g2_fill_1 FILLER_35_521 ();
 sg13g2_fill_1 FILLER_35_530 ();
 sg13g2_fill_2 FILLER_35_564 ();
 sg13g2_decap_4 FILLER_35_570 ();
 sg13g2_fill_2 FILLER_35_574 ();
 sg13g2_fill_2 FILLER_35_586 ();
 sg13g2_fill_1 FILLER_35_588 ();
 sg13g2_fill_1 FILLER_35_615 ();
 sg13g2_decap_4 FILLER_35_646 ();
 sg13g2_fill_2 FILLER_35_650 ();
 sg13g2_fill_1 FILLER_35_694 ();
 sg13g2_fill_2 FILLER_35_699 ();
 sg13g2_fill_1 FILLER_35_705 ();
 sg13g2_fill_1 FILLER_35_711 ();
 sg13g2_fill_1 FILLER_35_716 ();
 sg13g2_fill_1 FILLER_35_745 ();
 sg13g2_decap_8 FILLER_35_762 ();
 sg13g2_fill_1 FILLER_35_769 ();
 sg13g2_fill_1 FILLER_35_782 ();
 sg13g2_decap_8 FILLER_35_787 ();
 sg13g2_decap_8 FILLER_35_794 ();
 sg13g2_decap_8 FILLER_35_801 ();
 sg13g2_decap_8 FILLER_35_808 ();
 sg13g2_decap_8 FILLER_35_815 ();
 sg13g2_decap_8 FILLER_35_822 ();
 sg13g2_decap_8 FILLER_35_829 ();
 sg13g2_decap_8 FILLER_35_836 ();
 sg13g2_decap_8 FILLER_35_843 ();
 sg13g2_decap_8 FILLER_35_850 ();
 sg13g2_decap_8 FILLER_35_857 ();
 sg13g2_decap_8 FILLER_35_864 ();
 sg13g2_decap_8 FILLER_35_871 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_4 FILLER_36_133 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_decap_8 FILLER_36_164 ();
 sg13g2_decap_8 FILLER_36_171 ();
 sg13g2_fill_2 FILLER_36_178 ();
 sg13g2_decap_8 FILLER_36_184 ();
 sg13g2_decap_4 FILLER_36_191 ();
 sg13g2_fill_1 FILLER_36_195 ();
 sg13g2_decap_8 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_208 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_237 ();
 sg13g2_fill_1 FILLER_36_239 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_fill_1 FILLER_36_252 ();
 sg13g2_fill_1 FILLER_36_261 ();
 sg13g2_decap_4 FILLER_36_270 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_4 FILLER_36_329 ();
 sg13g2_fill_1 FILLER_36_361 ();
 sg13g2_decap_8 FILLER_36_389 ();
 sg13g2_fill_1 FILLER_36_396 ();
 sg13g2_fill_1 FILLER_36_403 ();
 sg13g2_fill_1 FILLER_36_409 ();
 sg13g2_fill_1 FILLER_36_417 ();
 sg13g2_fill_1 FILLER_36_427 ();
 sg13g2_fill_2 FILLER_36_432 ();
 sg13g2_fill_2 FILLER_36_470 ();
 sg13g2_fill_1 FILLER_36_472 ();
 sg13g2_fill_1 FILLER_36_512 ();
 sg13g2_fill_1 FILLER_36_517 ();
 sg13g2_fill_1 FILLER_36_523 ();
 sg13g2_fill_2 FILLER_36_541 ();
 sg13g2_fill_1 FILLER_36_548 ();
 sg13g2_decap_4 FILLER_36_563 ();
 sg13g2_fill_1 FILLER_36_571 ();
 sg13g2_fill_1 FILLER_36_581 ();
 sg13g2_fill_1 FILLER_36_591 ();
 sg13g2_fill_1 FILLER_36_597 ();
 sg13g2_fill_2 FILLER_36_633 ();
 sg13g2_fill_1 FILLER_36_635 ();
 sg13g2_decap_4 FILLER_36_640 ();
 sg13g2_decap_4 FILLER_36_648 ();
 sg13g2_fill_1 FILLER_36_652 ();
 sg13g2_fill_1 FILLER_36_679 ();
 sg13g2_fill_1 FILLER_36_691 ();
 sg13g2_fill_1 FILLER_36_711 ();
 sg13g2_fill_2 FILLER_36_734 ();
 sg13g2_fill_1 FILLER_36_736 ();
 sg13g2_fill_1 FILLER_36_759 ();
 sg13g2_fill_2 FILLER_36_764 ();
 sg13g2_fill_1 FILLER_36_779 ();
 sg13g2_decap_8 FILLER_36_788 ();
 sg13g2_decap_8 FILLER_36_795 ();
 sg13g2_decap_4 FILLER_36_802 ();
 sg13g2_fill_1 FILLER_36_806 ();
 sg13g2_decap_8 FILLER_36_810 ();
 sg13g2_decap_8 FILLER_36_817 ();
 sg13g2_decap_8 FILLER_36_824 ();
 sg13g2_decap_8 FILLER_36_831 ();
 sg13g2_decap_8 FILLER_36_838 ();
 sg13g2_decap_8 FILLER_36_845 ();
 sg13g2_decap_8 FILLER_36_852 ();
 sg13g2_decap_8 FILLER_36_859 ();
 sg13g2_decap_8 FILLER_36_866 ();
 sg13g2_decap_4 FILLER_36_873 ();
 sg13g2_fill_1 FILLER_36_877 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_116 ();
 sg13g2_decap_8 FILLER_37_123 ();
 sg13g2_decap_8 FILLER_37_130 ();
 sg13g2_decap_8 FILLER_37_137 ();
 sg13g2_fill_2 FILLER_37_144 ();
 sg13g2_decap_8 FILLER_37_150 ();
 sg13g2_decap_8 FILLER_37_157 ();
 sg13g2_decap_8 FILLER_37_164 ();
 sg13g2_decap_4 FILLER_37_171 ();
 sg13g2_fill_2 FILLER_37_175 ();
 sg13g2_fill_1 FILLER_37_207 ();
 sg13g2_fill_2 FILLER_37_243 ();
 sg13g2_fill_1 FILLER_37_245 ();
 sg13g2_fill_2 FILLER_37_259 ();
 sg13g2_fill_2 FILLER_37_275 ();
 sg13g2_fill_2 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_decap_4 FILLER_37_333 ();
 sg13g2_fill_2 FILLER_37_353 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_fill_1 FILLER_37_376 ();
 sg13g2_fill_2 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_fill_2 FILLER_37_435 ();
 sg13g2_fill_1 FILLER_37_437 ();
 sg13g2_fill_1 FILLER_37_451 ();
 sg13g2_decap_4 FILLER_37_456 ();
 sg13g2_fill_1 FILLER_37_460 ();
 sg13g2_fill_2 FILLER_37_479 ();
 sg13g2_fill_1 FILLER_37_485 ();
 sg13g2_fill_1 FILLER_37_494 ();
 sg13g2_fill_2 FILLER_37_521 ();
 sg13g2_fill_1 FILLER_37_549 ();
 sg13g2_decap_8 FILLER_37_581 ();
 sg13g2_fill_1 FILLER_37_597 ();
 sg13g2_decap_4 FILLER_37_603 ();
 sg13g2_fill_1 FILLER_37_611 ();
 sg13g2_fill_2 FILLER_37_630 ();
 sg13g2_fill_1 FILLER_37_632 ();
 sg13g2_fill_1 FILLER_37_641 ();
 sg13g2_fill_1 FILLER_37_683 ();
 sg13g2_fill_2 FILLER_37_706 ();
 sg13g2_fill_2 FILLER_37_722 ();
 sg13g2_decap_4 FILLER_37_782 ();
 sg13g2_fill_1 FILLER_37_794 ();
 sg13g2_fill_2 FILLER_37_818 ();
 sg13g2_fill_1 FILLER_37_825 ();
 sg13g2_decap_8 FILLER_37_831 ();
 sg13g2_decap_8 FILLER_37_838 ();
 sg13g2_decap_8 FILLER_37_845 ();
 sg13g2_decap_8 FILLER_37_852 ();
 sg13g2_decap_8 FILLER_37_859 ();
 sg13g2_decap_8 FILLER_37_866 ();
 sg13g2_decap_4 FILLER_37_873 ();
 sg13g2_fill_1 FILLER_37_877 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_4 FILLER_38_120 ();
 sg13g2_fill_2 FILLER_38_124 ();
 sg13g2_fill_1 FILLER_38_186 ();
 sg13g2_fill_2 FILLER_38_217 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_decap_4 FILLER_38_237 ();
 sg13g2_fill_2 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_293 ();
 sg13g2_decap_8 FILLER_38_299 ();
 sg13g2_fill_2 FILLER_38_306 ();
 sg13g2_fill_2 FILLER_38_322 ();
 sg13g2_decap_4 FILLER_38_329 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_fill_2 FILLER_38_349 ();
 sg13g2_fill_1 FILLER_38_351 ();
 sg13g2_fill_2 FILLER_38_362 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_fill_2 FILLER_38_379 ();
 sg13g2_fill_1 FILLER_38_381 ();
 sg13g2_decap_4 FILLER_38_387 ();
 sg13g2_fill_2 FILLER_38_422 ();
 sg13g2_fill_1 FILLER_38_427 ();
 sg13g2_decap_8 FILLER_38_432 ();
 sg13g2_fill_2 FILLER_38_439 ();
 sg13g2_decap_8 FILLER_38_453 ();
 sg13g2_fill_2 FILLER_38_460 ();
 sg13g2_fill_2 FILLER_38_474 ();
 sg13g2_fill_1 FILLER_38_497 ();
 sg13g2_fill_1 FILLER_38_524 ();
 sg13g2_decap_4 FILLER_38_530 ();
 sg13g2_fill_1 FILLER_38_534 ();
 sg13g2_decap_4 FILLER_38_540 ();
 sg13g2_fill_1 FILLER_38_544 ();
 sg13g2_decap_4 FILLER_38_563 ();
 sg13g2_fill_2 FILLER_38_567 ();
 sg13g2_decap_4 FILLER_38_574 ();
 sg13g2_fill_1 FILLER_38_598 ();
 sg13g2_fill_2 FILLER_38_603 ();
 sg13g2_fill_2 FILLER_38_610 ();
 sg13g2_fill_2 FILLER_38_617 ();
 sg13g2_fill_2 FILLER_38_675 ();
 sg13g2_decap_4 FILLER_38_681 ();
 sg13g2_fill_1 FILLER_38_685 ();
 sg13g2_fill_2 FILLER_38_714 ();
 sg13g2_decap_4 FILLER_38_731 ();
 sg13g2_fill_2 FILLER_38_780 ();
 sg13g2_decap_4 FILLER_38_792 ();
 sg13g2_fill_1 FILLER_38_796 ();
 sg13g2_decap_8 FILLER_38_844 ();
 sg13g2_decap_8 FILLER_38_851 ();
 sg13g2_decap_8 FILLER_38_858 ();
 sg13g2_decap_8 FILLER_38_865 ();
 sg13g2_decap_4 FILLER_38_872 ();
 sg13g2_fill_2 FILLER_38_876 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_4 FILLER_39_98 ();
 sg13g2_fill_1 FILLER_39_102 ();
 sg13g2_decap_4 FILLER_39_129 ();
 sg13g2_decap_4 FILLER_39_137 ();
 sg13g2_decap_4 FILLER_39_179 ();
 sg13g2_fill_2 FILLER_39_183 ();
 sg13g2_decap_4 FILLER_39_203 ();
 sg13g2_fill_1 FILLER_39_211 ();
 sg13g2_fill_2 FILLER_39_216 ();
 sg13g2_decap_4 FILLER_39_249 ();
 sg13g2_decap_4 FILLER_39_288 ();
 sg13g2_decap_8 FILLER_39_344 ();
 sg13g2_decap_8 FILLER_39_351 ();
 sg13g2_fill_2 FILLER_39_368 ();
 sg13g2_fill_1 FILLER_39_409 ();
 sg13g2_fill_1 FILLER_39_472 ();
 sg13g2_fill_1 FILLER_39_481 ();
 sg13g2_decap_4 FILLER_39_486 ();
 sg13g2_fill_1 FILLER_39_490 ();
 sg13g2_fill_2 FILLER_39_504 ();
 sg13g2_decap_8 FILLER_39_510 ();
 sg13g2_fill_2 FILLER_39_517 ();
 sg13g2_fill_1 FILLER_39_524 ();
 sg13g2_decap_8 FILLER_39_535 ();
 sg13g2_decap_8 FILLER_39_542 ();
 sg13g2_fill_1 FILLER_39_549 ();
 sg13g2_fill_2 FILLER_39_576 ();
 sg13g2_fill_1 FILLER_39_587 ();
 sg13g2_fill_1 FILLER_39_609 ();
 sg13g2_fill_1 FILLER_39_617 ();
 sg13g2_decap_8 FILLER_39_624 ();
 sg13g2_decap_4 FILLER_39_631 ();
 sg13g2_decap_4 FILLER_39_651 ();
 sg13g2_fill_1 FILLER_39_655 ();
 sg13g2_fill_2 FILLER_39_681 ();
 sg13g2_fill_1 FILLER_39_740 ();
 sg13g2_decap_4 FILLER_39_749 ();
 sg13g2_decap_4 FILLER_39_770 ();
 sg13g2_fill_2 FILLER_39_794 ();
 sg13g2_fill_1 FILLER_39_796 ();
 sg13g2_fill_2 FILLER_39_801 ();
 sg13g2_fill_1 FILLER_39_803 ();
 sg13g2_decap_4 FILLER_39_819 ();
 sg13g2_fill_1 FILLER_39_823 ();
 sg13g2_decap_8 FILLER_39_833 ();
 sg13g2_decap_8 FILLER_39_840 ();
 sg13g2_decap_8 FILLER_39_847 ();
 sg13g2_decap_8 FILLER_39_854 ();
 sg13g2_decap_8 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_39_868 ();
 sg13g2_fill_2 FILLER_39_875 ();
 sg13g2_fill_1 FILLER_39_877 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_4 FILLER_40_105 ();
 sg13g2_fill_2 FILLER_40_121 ();
 sg13g2_fill_1 FILLER_40_123 ();
 sg13g2_fill_2 FILLER_40_133 ();
 sg13g2_fill_2 FILLER_40_140 ();
 sg13g2_fill_1 FILLER_40_151 ();
 sg13g2_decap_4 FILLER_40_157 ();
 sg13g2_fill_2 FILLER_40_165 ();
 sg13g2_fill_2 FILLER_40_219 ();
 sg13g2_fill_2 FILLER_40_229 ();
 sg13g2_fill_1 FILLER_40_231 ();
 sg13g2_fill_2 FILLER_40_237 ();
 sg13g2_fill_2 FILLER_40_244 ();
 sg13g2_fill_2 FILLER_40_250 ();
 sg13g2_fill_2 FILLER_40_262 ();
 sg13g2_fill_1 FILLER_40_264 ();
 sg13g2_fill_1 FILLER_40_283 ();
 sg13g2_decap_8 FILLER_40_289 ();
 sg13g2_decap_8 FILLER_40_296 ();
 sg13g2_fill_2 FILLER_40_303 ();
 sg13g2_fill_2 FILLER_40_338 ();
 sg13g2_fill_2 FILLER_40_355 ();
 sg13g2_decap_8 FILLER_40_366 ();
 sg13g2_fill_2 FILLER_40_373 ();
 sg13g2_fill_1 FILLER_40_399 ();
 sg13g2_fill_2 FILLER_40_413 ();
 sg13g2_fill_1 FILLER_40_428 ();
 sg13g2_fill_1 FILLER_40_446 ();
 sg13g2_fill_1 FILLER_40_492 ();
 sg13g2_fill_2 FILLER_40_524 ();
 sg13g2_decap_8 FILLER_40_536 ();
 sg13g2_fill_2 FILLER_40_568 ();
 sg13g2_fill_2 FILLER_40_601 ();
 sg13g2_fill_1 FILLER_40_603 ();
 sg13g2_fill_2 FILLER_40_612 ();
 sg13g2_decap_4 FILLER_40_627 ();
 sg13g2_fill_1 FILLER_40_631 ();
 sg13g2_fill_2 FILLER_40_652 ();
 sg13g2_fill_1 FILLER_40_654 ();
 sg13g2_decap_4 FILLER_40_668 ();
 sg13g2_fill_2 FILLER_40_686 ();
 sg13g2_decap_8 FILLER_40_692 ();
 sg13g2_decap_8 FILLER_40_699 ();
 sg13g2_decap_4 FILLER_40_706 ();
 sg13g2_fill_1 FILLER_40_710 ();
 sg13g2_decap_4 FILLER_40_731 ();
 sg13g2_fill_2 FILLER_40_755 ();
 sg13g2_fill_1 FILLER_40_757 ();
 sg13g2_fill_2 FILLER_40_767 ();
 sg13g2_fill_1 FILLER_40_787 ();
 sg13g2_fill_1 FILLER_40_803 ();
 sg13g2_fill_1 FILLER_40_809 ();
 sg13g2_fill_1 FILLER_40_819 ();
 sg13g2_decap_8 FILLER_40_849 ();
 sg13g2_decap_8 FILLER_40_856 ();
 sg13g2_decap_8 FILLER_40_863 ();
 sg13g2_decap_8 FILLER_40_870 ();
 sg13g2_fill_1 FILLER_40_877 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_fill_2 FILLER_41_91 ();
 sg13g2_fill_2 FILLER_41_119 ();
 sg13g2_fill_1 FILLER_41_126 ();
 sg13g2_fill_2 FILLER_41_134 ();
 sg13g2_fill_1 FILLER_41_136 ();
 sg13g2_fill_2 FILLER_41_153 ();
 sg13g2_fill_1 FILLER_41_160 ();
 sg13g2_decap_4 FILLER_41_166 ();
 sg13g2_fill_2 FILLER_41_176 ();
 sg13g2_fill_1 FILLER_41_178 ();
 sg13g2_decap_4 FILLER_41_185 ();
 sg13g2_decap_8 FILLER_41_200 ();
 sg13g2_decap_8 FILLER_41_207 ();
 sg13g2_fill_2 FILLER_41_214 ();
 sg13g2_fill_2 FILLER_41_235 ();
 sg13g2_fill_1 FILLER_41_240 ();
 sg13g2_fill_2 FILLER_41_250 ();
 sg13g2_fill_1 FILLER_41_257 ();
 sg13g2_fill_1 FILLER_41_262 ();
 sg13g2_fill_1 FILLER_41_268 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_fill_1 FILLER_41_280 ();
 sg13g2_fill_1 FILLER_41_287 ();
 sg13g2_fill_2 FILLER_41_319 ();
 sg13g2_decap_8 FILLER_41_365 ();
 sg13g2_decap_4 FILLER_41_372 ();
 sg13g2_fill_1 FILLER_41_376 ();
 sg13g2_fill_1 FILLER_41_381 ();
 sg13g2_fill_1 FILLER_41_405 ();
 sg13g2_fill_1 FILLER_41_413 ();
 sg13g2_fill_2 FILLER_41_452 ();
 sg13g2_fill_2 FILLER_41_480 ();
 sg13g2_fill_1 FILLER_41_482 ();
 sg13g2_fill_1 FILLER_41_491 ();
 sg13g2_fill_1 FILLER_41_507 ();
 sg13g2_decap_4 FILLER_41_516 ();
 sg13g2_fill_2 FILLER_41_520 ();
 sg13g2_fill_2 FILLER_41_531 ();
 sg13g2_fill_2 FILLER_41_545 ();
 sg13g2_fill_1 FILLER_41_570 ();
 sg13g2_decap_4 FILLER_41_576 ();
 sg13g2_fill_1 FILLER_41_580 ();
 sg13g2_decap_4 FILLER_41_585 ();
 sg13g2_fill_2 FILLER_41_589 ();
 sg13g2_fill_2 FILLER_41_601 ();
 sg13g2_fill_2 FILLER_41_655 ();
 sg13g2_fill_2 FILLER_41_673 ();
 sg13g2_fill_2 FILLER_41_680 ();
 sg13g2_fill_1 FILLER_41_691 ();
 sg13g2_decap_8 FILLER_41_696 ();
 sg13g2_decap_8 FILLER_41_703 ();
 sg13g2_fill_2 FILLER_41_726 ();
 sg13g2_fill_1 FILLER_41_728 ();
 sg13g2_decap_4 FILLER_41_747 ();
 sg13g2_fill_1 FILLER_41_780 ();
 sg13g2_fill_1 FILLER_41_807 ();
 sg13g2_decap_4 FILLER_41_814 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_854 ();
 sg13g2_decap_8 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_41_868 ();
 sg13g2_fill_2 FILLER_41_875 ();
 sg13g2_fill_1 FILLER_41_877 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_fill_2 FILLER_42_70 ();
 sg13g2_fill_1 FILLER_42_72 ();
 sg13g2_fill_1 FILLER_42_80 ();
 sg13g2_fill_1 FILLER_42_89 ();
 sg13g2_fill_2 FILLER_42_94 ();
 sg13g2_fill_2 FILLER_42_122 ();
 sg13g2_fill_2 FILLER_42_128 ();
 sg13g2_fill_1 FILLER_42_130 ();
 sg13g2_decap_8 FILLER_42_148 ();
 sg13g2_fill_1 FILLER_42_161 ();
 sg13g2_fill_2 FILLER_42_170 ();
 sg13g2_fill_1 FILLER_42_172 ();
 sg13g2_fill_2 FILLER_42_185 ();
 sg13g2_fill_1 FILLER_42_187 ();
 sg13g2_decap_4 FILLER_42_240 ();
 sg13g2_fill_2 FILLER_42_244 ();
 sg13g2_fill_2 FILLER_42_250 ();
 sg13g2_fill_2 FILLER_42_261 ();
 sg13g2_fill_1 FILLER_42_263 ();
 sg13g2_fill_1 FILLER_42_269 ();
 sg13g2_decap_8 FILLER_42_275 ();
 sg13g2_fill_2 FILLER_42_282 ();
 sg13g2_fill_1 FILLER_42_284 ();
 sg13g2_fill_2 FILLER_42_298 ();
 sg13g2_fill_1 FILLER_42_304 ();
 sg13g2_fill_1 FILLER_42_309 ();
 sg13g2_fill_1 FILLER_42_315 ();
 sg13g2_fill_1 FILLER_42_320 ();
 sg13g2_decap_4 FILLER_42_325 ();
 sg13g2_decap_8 FILLER_42_333 ();
 sg13g2_decap_8 FILLER_42_340 ();
 sg13g2_fill_1 FILLER_42_370 ();
 sg13g2_fill_2 FILLER_42_375 ();
 sg13g2_fill_1 FILLER_42_386 ();
 sg13g2_fill_2 FILLER_42_392 ();
 sg13g2_fill_2 FILLER_42_420 ();
 sg13g2_decap_8 FILLER_42_444 ();
 sg13g2_decap_8 FILLER_42_482 ();
 sg13g2_decap_8 FILLER_42_489 ();
 sg13g2_fill_1 FILLER_42_496 ();
 sg13g2_decap_8 FILLER_42_501 ();
 sg13g2_fill_2 FILLER_42_508 ();
 sg13g2_fill_1 FILLER_42_529 ();
 sg13g2_fill_1 FILLER_42_535 ();
 sg13g2_fill_1 FILLER_42_541 ();
 sg13g2_fill_1 FILLER_42_552 ();
 sg13g2_fill_2 FILLER_42_557 ();
 sg13g2_decap_8 FILLER_42_570 ();
 sg13g2_decap_4 FILLER_42_577 ();
 sg13g2_fill_2 FILLER_42_610 ();
 sg13g2_fill_2 FILLER_42_616 ();
 sg13g2_fill_1 FILLER_42_618 ();
 sg13g2_decap_8 FILLER_42_629 ();
 sg13g2_decap_8 FILLER_42_636 ();
 sg13g2_decap_4 FILLER_42_643 ();
 sg13g2_fill_2 FILLER_42_652 ();
 sg13g2_fill_1 FILLER_42_659 ();
 sg13g2_fill_2 FILLER_42_665 ();
 sg13g2_fill_2 FILLER_42_672 ();
 sg13g2_fill_2 FILLER_42_678 ();
 sg13g2_fill_1 FILLER_42_680 ();
 sg13g2_fill_2 FILLER_42_707 ();
 sg13g2_fill_2 FILLER_42_725 ();
 sg13g2_fill_2 FILLER_42_731 ();
 sg13g2_fill_2 FILLER_42_743 ();
 sg13g2_fill_1 FILLER_42_745 ();
 sg13g2_fill_2 FILLER_42_787 ();
 sg13g2_fill_1 FILLER_42_789 ();
 sg13g2_fill_1 FILLER_42_799 ();
 sg13g2_fill_2 FILLER_42_813 ();
 sg13g2_decap_8 FILLER_42_848 ();
 sg13g2_decap_8 FILLER_42_855 ();
 sg13g2_decap_8 FILLER_42_862 ();
 sg13g2_decap_8 FILLER_42_869 ();
 sg13g2_fill_2 FILLER_42_876 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_fill_2 FILLER_43_72 ();
 sg13g2_fill_1 FILLER_43_74 ();
 sg13g2_fill_2 FILLER_43_98 ();
 sg13g2_fill_1 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_118 ();
 sg13g2_fill_2 FILLER_43_125 ();
 sg13g2_fill_2 FILLER_43_132 ();
 sg13g2_fill_1 FILLER_43_144 ();
 sg13g2_fill_2 FILLER_43_153 ();
 sg13g2_fill_2 FILLER_43_159 ();
 sg13g2_fill_2 FILLER_43_168 ();
 sg13g2_fill_1 FILLER_43_170 ();
 sg13g2_decap_8 FILLER_43_194 ();
 sg13g2_fill_2 FILLER_43_201 ();
 sg13g2_fill_1 FILLER_43_203 ();
 sg13g2_fill_1 FILLER_43_209 ();
 sg13g2_fill_1 FILLER_43_214 ();
 sg13g2_fill_1 FILLER_43_220 ();
 sg13g2_fill_1 FILLER_43_228 ();
 sg13g2_fill_2 FILLER_43_281 ();
 sg13g2_fill_2 FILLER_43_313 ();
 sg13g2_decap_8 FILLER_43_359 ();
 sg13g2_decap_4 FILLER_43_366 ();
 sg13g2_fill_2 FILLER_43_370 ();
 sg13g2_decap_4 FILLER_43_376 ();
 sg13g2_fill_2 FILLER_43_410 ();
 sg13g2_decap_4 FILLER_43_432 ();
 sg13g2_fill_2 FILLER_43_436 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_4 FILLER_43_448 ();
 sg13g2_decap_4 FILLER_43_474 ();
 sg13g2_fill_1 FILLER_43_483 ();
 sg13g2_decap_8 FILLER_43_512 ();
 sg13g2_fill_1 FILLER_43_519 ();
 sg13g2_decap_8 FILLER_43_525 ();
 sg13g2_fill_1 FILLER_43_532 ();
 sg13g2_fill_1 FILLER_43_568 ();
 sg13g2_fill_1 FILLER_43_603 ();
 sg13g2_fill_2 FILLER_43_613 ();
 sg13g2_fill_1 FILLER_43_615 ();
 sg13g2_fill_1 FILLER_43_643 ();
 sg13g2_decap_8 FILLER_43_649 ();
 sg13g2_decap_8 FILLER_43_662 ();
 sg13g2_fill_2 FILLER_43_669 ();
 sg13g2_fill_1 FILLER_43_671 ();
 sg13g2_decap_4 FILLER_43_681 ();
 sg13g2_decap_4 FILLER_43_753 ();
 sg13g2_fill_2 FILLER_43_810 ();
 sg13g2_fill_1 FILLER_43_812 ();
 sg13g2_fill_1 FILLER_43_827 ();
 sg13g2_decap_8 FILLER_43_833 ();
 sg13g2_decap_8 FILLER_43_840 ();
 sg13g2_decap_8 FILLER_43_847 ();
 sg13g2_decap_8 FILLER_43_854 ();
 sg13g2_decap_8 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_43_868 ();
 sg13g2_fill_2 FILLER_43_875 ();
 sg13g2_fill_1 FILLER_43_877 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_fill_2 FILLER_44_73 ();
 sg13g2_fill_1 FILLER_44_133 ();
 sg13g2_fill_2 FILLER_44_139 ();
 sg13g2_fill_1 FILLER_44_141 ();
 sg13g2_fill_2 FILLER_44_154 ();
 sg13g2_fill_1 FILLER_44_156 ();
 sg13g2_fill_1 FILLER_44_162 ();
 sg13g2_fill_1 FILLER_44_171 ();
 sg13g2_fill_1 FILLER_44_180 ();
 sg13g2_fill_1 FILLER_44_187 ();
 sg13g2_fill_2 FILLER_44_205 ();
 sg13g2_fill_2 FILLER_44_221 ();
 sg13g2_fill_2 FILLER_44_228 ();
 sg13g2_fill_1 FILLER_44_296 ();
 sg13g2_fill_1 FILLER_44_320 ();
 sg13g2_fill_1 FILLER_44_330 ();
 sg13g2_fill_2 FILLER_44_336 ();
 sg13g2_fill_1 FILLER_44_338 ();
 sg13g2_fill_1 FILLER_44_394 ();
 sg13g2_fill_1 FILLER_44_405 ();
 sg13g2_fill_1 FILLER_44_411 ();
 sg13g2_fill_1 FILLER_44_418 ();
 sg13g2_fill_2 FILLER_44_445 ();
 sg13g2_decap_4 FILLER_44_451 ();
 sg13g2_fill_2 FILLER_44_455 ();
 sg13g2_fill_1 FILLER_44_482 ();
 sg13g2_fill_2 FILLER_44_488 ();
 sg13g2_fill_1 FILLER_44_490 ();
 sg13g2_decap_4 FILLER_44_510 ();
 sg13g2_fill_1 FILLER_44_518 ();
 sg13g2_decap_8 FILLER_44_558 ();
 sg13g2_fill_1 FILLER_44_573 ();
 sg13g2_fill_2 FILLER_44_583 ();
 sg13g2_fill_1 FILLER_44_585 ();
 sg13g2_fill_1 FILLER_44_609 ();
 sg13g2_fill_1 FILLER_44_639 ();
 sg13g2_fill_1 FILLER_44_654 ();
 sg13g2_fill_2 FILLER_44_668 ();
 sg13g2_fill_1 FILLER_44_691 ();
 sg13g2_fill_1 FILLER_44_697 ();
 sg13g2_fill_1 FILLER_44_711 ();
 sg13g2_decap_4 FILLER_44_723 ();
 sg13g2_fill_2 FILLER_44_735 ();
 sg13g2_decap_4 FILLER_44_748 ();
 sg13g2_fill_1 FILLER_44_755 ();
 sg13g2_fill_2 FILLER_44_770 ();
 sg13g2_fill_1 FILLER_44_777 ();
 sg13g2_fill_2 FILLER_44_792 ();
 sg13g2_fill_1 FILLER_44_794 ();
 sg13g2_fill_2 FILLER_44_800 ();
 sg13g2_fill_2 FILLER_44_806 ();
 sg13g2_fill_1 FILLER_44_808 ();
 sg13g2_decap_8 FILLER_44_838 ();
 sg13g2_decap_8 FILLER_44_845 ();
 sg13g2_decap_8 FILLER_44_852 ();
 sg13g2_decap_8 FILLER_44_859 ();
 sg13g2_decap_8 FILLER_44_866 ();
 sg13g2_decap_4 FILLER_44_873 ();
 sg13g2_fill_1 FILLER_44_877 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_fill_2 FILLER_45_63 ();
 sg13g2_fill_1 FILLER_45_65 ();
 sg13g2_fill_2 FILLER_45_94 ();
 sg13g2_fill_1 FILLER_45_96 ();
 sg13g2_decap_8 FILLER_45_120 ();
 sg13g2_fill_2 FILLER_45_163 ();
 sg13g2_fill_2 FILLER_45_172 ();
 sg13g2_fill_1 FILLER_45_174 ();
 sg13g2_decap_8 FILLER_45_180 ();
 sg13g2_decap_8 FILLER_45_190 ();
 sg13g2_decap_4 FILLER_45_212 ();
 sg13g2_fill_1 FILLER_45_216 ();
 sg13g2_fill_1 FILLER_45_234 ();
 sg13g2_fill_1 FILLER_45_247 ();
 sg13g2_fill_2 FILLER_45_293 ();
 sg13g2_fill_2 FILLER_45_300 ();
 sg13g2_fill_1 FILLER_45_302 ();
 sg13g2_decap_4 FILLER_45_307 ();
 sg13g2_fill_1 FILLER_45_311 ();
 sg13g2_decap_4 FILLER_45_330 ();
 sg13g2_fill_1 FILLER_45_370 ();
 sg13g2_decap_4 FILLER_45_376 ();
 sg13g2_fill_2 FILLER_45_380 ();
 sg13g2_decap_8 FILLER_45_386 ();
 sg13g2_fill_1 FILLER_45_393 ();
 sg13g2_fill_2 FILLER_45_399 ();
 sg13g2_decap_4 FILLER_45_415 ();
 sg13g2_fill_1 FILLER_45_419 ();
 sg13g2_decap_4 FILLER_45_430 ();
 sg13g2_fill_2 FILLER_45_460 ();
 sg13g2_fill_1 FILLER_45_462 ();
 sg13g2_fill_2 FILLER_45_473 ();
 sg13g2_fill_1 FILLER_45_475 ();
 sg13g2_fill_2 FILLER_45_486 ();
 sg13g2_fill_1 FILLER_45_496 ();
 sg13g2_fill_1 FILLER_45_506 ();
 sg13g2_fill_1 FILLER_45_511 ();
 sg13g2_fill_2 FILLER_45_516 ();
 sg13g2_fill_2 FILLER_45_523 ();
 sg13g2_fill_1 FILLER_45_525 ();
 sg13g2_fill_2 FILLER_45_530 ();
 sg13g2_fill_1 FILLER_45_532 ();
 sg13g2_fill_2 FILLER_45_540 ();
 sg13g2_decap_8 FILLER_45_546 ();
 sg13g2_fill_1 FILLER_45_609 ();
 sg13g2_fill_1 FILLER_45_620 ();
 sg13g2_fill_2 FILLER_45_626 ();
 sg13g2_fill_1 FILLER_45_634 ();
 sg13g2_fill_2 FILLER_45_640 ();
 sg13g2_fill_1 FILLER_45_651 ();
 sg13g2_fill_2 FILLER_45_684 ();
 sg13g2_decap_4 FILLER_45_701 ();
 sg13g2_fill_2 FILLER_45_744 ();
 sg13g2_decap_4 FILLER_45_761 ();
 sg13g2_fill_1 FILLER_45_765 ();
 sg13g2_fill_1 FILLER_45_783 ();
 sg13g2_fill_2 FILLER_45_792 ();
 sg13g2_fill_1 FILLER_45_808 ();
 sg13g2_decap_4 FILLER_45_814 ();
 sg13g2_fill_2 FILLER_45_823 ();
 sg13g2_decap_8 FILLER_45_851 ();
 sg13g2_decap_8 FILLER_45_858 ();
 sg13g2_decap_8 FILLER_45_865 ();
 sg13g2_decap_4 FILLER_45_872 ();
 sg13g2_fill_2 FILLER_45_876 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_4 FILLER_46_63 ();
 sg13g2_fill_1 FILLER_46_67 ();
 sg13g2_fill_1 FILLER_46_83 ();
 sg13g2_fill_2 FILLER_46_89 ();
 sg13g2_fill_1 FILLER_46_116 ();
 sg13g2_decap_8 FILLER_46_121 ();
 sg13g2_fill_1 FILLER_46_128 ();
 sg13g2_fill_1 FILLER_46_152 ();
 sg13g2_fill_1 FILLER_46_177 ();
 sg13g2_decap_4 FILLER_46_183 ();
 sg13g2_fill_1 FILLER_46_187 ();
 sg13g2_fill_1 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_209 ();
 sg13g2_fill_1 FILLER_46_216 ();
 sg13g2_fill_1 FILLER_46_246 ();
 sg13g2_fill_1 FILLER_46_253 ();
 sg13g2_fill_1 FILLER_46_266 ();
 sg13g2_fill_2 FILLER_46_291 ();
 sg13g2_fill_1 FILLER_46_298 ();
 sg13g2_fill_1 FILLER_46_309 ();
 sg13g2_fill_1 FILLER_46_315 ();
 sg13g2_fill_1 FILLER_46_321 ();
 sg13g2_fill_2 FILLER_46_354 ();
 sg13g2_fill_1 FILLER_46_370 ();
 sg13g2_fill_1 FILLER_46_381 ();
 sg13g2_decap_8 FILLER_46_397 ();
 sg13g2_fill_2 FILLER_46_404 ();
 sg13g2_fill_1 FILLER_46_406 ();
 sg13g2_decap_4 FILLER_46_412 ();
 sg13g2_decap_4 FILLER_46_442 ();
 sg13g2_fill_1 FILLER_46_446 ();
 sg13g2_decap_4 FILLER_46_456 ();
 sg13g2_fill_1 FILLER_46_460 ();
 sg13g2_fill_2 FILLER_46_469 ();
 sg13g2_fill_2 FILLER_46_476 ();
 sg13g2_fill_1 FILLER_46_478 ();
 sg13g2_fill_2 FILLER_46_489 ();
 sg13g2_fill_1 FILLER_46_501 ();
 sg13g2_fill_2 FILLER_46_543 ();
 sg13g2_fill_2 FILLER_46_576 ();
 sg13g2_decap_8 FILLER_46_583 ();
 sg13g2_decap_4 FILLER_46_594 ();
 sg13g2_fill_2 FILLER_46_602 ();
 sg13g2_fill_1 FILLER_46_604 ();
 sg13g2_fill_1 FILLER_46_621 ();
 sg13g2_decap_4 FILLER_46_626 ();
 sg13g2_fill_2 FILLER_46_640 ();
 sg13g2_fill_1 FILLER_46_642 ();
 sg13g2_fill_1 FILLER_46_661 ();
 sg13g2_fill_1 FILLER_46_672 ();
 sg13g2_decap_8 FILLER_46_681 ();
 sg13g2_decap_8 FILLER_46_688 ();
 sg13g2_decap_8 FILLER_46_695 ();
 sg13g2_fill_2 FILLER_46_702 ();
 sg13g2_fill_1 FILLER_46_729 ();
 sg13g2_fill_1 FILLER_46_743 ();
 sg13g2_fill_2 FILLER_46_757 ();
 sg13g2_fill_1 FILLER_46_759 ();
 sg13g2_decap_4 FILLER_46_764 ();
 sg13g2_fill_1 FILLER_46_768 ();
 sg13g2_decap_4 FILLER_46_774 ();
 sg13g2_fill_1 FILLER_46_778 ();
 sg13g2_fill_2 FILLER_46_787 ();
 sg13g2_fill_1 FILLER_46_789 ();
 sg13g2_fill_2 FILLER_46_795 ();
 sg13g2_fill_1 FILLER_46_797 ();
 sg13g2_decap_8 FILLER_46_830 ();
 sg13g2_decap_8 FILLER_46_837 ();
 sg13g2_decap_8 FILLER_46_844 ();
 sg13g2_decap_8 FILLER_46_851 ();
 sg13g2_decap_8 FILLER_46_858 ();
 sg13g2_decap_8 FILLER_46_865 ();
 sg13g2_decap_4 FILLER_46_872 ();
 sg13g2_fill_2 FILLER_46_876 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_68 ();
 sg13g2_fill_2 FILLER_47_75 ();
 sg13g2_decap_4 FILLER_47_89 ();
 sg13g2_fill_1 FILLER_47_98 ();
 sg13g2_fill_2 FILLER_47_104 ();
 sg13g2_decap_4 FILLER_47_129 ();
 sg13g2_fill_2 FILLER_47_170 ();
 sg13g2_fill_2 FILLER_47_188 ();
 sg13g2_fill_2 FILLER_47_195 ();
 sg13g2_decap_4 FILLER_47_207 ();
 sg13g2_decap_8 FILLER_47_233 ();
 sg13g2_fill_1 FILLER_47_240 ();
 sg13g2_fill_1 FILLER_47_255 ();
 sg13g2_fill_2 FILLER_47_293 ();
 sg13g2_fill_1 FILLER_47_295 ();
 sg13g2_fill_2 FILLER_47_300 ();
 sg13g2_fill_1 FILLER_47_302 ();
 sg13g2_fill_1 FILLER_47_308 ();
 sg13g2_fill_1 FILLER_47_314 ();
 sg13g2_fill_1 FILLER_47_326 ();
 sg13g2_decap_4 FILLER_47_331 ();
 sg13g2_fill_2 FILLER_47_335 ();
 sg13g2_decap_4 FILLER_47_343 ();
 sg13g2_fill_2 FILLER_47_347 ();
 sg13g2_fill_2 FILLER_47_364 ();
 sg13g2_decap_4 FILLER_47_375 ();
 sg13g2_fill_2 FILLER_47_395 ();
 sg13g2_decap_4 FILLER_47_401 ();
 sg13g2_fill_1 FILLER_47_410 ();
 sg13g2_decap_4 FILLER_47_448 ();
 sg13g2_fill_2 FILLER_47_477 ();
 sg13g2_fill_1 FILLER_47_479 ();
 sg13g2_decap_4 FILLER_47_487 ();
 sg13g2_fill_1 FILLER_47_491 ();
 sg13g2_fill_2 FILLER_47_539 ();
 sg13g2_decap_4 FILLER_47_550 ();
 sg13g2_decap_8 FILLER_47_577 ();
 sg13g2_decap_8 FILLER_47_584 ();
 sg13g2_fill_1 FILLER_47_591 ();
 sg13g2_fill_1 FILLER_47_596 ();
 sg13g2_decap_8 FILLER_47_609 ();
 sg13g2_fill_2 FILLER_47_631 ();
 sg13g2_fill_1 FILLER_47_633 ();
 sg13g2_fill_1 FILLER_47_639 ();
 sg13g2_fill_1 FILLER_47_645 ();
 sg13g2_fill_1 FILLER_47_672 ();
 sg13g2_fill_2 FILLER_47_695 ();
 sg13g2_fill_2 FILLER_47_701 ();
 sg13g2_fill_2 FILLER_47_720 ();
 sg13g2_fill_1 FILLER_47_722 ();
 sg13g2_fill_2 FILLER_47_729 ();
 sg13g2_fill_1 FILLER_47_754 ();
 sg13g2_fill_1 FILLER_47_760 ();
 sg13g2_fill_1 FILLER_47_765 ();
 sg13g2_fill_1 FILLER_47_772 ();
 sg13g2_fill_1 FILLER_47_778 ();
 sg13g2_fill_1 FILLER_47_792 ();
 sg13g2_fill_1 FILLER_47_797 ();
 sg13g2_decap_4 FILLER_47_806 ();
 sg13g2_fill_2 FILLER_47_810 ();
 sg13g2_fill_1 FILLER_47_823 ();
 sg13g2_decap_8 FILLER_47_832 ();
 sg13g2_decap_8 FILLER_47_839 ();
 sg13g2_decap_8 FILLER_47_846 ();
 sg13g2_decap_8 FILLER_47_853 ();
 sg13g2_decap_8 FILLER_47_860 ();
 sg13g2_decap_8 FILLER_47_867 ();
 sg13g2_decap_4 FILLER_47_874 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_fill_2 FILLER_48_49 ();
 sg13g2_fill_1 FILLER_48_51 ();
 sg13g2_fill_2 FILLER_48_83 ();
 sg13g2_fill_2 FILLER_48_91 ();
 sg13g2_fill_1 FILLER_48_119 ();
 sg13g2_fill_2 FILLER_48_146 ();
 sg13g2_fill_1 FILLER_48_148 ();
 sg13g2_fill_2 FILLER_48_156 ();
 sg13g2_fill_1 FILLER_48_158 ();
 sg13g2_fill_1 FILLER_48_167 ();
 sg13g2_decap_4 FILLER_48_200 ();
 sg13g2_fill_2 FILLER_48_204 ();
 sg13g2_decap_4 FILLER_48_211 ();
 sg13g2_fill_2 FILLER_48_239 ();
 sg13g2_fill_1 FILLER_48_241 ();
 sg13g2_fill_2 FILLER_48_255 ();
 sg13g2_fill_1 FILLER_48_257 ();
 sg13g2_fill_1 FILLER_48_263 ();
 sg13g2_fill_1 FILLER_48_283 ();
 sg13g2_fill_2 FILLER_48_295 ();
 sg13g2_fill_2 FILLER_48_332 ();
 sg13g2_fill_1 FILLER_48_339 ();
 sg13g2_fill_1 FILLER_48_347 ();
 sg13g2_fill_1 FILLER_48_363 ();
 sg13g2_fill_1 FILLER_48_400 ();
 sg13g2_fill_1 FILLER_48_411 ();
 sg13g2_decap_4 FILLER_48_421 ();
 sg13g2_decap_8 FILLER_48_439 ();
 sg13g2_fill_2 FILLER_48_446 ();
 sg13g2_decap_4 FILLER_48_453 ();
 sg13g2_fill_1 FILLER_48_457 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_503 ();
 sg13g2_decap_8 FILLER_48_597 ();
 sg13g2_decap_4 FILLER_48_608 ();
 sg13g2_fill_2 FILLER_48_612 ();
 sg13g2_fill_2 FILLER_48_638 ();
 sg13g2_decap_4 FILLER_48_658 ();
 sg13g2_fill_1 FILLER_48_662 ();
 sg13g2_decap_4 FILLER_48_683 ();
 sg13g2_fill_1 FILLER_48_692 ();
 sg13g2_fill_2 FILLER_48_702 ();
 sg13g2_fill_1 FILLER_48_728 ();
 sg13g2_fill_1 FILLER_48_733 ();
 sg13g2_fill_2 FILLER_48_739 ();
 sg13g2_fill_2 FILLER_48_758 ();
 sg13g2_fill_1 FILLER_48_760 ();
 sg13g2_fill_1 FILLER_48_773 ();
 sg13g2_fill_1 FILLER_48_780 ();
 sg13g2_fill_1 FILLER_48_786 ();
 sg13g2_decap_8 FILLER_48_849 ();
 sg13g2_decap_8 FILLER_48_856 ();
 sg13g2_decap_8 FILLER_48_863 ();
 sg13g2_decap_8 FILLER_48_870 ();
 sg13g2_fill_1 FILLER_48_877 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_4 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_48 ();
 sg13g2_decap_4 FILLER_49_55 ();
 sg13g2_fill_1 FILLER_49_59 ();
 sg13g2_decap_4 FILLER_49_64 ();
 sg13g2_fill_1 FILLER_49_68 ();
 sg13g2_decap_4 FILLER_49_73 ();
 sg13g2_fill_2 FILLER_49_82 ();
 sg13g2_fill_1 FILLER_49_84 ();
 sg13g2_fill_2 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_99 ();
 sg13g2_decap_4 FILLER_49_104 ();
 sg13g2_fill_2 FILLER_49_108 ();
 sg13g2_fill_1 FILLER_49_116 ();
 sg13g2_decap_8 FILLER_49_127 ();
 sg13g2_fill_1 FILLER_49_134 ();
 sg13g2_decap_4 FILLER_49_165 ();
 sg13g2_fill_2 FILLER_49_169 ();
 sg13g2_fill_2 FILLER_49_176 ();
 sg13g2_fill_1 FILLER_49_178 ();
 sg13g2_fill_1 FILLER_49_187 ();
 sg13g2_fill_1 FILLER_49_204 ();
 sg13g2_fill_2 FILLER_49_209 ();
 sg13g2_fill_1 FILLER_49_221 ();
 sg13g2_fill_1 FILLER_49_255 ();
 sg13g2_fill_2 FILLER_49_282 ();
 sg13g2_fill_2 FILLER_49_288 ();
 sg13g2_fill_1 FILLER_49_290 ();
 sg13g2_fill_2 FILLER_49_328 ();
 sg13g2_fill_2 FILLER_49_335 ();
 sg13g2_fill_1 FILLER_49_342 ();
 sg13g2_fill_2 FILLER_49_364 ();
 sg13g2_fill_1 FILLER_49_366 ();
 sg13g2_decap_4 FILLER_49_462 ();
 sg13g2_fill_2 FILLER_49_512 ();
 sg13g2_fill_1 FILLER_49_514 ();
 sg13g2_fill_2 FILLER_49_538 ();
 sg13g2_fill_1 FILLER_49_540 ();
 sg13g2_fill_2 FILLER_49_546 ();
 sg13g2_fill_1 FILLER_49_548 ();
 sg13g2_fill_2 FILLER_49_561 ();
 sg13g2_fill_1 FILLER_49_563 ();
 sg13g2_fill_1 FILLER_49_568 ();
 sg13g2_fill_2 FILLER_49_599 ();
 sg13g2_fill_1 FILLER_49_601 ();
 sg13g2_decap_8 FILLER_49_607 ();
 sg13g2_fill_1 FILLER_49_614 ();
 sg13g2_decap_8 FILLER_49_620 ();
 sg13g2_decap_8 FILLER_49_627 ();
 sg13g2_decap_8 FILLER_49_634 ();
 sg13g2_decap_4 FILLER_49_641 ();
 sg13g2_fill_1 FILLER_49_662 ();
 sg13g2_decap_4 FILLER_49_667 ();
 sg13g2_fill_1 FILLER_49_680 ();
 sg13g2_fill_2 FILLER_49_693 ();
 sg13g2_fill_1 FILLER_49_695 ();
 sg13g2_fill_1 FILLER_49_700 ();
 sg13g2_decap_8 FILLER_49_732 ();
 sg13g2_decap_8 FILLER_49_739 ();
 sg13g2_fill_2 FILLER_49_746 ();
 sg13g2_fill_1 FILLER_49_748 ();
 sg13g2_fill_2 FILLER_49_753 ();
 sg13g2_fill_2 FILLER_49_764 ();
 sg13g2_fill_1 FILLER_49_766 ();
 sg13g2_fill_1 FILLER_49_772 ();
 sg13g2_fill_2 FILLER_49_777 ();
 sg13g2_fill_1 FILLER_49_779 ();
 sg13g2_fill_1 FILLER_49_792 ();
 sg13g2_fill_1 FILLER_49_809 ();
 sg13g2_fill_1 FILLER_49_813 ();
 sg13g2_decap_8 FILLER_49_840 ();
 sg13g2_decap_8 FILLER_49_847 ();
 sg13g2_decap_8 FILLER_49_854 ();
 sg13g2_decap_8 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_49_868 ();
 sg13g2_fill_2 FILLER_49_875 ();
 sg13g2_fill_1 FILLER_49_877 ();
 sg13g2_decap_4 FILLER_50_26 ();
 sg13g2_fill_1 FILLER_50_30 ();
 sg13g2_fill_2 FILLER_50_35 ();
 sg13g2_fill_2 FILLER_50_63 ();
 sg13g2_fill_1 FILLER_50_65 ();
 sg13g2_fill_2 FILLER_50_92 ();
 sg13g2_decap_8 FILLER_50_97 ();
 sg13g2_decap_8 FILLER_50_104 ();
 sg13g2_decap_4 FILLER_50_111 ();
 sg13g2_fill_1 FILLER_50_118 ();
 sg13g2_fill_1 FILLER_50_153 ();
 sg13g2_fill_1 FILLER_50_171 ();
 sg13g2_fill_1 FILLER_50_182 ();
 sg13g2_fill_2 FILLER_50_188 ();
 sg13g2_fill_1 FILLER_50_190 ();
 sg13g2_fill_2 FILLER_50_196 ();
 sg13g2_fill_2 FILLER_50_202 ();
 sg13g2_fill_1 FILLER_50_213 ();
 sg13g2_fill_2 FILLER_50_222 ();
 sg13g2_fill_2 FILLER_50_228 ();
 sg13g2_fill_2 FILLER_50_235 ();
 sg13g2_fill_1 FILLER_50_237 ();
 sg13g2_decap_8 FILLER_50_246 ();
 sg13g2_decap_4 FILLER_50_253 ();
 sg13g2_fill_2 FILLER_50_257 ();
 sg13g2_decap_4 FILLER_50_271 ();
 sg13g2_fill_2 FILLER_50_275 ();
 sg13g2_fill_2 FILLER_50_285 ();
 sg13g2_fill_1 FILLER_50_292 ();
 sg13g2_fill_1 FILLER_50_299 ();
 sg13g2_fill_2 FILLER_50_306 ();
 sg13g2_fill_2 FILLER_50_314 ();
 sg13g2_fill_1 FILLER_50_343 ();
 sg13g2_fill_1 FILLER_50_381 ();
 sg13g2_fill_2 FILLER_50_391 ();
 sg13g2_fill_1 FILLER_50_423 ();
 sg13g2_fill_2 FILLER_50_474 ();
 sg13g2_fill_2 FILLER_50_484 ();
 sg13g2_decap_8 FILLER_50_495 ();
 sg13g2_decap_4 FILLER_50_502 ();
 sg13g2_fill_2 FILLER_50_506 ();
 sg13g2_fill_1 FILLER_50_550 ();
 sg13g2_decap_4 FILLER_50_566 ();
 sg13g2_fill_1 FILLER_50_570 ();
 sg13g2_decap_8 FILLER_50_580 ();
 sg13g2_fill_2 FILLER_50_587 ();
 sg13g2_fill_2 FILLER_50_593 ();
 sg13g2_decap_4 FILLER_50_607 ();
 sg13g2_fill_2 FILLER_50_633 ();
 sg13g2_decap_4 FILLER_50_639 ();
 sg13g2_fill_2 FILLER_50_643 ();
 sg13g2_fill_1 FILLER_50_689 ();
 sg13g2_decap_4 FILLER_50_694 ();
 sg13g2_fill_1 FILLER_50_698 ();
 sg13g2_fill_1 FILLER_50_703 ();
 sg13g2_fill_1 FILLER_50_719 ();
 sg13g2_decap_8 FILLER_50_741 ();
 sg13g2_fill_1 FILLER_50_748 ();
 sg13g2_fill_2 FILLER_50_754 ();
 sg13g2_decap_8 FILLER_50_760 ();
 sg13g2_fill_2 FILLER_50_767 ();
 sg13g2_fill_2 FILLER_50_814 ();
 sg13g2_decap_8 FILLER_50_820 ();
 sg13g2_decap_8 FILLER_50_837 ();
 sg13g2_decap_8 FILLER_50_844 ();
 sg13g2_decap_8 FILLER_50_851 ();
 sg13g2_decap_8 FILLER_50_858 ();
 sg13g2_decap_8 FILLER_50_865 ();
 sg13g2_decap_4 FILLER_50_872 ();
 sg13g2_fill_2 FILLER_50_876 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_fill_2 FILLER_51_23 ();
 sg13g2_fill_1 FILLER_51_25 ();
 sg13g2_fill_1 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_59 ();
 sg13g2_decap_4 FILLER_51_66 ();
 sg13g2_fill_2 FILLER_51_82 ();
 sg13g2_fill_1 FILLER_51_89 ();
 sg13g2_fill_1 FILLER_51_94 ();
 sg13g2_fill_1 FILLER_51_99 ();
 sg13g2_fill_2 FILLER_51_108 ();
 sg13g2_fill_1 FILLER_51_126 ();
 sg13g2_fill_2 FILLER_51_162 ();
 sg13g2_fill_1 FILLER_51_164 ();
 sg13g2_fill_1 FILLER_51_195 ();
 sg13g2_decap_4 FILLER_51_205 ();
 sg13g2_fill_1 FILLER_51_209 ();
 sg13g2_fill_1 FILLER_51_225 ();
 sg13g2_decap_4 FILLER_51_234 ();
 sg13g2_fill_1 FILLER_51_238 ();
 sg13g2_decap_4 FILLER_51_265 ();
 sg13g2_fill_1 FILLER_51_273 ();
 sg13g2_fill_1 FILLER_51_282 ();
 sg13g2_fill_1 FILLER_51_287 ();
 sg13g2_fill_1 FILLER_51_293 ();
 sg13g2_fill_1 FILLER_51_306 ();
 sg13g2_fill_1 FILLER_51_315 ();
 sg13g2_fill_1 FILLER_51_321 ();
 sg13g2_fill_2 FILLER_51_330 ();
 sg13g2_decap_4 FILLER_51_340 ();
 sg13g2_fill_2 FILLER_51_348 ();
 sg13g2_fill_2 FILLER_51_358 ();
 sg13g2_decap_4 FILLER_51_364 ();
 sg13g2_fill_1 FILLER_51_422 ();
 sg13g2_fill_2 FILLER_51_436 ();
 sg13g2_fill_2 FILLER_51_458 ();
 sg13g2_fill_2 FILLER_51_469 ();
 sg13g2_fill_1 FILLER_51_471 ();
 sg13g2_decap_8 FILLER_51_497 ();
 sg13g2_fill_2 FILLER_51_504 ();
 sg13g2_decap_8 FILLER_51_510 ();
 sg13g2_fill_1 FILLER_51_517 ();
 sg13g2_fill_1 FILLER_51_530 ();
 sg13g2_fill_1 FILLER_51_559 ();
 sg13g2_fill_2 FILLER_51_572 ();
 sg13g2_fill_2 FILLER_51_587 ();
 sg13g2_fill_2 FILLER_51_599 ();
 sg13g2_fill_1 FILLER_51_601 ();
 sg13g2_fill_2 FILLER_51_611 ();
 sg13g2_fill_1 FILLER_51_613 ();
 sg13g2_decap_4 FILLER_51_632 ();
 sg13g2_fill_2 FILLER_51_636 ();
 sg13g2_fill_2 FILLER_51_643 ();
 sg13g2_fill_1 FILLER_51_645 ();
 sg13g2_fill_1 FILLER_51_655 ();
 sg13g2_fill_2 FILLER_51_688 ();
 sg13g2_fill_1 FILLER_51_700 ();
 sg13g2_decap_4 FILLER_51_711 ();
 sg13g2_fill_1 FILLER_51_715 ();
 sg13g2_fill_2 FILLER_51_741 ();
 sg13g2_fill_2 FILLER_51_764 ();
 sg13g2_fill_2 FILLER_51_776 ();
 sg13g2_fill_1 FILLER_51_783 ();
 sg13g2_decap_4 FILLER_51_788 ();
 sg13g2_fill_1 FILLER_51_796 ();
 sg13g2_fill_2 FILLER_51_802 ();
 sg13g2_fill_1 FILLER_51_809 ();
 sg13g2_fill_1 FILLER_51_814 ();
 sg13g2_fill_2 FILLER_51_819 ();
 sg13g2_fill_1 FILLER_51_821 ();
 sg13g2_fill_2 FILLER_51_826 ();
 sg13g2_decap_8 FILLER_51_832 ();
 sg13g2_decap_8 FILLER_51_839 ();
 sg13g2_decap_8 FILLER_51_846 ();
 sg13g2_decap_8 FILLER_51_853 ();
 sg13g2_decap_8 FILLER_51_860 ();
 sg13g2_decap_8 FILLER_51_867 ();
 sg13g2_decap_4 FILLER_51_874 ();
 sg13g2_fill_2 FILLER_52_26 ();
 sg13g2_fill_1 FILLER_52_28 ();
 sg13g2_fill_1 FILLER_52_44 ();
 sg13g2_fill_2 FILLER_52_50 ();
 sg13g2_fill_1 FILLER_52_52 ();
 sg13g2_fill_2 FILLER_52_68 ();
 sg13g2_fill_1 FILLER_52_82 ();
 sg13g2_fill_1 FILLER_52_87 ();
 sg13g2_fill_1 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_117 ();
 sg13g2_fill_2 FILLER_52_124 ();
 sg13g2_fill_2 FILLER_52_136 ();
 sg13g2_fill_2 FILLER_52_142 ();
 sg13g2_fill_1 FILLER_52_144 ();
 sg13g2_fill_1 FILLER_52_149 ();
 sg13g2_fill_2 FILLER_52_154 ();
 sg13g2_fill_1 FILLER_52_156 ();
 sg13g2_decap_4 FILLER_52_174 ();
 sg13g2_fill_2 FILLER_52_178 ();
 sg13g2_decap_4 FILLER_52_200 ();
 sg13g2_fill_1 FILLER_52_204 ();
 sg13g2_fill_2 FILLER_52_221 ();
 sg13g2_fill_1 FILLER_52_231 ();
 sg13g2_fill_1 FILLER_52_237 ();
 sg13g2_fill_1 FILLER_52_248 ();
 sg13g2_fill_2 FILLER_52_257 ();
 sg13g2_fill_2 FILLER_52_264 ();
 sg13g2_fill_1 FILLER_52_295 ();
 sg13g2_fill_1 FILLER_52_319 ();
 sg13g2_fill_2 FILLER_52_334 ();
 sg13g2_decap_4 FILLER_52_340 ();
 sg13g2_fill_1 FILLER_52_348 ();
 sg13g2_decap_8 FILLER_52_375 ();
 sg13g2_fill_1 FILLER_52_386 ();
 sg13g2_fill_2 FILLER_52_396 ();
 sg13g2_fill_1 FILLER_52_407 ();
 sg13g2_fill_2 FILLER_52_451 ();
 sg13g2_fill_2 FILLER_52_463 ();
 sg13g2_fill_1 FILLER_52_465 ();
 sg13g2_decap_4 FILLER_52_500 ();
 sg13g2_decap_4 FILLER_52_513 ();
 sg13g2_fill_1 FILLER_52_524 ();
 sg13g2_fill_1 FILLER_52_532 ();
 sg13g2_fill_1 FILLER_52_541 ();
 sg13g2_fill_2 FILLER_52_554 ();
 sg13g2_decap_8 FILLER_52_566 ();
 sg13g2_fill_2 FILLER_52_593 ();
 sg13g2_fill_1 FILLER_52_600 ();
 sg13g2_fill_1 FILLER_52_608 ();
 sg13g2_fill_1 FILLER_52_620 ();
 sg13g2_fill_1 FILLER_52_625 ();
 sg13g2_fill_2 FILLER_52_635 ();
 sg13g2_fill_1 FILLER_52_646 ();
 sg13g2_fill_2 FILLER_52_680 ();
 sg13g2_fill_1 FILLER_52_682 ();
 sg13g2_decap_4 FILLER_52_695 ();
 sg13g2_fill_1 FILLER_52_714 ();
 sg13g2_fill_1 FILLER_52_719 ();
 sg13g2_fill_1 FILLER_52_728 ();
 sg13g2_fill_2 FILLER_52_734 ();
 sg13g2_decap_4 FILLER_52_741 ();
 sg13g2_fill_1 FILLER_52_779 ();
 sg13g2_fill_2 FILLER_52_785 ();
 sg13g2_fill_1 FILLER_52_791 ();
 sg13g2_fill_1 FILLER_52_796 ();
 sg13g2_fill_2 FILLER_52_801 ();
 sg13g2_fill_1 FILLER_52_815 ();
 sg13g2_fill_1 FILLER_52_821 ();
 sg13g2_decap_8 FILLER_52_826 ();
 sg13g2_decap_8 FILLER_52_833 ();
 sg13g2_decap_8 FILLER_52_840 ();
 sg13g2_decap_8 FILLER_52_847 ();
 sg13g2_decap_8 FILLER_52_854 ();
 sg13g2_decap_8 FILLER_52_861 ();
 sg13g2_decap_8 FILLER_52_868 ();
 sg13g2_fill_2 FILLER_52_875 ();
 sg13g2_fill_1 FILLER_52_877 ();
 sg13g2_decap_4 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_4 ();
 sg13g2_fill_2 FILLER_53_22 ();
 sg13g2_fill_2 FILLER_53_27 ();
 sg13g2_fill_2 FILLER_53_34 ();
 sg13g2_decap_4 FILLER_53_58 ();
 sg13g2_fill_1 FILLER_53_62 ();
 sg13g2_decap_4 FILLER_53_66 ();
 sg13g2_fill_2 FILLER_53_70 ();
 sg13g2_fill_2 FILLER_53_103 ();
 sg13g2_fill_2 FILLER_53_115 ();
 sg13g2_fill_2 FILLER_53_122 ();
 sg13g2_fill_1 FILLER_53_124 ();
 sg13g2_decap_4 FILLER_53_133 ();
 sg13g2_fill_2 FILLER_53_159 ();
 sg13g2_decap_4 FILLER_53_173 ();
 sg13g2_fill_2 FILLER_53_180 ();
 sg13g2_fill_1 FILLER_53_182 ();
 sg13g2_fill_2 FILLER_53_188 ();
 sg13g2_fill_2 FILLER_53_203 ();
 sg13g2_fill_1 FILLER_53_205 ();
 sg13g2_fill_2 FILLER_53_225 ();
 sg13g2_fill_2 FILLER_53_232 ();
 sg13g2_fill_1 FILLER_53_239 ();
 sg13g2_fill_1 FILLER_53_245 ();
 sg13g2_fill_1 FILLER_53_251 ();
 sg13g2_fill_2 FILLER_53_260 ();
 sg13g2_fill_1 FILLER_53_292 ();
 sg13g2_fill_1 FILLER_53_326 ();
 sg13g2_decap_4 FILLER_53_340 ();
 sg13g2_decap_8 FILLER_53_349 ();
 sg13g2_fill_1 FILLER_53_356 ();
 sg13g2_fill_2 FILLER_53_361 ();
 sg13g2_fill_2 FILLER_53_366 ();
 sg13g2_decap_4 FILLER_53_373 ();
 sg13g2_fill_1 FILLER_53_377 ();
 sg13g2_decap_4 FILLER_53_418 ();
 sg13g2_fill_1 FILLER_53_422 ();
 sg13g2_fill_2 FILLER_53_427 ();
 sg13g2_fill_1 FILLER_53_437 ();
 sg13g2_fill_2 FILLER_53_448 ();
 sg13g2_fill_1 FILLER_53_450 ();
 sg13g2_fill_2 FILLER_53_456 ();
 sg13g2_fill_1 FILLER_53_458 ();
 sg13g2_decap_8 FILLER_53_475 ();
 sg13g2_decap_4 FILLER_53_482 ();
 sg13g2_fill_2 FILLER_53_525 ();
 sg13g2_fill_1 FILLER_53_536 ();
 sg13g2_fill_2 FILLER_53_541 ();
 sg13g2_fill_2 FILLER_53_552 ();
 sg13g2_fill_1 FILLER_53_554 ();
 sg13g2_decap_8 FILLER_53_561 ();
 sg13g2_fill_1 FILLER_53_568 ();
 sg13g2_fill_2 FILLER_53_578 ();
 sg13g2_fill_1 FILLER_53_580 ();
 sg13g2_fill_2 FILLER_53_586 ();
 sg13g2_fill_2 FILLER_53_625 ();
 sg13g2_fill_1 FILLER_53_637 ();
 sg13g2_fill_1 FILLER_53_685 ();
 sg13g2_fill_1 FILLER_53_696 ();
 sg13g2_decap_4 FILLER_53_707 ();
 sg13g2_fill_1 FILLER_53_711 ();
 sg13g2_fill_2 FILLER_53_721 ();
 sg13g2_decap_8 FILLER_53_738 ();
 sg13g2_fill_1 FILLER_53_745 ();
 sg13g2_decap_4 FILLER_53_766 ();
 sg13g2_fill_1 FILLER_53_770 ();
 sg13g2_fill_2 FILLER_53_776 ();
 sg13g2_fill_2 FILLER_53_783 ();
 sg13g2_fill_1 FILLER_53_785 ();
 sg13g2_fill_2 FILLER_53_790 ();
 sg13g2_fill_1 FILLER_53_792 ();
 sg13g2_fill_2 FILLER_53_798 ();
 sg13g2_fill_1 FILLER_53_805 ();
 sg13g2_decap_8 FILLER_53_836 ();
 sg13g2_decap_8 FILLER_53_843 ();
 sg13g2_decap_8 FILLER_53_850 ();
 sg13g2_decap_8 FILLER_53_857 ();
 sg13g2_decap_8 FILLER_53_864 ();
 sg13g2_decap_8 FILLER_53_871 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_7 ();
 sg13g2_fill_1 FILLER_54_16 ();
 sg13g2_fill_1 FILLER_54_27 ();
 sg13g2_fill_1 FILLER_54_89 ();
 sg13g2_fill_1 FILLER_54_110 ();
 sg13g2_fill_1 FILLER_54_121 ();
 sg13g2_fill_1 FILLER_54_138 ();
 sg13g2_fill_1 FILLER_54_147 ();
 sg13g2_fill_1 FILLER_54_161 ();
 sg13g2_fill_2 FILLER_54_167 ();
 sg13g2_fill_1 FILLER_54_169 ();
 sg13g2_decap_8 FILLER_54_179 ();
 sg13g2_fill_2 FILLER_54_202 ();
 sg13g2_fill_2 FILLER_54_214 ();
 sg13g2_fill_1 FILLER_54_216 ();
 sg13g2_fill_1 FILLER_54_221 ();
 sg13g2_fill_2 FILLER_54_231 ();
 sg13g2_fill_1 FILLER_54_237 ();
 sg13g2_fill_1 FILLER_54_243 ();
 sg13g2_fill_2 FILLER_54_249 ();
 sg13g2_fill_1 FILLER_54_256 ();
 sg13g2_fill_1 FILLER_54_286 ();
 sg13g2_fill_1 FILLER_54_293 ();
 sg13g2_fill_1 FILLER_54_299 ();
 sg13g2_fill_1 FILLER_54_305 ();
 sg13g2_fill_1 FILLER_54_311 ();
 sg13g2_fill_2 FILLER_54_316 ();
 sg13g2_fill_2 FILLER_54_329 ();
 sg13g2_decap_8 FILLER_54_339 ();
 sg13g2_fill_1 FILLER_54_346 ();
 sg13g2_decap_4 FILLER_54_351 ();
 sg13g2_decap_8 FILLER_54_381 ();
 sg13g2_decap_8 FILLER_54_392 ();
 sg13g2_decap_4 FILLER_54_408 ();
 sg13g2_fill_2 FILLER_54_412 ();
 sg13g2_fill_2 FILLER_54_440 ();
 sg13g2_fill_1 FILLER_54_447 ();
 sg13g2_decap_8 FILLER_54_462 ();
 sg13g2_decap_8 FILLER_54_469 ();
 sg13g2_fill_2 FILLER_54_476 ();
 sg13g2_fill_1 FILLER_54_478 ();
 sg13g2_fill_2 FILLER_54_491 ();
 sg13g2_fill_1 FILLER_54_493 ();
 sg13g2_fill_1 FILLER_54_498 ();
 sg13g2_fill_2 FILLER_54_503 ();
 sg13g2_fill_1 FILLER_54_505 ();
 sg13g2_decap_8 FILLER_54_510 ();
 sg13g2_fill_2 FILLER_54_517 ();
 sg13g2_fill_2 FILLER_54_541 ();
 sg13g2_fill_1 FILLER_54_563 ();
 sg13g2_fill_2 FILLER_54_572 ();
 sg13g2_fill_1 FILLER_54_578 ();
 sg13g2_decap_4 FILLER_54_588 ();
 sg13g2_fill_1 FILLER_54_602 ();
 sg13g2_fill_1 FILLER_54_621 ();
 sg13g2_fill_1 FILLER_54_674 ();
 sg13g2_decap_4 FILLER_54_699 ();
 sg13g2_fill_1 FILLER_54_703 ();
 sg13g2_fill_1 FILLER_54_709 ();
 sg13g2_decap_4 FILLER_54_721 ();
 sg13g2_fill_1 FILLER_54_735 ();
 sg13g2_fill_1 FILLER_54_740 ();
 sg13g2_fill_1 FILLER_54_748 ();
 sg13g2_fill_1 FILLER_54_754 ();
 sg13g2_decap_8 FILLER_54_759 ();
 sg13g2_fill_1 FILLER_54_780 ();
 sg13g2_fill_2 FILLER_54_808 ();
 sg13g2_fill_1 FILLER_54_838 ();
 sg13g2_decap_8 FILLER_54_848 ();
 sg13g2_decap_8 FILLER_54_855 ();
 sg13g2_decap_8 FILLER_54_862 ();
 sg13g2_decap_8 FILLER_54_869 ();
 sg13g2_fill_2 FILLER_54_876 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_14 ();
 sg13g2_fill_1 FILLER_55_16 ();
 sg13g2_fill_1 FILLER_55_43 ();
 sg13g2_fill_2 FILLER_55_49 ();
 sg13g2_decap_4 FILLER_55_66 ();
 sg13g2_fill_1 FILLER_55_70 ();
 sg13g2_fill_1 FILLER_55_82 ();
 sg13g2_fill_2 FILLER_55_97 ();
 sg13g2_fill_1 FILLER_55_104 ();
 sg13g2_decap_8 FILLER_55_108 ();
 sg13g2_fill_2 FILLER_55_120 ();
 sg13g2_fill_1 FILLER_55_122 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_4 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_157 ();
 sg13g2_fill_2 FILLER_55_164 ();
 sg13g2_fill_1 FILLER_55_166 ();
 sg13g2_fill_1 FILLER_55_182 ();
 sg13g2_fill_2 FILLER_55_211 ();
 sg13g2_fill_1 FILLER_55_217 ();
 sg13g2_decap_8 FILLER_55_222 ();
 sg13g2_fill_1 FILLER_55_229 ();
 sg13g2_fill_1 FILLER_55_235 ();
 sg13g2_decap_8 FILLER_55_255 ();
 sg13g2_decap_4 FILLER_55_262 ();
 sg13g2_fill_2 FILLER_55_269 ();
 sg13g2_fill_2 FILLER_55_276 ();
 sg13g2_fill_2 FILLER_55_283 ();
 sg13g2_fill_2 FILLER_55_290 ();
 sg13g2_fill_1 FILLER_55_296 ();
 sg13g2_fill_2 FILLER_55_304 ();
 sg13g2_fill_2 FILLER_55_311 ();
 sg13g2_decap_4 FILLER_55_321 ();
 sg13g2_decap_4 FILLER_55_330 ();
 sg13g2_decap_4 FILLER_55_381 ();
 sg13g2_fill_2 FILLER_55_393 ();
 sg13g2_fill_1 FILLER_55_395 ();
 sg13g2_decap_8 FILLER_55_431 ();
 sg13g2_fill_2 FILLER_55_438 ();
 sg13g2_fill_1 FILLER_55_440 ();
 sg13g2_decap_8 FILLER_55_465 ();
 sg13g2_fill_1 FILLER_55_480 ();
 sg13g2_fill_1 FILLER_55_512 ();
 sg13g2_fill_1 FILLER_55_518 ();
 sg13g2_fill_1 FILLER_55_524 ();
 sg13g2_fill_1 FILLER_55_539 ();
 sg13g2_fill_1 FILLER_55_568 ();
 sg13g2_fill_1 FILLER_55_597 ();
 sg13g2_fill_1 FILLER_55_609 ();
 sg13g2_fill_1 FILLER_55_615 ();
 sg13g2_fill_2 FILLER_55_621 ();
 sg13g2_fill_2 FILLER_55_627 ();
 sg13g2_fill_1 FILLER_55_664 ();
 sg13g2_decap_4 FILLER_55_671 ();
 sg13g2_fill_1 FILLER_55_680 ();
 sg13g2_decap_8 FILLER_55_698 ();
 sg13g2_fill_1 FILLER_55_735 ();
 sg13g2_fill_1 FILLER_55_746 ();
 sg13g2_fill_1 FILLER_55_761 ();
 sg13g2_fill_2 FILLER_55_773 ();
 sg13g2_fill_2 FILLER_55_821 ();
 sg13g2_fill_2 FILLER_55_831 ();
 sg13g2_fill_1 FILLER_55_833 ();
 sg13g2_decap_8 FILLER_55_856 ();
 sg13g2_decap_8 FILLER_55_863 ();
 sg13g2_decap_8 FILLER_55_870 ();
 sg13g2_fill_1 FILLER_55_877 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_4 ();
 sg13g2_fill_1 FILLER_56_22 ();
 sg13g2_fill_2 FILLER_56_28 ();
 sg13g2_fill_1 FILLER_56_36 ();
 sg13g2_fill_2 FILLER_56_42 ();
 sg13g2_fill_2 FILLER_56_54 ();
 sg13g2_fill_2 FILLER_56_111 ();
 sg13g2_fill_1 FILLER_56_113 ();
 sg13g2_decap_8 FILLER_56_123 ();
 sg13g2_fill_1 FILLER_56_130 ();
 sg13g2_fill_1 FILLER_56_154 ();
 sg13g2_fill_2 FILLER_56_160 ();
 sg13g2_fill_2 FILLER_56_170 ();
 sg13g2_fill_1 FILLER_56_191 ();
 sg13g2_fill_1 FILLER_56_196 ();
 sg13g2_fill_2 FILLER_56_202 ();
 sg13g2_decap_4 FILLER_56_246 ();
 sg13g2_fill_1 FILLER_56_250 ();
 sg13g2_decap_4 FILLER_56_261 ();
 sg13g2_fill_1 FILLER_56_265 ();
 sg13g2_fill_1 FILLER_56_269 ();
 sg13g2_fill_2 FILLER_56_274 ();
 sg13g2_decap_4 FILLER_56_280 ();
 sg13g2_fill_1 FILLER_56_289 ();
 sg13g2_fill_2 FILLER_56_309 ();
 sg13g2_fill_2 FILLER_56_341 ();
 sg13g2_fill_1 FILLER_56_343 ();
 sg13g2_decap_4 FILLER_56_349 ();
 sg13g2_fill_2 FILLER_56_353 ();
 sg13g2_fill_2 FILLER_56_363 ();
 sg13g2_decap_4 FILLER_56_377 ();
 sg13g2_decap_4 FILLER_56_405 ();
 sg13g2_fill_2 FILLER_56_444 ();
 sg13g2_decap_8 FILLER_56_462 ();
 sg13g2_fill_2 FILLER_56_480 ();
 sg13g2_decap_8 FILLER_56_493 ();
 sg13g2_decap_4 FILLER_56_500 ();
 sg13g2_fill_2 FILLER_56_504 ();
 sg13g2_decap_4 FILLER_56_524 ();
 sg13g2_decap_4 FILLER_56_532 ();
 sg13g2_fill_1 FILLER_56_561 ();
 sg13g2_fill_1 FILLER_56_583 ();
 sg13g2_fill_2 FILLER_56_621 ();
 sg13g2_fill_1 FILLER_56_643 ();
 sg13g2_fill_1 FILLER_56_649 ();
 sg13g2_fill_2 FILLER_56_672 ();
 sg13g2_fill_2 FILLER_56_695 ();
 sg13g2_fill_1 FILLER_56_701 ();
 sg13g2_fill_2 FILLER_56_712 ();
 sg13g2_fill_2 FILLER_56_720 ();
 sg13g2_fill_1 FILLER_56_722 ();
 sg13g2_fill_1 FILLER_56_728 ();
 sg13g2_fill_1 FILLER_56_739 ();
 sg13g2_fill_1 FILLER_56_746 ();
 sg13g2_fill_1 FILLER_56_759 ();
 sg13g2_fill_2 FILLER_56_765 ();
 sg13g2_fill_1 FILLER_56_767 ();
 sg13g2_fill_2 FILLER_56_802 ();
 sg13g2_fill_1 FILLER_56_809 ();
 sg13g2_fill_2 FILLER_56_819 ();
 sg13g2_fill_1 FILLER_56_821 ();
 sg13g2_decap_4 FILLER_56_835 ();
 sg13g2_fill_1 FILLER_56_852 ();
 sg13g2_decap_8 FILLER_56_858 ();
 sg13g2_decap_8 FILLER_56_865 ();
 sg13g2_decap_4 FILLER_56_872 ();
 sg13g2_fill_2 FILLER_56_876 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_4 ();
 sg13g2_fill_1 FILLER_57_43 ();
 sg13g2_fill_2 FILLER_57_73 ();
 sg13g2_fill_1 FILLER_57_85 ();
 sg13g2_fill_1 FILLER_57_102 ();
 sg13g2_fill_2 FILLER_57_108 ();
 sg13g2_fill_1 FILLER_57_110 ();
 sg13g2_fill_2 FILLER_57_124 ();
 sg13g2_fill_1 FILLER_57_126 ();
 sg13g2_fill_2 FILLER_57_142 ();
 sg13g2_fill_2 FILLER_57_149 ();
 sg13g2_fill_1 FILLER_57_151 ();
 sg13g2_fill_2 FILLER_57_158 ();
 sg13g2_fill_1 FILLER_57_160 ();
 sg13g2_fill_2 FILLER_57_166 ();
 sg13g2_fill_1 FILLER_57_168 ();
 sg13g2_fill_1 FILLER_57_182 ();
 sg13g2_fill_1 FILLER_57_191 ();
 sg13g2_fill_1 FILLER_57_205 ();
 sg13g2_fill_2 FILLER_57_217 ();
 sg13g2_fill_2 FILLER_57_245 ();
 sg13g2_fill_1 FILLER_57_273 ();
 sg13g2_decap_8 FILLER_57_284 ();
 sg13g2_fill_2 FILLER_57_314 ();
 sg13g2_fill_2 FILLER_57_320 ();
 sg13g2_fill_1 FILLER_57_326 ();
 sg13g2_fill_2 FILLER_57_337 ();
 sg13g2_fill_2 FILLER_57_369 ();
 sg13g2_decap_8 FILLER_57_375 ();
 sg13g2_fill_1 FILLER_57_382 ();
 sg13g2_decap_4 FILLER_57_390 ();
 sg13g2_fill_1 FILLER_57_405 ();
 sg13g2_decap_4 FILLER_57_419 ();
 sg13g2_fill_1 FILLER_57_423 ();
 sg13g2_fill_2 FILLER_57_428 ();
 sg13g2_fill_1 FILLER_57_430 ();
 sg13g2_decap_4 FILLER_57_441 ();
 sg13g2_fill_2 FILLER_57_464 ();
 sg13g2_fill_2 FILLER_57_505 ();
 sg13g2_fill_2 FILLER_57_519 ();
 sg13g2_fill_2 FILLER_57_526 ();
 sg13g2_fill_1 FILLER_57_537 ();
 sg13g2_fill_1 FILLER_57_551 ();
 sg13g2_fill_1 FILLER_57_557 ();
 sg13g2_fill_1 FILLER_57_562 ();
 sg13g2_fill_2 FILLER_57_567 ();
 sg13g2_fill_1 FILLER_57_596 ();
 sg13g2_fill_1 FILLER_57_601 ();
 sg13g2_fill_1 FILLER_57_609 ();
 sg13g2_fill_2 FILLER_57_641 ();
 sg13g2_fill_1 FILLER_57_643 ();
 sg13g2_fill_1 FILLER_57_656 ();
 sg13g2_fill_1 FILLER_57_671 ();
 sg13g2_fill_1 FILLER_57_682 ();
 sg13g2_fill_2 FILLER_57_687 ();
 sg13g2_fill_2 FILLER_57_711 ();
 sg13g2_fill_1 FILLER_57_713 ();
 sg13g2_fill_1 FILLER_57_719 ();
 sg13g2_fill_2 FILLER_57_726 ();
 sg13g2_fill_1 FILLER_57_742 ();
 sg13g2_fill_1 FILLER_57_770 ();
 sg13g2_decap_4 FILLER_57_794 ();
 sg13g2_fill_1 FILLER_57_798 ();
 sg13g2_fill_1 FILLER_57_819 ();
 sg13g2_fill_1 FILLER_57_829 ();
 sg13g2_fill_1 FILLER_57_840 ();
 sg13g2_fill_2 FILLER_57_845 ();
 sg13g2_decap_8 FILLER_57_852 ();
 sg13g2_decap_8 FILLER_57_859 ();
 sg13g2_decap_8 FILLER_57_866 ();
 sg13g2_decap_4 FILLER_57_873 ();
 sg13g2_fill_1 FILLER_57_877 ();
 sg13g2_fill_2 FILLER_58_42 ();
 sg13g2_decap_4 FILLER_58_47 ();
 sg13g2_fill_1 FILLER_58_65 ();
 sg13g2_fill_1 FILLER_58_71 ();
 sg13g2_fill_1 FILLER_58_81 ();
 sg13g2_fill_1 FILLER_58_92 ();
 sg13g2_fill_1 FILLER_58_99 ();
 sg13g2_fill_1 FILLER_58_105 ();
 sg13g2_fill_1 FILLER_58_114 ();
 sg13g2_fill_1 FILLER_58_128 ();
 sg13g2_fill_1 FILLER_58_139 ();
 sg13g2_decap_4 FILLER_58_146 ();
 sg13g2_decap_4 FILLER_58_160 ();
 sg13g2_fill_2 FILLER_58_164 ();
 sg13g2_fill_1 FILLER_58_174 ();
 sg13g2_fill_1 FILLER_58_180 ();
 sg13g2_fill_2 FILLER_58_209 ();
 sg13g2_fill_2 FILLER_58_217 ();
 sg13g2_fill_1 FILLER_58_219 ();
 sg13g2_fill_1 FILLER_58_233 ();
 sg13g2_fill_2 FILLER_58_255 ();
 sg13g2_fill_1 FILLER_58_257 ();
 sg13g2_fill_2 FILLER_58_274 ();
 sg13g2_fill_1 FILLER_58_276 ();
 sg13g2_fill_1 FILLER_58_282 ();
 sg13g2_decap_4 FILLER_58_292 ();
 sg13g2_fill_2 FILLER_58_296 ();
 sg13g2_fill_2 FILLER_58_315 ();
 sg13g2_fill_1 FILLER_58_317 ();
 sg13g2_fill_1 FILLER_58_323 ();
 sg13g2_fill_2 FILLER_58_329 ();
 sg13g2_fill_2 FILLER_58_361 ();
 sg13g2_fill_1 FILLER_58_363 ();
 sg13g2_fill_2 FILLER_58_395 ();
 sg13g2_fill_2 FILLER_58_405 ();
 sg13g2_fill_2 FILLER_58_457 ();
 sg13g2_fill_1 FILLER_58_464 ();
 sg13g2_fill_1 FILLER_58_469 ();
 sg13g2_fill_1 FILLER_58_480 ();
 sg13g2_decap_4 FILLER_58_507 ();
 sg13g2_fill_2 FILLER_58_511 ();
 sg13g2_fill_2 FILLER_58_519 ();
 sg13g2_fill_1 FILLER_58_521 ();
 sg13g2_fill_2 FILLER_58_526 ();
 sg13g2_fill_1 FILLER_58_532 ();
 sg13g2_fill_1 FILLER_58_547 ();
 sg13g2_fill_1 FILLER_58_566 ();
 sg13g2_decap_4 FILLER_58_628 ();
 sg13g2_fill_2 FILLER_58_651 ();
 sg13g2_fill_1 FILLER_58_663 ();
 sg13g2_fill_2 FILLER_58_678 ();
 sg13g2_fill_2 FILLER_58_713 ();
 sg13g2_fill_1 FILLER_58_715 ();
 sg13g2_fill_2 FILLER_58_748 ();
 sg13g2_decap_4 FILLER_58_755 ();
 sg13g2_fill_1 FILLER_58_759 ();
 sg13g2_fill_2 FILLER_58_770 ();
 sg13g2_fill_2 FILLER_58_791 ();
 sg13g2_fill_1 FILLER_58_834 ();
 sg13g2_fill_2 FILLER_58_844 ();
 sg13g2_fill_2 FILLER_58_850 ();
 sg13g2_decap_8 FILLER_58_860 ();
 sg13g2_decap_8 FILLER_58_867 ();
 sg13g2_decap_4 FILLER_58_874 ();
 sg13g2_decap_4 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_4 ();
 sg13g2_fill_2 FILLER_59_53 ();
 sg13g2_fill_1 FILLER_59_55 ();
 sg13g2_fill_2 FILLER_59_60 ();
 sg13g2_fill_1 FILLER_59_62 ();
 sg13g2_decap_8 FILLER_59_68 ();
 sg13g2_fill_2 FILLER_59_75 ();
 sg13g2_fill_1 FILLER_59_77 ();
 sg13g2_fill_1 FILLER_59_93 ();
 sg13g2_fill_1 FILLER_59_103 ();
 sg13g2_fill_2 FILLER_59_133 ();
 sg13g2_fill_1 FILLER_59_135 ();
 sg13g2_fill_2 FILLER_59_170 ();
 sg13g2_fill_1 FILLER_59_177 ();
 sg13g2_fill_1 FILLER_59_233 ();
 sg13g2_fill_2 FILLER_59_304 ();
 sg13g2_fill_1 FILLER_59_306 ();
 sg13g2_decap_4 FILLER_59_317 ();
 sg13g2_decap_4 FILLER_59_346 ();
 sg13g2_fill_2 FILLER_59_350 ();
 sg13g2_fill_1 FILLER_59_410 ();
 sg13g2_fill_2 FILLER_59_416 ();
 sg13g2_fill_2 FILLER_59_423 ();
 sg13g2_fill_1 FILLER_59_425 ();
 sg13g2_decap_8 FILLER_59_440 ();
 sg13g2_fill_2 FILLER_59_447 ();
 sg13g2_fill_1 FILLER_59_475 ();
 sg13g2_fill_2 FILLER_59_494 ();
 sg13g2_fill_2 FILLER_59_515 ();
 sg13g2_fill_1 FILLER_59_550 ();
 sg13g2_fill_2 FILLER_59_570 ();
 sg13g2_fill_2 FILLER_59_592 ();
 sg13g2_fill_2 FILLER_59_599 ();
 sg13g2_fill_1 FILLER_59_611 ();
 sg13g2_fill_1 FILLER_59_627 ();
 sg13g2_fill_2 FILLER_59_652 ();
 sg13g2_fill_1 FILLER_59_654 ();
 sg13g2_fill_1 FILLER_59_669 ();
 sg13g2_fill_1 FILLER_59_685 ();
 sg13g2_fill_2 FILLER_59_701 ();
 sg13g2_fill_2 FILLER_59_706 ();
 sg13g2_fill_1 FILLER_59_708 ();
 sg13g2_fill_2 FILLER_59_715 ();
 sg13g2_fill_1 FILLER_59_722 ();
 sg13g2_fill_1 FILLER_59_727 ();
 sg13g2_fill_2 FILLER_59_762 ();
 sg13g2_fill_2 FILLER_59_769 ();
 sg13g2_fill_2 FILLER_59_776 ();
 sg13g2_fill_1 FILLER_59_778 ();
 sg13g2_fill_2 FILLER_59_827 ();
 sg13g2_fill_2 FILLER_59_846 ();
 sg13g2_fill_1 FILLER_59_848 ();
 sg13g2_decap_8 FILLER_59_859 ();
 sg13g2_decap_8 FILLER_59_866 ();
 sg13g2_decap_4 FILLER_59_873 ();
 sg13g2_fill_1 FILLER_59_877 ();
 sg13g2_fill_1 FILLER_60_68 ();
 sg13g2_fill_1 FILLER_60_78 ();
 sg13g2_fill_1 FILLER_60_106 ();
 sg13g2_fill_1 FILLER_60_144 ();
 sg13g2_decap_4 FILLER_60_167 ();
 sg13g2_decap_4 FILLER_60_175 ();
 sg13g2_fill_1 FILLER_60_179 ();
 sg13g2_fill_2 FILLER_60_198 ();
 sg13g2_fill_2 FILLER_60_220 ();
 sg13g2_fill_1 FILLER_60_227 ();
 sg13g2_fill_2 FILLER_60_243 ();
 sg13g2_fill_1 FILLER_60_250 ();
 sg13g2_fill_1 FILLER_60_260 ();
 sg13g2_fill_1 FILLER_60_264 ();
 sg13g2_fill_2 FILLER_60_279 ();
 sg13g2_fill_1 FILLER_60_281 ();
 sg13g2_fill_2 FILLER_60_327 ();
 sg13g2_fill_2 FILLER_60_414 ();
 sg13g2_decap_4 FILLER_60_441 ();
 sg13g2_fill_1 FILLER_60_445 ();
 sg13g2_decap_4 FILLER_60_451 ();
 sg13g2_fill_2 FILLER_60_455 ();
 sg13g2_fill_2 FILLER_60_468 ();
 sg13g2_fill_1 FILLER_60_475 ();
 sg13g2_decap_8 FILLER_60_507 ();
 sg13g2_decap_4 FILLER_60_514 ();
 sg13g2_fill_2 FILLER_60_518 ();
 sg13g2_decap_4 FILLER_60_524 ();
 sg13g2_fill_1 FILLER_60_528 ();
 sg13g2_decap_8 FILLER_60_533 ();
 sg13g2_fill_1 FILLER_60_559 ();
 sg13g2_fill_2 FILLER_60_564 ();
 sg13g2_fill_1 FILLER_60_585 ();
 sg13g2_fill_1 FILLER_60_590 ();
 sg13g2_fill_1 FILLER_60_596 ();
 sg13g2_fill_1 FILLER_60_619 ();
 sg13g2_fill_1 FILLER_60_630 ();
 sg13g2_fill_1 FILLER_60_651 ();
 sg13g2_fill_1 FILLER_60_684 ();
 sg13g2_fill_2 FILLER_60_720 ();
 sg13g2_fill_1 FILLER_60_722 ();
 sg13g2_fill_2 FILLER_60_740 ();
 sg13g2_fill_2 FILLER_60_747 ();
 sg13g2_fill_1 FILLER_60_749 ();
 sg13g2_decap_8 FILLER_60_762 ();
 sg13g2_fill_1 FILLER_60_769 ();
 sg13g2_fill_1 FILLER_60_796 ();
 sg13g2_decap_4 FILLER_60_820 ();
 sg13g2_fill_1 FILLER_60_824 ();
 sg13g2_fill_2 FILLER_60_842 ();
 sg13g2_fill_1 FILLER_60_844 ();
 sg13g2_decap_4 FILLER_60_849 ();
 sg13g2_decap_8 FILLER_60_862 ();
 sg13g2_decap_8 FILLER_60_869 ();
 sg13g2_fill_2 FILLER_60_876 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_76 ();
 sg13g2_fill_1 FILLER_61_78 ();
 sg13g2_decap_4 FILLER_61_84 ();
 sg13g2_fill_1 FILLER_61_93 ();
 sg13g2_fill_2 FILLER_61_104 ();
 sg13g2_decap_4 FILLER_61_111 ();
 sg13g2_fill_2 FILLER_61_115 ();
 sg13g2_fill_2 FILLER_61_167 ();
 sg13g2_decap_4 FILLER_61_178 ();
 sg13g2_fill_1 FILLER_61_195 ();
 sg13g2_fill_2 FILLER_61_201 ();
 sg13g2_fill_1 FILLER_61_203 ();
 sg13g2_fill_1 FILLER_61_207 ();
 sg13g2_fill_2 FILLER_61_224 ();
 sg13g2_fill_1 FILLER_61_237 ();
 sg13g2_fill_2 FILLER_61_253 ();
 sg13g2_fill_1 FILLER_61_255 ();
 sg13g2_decap_8 FILLER_61_260 ();
 sg13g2_decap_8 FILLER_61_267 ();
 sg13g2_decap_8 FILLER_61_274 ();
 sg13g2_fill_1 FILLER_61_295 ();
 sg13g2_decap_8 FILLER_61_301 ();
 sg13g2_fill_1 FILLER_61_308 ();
 sg13g2_decap_4 FILLER_61_318 ();
 sg13g2_fill_1 FILLER_61_322 ();
 sg13g2_fill_2 FILLER_61_328 ();
 sg13g2_fill_1 FILLER_61_330 ();
 sg13g2_decap_4 FILLER_61_346 ();
 sg13g2_decap_4 FILLER_61_354 ();
 sg13g2_fill_1 FILLER_61_358 ();
 sg13g2_decap_4 FILLER_61_368 ();
 sg13g2_fill_1 FILLER_61_372 ();
 sg13g2_fill_2 FILLER_61_377 ();
 sg13g2_fill_2 FILLER_61_396 ();
 sg13g2_decap_4 FILLER_61_433 ();
 sg13g2_fill_2 FILLER_61_437 ();
 sg13g2_fill_1 FILLER_61_465 ();
 sg13g2_fill_1 FILLER_61_470 ();
 sg13g2_fill_1 FILLER_61_482 ();
 sg13g2_decap_8 FILLER_61_490 ();
 sg13g2_decap_4 FILLER_61_497 ();
 sg13g2_fill_1 FILLER_61_505 ();
 sg13g2_fill_1 FILLER_61_511 ();
 sg13g2_decap_4 FILLER_61_530 ();
 sg13g2_fill_2 FILLER_61_572 ();
 sg13g2_fill_1 FILLER_61_642 ();
 sg13g2_fill_1 FILLER_61_649 ();
 sg13g2_fill_1 FILLER_61_682 ();
 sg13g2_fill_2 FILLER_61_691 ();
 sg13g2_fill_1 FILLER_61_693 ();
 sg13g2_decap_4 FILLER_61_708 ();
 sg13g2_fill_1 FILLER_61_716 ();
 sg13g2_fill_1 FILLER_61_721 ();
 sg13g2_decap_4 FILLER_61_760 ();
 sg13g2_fill_1 FILLER_61_778 ();
 sg13g2_fill_1 FILLER_61_784 ();
 sg13g2_fill_1 FILLER_61_790 ();
 sg13g2_fill_2 FILLER_61_800 ();
 sg13g2_fill_1 FILLER_61_802 ();
 sg13g2_fill_2 FILLER_61_824 ();
 sg13g2_fill_2 FILLER_61_839 ();
 sg13g2_decap_8 FILLER_61_865 ();
 sg13g2_decap_4 FILLER_61_872 ();
 sg13g2_fill_2 FILLER_61_876 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_7 ();
 sg13g2_decap_4 FILLER_62_43 ();
 sg13g2_fill_1 FILLER_62_47 ();
 sg13g2_decap_4 FILLER_62_64 ();
 sg13g2_decap_4 FILLER_62_77 ();
 sg13g2_fill_1 FILLER_62_81 ();
 sg13g2_fill_2 FILLER_62_86 ();
 sg13g2_fill_1 FILLER_62_88 ();
 sg13g2_fill_1 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_121 ();
 sg13g2_fill_2 FILLER_62_132 ();
 sg13g2_fill_1 FILLER_62_134 ();
 sg13g2_fill_1 FILLER_62_157 ();
 sg13g2_fill_1 FILLER_62_163 ();
 sg13g2_fill_2 FILLER_62_168 ();
 sg13g2_fill_1 FILLER_62_175 ();
 sg13g2_fill_1 FILLER_62_181 ();
 sg13g2_fill_1 FILLER_62_216 ();
 sg13g2_fill_2 FILLER_62_221 ();
 sg13g2_decap_4 FILLER_62_227 ();
 sg13g2_fill_2 FILLER_62_236 ();
 sg13g2_decap_4 FILLER_62_281 ();
 sg13g2_fill_2 FILLER_62_289 ();
 sg13g2_fill_1 FILLER_62_291 ();
 sg13g2_fill_1 FILLER_62_302 ();
 sg13g2_decap_8 FILLER_62_313 ();
 sg13g2_decap_4 FILLER_62_320 ();
 sg13g2_decap_8 FILLER_62_333 ();
 sg13g2_decap_4 FILLER_62_340 ();
 sg13g2_fill_2 FILLER_62_344 ();
 sg13g2_fill_1 FILLER_62_351 ();
 sg13g2_fill_2 FILLER_62_378 ();
 sg13g2_fill_1 FILLER_62_380 ();
 sg13g2_decap_8 FILLER_62_390 ();
 sg13g2_decap_8 FILLER_62_397 ();
 sg13g2_fill_2 FILLER_62_415 ();
 sg13g2_fill_1 FILLER_62_417 ();
 sg13g2_decap_4 FILLER_62_423 ();
 sg13g2_fill_1 FILLER_62_427 ();
 sg13g2_decap_8 FILLER_62_432 ();
 sg13g2_fill_1 FILLER_62_439 ();
 sg13g2_decap_8 FILLER_62_445 ();
 sg13g2_decap_8 FILLER_62_457 ();
 sg13g2_fill_2 FILLER_62_479 ();
 sg13g2_fill_1 FILLER_62_481 ();
 sg13g2_fill_1 FILLER_62_498 ();
 sg13g2_fill_1 FILLER_62_504 ();
 sg13g2_fill_1 FILLER_62_512 ();
 sg13g2_decap_4 FILLER_62_530 ();
 sg13g2_fill_1 FILLER_62_557 ();
 sg13g2_decap_4 FILLER_62_596 ();
 sg13g2_fill_1 FILLER_62_600 ();
 sg13g2_fill_1 FILLER_62_613 ();
 sg13g2_fill_2 FILLER_62_620 ();
 sg13g2_fill_1 FILLER_62_622 ();
 sg13g2_decap_4 FILLER_62_628 ();
 sg13g2_fill_2 FILLER_62_652 ();
 sg13g2_fill_2 FILLER_62_657 ();
 sg13g2_fill_1 FILLER_62_659 ();
 sg13g2_fill_2 FILLER_62_665 ();
 sg13g2_fill_2 FILLER_62_681 ();
 sg13g2_decap_4 FILLER_62_693 ();
 sg13g2_fill_2 FILLER_62_697 ();
 sg13g2_fill_2 FILLER_62_704 ();
 sg13g2_fill_1 FILLER_62_706 ();
 sg13g2_fill_1 FILLER_62_712 ();
 sg13g2_fill_2 FILLER_62_717 ();
 sg13g2_fill_1 FILLER_62_722 ();
 sg13g2_fill_1 FILLER_62_729 ();
 sg13g2_decap_4 FILLER_62_734 ();
 sg13g2_fill_2 FILLER_62_738 ();
 sg13g2_fill_2 FILLER_62_746 ();
 sg13g2_fill_1 FILLER_62_748 ();
 sg13g2_fill_1 FILLER_62_753 ();
 sg13g2_fill_1 FILLER_62_793 ();
 sg13g2_fill_2 FILLER_62_799 ();
 sg13g2_fill_1 FILLER_62_805 ();
 sg13g2_fill_1 FILLER_62_813 ();
 sg13g2_fill_1 FILLER_62_825 ();
 sg13g2_fill_1 FILLER_62_833 ();
 sg13g2_fill_1 FILLER_62_844 ();
 sg13g2_fill_2 FILLER_62_850 ();
 sg13g2_decap_8 FILLER_62_867 ();
 sg13g2_decap_4 FILLER_62_874 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_4 FILLER_63_7 ();
 sg13g2_fill_2 FILLER_63_33 ();
 sg13g2_fill_1 FILLER_63_35 ();
 sg13g2_fill_1 FILLER_63_40 ();
 sg13g2_fill_1 FILLER_63_50 ();
 sg13g2_fill_1 FILLER_63_60 ();
 sg13g2_fill_1 FILLER_63_87 ();
 sg13g2_fill_1 FILLER_63_92 ();
 sg13g2_fill_2 FILLER_63_111 ();
 sg13g2_fill_1 FILLER_63_117 ();
 sg13g2_fill_2 FILLER_63_123 ();
 sg13g2_fill_1 FILLER_63_125 ();
 sg13g2_fill_2 FILLER_63_140 ();
 sg13g2_fill_2 FILLER_63_155 ();
 sg13g2_fill_1 FILLER_63_176 ();
 sg13g2_decap_4 FILLER_63_187 ();
 sg13g2_fill_1 FILLER_63_191 ();
 sg13g2_fill_2 FILLER_63_200 ();
 sg13g2_fill_1 FILLER_63_214 ();
 sg13g2_decap_8 FILLER_63_260 ();
 sg13g2_decap_8 FILLER_63_267 ();
 sg13g2_fill_2 FILLER_63_274 ();
 sg13g2_decap_4 FILLER_63_335 ();
 sg13g2_fill_1 FILLER_63_339 ();
 sg13g2_fill_1 FILLER_63_385 ();
 sg13g2_fill_1 FILLER_63_395 ();
 sg13g2_fill_2 FILLER_63_400 ();
 sg13g2_fill_1 FILLER_63_406 ();
 sg13g2_fill_1 FILLER_63_412 ();
 sg13g2_fill_2 FILLER_63_422 ();
 sg13g2_decap_8 FILLER_63_438 ();
 sg13g2_fill_1 FILLER_63_445 ();
 sg13g2_fill_1 FILLER_63_472 ();
 sg13g2_fill_1 FILLER_63_478 ();
 sg13g2_decap_8 FILLER_63_499 ();
 sg13g2_fill_2 FILLER_63_506 ();
 sg13g2_fill_1 FILLER_63_508 ();
 sg13g2_fill_2 FILLER_63_513 ();
 sg13g2_fill_1 FILLER_63_515 ();
 sg13g2_fill_1 FILLER_63_537 ();
 sg13g2_fill_2 FILLER_63_543 ();
 sg13g2_fill_2 FILLER_63_550 ();
 sg13g2_fill_2 FILLER_63_558 ();
 sg13g2_fill_1 FILLER_63_566 ();
 sg13g2_fill_2 FILLER_63_576 ();
 sg13g2_fill_1 FILLER_63_578 ();
 sg13g2_decap_8 FILLER_63_583 ();
 sg13g2_fill_1 FILLER_63_615 ();
 sg13g2_fill_2 FILLER_63_626 ();
 sg13g2_fill_1 FILLER_63_651 ();
 sg13g2_fill_2 FILLER_63_656 ();
 sg13g2_fill_2 FILLER_63_677 ();
 sg13g2_fill_2 FILLER_63_683 ();
 sg13g2_fill_1 FILLER_63_685 ();
 sg13g2_fill_1 FILLER_63_704 ();
 sg13g2_fill_2 FILLER_63_726 ();
 sg13g2_decap_4 FILLER_63_734 ();
 sg13g2_fill_2 FILLER_63_738 ();
 sg13g2_fill_1 FILLER_63_754 ();
 sg13g2_fill_1 FILLER_63_762 ();
 sg13g2_fill_2 FILLER_63_773 ();
 sg13g2_fill_2 FILLER_63_780 ();
 sg13g2_fill_2 FILLER_63_794 ();
 sg13g2_fill_1 FILLER_63_799 ();
 sg13g2_fill_2 FILLER_63_810 ();
 sg13g2_fill_1 FILLER_63_812 ();
 sg13g2_fill_2 FILLER_63_838 ();
 sg13g2_fill_1 FILLER_63_855 ();
 sg13g2_fill_2 FILLER_63_860 ();
 sg13g2_fill_1 FILLER_63_862 ();
 sg13g2_fill_1 FILLER_63_868 ();
 sg13g2_decap_4 FILLER_63_874 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_7 ();
 sg13g2_fill_1 FILLER_64_53 ();
 sg13g2_fill_1 FILLER_64_59 ();
 sg13g2_decap_4 FILLER_64_65 ();
 sg13g2_fill_1 FILLER_64_69 ();
 sg13g2_decap_4 FILLER_64_74 ();
 sg13g2_decap_8 FILLER_64_89 ();
 sg13g2_fill_1 FILLER_64_96 ();
 sg13g2_fill_1 FILLER_64_101 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_fill_1 FILLER_64_117 ();
 sg13g2_fill_1 FILLER_64_149 ();
 sg13g2_fill_1 FILLER_64_184 ();
 sg13g2_fill_2 FILLER_64_193 ();
 sg13g2_fill_1 FILLER_64_199 ();
 sg13g2_decap_8 FILLER_64_204 ();
 sg13g2_decap_4 FILLER_64_211 ();
 sg13g2_fill_1 FILLER_64_226 ();
 sg13g2_fill_2 FILLER_64_233 ();
 sg13g2_fill_1 FILLER_64_243 ();
 sg13g2_fill_1 FILLER_64_252 ();
 sg13g2_fill_2 FILLER_64_256 ();
 sg13g2_fill_2 FILLER_64_281 ();
 sg13g2_fill_2 FILLER_64_291 ();
 sg13g2_fill_1 FILLER_64_293 ();
 sg13g2_fill_1 FILLER_64_303 ();
 sg13g2_decap_8 FILLER_64_340 ();
 sg13g2_fill_1 FILLER_64_347 ();
 sg13g2_fill_2 FILLER_64_353 ();
 sg13g2_fill_2 FILLER_64_363 ();
 sg13g2_fill_1 FILLER_64_365 ();
 sg13g2_fill_2 FILLER_64_377 ();
 sg13g2_fill_1 FILLER_64_426 ();
 sg13g2_decap_4 FILLER_64_458 ();
 sg13g2_fill_2 FILLER_64_470 ();
 sg13g2_fill_2 FILLER_64_482 ();
 sg13g2_fill_1 FILLER_64_484 ();
 sg13g2_decap_8 FILLER_64_491 ();
 sg13g2_decap_8 FILLER_64_498 ();
 sg13g2_fill_2 FILLER_64_505 ();
 sg13g2_decap_8 FILLER_64_516 ();
 sg13g2_decap_4 FILLER_64_523 ();
 sg13g2_fill_2 FILLER_64_533 ();
 sg13g2_fill_1 FILLER_64_544 ();
 sg13g2_fill_1 FILLER_64_550 ();
 sg13g2_fill_1 FILLER_64_561 ();
 sg13g2_decap_4 FILLER_64_569 ();
 sg13g2_fill_1 FILLER_64_573 ();
 sg13g2_fill_1 FILLER_64_578 ();
 sg13g2_fill_1 FILLER_64_584 ();
 sg13g2_fill_1 FILLER_64_590 ();
 sg13g2_fill_1 FILLER_64_596 ();
 sg13g2_fill_1 FILLER_64_603 ();
 sg13g2_decap_4 FILLER_64_624 ();
 sg13g2_fill_1 FILLER_64_628 ();
 sg13g2_decap_4 FILLER_64_641 ();
 sg13g2_fill_2 FILLER_64_664 ();
 sg13g2_fill_2 FILLER_64_684 ();
 sg13g2_fill_1 FILLER_64_690 ();
 sg13g2_fill_2 FILLER_64_701 ();
 sg13g2_fill_1 FILLER_64_703 ();
 sg13g2_fill_1 FILLER_64_716 ();
 sg13g2_fill_1 FILLER_64_729 ();
 sg13g2_fill_1 FILLER_64_736 ();
 sg13g2_fill_1 FILLER_64_743 ();
 sg13g2_fill_1 FILLER_64_748 ();
 sg13g2_fill_1 FILLER_64_758 ();
 sg13g2_decap_4 FILLER_64_800 ();
 sg13g2_fill_2 FILLER_64_809 ();
 sg13g2_fill_1 FILLER_64_833 ();
 sg13g2_fill_2 FILLER_64_850 ();
 sg13g2_fill_1 FILLER_64_852 ();
 sg13g2_fill_2 FILLER_64_858 ();
 sg13g2_fill_1 FILLER_64_860 ();
 sg13g2_fill_2 FILLER_64_871 ();
 sg13g2_fill_1 FILLER_64_873 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_9 ();
 sg13g2_fill_1 FILLER_65_39 ();
 sg13g2_fill_1 FILLER_65_48 ();
 sg13g2_fill_1 FILLER_65_53 ();
 sg13g2_fill_2 FILLER_65_95 ();
 sg13g2_fill_1 FILLER_65_97 ();
 sg13g2_fill_1 FILLER_65_108 ();
 sg13g2_fill_2 FILLER_65_124 ();
 sg13g2_fill_1 FILLER_65_126 ();
 sg13g2_fill_1 FILLER_65_141 ();
 sg13g2_fill_2 FILLER_65_153 ();
 sg13g2_fill_1 FILLER_65_213 ();
 sg13g2_fill_1 FILLER_65_223 ();
 sg13g2_fill_2 FILLER_65_234 ();
 sg13g2_decap_4 FILLER_65_260 ();
 sg13g2_fill_1 FILLER_65_264 ();
 sg13g2_fill_2 FILLER_65_280 ();
 sg13g2_fill_1 FILLER_65_282 ();
 sg13g2_fill_2 FILLER_65_299 ();
 sg13g2_fill_2 FILLER_65_309 ();
 sg13g2_fill_2 FILLER_65_324 ();
 sg13g2_decap_8 FILLER_65_337 ();
 sg13g2_fill_1 FILLER_65_354 ();
 sg13g2_fill_1 FILLER_65_363 ();
 sg13g2_fill_2 FILLER_65_395 ();
 sg13g2_fill_1 FILLER_65_401 ();
 sg13g2_fill_2 FILLER_65_406 ();
 sg13g2_decap_4 FILLER_65_427 ();
 sg13g2_fill_2 FILLER_65_431 ();
 sg13g2_fill_1 FILLER_65_441 ();
 sg13g2_fill_2 FILLER_65_451 ();
 sg13g2_decap_8 FILLER_65_459 ();
 sg13g2_fill_2 FILLER_65_466 ();
 sg13g2_decap_4 FILLER_65_482 ();
 sg13g2_decap_4 FILLER_65_490 ();
 sg13g2_fill_2 FILLER_65_506 ();
 sg13g2_fill_1 FILLER_65_508 ();
 sg13g2_fill_2 FILLER_65_517 ();
 sg13g2_decap_4 FILLER_65_533 ();
 sg13g2_fill_2 FILLER_65_557 ();
 sg13g2_fill_1 FILLER_65_559 ();
 sg13g2_decap_8 FILLER_65_591 ();
 sg13g2_fill_1 FILLER_65_598 ();
 sg13g2_fill_1 FILLER_65_613 ();
 sg13g2_decap_8 FILLER_65_629 ();
 sg13g2_fill_2 FILLER_65_661 ();
 sg13g2_fill_1 FILLER_65_696 ();
 sg13g2_fill_1 FILLER_65_726 ();
 sg13g2_fill_2 FILLER_65_731 ();
 sg13g2_decap_4 FILLER_65_738 ();
 sg13g2_fill_2 FILLER_65_792 ();
 sg13g2_fill_1 FILLER_65_798 ();
 sg13g2_fill_2 FILLER_65_819 ();
 sg13g2_fill_1 FILLER_65_856 ();
 sg13g2_fill_2 FILLER_65_866 ();
 sg13g2_decap_4 FILLER_65_873 ();
 sg13g2_fill_1 FILLER_65_877 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_7 ();
 sg13g2_fill_2 FILLER_66_11 ();
 sg13g2_fill_2 FILLER_66_56 ();
 sg13g2_fill_1 FILLER_66_67 ();
 sg13g2_decap_4 FILLER_66_72 ();
 sg13g2_decap_4 FILLER_66_80 ();
 sg13g2_fill_2 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_90 ();
 sg13g2_decap_8 FILLER_66_97 ();
 sg13g2_fill_1 FILLER_66_104 ();
 sg13g2_fill_2 FILLER_66_126 ();
 sg13g2_fill_1 FILLER_66_128 ();
 sg13g2_fill_1 FILLER_66_148 ();
 sg13g2_fill_2 FILLER_66_190 ();
 sg13g2_fill_1 FILLER_66_203 ();
 sg13g2_fill_1 FILLER_66_209 ();
 sg13g2_fill_2 FILLER_66_247 ();
 sg13g2_fill_1 FILLER_66_257 ();
 sg13g2_fill_2 FILLER_66_299 ();
 sg13g2_fill_1 FILLER_66_374 ();
 sg13g2_fill_2 FILLER_66_379 ();
 sg13g2_fill_2 FILLER_66_385 ();
 sg13g2_fill_1 FILLER_66_392 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_fill_1 FILLER_66_414 ();
 sg13g2_fill_2 FILLER_66_419 ();
 sg13g2_fill_2 FILLER_66_439 ();
 sg13g2_fill_1 FILLER_66_441 ();
 sg13g2_fill_1 FILLER_66_473 ();
 sg13g2_fill_1 FILLER_66_503 ();
 sg13g2_decap_8 FILLER_66_512 ();
 sg13g2_fill_2 FILLER_66_524 ();
 sg13g2_fill_1 FILLER_66_526 ();
 sg13g2_fill_2 FILLER_66_553 ();
 sg13g2_fill_1 FILLER_66_559 ();
 sg13g2_decap_4 FILLER_66_565 ();
 sg13g2_fill_1 FILLER_66_569 ();
 sg13g2_fill_2 FILLER_66_575 ();
 sg13g2_fill_2 FILLER_66_620 ();
 sg13g2_fill_1 FILLER_66_643 ();
 sg13g2_fill_1 FILLER_66_652 ();
 sg13g2_fill_1 FILLER_66_658 ();
 sg13g2_fill_2 FILLER_66_664 ();
 sg13g2_fill_2 FILLER_66_670 ();
 sg13g2_fill_1 FILLER_66_672 ();
 sg13g2_fill_1 FILLER_66_685 ();
 sg13g2_fill_1 FILLER_66_702 ();
 sg13g2_fill_1 FILLER_66_729 ();
 sg13g2_decap_4 FILLER_66_754 ();
 sg13g2_fill_1 FILLER_66_758 ();
 sg13g2_fill_1 FILLER_66_764 ();
 sg13g2_fill_1 FILLER_66_786 ();
 sg13g2_fill_2 FILLER_66_807 ();
 sg13g2_fill_1 FILLER_66_814 ();
 sg13g2_fill_1 FILLER_66_819 ();
 sg13g2_decap_8 FILLER_66_870 ();
 sg13g2_fill_1 FILLER_66_877 ();
 sg13g2_fill_1 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_27 ();
 sg13g2_decap_8 FILLER_67_32 ();
 sg13g2_fill_2 FILLER_67_65 ();
 sg13g2_fill_1 FILLER_67_89 ();
 sg13g2_fill_1 FILLER_67_123 ();
 sg13g2_fill_1 FILLER_67_134 ();
 sg13g2_fill_1 FILLER_67_140 ();
 sg13g2_fill_1 FILLER_67_163 ();
 sg13g2_decap_4 FILLER_67_170 ();
 sg13g2_fill_1 FILLER_67_192 ();
 sg13g2_fill_2 FILLER_67_206 ();
 sg13g2_fill_2 FILLER_67_220 ();
 sg13g2_fill_1 FILLER_67_222 ();
 sg13g2_decap_8 FILLER_67_258 ();
 sg13g2_decap_4 FILLER_67_275 ();
 sg13g2_fill_2 FILLER_67_279 ();
 sg13g2_fill_2 FILLER_67_302 ();
 sg13g2_fill_1 FILLER_67_304 ();
 sg13g2_fill_1 FILLER_67_332 ();
 sg13g2_decap_4 FILLER_67_339 ();
 sg13g2_fill_2 FILLER_67_370 ();
 sg13g2_fill_1 FILLER_67_372 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_fill_2 FILLER_67_446 ();
 sg13g2_fill_1 FILLER_67_448 ();
 sg13g2_fill_1 FILLER_67_458 ();
 sg13g2_fill_2 FILLER_67_469 ();
 sg13g2_fill_1 FILLER_67_471 ();
 sg13g2_fill_2 FILLER_67_476 ();
 sg13g2_fill_1 FILLER_67_478 ();
 sg13g2_decap_4 FILLER_67_494 ();
 sg13g2_fill_2 FILLER_67_515 ();
 sg13g2_fill_1 FILLER_67_517 ();
 sg13g2_decap_4 FILLER_67_524 ();
 sg13g2_decap_4 FILLER_67_531 ();
 sg13g2_fill_2 FILLER_67_535 ();
 sg13g2_fill_2 FILLER_67_554 ();
 sg13g2_fill_1 FILLER_67_556 ();
 sg13g2_fill_1 FILLER_67_562 ();
 sg13g2_decap_4 FILLER_67_570 ();
 sg13g2_fill_2 FILLER_67_579 ();
 sg13g2_fill_1 FILLER_67_581 ();
 sg13g2_fill_2 FILLER_67_613 ();
 sg13g2_fill_1 FILLER_67_634 ();
 sg13g2_fill_2 FILLER_67_639 ();
 sg13g2_fill_2 FILLER_67_655 ();
 sg13g2_fill_2 FILLER_67_676 ();
 sg13g2_fill_1 FILLER_67_688 ();
 sg13g2_fill_1 FILLER_67_693 ();
 sg13g2_fill_2 FILLER_67_699 ();
 sg13g2_fill_1 FILLER_67_710 ();
 sg13g2_decap_8 FILLER_67_720 ();
 sg13g2_fill_2 FILLER_67_727 ();
 sg13g2_fill_1 FILLER_67_729 ();
 sg13g2_fill_2 FILLER_67_738 ();
 sg13g2_fill_2 FILLER_67_772 ();
 sg13g2_fill_1 FILLER_67_779 ();
 sg13g2_fill_1 FILLER_67_785 ();
 sg13g2_fill_1 FILLER_67_796 ();
 sg13g2_fill_1 FILLER_67_805 ();
 sg13g2_fill_2 FILLER_67_811 ();
 sg13g2_fill_1 FILLER_67_817 ();
 sg13g2_fill_1 FILLER_67_822 ();
 sg13g2_fill_2 FILLER_67_827 ();
 sg13g2_fill_2 FILLER_67_875 ();
 sg13g2_fill_1 FILLER_67_877 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_fill_1 FILLER_68_14 ();
 sg13g2_fill_1 FILLER_68_19 ();
 sg13g2_fill_1 FILLER_68_24 ();
 sg13g2_fill_2 FILLER_68_33 ();
 sg13g2_fill_1 FILLER_68_39 ();
 sg13g2_fill_2 FILLER_68_45 ();
 sg13g2_fill_1 FILLER_68_73 ();
 sg13g2_fill_1 FILLER_68_79 ();
 sg13g2_decap_8 FILLER_68_95 ();
 sg13g2_fill_1 FILLER_68_102 ();
 sg13g2_decap_4 FILLER_68_108 ();
 sg13g2_fill_1 FILLER_68_112 ();
 sg13g2_fill_1 FILLER_68_137 ();
 sg13g2_decap_4 FILLER_68_152 ();
 sg13g2_decap_4 FILLER_68_161 ();
 sg13g2_decap_4 FILLER_68_186 ();
 sg13g2_fill_2 FILLER_68_190 ();
 sg13g2_fill_1 FILLER_68_197 ();
 sg13g2_fill_1 FILLER_68_210 ();
 sg13g2_decap_4 FILLER_68_219 ();
 sg13g2_fill_1 FILLER_68_223 ();
 sg13g2_fill_2 FILLER_68_240 ();
 sg13g2_decap_8 FILLER_68_316 ();
 sg13g2_fill_2 FILLER_68_323 ();
 sg13g2_fill_1 FILLER_68_325 ();
 sg13g2_fill_1 FILLER_68_399 ();
 sg13g2_fill_2 FILLER_68_405 ();
 sg13g2_fill_2 FILLER_68_411 ();
 sg13g2_fill_2 FILLER_68_426 ();
 sg13g2_fill_1 FILLER_68_428 ();
 sg13g2_fill_2 FILLER_68_434 ();
 sg13g2_fill_1 FILLER_68_436 ();
 sg13g2_fill_1 FILLER_68_458 ();
 sg13g2_fill_1 FILLER_68_493 ();
 sg13g2_fill_1 FILLER_68_505 ();
 sg13g2_fill_1 FILLER_68_510 ();
 sg13g2_fill_1 FILLER_68_515 ();
 sg13g2_fill_2 FILLER_68_535 ();
 sg13g2_fill_1 FILLER_68_537 ();
 sg13g2_decap_8 FILLER_68_551 ();
 sg13g2_fill_2 FILLER_68_563 ();
 sg13g2_fill_1 FILLER_68_565 ();
 sg13g2_fill_2 FILLER_68_576 ();
 sg13g2_fill_2 FILLER_68_606 ();
 sg13g2_fill_2 FILLER_68_619 ();
 sg13g2_fill_2 FILLER_68_627 ();
 sg13g2_fill_1 FILLER_68_629 ();
 sg13g2_fill_1 FILLER_68_634 ();
 sg13g2_fill_1 FILLER_68_641 ();
 sg13g2_fill_1 FILLER_68_649 ();
 sg13g2_fill_1 FILLER_68_660 ();
 sg13g2_fill_1 FILLER_68_667 ();
 sg13g2_fill_1 FILLER_68_673 ();
 sg13g2_fill_2 FILLER_68_681 ();
 sg13g2_fill_1 FILLER_68_683 ();
 sg13g2_decap_4 FILLER_68_689 ();
 sg13g2_fill_1 FILLER_68_701 ();
 sg13g2_fill_2 FILLER_68_711 ();
 sg13g2_fill_1 FILLER_68_713 ();
 sg13g2_fill_1 FILLER_68_724 ();
 sg13g2_fill_1 FILLER_68_729 ();
 sg13g2_fill_1 FILLER_68_748 ();
 sg13g2_fill_2 FILLER_68_754 ();
 sg13g2_fill_1 FILLER_68_761 ();
 sg13g2_fill_2 FILLER_68_785 ();
 sg13g2_fill_2 FILLER_68_800 ();
 sg13g2_fill_1 FILLER_68_802 ();
 sg13g2_fill_1 FILLER_68_819 ();
 sg13g2_fill_1 FILLER_68_825 ();
 sg13g2_fill_1 FILLER_68_831 ();
 sg13g2_fill_2 FILLER_68_871 ();
 sg13g2_fill_1 FILLER_68_873 ();
 sg13g2_decap_4 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_4 ();
 sg13g2_fill_1 FILLER_69_28 ();
 sg13g2_fill_1 FILLER_69_37 ();
 sg13g2_fill_1 FILLER_69_48 ();
 sg13g2_fill_1 FILLER_69_55 ();
 sg13g2_fill_2 FILLER_69_74 ();
 sg13g2_fill_1 FILLER_69_81 ();
 sg13g2_fill_1 FILLER_69_87 ();
 sg13g2_fill_1 FILLER_69_114 ();
 sg13g2_fill_1 FILLER_69_123 ();
 sg13g2_fill_1 FILLER_69_129 ();
 sg13g2_fill_2 FILLER_69_142 ();
 sg13g2_fill_2 FILLER_69_149 ();
 sg13g2_fill_1 FILLER_69_151 ();
 sg13g2_decap_8 FILLER_69_157 ();
 sg13g2_decap_8 FILLER_69_164 ();
 sg13g2_decap_4 FILLER_69_171 ();
 sg13g2_fill_1 FILLER_69_175 ();
 sg13g2_decap_8 FILLER_69_186 ();
 sg13g2_fill_1 FILLER_69_206 ();
 sg13g2_decap_4 FILLER_69_212 ();
 sg13g2_fill_2 FILLER_69_216 ();
 sg13g2_decap_4 FILLER_69_226 ();
 sg13g2_fill_1 FILLER_69_230 ();
 sg13g2_fill_2 FILLER_69_248 ();
 sg13g2_fill_1 FILLER_69_254 ();
 sg13g2_fill_1 FILLER_69_296 ();
 sg13g2_fill_1 FILLER_69_301 ();
 sg13g2_fill_2 FILLER_69_306 ();
 sg13g2_decap_8 FILLER_69_320 ();
 sg13g2_fill_2 FILLER_69_327 ();
 sg13g2_decap_8 FILLER_69_334 ();
 sg13g2_decap_8 FILLER_69_341 ();
 sg13g2_fill_1 FILLER_69_348 ();
 sg13g2_fill_2 FILLER_69_363 ();
 sg13g2_fill_2 FILLER_69_373 ();
 sg13g2_fill_1 FILLER_69_375 ();
 sg13g2_fill_2 FILLER_69_386 ();
 sg13g2_decap_8 FILLER_69_406 ();
 sg13g2_decap_8 FILLER_69_418 ();
 sg13g2_decap_4 FILLER_69_425 ();
 sg13g2_fill_2 FILLER_69_429 ();
 sg13g2_decap_8 FILLER_69_435 ();
 sg13g2_fill_2 FILLER_69_446 ();
 sg13g2_fill_1 FILLER_69_448 ();
 sg13g2_fill_1 FILLER_69_457 ();
 sg13g2_decap_8 FILLER_69_466 ();
 sg13g2_decap_4 FILLER_69_473 ();
 sg13g2_decap_8 FILLER_69_494 ();
 sg13g2_fill_1 FILLER_69_501 ();
 sg13g2_fill_2 FILLER_69_506 ();
 sg13g2_fill_2 FILLER_69_548 ();
 sg13g2_fill_2 FILLER_69_559 ();
 sg13g2_fill_1 FILLER_69_561 ();
 sg13g2_fill_2 FILLER_69_581 ();
 sg13g2_fill_1 FILLER_69_583 ();
 sg13g2_fill_1 FILLER_69_590 ();
 sg13g2_fill_1 FILLER_69_595 ();
 sg13g2_fill_1 FILLER_69_609 ();
 sg13g2_fill_2 FILLER_69_615 ();
 sg13g2_fill_1 FILLER_69_632 ();
 sg13g2_fill_1 FILLER_69_678 ();
 sg13g2_fill_1 FILLER_69_699 ();
 sg13g2_fill_2 FILLER_69_712 ();
 sg13g2_fill_1 FILLER_69_714 ();
 sg13g2_fill_1 FILLER_69_726 ();
 sg13g2_fill_1 FILLER_69_732 ();
 sg13g2_fill_2 FILLER_69_738 ();
 sg13g2_fill_1 FILLER_69_754 ();
 sg13g2_fill_1 FILLER_69_759 ();
 sg13g2_fill_1 FILLER_69_772 ();
 sg13g2_fill_1 FILLER_69_777 ();
 sg13g2_fill_1 FILLER_69_781 ();
 sg13g2_fill_1 FILLER_69_786 ();
 sg13g2_fill_1 FILLER_69_792 ();
 sg13g2_fill_1 FILLER_69_802 ();
 sg13g2_fill_1 FILLER_69_838 ();
 sg13g2_fill_2 FILLER_69_860 ();
 sg13g2_fill_2 FILLER_69_875 ();
 sg13g2_fill_1 FILLER_69_877 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_17 ();
 sg13g2_decap_4 FILLER_70_35 ();
 sg13g2_fill_1 FILLER_70_39 ();
 sg13g2_fill_1 FILLER_70_67 ();
 sg13g2_fill_1 FILLER_70_80 ();
 sg13g2_fill_1 FILLER_70_98 ();
 sg13g2_fill_1 FILLER_70_111 ();
 sg13g2_decap_4 FILLER_70_132 ();
 sg13g2_fill_1 FILLER_70_139 ();
 sg13g2_fill_2 FILLER_70_154 ();
 sg13g2_fill_2 FILLER_70_161 ();
 sg13g2_fill_1 FILLER_70_163 ();
 sg13g2_fill_2 FILLER_70_198 ();
 sg13g2_fill_1 FILLER_70_200 ();
 sg13g2_fill_2 FILLER_70_209 ();
 sg13g2_fill_2 FILLER_70_226 ();
 sg13g2_fill_1 FILLER_70_228 ();
 sg13g2_decap_4 FILLER_70_239 ();
 sg13g2_fill_1 FILLER_70_243 ();
 sg13g2_decap_8 FILLER_70_267 ();
 sg13g2_fill_1 FILLER_70_274 ();
 sg13g2_fill_1 FILLER_70_284 ();
 sg13g2_decap_4 FILLER_70_309 ();
 sg13g2_decap_4 FILLER_70_339 ();
 sg13g2_fill_1 FILLER_70_343 ();
 sg13g2_fill_2 FILLER_70_360 ();
 sg13g2_fill_1 FILLER_70_362 ();
 sg13g2_fill_1 FILLER_70_370 ();
 sg13g2_decap_8 FILLER_70_417 ();
 sg13g2_decap_8 FILLER_70_428 ();
 sg13g2_decap_4 FILLER_70_435 ();
 sg13g2_fill_1 FILLER_70_439 ();
 sg13g2_fill_1 FILLER_70_475 ();
 sg13g2_fill_1 FILLER_70_488 ();
 sg13g2_decap_4 FILLER_70_498 ();
 sg13g2_fill_1 FILLER_70_502 ();
 sg13g2_fill_2 FILLER_70_532 ();
 sg13g2_fill_1 FILLER_70_538 ();
 sg13g2_fill_1 FILLER_70_566 ();
 sg13g2_fill_2 FILLER_70_573 ();
 sg13g2_fill_2 FILLER_70_599 ();
 sg13g2_fill_1 FILLER_70_622 ();
 sg13g2_fill_2 FILLER_70_634 ();
 sg13g2_fill_1 FILLER_70_645 ();
 sg13g2_fill_1 FILLER_70_652 ();
 sg13g2_decap_4 FILLER_70_661 ();
 sg13g2_fill_1 FILLER_70_670 ();
 sg13g2_fill_1 FILLER_70_676 ();
 sg13g2_fill_1 FILLER_70_681 ();
 sg13g2_fill_1 FILLER_70_687 ();
 sg13g2_fill_1 FILLER_70_710 ();
 sg13g2_fill_2 FILLER_70_731 ();
 sg13g2_fill_1 FILLER_70_738 ();
 sg13g2_fill_1 FILLER_70_757 ();
 sg13g2_fill_2 FILLER_70_788 ();
 sg13g2_fill_1 FILLER_70_808 ();
 sg13g2_fill_1 FILLER_70_823 ();
 sg13g2_fill_1 FILLER_70_829 ();
 sg13g2_fill_1 FILLER_70_833 ();
 sg13g2_fill_2 FILLER_70_846 ();
 sg13g2_fill_1 FILLER_70_853 ();
 sg13g2_decap_8 FILLER_70_867 ();
 sg13g2_decap_4 FILLER_70_874 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_7 ();
 sg13g2_decap_4 FILLER_71_34 ();
 sg13g2_fill_2 FILLER_71_60 ();
 sg13g2_fill_1 FILLER_71_62 ();
 sg13g2_fill_2 FILLER_71_71 ();
 sg13g2_fill_1 FILLER_71_73 ();
 sg13g2_decap_8 FILLER_71_100 ();
 sg13g2_decap_4 FILLER_71_107 ();
 sg13g2_fill_1 FILLER_71_111 ();
 sg13g2_fill_2 FILLER_71_116 ();
 sg13g2_fill_1 FILLER_71_118 ();
 sg13g2_decap_4 FILLER_71_128 ();
 sg13g2_fill_1 FILLER_71_132 ();
 sg13g2_fill_2 FILLER_71_148 ();
 sg13g2_fill_1 FILLER_71_160 ();
 sg13g2_fill_1 FILLER_71_166 ();
 sg13g2_decap_8 FILLER_71_176 ();
 sg13g2_decap_4 FILLER_71_261 ();
 sg13g2_fill_2 FILLER_71_265 ();
 sg13g2_fill_2 FILLER_71_271 ();
 sg13g2_fill_1 FILLER_71_277 ();
 sg13g2_fill_1 FILLER_71_295 ();
 sg13g2_fill_1 FILLER_71_314 ();
 sg13g2_decap_4 FILLER_71_341 ();
 sg13g2_fill_2 FILLER_71_376 ();
 sg13g2_decap_8 FILLER_71_383 ();
 sg13g2_fill_1 FILLER_71_399 ();
 sg13g2_fill_2 FILLER_71_405 ();
 sg13g2_fill_1 FILLER_71_407 ();
 sg13g2_fill_1 FILLER_71_413 ();
 sg13g2_fill_2 FILLER_71_418 ();
 sg13g2_fill_2 FILLER_71_463 ();
 sg13g2_decap_8 FILLER_71_509 ();
 sg13g2_decap_8 FILLER_71_516 ();
 sg13g2_decap_8 FILLER_71_523 ();
 sg13g2_fill_1 FILLER_71_530 ();
 sg13g2_fill_2 FILLER_71_553 ();
 sg13g2_fill_1 FILLER_71_564 ();
 sg13g2_decap_4 FILLER_71_581 ();
 sg13g2_fill_1 FILLER_71_585 ();
 sg13g2_fill_2 FILLER_71_609 ();
 sg13g2_fill_1 FILLER_71_616 ();
 sg13g2_decap_4 FILLER_71_631 ();
 sg13g2_fill_1 FILLER_71_635 ();
 sg13g2_fill_2 FILLER_71_641 ();
 sg13g2_fill_2 FILLER_71_657 ();
 sg13g2_fill_1 FILLER_71_659 ();
 sg13g2_fill_2 FILLER_71_681 ();
 sg13g2_fill_1 FILLER_71_687 ();
 sg13g2_fill_1 FILLER_71_692 ();
 sg13g2_fill_2 FILLER_71_698 ();
 sg13g2_decap_4 FILLER_71_714 ();
 sg13g2_fill_1 FILLER_71_718 ();
 sg13g2_fill_1 FILLER_71_746 ();
 sg13g2_fill_2 FILLER_71_772 ();
 sg13g2_fill_1 FILLER_71_778 ();
 sg13g2_fill_2 FILLER_71_802 ();
 sg13g2_fill_1 FILLER_71_808 ();
 sg13g2_fill_2 FILLER_71_814 ();
 sg13g2_decap_4 FILLER_71_846 ();
 sg13g2_fill_2 FILLER_71_859 ();
 sg13g2_decap_8 FILLER_71_866 ();
 sg13g2_decap_4 FILLER_71_873 ();
 sg13g2_fill_1 FILLER_71_877 ();
 sg13g2_fill_2 FILLER_72_60 ();
 sg13g2_fill_2 FILLER_72_82 ();
 sg13g2_fill_1 FILLER_72_84 ();
 sg13g2_decap_4 FILLER_72_90 ();
 sg13g2_fill_2 FILLER_72_94 ();
 sg13g2_decap_4 FILLER_72_126 ();
 sg13g2_fill_1 FILLER_72_130 ();
 sg13g2_decap_8 FILLER_72_135 ();
 sg13g2_decap_8 FILLER_72_142 ();
 sg13g2_fill_2 FILLER_72_149 ();
 sg13g2_fill_1 FILLER_72_156 ();
 sg13g2_fill_1 FILLER_72_177 ();
 sg13g2_fill_2 FILLER_72_193 ();
 sg13g2_fill_2 FILLER_72_206 ();
 sg13g2_fill_1 FILLER_72_208 ();
 sg13g2_fill_1 FILLER_72_214 ();
 sg13g2_decap_8 FILLER_72_229 ();
 sg13g2_decap_4 FILLER_72_250 ();
 sg13g2_fill_2 FILLER_72_308 ();
 sg13g2_fill_1 FILLER_72_310 ();
 sg13g2_decap_4 FILLER_72_316 ();
 sg13g2_fill_2 FILLER_72_333 ();
 sg13g2_decap_8 FILLER_72_340 ();
 sg13g2_decap_4 FILLER_72_347 ();
 sg13g2_fill_2 FILLER_72_351 ();
 sg13g2_fill_1 FILLER_72_364 ();
 sg13g2_fill_1 FILLER_72_374 ();
 sg13g2_decap_4 FILLER_72_379 ();
 sg13g2_fill_1 FILLER_72_390 ();
 sg13g2_decap_4 FILLER_72_417 ();
 sg13g2_fill_1 FILLER_72_421 ();
 sg13g2_decap_4 FILLER_72_430 ();
 sg13g2_fill_2 FILLER_72_434 ();
 sg13g2_fill_2 FILLER_72_443 ();
 sg13g2_fill_1 FILLER_72_445 ();
 sg13g2_decap_8 FILLER_72_466 ();
 sg13g2_decap_4 FILLER_72_473 ();
 sg13g2_fill_1 FILLER_72_481 ();
 sg13g2_fill_2 FILLER_72_486 ();
 sg13g2_fill_1 FILLER_72_502 ();
 sg13g2_fill_2 FILLER_72_507 ();
 sg13g2_fill_1 FILLER_72_514 ();
 sg13g2_decap_4 FILLER_72_521 ();
 sg13g2_fill_1 FILLER_72_525 ();
 sg13g2_fill_1 FILLER_72_535 ();
 sg13g2_fill_2 FILLER_72_539 ();
 sg13g2_decap_4 FILLER_72_545 ();
 sg13g2_decap_4 FILLER_72_559 ();
 sg13g2_decap_4 FILLER_72_572 ();
 sg13g2_fill_2 FILLER_72_576 ();
 sg13g2_decap_8 FILLER_72_583 ();
 sg13g2_fill_2 FILLER_72_590 ();
 sg13g2_fill_1 FILLER_72_596 ();
 sg13g2_decap_4 FILLER_72_611 ();
 sg13g2_fill_1 FILLER_72_615 ();
 sg13g2_fill_1 FILLER_72_646 ();
 sg13g2_fill_2 FILLER_72_660 ();
 sg13g2_fill_1 FILLER_72_662 ();
 sg13g2_fill_2 FILLER_72_670 ();
 sg13g2_fill_1 FILLER_72_672 ();
 sg13g2_fill_1 FILLER_72_683 ();
 sg13g2_fill_1 FILLER_72_690 ();
 sg13g2_fill_1 FILLER_72_705 ();
 sg13g2_fill_1 FILLER_72_711 ();
 sg13g2_fill_1 FILLER_72_731 ();
 sg13g2_fill_1 FILLER_72_743 ();
 sg13g2_fill_1 FILLER_72_758 ();
 sg13g2_fill_1 FILLER_72_764 ();
 sg13g2_fill_1 FILLER_72_774 ();
 sg13g2_fill_1 FILLER_72_780 ();
 sg13g2_fill_2 FILLER_72_790 ();
 sg13g2_fill_1 FILLER_72_812 ();
 sg13g2_fill_1 FILLER_72_820 ();
 sg13g2_fill_2 FILLER_72_841 ();
 sg13g2_decap_8 FILLER_72_861 ();
 sg13g2_decap_8 FILLER_72_868 ();
 sg13g2_fill_2 FILLER_72_875 ();
 sg13g2_fill_1 FILLER_72_877 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_12 ();
 sg13g2_fill_1 FILLER_73_14 ();
 sg13g2_fill_2 FILLER_73_45 ();
 sg13g2_decap_4 FILLER_73_57 ();
 sg13g2_fill_2 FILLER_73_61 ();
 sg13g2_fill_2 FILLER_73_89 ();
 sg13g2_decap_8 FILLER_73_95 ();
 sg13g2_decap_8 FILLER_73_102 ();
 sg13g2_fill_2 FILLER_73_114 ();
 sg13g2_fill_2 FILLER_73_188 ();
 sg13g2_fill_1 FILLER_73_195 ();
 sg13g2_decap_4 FILLER_73_209 ();
 sg13g2_decap_8 FILLER_73_227 ();
 sg13g2_decap_4 FILLER_73_234 ();
 sg13g2_fill_1 FILLER_73_238 ();
 sg13g2_fill_1 FILLER_73_257 ();
 sg13g2_decap_4 FILLER_73_265 ();
 sg13g2_fill_2 FILLER_73_269 ();
 sg13g2_decap_8 FILLER_73_281 ();
 sg13g2_decap_8 FILLER_73_292 ();
 sg13g2_decap_8 FILLER_73_299 ();
 sg13g2_decap_8 FILLER_73_306 ();
 sg13g2_fill_1 FILLER_73_313 ();
 sg13g2_fill_2 FILLER_73_326 ();
 sg13g2_fill_1 FILLER_73_359 ();
 sg13g2_fill_2 FILLER_73_405 ();
 sg13g2_fill_1 FILLER_73_407 ();
 sg13g2_fill_2 FILLER_73_512 ();
 sg13g2_fill_1 FILLER_73_514 ();
 sg13g2_fill_2 FILLER_73_520 ();
 sg13g2_fill_1 FILLER_73_522 ();
 sg13g2_decap_8 FILLER_73_554 ();
 sg13g2_decap_8 FILLER_73_561 ();
 sg13g2_decap_4 FILLER_73_568 ();
 sg13g2_fill_2 FILLER_73_572 ();
 sg13g2_fill_2 FILLER_73_578 ();
 sg13g2_fill_1 FILLER_73_580 ();
 sg13g2_decap_8 FILLER_73_607 ();
 sg13g2_decap_8 FILLER_73_614 ();
 sg13g2_decap_8 FILLER_73_621 ();
 sg13g2_decap_8 FILLER_73_628 ();
 sg13g2_decap_8 FILLER_73_635 ();
 sg13g2_fill_2 FILLER_73_642 ();
 sg13g2_fill_1 FILLER_73_644 ();
 sg13g2_decap_4 FILLER_73_650 ();
 sg13g2_fill_1 FILLER_73_654 ();
 sg13g2_fill_2 FILLER_73_660 ();
 sg13g2_fill_2 FILLER_73_675 ();
 sg13g2_fill_2 FILLER_73_704 ();
 sg13g2_fill_2 FILLER_73_710 ();
 sg13g2_decap_4 FILLER_73_751 ();
 sg13g2_fill_2 FILLER_73_755 ();
 sg13g2_decap_4 FILLER_73_770 ();
 sg13g2_fill_2 FILLER_73_791 ();
 sg13g2_fill_1 FILLER_73_811 ();
 sg13g2_fill_1 FILLER_73_817 ();
 sg13g2_decap_8 FILLER_73_847 ();
 sg13g2_decap_8 FILLER_73_854 ();
 sg13g2_decap_8 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_73_868 ();
 sg13g2_fill_2 FILLER_73_875 ();
 sg13g2_fill_1 FILLER_73_877 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_7 ();
 sg13g2_fill_1 FILLER_74_11 ();
 sg13g2_decap_4 FILLER_74_42 ();
 sg13g2_decap_4 FILLER_74_77 ();
 sg13g2_fill_2 FILLER_74_91 ();
 sg13g2_fill_1 FILLER_74_93 ();
 sg13g2_fill_1 FILLER_74_120 ();
 sg13g2_fill_1 FILLER_74_171 ();
 sg13g2_fill_1 FILLER_74_176 ();
 sg13g2_fill_1 FILLER_74_182 ();
 sg13g2_fill_2 FILLER_74_214 ();
 sg13g2_fill_2 FILLER_74_220 ();
 sg13g2_decap_4 FILLER_74_253 ();
 sg13g2_decap_4 FILLER_74_261 ();
 sg13g2_fill_1 FILLER_74_265 ();
 sg13g2_decap_8 FILLER_74_327 ();
 sg13g2_decap_8 FILLER_74_334 ();
 sg13g2_decap_8 FILLER_74_341 ();
 sg13g2_fill_1 FILLER_74_348 ();
 sg13g2_fill_2 FILLER_74_358 ();
 sg13g2_fill_1 FILLER_74_360 ();
 sg13g2_decap_4 FILLER_74_365 ();
 sg13g2_fill_2 FILLER_74_369 ();
 sg13g2_decap_4 FILLER_74_380 ();
 sg13g2_fill_1 FILLER_74_406 ();
 sg13g2_fill_1 FILLER_74_413 ();
 sg13g2_fill_1 FILLER_74_422 ();
 sg13g2_decap_8 FILLER_74_432 ();
 sg13g2_fill_1 FILLER_74_439 ();
 sg13g2_fill_1 FILLER_74_451 ();
 sg13g2_fill_1 FILLER_74_455 ();
 sg13g2_decap_8 FILLER_74_469 ();
 sg13g2_decap_8 FILLER_74_489 ();
 sg13g2_fill_1 FILLER_74_496 ();
 sg13g2_decap_8 FILLER_74_501 ();
 sg13g2_fill_1 FILLER_74_508 ();
 sg13g2_fill_2 FILLER_74_515 ();
 sg13g2_fill_1 FILLER_74_524 ();
 sg13g2_fill_1 FILLER_74_544 ();
 sg13g2_fill_2 FILLER_74_576 ();
 sg13g2_fill_2 FILLER_74_593 ();
 sg13g2_fill_1 FILLER_74_595 ();
 sg13g2_fill_1 FILLER_74_601 ();
 sg13g2_decap_4 FILLER_74_611 ();
 sg13g2_fill_2 FILLER_74_615 ();
 sg13g2_fill_2 FILLER_74_643 ();
 sg13g2_decap_8 FILLER_74_671 ();
 sg13g2_fill_2 FILLER_74_691 ();
 sg13g2_fill_2 FILLER_74_727 ();
 sg13g2_fill_2 FILLER_74_744 ();
 sg13g2_fill_1 FILLER_74_746 ();
 sg13g2_fill_2 FILLER_74_752 ();
 sg13g2_fill_1 FILLER_74_754 ();
 sg13g2_fill_2 FILLER_74_762 ();
 sg13g2_fill_2 FILLER_74_796 ();
 sg13g2_fill_2 FILLER_74_816 ();
 sg13g2_fill_1 FILLER_74_833 ();
 sg13g2_fill_1 FILLER_74_857 ();
 sg13g2_decap_8 FILLER_74_871 ();
 sg13g2_decap_4 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_4 ();
 sg13g2_fill_1 FILLER_75_35 ();
 sg13g2_fill_2 FILLER_75_46 ();
 sg13g2_fill_1 FILLER_75_48 ();
 sg13g2_decap_8 FILLER_75_69 ();
 sg13g2_fill_1 FILLER_75_76 ();
 sg13g2_decap_8 FILLER_75_81 ();
 sg13g2_fill_1 FILLER_75_88 ();
 sg13g2_fill_2 FILLER_75_93 ();
 sg13g2_fill_1 FILLER_75_95 ();
 sg13g2_fill_1 FILLER_75_101 ();
 sg13g2_decap_8 FILLER_75_139 ();
 sg13g2_fill_2 FILLER_75_146 ();
 sg13g2_fill_1 FILLER_75_148 ();
 sg13g2_decap_4 FILLER_75_152 ();
 sg13g2_fill_1 FILLER_75_178 ();
 sg13g2_decap_8 FILLER_75_191 ();
 sg13g2_fill_1 FILLER_75_203 ();
 sg13g2_fill_2 FILLER_75_241 ();
 sg13g2_fill_1 FILLER_75_251 ();
 sg13g2_fill_1 FILLER_75_257 ();
 sg13g2_fill_1 FILLER_75_265 ();
 sg13g2_decap_8 FILLER_75_292 ();
 sg13g2_decap_8 FILLER_75_299 ();
 sg13g2_decap_8 FILLER_75_306 ();
 sg13g2_decap_4 FILLER_75_323 ();
 sg13g2_fill_1 FILLER_75_327 ();
 sg13g2_decap_4 FILLER_75_332 ();
 sg13g2_fill_1 FILLER_75_399 ();
 sg13g2_decap_8 FILLER_75_406 ();
 sg13g2_fill_2 FILLER_75_417 ();
 sg13g2_fill_1 FILLER_75_429 ();
 sg13g2_decap_4 FILLER_75_438 ();
 sg13g2_decap_8 FILLER_75_468 ();
 sg13g2_decap_8 FILLER_75_475 ();
 sg13g2_decap_8 FILLER_75_482 ();
 sg13g2_fill_1 FILLER_75_489 ();
 sg13g2_decap_4 FILLER_75_494 ();
 sg13g2_fill_2 FILLER_75_498 ();
 sg13g2_fill_1 FILLER_75_504 ();
 sg13g2_fill_2 FILLER_75_510 ();
 sg13g2_fill_1 FILLER_75_512 ();
 sg13g2_decap_4 FILLER_75_544 ();
 sg13g2_fill_1 FILLER_75_569 ();
 sg13g2_fill_1 FILLER_75_573 ();
 sg13g2_fill_1 FILLER_75_580 ();
 sg13g2_fill_1 FILLER_75_588 ();
 sg13g2_fill_2 FILLER_75_605 ();
 sg13g2_decap_4 FILLER_75_643 ();
 sg13g2_fill_2 FILLER_75_647 ();
 sg13g2_decap_8 FILLER_75_659 ();
 sg13g2_decap_8 FILLER_75_666 ();
 sg13g2_decap_8 FILLER_75_673 ();
 sg13g2_fill_1 FILLER_75_680 ();
 sg13g2_decap_8 FILLER_75_691 ();
 sg13g2_decap_8 FILLER_75_698 ();
 sg13g2_fill_2 FILLER_75_715 ();
 sg13g2_fill_1 FILLER_75_722 ();
 sg13g2_fill_2 FILLER_75_728 ();
 sg13g2_fill_2 FILLER_75_739 ();
 sg13g2_fill_1 FILLER_75_741 ();
 sg13g2_fill_2 FILLER_75_772 ();
 sg13g2_fill_1 FILLER_75_774 ();
 sg13g2_fill_1 FILLER_75_780 ();
 sg13g2_fill_1 FILLER_75_789 ();
 sg13g2_fill_2 FILLER_75_816 ();
 sg13g2_decap_8 FILLER_75_833 ();
 sg13g2_decap_8 FILLER_75_840 ();
 sg13g2_decap_8 FILLER_75_847 ();
 sg13g2_decap_8 FILLER_75_854 ();
 sg13g2_decap_8 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_75_868 ();
 sg13g2_fill_2 FILLER_75_875 ();
 sg13g2_fill_1 FILLER_75_877 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_4 FILLER_76_21 ();
 sg13g2_fill_2 FILLER_76_25 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_4 FILLER_76_72 ();
 sg13g2_decap_8 FILLER_76_86 ();
 sg13g2_fill_1 FILLER_76_93 ();
 sg13g2_fill_2 FILLER_76_141 ();
 sg13g2_fill_1 FILLER_76_148 ();
 sg13g2_fill_1 FILLER_76_246 ();
 sg13g2_fill_1 FILLER_76_252 ();
 sg13g2_fill_1 FILLER_76_257 ();
 sg13g2_fill_1 FILLER_76_284 ();
 sg13g2_fill_1 FILLER_76_311 ();
 sg13g2_decap_4 FILLER_76_343 ();
 sg13g2_fill_1 FILLER_76_347 ();
 sg13g2_decap_4 FILLER_76_364 ();
 sg13g2_decap_4 FILLER_76_381 ();
 sg13g2_fill_2 FILLER_76_385 ();
 sg13g2_fill_2 FILLER_76_392 ();
 sg13g2_fill_1 FILLER_76_398 ();
 sg13g2_fill_1 FILLER_76_403 ();
 sg13g2_fill_1 FILLER_76_412 ();
 sg13g2_fill_2 FILLER_76_418 ();
 sg13g2_fill_1 FILLER_76_425 ();
 sg13g2_fill_2 FILLER_76_436 ();
 sg13g2_fill_2 FILLER_76_443 ();
 sg13g2_fill_2 FILLER_76_512 ();
 sg13g2_fill_1 FILLER_76_542 ();
 sg13g2_decap_8 FILLER_76_551 ();
 sg13g2_decap_4 FILLER_76_558 ();
 sg13g2_fill_1 FILLER_76_562 ();
 sg13g2_fill_1 FILLER_76_580 ();
 sg13g2_fill_2 FILLER_76_585 ();
 sg13g2_fill_1 FILLER_76_606 ();
 sg13g2_decap_8 FILLER_76_641 ();
 sg13g2_fill_1 FILLER_76_648 ();
 sg13g2_decap_4 FILLER_76_661 ();
 sg13g2_fill_2 FILLER_76_665 ();
 sg13g2_fill_2 FILLER_76_680 ();
 sg13g2_fill_1 FILLER_76_695 ();
 sg13g2_fill_2 FILLER_76_723 ();
 sg13g2_fill_2 FILLER_76_730 ();
 sg13g2_fill_2 FILLER_76_737 ();
 sg13g2_fill_1 FILLER_76_739 ();
 sg13g2_decap_8 FILLER_76_745 ();
 sg13g2_fill_2 FILLER_76_752 ();
 sg13g2_fill_1 FILLER_76_754 ();
 sg13g2_decap_8 FILLER_76_771 ();
 sg13g2_decap_4 FILLER_76_778 ();
 sg13g2_fill_2 FILLER_76_782 ();
 sg13g2_fill_1 FILLER_76_797 ();
 sg13g2_decap_8 FILLER_76_802 ();
 sg13g2_decap_8 FILLER_76_809 ();
 sg13g2_decap_8 FILLER_76_816 ();
 sg13g2_decap_8 FILLER_76_823 ();
 sg13g2_decap_8 FILLER_76_830 ();
 sg13g2_decap_8 FILLER_76_837 ();
 sg13g2_decap_8 FILLER_76_844 ();
 sg13g2_decap_8 FILLER_76_851 ();
 sg13g2_decap_8 FILLER_76_858 ();
 sg13g2_decap_8 FILLER_76_865 ();
 sg13g2_decap_4 FILLER_76_872 ();
 sg13g2_fill_2 FILLER_76_876 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_fill_2 FILLER_77_21 ();
 sg13g2_fill_2 FILLER_77_49 ();
 sg13g2_fill_1 FILLER_77_51 ();
 sg13g2_fill_2 FILLER_77_60 ();
 sg13g2_fill_1 FILLER_77_62 ();
 sg13g2_fill_1 FILLER_77_73 ();
 sg13g2_decap_8 FILLER_77_78 ();
 sg13g2_fill_2 FILLER_77_156 ();
 sg13g2_fill_2 FILLER_77_198 ();
 sg13g2_fill_2 FILLER_77_207 ();
 sg13g2_fill_2 FILLER_77_214 ();
 sg13g2_fill_1 FILLER_77_216 ();
 sg13g2_fill_2 FILLER_77_231 ();
 sg13g2_fill_1 FILLER_77_238 ();
 sg13g2_fill_2 FILLER_77_248 ();
 sg13g2_fill_1 FILLER_77_250 ();
 sg13g2_fill_2 FILLER_77_269 ();
 sg13g2_decap_8 FILLER_77_297 ();
 sg13g2_decap_8 FILLER_77_304 ();
 sg13g2_decap_4 FILLER_77_311 ();
 sg13g2_decap_8 FILLER_77_341 ();
 sg13g2_decap_4 FILLER_77_348 ();
 sg13g2_fill_2 FILLER_77_352 ();
 sg13g2_fill_2 FILLER_77_359 ();
 sg13g2_fill_1 FILLER_77_361 ();
 sg13g2_decap_4 FILLER_77_422 ();
 sg13g2_decap_4 FILLER_77_436 ();
 sg13g2_fill_2 FILLER_77_440 ();
 sg13g2_fill_2 FILLER_77_467 ();
 sg13g2_decap_8 FILLER_77_476 ();
 sg13g2_fill_2 FILLER_77_497 ();
 sg13g2_fill_2 FILLER_77_512 ();
 sg13g2_fill_2 FILLER_77_532 ();
 sg13g2_fill_1 FILLER_77_534 ();
 sg13g2_fill_1 FILLER_77_574 ();
 sg13g2_fill_1 FILLER_77_585 ();
 sg13g2_fill_2 FILLER_77_590 ();
 sg13g2_fill_1 FILLER_77_597 ();
 sg13g2_decap_4 FILLER_77_605 ();
 sg13g2_fill_1 FILLER_77_700 ();
 sg13g2_decap_8 FILLER_77_708 ();
 sg13g2_fill_1 FILLER_77_715 ();
 sg13g2_fill_2 FILLER_77_747 ();
 sg13g2_decap_4 FILLER_77_754 ();
 sg13g2_fill_1 FILLER_77_758 ();
 sg13g2_decap_8 FILLER_77_798 ();
 sg13g2_decap_8 FILLER_77_805 ();
 sg13g2_decap_8 FILLER_77_812 ();
 sg13g2_decap_8 FILLER_77_819 ();
 sg13g2_decap_8 FILLER_77_826 ();
 sg13g2_decap_8 FILLER_77_833 ();
 sg13g2_decap_8 FILLER_77_840 ();
 sg13g2_decap_8 FILLER_77_847 ();
 sg13g2_decap_8 FILLER_77_854 ();
 sg13g2_decap_8 FILLER_77_861 ();
 sg13g2_decap_8 FILLER_77_868 ();
 sg13g2_fill_2 FILLER_77_875 ();
 sg13g2_fill_1 FILLER_77_877 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_32 ();
 sg13g2_fill_2 FILLER_78_119 ();
 sg13g2_fill_1 FILLER_78_154 ();
 sg13g2_fill_1 FILLER_78_234 ();
 sg13g2_fill_2 FILLER_78_252 ();
 sg13g2_fill_2 FILLER_78_282 ();
 sg13g2_fill_2 FILLER_78_288 ();
 sg13g2_fill_1 FILLER_78_401 ();
 sg13g2_fill_1 FILLER_78_407 ();
 sg13g2_fill_1 FILLER_78_434 ();
 sg13g2_fill_2 FILLER_78_465 ();
 sg13g2_fill_1 FILLER_78_467 ();
 sg13g2_fill_2 FILLER_78_494 ();
 sg13g2_fill_2 FILLER_78_524 ();
 sg13g2_fill_1 FILLER_78_536 ();
 sg13g2_fill_2 FILLER_78_542 ();
 sg13g2_fill_1 FILLER_78_549 ();
 sg13g2_fill_2 FILLER_78_557 ();
 sg13g2_fill_2 FILLER_78_562 ();
 sg13g2_fill_2 FILLER_78_569 ();
 sg13g2_decap_8 FILLER_78_616 ();
 sg13g2_decap_8 FILLER_78_623 ();
 sg13g2_decap_8 FILLER_78_630 ();
 sg13g2_decap_8 FILLER_78_637 ();
 sg13g2_fill_1 FILLER_78_670 ();
 sg13g2_fill_2 FILLER_78_684 ();
 sg13g2_fill_2 FILLER_78_689 ();
 sg13g2_decap_8 FILLER_78_743 ();
 sg13g2_decap_8 FILLER_78_750 ();
 sg13g2_decap_8 FILLER_78_757 ();
 sg13g2_decap_8 FILLER_78_764 ();
 sg13g2_decap_8 FILLER_78_771 ();
 sg13g2_decap_8 FILLER_78_778 ();
 sg13g2_decap_8 FILLER_78_785 ();
 sg13g2_decap_8 FILLER_78_792 ();
 sg13g2_decap_8 FILLER_78_799 ();
 sg13g2_decap_8 FILLER_78_806 ();
 sg13g2_decap_8 FILLER_78_813 ();
 sg13g2_decap_8 FILLER_78_820 ();
 sg13g2_decap_8 FILLER_78_827 ();
 sg13g2_decap_8 FILLER_78_834 ();
 sg13g2_decap_8 FILLER_78_841 ();
 sg13g2_decap_8 FILLER_78_848 ();
 sg13g2_decap_8 FILLER_78_855 ();
 sg13g2_decap_8 FILLER_78_862 ();
 sg13g2_decap_8 FILLER_78_869 ();
 sg13g2_fill_2 FILLER_78_876 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_4 FILLER_79_21 ();
 sg13g2_fill_1 FILLER_79_25 ();
 sg13g2_fill_1 FILLER_79_52 ();
 sg13g2_fill_1 FILLER_79_123 ();
 sg13g2_fill_2 FILLER_79_228 ();
 sg13g2_fill_1 FILLER_79_240 ();
 sg13g2_fill_1 FILLER_79_330 ();
 sg13g2_fill_1 FILLER_79_345 ();
 sg13g2_fill_2 FILLER_79_398 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_fill_1 FILLER_79_454 ();
 sg13g2_fill_2 FILLER_79_458 ();
 sg13g2_fill_2 FILLER_79_476 ();
 sg13g2_fill_1 FILLER_79_478 ();
 sg13g2_fill_1 FILLER_79_542 ();
 sg13g2_fill_1 FILLER_79_605 ();
 sg13g2_decap_8 FILLER_79_610 ();
 sg13g2_decap_4 FILLER_79_617 ();
 sg13g2_decap_8 FILLER_79_626 ();
 sg13g2_decap_8 FILLER_79_633 ();
 sg13g2_fill_2 FILLER_79_640 ();
 sg13g2_fill_1 FILLER_79_642 ();
 sg13g2_decap_8 FILLER_79_651 ();
 sg13g2_decap_8 FILLER_79_658 ();
 sg13g2_decap_8 FILLER_79_665 ();
 sg13g2_decap_8 FILLER_79_711 ();
 sg13g2_decap_8 FILLER_79_718 ();
 sg13g2_decap_8 FILLER_79_725 ();
 sg13g2_decap_8 FILLER_79_732 ();
 sg13g2_decap_8 FILLER_79_739 ();
 sg13g2_decap_8 FILLER_79_746 ();
 sg13g2_fill_2 FILLER_79_753 ();
 sg13g2_decap_8 FILLER_79_758 ();
 sg13g2_decap_8 FILLER_79_765 ();
 sg13g2_decap_8 FILLER_79_772 ();
 sg13g2_decap_8 FILLER_79_779 ();
 sg13g2_decap_8 FILLER_79_786 ();
 sg13g2_decap_8 FILLER_79_793 ();
 sg13g2_decap_8 FILLER_79_800 ();
 sg13g2_decap_8 FILLER_79_807 ();
 sg13g2_decap_8 FILLER_79_814 ();
 sg13g2_decap_8 FILLER_79_821 ();
 sg13g2_decap_8 FILLER_79_828 ();
 sg13g2_decap_8 FILLER_79_835 ();
 sg13g2_decap_8 FILLER_79_842 ();
 sg13g2_decap_8 FILLER_79_849 ();
 sg13g2_decap_8 FILLER_79_856 ();
 sg13g2_decap_8 FILLER_79_863 ();
 sg13g2_decap_8 FILLER_79_870 ();
 sg13g2_fill_1 FILLER_79_877 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_4 FILLER_80_35 ();
 sg13g2_fill_1 FILLER_80_39 ();
 sg13g2_fill_1 FILLER_80_99 ();
 sg13g2_fill_2 FILLER_80_141 ();
 sg13g2_fill_2 FILLER_80_157 ();
 sg13g2_fill_1 FILLER_80_218 ();
 sg13g2_fill_2 FILLER_80_228 ();
 sg13g2_fill_2 FILLER_80_243 ();
 sg13g2_fill_1 FILLER_80_258 ();
 sg13g2_decap_4 FILLER_80_293 ();
 sg13g2_fill_1 FILLER_80_297 ();
 sg13g2_fill_2 FILLER_80_389 ();
 sg13g2_fill_1 FILLER_80_391 ();
 sg13g2_fill_1 FILLER_80_431 ();
 sg13g2_decap_8 FILLER_80_458 ();
 sg13g2_decap_8 FILLER_80_465 ();
 sg13g2_fill_2 FILLER_80_472 ();
 sg13g2_fill_2 FILLER_80_536 ();
 sg13g2_fill_1 FILLER_80_538 ();
 sg13g2_fill_2 FILLER_80_578 ();
 sg13g2_fill_1 FILLER_80_580 ();
 sg13g2_decap_8 FILLER_80_607 ();
 sg13g2_decap_8 FILLER_80_614 ();
 sg13g2_decap_8 FILLER_80_621 ();
 sg13g2_decap_8 FILLER_80_628 ();
 sg13g2_decap_8 FILLER_80_635 ();
 sg13g2_decap_8 FILLER_80_642 ();
 sg13g2_decap_8 FILLER_80_649 ();
 sg13g2_decap_8 FILLER_80_656 ();
 sg13g2_decap_8 FILLER_80_663 ();
 sg13g2_decap_8 FILLER_80_670 ();
 sg13g2_decap_8 FILLER_80_677 ();
 sg13g2_decap_4 FILLER_80_684 ();
 sg13g2_fill_2 FILLER_80_688 ();
 sg13g2_decap_8 FILLER_80_711 ();
 sg13g2_decap_8 FILLER_80_718 ();
 sg13g2_decap_8 FILLER_80_725 ();
 sg13g2_decap_8 FILLER_80_732 ();
 sg13g2_decap_8 FILLER_80_739 ();
 sg13g2_decap_8 FILLER_80_746 ();
 sg13g2_decap_8 FILLER_80_753 ();
 sg13g2_decap_8 FILLER_80_760 ();
 sg13g2_decap_8 FILLER_80_767 ();
 sg13g2_decap_8 FILLER_80_774 ();
 sg13g2_decap_8 FILLER_80_781 ();
 sg13g2_decap_8 FILLER_80_788 ();
 sg13g2_decap_8 FILLER_80_795 ();
 sg13g2_decap_8 FILLER_80_802 ();
 sg13g2_decap_8 FILLER_80_809 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_decap_8 FILLER_80_823 ();
 sg13g2_decap_8 FILLER_80_830 ();
 sg13g2_decap_8 FILLER_80_837 ();
 sg13g2_decap_8 FILLER_80_844 ();
 sg13g2_decap_8 FILLER_80_851 ();
 sg13g2_decap_8 FILLER_80_858 ();
 sg13g2_decap_8 FILLER_80_865 ();
 sg13g2_decap_4 FILLER_80_872 ();
 sg13g2_fill_2 FILLER_80_876 ();
endmodule
