module tt_um_kbeckmann_flame (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \LFSR[0] ;
 wire \LFSR[1] ;
 wire \LFSR[2] ;
 wire \LFSR[3] ;
 wire \LFSR[4] ;
 wire \LFSR[5] ;
 wire \VAL[0] ;
 wire \VAL[10] ;
 wire \VAL[11] ;
 wire \VAL[12] ;
 wire \VAL[13] ;
 wire \VAL[14] ;
 wire \VAL[15] ;
 wire \VAL[16] ;
 wire \VAL[17] ;
 wire \VAL[18] ;
 wire \VAL[19] ;
 wire \VAL[1] ;
 wire \VAL[20] ;
 wire \VAL[21] ;
 wire \VAL[22] ;
 wire \VAL[23] ;
 wire \VAL[2] ;
 wire \VAL[3] ;
 wire \VAL[4] ;
 wire \VAL[5] ;
 wire \VAL[6] ;
 wire \VAL[7] ;
 wire \VAL[8] ;
 wire \VAL[9] ;
 wire \Voice1.accumulator[0] ;
 wire \Voice1.accumulator[10] ;
 wire \Voice1.accumulator[11] ;
 wire \Voice1.accumulator[12] ;
 wire \Voice1.accumulator[13] ;
 wire \Voice1.accumulator[14] ;
 wire \Voice1.accumulator[15] ;
 wire \Voice1.accumulator[16] ;
 wire \Voice1.accumulator[17] ;
 wire \Voice1.accumulator[18] ;
 wire \Voice1.accumulator[19] ;
 wire \Voice1.accumulator[1] ;
 wire \Voice1.accumulator[20] ;
 wire \Voice1.accumulator[21] ;
 wire \Voice1.accumulator[22] ;
 wire \Voice1.accumulator[23] ;
 wire \Voice1.accumulator[2] ;
 wire \Voice1.accumulator[3] ;
 wire \Voice1.accumulator[4] ;
 wire \Voice1.accumulator[5] ;
 wire \Voice1.accumulator[6] ;
 wire \Voice1.accumulator[7] ;
 wire \Voice1.accumulator[8] ;
 wire \Voice1.accumulator[9] ;
 wire \Voice1.en ;
 wire \Voice1.pulse ;
 wire \Voice1.pulsewidth[0] ;
 wire \Voice1.pulsewidth[10] ;
 wire \Voice1.pulsewidth[1] ;
 wire \Voice1.pulsewidth[2] ;
 wire \Voice1.pulsewidth[3] ;
 wire \Voice1.pulsewidth[4] ;
 wire \Voice1.pulsewidth[5] ;
 wire \Voice1.pulsewidth[6] ;
 wire \Voice1.pulsewidth[7] ;
 wire \Voice1.pulsewidth[8] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire clknet_0_clk;
 wire net90;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \ctr_audio[0] ;
 wire \ctr_audio[19] ;
 wire \ctr_audio[1] ;
 wire \ctr_audio[20] ;
 wire \ctr_audio[21] ;
 wire \ctr_audio[22] ;
 wire \ctr_audio[2] ;
 wire \ctr_audio[3] ;
 wire \ctr_audio[4] ;
 wire \ctr_audio[5] ;
 wire \ctr_audio[6] ;
 wire \ctr_audio[7] ;
 wire \ctr_audio[8] ;
 wire \ctr_audio[9] ;
 wire \ctr_clkdiv25[0] ;
 wire \ctr_clkdiv25[1] ;
 wire \ctr_clkdiv25[2] ;
 wire \ctr_clkdiv25[3] ;
 wire \ctr_clkdiv25[4] ;
 wire \ctr_clkdiv25[5] ;
 wire \ctr_clkdiv25[6] ;
 wire \ctr_clkdiv25[7] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \xq[0] ;
 wire \xq[10] ;
 wire \xq[11] ;
 wire \xq[1] ;
 wire \xq[2] ;
 wire \xq[3] ;
 wire \xq[4] ;
 wire \xq[5] ;
 wire \xq[6] ;
 wire \xq[7] ;
 wire \xq[8] ;
 wire \xq[9] ;
 wire \xqo[0] ;
 wire \xqo[10] ;
 wire \xqo[11] ;
 wire \xqo[1] ;
 wire \xqo[2] ;
 wire \xqo[3] ;
 wire \xqo[4] ;
 wire \xqo[5] ;
 wire \xqo[6] ;
 wire \xqo[7] ;
 wire \xqo[8] ;
 wire \xqo[9] ;
 wire \yq[0] ;
 wire \yq[10] ;
 wire \yq[11] ;
 wire \yq[12] ;
 wire \yq[1] ;
 wire \yq[2] ;
 wire \yq[3] ;
 wire \yq[4] ;
 wire \yq[5] ;
 wire \yq[6] ;
 wire \yq[7] ;
 wire \yq[8] ;
 wire \yq[9] ;
 wire \yqo[0] ;
 wire \yqo[10] ;
 wire \yqo[11] ;
 wire \yqo[12] ;
 wire \yqo[1] ;
 wire \yqo[2] ;
 wire \yqo[3] ;
 wire \yqo[4] ;
 wire \yqo[5] ;
 wire \yqo[6] ;
 wire \yqo[7] ;
 wire \yqo[8] ;
 wire \yqo[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_dfrbp_1 \LFSR[0]$_SDFF_PP1_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net90),
    .D(_0019_),
    .Q_N(_1639_),
    .Q(\LFSR[0] ));
 sg13g2_dfrbp_1 \LFSR[1]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net91),
    .D(_0020_),
    .Q_N(_1638_),
    .Q(\LFSR[1] ));
 sg13g2_dfrbp_1 \LFSR[2]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net92),
    .D(_0021_),
    .Q_N(_1637_),
    .Q(\LFSR[2] ));
 sg13g2_dfrbp_1 \LFSR[3]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net93),
    .D(_0022_),
    .Q_N(_1636_),
    .Q(\LFSR[3] ));
 sg13g2_dfrbp_1 \LFSR[4]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net94),
    .D(_0023_),
    .Q_N(_1635_),
    .Q(\LFSR[4] ));
 sg13g2_dfrbp_1 \LFSR[5]$_SDFF_PP0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net95),
    .D(_0024_),
    .Q_N(_1634_),
    .Q(\LFSR[5] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[0]$_DFFE_PP_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net96),
    .D(_0025_),
    .Q_N(_1633_),
    .Q(\Voice1.accumulator[0] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[10]$_DFFE_PP_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net97),
    .D(_0026_),
    .Q_N(_1632_),
    .Q(\Voice1.accumulator[10] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[11]$_DFFE_PP_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net98),
    .D(_0027_),
    .Q_N(_1631_),
    .Q(\Voice1.accumulator[11] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[12]$_DFFE_PP_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net99),
    .D(_0028_),
    .Q_N(_1630_),
    .Q(\Voice1.accumulator[12] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[13]$_DFFE_PP_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net100),
    .D(_0029_),
    .Q_N(_0002_),
    .Q(\Voice1.accumulator[13] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[14]$_DFFE_PP_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net101),
    .D(_0030_),
    .Q_N(_1629_),
    .Q(\Voice1.accumulator[14] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[15]$_DFFE_PP_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net102),
    .D(_0031_),
    .Q_N(_1628_),
    .Q(\Voice1.accumulator[15] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[16]$_DFFE_PP_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net103),
    .D(_0032_),
    .Q_N(_1627_),
    .Q(\Voice1.accumulator[16] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[17]$_DFFE_PP_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net104),
    .D(_0033_),
    .Q_N(_1626_),
    .Q(\Voice1.accumulator[17] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[18]$_DFFE_PP_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net105),
    .D(_0034_),
    .Q_N(_1625_),
    .Q(\Voice1.accumulator[18] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[19]$_DFFE_PP_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net106),
    .D(_0035_),
    .Q_N(_1624_),
    .Q(\Voice1.accumulator[19] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[1]$_DFFE_PP_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net107),
    .D(_0036_),
    .Q_N(_1623_),
    .Q(\Voice1.accumulator[1] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[20]$_DFFE_PP_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net108),
    .D(_0037_),
    .Q_N(_1622_),
    .Q(\Voice1.accumulator[20] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[21]$_DFFE_PP_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net109),
    .D(_0038_),
    .Q_N(_0005_),
    .Q(\Voice1.accumulator[21] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[22]$_DFFE_PP_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net110),
    .D(_0039_),
    .Q_N(_1621_),
    .Q(\Voice1.accumulator[22] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[23]$_DFFE_PP_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net111),
    .D(_0040_),
    .Q_N(_0004_),
    .Q(\Voice1.accumulator[23] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[2]$_DFFE_PP_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net112),
    .D(_0041_),
    .Q_N(_1620_),
    .Q(\Voice1.accumulator[2] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[3]$_DFFE_PP_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net113),
    .D(_0042_),
    .Q_N(_1619_),
    .Q(\Voice1.accumulator[3] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[4]$_DFFE_PP_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net114),
    .D(_0043_),
    .Q_N(_1618_),
    .Q(\Voice1.accumulator[4] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[5]$_DFFE_PP_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net115),
    .D(_0044_),
    .Q_N(_1617_),
    .Q(\Voice1.accumulator[5] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[6]$_DFFE_PP_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net116),
    .D(_0045_),
    .Q_N(_1616_),
    .Q(\Voice1.accumulator[6] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[7]$_DFFE_PP_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net117),
    .D(_0046_),
    .Q_N(_1615_),
    .Q(\Voice1.accumulator[7] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[8]$_DFFE_PP_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net118),
    .D(_0047_),
    .Q_N(_1614_),
    .Q(\Voice1.accumulator[8] ));
 sg13g2_dfrbp_1 \Voice1.accumulator[9]$_DFFE_PP_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net119),
    .D(_0048_),
    .Q_N(_1613_),
    .Q(\Voice1.accumulator[9] ));
 sg13g2_dfrbp_1 \Voice1.pulse$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net120),
    .D(_0049_),
    .Q_N(_1612_),
    .Q(\Voice1.pulse ));
 sg13g2_buf_1 _1643_ (.A(\hvsync_gen.vpos[1] ),
    .X(_0923_));
 sg13g2_buf_8 _1644_ (.A(\hvsync_gen.vpos[2] ),
    .X(_0924_));
 sg13g2_buf_1 _1645_ (.A(\hvsync_gen.vpos[9] ),
    .X(_0925_));
 sg13g2_buf_1 _1646_ (.A(\hvsync_gen.vpos[5] ),
    .X(_0926_));
 sg13g2_buf_1 _1647_ (.A(net72),
    .X(_0927_));
 sg13g2_buf_1 _1648_ (.A(\hvsync_gen.vpos[7] ),
    .X(_0928_));
 sg13g2_buf_1 _1649_ (.A(_0928_),
    .X(_0929_));
 sg13g2_buf_1 _1650_ (.A(net61),
    .X(_0930_));
 sg13g2_buf_1 _1651_ (.A(\hvsync_gen.vpos[6] ),
    .X(_0931_));
 sg13g2_buf_1 _1652_ (.A(_0931_),
    .X(_0932_));
 sg13g2_buf_1 _1653_ (.A(net60),
    .X(_0933_));
 sg13g2_buf_1 _1654_ (.A(\hvsync_gen.vpos[8] ),
    .X(_0934_));
 sg13g2_buf_1 _1655_ (.A(_0934_),
    .X(_0935_));
 sg13g2_nand4_1 _1656_ (.B(net36),
    .C(net35),
    .A(net62),
    .Y(_0936_),
    .D(net59));
 sg13g2_buf_1 _1657_ (.A(_0936_),
    .X(_0937_));
 sg13g2_buf_8 _1658_ (.A(\hvsync_gen.vpos[3] ),
    .X(_0938_));
 sg13g2_buf_1 _1659_ (.A(_0938_),
    .X(_0939_));
 sg13g2_buf_8 _1660_ (.A(\hvsync_gen.vpos[4] ),
    .X(_0940_));
 sg13g2_buf_1 _1661_ (.A(net71),
    .X(_0941_));
 sg13g2_inv_1 _1662_ (.Y(_0942_),
    .A(net57));
 sg13g2_nand2_1 _1663_ (.Y(_0943_),
    .A(net58),
    .B(_0942_));
 sg13g2_nor4_1 _1664_ (.A(_0924_),
    .B(net73),
    .C(_0937_),
    .D(_0943_),
    .Y(_0944_));
 sg13g2_and2_1 _1665_ (.A(_0923_),
    .B(_0944_),
    .X(_0001_));
 sg13g2_buf_1 _1666_ (.A(\hvsync_gen.hpos[7] ),
    .X(_0945_));
 sg13g2_buf_2 _1667_ (.A(\hvsync_gen.hpos[8] ),
    .X(_0946_));
 sg13g2_buf_1 _1668_ (.A(_0946_),
    .X(_0947_));
 sg13g2_buf_1 _1669_ (.A(\hvsync_gen.hpos[9] ),
    .X(_0948_));
 sg13g2_buf_1 _1670_ (.A(_0948_),
    .X(_0949_));
 sg13g2_o21ai_1 _1671_ (.B1(_0949_),
    .Y(_0950_),
    .A1(net70),
    .A2(net56));
 sg13g2_buf_1 _1672_ (.A(\hvsync_gen.hpos[6] ),
    .X(_0951_));
 sg13g2_buf_1 _1673_ (.A(\hvsync_gen.hpos[5] ),
    .X(_0952_));
 sg13g2_buf_1 _1674_ (.A(_0952_),
    .X(_0953_));
 sg13g2_buf_1 _1675_ (.A(\hvsync_gen.hpos[4] ),
    .X(_0954_));
 sg13g2_nor4_1 _1676_ (.A(net56),
    .B(net68),
    .C(net54),
    .D(net67),
    .Y(_0955_));
 sg13g2_inv_2 _1677_ (.Y(_0956_),
    .A(_0946_));
 sg13g2_nand3_1 _1678_ (.B(net54),
    .C(net67),
    .A(net68),
    .Y(_0957_));
 sg13g2_a21oi_1 _1679_ (.A1(_0956_),
    .A2(_0957_),
    .Y(_0958_),
    .B1(_0006_));
 sg13g2_nor3_1 _1680_ (.A(_0950_),
    .B(_0955_),
    .C(_0958_),
    .Y(_0000_));
 sg13g2_buf_1 _1681_ (.A(rst_n),
    .X(_0959_));
 sg13g2_inv_1 _1682_ (.Y(_0960_),
    .A(_0959_));
 sg13g2_inv_1 _1683_ (.Y(_0961_),
    .A(\Voice1.en ));
 sg13g2_nor2_2 _1684_ (.A(_0960_),
    .B(_0961_),
    .Y(_0962_));
 sg13g2_buf_1 _1685_ (.A(\Voice1.pulsewidth[7] ),
    .X(_0963_));
 sg13g2_buf_2 _1686_ (.A(\ctr_audio[22] ),
    .X(_0964_));
 sg13g2_buf_2 _1687_ (.A(\ctr_audio[21] ),
    .X(_0965_));
 sg13g2_nand2b_1 _1688_ (.Y(_0966_),
    .B(_0965_),
    .A_N(_0964_));
 sg13g2_buf_1 _1689_ (.A(\ctr_audio[19] ),
    .X(_0967_));
 sg13g2_buf_1 _1690_ (.A(_0967_),
    .X(_0968_));
 sg13g2_a21o_1 _1691_ (.A2(_0966_),
    .A1(net66),
    .B1(net53),
    .X(_0969_));
 sg13g2_buf_1 _1692_ (.A(\Voice1.pulsewidth[10] ),
    .X(_0970_));
 sg13g2_buf_1 _1693_ (.A(_0970_),
    .X(_0971_));
 sg13g2_buf_8 _1694_ (.A(_0965_),
    .X(_0972_));
 sg13g2_and2_1 _1695_ (.A(net51),
    .B(_0964_),
    .X(_0973_));
 sg13g2_and2_1 _1696_ (.A(net66),
    .B(_0967_),
    .X(_0974_));
 sg13g2_buf_2 _1697_ (.A(_0974_),
    .X(_0975_));
 sg13g2_a22oi_1 _1698_ (.Y(_0976_),
    .B1(_0966_),
    .B2(_0975_),
    .A2(_0973_),
    .A1(net52));
 sg13g2_buf_2 _1699_ (.A(_0013_),
    .X(_0977_));
 sg13g2_a21oi_1 _1700_ (.A1(_0969_),
    .A2(_0976_),
    .Y(_0978_),
    .B1(_0977_));
 sg13g2_nand2_1 _1701_ (.Y(_0979_),
    .A(_0962_),
    .B(_0978_));
 sg13g2_xnor2_1 _1702_ (.Y(_0025_),
    .A(\Voice1.accumulator[0] ),
    .B(_0979_));
 sg13g2_inv_1 _1703_ (.Y(_0980_),
    .A(\Voice1.accumulator[7] ));
 sg13g2_inv_1 _1704_ (.Y(_0981_),
    .A(net53));
 sg13g2_buf_1 _1705_ (.A(_0963_),
    .X(_0982_));
 sg13g2_nand2b_1 _1706_ (.Y(_0983_),
    .B(_0964_),
    .A_N(_0970_));
 sg13g2_buf_8 _1707_ (.A(_0964_),
    .X(_0984_));
 sg13g2_nand2b_1 _1708_ (.Y(_0985_),
    .B(net66),
    .A_N(net49));
 sg13g2_o21ai_1 _1709_ (.B1(_0985_),
    .Y(_0986_),
    .A1(net50),
    .A2(_0983_));
 sg13g2_nand2_1 _1710_ (.Y(_0987_),
    .A(net53),
    .B(net49));
 sg13g2_nand2b_1 _1711_ (.Y(_0988_),
    .B(net66),
    .A_N(net53));
 sg13g2_nand2_1 _1712_ (.Y(_0989_),
    .A(_0987_),
    .B(_0988_));
 sg13g2_inv_1 _1713_ (.Y(_0990_),
    .A(net51));
 sg13g2_a221oi_1 _1714_ (.B2(net52),
    .C1(_0990_),
    .B1(_0989_),
    .A1(_0981_),
    .Y(_0991_),
    .A2(_0986_));
 sg13g2_nor2_1 _1715_ (.A(net51),
    .B(_0975_),
    .Y(_0992_));
 sg13g2_or3_1 _1716_ (.A(_0977_),
    .B(_0991_),
    .C(_0992_),
    .X(_0993_));
 sg13g2_buf_1 _1717_ (.A(_0993_),
    .X(_0994_));
 sg13g2_nand2_1 _1718_ (.Y(_0995_),
    .A(_0980_),
    .B(_0994_));
 sg13g2_inv_1 _1719_ (.Y(_0996_),
    .A(net50));
 sg13g2_nor2_1 _1720_ (.A(_0996_),
    .B(net49),
    .Y(_0997_));
 sg13g2_nand2b_1 _1721_ (.Y(_0998_),
    .B(net49),
    .A_N(net50));
 sg13g2_a21oi_1 _1722_ (.A1(_0998_),
    .A2(_0988_),
    .Y(_0999_),
    .B1(net52));
 sg13g2_o21ai_1 _1723_ (.B1(net51),
    .Y(_1000_),
    .A1(_0997_),
    .A2(_0999_));
 sg13g2_o21ai_1 _1724_ (.B1(_0975_),
    .Y(_1001_),
    .A1(net52),
    .A2(_0990_));
 sg13g2_a21oi_1 _1725_ (.A1(_1000_),
    .A2(_1001_),
    .Y(_1002_),
    .B1(_0977_));
 sg13g2_or2_1 _1726_ (.X(_1003_),
    .B(_1002_),
    .A(\Voice1.accumulator[6] ));
 sg13g2_nor2_1 _1727_ (.A(_0980_),
    .B(_0994_),
    .Y(_1004_));
 sg13g2_a21oi_1 _1728_ (.A1(_0995_),
    .A2(_1003_),
    .Y(_1005_),
    .B1(_1004_));
 sg13g2_a21o_1 _1729_ (.A2(_1002_),
    .A1(\Voice1.accumulator[6] ),
    .B1(_1004_),
    .X(_1006_));
 sg13g2_nor2b_2 _1730_ (.A(_1005_),
    .B_N(_1006_),
    .Y(_1007_));
 sg13g2_nor2_1 _1731_ (.A(_0967_),
    .B(net51),
    .Y(_1008_));
 sg13g2_and4_1 _1732_ (.A(_0970_),
    .B(_0967_),
    .C(_0965_),
    .D(_0964_),
    .X(_1009_));
 sg13g2_o21ai_1 _1733_ (.B1(net66),
    .Y(_1010_),
    .A1(_1008_),
    .A2(_1009_));
 sg13g2_nand2_2 _1734_ (.Y(_1011_),
    .A(_0965_),
    .B(_0964_));
 sg13g2_nor2b_1 _1735_ (.A(_0963_),
    .B_N(_0967_),
    .Y(_1012_));
 sg13g2_a21oi_1 _1736_ (.A1(_1011_),
    .A2(_1012_),
    .Y(_1013_),
    .B1(_0961_));
 sg13g2_and2_1 _1737_ (.A(_1010_),
    .B(_1013_),
    .X(_1014_));
 sg13g2_o21ai_1 _1738_ (.B1(net66),
    .Y(_1015_),
    .A1(net53),
    .A2(net51));
 sg13g2_a21oi_2 _1739_ (.B1(_0977_),
    .Y(_1016_),
    .A2(_1015_),
    .A1(_1011_));
 sg13g2_and2_1 _1740_ (.A(\Voice1.accumulator[2] ),
    .B(_1016_),
    .X(_1017_));
 sg13g2_a221oi_1 _1741_ (.B2(\Voice1.accumulator[1] ),
    .C1(_1017_),
    .B1(_1014_),
    .A1(\Voice1.accumulator[0] ),
    .Y(_1018_),
    .A2(_0978_));
 sg13g2_nor2_1 _1742_ (.A(\Voice1.accumulator[2] ),
    .B(_1016_),
    .Y(_1019_));
 sg13g2_a221oi_1 _1743_ (.B2(_1013_),
    .C1(\Voice1.accumulator[1] ),
    .B1(_1010_),
    .A1(\Voice1.accumulator[2] ),
    .Y(_1020_),
    .A2(_1016_));
 sg13g2_or2_1 _1744_ (.X(_1021_),
    .B(_1020_),
    .A(_1019_));
 sg13g2_nor2_2 _1745_ (.A(_1018_),
    .B(_1021_),
    .Y(_1022_));
 sg13g2_nand2b_1 _1746_ (.Y(_1023_),
    .B(_0968_),
    .A_N(net66));
 sg13g2_nand3_1 _1747_ (.B(_0981_),
    .C(net49),
    .A(net50),
    .Y(_1024_));
 sg13g2_a21oi_1 _1748_ (.A1(_1023_),
    .A2(_1024_),
    .Y(_1025_),
    .B1(net52));
 sg13g2_a21oi_1 _1749_ (.A1(net50),
    .A2(_1008_),
    .Y(_1026_),
    .B1(_0977_));
 sg13g2_o21ai_1 _1750_ (.B1(_1026_),
    .Y(_1027_),
    .A1(_0981_),
    .A2(_0966_));
 sg13g2_nand3_1 _1751_ (.B(net51),
    .C(net49),
    .A(_0971_),
    .Y(_1028_));
 sg13g2_mux2_1 _1752_ (.A0(_0972_),
    .A1(_1028_),
    .S(_0981_),
    .X(_1029_));
 sg13g2_nor2_1 _1753_ (.A(_0982_),
    .B(_1029_),
    .Y(_1030_));
 sg13g2_nor3_2 _1754_ (.A(_1025_),
    .B(_1027_),
    .C(_1030_),
    .Y(_1031_));
 sg13g2_nand2_1 _1755_ (.Y(_1032_),
    .A(net66),
    .B(net53));
 sg13g2_nor2_1 _1756_ (.A(_0984_),
    .B(_1032_),
    .Y(_1033_));
 sg13g2_a21oi_1 _1757_ (.A1(_0988_),
    .A2(_1023_),
    .Y(_1034_),
    .B1(_0983_));
 sg13g2_nor2_1 _1758_ (.A(_0990_),
    .B(_0977_),
    .Y(_1035_));
 sg13g2_o21ai_1 _1759_ (.B1(_1035_),
    .Y(_1036_),
    .A1(_1033_),
    .A2(_1034_));
 sg13g2_buf_1 _1760_ (.A(_1036_),
    .X(_1037_));
 sg13g2_nand2_1 _1761_ (.Y(_1038_),
    .A(_0971_),
    .B(_0984_));
 sg13g2_nand2b_1 _1762_ (.Y(_1039_),
    .B(_0972_),
    .A_N(_0977_));
 sg13g2_nor3_2 _1763_ (.A(_0975_),
    .B(_1038_),
    .C(_1039_),
    .Y(_1040_));
 sg13g2_nand2_1 _1764_ (.Y(_1041_),
    .A(\Voice1.accumulator[4] ),
    .B(_1040_));
 sg13g2_nand2_1 _1765_ (.Y(_1042_),
    .A(_1037_),
    .B(_1041_));
 sg13g2_nor3_1 _1766_ (.A(_1022_),
    .B(_1031_),
    .C(_1042_),
    .Y(_1043_));
 sg13g2_inv_1 _1767_ (.Y(_1044_),
    .A(\Voice1.accumulator[3] ));
 sg13g2_inv_1 _1768_ (.Y(_1045_),
    .A(\Voice1.accumulator[4] ));
 sg13g2_nor3_1 _1769_ (.A(_1044_),
    .B(_1045_),
    .C(_1037_),
    .Y(_1046_));
 sg13g2_a21oi_1 _1770_ (.A1(_1022_),
    .A2(_1046_),
    .Y(_1047_),
    .B1(\Voice1.accumulator[5] ));
 sg13g2_nor2_1 _1771_ (.A(\Voice1.accumulator[4] ),
    .B(_1040_),
    .Y(_1048_));
 sg13g2_nand2_1 _1772_ (.Y(_1049_),
    .A(_1037_),
    .B(_1048_));
 sg13g2_and3_1 _1773_ (.X(_1050_),
    .A(_1044_),
    .B(_1037_),
    .C(_1041_));
 sg13g2_nand2b_1 _1774_ (.Y(_1051_),
    .B(_1050_),
    .A_N(_1031_));
 sg13g2_o21ai_1 _1775_ (.B1(_1050_),
    .Y(_1052_),
    .A1(_1018_),
    .A2(_1021_));
 sg13g2_nand3_1 _1776_ (.B(_1051_),
    .C(_1052_),
    .A(_1049_),
    .Y(_1053_));
 sg13g2_nor4_2 _1777_ (.A(_1043_),
    .B(_1047_),
    .C(_1053_),
    .Y(_1054_),
    .D(_1005_));
 sg13g2_buf_1 _1778_ (.A(\Voice1.accumulator[9] ),
    .X(_1055_));
 sg13g2_nor3_2 _1779_ (.A(_0977_),
    .B(_1011_),
    .C(_1032_),
    .Y(_1056_));
 sg13g2_nand2_1 _1780_ (.Y(_1057_),
    .A(_1055_),
    .B(_1056_));
 sg13g2_nor2_1 _1781_ (.A(_0982_),
    .B(_0987_),
    .Y(_1058_));
 sg13g2_xnor2_1 _1782_ (.Y(_1059_),
    .A(_0968_),
    .B(net49));
 sg13g2_nor2_1 _1783_ (.A(_0996_),
    .B(_1059_),
    .Y(_1060_));
 sg13g2_o21ai_1 _1784_ (.B1(_1035_),
    .Y(_1061_),
    .A1(_1058_),
    .A2(_1060_));
 sg13g2_buf_1 _1785_ (.A(_1061_),
    .X(_1062_));
 sg13g2_nand2_1 _1786_ (.Y(_1063_),
    .A(_1057_),
    .B(_1062_));
 sg13g2_nor3_2 _1787_ (.A(_1007_),
    .B(_1054_),
    .C(_1063_),
    .Y(_1064_));
 sg13g2_a21oi_1 _1788_ (.A1(_1055_),
    .A2(_1056_),
    .Y(_1065_),
    .B1(\Voice1.accumulator[8] ));
 sg13g2_inv_1 _1789_ (.Y(_1066_),
    .A(_1065_));
 sg13g2_nor3_2 _1790_ (.A(_1007_),
    .B(_1054_),
    .C(_1066_),
    .Y(_1067_));
 sg13g2_nand2_1 _1791_ (.Y(_1068_),
    .A(_1062_),
    .B(_1065_));
 sg13g2_o21ai_1 _1792_ (.B1(_1068_),
    .Y(_1069_),
    .A1(_1055_),
    .A2(_1056_));
 sg13g2_nor3_2 _1793_ (.A(_1064_),
    .B(_1067_),
    .C(_1069_),
    .Y(_1070_));
 sg13g2_nand2_1 _1794_ (.Y(_1071_),
    .A(_1011_),
    .B(_1012_));
 sg13g2_nand3_1 _1795_ (.B(_1071_),
    .C(_1026_),
    .A(_1028_),
    .Y(_1072_));
 sg13g2_xnor2_1 _1796_ (.Y(_1073_),
    .A(_1070_),
    .B(_1072_));
 sg13g2_nand2_1 _1797_ (.Y(_1074_),
    .A(_0962_),
    .B(_1073_));
 sg13g2_xnor2_1 _1798_ (.Y(_0026_),
    .A(\Voice1.accumulator[10] ),
    .B(_1074_));
 sg13g2_and3_1 _1799_ (.X(_1075_),
    .A(_1028_),
    .B(_1071_),
    .C(_1026_));
 sg13g2_buf_1 _1800_ (.A(_1075_),
    .X(_1076_));
 sg13g2_nor2_1 _1801_ (.A(_1070_),
    .B(_1076_),
    .Y(_1077_));
 sg13g2_a21oi_1 _1802_ (.A1(_1070_),
    .A2(_1076_),
    .Y(_1078_),
    .B1(\Voice1.accumulator[10] ));
 sg13g2_or2_1 _1803_ (.X(_1079_),
    .B(_1039_),
    .A(_1038_));
 sg13g2_o21ai_1 _1804_ (.B1(_1079_),
    .Y(_1080_),
    .A1(_1077_),
    .A2(_1078_));
 sg13g2_nor2_1 _1805_ (.A(_1038_),
    .B(_1039_),
    .Y(_1081_));
 sg13g2_nand3_1 _1806_ (.B(_1081_),
    .C(_1070_),
    .A(\Voice1.accumulator[10] ),
    .Y(_1082_));
 sg13g2_nand3_1 _1807_ (.B(_1080_),
    .C(_1082_),
    .A(_0962_),
    .Y(_1083_));
 sg13g2_xnor2_1 _1808_ (.Y(_0027_),
    .A(\Voice1.accumulator[11] ),
    .B(_1083_));
 sg13g2_buf_1 _1809_ (.A(\Voice1.accumulator[12] ),
    .X(_1084_));
 sg13g2_or2_1 _1810_ (.X(_1085_),
    .B(_1081_),
    .A(\Voice1.accumulator[11] ));
 sg13g2_buf_1 _1811_ (.A(_1085_),
    .X(_1086_));
 sg13g2_o21ai_1 _1812_ (.B1(_1086_),
    .Y(_1087_),
    .A1(_1070_),
    .A2(_1076_));
 sg13g2_nand2_1 _1813_ (.Y(_1088_),
    .A(\Voice1.accumulator[11] ),
    .B(_1081_));
 sg13g2_o21ai_1 _1814_ (.B1(_1088_),
    .Y(_1089_),
    .A1(_1078_),
    .A2(_1087_));
 sg13g2_nand2_1 _1815_ (.Y(_1090_),
    .A(_0962_),
    .B(_1089_));
 sg13g2_xnor2_1 _1816_ (.Y(_0028_),
    .A(_1084_),
    .B(_1090_));
 sg13g2_buf_1 _1817_ (.A(_0959_),
    .X(_1091_));
 sg13g2_nand2_1 _1818_ (.Y(_1092_),
    .A(net65),
    .B(\Voice1.en ));
 sg13g2_buf_1 _1819_ (.A(_1092_),
    .X(_1093_));
 sg13g2_buf_1 _1820_ (.A(_1093_),
    .X(_1094_));
 sg13g2_nand3_1 _1821_ (.B(_1076_),
    .C(_1086_),
    .A(_1084_),
    .Y(_1095_));
 sg13g2_nor4_1 _1822_ (.A(_1064_),
    .B(_1067_),
    .C(_1069_),
    .D(_1095_),
    .Y(_1096_));
 sg13g2_nand3_1 _1823_ (.B(\Voice1.accumulator[10] ),
    .C(_1086_),
    .A(_1084_),
    .Y(_1097_));
 sg13g2_nor4_1 _1824_ (.A(_1064_),
    .B(_1067_),
    .C(_1069_),
    .D(_1097_),
    .Y(_1098_));
 sg13g2_nand3_1 _1825_ (.B(\Voice1.accumulator[11] ),
    .C(_1081_),
    .A(_1084_),
    .Y(_1099_));
 sg13g2_o21ai_1 _1826_ (.B1(_1099_),
    .Y(_1100_),
    .A1(_1072_),
    .A2(_1097_));
 sg13g2_nor3_2 _1827_ (.A(_1096_),
    .B(_1098_),
    .C(_1100_),
    .Y(_1101_));
 sg13g2_xnor2_1 _1828_ (.Y(_1102_),
    .A(_0002_),
    .B(_1101_));
 sg13g2_nand2_1 _1829_ (.Y(_1103_),
    .A(\Voice1.accumulator[13] ),
    .B(net23));
 sg13g2_o21ai_1 _1830_ (.B1(_1103_),
    .Y(_0029_),
    .A1(net23),
    .A2(_1102_));
 sg13g2_buf_1 _1831_ (.A(\Voice1.accumulator[14] ),
    .X(_1104_));
 sg13g2_or3_1 _1832_ (.A(_0002_),
    .B(_1093_),
    .C(_1101_),
    .X(_1105_));
 sg13g2_buf_2 _1833_ (.A(_1105_),
    .X(_1106_));
 sg13g2_xnor2_1 _1834_ (.Y(_0030_),
    .A(_1104_),
    .B(_1106_));
 sg13g2_buf_1 _1835_ (.A(\Voice1.accumulator[15] ),
    .X(_1107_));
 sg13g2_inv_1 _1836_ (.Y(_1108_),
    .A(\Voice1.accumulator[13] ));
 sg13g2_nor3_1 _1837_ (.A(_1108_),
    .B(_1093_),
    .C(_1101_),
    .Y(_1109_));
 sg13g2_nand2_1 _1838_ (.Y(_1110_),
    .A(_1104_),
    .B(_1109_));
 sg13g2_xnor2_1 _1839_ (.Y(_0031_),
    .A(_1107_),
    .B(_1110_));
 sg13g2_inv_1 _1840_ (.Y(_1111_),
    .A(\Voice1.accumulator[16] ));
 sg13g2_inv_1 _1841_ (.Y(_1112_),
    .A(_1107_));
 sg13g2_inv_1 _1842_ (.Y(_1113_),
    .A(_1104_));
 sg13g2_nor3_1 _1843_ (.A(_1112_),
    .B(_1113_),
    .C(_1106_),
    .Y(_1114_));
 sg13g2_xnor2_1 _1844_ (.Y(_0032_),
    .A(_1111_),
    .B(_1114_));
 sg13g2_inv_1 _1845_ (.Y(_1115_),
    .A(\Voice1.accumulator[17] ));
 sg13g2_nand3_1 _1846_ (.B(_1107_),
    .C(_1104_),
    .A(\Voice1.accumulator[16] ),
    .Y(_1116_));
 sg13g2_buf_1 _1847_ (.A(_1116_),
    .X(_1117_));
 sg13g2_nor4_1 _1848_ (.A(_1108_),
    .B(_1093_),
    .C(_1101_),
    .D(_1117_),
    .Y(_1118_));
 sg13g2_xnor2_1 _1849_ (.Y(_0033_),
    .A(_1115_),
    .B(_1118_));
 sg13g2_buf_1 _1850_ (.A(\Voice1.accumulator[18] ),
    .X(_1119_));
 sg13g2_nor3_1 _1851_ (.A(_1115_),
    .B(_1106_),
    .C(_1117_),
    .Y(_1120_));
 sg13g2_xor2_1 _1852_ (.B(_1120_),
    .A(_1119_),
    .X(_0034_));
 sg13g2_nand2_1 _1853_ (.Y(_1121_),
    .A(_1119_),
    .B(\Voice1.accumulator[17] ));
 sg13g2_nor2_1 _1854_ (.A(_1117_),
    .B(_1121_),
    .Y(_1122_));
 sg13g2_nand2_1 _1855_ (.Y(_1123_),
    .A(_1109_),
    .B(_1122_));
 sg13g2_xnor2_1 _1856_ (.Y(_0035_),
    .A(\Voice1.accumulator[19] ),
    .B(_1123_));
 sg13g2_nand2_1 _1857_ (.Y(_1124_),
    .A(\Voice1.accumulator[0] ),
    .B(_0978_));
 sg13g2_xnor2_1 _1858_ (.Y(_1125_),
    .A(_1124_),
    .B(_1014_));
 sg13g2_nand2_1 _1859_ (.Y(_1126_),
    .A(_0962_),
    .B(_1125_));
 sg13g2_xnor2_1 _1860_ (.Y(_0036_),
    .A(\Voice1.accumulator[1] ),
    .B(_1126_));
 sg13g2_buf_1 _1861_ (.A(\Voice1.accumulator[20] ),
    .X(_1127_));
 sg13g2_inv_1 _1862_ (.Y(_1128_),
    .A(\Voice1.accumulator[19] ));
 sg13g2_nor3_1 _1863_ (.A(_1128_),
    .B(_1117_),
    .C(_1121_),
    .Y(_1129_));
 sg13g2_nand2b_1 _1864_ (.Y(_1130_),
    .B(_1129_),
    .A_N(_1106_));
 sg13g2_xnor2_1 _1865_ (.Y(_0037_),
    .A(_1127_),
    .B(_1130_));
 sg13g2_nand2_1 _1866_ (.Y(_1131_),
    .A(_1127_),
    .B(_1129_));
 sg13g2_nor3_1 _1867_ (.A(_1108_),
    .B(_1101_),
    .C(_1131_),
    .Y(_1132_));
 sg13g2_xor2_1 _1868_ (.B(_1132_),
    .A(_0005_),
    .X(_1133_));
 sg13g2_nand2_1 _1869_ (.Y(_1134_),
    .A(\Voice1.accumulator[21] ),
    .B(net23));
 sg13g2_o21ai_1 _1870_ (.B1(_1134_),
    .Y(_0038_),
    .A1(net23),
    .A2(_1133_));
 sg13g2_inv_1 _1871_ (.Y(_1135_),
    .A(\Voice1.accumulator[22] ));
 sg13g2_nand3_1 _1872_ (.B(\Voice1.accumulator[21] ),
    .C(_1129_),
    .A(_1127_),
    .Y(_1136_));
 sg13g2_nor2_1 _1873_ (.A(_1106_),
    .B(_1136_),
    .Y(_1137_));
 sg13g2_xnor2_1 _1874_ (.Y(_0039_),
    .A(_1135_),
    .B(_1137_));
 sg13g2_inv_1 _1875_ (.Y(_1138_),
    .A(_0004_));
 sg13g2_nor4_1 _1876_ (.A(_1135_),
    .B(_1108_),
    .C(_1101_),
    .D(_1136_),
    .Y(_1139_));
 sg13g2_xnor2_1 _1877_ (.Y(_1140_),
    .A(_1138_),
    .B(_1139_));
 sg13g2_nand2_1 _1878_ (.Y(_1141_),
    .A(\Voice1.accumulator[23] ),
    .B(net23));
 sg13g2_o21ai_1 _1879_ (.B1(_1141_),
    .Y(_0040_),
    .A1(net23),
    .A2(_1140_));
 sg13g2_nand2_1 _1880_ (.Y(_1142_),
    .A(_1010_),
    .B(_1013_));
 sg13g2_nand2_1 _1881_ (.Y(_1143_),
    .A(_1124_),
    .B(_1142_));
 sg13g2_nor2_1 _1882_ (.A(_1124_),
    .B(_1142_),
    .Y(_1144_));
 sg13g2_a21oi_1 _1883_ (.A1(\Voice1.accumulator[1] ),
    .A2(_1143_),
    .Y(_1145_),
    .B1(_1144_));
 sg13g2_xor2_1 _1884_ (.B(_1145_),
    .A(_1016_),
    .X(_1146_));
 sg13g2_nor2_1 _1885_ (.A(net23),
    .B(_1146_),
    .Y(_1147_));
 sg13g2_xor2_1 _1886_ (.B(_1147_),
    .A(\Voice1.accumulator[2] ),
    .X(_0041_));
 sg13g2_xnor2_1 _1887_ (.Y(_1148_),
    .A(_1022_),
    .B(_1031_));
 sg13g2_nor2_1 _1888_ (.A(net23),
    .B(_1148_),
    .Y(_1149_));
 sg13g2_xnor2_1 _1889_ (.Y(_0042_),
    .A(_1044_),
    .B(_1149_));
 sg13g2_nor2_1 _1890_ (.A(_1022_),
    .B(_1031_),
    .Y(_1150_));
 sg13g2_a21oi_1 _1891_ (.A1(_1022_),
    .A2(_1031_),
    .Y(_1151_),
    .B1(\Voice1.accumulator[3] ));
 sg13g2_nor2_1 _1892_ (.A(_1150_),
    .B(_1151_),
    .Y(_1152_));
 sg13g2_xnor2_1 _1893_ (.Y(_1153_),
    .A(_1040_),
    .B(_1152_));
 sg13g2_nor2_1 _1894_ (.A(_1094_),
    .B(_1153_),
    .Y(_1154_));
 sg13g2_xnor2_1 _1895_ (.Y(_0043_),
    .A(_1045_),
    .B(_1154_));
 sg13g2_nand2_1 _1896_ (.Y(_1155_),
    .A(_1022_),
    .B(_1046_));
 sg13g2_o21ai_1 _1897_ (.B1(\Voice1.accumulator[4] ),
    .Y(_1156_),
    .A1(_1040_),
    .A2(_1152_));
 sg13g2_nand2_1 _1898_ (.Y(_1157_),
    .A(_1040_),
    .B(_1152_));
 sg13g2_nand3_1 _1899_ (.B(_1156_),
    .C(_1157_),
    .A(_1037_),
    .Y(_1158_));
 sg13g2_and3_1 _1900_ (.X(_1159_),
    .A(_0962_),
    .B(_1155_),
    .C(_1158_));
 sg13g2_xor2_1 _1901_ (.B(_1159_),
    .A(\Voice1.accumulator[5] ),
    .X(_0044_));
 sg13g2_inv_1 _1902_ (.Y(_1160_),
    .A(_1002_));
 sg13g2_or3_1 _1903_ (.A(_1043_),
    .B(_1047_),
    .C(_1053_),
    .X(_1161_));
 sg13g2_buf_1 _1904_ (.A(_1161_),
    .X(_1162_));
 sg13g2_xnor2_1 _1905_ (.Y(_1163_),
    .A(_1160_),
    .B(_1162_));
 sg13g2_nor2_1 _1906_ (.A(_1093_),
    .B(_1163_),
    .Y(_1164_));
 sg13g2_xor2_1 _1907_ (.B(_1164_),
    .A(\Voice1.accumulator[6] ),
    .X(_0045_));
 sg13g2_nand2_1 _1908_ (.Y(_1165_),
    .A(_1160_),
    .B(_1162_));
 sg13g2_nor2_1 _1909_ (.A(_1160_),
    .B(_1162_),
    .Y(_1166_));
 sg13g2_a21oi_1 _1910_ (.A1(\Voice1.accumulator[6] ),
    .A2(_1165_),
    .Y(_1167_),
    .B1(_1166_));
 sg13g2_xnor2_1 _1911_ (.Y(_1168_),
    .A(_0994_),
    .B(_1167_));
 sg13g2_nor2_1 _1912_ (.A(_1094_),
    .B(_1168_),
    .Y(_1169_));
 sg13g2_xnor2_1 _1913_ (.Y(_0046_),
    .A(_0980_),
    .B(_1169_));
 sg13g2_nor2_1 _1914_ (.A(_1007_),
    .B(_1054_),
    .Y(_1170_));
 sg13g2_xnor2_1 _1915_ (.Y(_1171_),
    .A(_1170_),
    .B(_1062_));
 sg13g2_nor2_1 _1916_ (.A(_1093_),
    .B(_1171_),
    .Y(_1172_));
 sg13g2_xor2_1 _1917_ (.B(_1172_),
    .A(\Voice1.accumulator[8] ),
    .X(_0047_));
 sg13g2_nand2_1 _1918_ (.Y(_1173_),
    .A(_1170_),
    .B(_1062_));
 sg13g2_nor2_1 _1919_ (.A(_1170_),
    .B(_1062_),
    .Y(_1174_));
 sg13g2_a21oi_1 _1920_ (.A1(\Voice1.accumulator[8] ),
    .A2(_1173_),
    .Y(_1175_),
    .B1(_1174_));
 sg13g2_xor2_1 _1921_ (.B(_1175_),
    .A(_1056_),
    .X(_1176_));
 sg13g2_nor2_1 _1922_ (.A(_1093_),
    .B(_1176_),
    .Y(_1177_));
 sg13g2_xor2_1 _1923_ (.B(_1177_),
    .A(_1055_),
    .X(_0048_));
 sg13g2_buf_1 _1924_ (.A(\hvsync_gen.vpos[0] ),
    .X(_1178_));
 sg13g2_buf_2 _1925_ (.A(\hvsync_gen.hpos[3] ),
    .X(_1179_));
 sg13g2_inv_1 _1926_ (.Y(_1180_),
    .A(_1179_));
 sg13g2_buf_2 _1927_ (.A(\hvsync_gen.hpos[2] ),
    .X(_1181_));
 sg13g2_nand3_1 _1928_ (.B(\hvsync_gen.hpos[1] ),
    .C(_1181_),
    .A(\hvsync_gen.hpos[0] ),
    .Y(_1182_));
 sg13g2_nor2_1 _1929_ (.A(_1180_),
    .B(_1182_),
    .Y(_1183_));
 sg13g2_and2_1 _1930_ (.A(net67),
    .B(_1183_),
    .X(_1184_));
 sg13g2_buf_1 _1931_ (.A(_1184_),
    .X(_1185_));
 sg13g2_nand2_1 _1932_ (.Y(_1186_),
    .A(net56),
    .B(net55));
 sg13g2_nor4_1 _1933_ (.A(net70),
    .B(net68),
    .C(net54),
    .D(_1186_),
    .Y(_1187_));
 sg13g2_and2_1 _1934_ (.A(_1185_),
    .B(_1187_),
    .X(_1188_));
 sg13g2_nor2_1 _1935_ (.A(_0960_),
    .B(_1188_),
    .Y(_1189_));
 sg13g2_buf_1 _1936_ (.A(_1189_),
    .X(_1190_));
 sg13g2_inv_2 _1937_ (.Y(_1191_),
    .A(net73));
 sg13g2_nor4_1 _1938_ (.A(_0923_),
    .B(net35),
    .C(net59),
    .D(_1191_),
    .Y(_1192_));
 sg13g2_nor2b_1 _1939_ (.A(_0943_),
    .B_N(_1192_),
    .Y(_1193_));
 sg13g2_inv_1 _1940_ (.Y(_1194_),
    .A(_0924_));
 sg13g2_nor4_1 _1941_ (.A(_1178_),
    .B(_1194_),
    .C(net72),
    .D(net36),
    .Y(_1195_));
 sg13g2_a21oi_2 _1942_ (.B1(_0960_),
    .Y(_1196_),
    .A2(_1195_),
    .A1(_1193_));
 sg13g2_and2_1 _1943_ (.A(_1188_),
    .B(_1196_),
    .X(_1197_));
 sg13g2_buf_2 _1944_ (.A(_1197_),
    .X(_1198_));
 sg13g2_a22oi_1 _1945_ (.Y(_1199_),
    .B1(_1198_),
    .B2(_0014_),
    .A2(net16),
    .A1(_1178_));
 sg13g2_inv_1 _1946_ (.Y(_0117_),
    .A(_1199_));
 sg13g2_nand2_1 _1947_ (.Y(_1200_),
    .A(_1178_),
    .B(_1198_));
 sg13g2_nor2b_1 _1948_ (.A(_1178_),
    .B_N(_1198_),
    .Y(_1201_));
 sg13g2_o21ai_1 _1949_ (.B1(_0923_),
    .Y(_1202_),
    .A1(net16),
    .A2(_1201_));
 sg13g2_o21ai_1 _1950_ (.B1(_1202_),
    .Y(_0118_),
    .A1(_0923_),
    .A2(_1200_));
 sg13g2_nand2_1 _1951_ (.Y(_1203_),
    .A(_0923_),
    .B(_1178_));
 sg13g2_nor3_1 _1952_ (.A(_0924_),
    .B(net16),
    .C(_1203_),
    .Y(_1204_));
 sg13g2_a21o_1 _1953_ (.A2(_1203_),
    .A1(_0924_),
    .B1(_1204_),
    .X(_1205_));
 sg13g2_a22oi_1 _1954_ (.Y(_1206_),
    .B1(_1196_),
    .B2(_1205_),
    .A2(_1190_),
    .A1(_0924_));
 sg13g2_inv_1 _1955_ (.Y(_0119_),
    .A(_1206_));
 sg13g2_nor2_1 _1956_ (.A(_1194_),
    .B(_1203_),
    .Y(_1207_));
 sg13g2_nand2_1 _1957_ (.Y(_1208_),
    .A(_1198_),
    .B(_1207_));
 sg13g2_inv_1 _1958_ (.Y(_1209_),
    .A(_1196_));
 sg13g2_nand2b_1 _1959_ (.Y(_1210_),
    .B(net65),
    .A_N(_1188_));
 sg13g2_buf_2 _1960_ (.A(_1210_),
    .X(_1211_));
 sg13g2_o21ai_1 _1961_ (.B1(_1211_),
    .Y(_1212_),
    .A1(_1209_),
    .A2(_1207_));
 sg13g2_nand2_1 _1962_ (.Y(_1213_),
    .A(net58),
    .B(_1212_));
 sg13g2_o21ai_1 _1963_ (.B1(_1213_),
    .Y(_0120_),
    .A1(net58),
    .A2(_1208_));
 sg13g2_a21oi_1 _1964_ (.A1(_0939_),
    .A2(_1207_),
    .Y(_1214_),
    .B1(_1209_));
 sg13g2_o21ai_1 _1965_ (.B1(_0941_),
    .Y(_1215_),
    .A1(net16),
    .A2(_1214_));
 sg13g2_o21ai_1 _1966_ (.B1(_1215_),
    .Y(_0121_),
    .A1(_0943_),
    .A2(_1208_));
 sg13g2_and3_1 _1967_ (.X(_1216_),
    .A(_0939_),
    .B(_0941_),
    .C(_1207_));
 sg13g2_buf_2 _1968_ (.A(_1216_),
    .X(_1217_));
 sg13g2_nand2_1 _1969_ (.Y(_1218_),
    .A(_1198_),
    .B(_1217_));
 sg13g2_o21ai_1 _1970_ (.B1(_1211_),
    .Y(_1219_),
    .A1(_1209_),
    .A2(_1217_));
 sg13g2_nand2_1 _1971_ (.Y(_1220_),
    .A(net62),
    .B(_1219_));
 sg13g2_o21ai_1 _1972_ (.B1(_1220_),
    .Y(_0122_),
    .A1(net62),
    .A2(_1218_));
 sg13g2_nand3_1 _1973_ (.B(_1198_),
    .C(_1217_),
    .A(net62),
    .Y(_1221_));
 sg13g2_a21oi_1 _1974_ (.A1(net62),
    .A2(_1217_),
    .Y(_1222_),
    .B1(_1209_));
 sg13g2_o21ai_1 _1975_ (.B1(net35),
    .Y(_1223_),
    .A1(net16),
    .A2(_1222_));
 sg13g2_o21ai_1 _1976_ (.B1(_1223_),
    .Y(_0123_),
    .A1(net35),
    .A2(_1221_));
 sg13g2_nand4_1 _1977_ (.B(net35),
    .C(_1198_),
    .A(net62),
    .Y(_1224_),
    .D(_1217_));
 sg13g2_nand3_1 _1978_ (.B(_0933_),
    .C(_1217_),
    .A(_0927_),
    .Y(_1225_));
 sg13g2_and2_1 _1979_ (.A(_1196_),
    .B(_1225_),
    .X(_1226_));
 sg13g2_o21ai_1 _1980_ (.B1(net36),
    .Y(_1227_),
    .A1(net16),
    .A2(_1226_));
 sg13g2_o21ai_1 _1981_ (.B1(_1227_),
    .Y(_0124_),
    .A1(net36),
    .A2(_1224_));
 sg13g2_nand2b_1 _1982_ (.Y(_1228_),
    .B(net36),
    .A_N(net59));
 sg13g2_nand4_1 _1983_ (.B(net36),
    .C(_0933_),
    .A(_0927_),
    .Y(_1229_),
    .D(_1217_));
 sg13g2_and2_1 _1984_ (.A(_1196_),
    .B(_1229_),
    .X(_1230_));
 sg13g2_o21ai_1 _1985_ (.B1(net59),
    .Y(_1231_),
    .A1(net16),
    .A2(_1230_));
 sg13g2_o21ai_1 _1986_ (.B1(_1231_),
    .Y(_0125_),
    .A1(_1224_),
    .A2(_1228_));
 sg13g2_nand2b_1 _1987_ (.Y(_1232_),
    .B(_1217_),
    .A_N(_0937_));
 sg13g2_a21oi_1 _1988_ (.A1(_1196_),
    .A2(_1232_),
    .Y(_1233_),
    .B1(net16));
 sg13g2_or3_1 _1989_ (.A(_0925_),
    .B(_0937_),
    .C(_1218_),
    .X(_1234_));
 sg13g2_o21ai_1 _1990_ (.B1(_1234_),
    .Y(_0126_),
    .A1(_1191_),
    .A2(_1233_));
 sg13g2_buf_1 _1991_ (.A(_0960_),
    .X(_1235_));
 sg13g2_nor2_1 _1992_ (.A(net48),
    .B(net74),
    .Y(_1236_));
 sg13g2_buf_1 _1993_ (.A(\LFSR[2] ),
    .X(_1237_));
 sg13g2_buf_1 _1994_ (.A(\LFSR[1] ),
    .X(_1238_));
 sg13g2_xnor2_1 _1995_ (.Y(_1239_),
    .A(_1237_),
    .B(_1238_));
 sg13g2_nand2_1 _1996_ (.Y(_0019_),
    .A(_1236_),
    .B(_1239_));
 sg13g2_inv_1 _1997_ (.Y(_1240_),
    .A(\LFSR[0] ));
 sg13g2_nand2b_1 _1998_ (.Y(_1241_),
    .B(net65),
    .A_N(net74));
 sg13g2_buf_1 _1999_ (.A(_1241_),
    .X(_1242_));
 sg13g2_buf_1 _2000_ (.A(_1242_),
    .X(_1243_));
 sg13g2_nor2_1 _2001_ (.A(_1240_),
    .B(net22),
    .Y(_0020_));
 sg13g2_and2_1 _2002_ (.A(_1238_),
    .B(_1236_),
    .X(_0021_));
 sg13g2_inv_1 _2003_ (.Y(_1244_),
    .A(_1237_));
 sg13g2_nor2_1 _2004_ (.A(_1244_),
    .B(net22),
    .Y(_0022_));
 sg13g2_buf_1 _2005_ (.A(\LFSR[3] ),
    .X(_1245_));
 sg13g2_and2_1 _2006_ (.A(_1245_),
    .B(_1236_),
    .X(_0023_));
 sg13g2_inv_1 _2007_ (.Y(_1246_),
    .A(\LFSR[4] ));
 sg13g2_nor2_1 _2008_ (.A(_1246_),
    .B(net22),
    .Y(_0024_));
 sg13g2_inv_1 _2009_ (.Y(_1247_),
    .A(_0016_));
 sg13g2_buf_2 _2010_ (.A(\ctr_clkdiv25[4] ),
    .X(_1248_));
 sg13g2_nor2b_1 _2011_ (.A(\ctr_clkdiv25[6] ),
    .B_N(_1248_),
    .Y(_1249_));
 sg13g2_and2_1 _2012_ (.A(\ctr_clkdiv25[0] ),
    .B(\ctr_clkdiv25[3] ),
    .X(_1250_));
 sg13g2_nor4_1 _2013_ (.A(\ctr_clkdiv25[1] ),
    .B(\ctr_clkdiv25[2] ),
    .C(\ctr_clkdiv25[5] ),
    .D(\ctr_clkdiv25[7] ),
    .Y(_1251_));
 sg13g2_and3_1 _2014_ (.X(_1252_),
    .A(_1249_),
    .B(_1250_),
    .C(_1251_));
 sg13g2_buf_1 _2015_ (.A(_1252_),
    .X(_1253_));
 sg13g2_nand2b_1 _2016_ (.Y(_1254_),
    .B(net65),
    .A_N(_1253_));
 sg13g2_buf_2 _2017_ (.A(_1254_),
    .X(_1255_));
 sg13g2_nor2_1 _2018_ (.A(_1247_),
    .B(_1255_),
    .Y(_0091_));
 sg13g2_xnor2_1 _2019_ (.Y(_1256_),
    .A(\ctr_clkdiv25[0] ),
    .B(\ctr_clkdiv25[1] ));
 sg13g2_nor2_1 _2020_ (.A(_1255_),
    .B(_1256_),
    .Y(_0092_));
 sg13g2_buf_1 _2021_ (.A(net48),
    .X(_1257_));
 sg13g2_nand2_1 _2022_ (.Y(_1258_),
    .A(\ctr_clkdiv25[0] ),
    .B(\ctr_clkdiv25[1] ));
 sg13g2_xor2_1 _2023_ (.B(_1258_),
    .A(\ctr_clkdiv25[2] ),
    .X(_1259_));
 sg13g2_nor2_1 _2024_ (.A(_1257_),
    .B(_1259_),
    .Y(_0093_));
 sg13g2_inv_1 _2025_ (.Y(_1260_),
    .A(\ctr_clkdiv25[3] ));
 sg13g2_nand3_1 _2026_ (.B(\ctr_clkdiv25[1] ),
    .C(\ctr_clkdiv25[2] ),
    .A(\ctr_clkdiv25[0] ),
    .Y(_1261_));
 sg13g2_xnor2_1 _2027_ (.Y(_1262_),
    .A(_1260_),
    .B(_1261_));
 sg13g2_nor2_1 _2028_ (.A(_1255_),
    .B(_1262_),
    .Y(_0094_));
 sg13g2_nor2_2 _2029_ (.A(_1260_),
    .B(_1261_),
    .Y(_1263_));
 sg13g2_xnor2_1 _2030_ (.Y(_1264_),
    .A(_1248_),
    .B(_1263_));
 sg13g2_nor2_1 _2031_ (.A(_1255_),
    .B(_1264_),
    .Y(_0095_));
 sg13g2_nand2_1 _2032_ (.Y(_1265_),
    .A(_1248_),
    .B(_1263_));
 sg13g2_xor2_1 _2033_ (.B(_1265_),
    .A(\ctr_clkdiv25[5] ),
    .X(_1266_));
 sg13g2_nor2_1 _2034_ (.A(_1255_),
    .B(_1266_),
    .Y(_0096_));
 sg13g2_nand3_1 _2035_ (.B(_1248_),
    .C(_1263_),
    .A(\ctr_clkdiv25[5] ),
    .Y(_1267_));
 sg13g2_xor2_1 _2036_ (.B(_1267_),
    .A(\ctr_clkdiv25[6] ),
    .X(_1268_));
 sg13g2_nor2_1 _2037_ (.A(_1255_),
    .B(_1268_),
    .Y(_0097_));
 sg13g2_nand4_1 _2038_ (.B(_1248_),
    .C(\ctr_clkdiv25[6] ),
    .A(\ctr_clkdiv25[5] ),
    .Y(_1269_),
    .D(_1263_));
 sg13g2_xor2_1 _2039_ (.B(_1269_),
    .A(\ctr_clkdiv25[7] ),
    .X(_1270_));
 sg13g2_nor2_1 _2040_ (.A(_1255_),
    .B(_1270_),
    .Y(_0098_));
 sg13g2_and2_1 _2041_ (.A(_0018_),
    .B(_1190_),
    .X(_0107_));
 sg13g2_xnor2_1 _2042_ (.Y(_1271_),
    .A(\hvsync_gen.hpos[0] ),
    .B(\hvsync_gen.hpos[1] ));
 sg13g2_nor2_1 _2043_ (.A(_1211_),
    .B(_1271_),
    .Y(_0108_));
 sg13g2_nand2_1 _2044_ (.Y(_1272_),
    .A(\hvsync_gen.hpos[0] ),
    .B(\hvsync_gen.hpos[1] ));
 sg13g2_xor2_1 _2045_ (.B(_1272_),
    .A(_1181_),
    .X(_1273_));
 sg13g2_nor2_1 _2046_ (.A(_1211_),
    .B(_1273_),
    .Y(_0109_));
 sg13g2_xnor2_1 _2047_ (.Y(_1274_),
    .A(_1180_),
    .B(_1182_));
 sg13g2_nor2_1 _2048_ (.A(net34),
    .B(_1274_),
    .Y(_0110_));
 sg13g2_xnor2_1 _2049_ (.Y(_1275_),
    .A(net67),
    .B(_1183_));
 sg13g2_nor2_1 _2050_ (.A(net34),
    .B(_1275_),
    .Y(_0111_));
 sg13g2_xnor2_1 _2051_ (.Y(_1276_),
    .A(net54),
    .B(_1185_));
 sg13g2_nor2_1 _2052_ (.A(_1211_),
    .B(_1276_),
    .Y(_0112_));
 sg13g2_inv_1 _2053_ (.Y(_1277_),
    .A(\hvsync_gen.hpos[6] ));
 sg13g2_nand2_1 _2054_ (.Y(_1278_),
    .A(net54),
    .B(_1185_));
 sg13g2_xnor2_1 _2055_ (.Y(_1279_),
    .A(_1277_),
    .B(_1278_));
 sg13g2_nor2_1 _2056_ (.A(net34),
    .B(_1279_),
    .Y(_0113_));
 sg13g2_nand3_1 _2057_ (.B(net54),
    .C(_1185_),
    .A(net68),
    .Y(_1280_));
 sg13g2_xor2_1 _2058_ (.B(_1280_),
    .A(net70),
    .X(_1281_));
 sg13g2_nor2_1 _2059_ (.A(net34),
    .B(_1281_),
    .Y(_0114_));
 sg13g2_nand4_1 _2060_ (.B(_0951_),
    .C(net54),
    .A(net70),
    .Y(_1282_),
    .D(_1185_));
 sg13g2_xnor2_1 _2061_ (.Y(_1283_),
    .A(_0956_),
    .B(_1282_));
 sg13g2_nor2_1 _2062_ (.A(_1211_),
    .B(_1283_),
    .Y(_0115_));
 sg13g2_inv_1 _2063_ (.Y(_1284_),
    .A(net69));
 sg13g2_or2_1 _2064_ (.X(_1285_),
    .B(_1282_),
    .A(_0956_));
 sg13g2_xnor2_1 _2065_ (.Y(_1286_),
    .A(net47),
    .B(_1285_));
 sg13g2_nor2_1 _2066_ (.A(_1211_),
    .B(_1286_),
    .Y(_0116_));
 sg13g2_buf_2 _2067_ (.A(hsync),
    .X(_1287_));
 sg13g2_nand2b_1 _2068_ (.Y(_1288_),
    .B(net65),
    .A_N(_1287_));
 sg13g2_inv_1 _2069_ (.Y(_1289_),
    .A(\xqo[0] ));
 sg13g2_buf_2 _2070_ (.A(\counter[3] ),
    .X(_1290_));
 sg13g2_inv_1 _2071_ (.Y(_1291_),
    .A(_1290_));
 sg13g2_buf_8 _2072_ (.A(\counter[2] ),
    .X(_1292_));
 sg13g2_nand2_1 _2073_ (.Y(_1293_),
    .A(_0952_),
    .B(net46));
 sg13g2_nor2_1 _2074_ (.A(_0952_),
    .B(net46),
    .Y(_1294_));
 sg13g2_buf_8 _2075_ (.A(\counter[1] ),
    .X(_1295_));
 sg13g2_nor2_1 _2076_ (.A(net67),
    .B(_1295_),
    .Y(_1296_));
 sg13g2_buf_8 _2077_ (.A(\counter[0] ),
    .X(_1297_));
 sg13g2_a22oi_1 _2078_ (.Y(_1298_),
    .B1(_1297_),
    .B2(_1179_),
    .A2(_1295_),
    .A1(_0954_));
 sg13g2_or3_1 _2079_ (.A(_1294_),
    .B(_1296_),
    .C(_1298_),
    .X(_1299_));
 sg13g2_a22oi_1 _2080_ (.Y(_1300_),
    .B1(_1293_),
    .B2(_1299_),
    .A2(_1291_),
    .A1(_1277_));
 sg13g2_buf_1 _2081_ (.A(_1300_),
    .X(_1301_));
 sg13g2_buf_1 _2082_ (.A(\counter[4] ),
    .X(_1302_));
 sg13g2_nand2_1 _2083_ (.Y(_1303_),
    .A(\hvsync_gen.hpos[7] ),
    .B(_1302_));
 sg13g2_o21ai_1 _2084_ (.B1(_1303_),
    .Y(_1304_),
    .A1(_1277_),
    .A2(_1291_));
 sg13g2_buf_1 _2085_ (.A(_1304_),
    .X(_1305_));
 sg13g2_buf_1 _2086_ (.A(_1302_),
    .X(_1306_));
 sg13g2_or2_1 _2087_ (.X(_1307_),
    .B(net33),
    .A(_0945_));
 sg13g2_o21ai_1 _2088_ (.B1(_1307_),
    .Y(_1308_),
    .A1(_1301_),
    .A2(_1305_));
 sg13g2_buf_1 _2089_ (.A(\counter[5] ),
    .X(_1309_));
 sg13g2_buf_1 _2090_ (.A(\counter[8] ),
    .X(_1310_));
 sg13g2_xnor2_1 _2091_ (.Y(_1311_),
    .A(net45),
    .B(net44));
 sg13g2_xnor2_1 _2092_ (.Y(_1312_),
    .A(_0946_),
    .B(_1311_));
 sg13g2_xnor2_1 _2093_ (.Y(_1313_),
    .A(_1308_),
    .B(_1312_));
 sg13g2_buf_1 _2094_ (.A(\counter[6] ),
    .X(_1314_));
 sg13g2_inv_1 _2095_ (.Y(_1315_),
    .A(_1314_));
 sg13g2_nor2_1 _2096_ (.A(_0945_),
    .B(_1302_),
    .Y(_1316_));
 sg13g2_nor2_1 _2097_ (.A(_0946_),
    .B(net45),
    .Y(_1317_));
 sg13g2_nor3_1 _2098_ (.A(_1315_),
    .B(_1316_),
    .C(_1317_),
    .Y(_1318_));
 sg13g2_o21ai_1 _2099_ (.B1(_1318_),
    .Y(_1319_),
    .A1(_1301_),
    .A2(_1305_));
 sg13g2_and2_1 _2100_ (.A(_0946_),
    .B(net45),
    .X(_1320_));
 sg13g2_buf_1 _2101_ (.A(_1320_),
    .X(_1321_));
 sg13g2_nand2_1 _2102_ (.Y(_1322_),
    .A(net43),
    .B(_1321_));
 sg13g2_buf_1 _2103_ (.A(\counter[7] ),
    .X(_1323_));
 sg13g2_inv_1 _2104_ (.Y(_1324_),
    .A(_1323_));
 sg13g2_a21o_1 _2105_ (.A2(_1322_),
    .A1(_1319_),
    .B1(_1324_),
    .X(_1325_));
 sg13g2_nor2_1 _2106_ (.A(_1316_),
    .B(_1317_),
    .Y(_1326_));
 sg13g2_o21ai_1 _2107_ (.B1(_1326_),
    .Y(_1327_),
    .A1(_1301_),
    .A2(_1305_));
 sg13g2_buf_2 _2108_ (.A(_1327_),
    .X(_1328_));
 sg13g2_nor2_1 _2109_ (.A(net43),
    .B(_1321_),
    .Y(_1329_));
 sg13g2_nand2_1 _2110_ (.Y(_1330_),
    .A(net69),
    .B(_1323_));
 sg13g2_a21o_1 _2111_ (.A2(_1329_),
    .A1(_1328_),
    .B1(_1330_),
    .X(_1331_));
 sg13g2_and2_1 _2112_ (.A(_1325_),
    .B(_1331_),
    .X(_1332_));
 sg13g2_xor2_1 _2113_ (.B(_1332_),
    .A(_1313_),
    .X(_1333_));
 sg13g2_and2_1 _2114_ (.A(_1289_),
    .B(_1333_),
    .X(_1334_));
 sg13g2_and4_1 _2115_ (.A(\xqo[0] ),
    .B(_1313_),
    .C(_1325_),
    .D(_1331_),
    .X(_1335_));
 sg13g2_nand2b_1 _2116_ (.Y(_1336_),
    .B(_1312_),
    .A_N(_1308_));
 sg13g2_or2_1 _2117_ (.X(_1337_),
    .B(_1305_),
    .A(_1301_));
 sg13g2_a21o_1 _2118_ (.A2(_1337_),
    .A1(_1307_),
    .B1(_1312_),
    .X(_1338_));
 sg13g2_a221oi_1 _2119_ (.B2(_1331_),
    .C1(_1289_),
    .B1(_1325_),
    .A1(_1336_),
    .Y(_1339_),
    .A2(_1338_));
 sg13g2_or2_1 _2120_ (.X(_1340_),
    .B(_1339_),
    .A(_1335_));
 sg13g2_buf_1 _2121_ (.A(_1340_),
    .X(_1341_));
 sg13g2_nor3_1 _2122_ (.A(_1288_),
    .B(_1334_),
    .C(_1341_),
    .Y(_0136_));
 sg13g2_buf_1 _2123_ (.A(_1288_),
    .X(_1342_));
 sg13g2_nand2_1 _2124_ (.Y(_1343_),
    .A(\xqo[8] ),
    .B(\xqo[9] ));
 sg13g2_nor3_1 _2125_ (.A(net44),
    .B(_1321_),
    .C(_1330_),
    .Y(_1344_));
 sg13g2_nor4_1 _2126_ (.A(net47),
    .B(net43),
    .C(net44),
    .D(_1321_),
    .Y(_1345_));
 sg13g2_o21ai_1 _2127_ (.B1(_1328_),
    .Y(_1346_),
    .A1(_1344_),
    .A2(_1345_));
 sg13g2_nor4_1 _2128_ (.A(net69),
    .B(_1315_),
    .C(net44),
    .D(_1321_),
    .Y(_1347_));
 sg13g2_nand2_2 _2129_ (.Y(_1348_),
    .A(_0946_),
    .B(net45));
 sg13g2_inv_1 _2130_ (.Y(_1349_),
    .A(net44));
 sg13g2_nor2_1 _2131_ (.A(_1323_),
    .B(_1349_),
    .Y(_1350_));
 sg13g2_and4_1 _2132_ (.A(net69),
    .B(net43),
    .C(_1348_),
    .D(_1350_),
    .X(_1351_));
 sg13g2_o21ai_1 _2133_ (.B1(_1328_),
    .Y(_1352_),
    .A1(_1347_),
    .A2(_1351_));
 sg13g2_nor2_1 _2134_ (.A(_1323_),
    .B(net44),
    .Y(_1353_));
 sg13g2_nand3_1 _2135_ (.B(net43),
    .C(_1353_),
    .A(net69),
    .Y(_1354_));
 sg13g2_nor2_1 _2136_ (.A(net69),
    .B(net43),
    .Y(_1355_));
 sg13g2_nand3_1 _2137_ (.B(_1348_),
    .C(_1355_),
    .A(net44),
    .Y(_1356_));
 sg13g2_mux2_1 _2138_ (.A0(_1354_),
    .A1(_1356_),
    .S(_1328_),
    .X(_1357_));
 sg13g2_nand2_1 _2139_ (.Y(_1358_),
    .A(_1349_),
    .B(_1355_));
 sg13g2_nor2_1 _2140_ (.A(net47),
    .B(net43),
    .Y(_1359_));
 sg13g2_nand2_1 _2141_ (.Y(_1360_),
    .A(_1359_),
    .B(_1350_));
 sg13g2_a21o_1 _2142_ (.A2(_1360_),
    .A1(_1358_),
    .B1(_1328_),
    .X(_1361_));
 sg13g2_nand4_1 _2143_ (.B(_1352_),
    .C(_1357_),
    .A(_1346_),
    .Y(_1362_),
    .D(_1361_));
 sg13g2_nor2_1 _2144_ (.A(net69),
    .B(_1315_),
    .Y(_1363_));
 sg13g2_nand2_1 _2145_ (.Y(_1364_),
    .A(_1363_),
    .B(_1350_));
 sg13g2_nand4_1 _2146_ (.B(net43),
    .C(_1323_),
    .A(net69),
    .Y(_1365_),
    .D(_1310_));
 sg13g2_a21oi_1 _2147_ (.A1(_1364_),
    .A2(_1365_),
    .Y(_1366_),
    .B1(_1328_));
 sg13g2_nand3_1 _2148_ (.B(_1321_),
    .C(_1355_),
    .A(_1349_),
    .Y(_1367_));
 sg13g2_o21ai_1 _2149_ (.B1(_1367_),
    .Y(_1368_),
    .A1(_1348_),
    .A2(_1354_));
 sg13g2_a21oi_1 _2150_ (.A1(_1360_),
    .A2(_1364_),
    .Y(_1369_),
    .B1(_1348_));
 sg13g2_nor2_1 _2151_ (.A(_1324_),
    .B(_1310_),
    .Y(_1370_));
 sg13g2_o21ai_1 _2152_ (.B1(_1370_),
    .Y(_1371_),
    .A1(_1359_),
    .A2(_1363_));
 sg13g2_o21ai_1 _2153_ (.B1(_1371_),
    .Y(_1372_),
    .A1(_1348_),
    .A2(_1365_));
 sg13g2_or4_1 _2154_ (.A(_1366_),
    .B(_1368_),
    .C(_1369_),
    .D(_1372_),
    .X(_1373_));
 sg13g2_or2_1 _2155_ (.X(_1374_),
    .B(_1373_),
    .A(_1362_));
 sg13g2_a21oi_1 _2156_ (.A1(_1328_),
    .A2(_1329_),
    .Y(_1375_),
    .B1(_1349_));
 sg13g2_nand3_1 _2157_ (.B(_1319_),
    .C(_1322_),
    .A(net47),
    .Y(_1376_));
 sg13g2_mux2_1 _2158_ (.A0(_1353_),
    .A1(_1375_),
    .S(_1376_),
    .X(_1377_));
 sg13g2_nand3_1 _2159_ (.B(_1329_),
    .C(_1353_),
    .A(_1328_),
    .Y(_1378_));
 sg13g2_o21ai_1 _2160_ (.B1(_1378_),
    .Y(_1379_),
    .A1(_1324_),
    .A2(_1349_));
 sg13g2_nor2_1 _2161_ (.A(_1377_),
    .B(_1379_),
    .Y(_1380_));
 sg13g2_buf_1 _2162_ (.A(\xqo[2] ),
    .X(_1381_));
 sg13g2_buf_1 _2163_ (.A(\xqo[3] ),
    .X(_1382_));
 sg13g2_a221oi_1 _2164_ (.B2(_1381_),
    .C1(_1382_),
    .B1(_1380_),
    .A1(_1341_),
    .Y(_1383_),
    .A2(_1374_));
 sg13g2_buf_2 _2165_ (.A(\xqo[1] ),
    .X(_1384_));
 sg13g2_nor2_1 _2166_ (.A(_1384_),
    .B(_1381_),
    .Y(_1385_));
 sg13g2_o21ai_1 _2167_ (.B1(_1385_),
    .Y(_1386_),
    .A1(_1377_),
    .A2(_1379_));
 sg13g2_or2_1 _2168_ (.X(_1387_),
    .B(_1382_),
    .A(_1384_));
 sg13g2_or4_1 _2169_ (.A(_1335_),
    .B(_1339_),
    .C(_1362_),
    .D(_1373_),
    .X(_1388_));
 sg13g2_buf_2 _2170_ (.A(_1388_),
    .X(_1389_));
 sg13g2_a21oi_1 _2171_ (.A1(_1386_),
    .A2(_1387_),
    .Y(_1390_),
    .B1(_1389_));
 sg13g2_or2_1 _2172_ (.X(_1391_),
    .B(_1382_),
    .A(_1381_));
 sg13g2_a21oi_1 _2173_ (.A1(_1391_),
    .A2(_1387_),
    .Y(_1392_),
    .B1(_1380_));
 sg13g2_nor3_1 _2174_ (.A(_1384_),
    .B(_1381_),
    .C(_1382_),
    .Y(_1393_));
 sg13g2_nor4_2 _2175_ (.A(_1383_),
    .B(_1390_),
    .C(_1392_),
    .Y(_1394_),
    .D(_1393_));
 sg13g2_and3_1 _2176_ (.X(_1395_),
    .A(\xqo[5] ),
    .B(\xqo[7] ),
    .C(\xqo[6] ));
 sg13g2_o21ai_1 _2177_ (.B1(_1395_),
    .Y(_1396_),
    .A1(\xqo[4] ),
    .A2(_1394_));
 sg13g2_nor2_1 _2178_ (.A(_1343_),
    .B(_1396_),
    .Y(_1397_));
 sg13g2_xnor2_1 _2179_ (.Y(_1398_),
    .A(\xqo[10] ),
    .B(_1397_));
 sg13g2_nor2_1 _2180_ (.A(net32),
    .B(_1398_),
    .Y(_0137_));
 sg13g2_nand2_1 _2181_ (.Y(_1399_),
    .A(\xqo[9] ),
    .B(\xqo[10] ));
 sg13g2_or2_1 _2182_ (.X(_1400_),
    .B(_1394_),
    .A(\xqo[4] ));
 sg13g2_buf_2 _2183_ (.A(_1400_),
    .X(_1401_));
 sg13g2_nor2b_1 _2184_ (.A(_0003_),
    .B_N(\xqo[5] ),
    .Y(_1402_));
 sg13g2_nand4_1 _2185_ (.B(\xqo[8] ),
    .C(_1401_),
    .A(\xqo[7] ),
    .Y(_1403_),
    .D(_1402_));
 sg13g2_o21ai_1 _2186_ (.B1(\xqo[11] ),
    .Y(_1404_),
    .A1(_1399_),
    .A2(_1403_));
 sg13g2_or3_1 _2187_ (.A(\xqo[11] ),
    .B(_1399_),
    .C(_1403_),
    .X(_1405_));
 sg13g2_a21oi_1 _2188_ (.A1(_1404_),
    .A2(_1405_),
    .Y(_0138_),
    .B1(net32));
 sg13g2_nand2_1 _2189_ (.Y(_1406_),
    .A(_1341_),
    .B(_1374_));
 sg13g2_and2_1 _2190_ (.A(_1406_),
    .B(_1389_),
    .X(_1407_));
 sg13g2_xor2_1 _2191_ (.B(_1407_),
    .A(_1384_),
    .X(_1408_));
 sg13g2_nor2_1 _2192_ (.A(net32),
    .B(_1408_),
    .Y(_0139_));
 sg13g2_mux2_1 _2193_ (.A0(_1389_),
    .A1(_1406_),
    .S(_1384_),
    .X(_1409_));
 sg13g2_xnor2_1 _2194_ (.Y(_1410_),
    .A(_1381_),
    .B(_1380_));
 sg13g2_xnor2_1 _2195_ (.Y(_1411_),
    .A(_1409_),
    .B(_1410_));
 sg13g2_nor2_1 _2196_ (.A(_1342_),
    .B(_1411_),
    .Y(_0140_));
 sg13g2_or2_1 _2197_ (.X(_1412_),
    .B(_1379_),
    .A(_1377_));
 sg13g2_a21oi_1 _2198_ (.A1(_1380_),
    .A2(_1389_),
    .Y(_1413_),
    .B1(_1384_));
 sg13g2_a21oi_1 _2199_ (.A1(_1406_),
    .A2(_1412_),
    .Y(_1414_),
    .B1(_1413_));
 sg13g2_nor2_1 _2200_ (.A(_1406_),
    .B(_1412_),
    .Y(_1415_));
 sg13g2_nor2_1 _2201_ (.A(_1389_),
    .B(_1386_),
    .Y(_1416_));
 sg13g2_a221oi_1 _2202_ (.B2(_1384_),
    .C1(_1416_),
    .B1(_1415_),
    .A1(_1381_),
    .Y(_1417_),
    .A2(_1414_));
 sg13g2_xnor2_1 _2203_ (.Y(_1418_),
    .A(_1382_),
    .B(_1417_));
 sg13g2_nor2_1 _2204_ (.A(net32),
    .B(_1418_),
    .Y(_0141_));
 sg13g2_nand2_1 _2205_ (.Y(_1419_),
    .A(\xqo[4] ),
    .B(_1394_));
 sg13g2_a21oi_1 _2206_ (.A1(_1401_),
    .A2(_1419_),
    .Y(_0142_),
    .B1(net32));
 sg13g2_xnor2_1 _2207_ (.Y(_1420_),
    .A(\xqo[5] ),
    .B(_1401_));
 sg13g2_nor2_1 _2208_ (.A(net32),
    .B(_1420_),
    .Y(_0143_));
 sg13g2_nand2_1 _2209_ (.Y(_1421_),
    .A(\xqo[5] ),
    .B(_1401_));
 sg13g2_xor2_1 _2210_ (.B(_1421_),
    .A(_0003_),
    .X(_1422_));
 sg13g2_nor2b_1 _2211_ (.A(_1342_),
    .B_N(_1422_),
    .Y(_0144_));
 sg13g2_o21ai_1 _2212_ (.B1(\xqo[7] ),
    .Y(_1423_),
    .A1(_0003_),
    .A2(_1421_));
 sg13g2_nand3b_1 _2213_ (.B(_1401_),
    .C(_1402_),
    .Y(_1424_),
    .A_N(\xqo[7] ));
 sg13g2_a21oi_1 _2214_ (.A1(_1423_),
    .A2(_1424_),
    .Y(_0145_),
    .B1(_1288_));
 sg13g2_xor2_1 _2215_ (.B(_1396_),
    .A(\xqo[8] ),
    .X(_1425_));
 sg13g2_nor2_1 _2216_ (.A(net32),
    .B(_1425_),
    .Y(_0146_));
 sg13g2_xor2_1 _2217_ (.B(_1403_),
    .A(\xqo[9] ),
    .X(_1426_));
 sg13g2_nor2_1 _2218_ (.A(net32),
    .B(_1426_),
    .Y(_0147_));
 sg13g2_buf_1 _2219_ (.A(_1287_),
    .X(_1427_));
 sg13g2_nand2b_1 _2220_ (.Y(_1428_),
    .B(\yq[0] ),
    .A_N(net42));
 sg13g2_buf_8 _2221_ (.A(_1287_),
    .X(_1429_));
 sg13g2_buf_1 _2222_ (.A(net41),
    .X(_1430_));
 sg13g2_nor2_1 _2223_ (.A(net72),
    .B(_1290_),
    .Y(_1431_));
 sg13g2_buf_1 _2224_ (.A(_1431_),
    .X(_1432_));
 sg13g2_or2_1 _2225_ (.X(_1433_),
    .B(_1292_),
    .A(net71));
 sg13g2_a21o_1 _2226_ (.A2(_1297_),
    .A1(_0924_),
    .B1(_1295_),
    .X(_1434_));
 sg13g2_and3_1 _2227_ (.X(_1435_),
    .A(_0924_),
    .B(_1295_),
    .C(_1297_));
 sg13g2_a21o_1 _2228_ (.A2(_1434_),
    .A1(_0938_),
    .B1(_1435_),
    .X(_1436_));
 sg13g2_and2_1 _2229_ (.A(net71),
    .B(net46),
    .X(_1437_));
 sg13g2_a221oi_1 _2230_ (.B2(_1436_),
    .C1(_1437_),
    .B1(_1433_),
    .A1(net72),
    .Y(_1438_),
    .A2(_1290_));
 sg13g2_buf_2 _2231_ (.A(_1438_),
    .X(_1439_));
 sg13g2_xnor2_1 _2232_ (.Y(_1440_),
    .A(_0934_),
    .B(_1314_));
 sg13g2_buf_2 _2233_ (.A(_1440_),
    .X(_1441_));
 sg13g2_a221oi_1 _2234_ (.B2(_0928_),
    .C1(_1441_),
    .B1(net45),
    .A1(_0931_),
    .Y(_1442_),
    .A2(net33));
 sg13g2_o21ai_1 _2235_ (.B1(_1442_),
    .Y(_1443_),
    .A1(net21),
    .A2(_1439_));
 sg13g2_nor2_1 _2236_ (.A(_0931_),
    .B(_1302_),
    .Y(_1444_));
 sg13g2_or2_1 _2237_ (.X(_1445_),
    .B(\counter[5] ),
    .A(_0928_));
 sg13g2_buf_1 _2238_ (.A(_1445_),
    .X(_1446_));
 sg13g2_nand3b_1 _2239_ (.B(_1441_),
    .C(_1446_),
    .Y(_1447_),
    .A_N(_1444_));
 sg13g2_or3_1 _2240_ (.A(net21),
    .B(_1439_),
    .C(_1447_),
    .X(_1448_));
 sg13g2_and2_1 _2241_ (.A(_0928_),
    .B(_1309_),
    .X(_1449_));
 sg13g2_nand4_1 _2242_ (.B(net33),
    .C(_1441_),
    .A(net60),
    .Y(_1450_),
    .D(_1446_));
 sg13g2_o21ai_1 _2243_ (.B1(_1450_),
    .Y(_1451_),
    .A1(_1441_),
    .A2(_1446_));
 sg13g2_a221oi_1 _2244_ (.B2(_1444_),
    .C1(_1451_),
    .B1(_1442_),
    .A1(_1449_),
    .Y(_1452_),
    .A2(_1441_));
 sg13g2_nand3_1 _2245_ (.B(_1448_),
    .C(_1452_),
    .A(_1443_),
    .Y(_1453_));
 sg13g2_buf_1 _2246_ (.A(_1453_),
    .X(_1454_));
 sg13g2_inv_2 _2247_ (.Y(_1455_),
    .A(\yqo[0] ));
 sg13g2_nand2_1 _2248_ (.Y(_1456_),
    .A(_0924_),
    .B(_1297_));
 sg13g2_xnor2_1 _2249_ (.Y(_1457_),
    .A(_0938_),
    .B(_1295_));
 sg13g2_xnor2_1 _2250_ (.Y(_1458_),
    .A(_1456_),
    .B(_1457_));
 sg13g2_xnor2_1 _2251_ (.Y(_1459_),
    .A(_1455_),
    .B(_1458_));
 sg13g2_xnor2_1 _2252_ (.Y(_1460_),
    .A(_1454_),
    .B(_1459_));
 sg13g2_nand2_1 _2253_ (.Y(_1461_),
    .A(net31),
    .B(_1460_));
 sg13g2_a21oi_1 _2254_ (.A1(_1428_),
    .A2(_1461_),
    .Y(_0160_),
    .B1(net22));
 sg13g2_nand2b_1 _2255_ (.Y(_1462_),
    .B(\yq[10] ),
    .A_N(net42));
 sg13g2_buf_1 _2256_ (.A(\yqo[10] ),
    .X(_1463_));
 sg13g2_buf_1 _2257_ (.A(\yqo[8] ),
    .X(_1464_));
 sg13g2_buf_8 _2258_ (.A(\yqo[9] ),
    .X(_1465_));
 sg13g2_nor2_1 _2259_ (.A(net64),
    .B(_1465_),
    .Y(_1466_));
 sg13g2_buf_8 _2260_ (.A(\yqo[7] ),
    .X(_1467_));
 sg13g2_xnor2_1 _2261_ (.Y(_1468_),
    .A(net60),
    .B(net33));
 sg13g2_o21ai_1 _2262_ (.B1(_1468_),
    .Y(_1469_),
    .A1(net21),
    .A2(_1439_));
 sg13g2_or3_1 _2263_ (.A(net21),
    .B(_1439_),
    .C(_1468_),
    .X(_1470_));
 sg13g2_buf_1 _2264_ (.A(_1470_),
    .X(_1471_));
 sg13g2_nor2_1 _2265_ (.A(net71),
    .B(net46),
    .Y(_1472_));
 sg13g2_a221oi_1 _2266_ (.B2(_0938_),
    .C1(_1435_),
    .B1(_1434_),
    .A1(net71),
    .Y(_1473_),
    .A2(net46));
 sg13g2_xnor2_1 _2267_ (.Y(_1474_),
    .A(_0926_),
    .B(_1290_));
 sg13g2_o21ai_1 _2268_ (.B1(_1474_),
    .Y(_1475_),
    .A1(_1472_),
    .A2(_1473_));
 sg13g2_or3_1 _2269_ (.A(_1472_),
    .B(_1473_),
    .C(_1474_),
    .X(_1476_));
 sg13g2_and2_1 _2270_ (.A(_1475_),
    .B(_1476_),
    .X(_1477_));
 sg13g2_buf_1 _2271_ (.A(_1477_),
    .X(_1478_));
 sg13g2_and3_1 _2272_ (.X(_1479_),
    .A(_1469_),
    .B(_1471_),
    .C(_1478_));
 sg13g2_a21oi_1 _2273_ (.A1(_1469_),
    .A2(_1471_),
    .Y(_1480_),
    .B1(_1478_));
 sg13g2_a22oi_1 _2274_ (.Y(_1481_),
    .B1(net33),
    .B2(net60),
    .A2(net46),
    .A1(net71));
 sg13g2_inv_1 _2275_ (.Y(_1482_),
    .A(_1481_));
 sg13g2_a221oi_1 _2276_ (.B2(_1436_),
    .C1(_1482_),
    .B1(_1433_),
    .A1(_0926_),
    .Y(_1483_),
    .A2(_1290_));
 sg13g2_nand2_1 _2277_ (.Y(_1484_),
    .A(_0932_),
    .B(_1306_));
 sg13g2_a21o_1 _2278_ (.A2(_1484_),
    .A1(net21),
    .B1(_1444_),
    .X(_1485_));
 sg13g2_xnor2_1 _2279_ (.Y(_1486_),
    .A(net45),
    .B(\yqo[4] ));
 sg13g2_xnor2_1 _2280_ (.Y(_1487_),
    .A(_0929_),
    .B(_1486_));
 sg13g2_or3_1 _2281_ (.A(_1483_),
    .B(_1485_),
    .C(_1487_),
    .X(_1488_));
 sg13g2_buf_1 _2282_ (.A(_1488_),
    .X(_0186_));
 sg13g2_o21ai_1 _2283_ (.B1(_1487_),
    .Y(_0187_),
    .A1(_1483_),
    .A2(_1485_));
 sg13g2_nand2_2 _2284_ (.Y(_0188_),
    .A(_0186_),
    .B(_0187_));
 sg13g2_mux2_1 _2285_ (.A0(_1479_),
    .A1(_1480_),
    .S(_0188_),
    .X(_0189_));
 sg13g2_buf_2 _2286_ (.A(\yqo[2] ),
    .X(_0190_));
 sg13g2_inv_1 _2287_ (.Y(_0191_),
    .A(_0190_));
 sg13g2_buf_1 _2288_ (.A(\yqo[3] ),
    .X(_0192_));
 sg13g2_nor2_1 _2289_ (.A(_0191_),
    .B(net63),
    .Y(_0193_));
 sg13g2_and2_1 _2290_ (.A(_0190_),
    .B(net63),
    .X(_0194_));
 sg13g2_and3_1 _2291_ (.X(_0195_),
    .A(_1478_),
    .B(_0186_),
    .C(_0187_));
 sg13g2_a21oi_1 _2292_ (.A1(_0186_),
    .A2(_0187_),
    .Y(_0196_),
    .B1(_1478_));
 sg13g2_mux2_1 _2293_ (.A0(_0195_),
    .A1(_0196_),
    .S(net15),
    .X(_0197_));
 sg13g2_a22oi_1 _2294_ (.Y(_0198_),
    .B1(_0194_),
    .B2(_0197_),
    .A2(_0193_),
    .A1(_0189_));
 sg13g2_nand2_1 _2295_ (.Y(_0199_),
    .A(_1469_),
    .B(_1471_));
 sg13g2_nand2_1 _2296_ (.Y(_0200_),
    .A(_0199_),
    .B(_0188_));
 sg13g2_or2_1 _2297_ (.X(_0201_),
    .B(_0188_),
    .A(_0199_));
 sg13g2_and3_1 _2298_ (.X(_0202_),
    .A(_1443_),
    .B(_1448_),
    .C(_1452_));
 sg13g2_buf_1 _2299_ (.A(_0202_),
    .X(_0203_));
 sg13g2_buf_8 _2300_ (.A(_0203_),
    .X(_0204_));
 sg13g2_xnor2_1 _2301_ (.Y(_0205_),
    .A(net63),
    .B(net13));
 sg13g2_mux2_1 _2302_ (.A0(_0200_),
    .A1(_0201_),
    .S(_0205_),
    .X(_0206_));
 sg13g2_buf_8 _2303_ (.A(\yqo[1] ),
    .X(_0207_));
 sg13g2_xor2_1 _2304_ (.B(net46),
    .A(_0940_),
    .X(_0208_));
 sg13g2_xnor2_1 _2305_ (.Y(_0209_),
    .A(_1436_),
    .B(_0208_));
 sg13g2_xnor2_1 _2306_ (.Y(_0210_),
    .A(_0207_),
    .B(_0209_));
 sg13g2_nor2b_1 _2307_ (.A(_0207_),
    .B_N(_0209_),
    .Y(_0211_));
 sg13g2_or4_1 _2308_ (.A(_1455_),
    .B(_1458_),
    .C(_0210_),
    .D(_0211_),
    .X(_0212_));
 sg13g2_a21o_1 _2309_ (.A2(_1476_),
    .A1(_1475_),
    .B1(_0191_),
    .X(_0213_));
 sg13g2_buf_1 _2310_ (.A(_0213_),
    .X(_0214_));
 sg13g2_nand3_1 _2311_ (.B(_1475_),
    .C(_1476_),
    .A(_0191_),
    .Y(_0215_));
 sg13g2_a21o_1 _2312_ (.A2(_0215_),
    .A1(_0214_),
    .B1(_0211_),
    .X(_0216_));
 sg13g2_a21oi_1 _2313_ (.A1(_0212_),
    .A2(_0216_),
    .Y(_0217_),
    .B1(net15));
 sg13g2_nand2_1 _2314_ (.Y(_0218_),
    .A(_0214_),
    .B(_0215_));
 sg13g2_nor3_1 _2315_ (.A(_1455_),
    .B(_1458_),
    .C(_0210_),
    .Y(_0219_));
 sg13g2_and3_1 _2316_ (.X(_0220_),
    .A(_0203_),
    .B(_0218_),
    .C(_0219_));
 sg13g2_and2_1 _2317_ (.A(\yqo[0] ),
    .B(_1458_),
    .X(_0221_));
 sg13g2_nand3_1 _2318_ (.B(_0221_),
    .C(_0209_),
    .A(_0207_),
    .Y(_0222_));
 sg13g2_nand4_1 _2319_ (.B(_0214_),
    .C(_0215_),
    .A(_0221_),
    .Y(_0223_),
    .D(_0210_));
 sg13g2_a21oi_1 _2320_ (.A1(_0222_),
    .A2(_0223_),
    .Y(_0224_),
    .B1(net13));
 sg13g2_nor2_1 _2321_ (.A(_0207_),
    .B(_0209_),
    .Y(_0225_));
 sg13g2_nor3_1 _2322_ (.A(net13),
    .B(_0218_),
    .C(_0225_),
    .Y(_0226_));
 sg13g2_nor4_2 _2323_ (.A(_0217_),
    .B(_0220_),
    .C(_0224_),
    .Y(_0227_),
    .D(_0226_));
 sg13g2_xor2_1 _2324_ (.B(_1306_),
    .A(_0932_),
    .X(_0228_));
 sg13g2_and2_1 _2325_ (.A(_0192_),
    .B(_0228_),
    .X(_0229_));
 sg13g2_o21ai_1 _2326_ (.B1(_0229_),
    .Y(_0230_),
    .A1(net21),
    .A2(_1439_));
 sg13g2_or4_1 _2327_ (.A(net63),
    .B(net21),
    .C(_1439_),
    .D(_1468_),
    .X(_0231_));
 sg13g2_nor2_1 _2328_ (.A(_0192_),
    .B(_0228_),
    .Y(_0232_));
 sg13g2_o21ai_1 _2329_ (.B1(_0232_),
    .Y(_0233_),
    .A1(net21),
    .A2(_1439_));
 sg13g2_nand2_1 _2330_ (.Y(_0234_),
    .A(\yqo[3] ),
    .B(_1468_));
 sg13g2_or3_1 _2331_ (.A(_1432_),
    .B(_1439_),
    .C(_0234_),
    .X(_0235_));
 sg13g2_nand4_1 _2332_ (.B(_0231_),
    .C(_0233_),
    .A(_0230_),
    .Y(_0236_),
    .D(_0235_));
 sg13g2_buf_2 _2333_ (.A(_0236_),
    .X(_0237_));
 sg13g2_and3_1 _2334_ (.X(_0238_),
    .A(net13),
    .B(_1478_),
    .C(_0237_));
 sg13g2_nor3_1 _2335_ (.A(net13),
    .B(_1478_),
    .C(_0237_),
    .Y(_0239_));
 sg13g2_o21ai_1 _2336_ (.B1(_0190_),
    .Y(_0240_),
    .A1(_0238_),
    .A2(_0239_));
 sg13g2_a22oi_1 _2337_ (.Y(_0241_),
    .B1(_0227_),
    .B2(_0240_),
    .A2(_0206_),
    .A1(_0198_));
 sg13g2_buf_2 _2338_ (.A(_0241_),
    .X(_0242_));
 sg13g2_nand2_1 _2339_ (.Y(_0243_),
    .A(_0929_),
    .B(net45));
 sg13g2_nor2_1 _2340_ (.A(_1483_),
    .B(_1485_),
    .Y(_0244_));
 sg13g2_mux2_1 _2341_ (.A0(_1446_),
    .A1(_0243_),
    .S(_0244_),
    .X(_0245_));
 sg13g2_xnor2_1 _2342_ (.Y(_0246_),
    .A(_1441_),
    .B(_0245_));
 sg13g2_nand2_2 _2343_ (.Y(_0247_),
    .A(\yqo[4] ),
    .B(_0246_));
 sg13g2_xnor2_1 _2344_ (.Y(_0248_),
    .A(net15),
    .B(_0199_));
 sg13g2_xnor2_1 _2345_ (.Y(_0249_),
    .A(net13),
    .B(_0188_));
 sg13g2_o21ai_1 _2346_ (.B1(_0249_),
    .Y(_0250_),
    .A1(net63),
    .A2(_0248_));
 sg13g2_nand2_1 _2347_ (.Y(_0251_),
    .A(_0247_),
    .B(_0250_));
 sg13g2_buf_2 _2348_ (.A(\yqo[5] ),
    .X(_0252_));
 sg13g2_buf_8 _2349_ (.A(\yqo[6] ),
    .X(_0253_));
 sg13g2_or2_1 _2350_ (.X(_0254_),
    .B(_0253_),
    .A(_0252_));
 sg13g2_nor4_2 _2351_ (.A(_1467_),
    .B(_0242_),
    .C(_0251_),
    .Y(_0255_),
    .D(_0254_));
 sg13g2_and2_1 _2352_ (.A(net64),
    .B(_1465_),
    .X(_0256_));
 sg13g2_inv_1 _2353_ (.Y(_0257_),
    .A(_0247_));
 sg13g2_and3_1 _2354_ (.X(_0258_),
    .A(_0252_),
    .B(_0253_),
    .C(_1467_));
 sg13g2_and3_1 _2355_ (.X(_0259_),
    .A(_0257_),
    .B(_0242_),
    .C(_0258_));
 sg13g2_buf_1 _2356_ (.A(_0259_),
    .X(_0260_));
 sg13g2_a22oi_1 _2357_ (.Y(_0261_),
    .B1(_0256_),
    .B2(_0260_),
    .A2(_0255_),
    .A1(_1466_));
 sg13g2_xnor2_1 _2358_ (.Y(_0262_),
    .A(_1463_),
    .B(_0261_));
 sg13g2_nand2_1 _2359_ (.Y(_0263_),
    .A(net31),
    .B(_0262_));
 sg13g2_a21oi_1 _2360_ (.A1(_1462_),
    .A2(_0263_),
    .Y(_0161_),
    .B1(net22));
 sg13g2_nand2b_1 _2361_ (.Y(_0264_),
    .B(\yq[11] ),
    .A_N(net42));
 sg13g2_nor3_1 _2362_ (.A(net64),
    .B(_1465_),
    .C(_1463_),
    .Y(_0265_));
 sg13g2_nand4_1 _2363_ (.B(_1465_),
    .C(_1463_),
    .A(net64),
    .Y(_0266_),
    .D(_0258_));
 sg13g2_nor2_1 _2364_ (.A(_0247_),
    .B(_0266_),
    .Y(_0267_));
 sg13g2_nand2b_1 _2365_ (.Y(_0268_),
    .B(_0250_),
    .A_N(_0242_));
 sg13g2_a22oi_1 _2366_ (.Y(_0269_),
    .B1(_0267_),
    .B2(_0268_),
    .A2(_0265_),
    .A1(_0255_));
 sg13g2_xnor2_1 _2367_ (.Y(_0270_),
    .A(\yqo[11] ),
    .B(_0269_));
 sg13g2_nand2_1 _2368_ (.Y(_0271_),
    .A(net31),
    .B(_0270_));
 sg13g2_a21oi_1 _2369_ (.A1(_0264_),
    .A2(_0271_),
    .Y(_0162_),
    .B1(net22));
 sg13g2_nand2b_1 _2370_ (.Y(_0272_),
    .B(\yq[12] ),
    .A_N(net42));
 sg13g2_nor4_1 _2371_ (.A(net64),
    .B(_1465_),
    .C(_1463_),
    .D(\yqo[11] ),
    .Y(_0273_));
 sg13g2_and4_1 _2372_ (.A(_0252_),
    .B(_1467_),
    .C(_1465_),
    .D(_1463_),
    .X(_0274_));
 sg13g2_nand4_1 _2373_ (.B(_1464_),
    .C(\yqo[11] ),
    .A(_0253_),
    .Y(_0275_),
    .D(_0274_));
 sg13g2_nor2_1 _2374_ (.A(_0247_),
    .B(_0275_),
    .Y(_0276_));
 sg13g2_a22oi_1 _2375_ (.Y(_0277_),
    .B1(_0276_),
    .B2(_0268_),
    .A2(_0273_),
    .A1(_0255_));
 sg13g2_xnor2_1 _2376_ (.Y(_0278_),
    .A(\yqo[12] ),
    .B(_0277_));
 sg13g2_nand2_1 _2377_ (.Y(_0279_),
    .A(net31),
    .B(_0278_));
 sg13g2_a21oi_1 _2378_ (.A1(_0272_),
    .A2(_0279_),
    .Y(_0163_),
    .B1(net22));
 sg13g2_nand2b_1 _2379_ (.Y(_0280_),
    .B(\yq[1] ),
    .A_N(net41));
 sg13g2_a21o_1 _2380_ (.A2(net13),
    .A1(_1455_),
    .B1(_0221_),
    .X(_0281_));
 sg13g2_xor2_1 _2381_ (.B(_0281_),
    .A(_0210_),
    .X(_0282_));
 sg13g2_nand2_1 _2382_ (.Y(_0283_),
    .A(net31),
    .B(_0282_));
 sg13g2_a21oi_1 _2383_ (.A1(_0280_),
    .A2(_0283_),
    .Y(_0164_),
    .B1(net22));
 sg13g2_nand2b_1 _2384_ (.Y(_0284_),
    .B(\yq[2] ),
    .A_N(_1429_));
 sg13g2_and3_1 _2385_ (.X(_0285_),
    .A(net15),
    .B(_1458_),
    .C(_0210_));
 sg13g2_nor3_1 _2386_ (.A(net15),
    .B(_1458_),
    .C(_0210_),
    .Y(_0286_));
 sg13g2_o21ai_1 _2387_ (.B1(\yqo[0] ),
    .Y(_0287_),
    .A1(_0285_),
    .A2(_0286_));
 sg13g2_a21oi_1 _2388_ (.A1(_0207_),
    .A2(_0204_),
    .Y(_0288_),
    .B1(_0225_));
 sg13g2_xnor2_1 _2389_ (.Y(_0289_),
    .A(_0218_),
    .B(_0288_));
 sg13g2_xnor2_1 _2390_ (.Y(_0290_),
    .A(_0287_),
    .B(_0289_));
 sg13g2_nand2_1 _2391_ (.Y(_0291_),
    .A(_1430_),
    .B(_0290_));
 sg13g2_a21oi_1 _2392_ (.A1(_0284_),
    .A2(_0291_),
    .Y(_0165_),
    .B1(_1243_));
 sg13g2_nand2b_1 _2393_ (.Y(_0292_),
    .B(\yq[3] ),
    .A_N(_1429_));
 sg13g2_o21ai_1 _2394_ (.B1(_0214_),
    .Y(_0293_),
    .A1(_0190_),
    .A2(net15));
 sg13g2_xnor2_1 _2395_ (.Y(_0294_),
    .A(_0237_),
    .B(_0293_));
 sg13g2_xnor2_1 _2396_ (.Y(_0295_),
    .A(_0227_),
    .B(_0294_));
 sg13g2_nand2_1 _2397_ (.Y(_0296_),
    .A(_1430_),
    .B(_0295_));
 sg13g2_a21oi_1 _2398_ (.A1(_0292_),
    .A2(_0296_),
    .Y(_0166_),
    .B1(_1243_));
 sg13g2_nand2b_1 _2399_ (.Y(_0297_),
    .B(\yq[4] ),
    .A_N(net41));
 sg13g2_buf_8 _2400_ (.A(_1287_),
    .X(_0298_));
 sg13g2_xnor2_1 _2401_ (.Y(_0299_),
    .A(net15),
    .B(_0237_));
 sg13g2_nand2b_1 _2402_ (.Y(_0300_),
    .B(_0227_),
    .A_N(_0237_));
 sg13g2_nand2_1 _2403_ (.Y(_0301_),
    .A(_0190_),
    .B(_1478_));
 sg13g2_nor2_1 _2404_ (.A(net15),
    .B(_0301_),
    .Y(_0302_));
 sg13g2_nor2_1 _2405_ (.A(_0204_),
    .B(_0214_),
    .Y(_0303_));
 sg13g2_nand2_1 _2406_ (.Y(_0304_),
    .A(_0227_),
    .B(_0237_));
 sg13g2_a22oi_1 _2407_ (.Y(_0305_),
    .B1(_0303_),
    .B2(_0304_),
    .A2(_0302_),
    .A1(_0300_));
 sg13g2_o21ai_1 _2408_ (.B1(_0305_),
    .Y(_0306_),
    .A1(_0227_),
    .A2(_0299_));
 sg13g2_nor2_1 _2409_ (.A(net63),
    .B(_0199_),
    .Y(_0307_));
 sg13g2_a21oi_1 _2410_ (.A1(net63),
    .A2(net13),
    .Y(_0308_),
    .B1(_0307_));
 sg13g2_xor2_1 _2411_ (.B(_0188_),
    .A(_0308_),
    .X(_0309_));
 sg13g2_xnor2_1 _2412_ (.Y(_0310_),
    .A(_0306_),
    .B(_0309_));
 sg13g2_nand2_1 _2413_ (.Y(_0311_),
    .A(_0298_),
    .B(_0310_));
 sg13g2_buf_8 _2414_ (.A(_1242_),
    .X(_0312_));
 sg13g2_buf_1 _2415_ (.A(net20),
    .X(_0313_));
 sg13g2_a21oi_1 _2416_ (.A1(_0297_),
    .A2(_0311_),
    .Y(_0167_),
    .B1(_0313_));
 sg13g2_nand2b_1 _2417_ (.Y(_0314_),
    .B(\yq[5] ),
    .A_N(net41));
 sg13g2_xnor2_1 _2418_ (.Y(_0315_),
    .A(_0252_),
    .B(_0247_));
 sg13g2_xnor2_1 _2419_ (.Y(_0316_),
    .A(_0268_),
    .B(_0315_));
 sg13g2_nand2_1 _2420_ (.Y(_0317_),
    .A(_0298_),
    .B(_0316_));
 sg13g2_a21oi_1 _2421_ (.A1(_0314_),
    .A2(_0317_),
    .Y(_0168_),
    .B1(net18));
 sg13g2_buf_1 _2422_ (.A(\yq[6] ),
    .X(_0318_));
 sg13g2_nand2b_1 _2423_ (.Y(_0319_),
    .B(_0318_),
    .A_N(net41));
 sg13g2_or2_1 _2424_ (.X(_0320_),
    .B(_0251_),
    .A(_0242_));
 sg13g2_nand3_1 _2425_ (.B(_0257_),
    .C(_0242_),
    .A(_0252_),
    .Y(_0321_));
 sg13g2_o21ai_1 _2426_ (.B1(_0321_),
    .Y(_0322_),
    .A1(_0252_),
    .A2(_0320_));
 sg13g2_xor2_1 _2427_ (.B(_0322_),
    .A(_0253_),
    .X(_0323_));
 sg13g2_nand2_1 _2428_ (.Y(_0324_),
    .A(net40),
    .B(_0323_));
 sg13g2_a21oi_1 _2429_ (.A1(_0319_),
    .A2(_0324_),
    .Y(_0169_),
    .B1(net18));
 sg13g2_buf_2 _2430_ (.A(\yq[7] ),
    .X(_0325_));
 sg13g2_nand2b_1 _2431_ (.Y(_0326_),
    .B(_0325_),
    .A_N(net41));
 sg13g2_nand4_1 _2432_ (.B(_0253_),
    .C(_0257_),
    .A(_0252_),
    .Y(_0327_),
    .D(_0242_));
 sg13g2_o21ai_1 _2433_ (.B1(_0327_),
    .Y(_0328_),
    .A1(_0320_),
    .A2(_0254_));
 sg13g2_xor2_1 _2434_ (.B(_0328_),
    .A(_1467_),
    .X(_0329_));
 sg13g2_nand2_1 _2435_ (.Y(_0330_),
    .A(net40),
    .B(_0329_));
 sg13g2_a21oi_1 _2436_ (.A1(_0326_),
    .A2(_0330_),
    .Y(_0170_),
    .B1(net18));
 sg13g2_buf_2 _2437_ (.A(\yq[8] ),
    .X(_0331_));
 sg13g2_nand2b_1 _2438_ (.Y(_0332_),
    .B(_0331_),
    .A_N(net41));
 sg13g2_nor2_1 _2439_ (.A(_0255_),
    .B(_0260_),
    .Y(_0333_));
 sg13g2_xnor2_1 _2440_ (.Y(_0334_),
    .A(net64),
    .B(_0333_));
 sg13g2_nand2_1 _2441_ (.Y(_0335_),
    .A(net40),
    .B(_0334_));
 sg13g2_a21oi_1 _2442_ (.A1(_0332_),
    .A2(_0335_),
    .Y(_0171_),
    .B1(net18));
 sg13g2_buf_8 _2443_ (.A(\yq[9] ),
    .X(_0336_));
 sg13g2_nand2b_1 _2444_ (.Y(_0337_),
    .B(_0336_),
    .A_N(net41));
 sg13g2_mux2_1 _2445_ (.A0(_0255_),
    .A1(_0260_),
    .S(net64),
    .X(_0338_));
 sg13g2_xor2_1 _2446_ (.B(_0338_),
    .A(_1465_),
    .X(_0339_));
 sg13g2_nand2_1 _2447_ (.Y(_0340_),
    .A(net40),
    .B(_0339_));
 sg13g2_a21oi_1 _2448_ (.A1(_0337_),
    .A2(_0340_),
    .Y(_0172_),
    .B1(net18));
 sg13g2_nand2_1 _2449_ (.Y(_0341_),
    .A(net42),
    .B(\yqo[0] ));
 sg13g2_a21oi_1 _2450_ (.A1(_1428_),
    .A2(_0341_),
    .Y(_0173_),
    .B1(_0313_));
 sg13g2_nand2_1 _2451_ (.Y(_0342_),
    .A(net31),
    .B(_1463_));
 sg13g2_a21oi_1 _2452_ (.A1(_1462_),
    .A2(_0342_),
    .Y(_0174_),
    .B1(net18));
 sg13g2_nand2_1 _2453_ (.Y(_0343_),
    .A(net31),
    .B(\yqo[11] ));
 sg13g2_a21oi_1 _2454_ (.A1(_0264_),
    .A2(_0343_),
    .Y(_0175_),
    .B1(net18));
 sg13g2_nand2_1 _2455_ (.Y(_0344_),
    .A(net31),
    .B(\yqo[12] ));
 sg13g2_a21oi_1 _2456_ (.A1(_0272_),
    .A2(_0344_),
    .Y(_0176_),
    .B1(net18));
 sg13g2_nand2_1 _2457_ (.Y(_0345_),
    .A(net42),
    .B(_0207_));
 sg13g2_a21oi_1 _2458_ (.A1(_0280_),
    .A2(_0345_),
    .Y(_0177_),
    .B1(net20));
 sg13g2_nand2_1 _2459_ (.Y(_0346_),
    .A(_1427_),
    .B(_0190_));
 sg13g2_a21oi_1 _2460_ (.A1(_0284_),
    .A2(_0346_),
    .Y(_0178_),
    .B1(net20));
 sg13g2_nand2_1 _2461_ (.Y(_0347_),
    .A(_1427_),
    .B(net63));
 sg13g2_a21oi_1 _2462_ (.A1(_0292_),
    .A2(_0347_),
    .Y(_0179_),
    .B1(_0312_));
 sg13g2_nand2_1 _2463_ (.Y(_0348_),
    .A(net42),
    .B(\yqo[4] ));
 sg13g2_a21oi_1 _2464_ (.A1(_0297_),
    .A2(_0348_),
    .Y(_0180_),
    .B1(_0312_));
 sg13g2_nand2_1 _2465_ (.Y(_0349_),
    .A(net42),
    .B(_0252_));
 sg13g2_a21oi_1 _2466_ (.A1(_0314_),
    .A2(_0349_),
    .Y(_0181_),
    .B1(net20));
 sg13g2_nand2_1 _2467_ (.Y(_0350_),
    .A(net40),
    .B(_0253_));
 sg13g2_a21oi_1 _2468_ (.A1(_0319_),
    .A2(_0350_),
    .Y(_0182_),
    .B1(net20));
 sg13g2_nand2_1 _2469_ (.Y(_0351_),
    .A(net40),
    .B(_1467_));
 sg13g2_a21oi_1 _2470_ (.A1(_0326_),
    .A2(_0351_),
    .Y(_0183_),
    .B1(net20));
 sg13g2_nand2_1 _2471_ (.Y(_0352_),
    .A(net40),
    .B(net64));
 sg13g2_a21oi_1 _2472_ (.A1(_0332_),
    .A2(_0352_),
    .Y(_0184_),
    .B1(net20));
 sg13g2_nand2_1 _2473_ (.Y(_0353_),
    .A(net40),
    .B(_1465_));
 sg13g2_a21oi_1 _2474_ (.A1(_0337_),
    .A2(_0353_),
    .Y(_0185_),
    .B1(net20));
 sg13g2_inv_1 _2475_ (.Y(_0354_),
    .A(\Voice1.pulsewidth[8] ));
 sg13g2_nor2_1 _2476_ (.A(_1127_),
    .B(_0354_),
    .Y(_0355_));
 sg13g2_inv_1 _2477_ (.Y(_0356_),
    .A(\Voice1.pulsewidth[5] ));
 sg13g2_inv_1 _2478_ (.Y(_0357_),
    .A(\Voice1.pulsewidth[4] ));
 sg13g2_inv_1 _2479_ (.Y(_0358_),
    .A(\Voice1.pulsewidth[3] ));
 sg13g2_inv_1 _2480_ (.Y(_0359_),
    .A(\Voice1.pulsewidth[2] ));
 sg13g2_buf_1 _2481_ (.A(\Voice1.pulsewidth[1] ),
    .X(_0360_));
 sg13g2_inv_1 _2482_ (.Y(_0361_),
    .A(_0360_));
 sg13g2_nand2b_1 _2483_ (.Y(_0362_),
    .B(\Voice1.pulsewidth[0] ),
    .A_N(_1084_));
 sg13g2_nand2_1 _2484_ (.Y(_0363_),
    .A(_0361_),
    .B(_0362_));
 sg13g2_o21ai_1 _2485_ (.B1(\Voice1.accumulator[13] ),
    .Y(_0364_),
    .A1(_0361_),
    .A2(_0362_));
 sg13g2_a22oi_1 _2486_ (.Y(_0365_),
    .B1(_0363_),
    .B2(_0364_),
    .A2(\Voice1.pulsewidth[2] ),
    .A1(_1113_));
 sg13g2_a221oi_1 _2487_ (.B2(_0359_),
    .C1(_0365_),
    .B1(_1104_),
    .A1(_1107_),
    .Y(_0366_),
    .A2(_0358_));
 sg13g2_a221oi_1 _2488_ (.B2(\Voice1.pulsewidth[3] ),
    .C1(_0366_),
    .B1(_1112_),
    .A1(_1111_),
    .Y(_0367_),
    .A2(\Voice1.pulsewidth[4] ));
 sg13g2_a21o_1 _2489_ (.A2(_0357_),
    .A1(\Voice1.accumulator[16] ),
    .B1(_0367_),
    .X(_0368_));
 sg13g2_o21ai_1 _2490_ (.B1(_0368_),
    .Y(_0369_),
    .A1(\Voice1.accumulator[17] ),
    .A2(_0356_));
 sg13g2_buf_1 _2491_ (.A(\Voice1.pulsewidth[6] ),
    .X(_0370_));
 sg13g2_inv_1 _2492_ (.Y(_0371_),
    .A(_0370_));
 sg13g2_a22oi_1 _2493_ (.Y(_0372_),
    .B1(\Voice1.accumulator[17] ),
    .B2(_0356_),
    .A2(_0371_),
    .A1(_1119_));
 sg13g2_nor2_1 _2494_ (.A(_1119_),
    .B(_0371_),
    .Y(_0373_));
 sg13g2_a221oi_1 _2495_ (.B2(_0372_),
    .C1(_0373_),
    .B1(_0369_),
    .A1(_1128_),
    .Y(_0374_),
    .A2(net50));
 sg13g2_a221oi_1 _2496_ (.B2(_0996_),
    .C1(_0374_),
    .B1(\Voice1.accumulator[19] ),
    .A1(_1127_),
    .Y(_0375_),
    .A2(_0354_));
 sg13g2_or4_1 _2497_ (.A(_1138_),
    .B(_0005_),
    .C(_0355_),
    .D(_0375_),
    .X(_0376_));
 sg13g2_nand2_1 _2498_ (.Y(_0377_),
    .A(net52),
    .B(_0376_));
 sg13g2_o21ai_1 _2499_ (.B1(_1135_),
    .Y(_0378_),
    .A1(net52),
    .A2(_0376_));
 sg13g2_a21oi_1 _2500_ (.A1(_0377_),
    .A2(_0378_),
    .Y(_0379_),
    .B1(\Voice1.accumulator[23] ));
 sg13g2_o21ai_1 _2501_ (.B1(net65),
    .Y(_0380_),
    .A1(\Voice1.en ),
    .A2(\Voice1.pulse ));
 sg13g2_a21oi_1 _2502_ (.A1(\Voice1.en ),
    .A2(_0379_),
    .Y(_0049_),
    .B1(_0380_));
 sg13g2_buf_1 _2503_ (.A(\VAL[8] ),
    .X(_0381_));
 sg13g2_xnor2_1 _2504_ (.Y(_0382_),
    .A(net57),
    .B(_0381_));
 sg13g2_nor2_1 _2505_ (.A(net34),
    .B(_0382_),
    .Y(_0050_));
 sg13g2_nand2_1 _2506_ (.Y(_0383_),
    .A(net57),
    .B(_0381_));
 sg13g2_buf_1 _2507_ (.A(\VAL[9] ),
    .X(_0384_));
 sg13g2_xnor2_1 _2508_ (.Y(_0385_),
    .A(net62),
    .B(_0384_));
 sg13g2_xnor2_1 _2509_ (.Y(_0386_),
    .A(_0383_),
    .B(_0385_));
 sg13g2_nor2_1 _2510_ (.A(net34),
    .B(_0386_),
    .Y(_0051_));
 sg13g2_inv_1 _2511_ (.Y(_0387_),
    .A(net72));
 sg13g2_a21oi_1 _2512_ (.A1(net57),
    .A2(_0381_),
    .Y(_0388_),
    .B1(_0384_));
 sg13g2_nand3_1 _2513_ (.B(_0384_),
    .C(_0381_),
    .A(net57),
    .Y(_0389_));
 sg13g2_o21ai_1 _2514_ (.B1(_0389_),
    .Y(_0390_),
    .A1(_0387_),
    .A2(_0388_));
 sg13g2_buf_1 _2515_ (.A(\VAL[10] ),
    .X(_0391_));
 sg13g2_xor2_1 _2516_ (.B(_0391_),
    .A(net35),
    .X(_0392_));
 sg13g2_xnor2_1 _2517_ (.Y(_0393_),
    .A(_0390_),
    .B(_0392_));
 sg13g2_nor2_1 _2518_ (.A(net34),
    .B(_0393_),
    .Y(_0052_));
 sg13g2_nor2_1 _2519_ (.A(_0391_),
    .B(_0390_),
    .Y(_0394_));
 sg13g2_a21oi_1 _2520_ (.A1(_0391_),
    .A2(_0390_),
    .Y(_0395_),
    .B1(net60));
 sg13g2_nor2_1 _2521_ (.A(_0394_),
    .B(_0395_),
    .Y(_0396_));
 sg13g2_buf_1 _2522_ (.A(\VAL[11] ),
    .X(_0397_));
 sg13g2_xor2_1 _2523_ (.B(_0397_),
    .A(_0930_),
    .X(_0398_));
 sg13g2_xnor2_1 _2524_ (.Y(_0399_),
    .A(_0396_),
    .B(_0398_));
 sg13g2_nor2_1 _2525_ (.A(net34),
    .B(_0399_),
    .Y(_0053_));
 sg13g2_a21o_1 _2526_ (.A2(_0396_),
    .A1(_0397_),
    .B1(net61),
    .X(_0400_));
 sg13g2_o21ai_1 _2527_ (.B1(_0400_),
    .Y(_0401_),
    .A1(_0397_),
    .A2(_0396_));
 sg13g2_xnor2_1 _2528_ (.Y(_0402_),
    .A(net59),
    .B(\VAL[12] ));
 sg13g2_xnor2_1 _2529_ (.Y(_0403_),
    .A(_0401_),
    .B(_0402_));
 sg13g2_nor2_1 _2530_ (.A(_1257_),
    .B(_0403_),
    .Y(_0054_));
 sg13g2_inv_1 _2531_ (.Y(_0404_),
    .A(\VAL[12] ));
 sg13g2_inv_1 _2532_ (.Y(_0405_),
    .A(_0401_));
 sg13g2_a21oi_1 _2533_ (.A1(\VAL[12] ),
    .A2(_0405_),
    .Y(_0406_),
    .B1(net59));
 sg13g2_a21oi_1 _2534_ (.A1(_0404_),
    .A2(_0401_),
    .Y(_0407_),
    .B1(_0406_));
 sg13g2_nand2b_1 _2535_ (.Y(_0408_),
    .B(_0407_),
    .A_N(_0012_));
 sg13g2_nand2b_1 _2536_ (.Y(_0409_),
    .B(_0012_),
    .A_N(_0407_));
 sg13g2_and3_1 _2537_ (.X(_0055_),
    .A(_1091_),
    .B(_0408_),
    .C(_0409_));
 sg13g2_buf_1 _2538_ (.A(net48),
    .X(_0410_));
 sg13g2_xnor2_1 _2539_ (.Y(_0411_),
    .A(_0009_),
    .B(_0408_));
 sg13g2_nor2_1 _2540_ (.A(net30),
    .B(_0411_),
    .Y(_0056_));
 sg13g2_nand3_1 _2541_ (.B(\VAL[14] ),
    .C(_0407_),
    .A(\VAL[13] ),
    .Y(_0412_));
 sg13g2_xnor2_1 _2542_ (.Y(_0413_),
    .A(_0010_),
    .B(_0412_));
 sg13g2_nor2_1 _2543_ (.A(net30),
    .B(_0413_),
    .Y(_0057_));
 sg13g2_buf_1 _2544_ (.A(net65),
    .X(_0414_));
 sg13g2_and2_1 _2545_ (.A(_0414_),
    .B(_0015_),
    .X(_0058_));
 sg13g2_xnor2_1 _2546_ (.Y(_0415_),
    .A(_1295_),
    .B(_1297_));
 sg13g2_nor2_1 _2547_ (.A(_0410_),
    .B(_0415_),
    .Y(_0059_));
 sg13g2_nand2_1 _2548_ (.Y(_0416_),
    .A(_1295_),
    .B(_1297_));
 sg13g2_xor2_1 _2549_ (.B(_0416_),
    .A(_1292_),
    .X(_0417_));
 sg13g2_nor2_1 _2550_ (.A(net30),
    .B(_0417_),
    .Y(_0060_));
 sg13g2_nand3_1 _2551_ (.B(_1297_),
    .C(net46),
    .A(_1295_),
    .Y(_0418_));
 sg13g2_xnor2_1 _2552_ (.Y(_0419_),
    .A(_1291_),
    .B(_0418_));
 sg13g2_nor2_1 _2553_ (.A(_0410_),
    .B(_0419_),
    .Y(_0061_));
 sg13g2_nor2_1 _2554_ (.A(_1291_),
    .B(_0418_),
    .Y(_0420_));
 sg13g2_xnor2_1 _2555_ (.Y(_0421_),
    .A(net33),
    .B(_0420_));
 sg13g2_nor2_1 _2556_ (.A(net30),
    .B(_0421_),
    .Y(_0062_));
 sg13g2_nand2_1 _2557_ (.Y(_0422_),
    .A(net33),
    .B(_0420_));
 sg13g2_xor2_1 _2558_ (.B(_0422_),
    .A(_1309_),
    .X(_0423_));
 sg13g2_nor2_1 _2559_ (.A(net30),
    .B(_0423_),
    .Y(_0063_));
 sg13g2_nand3_1 _2560_ (.B(net45),
    .C(_0420_),
    .A(net33),
    .Y(_0424_));
 sg13g2_xnor2_1 _2561_ (.Y(_0425_),
    .A(_1315_),
    .B(_0424_));
 sg13g2_nor2_1 _2562_ (.A(net30),
    .B(_0425_),
    .Y(_0064_));
 sg13g2_or2_1 _2563_ (.X(_0426_),
    .B(_0424_),
    .A(_1315_));
 sg13g2_xnor2_1 _2564_ (.Y(_0427_),
    .A(_1324_),
    .B(_0426_));
 sg13g2_nor2_1 _2565_ (.A(net30),
    .B(_0427_),
    .Y(_0065_));
 sg13g2_nor2_1 _2566_ (.A(_1324_),
    .B(_0426_),
    .Y(_0428_));
 sg13g2_xnor2_1 _2567_ (.Y(_0429_),
    .A(net44),
    .B(_0428_));
 sg13g2_nor2_1 _2568_ (.A(net30),
    .B(_0429_),
    .Y(_0066_));
 sg13g2_nand2_1 _2569_ (.Y(_0430_),
    .A(_0017_),
    .B(_1253_));
 sg13g2_buf_2 _2570_ (.A(\ctr_audio[0] ),
    .X(_0431_));
 sg13g2_nand2b_1 _2571_ (.Y(_0432_),
    .B(_0431_),
    .A_N(_1253_));
 sg13g2_a21oi_1 _2572_ (.A1(_0430_),
    .A2(_0432_),
    .Y(_0067_),
    .B1(net48));
 sg13g2_buf_1 _2573_ (.A(net48),
    .X(_0433_));
 sg13g2_inv_1 _2574_ (.Y(_0434_),
    .A(\ctr_audio[7] ));
 sg13g2_inv_1 _2575_ (.Y(_0435_),
    .A(\ctr_audio[8] ));
 sg13g2_and4_1 _2576_ (.A(\ctr_audio[1] ),
    .B(_0431_),
    .C(\ctr_audio[2] ),
    .D(\ctr_audio[3] ),
    .X(_0436_));
 sg13g2_and4_1 _2577_ (.A(_1249_),
    .B(_1250_),
    .C(_1251_),
    .D(_0436_),
    .X(_0437_));
 sg13g2_buf_2 _2578_ (.A(_0437_),
    .X(_0438_));
 sg13g2_nand4_1 _2579_ (.B(\ctr_audio[5] ),
    .C(\ctr_audio[6] ),
    .A(\ctr_audio[4] ),
    .Y(_0439_),
    .D(_0438_));
 sg13g2_nor3_2 _2580_ (.A(_0434_),
    .B(_0435_),
    .C(_0439_),
    .Y(_0440_));
 sg13g2_nand2_1 _2581_ (.Y(_0441_),
    .A(\ctr_audio[9] ),
    .B(_0440_));
 sg13g2_xor2_1 _2582_ (.B(_0441_),
    .A(\Voice1.pulsewidth[0] ),
    .X(_0442_));
 sg13g2_nor2_1 _2583_ (.A(net29),
    .B(_0442_),
    .Y(_0068_));
 sg13g2_and3_1 _2584_ (.X(_0443_),
    .A(\Voice1.pulsewidth[0] ),
    .B(\ctr_audio[9] ),
    .C(_0440_));
 sg13g2_buf_1 _2585_ (.A(_0443_),
    .X(_0444_));
 sg13g2_xnor2_1 _2586_ (.Y(_0445_),
    .A(_0360_),
    .B(_0444_));
 sg13g2_nor2_1 _2587_ (.A(net29),
    .B(_0445_),
    .Y(_0069_));
 sg13g2_nand2_1 _2588_ (.Y(_0446_),
    .A(_0360_),
    .B(_0444_));
 sg13g2_xnor2_1 _2589_ (.Y(_0447_),
    .A(_0359_),
    .B(_0446_));
 sg13g2_nor2_1 _2590_ (.A(net29),
    .B(_0447_),
    .Y(_0070_));
 sg13g2_and3_1 _2591_ (.X(_0448_),
    .A(\Voice1.pulsewidth[2] ),
    .B(_0360_),
    .C(_0444_));
 sg13g2_xnor2_1 _2592_ (.Y(_0449_),
    .A(\Voice1.pulsewidth[3] ),
    .B(_0448_));
 sg13g2_nor2_1 _2593_ (.A(net29),
    .B(_0449_),
    .Y(_0071_));
 sg13g2_nand4_1 _2594_ (.B(\Voice1.pulsewidth[2] ),
    .C(_0360_),
    .A(\Voice1.pulsewidth[3] ),
    .Y(_0450_),
    .D(_0444_));
 sg13g2_buf_1 _2595_ (.A(_0450_),
    .X(_0451_));
 sg13g2_xnor2_1 _2596_ (.Y(_0452_),
    .A(_0357_),
    .B(_0451_));
 sg13g2_nor2_1 _2597_ (.A(net29),
    .B(_0452_),
    .Y(_0072_));
 sg13g2_nor2_1 _2598_ (.A(_0357_),
    .B(_0451_),
    .Y(_0453_));
 sg13g2_xnor2_1 _2599_ (.Y(_0454_),
    .A(\Voice1.pulsewidth[5] ),
    .B(_0453_));
 sg13g2_nor2_1 _2600_ (.A(net29),
    .B(_0454_),
    .Y(_0073_));
 sg13g2_nor3_2 _2601_ (.A(_0356_),
    .B(_0357_),
    .C(_0451_),
    .Y(_0455_));
 sg13g2_xnor2_1 _2602_ (.Y(_0456_),
    .A(_0370_),
    .B(_0455_));
 sg13g2_nor2_1 _2603_ (.A(net29),
    .B(_0456_),
    .Y(_0074_));
 sg13g2_nand2_1 _2604_ (.Y(_0457_),
    .A(_0370_),
    .B(_0455_));
 sg13g2_xnor2_1 _2605_ (.Y(_0458_),
    .A(_0996_),
    .B(_0457_));
 sg13g2_nor2_1 _2606_ (.A(net29),
    .B(_0458_),
    .Y(_0075_));
 sg13g2_nand3_1 _2607_ (.B(_0370_),
    .C(_0455_),
    .A(net50),
    .Y(_0459_));
 sg13g2_xnor2_1 _2608_ (.Y(_0460_),
    .A(_0354_),
    .B(_0459_));
 sg13g2_nor2_1 _2609_ (.A(_0433_),
    .B(_0460_),
    .Y(_0076_));
 sg13g2_and4_1 _2610_ (.A(\Voice1.pulsewidth[8] ),
    .B(net50),
    .C(_0370_),
    .D(_0455_),
    .X(_0461_));
 sg13g2_xnor2_1 _2611_ (.Y(_0462_),
    .A(net53),
    .B(_0461_));
 sg13g2_nor2_1 _2612_ (.A(_0433_),
    .B(_0462_),
    .Y(_0077_));
 sg13g2_buf_1 _2613_ (.A(_1235_),
    .X(_0463_));
 sg13g2_nand2_1 _2614_ (.Y(_0464_),
    .A(_0431_),
    .B(_1253_));
 sg13g2_xor2_1 _2615_ (.B(_0464_),
    .A(\ctr_audio[1] ),
    .X(_0465_));
 sg13g2_nor2_1 _2616_ (.A(net28),
    .B(_0465_),
    .Y(_0078_));
 sg13g2_and2_1 _2617_ (.A(net53),
    .B(_0461_),
    .X(_0466_));
 sg13g2_buf_1 _2618_ (.A(_0466_),
    .X(_0467_));
 sg13g2_xnor2_1 _2619_ (.Y(_0468_),
    .A(\ctr_audio[20] ),
    .B(_0467_));
 sg13g2_nor2_1 _2620_ (.A(net28),
    .B(_0468_),
    .Y(_0079_));
 sg13g2_nand2_1 _2621_ (.Y(_0469_),
    .A(\ctr_audio[20] ),
    .B(_0467_));
 sg13g2_xnor2_1 _2622_ (.Y(_0470_),
    .A(_0990_),
    .B(_0469_));
 sg13g2_nor2_1 _2623_ (.A(net28),
    .B(_0470_),
    .Y(_0080_));
 sg13g2_nand3_1 _2624_ (.B(net51),
    .C(_0467_),
    .A(\ctr_audio[20] ),
    .Y(_0471_));
 sg13g2_xor2_1 _2625_ (.B(_0471_),
    .A(net49),
    .X(_0472_));
 sg13g2_nor2_1 _2626_ (.A(_0463_),
    .B(_0472_),
    .Y(_0081_));
 sg13g2_nor2_1 _2627_ (.A(_1011_),
    .B(_0469_),
    .Y(_0473_));
 sg13g2_xnor2_1 _2628_ (.Y(_0474_),
    .A(net52),
    .B(_0473_));
 sg13g2_nor2_1 _2629_ (.A(_0463_),
    .B(_0474_),
    .Y(_0082_));
 sg13g2_nand3_1 _2630_ (.B(_0431_),
    .C(_1253_),
    .A(\ctr_audio[1] ),
    .Y(_0475_));
 sg13g2_xor2_1 _2631_ (.B(_0475_),
    .A(\ctr_audio[2] ),
    .X(_0476_));
 sg13g2_nor2_1 _2632_ (.A(net28),
    .B(_0476_),
    .Y(_0083_));
 sg13g2_nand4_1 _2633_ (.B(_0431_),
    .C(\ctr_audio[2] ),
    .A(\ctr_audio[1] ),
    .Y(_0477_),
    .D(_1253_));
 sg13g2_xor2_1 _2634_ (.B(_0477_),
    .A(\ctr_audio[3] ),
    .X(_0478_));
 sg13g2_nor2_1 _2635_ (.A(net28),
    .B(_0478_),
    .Y(_0084_));
 sg13g2_xnor2_1 _2636_ (.Y(_0479_),
    .A(\ctr_audio[4] ),
    .B(_0438_));
 sg13g2_nor2_1 _2637_ (.A(net28),
    .B(_0479_),
    .Y(_0085_));
 sg13g2_nand2_1 _2638_ (.Y(_0480_),
    .A(\ctr_audio[4] ),
    .B(_0438_));
 sg13g2_xor2_1 _2639_ (.B(_0480_),
    .A(\ctr_audio[5] ),
    .X(_0481_));
 sg13g2_nor2_1 _2640_ (.A(net28),
    .B(_0481_),
    .Y(_0086_));
 sg13g2_nand3_1 _2641_ (.B(\ctr_audio[5] ),
    .C(_0438_),
    .A(\ctr_audio[4] ),
    .Y(_0482_));
 sg13g2_xor2_1 _2642_ (.B(_0482_),
    .A(\ctr_audio[6] ),
    .X(_0483_));
 sg13g2_nor2_1 _2643_ (.A(net28),
    .B(_0483_),
    .Y(_0087_));
 sg13g2_buf_1 _2644_ (.A(_1235_),
    .X(_0484_));
 sg13g2_xnor2_1 _2645_ (.Y(_0485_),
    .A(_0434_),
    .B(_0439_));
 sg13g2_nor2_1 _2646_ (.A(net27),
    .B(_0485_),
    .Y(_0088_));
 sg13g2_nor2_1 _2647_ (.A(_0434_),
    .B(_0439_),
    .Y(_0486_));
 sg13g2_xnor2_1 _2648_ (.Y(_0487_),
    .A(\ctr_audio[8] ),
    .B(_0486_));
 sg13g2_nor2_1 _2649_ (.A(net27),
    .B(_0487_),
    .Y(_0089_));
 sg13g2_xnor2_1 _2650_ (.Y(_0488_),
    .A(\ctr_audio[9] ),
    .B(_0440_));
 sg13g2_nor2_1 _2651_ (.A(net27),
    .B(_0488_),
    .Y(_0090_));
 sg13g2_buf_1 _2652_ (.A(\VAL[0] ),
    .X(_0489_));
 sg13g2_xnor2_1 _2653_ (.Y(_0490_),
    .A(net57),
    .B(_0489_));
 sg13g2_nor2_1 _2654_ (.A(net27),
    .B(_0490_),
    .Y(_0099_));
 sg13g2_nand2_1 _2655_ (.Y(_0491_),
    .A(net57),
    .B(_0489_));
 sg13g2_xnor2_1 _2656_ (.Y(_0492_),
    .A(net62),
    .B(\VAL[1] ));
 sg13g2_xnor2_1 _2657_ (.Y(_0493_),
    .A(_0491_),
    .B(_0492_));
 sg13g2_nor2_1 _2658_ (.A(net27),
    .B(_0493_),
    .Y(_0100_));
 sg13g2_a21oi_1 _2659_ (.A1(net71),
    .A2(_0489_),
    .Y(_0494_),
    .B1(\VAL[1] ));
 sg13g2_nand3_1 _2660_ (.B(\VAL[1] ),
    .C(_0489_),
    .A(net57),
    .Y(_0495_));
 sg13g2_o21ai_1 _2661_ (.B1(_0495_),
    .Y(_0496_),
    .A1(_0387_),
    .A2(_0494_));
 sg13g2_buf_1 _2662_ (.A(\VAL[2] ),
    .X(_0497_));
 sg13g2_xor2_1 _2663_ (.B(_0497_),
    .A(net35),
    .X(_0498_));
 sg13g2_xnor2_1 _2664_ (.Y(_0499_),
    .A(_0496_),
    .B(_0498_));
 sg13g2_nor2_1 _2665_ (.A(net27),
    .B(_0499_),
    .Y(_0101_));
 sg13g2_nor2_1 _2666_ (.A(_0497_),
    .B(_0496_),
    .Y(_0500_));
 sg13g2_a21oi_1 _2667_ (.A1(_0497_),
    .A2(_0496_),
    .Y(_0501_),
    .B1(net60));
 sg13g2_nor2_1 _2668_ (.A(_0500_),
    .B(_0501_),
    .Y(_0502_));
 sg13g2_xor2_1 _2669_ (.B(\VAL[3] ),
    .A(_0930_),
    .X(_0503_));
 sg13g2_xnor2_1 _2670_ (.Y(_0504_),
    .A(_0502_),
    .B(_0503_));
 sg13g2_nor2_1 _2671_ (.A(net27),
    .B(_0504_),
    .Y(_0102_));
 sg13g2_a21o_1 _2672_ (.A2(_0502_),
    .A1(\VAL[3] ),
    .B1(net61),
    .X(_0505_));
 sg13g2_o21ai_1 _2673_ (.B1(_0505_),
    .Y(_0506_),
    .A1(\VAL[3] ),
    .A2(_0502_));
 sg13g2_xnor2_1 _2674_ (.Y(_0507_),
    .A(_0935_),
    .B(\VAL[4] ));
 sg13g2_xnor2_1 _2675_ (.Y(_0508_),
    .A(_0506_),
    .B(_0507_));
 sg13g2_nor2_1 _2676_ (.A(net27),
    .B(_0508_),
    .Y(_0103_));
 sg13g2_inv_1 _2677_ (.Y(_0509_),
    .A(\VAL[4] ));
 sg13g2_inv_1 _2678_ (.Y(_0510_),
    .A(_0506_));
 sg13g2_a21oi_1 _2679_ (.A1(\VAL[4] ),
    .A2(_0510_),
    .Y(_0511_),
    .B1(_0935_));
 sg13g2_a21oi_1 _2680_ (.A1(_0509_),
    .A2(_0506_),
    .Y(_0512_),
    .B1(_0511_));
 sg13g2_nand2b_1 _2681_ (.Y(_0513_),
    .B(_0512_),
    .A_N(_0011_));
 sg13g2_nand2b_1 _2682_ (.Y(_0514_),
    .B(_0011_),
    .A_N(_0512_));
 sg13g2_and3_1 _2683_ (.X(_0104_),
    .A(_1091_),
    .B(_0513_),
    .C(_0514_));
 sg13g2_xnor2_1 _2684_ (.Y(_0515_),
    .A(_0008_),
    .B(_0513_));
 sg13g2_nor2_1 _2685_ (.A(_0484_),
    .B(_0515_),
    .Y(_0105_));
 sg13g2_nand3_1 _2686_ (.B(\VAL[6] ),
    .C(_0512_),
    .A(\VAL[5] ),
    .Y(_0516_));
 sg13g2_xnor2_1 _2687_ (.Y(_0517_),
    .A(_0007_),
    .B(_0516_));
 sg13g2_nor2_1 _2688_ (.A(_0484_),
    .B(_0517_),
    .Y(_0106_));
 sg13g2_and2_1 _2689_ (.A(_0414_),
    .B(_1253_),
    .X(_0127_));
 sg13g2_nand2_1 _2690_ (.Y(_0518_),
    .A(_0959_),
    .B(_0006_));
 sg13g2_nand2_1 _2691_ (.Y(_0519_),
    .A(net70),
    .B(_0951_));
 sg13g2_xnor2_1 _2692_ (.Y(_0520_),
    .A(_0956_),
    .B(_0519_));
 sg13g2_or2_1 _2693_ (.X(_0521_),
    .B(_0520_),
    .A(_0518_));
 sg13g2_buf_1 _2694_ (.A(_0521_),
    .X(_0522_));
 sg13g2_xor2_1 _2695_ (.B(\yq[12] ),
    .A(\xq[11] ),
    .X(_0523_));
 sg13g2_buf_1 _2696_ (.A(_0523_),
    .X(_0524_));
 sg13g2_nor2b_1 _2697_ (.A(\xq[10] ),
    .B_N(\yq[11] ),
    .Y(_0525_));
 sg13g2_buf_1 _2698_ (.A(\xq[9] ),
    .X(_0526_));
 sg13g2_inv_1 _2699_ (.Y(_0527_),
    .A(_0526_));
 sg13g2_nor2b_1 _2700_ (.A(\xq[4] ),
    .B_N(\yq[5] ),
    .Y(_0528_));
 sg13g2_buf_2 _2701_ (.A(\xq[5] ),
    .X(_0529_));
 sg13g2_nor2b_1 _2702_ (.A(_0529_),
    .B_N(_0318_),
    .Y(_0530_));
 sg13g2_nand2b_1 _2703_ (.Y(_0531_),
    .B(_0529_),
    .A_N(_0318_));
 sg13g2_o21ai_1 _2704_ (.B1(_0531_),
    .Y(_0532_),
    .A1(_0528_),
    .A2(_0530_));
 sg13g2_buf_2 _2705_ (.A(_0532_),
    .X(_0533_));
 sg13g2_buf_8 _2706_ (.A(\xq[7] ),
    .X(_0534_));
 sg13g2_inv_2 _2707_ (.Y(_0535_),
    .A(_0534_));
 sg13g2_buf_2 _2708_ (.A(\xq[8] ),
    .X(_0536_));
 sg13g2_nor2b_1 _2709_ (.A(_0536_),
    .B_N(_0336_),
    .Y(_0537_));
 sg13g2_buf_1 _2710_ (.A(\xq[6] ),
    .X(_0538_));
 sg13g2_nor2b_1 _2711_ (.A(_0538_),
    .B_N(_0325_),
    .Y(_0539_));
 sg13g2_nor3_1 _2712_ (.A(_0535_),
    .B(_0537_),
    .C(_0539_),
    .Y(_0540_));
 sg13g2_inv_1 _2713_ (.Y(_0541_),
    .A(_0536_));
 sg13g2_nand2b_1 _2714_ (.Y(_0542_),
    .B(_0538_),
    .A_N(_0325_));
 sg13g2_a221oi_1 _2715_ (.B2(_0535_),
    .C1(_0542_),
    .B1(_0331_),
    .A1(_0336_),
    .Y(_0543_),
    .A2(_0541_));
 sg13g2_a21oi_1 _2716_ (.A1(_0533_),
    .A2(_0540_),
    .Y(_0544_),
    .B1(_0543_));
 sg13g2_nand2b_1 _2717_ (.Y(_0545_),
    .B(_0336_),
    .A_N(_0536_));
 sg13g2_nor2_1 _2718_ (.A(_0331_),
    .B(_0535_),
    .Y(_0546_));
 sg13g2_nor3_1 _2719_ (.A(_0331_),
    .B(_0537_),
    .C(_0539_),
    .Y(_0547_));
 sg13g2_a22oi_1 _2720_ (.Y(_0548_),
    .B1(_0547_),
    .B2(_0533_),
    .A2(_0546_),
    .A1(_0545_));
 sg13g2_buf_1 _2721_ (.A(_0548_),
    .X(_0549_));
 sg13g2_nor2b_1 _2722_ (.A(\yq[11] ),
    .B_N(\xq[10] ),
    .Y(_0550_));
 sg13g2_nor2b_1 _2723_ (.A(_0336_),
    .B_N(_0536_),
    .Y(_0551_));
 sg13g2_nor2_1 _2724_ (.A(_0550_),
    .B(_0551_),
    .Y(_0552_));
 sg13g2_and4_1 _2725_ (.A(_0527_),
    .B(_0544_),
    .C(_0549_),
    .D(_0552_),
    .X(_0553_));
 sg13g2_and4_1 _2726_ (.A(\yq[10] ),
    .B(_0544_),
    .C(_0549_),
    .D(_0552_),
    .X(_0554_));
 sg13g2_inv_1 _2727_ (.Y(_0555_),
    .A(\yq[10] ));
 sg13g2_nor3_1 _2728_ (.A(_0555_),
    .B(_0526_),
    .C(_0550_),
    .Y(_0556_));
 sg13g2_or4_1 _2729_ (.A(_0525_),
    .B(_0553_),
    .C(_0554_),
    .D(_0556_),
    .X(_0557_));
 sg13g2_buf_2 _2730_ (.A(_0557_),
    .X(_0558_));
 sg13g2_xnor2_1 _2731_ (.Y(_0559_),
    .A(net38),
    .B(_0558_));
 sg13g2_buf_2 _2732_ (.A(_0559_),
    .X(_0560_));
 sg13g2_xor2_1 _2733_ (.B(\yq[5] ),
    .A(\xq[4] ),
    .X(_0561_));
 sg13g2_xor2_1 _2734_ (.B(_1181_),
    .A(net58),
    .X(_0562_));
 sg13g2_xnor2_1 _2735_ (.Y(_0563_),
    .A(_0561_),
    .B(_0562_));
 sg13g2_xnor2_1 _2736_ (.Y(_0564_),
    .A(_0560_),
    .B(_0563_));
 sg13g2_nor2_1 _2737_ (.A(net17),
    .B(_0564_),
    .Y(_0128_));
 sg13g2_xor2_1 _2738_ (.B(_0529_),
    .A(_0318_),
    .X(_0565_));
 sg13g2_xnor2_1 _2739_ (.Y(_0566_),
    .A(_0528_),
    .B(_0565_));
 sg13g2_xor2_1 _2740_ (.B(_1179_),
    .A(net71),
    .X(_0567_));
 sg13g2_xnor2_1 _2741_ (.Y(_0568_),
    .A(_0566_),
    .B(_0567_));
 sg13g2_buf_2 _2742_ (.A(_0568_),
    .X(_0569_));
 sg13g2_nor2_1 _2743_ (.A(_1181_),
    .B(_0560_),
    .Y(_0570_));
 sg13g2_a21oi_1 _2744_ (.A1(_1181_),
    .A2(_0561_),
    .Y(_0571_),
    .B1(_0570_));
 sg13g2_mux2_1 _2745_ (.A0(_0561_),
    .A1(_0560_),
    .S(_1181_),
    .X(_0572_));
 sg13g2_nand2_1 _2746_ (.Y(_0573_),
    .A(net58),
    .B(_0572_));
 sg13g2_o21ai_1 _2747_ (.B1(_0573_),
    .Y(_0574_),
    .A1(net58),
    .A2(_0571_));
 sg13g2_xnor2_1 _2748_ (.Y(_0575_),
    .A(_0569_),
    .B(_0574_));
 sg13g2_nor2_1 _2749_ (.A(net17),
    .B(_0575_),
    .Y(_0129_));
 sg13g2_inv_1 _2750_ (.Y(_0576_),
    .A(_0566_));
 sg13g2_nor2_1 _2751_ (.A(_1180_),
    .B(_0576_),
    .Y(_0577_));
 sg13g2_nor2_1 _2752_ (.A(_1180_),
    .B(_0566_),
    .Y(_0578_));
 sg13g2_mux2_1 _2753_ (.A0(_0577_),
    .A1(_0578_),
    .S(_0560_),
    .X(_0579_));
 sg13g2_buf_2 _2754_ (.A(_0579_),
    .X(_0580_));
 sg13g2_xnor2_1 _2755_ (.Y(_0581_),
    .A(\xq[11] ),
    .B(\yq[12] ));
 sg13g2_buf_1 _2756_ (.A(_0581_),
    .X(_0582_));
 sg13g2_buf_1 _2757_ (.A(net37),
    .X(_0583_));
 sg13g2_nor4_2 _2758_ (.A(_0525_),
    .B(_0553_),
    .C(_0554_),
    .Y(_0584_),
    .D(_0556_));
 sg13g2_buf_8 _2759_ (.A(_0584_),
    .X(_0585_));
 sg13g2_nor4_1 _2760_ (.A(_1179_),
    .B(net26),
    .C(net14),
    .D(_0576_),
    .Y(_0586_));
 sg13g2_buf_1 _2761_ (.A(net38),
    .X(_0587_));
 sg13g2_buf_8 _2762_ (.A(_0558_),
    .X(_0588_));
 sg13g2_nor4_1 _2763_ (.A(_1179_),
    .B(_0587_),
    .C(net12),
    .D(_0576_),
    .Y(_0589_));
 sg13g2_nor3_1 _2764_ (.A(_1179_),
    .B(net37),
    .C(_0566_),
    .Y(_0590_));
 sg13g2_nor3_1 _2765_ (.A(_1179_),
    .B(net38),
    .C(_0566_),
    .Y(_0591_));
 sg13g2_mux2_1 _2766_ (.A0(_0590_),
    .A1(_0591_),
    .S(_0558_),
    .X(_0592_));
 sg13g2_nor4_2 _2767_ (.A(_0942_),
    .B(_0586_),
    .C(_0589_),
    .Y(_0593_),
    .D(_0592_));
 sg13g2_nor2_2 _2768_ (.A(_0580_),
    .B(_0593_),
    .Y(_0594_));
 sg13g2_and2_1 _2769_ (.A(net58),
    .B(_1181_),
    .X(_0595_));
 sg13g2_buf_1 _2770_ (.A(_0595_),
    .X(_0596_));
 sg13g2_inv_1 _2771_ (.Y(_0597_),
    .A(_0569_));
 sg13g2_nand3_1 _2772_ (.B(_0596_),
    .C(_0597_),
    .A(net38),
    .Y(_0598_));
 sg13g2_nand3_1 _2773_ (.B(_0596_),
    .C(_0597_),
    .A(net37),
    .Y(_0599_));
 sg13g2_mux2_1 _2774_ (.A0(_0598_),
    .A1(_0599_),
    .S(_0558_),
    .X(_0600_));
 sg13g2_nand3_1 _2775_ (.B(_0596_),
    .C(_0569_),
    .A(net38),
    .Y(_0601_));
 sg13g2_nand3_1 _2776_ (.B(_0596_),
    .C(_0569_),
    .A(net37),
    .Y(_0602_));
 sg13g2_mux2_1 _2777_ (.A0(_0601_),
    .A1(_0602_),
    .S(_0584_),
    .X(_0603_));
 sg13g2_or2_1 _2778_ (.X(_0604_),
    .B(_1181_),
    .A(net58));
 sg13g2_buf_1 _2779_ (.A(_0604_),
    .X(_0605_));
 sg13g2_nor2_1 _2780_ (.A(_0561_),
    .B(_0569_),
    .Y(_0606_));
 sg13g2_nand3_1 _2781_ (.B(_0605_),
    .C(_0606_),
    .A(_0524_),
    .Y(_0607_));
 sg13g2_nand3_1 _2782_ (.B(_0605_),
    .C(_0606_),
    .A(_0582_),
    .Y(_0608_));
 sg13g2_mux2_1 _2783_ (.A0(_0607_),
    .A1(_0608_),
    .S(_0558_),
    .X(_0609_));
 sg13g2_nand4_1 _2784_ (.B(_0561_),
    .C(_0605_),
    .A(_0524_),
    .Y(_0610_),
    .D(_0569_));
 sg13g2_nand4_1 _2785_ (.B(_0561_),
    .C(_0605_),
    .A(_0582_),
    .Y(_0611_),
    .D(_0569_));
 sg13g2_mux2_1 _2786_ (.A0(_0610_),
    .A1(_0611_),
    .S(_0584_),
    .X(_0612_));
 sg13g2_nand4_1 _2787_ (.B(_0603_),
    .C(_0609_),
    .A(_0600_),
    .Y(_0613_),
    .D(_0612_));
 sg13g2_buf_1 _2788_ (.A(_0613_),
    .X(_0614_));
 sg13g2_nor2b_1 _2789_ (.A(_0325_),
    .B_N(_0538_),
    .Y(_0615_));
 sg13g2_nor2_1 _2790_ (.A(_0615_),
    .B(_0539_),
    .Y(_0616_));
 sg13g2_xnor2_1 _2791_ (.Y(_0617_),
    .A(_0533_),
    .B(_0616_));
 sg13g2_xor2_1 _2792_ (.B(_0617_),
    .A(_0560_),
    .X(_0618_));
 sg13g2_buf_2 _2793_ (.A(_0618_),
    .X(_0619_));
 sg13g2_xor2_1 _2794_ (.B(net67),
    .A(net72),
    .X(_0620_));
 sg13g2_xnor2_1 _2795_ (.Y(_0621_),
    .A(_0619_),
    .B(_0620_));
 sg13g2_xnor2_1 _2796_ (.Y(_0622_),
    .A(_0614_),
    .B(_0621_));
 sg13g2_xnor2_1 _2797_ (.Y(_0623_),
    .A(_0594_),
    .B(_0622_));
 sg13g2_nor2_1 _2798_ (.A(net17),
    .B(_0623_),
    .Y(_0130_));
 sg13g2_xnor2_1 _2799_ (.Y(_0624_),
    .A(net60),
    .B(net54));
 sg13g2_buf_2 _2800_ (.A(_0624_),
    .X(_0625_));
 sg13g2_nor2_2 _2801_ (.A(net72),
    .B(net67),
    .Y(_0626_));
 sg13g2_xor2_1 _2802_ (.B(_0626_),
    .A(_0625_),
    .X(_0627_));
 sg13g2_nand2b_1 _2803_ (.Y(_0628_),
    .B(_0325_),
    .A_N(_0538_));
 sg13g2_a21oi_2 _2804_ (.B1(_0615_),
    .Y(_0629_),
    .A2(_0628_),
    .A1(_0533_));
 sg13g2_nor2b_1 _2805_ (.A(_0534_),
    .B_N(_0331_),
    .Y(_0630_));
 sg13g2_nor2_1 _2806_ (.A(_0546_),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_xnor2_1 _2807_ (.Y(_0632_),
    .A(_0629_),
    .B(_0631_));
 sg13g2_buf_2 _2808_ (.A(_0632_),
    .X(_0633_));
 sg13g2_nor3_1 _2809_ (.A(net26),
    .B(_0627_),
    .C(_0633_),
    .Y(_0634_));
 sg13g2_nor3_1 _2810_ (.A(net25),
    .B(_0627_),
    .C(_0633_),
    .Y(_0635_));
 sg13g2_mux2_1 _2811_ (.A0(_0634_),
    .A1(_0635_),
    .S(net12),
    .X(_0636_));
 sg13g2_xor2_1 _2812_ (.B(_0631_),
    .A(_0629_),
    .X(_0637_));
 sg13g2_buf_2 _2813_ (.A(_0637_),
    .X(_0638_));
 sg13g2_nor3_1 _2814_ (.A(net26),
    .B(_0627_),
    .C(_0638_),
    .Y(_0639_));
 sg13g2_nor3_1 _2815_ (.A(net25),
    .B(_0627_),
    .C(_0638_),
    .Y(_0640_));
 sg13g2_mux2_1 _2816_ (.A0(_0639_),
    .A1(_0640_),
    .S(net14),
    .X(_0641_));
 sg13g2_xnor2_1 _2817_ (.Y(_0642_),
    .A(_0625_),
    .B(_0626_));
 sg13g2_nor3_1 _2818_ (.A(net26),
    .B(_0642_),
    .C(_0633_),
    .Y(_0643_));
 sg13g2_nor3_1 _2819_ (.A(net25),
    .B(_0642_),
    .C(_0633_),
    .Y(_0644_));
 sg13g2_mux2_1 _2820_ (.A0(_0643_),
    .A1(_0644_),
    .S(net14),
    .X(_0645_));
 sg13g2_nor3_1 _2821_ (.A(net26),
    .B(_0642_),
    .C(_0638_),
    .Y(_0646_));
 sg13g2_nor3_1 _2822_ (.A(_0587_),
    .B(_0642_),
    .C(_0638_),
    .Y(_0647_));
 sg13g2_mux2_1 _2823_ (.A0(_0646_),
    .A1(_0647_),
    .S(net12),
    .X(_0648_));
 sg13g2_nor4_2 _2824_ (.A(_0636_),
    .B(_0641_),
    .C(_0645_),
    .Y(_0649_),
    .D(_0648_));
 sg13g2_xnor2_1 _2825_ (.Y(_0650_),
    .A(net72),
    .B(net67));
 sg13g2_nor2_1 _2826_ (.A(_0619_),
    .B(_0650_),
    .Y(_0651_));
 sg13g2_nor2_1 _2827_ (.A(_0594_),
    .B(_0620_),
    .Y(_0652_));
 sg13g2_nand2_1 _2828_ (.Y(_0653_),
    .A(_0594_),
    .B(_0620_));
 sg13g2_o21ai_1 _2829_ (.B1(_0653_),
    .Y(_0654_),
    .A1(_0619_),
    .A2(_0652_));
 sg13g2_and4_1 _2830_ (.A(_0600_),
    .B(_0603_),
    .C(_0609_),
    .D(_0612_),
    .X(_0655_));
 sg13g2_and3_1 _2831_ (.X(_0656_),
    .A(_0614_),
    .B(_0619_),
    .C(_0652_));
 sg13g2_a221oi_1 _2832_ (.B2(_0655_),
    .C1(_0656_),
    .B1(_0654_),
    .A1(_0594_),
    .Y(_0657_),
    .A2(_0651_));
 sg13g2_xnor2_1 _2833_ (.Y(_0658_),
    .A(_0649_),
    .B(_0657_));
 sg13g2_nor2_1 _2834_ (.A(net17),
    .B(_0658_),
    .Y(_0131_));
 sg13g2_nor3_1 _2835_ (.A(_0580_),
    .B(_0593_),
    .C(_0649_),
    .Y(_0659_));
 sg13g2_a21oi_1 _2836_ (.A1(_0614_),
    .A2(_0650_),
    .Y(_0660_),
    .B1(_0649_));
 sg13g2_nor4_1 _2837_ (.A(_0580_),
    .B(_0593_),
    .C(_0614_),
    .D(_0650_),
    .Y(_0661_));
 sg13g2_nor4_1 _2838_ (.A(_0580_),
    .B(_0593_),
    .C(_0614_),
    .D(_0619_),
    .Y(_0662_));
 sg13g2_nor4_2 _2839_ (.A(_0659_),
    .B(_0660_),
    .C(_0661_),
    .Y(_0663_),
    .D(_0662_));
 sg13g2_nor2_1 _2840_ (.A(_0614_),
    .B(_0619_),
    .Y(_0664_));
 sg13g2_nor2_1 _2841_ (.A(_0619_),
    .B(_0649_),
    .Y(_0665_));
 sg13g2_a221oi_1 _2842_ (.B2(_0620_),
    .C1(_0665_),
    .B1(_0664_),
    .A1(_0594_),
    .Y(_0666_),
    .A2(_0651_));
 sg13g2_buf_1 _2843_ (.A(_0666_),
    .X(_0667_));
 sg13g2_and2_1 _2844_ (.A(_0663_),
    .B(_0667_),
    .X(_0668_));
 sg13g2_buf_1 _2845_ (.A(net38),
    .X(_0669_));
 sg13g2_nand2_1 _2846_ (.Y(_0670_),
    .A(net24),
    .B(_0638_));
 sg13g2_nand2_1 _2847_ (.Y(_0671_),
    .A(net26),
    .B(_0638_));
 sg13g2_mux2_1 _2848_ (.A0(_0670_),
    .A1(_0671_),
    .S(_0585_),
    .X(_0672_));
 sg13g2_nand2_1 _2849_ (.Y(_0673_),
    .A(net25),
    .B(_0633_));
 sg13g2_nand2_1 _2850_ (.Y(_0674_),
    .A(_0583_),
    .B(_0633_));
 sg13g2_mux2_1 _2851_ (.A0(_0673_),
    .A1(_0674_),
    .S(net12),
    .X(_0675_));
 sg13g2_a21o_1 _2852_ (.A2(_0675_),
    .A1(_0672_),
    .B1(_0625_),
    .X(_0676_));
 sg13g2_buf_1 _2853_ (.A(_0676_),
    .X(_0677_));
 sg13g2_nand3_1 _2854_ (.B(_0625_),
    .C(_0638_),
    .A(net25),
    .Y(_0678_));
 sg13g2_nand3_1 _2855_ (.B(_0625_),
    .C(_0638_),
    .A(net26),
    .Y(_0679_));
 sg13g2_mux2_1 _2856_ (.A0(_0678_),
    .A1(_0679_),
    .S(_0588_),
    .X(_0680_));
 sg13g2_nand4_1 _2857_ (.B(_0588_),
    .C(_0625_),
    .A(net24),
    .Y(_0681_),
    .D(_0633_));
 sg13g2_buf_1 _2858_ (.A(net26),
    .X(_0682_));
 sg13g2_nand4_1 _2859_ (.B(_0585_),
    .C(_0625_),
    .A(net19),
    .Y(_0683_),
    .D(_0633_));
 sg13g2_nand4_1 _2860_ (.B(_0680_),
    .C(_0681_),
    .A(_0626_),
    .Y(_0684_),
    .D(_0683_));
 sg13g2_buf_1 _2861_ (.A(_0684_),
    .X(_0685_));
 sg13g2_nand2_1 _2862_ (.Y(_0686_),
    .A(_0677_),
    .B(_0685_));
 sg13g2_nand2b_1 _2863_ (.Y(_0687_),
    .B(_0534_),
    .A_N(_0331_));
 sg13g2_or3_1 _2864_ (.A(_0528_),
    .B(_0530_),
    .C(_0539_),
    .X(_0688_));
 sg13g2_nor2b_1 _2865_ (.A(_0318_),
    .B_N(_0529_),
    .Y(_0689_));
 sg13g2_a21oi_1 _2866_ (.A1(_0689_),
    .A2(_0628_),
    .Y(_0690_),
    .B1(_0615_));
 sg13g2_a21o_1 _2867_ (.A2(_0690_),
    .A1(_0688_),
    .B1(_0630_),
    .X(_0691_));
 sg13g2_nand2b_1 _2868_ (.Y(_0692_),
    .B(_0536_),
    .A_N(_0336_));
 sg13g2_nand2_1 _2869_ (.Y(_0693_),
    .A(_0545_),
    .B(_0692_));
 sg13g2_a21oi_1 _2870_ (.A1(_0687_),
    .A2(_0691_),
    .Y(_0694_),
    .B1(_0693_));
 sg13g2_buf_2 _2871_ (.A(_0694_),
    .X(_0695_));
 sg13g2_a21oi_1 _2872_ (.A1(_0688_),
    .A2(_0690_),
    .Y(_0696_),
    .B1(_0630_));
 sg13g2_nor2_1 _2873_ (.A(_0537_),
    .B(_0551_),
    .Y(_0697_));
 sg13g2_nor3_1 _2874_ (.A(_0546_),
    .B(_0696_),
    .C(_0697_),
    .Y(_0698_));
 sg13g2_buf_2 _2875_ (.A(_0698_),
    .X(_0699_));
 sg13g2_xor2_1 _2876_ (.B(net61),
    .A(net68),
    .X(_0700_));
 sg13g2_nor2_1 _2877_ (.A(net37),
    .B(_0700_),
    .Y(_0701_));
 sg13g2_o21ai_1 _2878_ (.B1(_0701_),
    .Y(_0702_),
    .A1(_0695_),
    .A2(_0699_));
 sg13g2_nor2_1 _2879_ (.A(net38),
    .B(_0700_),
    .Y(_0703_));
 sg13g2_o21ai_1 _2880_ (.B1(_0703_),
    .Y(_0704_),
    .A1(_0695_),
    .A2(_0699_));
 sg13g2_mux2_1 _2881_ (.A0(_0702_),
    .A1(_0704_),
    .S(net12),
    .X(_0705_));
 sg13g2_o21ai_1 _2882_ (.B1(_0697_),
    .Y(_0706_),
    .A1(_0546_),
    .A2(_0696_));
 sg13g2_buf_2 _2883_ (.A(_0706_),
    .X(_0707_));
 sg13g2_nand3_1 _2884_ (.B(_0691_),
    .C(_0693_),
    .A(_0687_),
    .Y(_0708_));
 sg13g2_buf_2 _2885_ (.A(_0708_),
    .X(_0709_));
 sg13g2_nand3_1 _2886_ (.B(_0709_),
    .C(_0701_),
    .A(_0707_),
    .Y(_0710_));
 sg13g2_nand3_1 _2887_ (.B(_0709_),
    .C(_0703_),
    .A(_0707_),
    .Y(_0711_));
 sg13g2_mux2_1 _2888_ (.A0(_0710_),
    .A1(_0711_),
    .S(net14),
    .X(_0712_));
 sg13g2_xnor2_1 _2889_ (.Y(_0713_),
    .A(net68),
    .B(net61));
 sg13g2_nor2_1 _2890_ (.A(net37),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_o21ai_1 _2891_ (.B1(_0714_),
    .Y(_0715_),
    .A1(_0695_),
    .A2(_0699_));
 sg13g2_nor2_1 _2892_ (.A(net38),
    .B(_0713_),
    .Y(_0716_));
 sg13g2_o21ai_1 _2893_ (.B1(_0716_),
    .Y(_0717_),
    .A1(_0695_),
    .A2(_0699_));
 sg13g2_mux2_1 _2894_ (.A0(_0715_),
    .A1(_0717_),
    .S(net14),
    .X(_0718_));
 sg13g2_nand3_1 _2895_ (.B(_0709_),
    .C(_0714_),
    .A(_0707_),
    .Y(_0719_));
 sg13g2_nand3_1 _2896_ (.B(_0709_),
    .C(_0716_),
    .A(_0707_),
    .Y(_0720_));
 sg13g2_mux2_1 _2897_ (.A0(_0719_),
    .A1(_0720_),
    .S(net12),
    .X(_0721_));
 sg13g2_nand4_1 _2898_ (.B(_0712_),
    .C(_0718_),
    .A(_0705_),
    .Y(_0722_),
    .D(_0721_));
 sg13g2_buf_1 _2899_ (.A(_0722_),
    .X(_0723_));
 sg13g2_nor2_1 _2900_ (.A(net35),
    .B(_0953_),
    .Y(_0724_));
 sg13g2_xnor2_1 _2901_ (.Y(_0725_),
    .A(_0723_),
    .B(_0724_));
 sg13g2_xnor2_1 _2902_ (.Y(_0726_),
    .A(_0686_),
    .B(_0725_));
 sg13g2_xnor2_1 _2903_ (.Y(_0727_),
    .A(_0668_),
    .B(_0726_));
 sg13g2_nor2_1 _2904_ (.A(_0522_),
    .B(_0727_),
    .Y(_0132_));
 sg13g2_a21oi_1 _2905_ (.A1(_0677_),
    .A2(_0685_),
    .Y(_0728_),
    .B1(_0723_));
 sg13g2_o21ai_1 _2906_ (.B1(net25),
    .Y(_0729_),
    .A1(_0695_),
    .A2(_0699_));
 sg13g2_o21ai_1 _2907_ (.B1(_0583_),
    .Y(_0730_),
    .A1(_0695_),
    .A2(_0699_));
 sg13g2_mux2_1 _2908_ (.A0(_0729_),
    .A1(_0730_),
    .S(net14),
    .X(_0731_));
 sg13g2_buf_1 _2909_ (.A(_0731_),
    .X(_0732_));
 sg13g2_nand3_1 _2910_ (.B(_0707_),
    .C(_0709_),
    .A(net25),
    .Y(_0733_));
 sg13g2_nand3_1 _2911_ (.B(_0707_),
    .C(_0709_),
    .A(net37),
    .Y(_0734_));
 sg13g2_mux2_1 _2912_ (.A0(_0733_),
    .A1(_0734_),
    .S(net12),
    .X(_0735_));
 sg13g2_buf_1 _2913_ (.A(_0735_),
    .X(_0736_));
 sg13g2_nand3_1 _2914_ (.B(_0732_),
    .C(_0736_),
    .A(_0700_),
    .Y(_0737_));
 sg13g2_a21o_1 _2915_ (.A2(_0736_),
    .A1(_0732_),
    .B1(_0700_),
    .X(_0738_));
 sg13g2_nand2_1 _2916_ (.Y(_0739_),
    .A(_0737_),
    .B(_0738_));
 sg13g2_nor2_1 _2917_ (.A(_0686_),
    .B(_0739_),
    .Y(_0740_));
 sg13g2_a21oi_1 _2918_ (.A1(_0663_),
    .A2(_0667_),
    .Y(_0741_),
    .B1(_0740_));
 sg13g2_o21ai_1 _2919_ (.B1(_0724_),
    .Y(_0742_),
    .A1(_0728_),
    .A2(_0741_));
 sg13g2_or2_1 _2920_ (.X(_0743_),
    .B(_0953_),
    .A(net60));
 sg13g2_buf_1 _2921_ (.A(_0743_),
    .X(_0744_));
 sg13g2_nand4_1 _2922_ (.B(_0685_),
    .C(_0723_),
    .A(_0677_),
    .Y(_0745_),
    .D(_0744_));
 sg13g2_nand3_1 _2923_ (.B(_0667_),
    .C(_0745_),
    .A(_0663_),
    .Y(_0746_));
 sg13g2_o21ai_1 _2924_ (.B1(_0746_),
    .Y(_0747_),
    .A1(_0668_),
    .A2(_0728_));
 sg13g2_nor2_1 _2925_ (.A(net61),
    .B(net37),
    .Y(_0748_));
 sg13g2_o21ai_1 _2926_ (.B1(_0748_),
    .Y(_0749_),
    .A1(_0695_),
    .A2(_0699_));
 sg13g2_nor2_1 _2927_ (.A(net61),
    .B(net25),
    .Y(_0750_));
 sg13g2_o21ai_1 _2928_ (.B1(_0750_),
    .Y(_0751_),
    .A1(_0695_),
    .A2(_0699_));
 sg13g2_mux2_1 _2929_ (.A0(_0749_),
    .A1(_0751_),
    .S(net14),
    .X(_0752_));
 sg13g2_nand4_1 _2930_ (.B(_0707_),
    .C(_0709_),
    .A(net14),
    .Y(_0753_),
    .D(_0748_));
 sg13g2_nand4_1 _2931_ (.B(_0707_),
    .C(_0709_),
    .A(net12),
    .Y(_0754_),
    .D(_0750_));
 sg13g2_nand4_1 _2932_ (.B(_0752_),
    .C(_0753_),
    .A(net68),
    .Y(_0755_),
    .D(_0754_));
 sg13g2_nand3_1 _2933_ (.B(_0732_),
    .C(_0736_),
    .A(net61),
    .Y(_0756_));
 sg13g2_nand2_1 _2934_ (.Y(_0757_),
    .A(_0755_),
    .B(_0756_));
 sg13g2_xor2_1 _2935_ (.B(_0934_),
    .A(net70),
    .X(_0758_));
 sg13g2_inv_1 _2936_ (.Y(_0759_),
    .A(_0758_));
 sg13g2_nand3_1 _2937_ (.B(_0549_),
    .C(_0692_),
    .A(_0544_),
    .Y(_0760_));
 sg13g2_xnor2_1 _2938_ (.Y(_0761_),
    .A(\yq[10] ),
    .B(_0526_));
 sg13g2_xnor2_1 _2939_ (.Y(_0762_),
    .A(_0760_),
    .B(_0761_));
 sg13g2_xnor2_1 _2940_ (.Y(_0763_),
    .A(_0759_),
    .B(_0762_));
 sg13g2_xnor2_1 _2941_ (.Y(_0764_),
    .A(_0560_),
    .B(_0763_));
 sg13g2_xnor2_1 _2942_ (.Y(_0765_),
    .A(_0757_),
    .B(_0764_));
 sg13g2_nor2_2 _2943_ (.A(_0518_),
    .B(_0520_),
    .Y(_0766_));
 sg13g2_nand2b_1 _2944_ (.Y(_0767_),
    .B(_0766_),
    .A_N(_0765_));
 sg13g2_a21oi_1 _2945_ (.A1(_0742_),
    .A2(_0747_),
    .Y(_0768_),
    .B1(_0767_));
 sg13g2_nand4_1 _2946_ (.B(_0742_),
    .C(_0747_),
    .A(_0766_),
    .Y(_0769_),
    .D(_0765_));
 sg13g2_nand2b_1 _2947_ (.Y(_0133_),
    .B(_0769_),
    .A_N(_0768_));
 sg13g2_nand2_1 _2948_ (.Y(_0770_),
    .A(_0723_),
    .B(_0744_));
 sg13g2_a21o_1 _2949_ (.A2(_0724_),
    .A1(_0739_),
    .B1(_0686_),
    .X(_0771_));
 sg13g2_a21oi_2 _2950_ (.B1(_0765_),
    .Y(_0772_),
    .A2(_0771_),
    .A1(_0770_));
 sg13g2_and2_1 _2951_ (.A(_0755_),
    .B(_0756_),
    .X(_0773_));
 sg13g2_a21oi_1 _2952_ (.A1(_0723_),
    .A2(_0744_),
    .Y(_0774_),
    .B1(_0764_));
 sg13g2_and2_1 _2953_ (.A(_0732_),
    .B(_0736_),
    .X(_0775_));
 sg13g2_and4_1 _2954_ (.A(net68),
    .B(_0752_),
    .C(_0753_),
    .D(_0754_),
    .X(_0776_));
 sg13g2_a221oi_1 _2955_ (.B2(net36),
    .C1(_0776_),
    .B1(_0775_),
    .A1(_0677_),
    .Y(_0777_),
    .A2(_0685_));
 sg13g2_xor2_1 _2956_ (.B(_0763_),
    .A(_0560_),
    .X(_0778_));
 sg13g2_a221oi_1 _2957_ (.B2(_0738_),
    .C1(_0744_),
    .B1(_0737_),
    .A1(_0677_),
    .Y(_0779_),
    .A2(_0685_));
 sg13g2_a221oi_1 _2958_ (.B2(_0778_),
    .C1(_0779_),
    .B1(_0777_),
    .A1(_0773_),
    .Y(_0780_),
    .A2(_0774_));
 sg13g2_a21oi_1 _2959_ (.A1(_0723_),
    .A2(_0744_),
    .Y(_0781_),
    .B1(_0778_));
 sg13g2_a22oi_1 _2960_ (.Y(_0782_),
    .B1(_0755_),
    .B2(_0756_),
    .A2(_0685_),
    .A1(_0677_));
 sg13g2_a22oi_1 _2961_ (.Y(_0783_),
    .B1(_0782_),
    .B2(_0764_),
    .A2(_0781_),
    .A1(_0757_));
 sg13g2_nand4_1 _2962_ (.B(_0667_),
    .C(_0780_),
    .A(_0663_),
    .Y(_0784_),
    .D(_0783_));
 sg13g2_buf_2 _2963_ (.A(_0784_),
    .X(_0785_));
 sg13g2_nand2b_1 _2964_ (.Y(_0786_),
    .B(_0785_),
    .A_N(_0772_));
 sg13g2_xor2_1 _2965_ (.B(_0762_),
    .A(_0560_),
    .X(_0787_));
 sg13g2_nor2_1 _2966_ (.A(_0759_),
    .B(_0787_),
    .Y(_0788_));
 sg13g2_a221oi_1 _2967_ (.B2(_0787_),
    .C1(_0776_),
    .B1(_0759_),
    .A1(net36),
    .Y(_0789_),
    .A2(_0775_));
 sg13g2_nor2_2 _2968_ (.A(_0788_),
    .B(_0789_),
    .Y(_0790_));
 sg13g2_nand4_1 _2969_ (.B(_0544_),
    .C(_0549_),
    .A(_0527_),
    .Y(_0791_),
    .D(_0692_));
 sg13g2_nand3_1 _2970_ (.B(_0534_),
    .C(_0545_),
    .A(_0526_),
    .Y(_0792_));
 sg13g2_nand3b_1 _2971_ (.B(_0545_),
    .C(_0526_),
    .Y(_0793_),
    .A_N(_0331_));
 sg13g2_a22oi_1 _2972_ (.Y(_0794_),
    .B1(_0792_),
    .B2(_0793_),
    .A2(_0690_),
    .A1(_0688_));
 sg13g2_nand2_1 _2973_ (.Y(_0795_),
    .A(_0526_),
    .B(_0551_));
 sg13g2_o21ai_1 _2974_ (.B1(_0795_),
    .Y(_0796_),
    .A1(_0535_),
    .A2(_0793_));
 sg13g2_or3_1 _2975_ (.A(_0555_),
    .B(_0794_),
    .C(_0796_),
    .X(_0797_));
 sg13g2_nand3_1 _2976_ (.B(_0791_),
    .C(_0797_),
    .A(_0550_),
    .Y(_0798_));
 sg13g2_buf_1 _2977_ (.A(_0798_),
    .X(_0799_));
 sg13g2_nand2b_1 _2978_ (.Y(_0800_),
    .B(\yq[11] ),
    .A_N(\xq[10] ));
 sg13g2_a21o_1 _2979_ (.A2(_0797_),
    .A1(_0791_),
    .B1(_0800_),
    .X(_0801_));
 sg13g2_buf_1 _2980_ (.A(_0801_),
    .X(_0802_));
 sg13g2_nand2_1 _2981_ (.Y(_0803_),
    .A(_0799_),
    .B(_0802_));
 sg13g2_xnor2_1 _2982_ (.Y(_0804_),
    .A(net19),
    .B(_0803_));
 sg13g2_or2_1 _2983_ (.X(_0805_),
    .B(net59),
    .A(net70));
 sg13g2_buf_1 _2984_ (.A(_0805_),
    .X(_0806_));
 sg13g2_nor2_1 _2985_ (.A(_0956_),
    .B(net73),
    .Y(_0807_));
 sg13g2_nor2_1 _2986_ (.A(_0947_),
    .B(_1191_),
    .Y(_0808_));
 sg13g2_nor2_1 _2987_ (.A(_0807_),
    .B(_0808_),
    .Y(_0809_));
 sg13g2_xnor2_1 _2988_ (.Y(_0810_),
    .A(_0806_),
    .B(_0809_));
 sg13g2_xnor2_1 _2989_ (.Y(_0811_),
    .A(_0804_),
    .B(_0810_));
 sg13g2_xor2_1 _2990_ (.B(_0811_),
    .A(_0790_),
    .X(_0812_));
 sg13g2_xnor2_1 _2991_ (.Y(_0813_),
    .A(_0786_),
    .B(_0812_));
 sg13g2_nor2_1 _2992_ (.A(net17),
    .B(_0813_),
    .Y(_0134_));
 sg13g2_nand4_1 _2993_ (.B(net73),
    .C(_1284_),
    .A(_0947_),
    .Y(_0814_),
    .D(_0806_));
 sg13g2_nor2_1 _2994_ (.A(net56),
    .B(net73),
    .Y(_0815_));
 sg13g2_nand3_1 _2995_ (.B(_0806_),
    .C(_0815_),
    .A(_0949_),
    .Y(_0816_));
 sg13g2_nor2_2 _2996_ (.A(net70),
    .B(net59),
    .Y(_0817_));
 sg13g2_nand3_1 _2997_ (.B(_0817_),
    .C(_0807_),
    .A(net55),
    .Y(_0818_));
 sg13g2_nand3_1 _2998_ (.B(_0817_),
    .C(_0808_),
    .A(net55),
    .Y(_0819_));
 sg13g2_nand4_1 _2999_ (.B(_0816_),
    .C(_0818_),
    .A(_0814_),
    .Y(_0820_),
    .D(_0819_));
 sg13g2_buf_1 _3000_ (.A(_0799_),
    .X(_0821_));
 sg13g2_buf_1 _3001_ (.A(_0802_),
    .X(_0822_));
 sg13g2_nor3_1 _3002_ (.A(_1191_),
    .B(_0948_),
    .C(_0817_),
    .Y(_0823_));
 sg13g2_nand2_1 _3003_ (.Y(_0824_),
    .A(net19),
    .B(_0823_));
 sg13g2_nor3_1 _3004_ (.A(_0956_),
    .B(net55),
    .C(_0817_),
    .Y(_0825_));
 sg13g2_nand2_1 _3005_ (.Y(_0826_),
    .A(net19),
    .B(_0825_));
 sg13g2_a22oi_1 _3006_ (.Y(_0827_),
    .B1(_0824_),
    .B2(_0826_),
    .A2(net10),
    .A1(net11));
 sg13g2_nand4_1 _3007_ (.B(_0821_),
    .C(net10),
    .A(net24),
    .Y(_0828_),
    .D(_0823_));
 sg13g2_nand4_1 _3008_ (.B(net11),
    .C(_0822_),
    .A(net24),
    .Y(_0829_),
    .D(_0825_));
 sg13g2_nand3b_1 _3009_ (.B(_0828_),
    .C(_0829_),
    .Y(_0830_),
    .A_N(_0827_));
 sg13g2_nand4_1 _3010_ (.B(net24),
    .C(_0817_),
    .A(_1284_),
    .Y(_0831_),
    .D(_0815_));
 sg13g2_nand4_1 _3011_ (.B(net55),
    .C(net24),
    .A(net56),
    .Y(_0832_),
    .D(_0817_));
 sg13g2_a22oi_1 _3012_ (.Y(_0833_),
    .B1(_0831_),
    .B2(_0832_),
    .A2(net10),
    .A1(net11));
 sg13g2_nand2_1 _3013_ (.Y(_0834_),
    .A(_0956_),
    .B(_1191_));
 sg13g2_nor4_1 _3014_ (.A(net55),
    .B(net24),
    .C(_0806_),
    .D(_0834_),
    .Y(_0835_));
 sg13g2_nand3_1 _3015_ (.B(net10),
    .C(_0835_),
    .A(net11),
    .Y(_0836_));
 sg13g2_or4_1 _3016_ (.A(_1186_),
    .B(net24),
    .C(_0803_),
    .D(_0806_),
    .X(_0837_));
 sg13g2_nand3b_1 _3017_ (.B(_0836_),
    .C(_0837_),
    .Y(_0838_),
    .A_N(_0833_));
 sg13g2_nor3_1 _3018_ (.A(_0956_),
    .B(net73),
    .C(net47),
    .Y(_0839_));
 sg13g2_nand2_1 _3019_ (.Y(_0840_),
    .A(_0669_),
    .B(_0839_));
 sg13g2_nor3_1 _3020_ (.A(net56),
    .B(_1191_),
    .C(net47),
    .Y(_0841_));
 sg13g2_nand2_1 _3021_ (.Y(_0842_),
    .A(_0669_),
    .B(_0841_));
 sg13g2_a22oi_1 _3022_ (.Y(_0843_),
    .B1(_0840_),
    .B2(_0842_),
    .A2(_0822_),
    .A1(_0821_));
 sg13g2_nand4_1 _3023_ (.B(net73),
    .C(net47),
    .A(net56),
    .Y(_0844_),
    .D(net19));
 sg13g2_nand3_1 _3024_ (.B(net19),
    .C(_0815_),
    .A(net55),
    .Y(_0845_));
 sg13g2_a22oi_1 _3025_ (.Y(_0846_),
    .B1(_0844_),
    .B2(_0845_),
    .A2(net10),
    .A1(net11));
 sg13g2_nand2_1 _3026_ (.Y(_0847_),
    .A(net56),
    .B(net73));
 sg13g2_nor3_1 _3027_ (.A(net55),
    .B(net19),
    .C(_0847_),
    .Y(_0848_));
 sg13g2_nand3_1 _3028_ (.B(net10),
    .C(_0848_),
    .A(net11),
    .Y(_0849_));
 sg13g2_nor3_1 _3029_ (.A(net47),
    .B(_0682_),
    .C(_0834_),
    .Y(_0850_));
 sg13g2_nand3_1 _3030_ (.B(net10),
    .C(_0850_),
    .A(net11),
    .Y(_0851_));
 sg13g2_nand4_1 _3031_ (.B(net11),
    .C(net10),
    .A(_0682_),
    .Y(_0852_),
    .D(_0839_));
 sg13g2_nand4_1 _3032_ (.B(_0799_),
    .C(_0802_),
    .A(net19),
    .Y(_0853_),
    .D(_0841_));
 sg13g2_nand4_1 _3033_ (.B(_0851_),
    .C(_0852_),
    .A(_0849_),
    .Y(_0854_),
    .D(_0853_));
 sg13g2_or3_1 _3034_ (.A(_0843_),
    .B(_0846_),
    .C(_0854_),
    .X(_0855_));
 sg13g2_nor4_1 _3035_ (.A(_0820_),
    .B(_0830_),
    .C(_0838_),
    .D(_0855_),
    .Y(_0856_));
 sg13g2_buf_1 _3036_ (.A(_0856_),
    .X(_0857_));
 sg13g2_and2_1 _3037_ (.A(_0766_),
    .B(_0811_),
    .X(_0858_));
 sg13g2_buf_1 _3038_ (.A(_0858_),
    .X(_0859_));
 sg13g2_nand3b_1 _3039_ (.B(_0857_),
    .C(_0859_),
    .Y(_0860_),
    .A_N(_0785_));
 sg13g2_nand3_1 _3040_ (.B(_0857_),
    .C(_0859_),
    .A(_0790_),
    .Y(_0861_));
 sg13g2_nand3_1 _3041_ (.B(_0857_),
    .C(_0859_),
    .A(_0772_),
    .Y(_0862_));
 sg13g2_nand4_1 _3042_ (.B(_0772_),
    .C(_0790_),
    .A(_0766_),
    .Y(_0863_),
    .D(_0857_));
 sg13g2_and4_1 _3043_ (.A(_0860_),
    .B(_0861_),
    .C(_0862_),
    .D(_0863_),
    .X(_0864_));
 sg13g2_nand3_1 _3044_ (.B(_0790_),
    .C(_0857_),
    .A(_0766_),
    .Y(_0865_));
 sg13g2_or2_1 _3045_ (.X(_0866_),
    .B(_0865_),
    .A(_0785_));
 sg13g2_nor4_1 _3046_ (.A(net17),
    .B(_0772_),
    .C(_0811_),
    .D(_0857_),
    .Y(_0867_));
 sg13g2_nand2_1 _3047_ (.Y(_0868_),
    .A(_0785_),
    .B(_0867_));
 sg13g2_or2_1 _3048_ (.X(_0869_),
    .B(_0857_),
    .A(_0790_));
 sg13g2_nor3_1 _3049_ (.A(net17),
    .B(_0772_),
    .C(_0869_),
    .Y(_0870_));
 sg13g2_nor3_1 _3050_ (.A(net17),
    .B(_0811_),
    .C(_0869_),
    .Y(_0871_));
 sg13g2_a21oi_1 _3051_ (.A1(_0785_),
    .A2(_0870_),
    .Y(_0872_),
    .B1(_0871_));
 sg13g2_nand4_1 _3052_ (.B(_0866_),
    .C(_0868_),
    .A(_0864_),
    .Y(_0135_),
    .D(_0872_));
 sg13g2_and2_1 _3053_ (.A(net39),
    .B(\xq[0] ),
    .X(_0148_));
 sg13g2_and2_1 _3054_ (.A(net39),
    .B(\xq[10] ),
    .X(_0149_));
 sg13g2_and2_1 _3055_ (.A(net39),
    .B(\xq[11] ),
    .X(_0150_));
 sg13g2_and2_1 _3056_ (.A(net39),
    .B(\xq[1] ),
    .X(_0151_));
 sg13g2_and2_1 _3057_ (.A(net39),
    .B(\xq[2] ),
    .X(_0152_));
 sg13g2_and2_1 _3058_ (.A(net39),
    .B(\xq[3] ),
    .X(_0153_));
 sg13g2_and2_1 _3059_ (.A(net39),
    .B(\xq[4] ),
    .X(_0154_));
 sg13g2_and2_1 _3060_ (.A(net39),
    .B(_0529_),
    .X(_0155_));
 sg13g2_and2_1 _3061_ (.A(net65),
    .B(_0538_),
    .X(_0156_));
 sg13g2_nor2_1 _3062_ (.A(net48),
    .B(_0535_),
    .Y(_0157_));
 sg13g2_nor2_1 _3063_ (.A(net48),
    .B(_0541_),
    .Y(_0158_));
 sg13g2_nor2_1 _3064_ (.A(net48),
    .B(_0527_),
    .Y(_0159_));
 sg13g2_nand3_1 _3065_ (.B(_0937_),
    .C(_0950_),
    .A(_1191_),
    .Y(_0873_));
 sg13g2_buf_1 _3066_ (.A(_0873_),
    .X(_0874_));
 sg13g2_inv_1 _3067_ (.Y(_0875_),
    .A(\LFSR[5] ));
 sg13g2_inv_1 _3068_ (.Y(_0876_),
    .A(\VAL[5] ));
 sg13g2_inv_1 _3069_ (.Y(_0877_),
    .A(_0497_));
 sg13g2_nand2_1 _3070_ (.Y(_0878_),
    .A(_0489_),
    .B(_1240_));
 sg13g2_nor2_1 _3071_ (.A(_1238_),
    .B(_0878_),
    .Y(_0879_));
 sg13g2_nor2_1 _3072_ (.A(\VAL[1] ),
    .B(_0879_),
    .Y(_0880_));
 sg13g2_a221oi_1 _3073_ (.B2(_0878_),
    .C1(_0880_),
    .B1(_1238_),
    .A1(_1237_),
    .Y(_0881_),
    .A2(_0877_));
 sg13g2_a21oi_1 _3074_ (.A1(_1244_),
    .A2(_0497_),
    .Y(_0882_),
    .B1(_0881_));
 sg13g2_nand2_1 _3075_ (.Y(_0883_),
    .A(_1245_),
    .B(_0882_));
 sg13g2_inv_1 _3076_ (.Y(_0884_),
    .A(\VAL[3] ));
 sg13g2_o21ai_1 _3077_ (.B1(_0884_),
    .Y(_0885_),
    .A1(_1245_),
    .A2(_0882_));
 sg13g2_a22oi_1 _3078_ (.Y(_0886_),
    .B1(_0883_),
    .B2(_0885_),
    .A2(_1246_),
    .A1(\VAL[4] ));
 sg13g2_a221oi_1 _3079_ (.B2(\LFSR[4] ),
    .C1(_0886_),
    .B1(_0509_),
    .A1(\LFSR[5] ),
    .Y(_0887_),
    .A2(_0876_));
 sg13g2_a21oi_1 _3080_ (.A1(_0875_),
    .A2(\VAL[5] ),
    .Y(_0888_),
    .B1(_0887_));
 sg13g2_nor2_1 _3081_ (.A(_0008_),
    .B(_0888_),
    .Y(_0889_));
 sg13g2_xor2_1 _3082_ (.B(_0889_),
    .A(_0007_),
    .X(_0890_));
 sg13g2_nor2_1 _3083_ (.A(_0874_),
    .B(_0890_),
    .Y(net2));
 sg13g2_inv_1 _3084_ (.Y(_0891_),
    .A(\VAL[13] ));
 sg13g2_inv_1 _3085_ (.Y(_0892_),
    .A(_0391_));
 sg13g2_a21oi_1 _3086_ (.A1(_1240_),
    .A2(_0381_),
    .Y(_0893_),
    .B1(_0384_));
 sg13g2_nand3_1 _3087_ (.B(_0384_),
    .C(_0381_),
    .A(_1240_),
    .Y(_0894_));
 sg13g2_o21ai_1 _3088_ (.B1(_0894_),
    .Y(_0895_),
    .A1(_1238_),
    .A2(_0893_));
 sg13g2_a21oi_1 _3089_ (.A1(_1244_),
    .A2(_0391_),
    .Y(_0896_),
    .B1(_0895_));
 sg13g2_a21oi_1 _3090_ (.A1(_1237_),
    .A2(_0892_),
    .Y(_0897_),
    .B1(_0896_));
 sg13g2_nor2_1 _3091_ (.A(_0397_),
    .B(_0897_),
    .Y(_0898_));
 sg13g2_nor2_1 _3092_ (.A(_1245_),
    .B(_0898_),
    .Y(_0899_));
 sg13g2_a221oi_1 _3093_ (.B2(_0897_),
    .C1(_0899_),
    .B1(_0397_),
    .A1(_1246_),
    .Y(_0900_),
    .A2(\VAL[12] ));
 sg13g2_a221oi_1 _3094_ (.B2(\LFSR[4] ),
    .C1(_0900_),
    .B1(_0404_),
    .A1(\LFSR[5] ),
    .Y(_0901_),
    .A2(_0891_));
 sg13g2_a21oi_1 _3095_ (.A1(_0875_),
    .A2(\VAL[13] ),
    .Y(_0902_),
    .B1(_0901_));
 sg13g2_nor2_1 _3096_ (.A(_0009_),
    .B(_0902_),
    .Y(_0903_));
 sg13g2_xor2_1 _3097_ (.B(_0903_),
    .A(_0010_),
    .X(_0904_));
 sg13g2_nor2_1 _3098_ (.A(_0874_),
    .B(_0904_),
    .Y(net3));
 sg13g2_inv_1 _3099_ (.Y(_0905_),
    .A(\VAL[21] ));
 sg13g2_inv_1 _3100_ (.Y(_0906_),
    .A(\VAL[20] ));
 sg13g2_inv_1 _3101_ (.Y(_0907_),
    .A(\VAL[18] ));
 sg13g2_a21oi_1 _3102_ (.A1(_1240_),
    .A2(\VAL[16] ),
    .Y(_0908_),
    .B1(\VAL[17] ));
 sg13g2_nand3_1 _3103_ (.B(\VAL[17] ),
    .C(\VAL[16] ),
    .A(_1240_),
    .Y(_0909_));
 sg13g2_o21ai_1 _3104_ (.B1(_0909_),
    .Y(_0910_),
    .A1(_1238_),
    .A2(_0908_));
 sg13g2_a21oi_1 _3105_ (.A1(_1244_),
    .A2(\VAL[18] ),
    .Y(_0911_),
    .B1(_0910_));
 sg13g2_a21oi_1 _3106_ (.A1(_1237_),
    .A2(_0907_),
    .Y(_0912_),
    .B1(_0911_));
 sg13g2_nor2_1 _3107_ (.A(\VAL[19] ),
    .B(_0912_),
    .Y(_0913_));
 sg13g2_nor2_1 _3108_ (.A(_1245_),
    .B(_0913_),
    .Y(_0914_));
 sg13g2_a221oi_1 _3109_ (.B2(_0912_),
    .C1(_0914_),
    .B1(\VAL[19] ),
    .A1(_1246_),
    .Y(_0915_),
    .A2(\VAL[20] ));
 sg13g2_a221oi_1 _3110_ (.B2(\LFSR[4] ),
    .C1(_0915_),
    .B1(_0906_),
    .A1(\LFSR[5] ),
    .Y(_0916_),
    .A2(_0905_));
 sg13g2_a21oi_1 _3111_ (.A1(_0875_),
    .A2(\VAL[21] ),
    .Y(_0917_),
    .B1(_0916_));
 sg13g2_nor2b_1 _3112_ (.A(_0917_),
    .B_N(\VAL[22] ),
    .Y(_0918_));
 sg13g2_xnor2_1 _3113_ (.Y(_0919_),
    .A(\VAL[23] ),
    .B(_0918_));
 sg13g2_nor2_1 _3114_ (.A(_0874_),
    .B(_0919_),
    .Y(net4));
 sg13g2_xor2_1 _3115_ (.B(_0888_),
    .A(\VAL[6] ),
    .X(_0920_));
 sg13g2_nor2_1 _3116_ (.A(_0874_),
    .B(_0920_),
    .Y(net6));
 sg13g2_and2_1 _3117_ (.A(_0009_),
    .B(_0902_),
    .X(_0921_));
 sg13g2_nor3_1 _3118_ (.A(_0874_),
    .B(_0903_),
    .C(_0921_),
    .Y(net7));
 sg13g2_xor2_1 _3119_ (.B(_0917_),
    .A(\VAL[22] ),
    .X(_0922_));
 sg13g2_nor2_1 _3120_ (.A(_0874_),
    .B(_0922_),
    .Y(net8));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \LFSR[0]$_SDFF_PP1__90  (.L_HI(net90));
 sg13g2_buf_1 _3123_ (.A(net76),
    .X(uio_oe[0]));
 sg13g2_buf_1 _3124_ (.A(net77),
    .X(uio_oe[1]));
 sg13g2_buf_1 _3125_ (.A(net78),
    .X(uio_oe[2]));
 sg13g2_buf_1 _3126_ (.A(net79),
    .X(uio_oe[3]));
 sg13g2_buf_1 _3127_ (.A(net80),
    .X(uio_oe[4]));
 sg13g2_buf_1 _3128_ (.A(net81),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3129_ (.A(net82),
    .X(uio_oe[6]));
 sg13g2_buf_1 _3130_ (.A(net121),
    .X(uio_oe[7]));
 sg13g2_buf_1 _3131_ (.A(net83),
    .X(uio_out[0]));
 sg13g2_buf_1 _3132_ (.A(net84),
    .X(uio_out[1]));
 sg13g2_buf_1 _3133_ (.A(net85),
    .X(uio_out[2]));
 sg13g2_buf_1 _3134_ (.A(net86),
    .X(uio_out[3]));
 sg13g2_buf_1 _3135_ (.A(net87),
    .X(uio_out[4]));
 sg13g2_buf_1 _3136_ (.A(net88),
    .X(uio_out[5]));
 sg13g2_buf_1 _3137_ (.A(net89),
    .X(uio_out[6]));
 sg13g2_buf_1 _3138_ (.A(\Voice1.pulse ),
    .X(net1));
 sg13g2_buf_1 _3139_ (.A(net75),
    .X(net5));
 sg13g2_buf_1 _3140_ (.A(hsync),
    .X(net9));
 sg13g2_dfrbp_1 \b[0]$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net122),
    .D(_0050_),
    .Q_N(_1611_),
    .Q(\VAL[16] ));
 sg13g2_dfrbp_1 \b[1]$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net123),
    .D(_0051_),
    .Q_N(_1610_),
    .Q(\VAL[17] ));
 sg13g2_dfrbp_1 \b[2]$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net124),
    .D(_0052_),
    .Q_N(_1609_),
    .Q(\VAL[18] ));
 sg13g2_dfrbp_1 \b[3]$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net125),
    .D(_0053_),
    .Q_N(_1608_),
    .Q(\VAL[19] ));
 sg13g2_dfrbp_1 \b[4]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net126),
    .D(_0054_),
    .Q_N(_1607_),
    .Q(\VAL[20] ));
 sg13g2_dfrbp_1 \b[5]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net127),
    .D(_0055_),
    .Q_N(_1606_),
    .Q(\VAL[21] ));
 sg13g2_dfrbp_1 \b[6]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net128),
    .D(_0056_),
    .Q_N(_1605_),
    .Q(\VAL[22] ));
 sg13g2_dfrbp_1 \b[7]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net129),
    .D(_0057_),
    .Q_N(_1604_),
    .Q(\VAL[23] ));
 sg13g2_dfrbp_1 \counter[0]$_SDFF_PN0_  (.CLK(net74),
    .RESET_B(net130),
    .D(_0058_),
    .Q_N(_0015_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 \counter[1]$_SDFF_PN0_  (.CLK(net75),
    .RESET_B(net131),
    .D(_0059_),
    .Q_N(_1603_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 \counter[2]$_SDFF_PN0_  (.CLK(net75),
    .RESET_B(net132),
    .D(_0060_),
    .Q_N(_1602_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 \counter[3]$_SDFF_PN0_  (.CLK(net75),
    .RESET_B(net133),
    .D(_0061_),
    .Q_N(_1601_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 \counter[4]$_SDFF_PN0_  (.CLK(net74),
    .RESET_B(net134),
    .D(_0062_),
    .Q_N(_1600_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 \counter[5]$_SDFF_PN0_  (.CLK(net74),
    .RESET_B(net135),
    .D(_0063_),
    .Q_N(_1599_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 \counter[6]$_SDFF_PN0_  (.CLK(net74),
    .RESET_B(net136),
    .D(_0064_),
    .Q_N(_1598_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 \counter[7]$_SDFF_PN0_  (.CLK(net74),
    .RESET_B(net137),
    .D(_0065_),
    .Q_N(_1597_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 \counter[8]$_SDFF_PN0_  (.CLK(net74),
    .RESET_B(net138),
    .D(_0066_),
    .Q_N(_1596_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 \ctr_audio[0]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net139),
    .D(_0067_),
    .Q_N(_0017_),
    .Q(\ctr_audio[0] ));
 sg13g2_dfrbp_1 \ctr_audio[10]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net140),
    .D(_0068_),
    .Q_N(_1595_),
    .Q(\Voice1.pulsewidth[0] ));
 sg13g2_dfrbp_1 \ctr_audio[11]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net141),
    .D(_0069_),
    .Q_N(_1594_),
    .Q(\Voice1.pulsewidth[1] ));
 sg13g2_dfrbp_1 \ctr_audio[12]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net142),
    .D(_0070_),
    .Q_N(_1593_),
    .Q(\Voice1.pulsewidth[2] ));
 sg13g2_dfrbp_1 \ctr_audio[13]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net143),
    .D(_0071_),
    .Q_N(_1592_),
    .Q(\Voice1.pulsewidth[3] ));
 sg13g2_dfrbp_1 \ctr_audio[14]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net144),
    .D(_0072_),
    .Q_N(_1591_),
    .Q(\Voice1.pulsewidth[4] ));
 sg13g2_dfrbp_1 \ctr_audio[15]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net145),
    .D(_0073_),
    .Q_N(_1590_),
    .Q(\Voice1.pulsewidth[5] ));
 sg13g2_dfrbp_1 \ctr_audio[16]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net146),
    .D(_0074_),
    .Q_N(_1589_),
    .Q(\Voice1.pulsewidth[6] ));
 sg13g2_dfrbp_1 \ctr_audio[17]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net147),
    .D(_0075_),
    .Q_N(_1588_),
    .Q(\Voice1.pulsewidth[7] ));
 sg13g2_dfrbp_1 \ctr_audio[18]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net148),
    .D(_0076_),
    .Q_N(_1587_),
    .Q(\Voice1.pulsewidth[8] ));
 sg13g2_dfrbp_1 \ctr_audio[19]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net149),
    .D(_0077_),
    .Q_N(_1586_),
    .Q(\ctr_audio[19] ));
 sg13g2_dfrbp_1 \ctr_audio[1]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net150),
    .D(_0078_),
    .Q_N(_1585_),
    .Q(\ctr_audio[1] ));
 sg13g2_dfrbp_1 \ctr_audio[20]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net151),
    .D(_0079_),
    .Q_N(_1584_),
    .Q(\ctr_audio[20] ));
 sg13g2_dfrbp_1 \ctr_audio[21]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net152),
    .D(_0080_),
    .Q_N(_1583_),
    .Q(\ctr_audio[21] ));
 sg13g2_dfrbp_1 \ctr_audio[22]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net153),
    .D(_0081_),
    .Q_N(_1582_),
    .Q(\ctr_audio[22] ));
 sg13g2_dfrbp_1 \ctr_audio[23]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net154),
    .D(_0082_),
    .Q_N(_1581_),
    .Q(\Voice1.pulsewidth[10] ));
 sg13g2_dfrbp_1 \ctr_audio[2]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net155),
    .D(_0083_),
    .Q_N(_1580_),
    .Q(\ctr_audio[2] ));
 sg13g2_dfrbp_1 \ctr_audio[3]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net156),
    .D(_0084_),
    .Q_N(_1579_),
    .Q(\ctr_audio[3] ));
 sg13g2_dfrbp_1 \ctr_audio[4]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net157),
    .D(_0085_),
    .Q_N(_1578_),
    .Q(\ctr_audio[4] ));
 sg13g2_dfrbp_1 \ctr_audio[5]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net158),
    .D(_0086_),
    .Q_N(_1577_),
    .Q(\ctr_audio[5] ));
 sg13g2_dfrbp_1 \ctr_audio[6]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net159),
    .D(_0087_),
    .Q_N(_1576_),
    .Q(\ctr_audio[6] ));
 sg13g2_dfrbp_1 \ctr_audio[7]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net160),
    .D(_0088_),
    .Q_N(_1575_),
    .Q(\ctr_audio[7] ));
 sg13g2_dfrbp_1 \ctr_audio[8]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net161),
    .D(_0089_),
    .Q_N(_1574_),
    .Q(\ctr_audio[8] ));
 sg13g2_dfrbp_1 \ctr_audio[9]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net162),
    .D(_0090_),
    .Q_N(_1573_),
    .Q(\ctr_audio[9] ));
 sg13g2_dfrbp_1 \ctr_clkdiv25[0]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net163),
    .D(_0091_),
    .Q_N(_0016_),
    .Q(\ctr_clkdiv25[0] ));
 sg13g2_dfrbp_1 \ctr_clkdiv25[1]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net164),
    .D(_0092_),
    .Q_N(_1572_),
    .Q(\ctr_clkdiv25[1] ));
 sg13g2_dfrbp_1 \ctr_clkdiv25[2]$_SDFF_PP0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net165),
    .D(_0093_),
    .Q_N(_1571_),
    .Q(\ctr_clkdiv25[2] ));
 sg13g2_dfrbp_1 \ctr_clkdiv25[3]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net166),
    .D(_0094_),
    .Q_N(_1570_),
    .Q(\ctr_clkdiv25[3] ));
 sg13g2_dfrbp_1 \ctr_clkdiv25[4]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net167),
    .D(_0095_),
    .Q_N(_1569_),
    .Q(\ctr_clkdiv25[4] ));
 sg13g2_dfrbp_1 \ctr_clkdiv25[5]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net168),
    .D(_0096_),
    .Q_N(_1568_),
    .Q(\ctr_clkdiv25[5] ));
 sg13g2_dfrbp_1 \ctr_clkdiv25[6]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net169),
    .D(_0097_),
    .Q_N(_1567_),
    .Q(\ctr_clkdiv25[6] ));
 sg13g2_dfrbp_1 \ctr_clkdiv25[7]$_SDFF_PP0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net170),
    .D(_0098_),
    .Q_N(_1566_),
    .Q(\ctr_clkdiv25[7] ));
 sg13g2_dfrbp_1 \g[0]$_SDFF_PN0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net171),
    .D(_0099_),
    .Q_N(_1565_),
    .Q(\VAL[8] ));
 sg13g2_dfrbp_1 \g[1]$_SDFF_PN0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net172),
    .D(_0100_),
    .Q_N(_1564_),
    .Q(\VAL[9] ));
 sg13g2_dfrbp_1 \g[2]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net173),
    .D(_0101_),
    .Q_N(_1563_),
    .Q(\VAL[10] ));
 sg13g2_dfrbp_1 \g[3]$_SDFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net174),
    .D(_0102_),
    .Q_N(_1562_),
    .Q(\VAL[11] ));
 sg13g2_dfrbp_1 \g[4]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net175),
    .D(_0103_),
    .Q_N(_1561_),
    .Q(\VAL[12] ));
 sg13g2_dfrbp_1 \g[5]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net176),
    .D(_0104_),
    .Q_N(_0012_),
    .Q(\VAL[13] ));
 sg13g2_dfrbp_1 \g[6]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net177),
    .D(_0105_),
    .Q_N(_0009_),
    .Q(\VAL[14] ));
 sg13g2_dfrbp_1 \g[7]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net178),
    .D(_0106_),
    .Q_N(_0010_),
    .Q(\VAL[15] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[0]$_SDFF_PP0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net179),
    .D(_0107_),
    .Q_N(_0018_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[1]$_SDFF_PP0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net180),
    .D(_0108_),
    .Q_N(_1560_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[2]$_SDFF_PP0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net181),
    .D(_0109_),
    .Q_N(_1559_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[3]$_SDFF_PP0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net182),
    .D(_0110_),
    .Q_N(_1558_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[4]$_SDFF_PP0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net183),
    .D(_0111_),
    .Q_N(_1557_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[5]$_SDFF_PP0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net184),
    .D(_0112_),
    .Q_N(_1556_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[6]$_SDFF_PP0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net185),
    .D(_0113_),
    .Q_N(_1555_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[7]$_SDFF_PP0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net186),
    .D(_0114_),
    .Q_N(_1554_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[8]$_SDFF_PP0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net187),
    .D(_0115_),
    .Q_N(_1553_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[9]$_SDFF_PP0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net188),
    .D(_0116_),
    .Q_N(_0006_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.hsync$_DFF_P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net189),
    .D(_0000_),
    .Q_N(_1552_),
    .Q(hsync));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[0]$_SDFFCE_PP0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net190),
    .D(_0117_),
    .Q_N(_0014_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[1]$_SDFFCE_PP0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net191),
    .D(_0118_),
    .Q_N(_1551_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[2]$_SDFFCE_PP0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net192),
    .D(_0119_),
    .Q_N(_1550_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[3]$_SDFFCE_PP0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net193),
    .D(_0120_),
    .Q_N(_1549_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[4]$_SDFFCE_PP0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net194),
    .D(_0121_),
    .Q_N(_1548_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[5]$_SDFFCE_PP0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net195),
    .D(_0122_),
    .Q_N(_1547_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[6]$_SDFFCE_PP0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net196),
    .D(_0123_),
    .Q_N(_1546_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[7]$_SDFFCE_PP0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net197),
    .D(_0124_),
    .Q_N(_1545_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[8]$_SDFFCE_PP0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net198),
    .D(_0125_),
    .Q_N(_1544_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[9]$_SDFFCE_PP0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net199),
    .D(_0126_),
    .Q_N(_1640_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.vsync$_DFF_P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net200),
    .D(_0001_),
    .Q_N(_1543_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 \pulse_1MHz$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net201),
    .D(_0127_),
    .Q_N(_0013_),
    .Q(\Voice1.en ));
 sg13g2_dfrbp_1 \r[0]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net202),
    .D(_0128_),
    .Q_N(_1542_),
    .Q(\VAL[0] ));
 sg13g2_dfrbp_1 \r[1]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net203),
    .D(_0129_),
    .Q_N(_1541_),
    .Q(\VAL[1] ));
 sg13g2_dfrbp_1 \r[2]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net204),
    .D(_0130_),
    .Q_N(_1540_),
    .Q(\VAL[2] ));
 sg13g2_dfrbp_1 \r[3]$_SDFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net205),
    .D(_0131_),
    .Q_N(_1539_),
    .Q(\VAL[3] ));
 sg13g2_dfrbp_1 \r[4]$_SDFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net206),
    .D(_0132_),
    .Q_N(_1538_),
    .Q(\VAL[4] ));
 sg13g2_dfrbp_1 \r[5]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net207),
    .D(_0133_),
    .Q_N(_0011_),
    .Q(\VAL[5] ));
 sg13g2_dfrbp_1 \r[6]$_SDFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net208),
    .D(_0134_),
    .Q_N(_0008_),
    .Q(\VAL[6] ));
 sg13g2_dfrbp_1 \r[7]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net209),
    .D(_0135_),
    .Q_N(_0007_),
    .Q(\VAL[7] ));
 sg13g2_dfrbp_1 \xq[0]$_SDFF_PP0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net210),
    .D(_0136_),
    .Q_N(_1537_),
    .Q(\xq[0] ));
 sg13g2_dfrbp_1 \xq[10]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net211),
    .D(_0137_),
    .Q_N(_1536_),
    .Q(\xq[10] ));
 sg13g2_dfrbp_1 \xq[11]$_SDFF_PP0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net212),
    .D(_0138_),
    .Q_N(_1535_),
    .Q(\xq[11] ));
 sg13g2_dfrbp_1 \xq[1]$_SDFF_PP0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net213),
    .D(_0139_),
    .Q_N(_1534_),
    .Q(\xq[1] ));
 sg13g2_dfrbp_1 \xq[2]$_SDFF_PP0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net214),
    .D(_0140_),
    .Q_N(_1533_),
    .Q(\xq[2] ));
 sg13g2_dfrbp_1 \xq[3]$_SDFF_PP0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net215),
    .D(_0141_),
    .Q_N(_1532_),
    .Q(\xq[3] ));
 sg13g2_dfrbp_1 \xq[4]$_SDFF_PP0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net216),
    .D(_0142_),
    .Q_N(_1531_),
    .Q(\xq[4] ));
 sg13g2_dfrbp_1 \xq[5]$_SDFF_PP0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net217),
    .D(_0143_),
    .Q_N(_1530_),
    .Q(\xq[5] ));
 sg13g2_dfrbp_1 \xq[6]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net218),
    .D(_0144_),
    .Q_N(_1529_),
    .Q(\xq[6] ));
 sg13g2_dfrbp_1 \xq[7]$_SDFF_PP0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net219),
    .D(_0145_),
    .Q_N(_1528_),
    .Q(\xq[7] ));
 sg13g2_dfrbp_1 \xq[8]$_SDFF_PP0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net220),
    .D(_0146_),
    .Q_N(_1527_),
    .Q(\xq[8] ));
 sg13g2_dfrbp_1 \xq[9]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net221),
    .D(_0147_),
    .Q_N(_1526_),
    .Q(\xq[9] ));
 sg13g2_dfrbp_1 \xqo[0]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net222),
    .D(_0148_),
    .Q_N(_1525_),
    .Q(\xqo[0] ));
 sg13g2_dfrbp_1 \xqo[10]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net223),
    .D(_0149_),
    .Q_N(_1524_),
    .Q(\xqo[10] ));
 sg13g2_dfrbp_1 \xqo[11]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net224),
    .D(_0150_),
    .Q_N(_1523_),
    .Q(\xqo[11] ));
 sg13g2_dfrbp_1 \xqo[1]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net225),
    .D(_0151_),
    .Q_N(_1522_),
    .Q(\xqo[1] ));
 sg13g2_dfrbp_1 \xqo[2]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net226),
    .D(_0152_),
    .Q_N(_1521_),
    .Q(\xqo[2] ));
 sg13g2_dfrbp_1 \xqo[3]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net227),
    .D(_0153_),
    .Q_N(_1520_),
    .Q(\xqo[3] ));
 sg13g2_dfrbp_1 \xqo[4]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net228),
    .D(_0154_),
    .Q_N(_1519_),
    .Q(\xqo[4] ));
 sg13g2_dfrbp_1 \xqo[5]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net229),
    .D(_0155_),
    .Q_N(_1518_),
    .Q(\xqo[5] ));
 sg13g2_dfrbp_1 \xqo[6]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net230),
    .D(_0156_),
    .Q_N(_0003_),
    .Q(\xqo[6] ));
 sg13g2_dfrbp_1 \xqo[7]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net231),
    .D(_0157_),
    .Q_N(_1517_),
    .Q(\xqo[7] ));
 sg13g2_dfrbp_1 \xqo[8]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net232),
    .D(_0158_),
    .Q_N(_1516_),
    .Q(\xqo[8] ));
 sg13g2_dfrbp_1 \xqo[9]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net233),
    .D(_0159_),
    .Q_N(_1515_),
    .Q(\xqo[9] ));
 sg13g2_dfrbp_1 \yq[0]$_SDFFE_PP0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net234),
    .D(_0160_),
    .Q_N(_1514_),
    .Q(\yq[0] ));
 sg13g2_dfrbp_1 \yq[10]$_SDFFE_PP0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net235),
    .D(_0161_),
    .Q_N(_1513_),
    .Q(\yq[10] ));
 sg13g2_dfrbp_1 \yq[11]$_SDFFE_PP0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net236),
    .D(_0162_),
    .Q_N(_1512_),
    .Q(\yq[11] ));
 sg13g2_dfrbp_1 \yq[12]$_SDFFE_PP0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net237),
    .D(_0163_),
    .Q_N(_1511_),
    .Q(\yq[12] ));
 sg13g2_dfrbp_1 \yq[1]$_SDFFE_PP0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net238),
    .D(_0164_),
    .Q_N(_1510_),
    .Q(\yq[1] ));
 sg13g2_dfrbp_1 \yq[2]$_SDFFE_PP0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net239),
    .D(_0165_),
    .Q_N(_1509_),
    .Q(\yq[2] ));
 sg13g2_dfrbp_1 \yq[3]$_SDFFE_PP0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net240),
    .D(_0166_),
    .Q_N(_1508_),
    .Q(\yq[3] ));
 sg13g2_dfrbp_1 \yq[4]$_SDFFE_PP0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net241),
    .D(_0167_),
    .Q_N(_1507_),
    .Q(\yq[4] ));
 sg13g2_dfrbp_1 \yq[5]$_SDFFE_PP0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net242),
    .D(_0168_),
    .Q_N(_1506_),
    .Q(\yq[5] ));
 sg13g2_dfrbp_1 \yq[6]$_SDFFE_PP0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net243),
    .D(_0169_),
    .Q_N(_1505_),
    .Q(\yq[6] ));
 sg13g2_dfrbp_1 \yq[7]$_SDFFE_PP0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net244),
    .D(_0170_),
    .Q_N(_1504_),
    .Q(\yq[7] ));
 sg13g2_dfrbp_1 \yq[8]$_SDFFE_PP0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net245),
    .D(_0171_),
    .Q_N(_1503_),
    .Q(\yq[8] ));
 sg13g2_dfrbp_1 \yq[9]$_SDFFE_PP0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net246),
    .D(_0172_),
    .Q_N(_1502_),
    .Q(\yq[9] ));
 sg13g2_dfrbp_1 \yqo[0]$_SDFFE_PP0N_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net247),
    .D(_0173_),
    .Q_N(_1501_),
    .Q(\yqo[0] ));
 sg13g2_dfrbp_1 \yqo[10]$_SDFFE_PP0N_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net248),
    .D(_0174_),
    .Q_N(_1500_),
    .Q(\yqo[10] ));
 sg13g2_dfrbp_1 \yqo[11]$_SDFFE_PP0N_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net249),
    .D(_0175_),
    .Q_N(_1499_),
    .Q(\yqo[11] ));
 sg13g2_dfrbp_1 \yqo[12]$_SDFFE_PP0N_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net250),
    .D(_0176_),
    .Q_N(_1498_),
    .Q(\yqo[12] ));
 sg13g2_dfrbp_1 \yqo[1]$_SDFFE_PP0N_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net251),
    .D(_0177_),
    .Q_N(_1497_),
    .Q(\yqo[1] ));
 sg13g2_dfrbp_1 \yqo[2]$_SDFFE_PP0N_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net252),
    .D(_0178_),
    .Q_N(_1496_),
    .Q(\yqo[2] ));
 sg13g2_dfrbp_1 \yqo[3]$_SDFFE_PP0N_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net253),
    .D(_0179_),
    .Q_N(_1495_),
    .Q(\yqo[3] ));
 sg13g2_dfrbp_1 \yqo[4]$_SDFFE_PP0N_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net254),
    .D(_0180_),
    .Q_N(_1494_),
    .Q(\yqo[4] ));
 sg13g2_dfrbp_1 \yqo[5]$_SDFFE_PP0N_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net255),
    .D(_0181_),
    .Q_N(_1493_),
    .Q(\yqo[5] ));
 sg13g2_dfrbp_1 \yqo[6]$_SDFFE_PP0N_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net256),
    .D(_0182_),
    .Q_N(_1492_),
    .Q(\yqo[6] ));
 sg13g2_dfrbp_1 \yqo[7]$_SDFFE_PP0N_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net257),
    .D(_0183_),
    .Q_N(_1491_),
    .Q(\yqo[7] ));
 sg13g2_dfrbp_1 \yqo[8]$_SDFFE_PP0N_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net258),
    .D(_0184_),
    .Q_N(_1490_),
    .Q(\yqo[8] ));
 sg13g2_dfrbp_1 \yqo[9]$_SDFFE_PP0N_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net259),
    .D(_0185_),
    .Q_N(_1489_),
    .Q(\yqo[9] ));
 sg13g2_buf_1 output1 (.A(net1),
    .X(uio_out[7]));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[3]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[4]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[5]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[6]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout10 (.A(_0822_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_0821_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_0588_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0204_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_0585_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_1454_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_1190_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0522_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0313_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0682_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0312_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_1432_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_1243_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_1094_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0669_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0587_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0583_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0484_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0463_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0433_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0410_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1430_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_1342_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1306_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1257_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0933_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0930_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0582_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0524_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0414_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0298_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1429_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1427_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1314_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1310_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1309_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1292_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1284_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1235_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0984_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0982_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0972_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0971_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0968_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0953_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0949_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0947_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0941_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0939_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0935_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0932_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0929_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0927_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0192_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1464_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1091_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0963_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0954_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0951_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0948_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0945_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0940_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0926_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0925_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(\hvsync_gen.vsync ),
    .X(net74));
 sg13g2_buf_1 fanout75 (.A(\hvsync_gen.vsync ),
    .X(net75));
 sg13g2_tielo _3123__76 (.L_LO(net76));
 sg13g2_tielo _3124__77 (.L_LO(net77));
 sg13g2_tielo _3125__78 (.L_LO(net78));
 sg13g2_tielo _3126__79 (.L_LO(net79));
 sg13g2_tielo _3127__80 (.L_LO(net80));
 sg13g2_tielo _3128__81 (.L_LO(net81));
 sg13g2_tielo _3129__82 (.L_LO(net82));
 sg13g2_tielo _3131__83 (.L_LO(net83));
 sg13g2_tielo _3132__84 (.L_LO(net84));
 sg13g2_tielo _3133__85 (.L_LO(net85));
 sg13g2_tielo _3134__86 (.L_LO(net86));
 sg13g2_tielo _3135__87 (.L_LO(net87));
 sg13g2_tielo _3136__88 (.L_LO(net88));
 sg13g2_tielo _3137__89 (.L_LO(net89));
 sg13g2_tiehi \LFSR[1]$_SDFF_PP0__91  (.L_HI(net91));
 sg13g2_tiehi \LFSR[2]$_SDFF_PP0__92  (.L_HI(net92));
 sg13g2_tiehi \LFSR[3]$_SDFF_PP0__93  (.L_HI(net93));
 sg13g2_tiehi \LFSR[4]$_SDFF_PP0__94  (.L_HI(net94));
 sg13g2_tiehi \LFSR[5]$_SDFF_PP0__95  (.L_HI(net95));
 sg13g2_tiehi \Voice1.accumulator[0]$_DFFE_PP__96  (.L_HI(net96));
 sg13g2_tiehi \Voice1.accumulator[10]$_DFFE_PP__97  (.L_HI(net97));
 sg13g2_tiehi \Voice1.accumulator[11]$_DFFE_PP__98  (.L_HI(net98));
 sg13g2_tiehi \Voice1.accumulator[12]$_DFFE_PP__99  (.L_HI(net99));
 sg13g2_tiehi \Voice1.accumulator[13]$_DFFE_PP__100  (.L_HI(net100));
 sg13g2_tiehi \Voice1.accumulator[14]$_DFFE_PP__101  (.L_HI(net101));
 sg13g2_tiehi \Voice1.accumulator[15]$_DFFE_PP__102  (.L_HI(net102));
 sg13g2_tiehi \Voice1.accumulator[16]$_DFFE_PP__103  (.L_HI(net103));
 sg13g2_tiehi \Voice1.accumulator[17]$_DFFE_PP__104  (.L_HI(net104));
 sg13g2_tiehi \Voice1.accumulator[18]$_DFFE_PP__105  (.L_HI(net105));
 sg13g2_tiehi \Voice1.accumulator[19]$_DFFE_PP__106  (.L_HI(net106));
 sg13g2_tiehi \Voice1.accumulator[1]$_DFFE_PP__107  (.L_HI(net107));
 sg13g2_tiehi \Voice1.accumulator[20]$_DFFE_PP__108  (.L_HI(net108));
 sg13g2_tiehi \Voice1.accumulator[21]$_DFFE_PP__109  (.L_HI(net109));
 sg13g2_tiehi \Voice1.accumulator[22]$_DFFE_PP__110  (.L_HI(net110));
 sg13g2_tiehi \Voice1.accumulator[23]$_DFFE_PP__111  (.L_HI(net111));
 sg13g2_tiehi \Voice1.accumulator[2]$_DFFE_PP__112  (.L_HI(net112));
 sg13g2_tiehi \Voice1.accumulator[3]$_DFFE_PP__113  (.L_HI(net113));
 sg13g2_tiehi \Voice1.accumulator[4]$_DFFE_PP__114  (.L_HI(net114));
 sg13g2_tiehi \Voice1.accumulator[5]$_DFFE_PP__115  (.L_HI(net115));
 sg13g2_tiehi \Voice1.accumulator[6]$_DFFE_PP__116  (.L_HI(net116));
 sg13g2_tiehi \Voice1.accumulator[7]$_DFFE_PP__117  (.L_HI(net117));
 sg13g2_tiehi \Voice1.accumulator[8]$_DFFE_PP__118  (.L_HI(net118));
 sg13g2_tiehi \Voice1.accumulator[9]$_DFFE_PP__119  (.L_HI(net119));
 sg13g2_tiehi \Voice1.pulse$_SDFFE_PN0P__120  (.L_HI(net120));
 sg13g2_tiehi _3130__121 (.L_HI(net121));
 sg13g2_tiehi \b[0]$_SDFF_PN0__122  (.L_HI(net122));
 sg13g2_tiehi \b[1]$_SDFF_PN0__123  (.L_HI(net123));
 sg13g2_tiehi \b[2]$_SDFF_PN0__124  (.L_HI(net124));
 sg13g2_tiehi \b[3]$_SDFF_PN0__125  (.L_HI(net125));
 sg13g2_tiehi \b[4]$_SDFF_PN0__126  (.L_HI(net126));
 sg13g2_tiehi \b[5]$_SDFF_PN0__127  (.L_HI(net127));
 sg13g2_tiehi \b[6]$_SDFF_PN0__128  (.L_HI(net128));
 sg13g2_tiehi \b[7]$_SDFF_PN0__129  (.L_HI(net129));
 sg13g2_tiehi \counter[0]$_SDFF_PN0__130  (.L_HI(net130));
 sg13g2_tiehi \counter[1]$_SDFF_PN0__131  (.L_HI(net131));
 sg13g2_tiehi \counter[2]$_SDFF_PN0__132  (.L_HI(net132));
 sg13g2_tiehi \counter[3]$_SDFF_PN0__133  (.L_HI(net133));
 sg13g2_tiehi \counter[4]$_SDFF_PN0__134  (.L_HI(net134));
 sg13g2_tiehi \counter[5]$_SDFF_PN0__135  (.L_HI(net135));
 sg13g2_tiehi \counter[6]$_SDFF_PN0__136  (.L_HI(net136));
 sg13g2_tiehi \counter[7]$_SDFF_PN0__137  (.L_HI(net137));
 sg13g2_tiehi \counter[8]$_SDFF_PN0__138  (.L_HI(net138));
 sg13g2_tiehi \ctr_audio[0]$_SDFFE_PN0P__139  (.L_HI(net139));
 sg13g2_tiehi \ctr_audio[10]$_SDFFE_PN0P__140  (.L_HI(net140));
 sg13g2_tiehi \ctr_audio[11]$_SDFFE_PN0P__141  (.L_HI(net141));
 sg13g2_tiehi \ctr_audio[12]$_SDFFE_PN0P__142  (.L_HI(net142));
 sg13g2_tiehi \ctr_audio[13]$_SDFFE_PN0P__143  (.L_HI(net143));
 sg13g2_tiehi \ctr_audio[14]$_SDFFE_PN0P__144  (.L_HI(net144));
 sg13g2_tiehi \ctr_audio[15]$_SDFFE_PN0P__145  (.L_HI(net145));
 sg13g2_tiehi \ctr_audio[16]$_SDFFE_PN0P__146  (.L_HI(net146));
 sg13g2_tiehi \ctr_audio[17]$_SDFFE_PN0P__147  (.L_HI(net147));
 sg13g2_tiehi \ctr_audio[18]$_SDFFE_PN0P__148  (.L_HI(net148));
 sg13g2_tiehi \ctr_audio[19]$_SDFFE_PN0P__149  (.L_HI(net149));
 sg13g2_tiehi \ctr_audio[1]$_SDFFE_PN0P__150  (.L_HI(net150));
 sg13g2_tiehi \ctr_audio[20]$_SDFFE_PN0P__151  (.L_HI(net151));
 sg13g2_tiehi \ctr_audio[21]$_SDFFE_PN0P__152  (.L_HI(net152));
 sg13g2_tiehi \ctr_audio[22]$_SDFFE_PN0P__153  (.L_HI(net153));
 sg13g2_tiehi \ctr_audio[23]$_SDFFE_PN0P__154  (.L_HI(net154));
 sg13g2_tiehi \ctr_audio[2]$_SDFFE_PN0P__155  (.L_HI(net155));
 sg13g2_tiehi \ctr_audio[3]$_SDFFE_PN0P__156  (.L_HI(net156));
 sg13g2_tiehi \ctr_audio[4]$_SDFFE_PN0P__157  (.L_HI(net157));
 sg13g2_tiehi \ctr_audio[5]$_SDFFE_PN0P__158  (.L_HI(net158));
 sg13g2_tiehi \ctr_audio[6]$_SDFFE_PN0P__159  (.L_HI(net159));
 sg13g2_tiehi \ctr_audio[7]$_SDFFE_PN0P__160  (.L_HI(net160));
 sg13g2_tiehi \ctr_audio[8]$_SDFFE_PN0P__161  (.L_HI(net161));
 sg13g2_tiehi \ctr_audio[9]$_SDFFE_PN0P__162  (.L_HI(net162));
 sg13g2_tiehi \ctr_clkdiv25[0]$_SDFF_PP0__163  (.L_HI(net163));
 sg13g2_tiehi \ctr_clkdiv25[1]$_SDFF_PP0__164  (.L_HI(net164));
 sg13g2_tiehi \ctr_clkdiv25[2]$_SDFF_PP0__165  (.L_HI(net165));
 sg13g2_tiehi \ctr_clkdiv25[3]$_SDFF_PP0__166  (.L_HI(net166));
 sg13g2_tiehi \ctr_clkdiv25[4]$_SDFF_PP0__167  (.L_HI(net167));
 sg13g2_tiehi \ctr_clkdiv25[5]$_SDFF_PP0__168  (.L_HI(net168));
 sg13g2_tiehi \ctr_clkdiv25[6]$_SDFF_PP0__169  (.L_HI(net169));
 sg13g2_tiehi \ctr_clkdiv25[7]$_SDFF_PP0__170  (.L_HI(net170));
 sg13g2_tiehi \g[0]$_SDFF_PN0__171  (.L_HI(net171));
 sg13g2_tiehi \g[1]$_SDFF_PN0__172  (.L_HI(net172));
 sg13g2_tiehi \g[2]$_SDFF_PN0__173  (.L_HI(net173));
 sg13g2_tiehi \g[3]$_SDFF_PN0__174  (.L_HI(net174));
 sg13g2_tiehi \g[4]$_SDFF_PN0__175  (.L_HI(net175));
 sg13g2_tiehi \g[5]$_SDFF_PN0__176  (.L_HI(net176));
 sg13g2_tiehi \g[6]$_SDFF_PN0__177  (.L_HI(net177));
 sg13g2_tiehi \g[7]$_SDFF_PN0__178  (.L_HI(net178));
 sg13g2_tiehi \hvsync_gen.hpos[0]$_SDFF_PP0__179  (.L_HI(net179));
 sg13g2_tiehi \hvsync_gen.hpos[1]$_SDFF_PP0__180  (.L_HI(net180));
 sg13g2_tiehi \hvsync_gen.hpos[2]$_SDFF_PP0__181  (.L_HI(net181));
 sg13g2_tiehi \hvsync_gen.hpos[3]$_SDFF_PP0__182  (.L_HI(net182));
 sg13g2_tiehi \hvsync_gen.hpos[4]$_SDFF_PP0__183  (.L_HI(net183));
 sg13g2_tiehi \hvsync_gen.hpos[5]$_SDFF_PP0__184  (.L_HI(net184));
 sg13g2_tiehi \hvsync_gen.hpos[6]$_SDFF_PP0__185  (.L_HI(net185));
 sg13g2_tiehi \hvsync_gen.hpos[7]$_SDFF_PP0__186  (.L_HI(net186));
 sg13g2_tiehi \hvsync_gen.hpos[8]$_SDFF_PP0__187  (.L_HI(net187));
 sg13g2_tiehi \hvsync_gen.hpos[9]$_SDFF_PP0__188  (.L_HI(net188));
 sg13g2_tiehi \hvsync_gen.hsync$_DFF_P__189  (.L_HI(net189));
 sg13g2_tiehi \hvsync_gen.vpos[0]$_SDFFCE_PP0P__190  (.L_HI(net190));
 sg13g2_tiehi \hvsync_gen.vpos[1]$_SDFFCE_PP0P__191  (.L_HI(net191));
 sg13g2_tiehi \hvsync_gen.vpos[2]$_SDFFCE_PP0P__192  (.L_HI(net192));
 sg13g2_tiehi \hvsync_gen.vpos[3]$_SDFFCE_PP0P__193  (.L_HI(net193));
 sg13g2_tiehi \hvsync_gen.vpos[4]$_SDFFCE_PP0P__194  (.L_HI(net194));
 sg13g2_tiehi \hvsync_gen.vpos[5]$_SDFFCE_PP0P__195  (.L_HI(net195));
 sg13g2_tiehi \hvsync_gen.vpos[6]$_SDFFCE_PP0P__196  (.L_HI(net196));
 sg13g2_tiehi \hvsync_gen.vpos[7]$_SDFFCE_PP0P__197  (.L_HI(net197));
 sg13g2_tiehi \hvsync_gen.vpos[8]$_SDFFCE_PP0P__198  (.L_HI(net198));
 sg13g2_tiehi \hvsync_gen.vpos[9]$_SDFFCE_PP0P__199  (.L_HI(net199));
 sg13g2_tiehi \hvsync_gen.vsync$_DFF_P__200  (.L_HI(net200));
 sg13g2_tiehi \pulse_1MHz$_SDFF_PN0__201  (.L_HI(net201));
 sg13g2_tiehi \r[0]$_SDFF_PN0__202  (.L_HI(net202));
 sg13g2_tiehi \r[1]$_SDFF_PN0__203  (.L_HI(net203));
 sg13g2_tiehi \r[2]$_SDFF_PN0__204  (.L_HI(net204));
 sg13g2_tiehi \r[3]$_SDFF_PN0__205  (.L_HI(net205));
 sg13g2_tiehi \r[4]$_SDFF_PN0__206  (.L_HI(net206));
 sg13g2_tiehi \r[5]$_SDFF_PN0__207  (.L_HI(net207));
 sg13g2_tiehi \r[6]$_SDFF_PN0__208  (.L_HI(net208));
 sg13g2_tiehi \r[7]$_SDFF_PN0__209  (.L_HI(net209));
 sg13g2_tiehi \xq[0]$_SDFF_PP0__210  (.L_HI(net210));
 sg13g2_tiehi \xq[10]$_SDFF_PP0__211  (.L_HI(net211));
 sg13g2_tiehi \xq[11]$_SDFF_PP0__212  (.L_HI(net212));
 sg13g2_tiehi \xq[1]$_SDFF_PP0__213  (.L_HI(net213));
 sg13g2_tiehi \xq[2]$_SDFF_PP0__214  (.L_HI(net214));
 sg13g2_tiehi \xq[3]$_SDFF_PP0__215  (.L_HI(net215));
 sg13g2_tiehi \xq[4]$_SDFF_PP0__216  (.L_HI(net216));
 sg13g2_tiehi \xq[5]$_SDFF_PP0__217  (.L_HI(net217));
 sg13g2_tiehi \xq[6]$_SDFF_PP0__218  (.L_HI(net218));
 sg13g2_tiehi \xq[7]$_SDFF_PP0__219  (.L_HI(net219));
 sg13g2_tiehi \xq[8]$_SDFF_PP0__220  (.L_HI(net220));
 sg13g2_tiehi \xq[9]$_SDFF_PP0__221  (.L_HI(net221));
 sg13g2_tiehi \xqo[0]$_SDFF_PN0__222  (.L_HI(net222));
 sg13g2_tiehi \xqo[10]$_SDFF_PN0__223  (.L_HI(net223));
 sg13g2_tiehi \xqo[11]$_SDFF_PN0__224  (.L_HI(net224));
 sg13g2_tiehi \xqo[1]$_SDFF_PN0__225  (.L_HI(net225));
 sg13g2_tiehi \xqo[2]$_SDFF_PN0__226  (.L_HI(net226));
 sg13g2_tiehi \xqo[3]$_SDFF_PN0__227  (.L_HI(net227));
 sg13g2_tiehi \xqo[4]$_SDFF_PN0__228  (.L_HI(net228));
 sg13g2_tiehi \xqo[5]$_SDFF_PN0__229  (.L_HI(net229));
 sg13g2_tiehi \xqo[6]$_SDFF_PN0__230  (.L_HI(net230));
 sg13g2_tiehi \xqo[7]$_SDFF_PN0__231  (.L_HI(net231));
 sg13g2_tiehi \xqo[8]$_SDFF_PN0__232  (.L_HI(net232));
 sg13g2_tiehi \xqo[9]$_SDFF_PN0__233  (.L_HI(net233));
 sg13g2_tiehi \yq[0]$_SDFFE_PP0P__234  (.L_HI(net234));
 sg13g2_tiehi \yq[10]$_SDFFE_PP0P__235  (.L_HI(net235));
 sg13g2_tiehi \yq[11]$_SDFFE_PP0P__236  (.L_HI(net236));
 sg13g2_tiehi \yq[12]$_SDFFE_PP0P__237  (.L_HI(net237));
 sg13g2_tiehi \yq[1]$_SDFFE_PP0P__238  (.L_HI(net238));
 sg13g2_tiehi \yq[2]$_SDFFE_PP0P__239  (.L_HI(net239));
 sg13g2_tiehi \yq[3]$_SDFFE_PP0P__240  (.L_HI(net240));
 sg13g2_tiehi \yq[4]$_SDFFE_PP0P__241  (.L_HI(net241));
 sg13g2_tiehi \yq[5]$_SDFFE_PP0P__242  (.L_HI(net242));
 sg13g2_tiehi \yq[6]$_SDFFE_PP0P__243  (.L_HI(net243));
 sg13g2_tiehi \yq[7]$_SDFFE_PP0P__244  (.L_HI(net244));
 sg13g2_tiehi \yq[8]$_SDFFE_PP0P__245  (.L_HI(net245));
 sg13g2_tiehi \yq[9]$_SDFFE_PP0P__246  (.L_HI(net246));
 sg13g2_tiehi \yqo[0]$_SDFFE_PP0N__247  (.L_HI(net247));
 sg13g2_tiehi \yqo[10]$_SDFFE_PP0N__248  (.L_HI(net248));
 sg13g2_tiehi \yqo[11]$_SDFFE_PP0N__249  (.L_HI(net249));
 sg13g2_tiehi \yqo[12]$_SDFFE_PP0N__250  (.L_HI(net250));
 sg13g2_tiehi \yqo[1]$_SDFFE_PP0N__251  (.L_HI(net251));
 sg13g2_tiehi \yqo[2]$_SDFFE_PP0N__252  (.L_HI(net252));
 sg13g2_tiehi \yqo[3]$_SDFFE_PP0N__253  (.L_HI(net253));
 sg13g2_tiehi \yqo[4]$_SDFFE_PP0N__254  (.L_HI(net254));
 sg13g2_tiehi \yqo[5]$_SDFFE_PP0N__255  (.L_HI(net255));
 sg13g2_tiehi \yqo[6]$_SDFFE_PP0N__256  (.L_HI(net256));
 sg13g2_tiehi \yqo[7]$_SDFFE_PP0N__257  (.L_HI(net257));
 sg13g2_tiehi \yqo[8]$_SDFFE_PP0N__258  (.L_HI(net258));
 sg13g2_tiehi \yqo[9]$_SDFFE_PP0N__259  (.L_HI(net259));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_fill_2 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_decap_8 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_297 ();
 sg13g2_decap_8 FILLER_17_304 ();
 sg13g2_decap_8 FILLER_17_311 ();
 sg13g2_decap_8 FILLER_17_318 ();
 sg13g2_decap_8 FILLER_17_325 ();
 sg13g2_decap_8 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_17_409 ();
 sg13g2_decap_8 FILLER_17_416 ();
 sg13g2_decap_8 FILLER_17_423 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_4 FILLER_18_224 ();
 sg13g2_fill_2 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_fill_2 FILLER_18_427 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_4 FILLER_19_217 ();
 sg13g2_fill_2 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_254 ();
 sg13g2_fill_2 FILLER_19_261 ();
 sg13g2_fill_1 FILLER_19_303 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_4 FILLER_19_315 ();
 sg13g2_fill_2 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_8 FILLER_19_403 ();
 sg13g2_decap_8 FILLER_19_410 ();
 sg13g2_decap_8 FILLER_19_417 ();
 sg13g2_decap_4 FILLER_19_424 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_4 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_243 ();
 sg13g2_decap_4 FILLER_20_248 ();
 sg13g2_fill_1 FILLER_20_252 ();
 sg13g2_fill_2 FILLER_20_322 ();
 sg13g2_fill_1 FILLER_20_328 ();
 sg13g2_fill_2 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_366 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_decap_8 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_20_415 ();
 sg13g2_decap_8 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_253 ();
 sg13g2_decap_8 FILLER_21_264 ();
 sg13g2_decap_4 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_275 ();
 sg13g2_decap_8 FILLER_21_282 ();
 sg13g2_fill_2 FILLER_21_289 ();
 sg13g2_fill_1 FILLER_21_291 ();
 sg13g2_decap_4 FILLER_21_331 ();
 sg13g2_fill_1 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_353 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_decap_8 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_21_414 ();
 sg13g2_decap_8 FILLER_21_421 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_4 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_4 FILLER_22_295 ();
 sg13g2_fill_1 FILLER_22_304 ();
 sg13g2_fill_2 FILLER_22_310 ();
 sg13g2_fill_2 FILLER_22_316 ();
 sg13g2_fill_2 FILLER_22_344 ();
 sg13g2_fill_1 FILLER_22_346 ();
 sg13g2_decap_8 FILLER_22_373 ();
 sg13g2_decap_8 FILLER_22_380 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_decap_8 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_22_415 ();
 sg13g2_decap_8 FILLER_22_422 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_4 FILLER_23_98 ();
 sg13g2_fill_2 FILLER_23_102 ();
 sg13g2_decap_8 FILLER_23_108 ();
 sg13g2_decap_8 FILLER_23_115 ();
 sg13g2_decap_8 FILLER_23_122 ();
 sg13g2_decap_8 FILLER_23_129 ();
 sg13g2_decap_8 FILLER_23_136 ();
 sg13g2_decap_8 FILLER_23_143 ();
 sg13g2_decap_8 FILLER_23_150 ();
 sg13g2_decap_8 FILLER_23_157 ();
 sg13g2_decap_8 FILLER_23_164 ();
 sg13g2_decap_8 FILLER_23_171 ();
 sg13g2_decap_8 FILLER_23_178 ();
 sg13g2_decap_8 FILLER_23_185 ();
 sg13g2_decap_8 FILLER_23_192 ();
 sg13g2_decap_8 FILLER_23_199 ();
 sg13g2_fill_1 FILLER_23_206 ();
 sg13g2_fill_1 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_216 ();
 sg13g2_fill_1 FILLER_23_243 ();
 sg13g2_fill_1 FILLER_23_249 ();
 sg13g2_fill_1 FILLER_23_258 ();
 sg13g2_fill_1 FILLER_23_302 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_346 ();
 sg13g2_fill_1 FILLER_23_353 ();
 sg13g2_fill_2 FILLER_23_358 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_fill_2 FILLER_23_365 ();
 sg13g2_fill_1 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_decap_8 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_23_414 ();
 sg13g2_decap_8 FILLER_23_421 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_4 FILLER_24_91 ();
 sg13g2_fill_2 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_123 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_decap_8 FILLER_24_137 ();
 sg13g2_decap_8 FILLER_24_144 ();
 sg13g2_decap_8 FILLER_24_151 ();
 sg13g2_decap_8 FILLER_24_158 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_172 ();
 sg13g2_decap_8 FILLER_24_179 ();
 sg13g2_decap_8 FILLER_24_186 ();
 sg13g2_decap_8 FILLER_24_193 ();
 sg13g2_fill_1 FILLER_24_265 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_decap_4 FILLER_24_300 ();
 sg13g2_decap_4 FILLER_24_311 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_fill_2 FILLER_24_322 ();
 sg13g2_fill_1 FILLER_24_324 ();
 sg13g2_fill_2 FILLER_24_341 ();
 sg13g2_fill_1 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_8 FILLER_24_403 ();
 sg13g2_decap_8 FILLER_24_410 ();
 sg13g2_decap_8 FILLER_24_417 ();
 sg13g2_decap_4 FILLER_24_424 ();
 sg13g2_fill_2 FILLER_24_428 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_103 ();
 sg13g2_decap_8 FILLER_25_110 ();
 sg13g2_fill_2 FILLER_25_122 ();
 sg13g2_fill_1 FILLER_25_124 ();
 sg13g2_decap_8 FILLER_25_129 ();
 sg13g2_decap_8 FILLER_25_136 ();
 sg13g2_decap_8 FILLER_25_143 ();
 sg13g2_decap_8 FILLER_25_150 ();
 sg13g2_decap_8 FILLER_25_157 ();
 sg13g2_decap_8 FILLER_25_164 ();
 sg13g2_decap_8 FILLER_25_171 ();
 sg13g2_decap_4 FILLER_25_178 ();
 sg13g2_fill_2 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_188 ();
 sg13g2_decap_8 FILLER_25_195 ();
 sg13g2_decap_8 FILLER_25_202 ();
 sg13g2_decap_8 FILLER_25_209 ();
 sg13g2_decap_8 FILLER_25_216 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_decap_8 FILLER_25_254 ();
 sg13g2_decap_8 FILLER_25_261 ();
 sg13g2_decap_4 FILLER_25_268 ();
 sg13g2_fill_2 FILLER_25_272 ();
 sg13g2_fill_1 FILLER_25_309 ();
 sg13g2_decap_8 FILLER_25_327 ();
 sg13g2_fill_2 FILLER_25_334 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_366 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_380 ();
 sg13g2_decap_8 FILLER_25_387 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_decap_8 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_25_415 ();
 sg13g2_decap_8 FILLER_25_422 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_fill_2 FILLER_26_106 ();
 sg13g2_decap_8 FILLER_26_146 ();
 sg13g2_decap_8 FILLER_26_153 ();
 sg13g2_decap_8 FILLER_26_160 ();
 sg13g2_decap_8 FILLER_26_167 ();
 sg13g2_decap_8 FILLER_26_174 ();
 sg13g2_decap_8 FILLER_26_181 ();
 sg13g2_decap_8 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_195 ();
 sg13g2_decap_8 FILLER_26_202 ();
 sg13g2_decap_8 FILLER_26_209 ();
 sg13g2_fill_1 FILLER_26_216 ();
 sg13g2_decap_8 FILLER_26_225 ();
 sg13g2_decap_8 FILLER_26_237 ();
 sg13g2_decap_8 FILLER_26_244 ();
 sg13g2_decap_8 FILLER_26_251 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_fill_2 FILLER_26_294 ();
 sg13g2_decap_4 FILLER_26_326 ();
 sg13g2_fill_2 FILLER_26_338 ();
 sg13g2_decap_4 FILLER_26_348 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_fill_2 FILLER_26_427 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_4 FILLER_27_84 ();
 sg13g2_fill_1 FILLER_27_88 ();
 sg13g2_decap_4 FILLER_27_93 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_fill_2 FILLER_27_115 ();
 sg13g2_fill_2 FILLER_27_122 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_fill_2 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_195 ();
 sg13g2_decap_8 FILLER_27_202 ();
 sg13g2_fill_2 FILLER_27_209 ();
 sg13g2_fill_1 FILLER_27_211 ();
 sg13g2_decap_8 FILLER_27_228 ();
 sg13g2_decap_8 FILLER_27_239 ();
 sg13g2_decap_8 FILLER_27_246 ();
 sg13g2_decap_8 FILLER_27_253 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_decap_8 FILLER_27_274 ();
 sg13g2_decap_8 FILLER_27_281 ();
 sg13g2_decap_8 FILLER_27_288 ();
 sg13g2_decap_8 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_decap_8 FILLER_27_309 ();
 sg13g2_decap_8 FILLER_27_316 ();
 sg13g2_fill_2 FILLER_27_323 ();
 sg13g2_fill_1 FILLER_27_325 ();
 sg13g2_fill_2 FILLER_27_341 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_decap_8 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_27_415 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_4 FILLER_28_77 ();
 sg13g2_decap_4 FILLER_28_118 ();
 sg13g2_decap_4 FILLER_28_130 ();
 sg13g2_fill_1 FILLER_28_134 ();
 sg13g2_decap_8 FILLER_28_139 ();
 sg13g2_decap_8 FILLER_28_146 ();
 sg13g2_decap_8 FILLER_28_153 ();
 sg13g2_decap_8 FILLER_28_160 ();
 sg13g2_decap_8 FILLER_28_167 ();
 sg13g2_decap_8 FILLER_28_174 ();
 sg13g2_decap_8 FILLER_28_181 ();
 sg13g2_decap_8 FILLER_28_188 ();
 sg13g2_decap_8 FILLER_28_195 ();
 sg13g2_decap_8 FILLER_28_202 ();
 sg13g2_fill_1 FILLER_28_209 ();
 sg13g2_fill_2 FILLER_28_219 ();
 sg13g2_fill_1 FILLER_28_221 ();
 sg13g2_fill_1 FILLER_28_227 ();
 sg13g2_decap_4 FILLER_28_238 ();
 sg13g2_fill_1 FILLER_28_242 ();
 sg13g2_decap_4 FILLER_28_252 ();
 sg13g2_fill_1 FILLER_28_256 ();
 sg13g2_decap_8 FILLER_28_272 ();
 sg13g2_fill_2 FILLER_28_279 ();
 sg13g2_decap_8 FILLER_28_307 ();
 sg13g2_decap_8 FILLER_28_314 ();
 sg13g2_decap_4 FILLER_28_321 ();
 sg13g2_fill_1 FILLER_28_325 ();
 sg13g2_decap_8 FILLER_28_365 ();
 sg13g2_decap_8 FILLER_28_372 ();
 sg13g2_fill_2 FILLER_28_379 ();
 sg13g2_fill_1 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_420 ();
 sg13g2_fill_2 FILLER_28_427 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_118 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_fill_1 FILLER_29_130 ();
 sg13g2_decap_8 FILLER_29_139 ();
 sg13g2_decap_8 FILLER_29_146 ();
 sg13g2_decap_8 FILLER_29_153 ();
 sg13g2_decap_8 FILLER_29_160 ();
 sg13g2_decap_8 FILLER_29_167 ();
 sg13g2_decap_8 FILLER_29_174 ();
 sg13g2_decap_4 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_fill_1 FILLER_29_206 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_4 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_234 ();
 sg13g2_fill_2 FILLER_29_241 ();
 sg13g2_fill_1 FILLER_29_243 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_fill_1 FILLER_29_257 ();
 sg13g2_decap_4 FILLER_29_276 ();
 sg13g2_fill_2 FILLER_29_285 ();
 sg13g2_fill_1 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_292 ();
 sg13g2_decap_4 FILLER_29_299 ();
 sg13g2_fill_1 FILLER_29_303 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_decap_8 FILLER_29_320 ();
 sg13g2_fill_2 FILLER_29_327 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_decap_4 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_29_375 ();
 sg13g2_decap_4 FILLER_29_382 ();
 sg13g2_fill_2 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_fill_2 FILLER_29_427 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_decap_4 FILLER_30_97 ();
 sg13g2_decap_8 FILLER_30_104 ();
 sg13g2_decap_4 FILLER_30_123 ();
 sg13g2_fill_2 FILLER_30_127 ();
 sg13g2_fill_2 FILLER_30_152 ();
 sg13g2_fill_1 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_160 ();
 sg13g2_decap_8 FILLER_30_167 ();
 sg13g2_decap_8 FILLER_30_174 ();
 sg13g2_decap_4 FILLER_30_181 ();
 sg13g2_decap_8 FILLER_30_204 ();
 sg13g2_decap_4 FILLER_30_226 ();
 sg13g2_fill_1 FILLER_30_230 ();
 sg13g2_decap_4 FILLER_30_236 ();
 sg13g2_fill_1 FILLER_30_259 ();
 sg13g2_fill_1 FILLER_30_264 ();
 sg13g2_fill_2 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_287 ();
 sg13g2_decap_4 FILLER_30_293 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_decap_4 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_338 ();
 sg13g2_decap_8 FILLER_30_345 ();
 sg13g2_decap_8 FILLER_30_352 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_8 FILLER_30_405 ();
 sg13g2_decap_4 FILLER_30_412 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_4 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_88 ();
 sg13g2_fill_1 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_fill_1 FILLER_31_182 ();
 sg13g2_fill_1 FILLER_31_218 ();
 sg13g2_fill_1 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_255 ();
 sg13g2_fill_1 FILLER_31_291 ();
 sg13g2_decap_4 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_4 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_361 ();
 sg13g2_decap_4 FILLER_31_373 ();
 sg13g2_fill_1 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_decap_4 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_4 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_88 ();
 sg13g2_decap_4 FILLER_32_120 ();
 sg13g2_fill_2 FILLER_32_153 ();
 sg13g2_decap_8 FILLER_32_159 ();
 sg13g2_decap_8 FILLER_32_166 ();
 sg13g2_decap_8 FILLER_32_173 ();
 sg13g2_decap_8 FILLER_32_180 ();
 sg13g2_decap_8 FILLER_32_187 ();
 sg13g2_decap_8 FILLER_32_194 ();
 sg13g2_decap_4 FILLER_32_201 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_4 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_244 ();
 sg13g2_decap_8 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_fill_1 FILLER_32_263 ();
 sg13g2_fill_2 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_281 ();
 sg13g2_decap_4 FILLER_32_300 ();
 sg13g2_fill_2 FILLER_32_304 ();
 sg13g2_decap_8 FILLER_32_323 ();
 sg13g2_fill_2 FILLER_32_348 ();
 sg13g2_fill_1 FILLER_32_350 ();
 sg13g2_fill_2 FILLER_32_377 ();
 sg13g2_fill_2 FILLER_32_383 ();
 sg13g2_fill_2 FILLER_32_389 ();
 sg13g2_fill_2 FILLER_32_400 ();
 sg13g2_fill_1 FILLER_32_402 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_104 ();
 sg13g2_decap_8 FILLER_33_111 ();
 sg13g2_fill_1 FILLER_33_118 ();
 sg13g2_decap_8 FILLER_33_132 ();
 sg13g2_decap_8 FILLER_33_139 ();
 sg13g2_decap_8 FILLER_33_146 ();
 sg13g2_decap_8 FILLER_33_153 ();
 sg13g2_decap_8 FILLER_33_160 ();
 sg13g2_decap_8 FILLER_33_167 ();
 sg13g2_decap_4 FILLER_33_174 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_decap_8 FILLER_33_188 ();
 sg13g2_decap_4 FILLER_33_195 ();
 sg13g2_fill_2 FILLER_33_199 ();
 sg13g2_decap_4 FILLER_33_211 ();
 sg13g2_fill_2 FILLER_33_215 ();
 sg13g2_decap_8 FILLER_33_222 ();
 sg13g2_decap_8 FILLER_33_229 ();
 sg13g2_decap_8 FILLER_33_236 ();
 sg13g2_fill_2 FILLER_33_243 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_decap_4 FILLER_33_260 ();
 sg13g2_fill_1 FILLER_33_264 ();
 sg13g2_decap_4 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_277 ();
 sg13g2_fill_2 FILLER_33_283 ();
 sg13g2_fill_1 FILLER_33_285 ();
 sg13g2_decap_8 FILLER_33_299 ();
 sg13g2_fill_2 FILLER_33_306 ();
 sg13g2_decap_4 FILLER_33_329 ();
 sg13g2_fill_2 FILLER_33_333 ();
 sg13g2_fill_2 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_fill_2 FILLER_33_355 ();
 sg13g2_fill_1 FILLER_33_357 ();
 sg13g2_fill_2 FILLER_33_362 ();
 sg13g2_fill_2 FILLER_33_369 ();
 sg13g2_fill_2 FILLER_33_375 ();
 sg13g2_fill_1 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_fill_1 FILLER_33_409 ();
 sg13g2_fill_2 FILLER_33_414 ();
 sg13g2_fill_2 FILLER_33_420 ();
 sg13g2_decap_4 FILLER_33_426 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_177 ();
 sg13g2_decap_4 FILLER_34_184 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_decap_8 FILLER_34_232 ();
 sg13g2_fill_2 FILLER_34_239 ();
 sg13g2_decap_4 FILLER_34_249 ();
 sg13g2_decap_8 FILLER_34_263 ();
 sg13g2_decap_8 FILLER_34_270 ();
 sg13g2_decap_8 FILLER_34_277 ();
 sg13g2_decap_8 FILLER_34_297 ();
 sg13g2_decap_8 FILLER_34_304 ();
 sg13g2_decap_4 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_328 ();
 sg13g2_fill_2 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_348 ();
 sg13g2_decap_8 FILLER_34_355 ();
 sg13g2_decap_4 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_4 FILLER_34_387 ();
 sg13g2_fill_2 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_2 FILLER_34_412 ();
 sg13g2_decap_8 FILLER_34_419 ();
 sg13g2_decap_4 FILLER_34_426 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_4 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_88 ();
 sg13g2_decap_8 FILLER_35_116 ();
 sg13g2_decap_8 FILLER_35_132 ();
 sg13g2_decap_8 FILLER_35_139 ();
 sg13g2_fill_1 FILLER_35_146 ();
 sg13g2_fill_1 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_176 ();
 sg13g2_fill_2 FILLER_35_195 ();
 sg13g2_fill_2 FILLER_35_202 ();
 sg13g2_fill_1 FILLER_35_216 ();
 sg13g2_fill_1 FILLER_35_222 ();
 sg13g2_fill_1 FILLER_35_237 ();
 sg13g2_fill_1 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_265 ();
 sg13g2_decap_8 FILLER_35_272 ();
 sg13g2_decap_8 FILLER_35_279 ();
 sg13g2_decap_4 FILLER_35_286 ();
 sg13g2_fill_2 FILLER_35_290 ();
 sg13g2_decap_8 FILLER_35_300 ();
 sg13g2_decap_8 FILLER_35_307 ();
 sg13g2_decap_4 FILLER_35_314 ();
 sg13g2_fill_1 FILLER_35_318 ();
 sg13g2_decap_8 FILLER_35_351 ();
 sg13g2_decap_8 FILLER_35_358 ();
 sg13g2_fill_2 FILLER_35_391 ();
 sg13g2_fill_1 FILLER_35_397 ();
 sg13g2_decap_8 FILLER_35_412 ();
 sg13g2_decap_8 FILLER_35_419 ();
 sg13g2_decap_4 FILLER_35_426 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_4 FILLER_36_56 ();
 sg13g2_decap_4 FILLER_36_90 ();
 sg13g2_fill_1 FILLER_36_94 ();
 sg13g2_fill_1 FILLER_36_103 ();
 sg13g2_fill_2 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_114 ();
 sg13g2_fill_2 FILLER_36_182 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_fill_2 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_4 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_264 ();
 sg13g2_decap_8 FILLER_36_274 ();
 sg13g2_decap_8 FILLER_36_281 ();
 sg13g2_decap_8 FILLER_36_288 ();
 sg13g2_decap_8 FILLER_36_295 ();
 sg13g2_decap_4 FILLER_36_302 ();
 sg13g2_decap_8 FILLER_36_319 ();
 sg13g2_fill_2 FILLER_36_326 ();
 sg13g2_fill_1 FILLER_36_328 ();
 sg13g2_fill_2 FILLER_36_382 ();
 sg13g2_fill_1 FILLER_36_384 ();
 sg13g2_fill_1 FILLER_36_398 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_fill_2 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_41 ();
 sg13g2_decap_8 FILLER_37_48 ();
 sg13g2_fill_2 FILLER_37_55 ();
 sg13g2_fill_1 FILLER_37_65 ();
 sg13g2_decap_8 FILLER_37_78 ();
 sg13g2_decap_8 FILLER_37_85 ();
 sg13g2_decap_4 FILLER_37_96 ();
 sg13g2_decap_4 FILLER_37_104 ();
 sg13g2_fill_2 FILLER_37_108 ();
 sg13g2_decap_4 FILLER_37_118 ();
 sg13g2_fill_1 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_179 ();
 sg13g2_decap_8 FILLER_37_186 ();
 sg13g2_decap_8 FILLER_37_198 ();
 sg13g2_decap_4 FILLER_37_205 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_4 FILLER_37_231 ();
 sg13g2_fill_2 FILLER_37_235 ();
 sg13g2_decap_4 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_246 ();
 sg13g2_fill_1 FILLER_37_295 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_4 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_fill_1 FILLER_37_329 ();
 sg13g2_fill_2 FILLER_37_334 ();
 sg13g2_fill_1 FILLER_37_336 ();
 sg13g2_fill_2 FILLER_37_363 ();
 sg13g2_fill_1 FILLER_37_365 ();
 sg13g2_fill_1 FILLER_37_371 ();
 sg13g2_fill_1 FILLER_37_377 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_fill_1 FILLER_37_387 ();
 sg13g2_decap_4 FILLER_37_393 ();
 sg13g2_fill_2 FILLER_37_397 ();
 sg13g2_fill_1 FILLER_37_416 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_82 ();
 sg13g2_fill_1 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_122 ();
 sg13g2_fill_1 FILLER_38_128 ();
 sg13g2_decap_4 FILLER_38_155 ();
 sg13g2_fill_2 FILLER_38_159 ();
 sg13g2_decap_8 FILLER_38_173 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_256 ();
 sg13g2_fill_1 FILLER_38_284 ();
 sg13g2_decap_4 FILLER_38_302 ();
 sg13g2_fill_2 FILLER_38_306 ();
 sg13g2_decap_4 FILLER_38_323 ();
 sg13g2_fill_2 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_337 ();
 sg13g2_decap_8 FILLER_38_352 ();
 sg13g2_fill_2 FILLER_38_359 ();
 sg13g2_decap_8 FILLER_38_365 ();
 sg13g2_decap_4 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_fill_2 FILLER_38_427 ();
 sg13g2_fill_1 FILLER_38_429 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_83 ();
 sg13g2_decap_8 FILLER_39_90 ();
 sg13g2_fill_1 FILLER_39_97 ();
 sg13g2_decap_8 FILLER_39_118 ();
 sg13g2_decap_8 FILLER_39_125 ();
 sg13g2_decap_8 FILLER_39_132 ();
 sg13g2_decap_8 FILLER_39_139 ();
 sg13g2_decap_4 FILLER_39_146 ();
 sg13g2_fill_1 FILLER_39_150 ();
 sg13g2_fill_1 FILLER_39_159 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_fill_1 FILLER_39_182 ();
 sg13g2_fill_2 FILLER_39_188 ();
 sg13g2_fill_1 FILLER_39_190 ();
 sg13g2_fill_1 FILLER_39_231 ();
 sg13g2_decap_4 FILLER_39_236 ();
 sg13g2_fill_2 FILLER_39_240 ();
 sg13g2_fill_2 FILLER_39_258 ();
 sg13g2_fill_1 FILLER_39_260 ();
 sg13g2_fill_1 FILLER_39_266 ();
 sg13g2_fill_2 FILLER_39_310 ();
 sg13g2_fill_2 FILLER_39_322 ();
 sg13g2_decap_8 FILLER_39_351 ();
 sg13g2_decap_8 FILLER_39_358 ();
 sg13g2_decap_8 FILLER_39_365 ();
 sg13g2_decap_8 FILLER_39_372 ();
 sg13g2_fill_1 FILLER_39_379 ();
 sg13g2_decap_4 FILLER_39_399 ();
 sg13g2_fill_2 FILLER_39_403 ();
 sg13g2_decap_8 FILLER_39_410 ();
 sg13g2_decap_8 FILLER_39_417 ();
 sg13g2_decap_4 FILLER_39_424 ();
 sg13g2_fill_2 FILLER_39_428 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_fill_1 FILLER_40_67 ();
 sg13g2_fill_1 FILLER_40_98 ();
 sg13g2_decap_4 FILLER_40_129 ();
 sg13g2_fill_1 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_146 ();
 sg13g2_decap_8 FILLER_40_153 ();
 sg13g2_fill_1 FILLER_40_160 ();
 sg13g2_decap_8 FILLER_40_171 ();
 sg13g2_fill_1 FILLER_40_193 ();
 sg13g2_fill_1 FILLER_40_226 ();
 sg13g2_fill_1 FILLER_40_237 ();
 sg13g2_decap_8 FILLER_40_242 ();
 sg13g2_fill_2 FILLER_40_249 ();
 sg13g2_fill_1 FILLER_40_251 ();
 sg13g2_fill_1 FILLER_40_257 ();
 sg13g2_fill_2 FILLER_40_283 ();
 sg13g2_decap_8 FILLER_40_305 ();
 sg13g2_decap_4 FILLER_40_312 ();
 sg13g2_fill_2 FILLER_40_321 ();
 sg13g2_fill_1 FILLER_40_328 ();
 sg13g2_decap_4 FILLER_40_333 ();
 sg13g2_fill_2 FILLER_40_346 ();
 sg13g2_decap_8 FILLER_40_353 ();
 sg13g2_decap_4 FILLER_40_360 ();
 sg13g2_fill_2 FILLER_40_364 ();
 sg13g2_fill_2 FILLER_40_376 ();
 sg13g2_fill_1 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_4 FILLER_41_21 ();
 sg13g2_fill_2 FILLER_41_25 ();
 sg13g2_decap_8 FILLER_41_31 ();
 sg13g2_decap_8 FILLER_41_38 ();
 sg13g2_decap_8 FILLER_41_45 ();
 sg13g2_decap_4 FILLER_41_52 ();
 sg13g2_fill_1 FILLER_41_56 ();
 sg13g2_fill_2 FILLER_41_63 ();
 sg13g2_fill_2 FILLER_41_72 ();
 sg13g2_fill_1 FILLER_41_74 ();
 sg13g2_decap_8 FILLER_41_79 ();
 sg13g2_decap_8 FILLER_41_86 ();
 sg13g2_fill_2 FILLER_41_93 ();
 sg13g2_decap_8 FILLER_41_99 ();
 sg13g2_fill_2 FILLER_41_106 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_fill_2 FILLER_41_119 ();
 sg13g2_decap_4 FILLER_41_147 ();
 sg13g2_fill_2 FILLER_41_156 ();
 sg13g2_fill_1 FILLER_41_158 ();
 sg13g2_decap_4 FILLER_41_168 ();
 sg13g2_fill_2 FILLER_41_172 ();
 sg13g2_fill_2 FILLER_41_184 ();
 sg13g2_decap_8 FILLER_41_232 ();
 sg13g2_fill_2 FILLER_41_239 ();
 sg13g2_fill_1 FILLER_41_254 ();
 sg13g2_fill_1 FILLER_41_263 ();
 sg13g2_fill_1 FILLER_41_269 ();
 sg13g2_fill_1 FILLER_41_276 ();
 sg13g2_decap_4 FILLER_41_293 ();
 sg13g2_fill_2 FILLER_41_301 ();
 sg13g2_fill_1 FILLER_41_303 ();
 sg13g2_decap_8 FILLER_41_421 ();
 sg13g2_fill_2 FILLER_41_428 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_4 FILLER_42_28 ();
 sg13g2_fill_1 FILLER_42_32 ();
 sg13g2_fill_1 FILLER_42_37 ();
 sg13g2_fill_1 FILLER_42_59 ();
 sg13g2_decap_8 FILLER_42_66 ();
 sg13g2_fill_1 FILLER_42_73 ();
 sg13g2_decap_8 FILLER_42_80 ();
 sg13g2_decap_8 FILLER_42_87 ();
 sg13g2_decap_8 FILLER_42_94 ();
 sg13g2_decap_4 FILLER_42_101 ();
 sg13g2_decap_8 FILLER_42_109 ();
 sg13g2_decap_8 FILLER_42_116 ();
 sg13g2_fill_1 FILLER_42_123 ();
 sg13g2_decap_4 FILLER_42_155 ();
 sg13g2_fill_1 FILLER_42_159 ();
 sg13g2_decap_4 FILLER_42_168 ();
 sg13g2_fill_1 FILLER_42_172 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_196 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_fill_2 FILLER_42_217 ();
 sg13g2_fill_1 FILLER_42_219 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_4 FILLER_42_231 ();
 sg13g2_fill_1 FILLER_42_235 ();
 sg13g2_decap_8 FILLER_42_241 ();
 sg13g2_decap_8 FILLER_42_248 ();
 sg13g2_decap_8 FILLER_42_255 ();
 sg13g2_fill_2 FILLER_42_262 ();
 sg13g2_decap_4 FILLER_42_268 ();
 sg13g2_fill_2 FILLER_42_272 ();
 sg13g2_fill_2 FILLER_42_279 ();
 sg13g2_fill_1 FILLER_42_281 ();
 sg13g2_decap_8 FILLER_42_291 ();
 sg13g2_decap_8 FILLER_42_298 ();
 sg13g2_fill_2 FILLER_42_305 ();
 sg13g2_fill_2 FILLER_42_312 ();
 sg13g2_fill_1 FILLER_42_314 ();
 sg13g2_decap_4 FILLER_42_329 ();
 sg13g2_fill_1 FILLER_42_333 ();
 sg13g2_fill_2 FILLER_42_338 ();
 sg13g2_decap_8 FILLER_42_349 ();
 sg13g2_fill_2 FILLER_42_356 ();
 sg13g2_fill_1 FILLER_42_358 ();
 sg13g2_fill_1 FILLER_42_367 ();
 sg13g2_fill_2 FILLER_42_372 ();
 sg13g2_decap_4 FILLER_42_382 ();
 sg13g2_fill_2 FILLER_42_386 ();
 sg13g2_decap_4 FILLER_42_426 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_4 FILLER_43_21 ();
 sg13g2_fill_1 FILLER_43_25 ();
 sg13g2_fill_2 FILLER_43_72 ();
 sg13g2_decap_8 FILLER_43_78 ();
 sg13g2_decap_4 FILLER_43_119 ();
 sg13g2_fill_1 FILLER_43_123 ();
 sg13g2_fill_1 FILLER_43_145 ();
 sg13g2_decap_8 FILLER_43_151 ();
 sg13g2_decap_4 FILLER_43_158 ();
 sg13g2_fill_1 FILLER_43_162 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_fill_2 FILLER_43_175 ();
 sg13g2_fill_2 FILLER_43_180 ();
 sg13g2_fill_1 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_195 ();
 sg13g2_fill_2 FILLER_43_202 ();
 sg13g2_fill_1 FILLER_43_208 ();
 sg13g2_decap_8 FILLER_43_213 ();
 sg13g2_decap_4 FILLER_43_220 ();
 sg13g2_decap_8 FILLER_43_228 ();
 sg13g2_decap_8 FILLER_43_235 ();
 sg13g2_decap_8 FILLER_43_242 ();
 sg13g2_decap_8 FILLER_43_249 ();
 sg13g2_decap_8 FILLER_43_256 ();
 sg13g2_fill_1 FILLER_43_263 ();
 sg13g2_decap_4 FILLER_43_284 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_fill_1 FILLER_43_329 ();
 sg13g2_decap_4 FILLER_43_336 ();
 sg13g2_fill_1 FILLER_43_340 ();
 sg13g2_fill_2 FILLER_43_346 ();
 sg13g2_fill_1 FILLER_43_348 ();
 sg13g2_fill_1 FILLER_43_354 ();
 sg13g2_decap_8 FILLER_43_359 ();
 sg13g2_decap_4 FILLER_43_366 ();
 sg13g2_fill_1 FILLER_43_370 ();
 sg13g2_fill_1 FILLER_43_383 ();
 sg13g2_decap_8 FILLER_43_398 ();
 sg13g2_decap_4 FILLER_43_405 ();
 sg13g2_fill_1 FILLER_43_409 ();
 sg13g2_decap_8 FILLER_43_418 ();
 sg13g2_decap_4 FILLER_43_425 ();
 sg13g2_fill_1 FILLER_43_429 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_fill_1 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_115 ();
 sg13g2_decap_8 FILLER_44_122 ();
 sg13g2_decap_8 FILLER_44_129 ();
 sg13g2_decap_8 FILLER_44_136 ();
 sg13g2_decap_4 FILLER_44_143 ();
 sg13g2_fill_2 FILLER_44_164 ();
 sg13g2_fill_1 FILLER_44_171 ();
 sg13g2_decap_8 FILLER_44_180 ();
 sg13g2_decap_8 FILLER_44_187 ();
 sg13g2_decap_4 FILLER_44_194 ();
 sg13g2_fill_1 FILLER_44_198 ();
 sg13g2_decap_4 FILLER_44_207 ();
 sg13g2_fill_2 FILLER_44_225 ();
 sg13g2_fill_1 FILLER_44_227 ();
 sg13g2_decap_8 FILLER_44_234 ();
 sg13g2_decap_4 FILLER_44_241 ();
 sg13g2_fill_2 FILLER_44_245 ();
 sg13g2_fill_1 FILLER_44_263 ();
 sg13g2_fill_1 FILLER_44_268 ();
 sg13g2_decap_8 FILLER_44_279 ();
 sg13g2_decap_8 FILLER_44_286 ();
 sg13g2_fill_1 FILLER_44_293 ();
 sg13g2_decap_4 FILLER_44_298 ();
 sg13g2_fill_1 FILLER_44_302 ();
 sg13g2_decap_8 FILLER_44_311 ();
 sg13g2_decap_8 FILLER_44_318 ();
 sg13g2_fill_2 FILLER_44_325 ();
 sg13g2_fill_1 FILLER_44_327 ();
 sg13g2_decap_8 FILLER_44_336 ();
 sg13g2_decap_8 FILLER_44_343 ();
 sg13g2_decap_8 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_4 FILLER_44_364 ();
 sg13g2_fill_1 FILLER_44_368 ();
 sg13g2_decap_8 FILLER_44_400 ();
 sg13g2_decap_4 FILLER_44_407 ();
 sg13g2_decap_8 FILLER_44_415 ();
 sg13g2_decap_8 FILLER_44_422 ();
 sg13g2_fill_1 FILLER_44_429 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_4 FILLER_45_14 ();
 sg13g2_fill_2 FILLER_45_18 ();
 sg13g2_decap_4 FILLER_45_24 ();
 sg13g2_fill_2 FILLER_45_28 ();
 sg13g2_decap_4 FILLER_45_38 ();
 sg13g2_fill_2 FILLER_45_42 ();
 sg13g2_fill_2 FILLER_45_56 ();
 sg13g2_fill_1 FILLER_45_65 ();
 sg13g2_fill_1 FILLER_45_75 ();
 sg13g2_fill_1 FILLER_45_80 ();
 sg13g2_decap_8 FILLER_45_86 ();
 sg13g2_decap_8 FILLER_45_93 ();
 sg13g2_fill_2 FILLER_45_100 ();
 sg13g2_fill_1 FILLER_45_110 ();
 sg13g2_fill_1 FILLER_45_120 ();
 sg13g2_fill_1 FILLER_45_125 ();
 sg13g2_decap_8 FILLER_45_129 ();
 sg13g2_decap_4 FILLER_45_136 ();
 sg13g2_fill_2 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_4 FILLER_45_196 ();
 sg13g2_fill_1 FILLER_45_200 ();
 sg13g2_decap_4 FILLER_45_218 ();
 sg13g2_fill_2 FILLER_45_233 ();
 sg13g2_fill_1 FILLER_45_235 ();
 sg13g2_fill_1 FILLER_45_256 ();
 sg13g2_fill_1 FILLER_45_270 ();
 sg13g2_fill_2 FILLER_45_309 ();
 sg13g2_fill_1 FILLER_45_311 ();
 sg13g2_fill_2 FILLER_45_317 ();
 sg13g2_fill_2 FILLER_45_361 ();
 sg13g2_fill_1 FILLER_45_363 ();
 sg13g2_decap_8 FILLER_45_368 ();
 sg13g2_decap_8 FILLER_45_375 ();
 sg13g2_decap_4 FILLER_45_382 ();
 sg13g2_fill_1 FILLER_45_390 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_fill_2 FILLER_46_42 ();
 sg13g2_fill_1 FILLER_46_44 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_4 FILLER_46_77 ();
 sg13g2_fill_2 FILLER_46_81 ();
 sg13g2_fill_1 FILLER_46_87 ();
 sg13g2_fill_2 FILLER_46_148 ();
 sg13g2_fill_2 FILLER_46_166 ();
 sg13g2_fill_2 FILLER_46_176 ();
 sg13g2_fill_2 FILLER_46_183 ();
 sg13g2_fill_1 FILLER_46_185 ();
 sg13g2_decap_8 FILLER_46_192 ();
 sg13g2_decap_8 FILLER_46_199 ();
 sg13g2_fill_2 FILLER_46_206 ();
 sg13g2_fill_1 FILLER_46_208 ();
 sg13g2_decap_4 FILLER_46_221 ();
 sg13g2_decap_8 FILLER_46_262 ();
 sg13g2_fill_2 FILLER_46_269 ();
 sg13g2_fill_2 FILLER_46_292 ();
 sg13g2_decap_4 FILLER_46_298 ();
 sg13g2_fill_2 FILLER_46_302 ();
 sg13g2_fill_1 FILLER_46_330 ();
 sg13g2_fill_1 FILLER_46_335 ();
 sg13g2_decap_8 FILLER_46_366 ();
 sg13g2_decap_4 FILLER_46_373 ();
 sg13g2_fill_1 FILLER_46_386 ();
 sg13g2_fill_1 FILLER_46_391 ();
 sg13g2_fill_1 FILLER_46_397 ();
 sg13g2_fill_1 FILLER_46_403 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_fill_2 FILLER_47_42 ();
 sg13g2_decap_4 FILLER_47_52 ();
 sg13g2_fill_1 FILLER_47_56 ();
 sg13g2_decap_4 FILLER_47_62 ();
 sg13g2_fill_1 FILLER_47_66 ();
 sg13g2_fill_2 FILLER_47_71 ();
 sg13g2_fill_1 FILLER_47_73 ();
 sg13g2_fill_2 FILLER_47_82 ();
 sg13g2_decap_8 FILLER_47_88 ();
 sg13g2_decap_8 FILLER_47_95 ();
 sg13g2_fill_2 FILLER_47_102 ();
 sg13g2_fill_1 FILLER_47_104 ();
 sg13g2_fill_2 FILLER_47_109 ();
 sg13g2_decap_4 FILLER_47_115 ();
 sg13g2_fill_1 FILLER_47_123 ();
 sg13g2_fill_2 FILLER_47_132 ();
 sg13g2_decap_8 FILLER_47_138 ();
 sg13g2_decap_4 FILLER_47_145 ();
 sg13g2_decap_8 FILLER_47_157 ();
 sg13g2_decap_8 FILLER_47_164 ();
 sg13g2_fill_2 FILLER_47_171 ();
 sg13g2_fill_1 FILLER_47_173 ();
 sg13g2_fill_1 FILLER_47_179 ();
 sg13g2_fill_1 FILLER_47_185 ();
 sg13g2_decap_8 FILLER_47_204 ();
 sg13g2_decap_8 FILLER_47_211 ();
 sg13g2_decap_8 FILLER_47_218 ();
 sg13g2_fill_2 FILLER_47_238 ();
 sg13g2_decap_4 FILLER_47_248 ();
 sg13g2_decap_4 FILLER_47_269 ();
 sg13g2_fill_1 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_279 ();
 sg13g2_decap_8 FILLER_47_286 ();
 sg13g2_decap_4 FILLER_47_293 ();
 sg13g2_fill_2 FILLER_47_297 ();
 sg13g2_fill_2 FILLER_47_303 ();
 sg13g2_decap_4 FILLER_47_309 ();
 sg13g2_fill_2 FILLER_47_313 ();
 sg13g2_decap_8 FILLER_47_320 ();
 sg13g2_decap_8 FILLER_47_327 ();
 sg13g2_decap_8 FILLER_47_334 ();
 sg13g2_decap_4 FILLER_47_341 ();
 sg13g2_fill_1 FILLER_47_345 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_4 FILLER_47_364 ();
 sg13g2_fill_1 FILLER_47_368 ();
 sg13g2_decap_8 FILLER_47_422 ();
 sg13g2_fill_1 FILLER_47_429 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_4 FILLER_48_14 ();
 sg13g2_fill_2 FILLER_48_18 ();
 sg13g2_decap_8 FILLER_48_24 ();
 sg13g2_decap_4 FILLER_48_31 ();
 sg13g2_fill_2 FILLER_48_46 ();
 sg13g2_fill_2 FILLER_48_104 ();
 sg13g2_fill_1 FILLER_48_106 ();
 sg13g2_fill_1 FILLER_48_137 ();
 sg13g2_decap_8 FILLER_48_143 ();
 sg13g2_decap_8 FILLER_48_150 ();
 sg13g2_decap_8 FILLER_48_157 ();
 sg13g2_decap_4 FILLER_48_164 ();
 sg13g2_fill_1 FILLER_48_168 ();
 sg13g2_fill_2 FILLER_48_184 ();
 sg13g2_fill_1 FILLER_48_186 ();
 sg13g2_decap_8 FILLER_48_202 ();
 sg13g2_decap_8 FILLER_48_209 ();
 sg13g2_decap_4 FILLER_48_216 ();
 sg13g2_fill_2 FILLER_48_228 ();
 sg13g2_fill_1 FILLER_48_230 ();
 sg13g2_decap_8 FILLER_48_237 ();
 sg13g2_decap_8 FILLER_48_244 ();
 sg13g2_fill_2 FILLER_48_251 ();
 sg13g2_fill_2 FILLER_48_256 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_fill_2 FILLER_48_273 ();
 sg13g2_fill_1 FILLER_48_275 ();
 sg13g2_fill_2 FILLER_48_287 ();
 sg13g2_decap_4 FILLER_48_293 ();
 sg13g2_fill_2 FILLER_48_327 ();
 sg13g2_decap_8 FILLER_48_333 ();
 sg13g2_decap_4 FILLER_48_340 ();
 sg13g2_fill_1 FILLER_48_344 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_fill_2 FILLER_48_385 ();
 sg13g2_fill_1 FILLER_48_392 ();
 sg13g2_fill_2 FILLER_48_398 ();
 sg13g2_fill_1 FILLER_48_409 ();
 sg13g2_fill_1 FILLER_48_414 ();
 sg13g2_decap_4 FILLER_48_419 ();
 sg13g2_fill_2 FILLER_48_427 ();
 sg13g2_fill_1 FILLER_48_429 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_fill_2 FILLER_49_40 ();
 sg13g2_fill_1 FILLER_49_42 ();
 sg13g2_fill_2 FILLER_49_48 ();
 sg13g2_fill_1 FILLER_49_50 ();
 sg13g2_fill_2 FILLER_49_69 ();
 sg13g2_fill_1 FILLER_49_74 ();
 sg13g2_decap_8 FILLER_49_79 ();
 sg13g2_decap_8 FILLER_49_86 ();
 sg13g2_decap_8 FILLER_49_93 ();
 sg13g2_decap_8 FILLER_49_100 ();
 sg13g2_decap_8 FILLER_49_107 ();
 sg13g2_decap_8 FILLER_49_114 ();
 sg13g2_decap_8 FILLER_49_121 ();
 sg13g2_decap_8 FILLER_49_128 ();
 sg13g2_decap_8 FILLER_49_135 ();
 sg13g2_decap_8 FILLER_49_142 ();
 sg13g2_decap_8 FILLER_49_149 ();
 sg13g2_fill_1 FILLER_49_176 ();
 sg13g2_decap_4 FILLER_49_209 ();
 sg13g2_fill_2 FILLER_49_225 ();
 sg13g2_fill_1 FILLER_49_227 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_242 ();
 sg13g2_decap_8 FILLER_49_249 ();
 sg13g2_fill_2 FILLER_49_262 ();
 sg13g2_fill_2 FILLER_49_269 ();
 sg13g2_fill_1 FILLER_49_271 ();
 sg13g2_fill_1 FILLER_49_276 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_fill_1 FILLER_49_315 ();
 sg13g2_fill_1 FILLER_49_429 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_4 FILLER_50_35 ();
 sg13g2_fill_1 FILLER_50_39 ();
 sg13g2_fill_1 FILLER_50_48 ();
 sg13g2_decap_8 FILLER_50_65 ();
 sg13g2_decap_4 FILLER_50_72 ();
 sg13g2_fill_2 FILLER_50_76 ();
 sg13g2_decap_8 FILLER_50_87 ();
 sg13g2_fill_2 FILLER_50_94 ();
 sg13g2_decap_4 FILLER_50_100 ();
 sg13g2_decap_8 FILLER_50_108 ();
 sg13g2_fill_1 FILLER_50_115 ();
 sg13g2_decap_4 FILLER_50_120 ();
 sg13g2_fill_1 FILLER_50_124 ();
 sg13g2_decap_8 FILLER_50_193 ();
 sg13g2_decap_8 FILLER_50_200 ();
 sg13g2_decap_4 FILLER_50_207 ();
 sg13g2_fill_1 FILLER_50_215 ();
 sg13g2_decap_8 FILLER_50_241 ();
 sg13g2_decap_8 FILLER_50_248 ();
 sg13g2_fill_2 FILLER_50_255 ();
 sg13g2_fill_1 FILLER_50_257 ();
 sg13g2_fill_1 FILLER_50_286 ();
 sg13g2_fill_2 FILLER_50_292 ();
 sg13g2_fill_1 FILLER_50_294 ();
 sg13g2_decap_8 FILLER_50_299 ();
 sg13g2_decap_4 FILLER_50_306 ();
 sg13g2_decap_8 FILLER_50_314 ();
 sg13g2_fill_2 FILLER_50_321 ();
 sg13g2_decap_4 FILLER_50_331 ();
 sg13g2_fill_2 FILLER_50_335 ();
 sg13g2_fill_1 FILLER_50_342 ();
 sg13g2_decap_8 FILLER_50_347 ();
 sg13g2_decap_8 FILLER_50_362 ();
 sg13g2_fill_1 FILLER_50_369 ();
 sg13g2_decap_4 FILLER_50_396 ();
 sg13g2_decap_8 FILLER_50_422 ();
 sg13g2_fill_1 FILLER_50_429 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_48 ();
 sg13g2_decap_8 FILLER_51_55 ();
 sg13g2_fill_1 FILLER_51_62 ();
 sg13g2_fill_1 FILLER_51_74 ();
 sg13g2_fill_1 FILLER_51_83 ();
 sg13g2_fill_1 FILLER_51_88 ();
 sg13g2_fill_2 FILLER_51_115 ();
 sg13g2_fill_1 FILLER_51_117 ();
 sg13g2_fill_1 FILLER_51_127 ();
 sg13g2_decap_8 FILLER_51_167 ();
 sg13g2_decap_8 FILLER_51_177 ();
 sg13g2_decap_8 FILLER_51_184 ();
 sg13g2_decap_8 FILLER_51_191 ();
 sg13g2_decap_8 FILLER_51_198 ();
 sg13g2_fill_2 FILLER_51_205 ();
 sg13g2_fill_2 FILLER_51_235 ();
 sg13g2_fill_2 FILLER_51_241 ();
 sg13g2_fill_1 FILLER_51_243 ();
 sg13g2_decap_4 FILLER_51_253 ();
 sg13g2_fill_2 FILLER_51_257 ();
 sg13g2_decap_4 FILLER_51_276 ();
 sg13g2_fill_2 FILLER_51_280 ();
 sg13g2_fill_2 FILLER_51_312 ();
 sg13g2_fill_1 FILLER_51_314 ();
 sg13g2_decap_8 FILLER_51_319 ();
 sg13g2_decap_8 FILLER_51_331 ();
 sg13g2_decap_8 FILLER_51_338 ();
 sg13g2_decap_8 FILLER_51_345 ();
 sg13g2_fill_1 FILLER_51_352 ();
 sg13g2_fill_1 FILLER_51_392 ();
 sg13g2_fill_2 FILLER_51_402 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_fill_1 FILLER_52_21 ();
 sg13g2_decap_4 FILLER_52_26 ();
 sg13g2_fill_2 FILLER_52_30 ();
 sg13g2_decap_8 FILLER_52_44 ();
 sg13g2_decap_4 FILLER_52_51 ();
 sg13g2_fill_1 FILLER_52_55 ();
 sg13g2_fill_1 FILLER_52_95 ();
 sg13g2_fill_2 FILLER_52_130 ();
 sg13g2_fill_1 FILLER_52_140 ();
 sg13g2_fill_1 FILLER_52_145 ();
 sg13g2_fill_1 FILLER_52_154 ();
 sg13g2_fill_1 FILLER_52_159 ();
 sg13g2_fill_1 FILLER_52_168 ();
 sg13g2_fill_1 FILLER_52_173 ();
 sg13g2_fill_1 FILLER_52_182 ();
 sg13g2_fill_2 FILLER_52_191 ();
 sg13g2_fill_1 FILLER_52_193 ();
 sg13g2_decap_4 FILLER_52_204 ();
 sg13g2_fill_1 FILLER_52_208 ();
 sg13g2_fill_2 FILLER_52_241 ();
 sg13g2_fill_1 FILLER_52_243 ();
 sg13g2_fill_1 FILLER_52_274 ();
 sg13g2_decap_4 FILLER_52_279 ();
 sg13g2_decap_8 FILLER_52_286 ();
 sg13g2_decap_8 FILLER_52_293 ();
 sg13g2_decap_8 FILLER_52_300 ();
 sg13g2_decap_4 FILLER_52_307 ();
 sg13g2_decap_8 FILLER_52_322 ();
 sg13g2_decap_4 FILLER_52_329 ();
 sg13g2_fill_1 FILLER_52_333 ();
 sg13g2_fill_2 FILLER_52_342 ();
 sg13g2_fill_1 FILLER_52_344 ();
 sg13g2_decap_4 FILLER_52_353 ();
 sg13g2_fill_2 FILLER_52_357 ();
 sg13g2_decap_8 FILLER_52_365 ();
 sg13g2_fill_1 FILLER_52_372 ();
 sg13g2_decap_8 FILLER_52_381 ();
 sg13g2_decap_8 FILLER_52_388 ();
 sg13g2_decap_4 FILLER_52_395 ();
 sg13g2_fill_2 FILLER_52_399 ();
 sg13g2_decap_8 FILLER_52_414 ();
 sg13g2_decap_8 FILLER_52_421 ();
 sg13g2_fill_2 FILLER_52_428 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_fill_1 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_59 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_4 FILLER_53_105 ();
 sg13g2_fill_1 FILLER_53_109 ();
 sg13g2_decap_8 FILLER_53_114 ();
 sg13g2_decap_8 FILLER_53_125 ();
 sg13g2_decap_8 FILLER_53_132 ();
 sg13g2_decap_8 FILLER_53_139 ();
 sg13g2_decap_8 FILLER_53_146 ();
 sg13g2_fill_2 FILLER_53_153 ();
 sg13g2_decap_4 FILLER_53_159 ();
 sg13g2_fill_1 FILLER_53_163 ();
 sg13g2_decap_4 FILLER_53_169 ();
 sg13g2_fill_2 FILLER_53_173 ();
 sg13g2_fill_1 FILLER_53_179 ();
 sg13g2_decap_4 FILLER_53_218 ();
 sg13g2_fill_2 FILLER_53_222 ();
 sg13g2_decap_8 FILLER_53_235 ();
 sg13g2_fill_2 FILLER_53_242 ();
 sg13g2_decap_4 FILLER_53_295 ();
 sg13g2_decap_8 FILLER_53_316 ();
 sg13g2_decap_8 FILLER_53_323 ();
 sg13g2_decap_4 FILLER_53_330 ();
 sg13g2_fill_1 FILLER_53_334 ();
 sg13g2_decap_8 FILLER_53_343 ();
 sg13g2_decap_8 FILLER_53_350 ();
 sg13g2_decap_8 FILLER_53_357 ();
 sg13g2_decap_8 FILLER_53_364 ();
 sg13g2_decap_8 FILLER_53_371 ();
 sg13g2_decap_8 FILLER_53_378 ();
 sg13g2_decap_8 FILLER_53_385 ();
 sg13g2_decap_4 FILLER_53_392 ();
 sg13g2_decap_8 FILLER_53_422 ();
 sg13g2_fill_1 FILLER_53_429 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_fill_2 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_51 ();
 sg13g2_decap_4 FILLER_54_58 ();
 sg13g2_fill_1 FILLER_54_62 ();
 sg13g2_decap_4 FILLER_54_67 ();
 sg13g2_decap_8 FILLER_54_75 ();
 sg13g2_decap_4 FILLER_54_82 ();
 sg13g2_fill_2 FILLER_54_86 ();
 sg13g2_decap_8 FILLER_54_93 ();
 sg13g2_fill_2 FILLER_54_100 ();
 sg13g2_decap_8 FILLER_54_114 ();
 sg13g2_decap_8 FILLER_54_121 ();
 sg13g2_decap_8 FILLER_54_128 ();
 sg13g2_decap_8 FILLER_54_135 ();
 sg13g2_decap_8 FILLER_54_142 ();
 sg13g2_decap_4 FILLER_54_149 ();
 sg13g2_fill_2 FILLER_54_153 ();
 sg13g2_decap_8 FILLER_54_190 ();
 sg13g2_decap_8 FILLER_54_197 ();
 sg13g2_decap_8 FILLER_54_204 ();
 sg13g2_fill_2 FILLER_54_211 ();
 sg13g2_decap_4 FILLER_54_217 ();
 sg13g2_decap_8 FILLER_54_230 ();
 sg13g2_decap_8 FILLER_54_237 ();
 sg13g2_decap_4 FILLER_54_244 ();
 sg13g2_fill_1 FILLER_54_248 ();
 sg13g2_fill_1 FILLER_54_273 ();
 sg13g2_fill_2 FILLER_54_308 ();
 sg13g2_fill_1 FILLER_54_310 ();
 sg13g2_decap_8 FILLER_54_319 ();
 sg13g2_fill_1 FILLER_54_326 ();
 sg13g2_fill_1 FILLER_54_357 ();
 sg13g2_decap_8 FILLER_54_362 ();
 sg13g2_decap_4 FILLER_54_369 ();
 sg13g2_fill_2 FILLER_54_373 ();
 sg13g2_decap_4 FILLER_54_379 ();
 sg13g2_decap_8 FILLER_54_388 ();
 sg13g2_fill_1 FILLER_54_395 ();
 sg13g2_fill_1 FILLER_54_400 ();
 sg13g2_decap_8 FILLER_54_410 ();
 sg13g2_decap_8 FILLER_54_417 ();
 sg13g2_decap_4 FILLER_54_424 ();
 sg13g2_fill_2 FILLER_54_428 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_4 FILLER_55_28 ();
 sg13g2_decap_4 FILLER_55_36 ();
 sg13g2_fill_1 FILLER_55_40 ();
 sg13g2_fill_2 FILLER_55_45 ();
 sg13g2_fill_2 FILLER_55_61 ();
 sg13g2_decap_4 FILLER_55_71 ();
 sg13g2_decap_4 FILLER_55_78 ();
 sg13g2_decap_4 FILLER_55_87 ();
 sg13g2_fill_2 FILLER_55_159 ();
 sg13g2_fill_1 FILLER_55_161 ();
 sg13g2_decap_8 FILLER_55_166 ();
 sg13g2_decap_8 FILLER_55_173 ();
 sg13g2_decap_8 FILLER_55_210 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_decap_4 FILLER_55_229 ();
 sg13g2_fill_2 FILLER_55_233 ();
 sg13g2_fill_1 FILLER_55_268 ();
 sg13g2_decap_8 FILLER_55_274 ();
 sg13g2_fill_2 FILLER_55_281 ();
 sg13g2_fill_1 FILLER_55_283 ();
 sg13g2_decap_8 FILLER_55_288 ();
 sg13g2_decap_4 FILLER_55_295 ();
 sg13g2_fill_1 FILLER_55_299 ();
 sg13g2_decap_8 FILLER_55_304 ();
 sg13g2_decap_8 FILLER_55_311 ();
 sg13g2_decap_8 FILLER_55_318 ();
 sg13g2_fill_2 FILLER_55_325 ();
 sg13g2_fill_1 FILLER_55_327 ();
 sg13g2_decap_8 FILLER_55_337 ();
 sg13g2_decap_8 FILLER_55_348 ();
 sg13g2_fill_1 FILLER_55_355 ();
 sg13g2_fill_2 FILLER_55_374 ();
 sg13g2_decap_4 FILLER_55_400 ();
 sg13g2_decap_8 FILLER_55_413 ();
 sg13g2_decap_8 FILLER_55_420 ();
 sg13g2_fill_2 FILLER_55_427 ();
 sg13g2_fill_1 FILLER_55_429 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_fill_2 FILLER_56_14 ();
 sg13g2_fill_2 FILLER_56_47 ();
 sg13g2_fill_1 FILLER_56_49 ();
 sg13g2_fill_1 FILLER_56_90 ();
 sg13g2_fill_1 FILLER_56_138 ();
 sg13g2_fill_2 FILLER_56_143 ();
 sg13g2_fill_1 FILLER_56_149 ();
 sg13g2_decap_8 FILLER_56_159 ();
 sg13g2_decap_8 FILLER_56_170 ();
 sg13g2_decap_8 FILLER_56_177 ();
 sg13g2_decap_8 FILLER_56_184 ();
 sg13g2_fill_2 FILLER_56_195 ();
 sg13g2_fill_1 FILLER_56_197 ();
 sg13g2_fill_1 FILLER_56_228 ();
 sg13g2_fill_2 FILLER_56_234 ();
 sg13g2_fill_1 FILLER_56_241 ();
 sg13g2_fill_2 FILLER_56_254 ();
 sg13g2_fill_1 FILLER_56_256 ();
 sg13g2_decap_8 FILLER_56_271 ();
 sg13g2_decap_4 FILLER_56_278 ();
 sg13g2_fill_2 FILLER_56_282 ();
 sg13g2_decap_8 FILLER_56_288 ();
 sg13g2_decap_4 FILLER_56_295 ();
 sg13g2_fill_2 FILLER_56_299 ();
 sg13g2_fill_2 FILLER_56_317 ();
 sg13g2_fill_1 FILLER_56_319 ();
 sg13g2_fill_2 FILLER_56_334 ();
 sg13g2_decap_8 FILLER_56_350 ();
 sg13g2_fill_2 FILLER_56_357 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_fill_2 FILLER_57_21 ();
 sg13g2_decap_4 FILLER_57_27 ();
 sg13g2_fill_1 FILLER_57_31 ();
 sg13g2_fill_1 FILLER_57_37 ();
 sg13g2_fill_1 FILLER_57_46 ();
 sg13g2_fill_1 FILLER_57_51 ();
 sg13g2_fill_2 FILLER_57_92 ();
 sg13g2_fill_2 FILLER_57_116 ();
 sg13g2_fill_1 FILLER_57_123 ();
 sg13g2_fill_2 FILLER_57_128 ();
 sg13g2_fill_1 FILLER_57_130 ();
 sg13g2_fill_2 FILLER_57_136 ();
 sg13g2_fill_2 FILLER_57_164 ();
 sg13g2_fill_1 FILLER_57_166 ();
 sg13g2_decap_8 FILLER_57_193 ();
 sg13g2_decap_8 FILLER_57_200 ();
 sg13g2_decap_8 FILLER_57_207 ();
 sg13g2_decap_8 FILLER_57_218 ();
 sg13g2_fill_1 FILLER_57_225 ();
 sg13g2_fill_2 FILLER_57_230 ();
 sg13g2_fill_1 FILLER_57_232 ();
 sg13g2_decap_8 FILLER_57_241 ();
 sg13g2_decap_4 FILLER_57_248 ();
 sg13g2_fill_2 FILLER_57_258 ();
 sg13g2_fill_2 FILLER_57_265 ();
 sg13g2_fill_1 FILLER_57_267 ();
 sg13g2_decap_4 FILLER_57_273 ();
 sg13g2_decap_4 FILLER_57_349 ();
 sg13g2_fill_1 FILLER_57_353 ();
 sg13g2_fill_1 FILLER_57_361 ();
 sg13g2_fill_2 FILLER_57_382 ();
 sg13g2_decap_4 FILLER_57_394 ();
 sg13g2_fill_1 FILLER_57_398 ();
 sg13g2_fill_1 FILLER_57_429 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_fill_2 FILLER_58_42 ();
 sg13g2_fill_1 FILLER_58_57 ();
 sg13g2_fill_1 FILLER_58_62 ();
 sg13g2_fill_2 FILLER_58_72 ();
 sg13g2_fill_1 FILLER_58_74 ();
 sg13g2_fill_2 FILLER_58_78 ();
 sg13g2_fill_1 FILLER_58_80 ();
 sg13g2_fill_2 FILLER_58_85 ();
 sg13g2_fill_1 FILLER_58_87 ();
 sg13g2_fill_2 FILLER_58_108 ();
 sg13g2_decap_8 FILLER_58_114 ();
 sg13g2_decap_4 FILLER_58_121 ();
 sg13g2_fill_2 FILLER_58_125 ();
 sg13g2_decap_8 FILLER_58_132 ();
 sg13g2_decap_8 FILLER_58_139 ();
 sg13g2_fill_2 FILLER_58_146 ();
 sg13g2_decap_8 FILLER_58_152 ();
 sg13g2_fill_2 FILLER_58_159 ();
 sg13g2_fill_1 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_166 ();
 sg13g2_fill_2 FILLER_58_173 ();
 sg13g2_fill_1 FILLER_58_175 ();
 sg13g2_decap_8 FILLER_58_180 ();
 sg13g2_fill_2 FILLER_58_187 ();
 sg13g2_decap_8 FILLER_58_201 ();
 sg13g2_decap_8 FILLER_58_208 ();
 sg13g2_decap_8 FILLER_58_215 ();
 sg13g2_decap_8 FILLER_58_222 ();
 sg13g2_decap_8 FILLER_58_229 ();
 sg13g2_fill_2 FILLER_58_236 ();
 sg13g2_decap_4 FILLER_58_243 ();
 sg13g2_fill_2 FILLER_58_262 ();
 sg13g2_fill_2 FILLER_58_322 ();
 sg13g2_decap_8 FILLER_58_369 ();
 sg13g2_decap_8 FILLER_58_376 ();
 sg13g2_fill_1 FILLER_58_383 ();
 sg13g2_decap_8 FILLER_58_394 ();
 sg13g2_fill_1 FILLER_58_401 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_fill_1 FILLER_58_409 ();
 sg13g2_decap_8 FILLER_58_419 ();
 sg13g2_decap_4 FILLER_58_426 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_fill_1 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_55 ();
 sg13g2_decap_8 FILLER_59_62 ();
 sg13g2_decap_8 FILLER_59_69 ();
 sg13g2_decap_4 FILLER_59_76 ();
 sg13g2_fill_2 FILLER_59_85 ();
 sg13g2_fill_1 FILLER_59_87 ();
 sg13g2_decap_8 FILLER_59_93 ();
 sg13g2_decap_8 FILLER_59_100 ();
 sg13g2_fill_1 FILLER_59_107 ();
 sg13g2_fill_1 FILLER_59_112 ();
 sg13g2_fill_2 FILLER_59_139 ();
 sg13g2_decap_4 FILLER_59_167 ();
 sg13g2_fill_2 FILLER_59_171 ();
 sg13g2_decap_8 FILLER_59_203 ();
 sg13g2_fill_1 FILLER_59_222 ();
 sg13g2_fill_1 FILLER_59_231 ();
 sg13g2_decap_4 FILLER_59_240 ();
 sg13g2_fill_1 FILLER_59_253 ();
 sg13g2_fill_1 FILLER_59_258 ();
 sg13g2_fill_1 FILLER_59_281 ();
 sg13g2_fill_2 FILLER_59_292 ();
 sg13g2_fill_1 FILLER_59_294 ();
 sg13g2_decap_8 FILLER_59_299 ();
 sg13g2_decap_8 FILLER_59_306 ();
 sg13g2_decap_4 FILLER_59_313 ();
 sg13g2_fill_1 FILLER_59_317 ();
 sg13g2_decap_4 FILLER_59_327 ();
 sg13g2_fill_1 FILLER_59_331 ();
 sg13g2_decap_8 FILLER_59_336 ();
 sg13g2_decap_8 FILLER_59_343 ();
 sg13g2_decap_8 FILLER_59_357 ();
 sg13g2_decap_8 FILLER_59_364 ();
 sg13g2_fill_2 FILLER_59_371 ();
 sg13g2_fill_1 FILLER_59_373 ();
 sg13g2_decap_4 FILLER_59_380 ();
 sg13g2_decap_8 FILLER_59_390 ();
 sg13g2_fill_2 FILLER_59_397 ();
 sg13g2_fill_1 FILLER_59_399 ();
 sg13g2_decap_8 FILLER_59_404 ();
 sg13g2_decap_8 FILLER_59_411 ();
 sg13g2_decap_8 FILLER_59_418 ();
 sg13g2_decap_4 FILLER_59_425 ();
 sg13g2_fill_1 FILLER_59_429 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_4 FILLER_60_21 ();
 sg13g2_fill_2 FILLER_60_25 ();
 sg13g2_decap_8 FILLER_60_53 ();
 sg13g2_decap_8 FILLER_60_60 ();
 sg13g2_decap_8 FILLER_60_67 ();
 sg13g2_fill_2 FILLER_60_91 ();
 sg13g2_fill_1 FILLER_60_93 ();
 sg13g2_decap_4 FILLER_60_99 ();
 sg13g2_fill_2 FILLER_60_103 ();
 sg13g2_fill_1 FILLER_60_139 ();
 sg13g2_decap_4 FILLER_60_144 ();
 sg13g2_fill_1 FILLER_60_148 ();
 sg13g2_decap_4 FILLER_60_153 ();
 sg13g2_fill_1 FILLER_60_173 ();
 sg13g2_fill_1 FILLER_60_182 ();
 sg13g2_decap_8 FILLER_60_187 ();
 sg13g2_fill_1 FILLER_60_199 ();
 sg13g2_decap_4 FILLER_60_217 ();
 sg13g2_fill_2 FILLER_60_221 ();
 sg13g2_decap_8 FILLER_60_249 ();
 sg13g2_fill_2 FILLER_60_256 ();
 sg13g2_fill_2 FILLER_60_279 ();
 sg13g2_fill_2 FILLER_60_287 ();
 sg13g2_fill_1 FILLER_60_289 ();
 sg13g2_decap_8 FILLER_60_320 ();
 sg13g2_decap_4 FILLER_60_327 ();
 sg13g2_decap_4 FILLER_60_339 ();
 sg13g2_fill_2 FILLER_60_378 ();
 sg13g2_fill_1 FILLER_60_385 ();
 sg13g2_fill_2 FILLER_60_394 ();
 sg13g2_fill_1 FILLER_60_396 ();
 sg13g2_fill_2 FILLER_60_401 ();
 sg13g2_fill_1 FILLER_60_403 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_4 FILLER_61_35 ();
 sg13g2_fill_1 FILLER_61_39 ();
 sg13g2_decap_8 FILLER_61_54 ();
 sg13g2_fill_2 FILLER_61_61 ();
 sg13g2_fill_1 FILLER_61_63 ();
 sg13g2_fill_1 FILLER_61_95 ();
 sg13g2_decap_8 FILLER_61_100 ();
 sg13g2_fill_1 FILLER_61_107 ();
 sg13g2_decap_4 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_132 ();
 sg13g2_fill_1 FILLER_61_139 ();
 sg13g2_decap_8 FILLER_61_170 ();
 sg13g2_decap_8 FILLER_61_187 ();
 sg13g2_fill_2 FILLER_61_194 ();
 sg13g2_fill_1 FILLER_61_196 ();
 sg13g2_fill_2 FILLER_61_205 ();
 sg13g2_fill_2 FILLER_61_219 ();
 sg13g2_fill_1 FILLER_61_221 ();
 sg13g2_fill_2 FILLER_61_230 ();
 sg13g2_decap_4 FILLER_61_236 ();
 sg13g2_fill_1 FILLER_61_244 ();
 sg13g2_decap_8 FILLER_61_249 ();
 sg13g2_decap_8 FILLER_61_256 ();
 sg13g2_decap_8 FILLER_61_263 ();
 sg13g2_fill_1 FILLER_61_270 ();
 sg13g2_decap_8 FILLER_61_286 ();
 sg13g2_decap_4 FILLER_61_293 ();
 sg13g2_decap_8 FILLER_61_301 ();
 sg13g2_decap_8 FILLER_61_308 ();
 sg13g2_decap_8 FILLER_61_320 ();
 sg13g2_fill_1 FILLER_61_327 ();
 sg13g2_decap_8 FILLER_61_339 ();
 sg13g2_fill_2 FILLER_61_346 ();
 sg13g2_fill_1 FILLER_61_348 ();
 sg13g2_fill_1 FILLER_61_398 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_fill_2 FILLER_62_28 ();
 sg13g2_fill_1 FILLER_62_30 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_fill_2 FILLER_62_42 ();
 sg13g2_fill_1 FILLER_62_44 ();
 sg13g2_decap_8 FILLER_62_53 ();
 sg13g2_decap_8 FILLER_62_60 ();
 sg13g2_decap_4 FILLER_62_72 ();
 sg13g2_decap_4 FILLER_62_94 ();
 sg13g2_decap_8 FILLER_62_103 ();
 sg13g2_decap_8 FILLER_62_118 ();
 sg13g2_decap_8 FILLER_62_125 ();
 sg13g2_decap_8 FILLER_62_132 ();
 sg13g2_decap_8 FILLER_62_139 ();
 sg13g2_decap_8 FILLER_62_150 ();
 sg13g2_fill_2 FILLER_62_157 ();
 sg13g2_decap_8 FILLER_62_167 ();
 sg13g2_decap_4 FILLER_62_174 ();
 sg13g2_fill_2 FILLER_62_178 ();
 sg13g2_decap_8 FILLER_62_188 ();
 sg13g2_fill_1 FILLER_62_195 ();
 sg13g2_decap_4 FILLER_62_209 ();
 sg13g2_decap_8 FILLER_62_260 ();
 sg13g2_fill_1 FILLER_62_267 ();
 sg13g2_fill_1 FILLER_62_286 ();
 sg13g2_fill_2 FILLER_62_321 ();
 sg13g2_fill_1 FILLER_62_327 ();
 sg13g2_decap_4 FILLER_62_331 ();
 sg13g2_fill_1 FILLER_62_335 ();
 sg13g2_fill_1 FILLER_62_348 ();
 sg13g2_decap_4 FILLER_62_353 ();
 sg13g2_fill_1 FILLER_62_357 ();
 sg13g2_fill_1 FILLER_62_388 ();
 sg13g2_decap_4 FILLER_62_397 ();
 sg13g2_fill_1 FILLER_62_401 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_decap_8 FILLER_62_418 ();
 sg13g2_decap_4 FILLER_62_425 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_fill_2 FILLER_63_21 ();
 sg13g2_fill_1 FILLER_63_23 ();
 sg13g2_fill_2 FILLER_63_58 ();
 sg13g2_fill_1 FILLER_63_60 ();
 sg13g2_fill_2 FILLER_63_65 ();
 sg13g2_fill_1 FILLER_63_67 ();
 sg13g2_fill_1 FILLER_63_77 ();
 sg13g2_fill_1 FILLER_63_95 ();
 sg13g2_fill_2 FILLER_63_101 ();
 sg13g2_fill_1 FILLER_63_103 ();
 sg13g2_decap_4 FILLER_63_127 ();
 sg13g2_fill_1 FILLER_63_131 ();
 sg13g2_fill_1 FILLER_63_136 ();
 sg13g2_decap_8 FILLER_63_141 ();
 sg13g2_decap_8 FILLER_63_148 ();
 sg13g2_fill_1 FILLER_63_155 ();
 sg13g2_decap_4 FILLER_63_164 ();
 sg13g2_fill_2 FILLER_63_183 ();
 sg13g2_fill_1 FILLER_63_185 ();
 sg13g2_fill_2 FILLER_63_194 ();
 sg13g2_fill_2 FILLER_63_217 ();
 sg13g2_fill_2 FILLER_63_223 ();
 sg13g2_fill_1 FILLER_63_225 ();
 sg13g2_fill_2 FILLER_63_234 ();
 sg13g2_fill_2 FILLER_63_244 ();
 sg13g2_fill_1 FILLER_63_252 ();
 sg13g2_fill_2 FILLER_63_257 ();
 sg13g2_fill_1 FILLER_63_259 ();
 sg13g2_fill_2 FILLER_63_265 ();
 sg13g2_fill_1 FILLER_63_267 ();
 sg13g2_fill_1 FILLER_63_274 ();
 sg13g2_fill_2 FILLER_63_282 ();
 sg13g2_decap_8 FILLER_63_314 ();
 sg13g2_decap_8 FILLER_63_321 ();
 sg13g2_fill_1 FILLER_63_328 ();
 sg13g2_decap_8 FILLER_63_350 ();
 sg13g2_decap_8 FILLER_63_357 ();
 sg13g2_decap_8 FILLER_63_364 ();
 sg13g2_decap_4 FILLER_63_371 ();
 sg13g2_fill_2 FILLER_63_375 ();
 sg13g2_fill_2 FILLER_63_385 ();
 sg13g2_decap_8 FILLER_63_397 ();
 sg13g2_decap_8 FILLER_63_404 ();
 sg13g2_fill_2 FILLER_63_411 ();
 sg13g2_decap_8 FILLER_63_417 ();
 sg13g2_decap_4 FILLER_63_424 ();
 sg13g2_fill_2 FILLER_63_428 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_4 FILLER_64_28 ();
 sg13g2_fill_2 FILLER_64_32 ();
 sg13g2_fill_2 FILLER_64_46 ();
 sg13g2_fill_1 FILLER_64_48 ();
 sg13g2_decap_8 FILLER_64_61 ();
 sg13g2_fill_1 FILLER_64_68 ();
 sg13g2_fill_2 FILLER_64_95 ();
 sg13g2_fill_2 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_124 ();
 sg13g2_fill_2 FILLER_64_131 ();
 sg13g2_fill_1 FILLER_64_163 ();
 sg13g2_fill_1 FILLER_64_177 ();
 sg13g2_decap_4 FILLER_64_186 ();
 sg13g2_fill_2 FILLER_64_190 ();
 sg13g2_decap_8 FILLER_64_195 ();
 sg13g2_decap_4 FILLER_64_202 ();
 sg13g2_fill_1 FILLER_64_206 ();
 sg13g2_decap_8 FILLER_64_211 ();
 sg13g2_decap_4 FILLER_64_218 ();
 sg13g2_decap_8 FILLER_64_232 ();
 sg13g2_decap_4 FILLER_64_239 ();
 sg13g2_fill_1 FILLER_64_243 ();
 sg13g2_decap_8 FILLER_64_255 ();
 sg13g2_fill_1 FILLER_64_288 ();
 sg13g2_fill_2 FILLER_64_306 ();
 sg13g2_decap_8 FILLER_64_312 ();
 sg13g2_decap_4 FILLER_64_319 ();
 sg13g2_fill_2 FILLER_64_323 ();
 sg13g2_fill_1 FILLER_64_338 ();
 sg13g2_decap_8 FILLER_64_344 ();
 sg13g2_decap_8 FILLER_64_351 ();
 sg13g2_decap_8 FILLER_64_358 ();
 sg13g2_decap_4 FILLER_64_365 ();
 sg13g2_fill_1 FILLER_64_376 ();
 sg13g2_fill_1 FILLER_64_386 ();
 sg13g2_fill_2 FILLER_64_395 ();
 sg13g2_fill_2 FILLER_64_401 ();
 sg13g2_fill_1 FILLER_64_403 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_4 FILLER_65_14 ();
 sg13g2_fill_1 FILLER_65_18 ();
 sg13g2_fill_2 FILLER_65_45 ();
 sg13g2_fill_1 FILLER_65_47 ();
 sg13g2_decap_8 FILLER_65_61 ();
 sg13g2_fill_2 FILLER_65_77 ();
 sg13g2_fill_1 FILLER_65_79 ();
 sg13g2_fill_2 FILLER_65_85 ();
 sg13g2_fill_1 FILLER_65_119 ();
 sg13g2_decap_4 FILLER_65_125 ();
 sg13g2_fill_1 FILLER_65_129 ();
 sg13g2_decap_4 FILLER_65_135 ();
 sg13g2_decap_4 FILLER_65_143 ();
 sg13g2_fill_2 FILLER_65_147 ();
 sg13g2_fill_1 FILLER_65_165 ();
 sg13g2_fill_2 FILLER_65_170 ();
 sg13g2_fill_1 FILLER_65_185 ();
 sg13g2_decap_4 FILLER_65_202 ();
 sg13g2_fill_2 FILLER_65_206 ();
 sg13g2_decap_8 FILLER_65_234 ();
 sg13g2_fill_1 FILLER_65_241 ();
 sg13g2_fill_2 FILLER_65_247 ();
 sg13g2_fill_1 FILLER_65_249 ();
 sg13g2_fill_2 FILLER_65_258 ();
 sg13g2_fill_1 FILLER_65_260 ();
 sg13g2_decap_8 FILLER_65_283 ();
 sg13g2_decap_8 FILLER_65_290 ();
 sg13g2_decap_4 FILLER_65_297 ();
 sg13g2_decap_8 FILLER_65_332 ();
 sg13g2_decap_4 FILLER_65_339 ();
 sg13g2_fill_2 FILLER_65_343 ();
 sg13g2_fill_2 FILLER_65_353 ();
 sg13g2_decap_8 FILLER_65_371 ();
 sg13g2_decap_4 FILLER_65_378 ();
 sg13g2_fill_2 FILLER_65_382 ();
 sg13g2_decap_8 FILLER_65_391 ();
 sg13g2_fill_1 FILLER_65_398 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_4 FILLER_66_21 ();
 sg13g2_fill_2 FILLER_66_25 ();
 sg13g2_decap_8 FILLER_66_31 ();
 sg13g2_decap_8 FILLER_66_38 ();
 sg13g2_fill_1 FILLER_66_58 ();
 sg13g2_decap_4 FILLER_66_68 ();
 sg13g2_fill_1 FILLER_66_72 ();
 sg13g2_fill_2 FILLER_66_102 ();
 sg13g2_fill_1 FILLER_66_104 ();
 sg13g2_fill_1 FILLER_66_113 ();
 sg13g2_fill_2 FILLER_66_119 ();
 sg13g2_fill_1 FILLER_66_121 ();
 sg13g2_decap_4 FILLER_66_148 ();
 sg13g2_decap_4 FILLER_66_156 ();
 sg13g2_decap_4 FILLER_66_164 ();
 sg13g2_fill_1 FILLER_66_168 ();
 sg13g2_fill_2 FILLER_66_173 ();
 sg13g2_fill_1 FILLER_66_175 ();
 sg13g2_decap_8 FILLER_66_181 ();
 sg13g2_fill_2 FILLER_66_188 ();
 sg13g2_decap_8 FILLER_66_203 ();
 sg13g2_fill_2 FILLER_66_210 ();
 sg13g2_fill_1 FILLER_66_221 ();
 sg13g2_fill_1 FILLER_66_225 ();
 sg13g2_decap_8 FILLER_66_230 ();
 sg13g2_decap_4 FILLER_66_237 ();
 sg13g2_fill_1 FILLER_66_241 ();
 sg13g2_decap_4 FILLER_66_254 ();
 sg13g2_fill_2 FILLER_66_258 ();
 sg13g2_fill_1 FILLER_66_267 ();
 sg13g2_fill_1 FILLER_66_273 ();
 sg13g2_decap_8 FILLER_66_286 ();
 sg13g2_decap_4 FILLER_66_293 ();
 sg13g2_decap_8 FILLER_66_311 ();
 sg13g2_decap_8 FILLER_66_318 ();
 sg13g2_fill_2 FILLER_66_325 ();
 sg13g2_fill_1 FILLER_66_327 ();
 sg13g2_decap_4 FILLER_66_335 ();
 sg13g2_fill_2 FILLER_66_339 ();
 sg13g2_fill_1 FILLER_66_357 ();
 sg13g2_fill_2 FILLER_66_362 ();
 sg13g2_decap_4 FILLER_66_374 ();
 sg13g2_fill_2 FILLER_66_378 ();
 sg13g2_fill_1 FILLER_66_393 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_fill_2 FILLER_66_418 ();
 sg13g2_decap_4 FILLER_66_425 ();
 sg13g2_fill_1 FILLER_66_429 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_fill_1 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_47 ();
 sg13g2_fill_2 FILLER_67_54 ();
 sg13g2_fill_1 FILLER_67_60 ();
 sg13g2_decap_4 FILLER_67_65 ();
 sg13g2_fill_2 FILLER_67_69 ();
 sg13g2_decap_4 FILLER_67_84 ();
 sg13g2_fill_1 FILLER_67_88 ();
 sg13g2_fill_1 FILLER_67_101 ();
 sg13g2_fill_1 FILLER_67_106 ();
 sg13g2_fill_1 FILLER_67_112 ();
 sg13g2_fill_2 FILLER_67_118 ();
 sg13g2_fill_2 FILLER_67_131 ();
 sg13g2_decap_8 FILLER_67_141 ();
 sg13g2_decap_4 FILLER_67_148 ();
 sg13g2_fill_1 FILLER_67_183 ();
 sg13g2_decap_8 FILLER_67_188 ();
 sg13g2_decap_8 FILLER_67_195 ();
 sg13g2_decap_8 FILLER_67_202 ();
 sg13g2_fill_2 FILLER_67_209 ();
 sg13g2_fill_2 FILLER_67_221 ();
 sg13g2_fill_1 FILLER_67_223 ();
 sg13g2_decap_8 FILLER_67_236 ();
 sg13g2_decap_4 FILLER_67_243 ();
 sg13g2_fill_1 FILLER_67_247 ();
 sg13g2_decap_8 FILLER_67_252 ();
 sg13g2_fill_2 FILLER_67_259 ();
 sg13g2_fill_1 FILLER_67_261 ();
 sg13g2_fill_2 FILLER_67_312 ();
 sg13g2_fill_2 FILLER_67_327 ();
 sg13g2_fill_2 FILLER_67_336 ();
 sg13g2_decap_8 FILLER_67_346 ();
 sg13g2_decap_8 FILLER_67_353 ();
 sg13g2_fill_2 FILLER_67_360 ();
 sg13g2_fill_1 FILLER_67_362 ();
 sg13g2_fill_2 FILLER_67_374 ();
 sg13g2_fill_2 FILLER_67_381 ();
 sg13g2_fill_1 FILLER_67_383 ();
 sg13g2_fill_1 FILLER_67_393 ();
 sg13g2_decap_8 FILLER_67_402 ();
 sg13g2_fill_2 FILLER_67_409 ();
 sg13g2_decap_8 FILLER_67_415 ();
 sg13g2_decap_8 FILLER_67_422 ();
 sg13g2_fill_1 FILLER_67_429 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_fill_2 FILLER_68_14 ();
 sg13g2_fill_1 FILLER_68_16 ();
 sg13g2_decap_4 FILLER_68_51 ();
 sg13g2_fill_2 FILLER_68_55 ();
 sg13g2_decap_8 FILLER_68_60 ();
 sg13g2_decap_8 FILLER_68_67 ();
 sg13g2_fill_2 FILLER_68_74 ();
 sg13g2_fill_1 FILLER_68_76 ();
 sg13g2_decap_8 FILLER_68_86 ();
 sg13g2_fill_2 FILLER_68_93 ();
 sg13g2_fill_1 FILLER_68_95 ();
 sg13g2_decap_8 FILLER_68_100 ();
 sg13g2_decap_8 FILLER_68_107 ();
 sg13g2_decap_8 FILLER_68_114 ();
 sg13g2_fill_2 FILLER_68_121 ();
 sg13g2_fill_1 FILLER_68_123 ();
 sg13g2_decap_4 FILLER_68_132 ();
 sg13g2_fill_1 FILLER_68_136 ();
 sg13g2_decap_8 FILLER_68_142 ();
 sg13g2_fill_2 FILLER_68_149 ();
 sg13g2_decap_8 FILLER_68_203 ();
 sg13g2_decap_8 FILLER_68_210 ();
 sg13g2_decap_4 FILLER_68_217 ();
 sg13g2_fill_1 FILLER_68_221 ();
 sg13g2_fill_2 FILLER_68_238 ();
 sg13g2_fill_1 FILLER_68_240 ();
 sg13g2_decap_4 FILLER_68_271 ();
 sg13g2_fill_2 FILLER_68_357 ();
 sg13g2_fill_2 FILLER_68_389 ();
 sg13g2_decap_4 FILLER_68_399 ();
 sg13g2_fill_2 FILLER_68_403 ();
 sg13g2_decap_8 FILLER_68_409 ();
 sg13g2_decap_8 FILLER_68_416 ();
 sg13g2_decap_8 FILLER_68_423 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_fill_2 FILLER_69_21 ();
 sg13g2_fill_1 FILLER_69_23 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_fill_2 FILLER_69_75 ();
 sg13g2_fill_1 FILLER_69_77 ();
 sg13g2_fill_1 FILLER_69_93 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_4 FILLER_69_119 ();
 sg13g2_fill_2 FILLER_69_123 ();
 sg13g2_decap_4 FILLER_69_151 ();
 sg13g2_fill_2 FILLER_69_159 ();
 sg13g2_decap_4 FILLER_69_165 ();
 sg13g2_fill_1 FILLER_69_169 ();
 sg13g2_decap_8 FILLER_69_180 ();
 sg13g2_fill_1 FILLER_69_187 ();
 sg13g2_fill_1 FILLER_69_197 ();
 sg13g2_decap_8 FILLER_69_206 ();
 sg13g2_fill_2 FILLER_69_213 ();
 sg13g2_fill_2 FILLER_69_219 ();
 sg13g2_fill_1 FILLER_69_225 ();
 sg13g2_decap_4 FILLER_69_233 ();
 sg13g2_fill_2 FILLER_69_237 ();
 sg13g2_decap_8 FILLER_69_253 ();
 sg13g2_decap_8 FILLER_69_260 ();
 sg13g2_decap_8 FILLER_69_267 ();
 sg13g2_fill_2 FILLER_69_274 ();
 sg13g2_fill_1 FILLER_69_276 ();
 sg13g2_decap_4 FILLER_69_289 ();
 sg13g2_decap_8 FILLER_69_301 ();
 sg13g2_decap_4 FILLER_69_308 ();
 sg13g2_fill_1 FILLER_69_325 ();
 sg13g2_decap_4 FILLER_69_350 ();
 sg13g2_fill_2 FILLER_69_354 ();
 sg13g2_fill_2 FILLER_69_369 ();
 sg13g2_fill_1 FILLER_69_383 ();
 sg13g2_fill_2 FILLER_69_397 ();
 sg13g2_decap_4 FILLER_69_409 ();
 sg13g2_fill_1 FILLER_69_413 ();
 sg13g2_fill_2 FILLER_69_427 ();
 sg13g2_fill_1 FILLER_69_429 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_4 FILLER_70_28 ();
 sg13g2_fill_1 FILLER_70_32 ();
 sg13g2_fill_2 FILLER_70_48 ();
 sg13g2_fill_1 FILLER_70_50 ();
 sg13g2_fill_1 FILLER_70_70 ();
 sg13g2_decap_4 FILLER_70_77 ();
 sg13g2_fill_1 FILLER_70_134 ();
 sg13g2_decap_8 FILLER_70_139 ();
 sg13g2_decap_8 FILLER_70_146 ();
 sg13g2_decap_8 FILLER_70_153 ();
 sg13g2_decap_8 FILLER_70_160 ();
 sg13g2_fill_2 FILLER_70_167 ();
 sg13g2_fill_1 FILLER_70_169 ();
 sg13g2_decap_8 FILLER_70_173 ();
 sg13g2_fill_2 FILLER_70_219 ();
 sg13g2_decap_8 FILLER_70_262 ();
 sg13g2_decap_8 FILLER_70_269 ();
 sg13g2_decap_8 FILLER_70_276 ();
 sg13g2_decap_4 FILLER_70_283 ();
 sg13g2_fill_1 FILLER_70_287 ();
 sg13g2_decap_8 FILLER_70_291 ();
 sg13g2_decap_8 FILLER_70_298 ();
 sg13g2_decap_8 FILLER_70_305 ();
 sg13g2_decap_8 FILLER_70_312 ();
 sg13g2_decap_8 FILLER_70_319 ();
 sg13g2_decap_8 FILLER_70_326 ();
 sg13g2_decap_8 FILLER_70_333 ();
 sg13g2_decap_8 FILLER_70_340 ();
 sg13g2_decap_8 FILLER_70_347 ();
 sg13g2_decap_8 FILLER_70_354 ();
 sg13g2_fill_2 FILLER_70_361 ();
 sg13g2_fill_1 FILLER_70_363 ();
 sg13g2_fill_1 FILLER_70_381 ();
 sg13g2_fill_2 FILLER_70_395 ();
 sg13g2_fill_2 FILLER_70_401 ();
 sg13g2_fill_1 FILLER_70_403 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_4 FILLER_71_21 ();
 sg13g2_decap_4 FILLER_71_61 ();
 sg13g2_fill_1 FILLER_71_65 ();
 sg13g2_fill_1 FILLER_71_88 ();
 sg13g2_fill_2 FILLER_71_132 ();
 sg13g2_fill_1 FILLER_71_134 ();
 sg13g2_decap_8 FILLER_71_139 ();
 sg13g2_fill_2 FILLER_71_172 ();
 sg13g2_fill_2 FILLER_71_187 ();
 sg13g2_fill_1 FILLER_71_189 ();
 sg13g2_fill_2 FILLER_71_233 ();
 sg13g2_fill_1 FILLER_71_235 ();
 sg13g2_fill_2 FILLER_71_249 ();
 sg13g2_decap_8 FILLER_71_256 ();
 sg13g2_fill_2 FILLER_71_263 ();
 sg13g2_fill_1 FILLER_71_272 ();
 sg13g2_fill_1 FILLER_71_279 ();
 sg13g2_fill_1 FILLER_71_289 ();
 sg13g2_decap_8 FILLER_71_316 ();
 sg13g2_fill_2 FILLER_71_331 ();
 sg13g2_decap_4 FILLER_71_345 ();
 sg13g2_decap_8 FILLER_71_362 ();
 sg13g2_decap_8 FILLER_71_369 ();
 sg13g2_fill_1 FILLER_71_376 ();
 sg13g2_decap_8 FILLER_71_382 ();
 sg13g2_decap_8 FILLER_71_420 ();
 sg13g2_fill_2 FILLER_71_427 ();
 sg13g2_fill_1 FILLER_71_429 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_4 FILLER_72_21 ();
 sg13g2_fill_1 FILLER_72_25 ();
 sg13g2_decap_4 FILLER_72_38 ();
 sg13g2_decap_8 FILLER_72_67 ();
 sg13g2_decap_4 FILLER_72_74 ();
 sg13g2_fill_1 FILLER_72_78 ();
 sg13g2_decap_8 FILLER_72_102 ();
 sg13g2_fill_2 FILLER_72_113 ();
 sg13g2_fill_1 FILLER_72_115 ();
 sg13g2_decap_8 FILLER_72_120 ();
 sg13g2_decap_8 FILLER_72_127 ();
 sg13g2_decap_8 FILLER_72_134 ();
 sg13g2_decap_8 FILLER_72_141 ();
 sg13g2_decap_8 FILLER_72_148 ();
 sg13g2_fill_2 FILLER_72_193 ();
 sg13g2_fill_1 FILLER_72_195 ();
 sg13g2_decap_4 FILLER_72_200 ();
 sg13g2_fill_2 FILLER_72_204 ();
 sg13g2_decap_8 FILLER_72_210 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_fill_2 FILLER_72_224 ();
 sg13g2_fill_1 FILLER_72_226 ();
 sg13g2_decap_8 FILLER_72_235 ();
 sg13g2_fill_2 FILLER_72_242 ();
 sg13g2_fill_2 FILLER_72_249 ();
 sg13g2_fill_1 FILLER_72_251 ();
 sg13g2_fill_2 FILLER_72_259 ();
 sg13g2_fill_1 FILLER_72_261 ();
 sg13g2_decap_4 FILLER_72_293 ();
 sg13g2_decap_8 FILLER_72_301 ();
 sg13g2_fill_2 FILLER_72_308 ();
 sg13g2_decap_8 FILLER_72_318 ();
 sg13g2_decap_4 FILLER_72_325 ();
 sg13g2_fill_2 FILLER_72_329 ();
 sg13g2_decap_8 FILLER_72_357 ();
 sg13g2_decap_8 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_371 ();
 sg13g2_decap_8 FILLER_72_378 ();
 sg13g2_decap_8 FILLER_72_385 ();
 sg13g2_decap_8 FILLER_72_392 ();
 sg13g2_fill_2 FILLER_72_399 ();
 sg13g2_decap_8 FILLER_72_405 ();
 sg13g2_decap_8 FILLER_72_416 ();
 sg13g2_decap_8 FILLER_72_423 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_fill_2 FILLER_73_14 ();
 sg13g2_fill_1 FILLER_73_45 ();
 sg13g2_decap_4 FILLER_73_50 ();
 sg13g2_decap_8 FILLER_73_61 ();
 sg13g2_decap_8 FILLER_73_68 ();
 sg13g2_decap_8 FILLER_73_75 ();
 sg13g2_fill_1 FILLER_73_82 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_124 ();
 sg13g2_decap_8 FILLER_73_131 ();
 sg13g2_decap_8 FILLER_73_138 ();
 sg13g2_decap_8 FILLER_73_145 ();
 sg13g2_decap_8 FILLER_73_152 ();
 sg13g2_decap_8 FILLER_73_159 ();
 sg13g2_decap_4 FILLER_73_170 ();
 sg13g2_decap_4 FILLER_73_200 ();
 sg13g2_decap_8 FILLER_73_208 ();
 sg13g2_decap_8 FILLER_73_215 ();
 sg13g2_fill_1 FILLER_73_222 ();
 sg13g2_decap_4 FILLER_73_280 ();
 sg13g2_decap_8 FILLER_73_301 ();
 sg13g2_fill_2 FILLER_73_308 ();
 sg13g2_fill_1 FILLER_73_310 ();
 sg13g2_decap_8 FILLER_73_315 ();
 sg13g2_decap_8 FILLER_73_322 ();
 sg13g2_decap_8 FILLER_73_329 ();
 sg13g2_fill_2 FILLER_73_336 ();
 sg13g2_fill_1 FILLER_73_338 ();
 sg13g2_decap_8 FILLER_73_343 ();
 sg13g2_decap_8 FILLER_73_350 ();
 sg13g2_decap_8 FILLER_73_357 ();
 sg13g2_decap_8 FILLER_73_364 ();
 sg13g2_decap_8 FILLER_73_371 ();
 sg13g2_decap_8 FILLER_73_378 ();
 sg13g2_decap_8 FILLER_73_385 ();
 sg13g2_decap_8 FILLER_73_392 ();
 sg13g2_decap_8 FILLER_73_399 ();
 sg13g2_decap_8 FILLER_73_406 ();
 sg13g2_decap_8 FILLER_73_413 ();
 sg13g2_decap_8 FILLER_73_420 ();
 sg13g2_fill_2 FILLER_73_427 ();
 sg13g2_fill_1 FILLER_73_429 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_fill_2 FILLER_74_21 ();
 sg13g2_fill_1 FILLER_74_23 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_4 FILLER_74_74 ();
 sg13g2_fill_1 FILLER_74_86 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_fill_1 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_124 ();
 sg13g2_fill_2 FILLER_74_131 ();
 sg13g2_decap_8 FILLER_74_137 ();
 sg13g2_decap_8 FILLER_74_144 ();
 sg13g2_decap_8 FILLER_74_151 ();
 sg13g2_decap_8 FILLER_74_158 ();
 sg13g2_decap_8 FILLER_74_165 ();
 sg13g2_decap_8 FILLER_74_172 ();
 sg13g2_fill_1 FILLER_74_179 ();
 sg13g2_decap_8 FILLER_74_184 ();
 sg13g2_decap_4 FILLER_74_191 ();
 sg13g2_fill_2 FILLER_74_195 ();
 sg13g2_fill_2 FILLER_74_228 ();
 sg13g2_fill_2 FILLER_74_237 ();
 sg13g2_fill_2 FILLER_74_243 ();
 sg13g2_fill_1 FILLER_74_245 ();
 sg13g2_fill_2 FILLER_74_261 ();
 sg13g2_fill_1 FILLER_74_263 ();
 sg13g2_fill_2 FILLER_74_268 ();
 sg13g2_fill_1 FILLER_74_279 ();
 sg13g2_fill_1 FILLER_74_284 ();
 sg13g2_decap_4 FILLER_74_311 ();
 sg13g2_fill_1 FILLER_74_315 ();
 sg13g2_decap_8 FILLER_74_355 ();
 sg13g2_decap_8 FILLER_74_362 ();
 sg13g2_decap_8 FILLER_74_369 ();
 sg13g2_decap_8 FILLER_74_376 ();
 sg13g2_decap_8 FILLER_74_383 ();
 sg13g2_decap_8 FILLER_74_390 ();
 sg13g2_decap_8 FILLER_74_397 ();
 sg13g2_decap_8 FILLER_74_404 ();
 sg13g2_decap_8 FILLER_74_411 ();
 sg13g2_decap_8 FILLER_74_418 ();
 sg13g2_decap_4 FILLER_74_425 ();
 sg13g2_fill_1 FILLER_74_429 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_4 FILLER_75_35 ();
 sg13g2_decap_4 FILLER_75_47 ();
 sg13g2_fill_1 FILLER_75_51 ();
 sg13g2_fill_2 FILLER_75_107 ();
 sg13g2_fill_1 FILLER_75_109 ();
 sg13g2_fill_2 FILLER_75_115 ();
 sg13g2_fill_1 FILLER_75_117 ();
 sg13g2_decap_8 FILLER_75_152 ();
 sg13g2_decap_8 FILLER_75_159 ();
 sg13g2_decap_8 FILLER_75_166 ();
 sg13g2_decap_8 FILLER_75_173 ();
 sg13g2_decap_8 FILLER_75_180 ();
 sg13g2_decap_8 FILLER_75_191 ();
 sg13g2_decap_8 FILLER_75_198 ();
 sg13g2_decap_8 FILLER_75_205 ();
 sg13g2_fill_1 FILLER_75_212 ();
 sg13g2_fill_1 FILLER_75_225 ();
 sg13g2_decap_4 FILLER_75_260 ();
 sg13g2_decap_8 FILLER_75_268 ();
 sg13g2_decap_4 FILLER_75_280 ();
 sg13g2_fill_1 FILLER_75_284 ();
 sg13g2_decap_8 FILLER_75_315 ();
 sg13g2_fill_1 FILLER_75_322 ();
 sg13g2_decap_8 FILLER_75_327 ();
 sg13g2_decap_8 FILLER_75_334 ();
 sg13g2_decap_8 FILLER_75_341 ();
 sg13g2_decap_8 FILLER_75_348 ();
 sg13g2_decap_8 FILLER_75_355 ();
 sg13g2_decap_8 FILLER_75_362 ();
 sg13g2_decap_8 FILLER_75_369 ();
 sg13g2_decap_8 FILLER_75_376 ();
 sg13g2_decap_8 FILLER_75_383 ();
 sg13g2_decap_8 FILLER_75_390 ();
 sg13g2_decap_8 FILLER_75_397 ();
 sg13g2_decap_8 FILLER_75_404 ();
 sg13g2_decap_8 FILLER_75_411 ();
 sg13g2_decap_8 FILLER_75_418 ();
 sg13g2_decap_4 FILLER_75_425 ();
 sg13g2_fill_1 FILLER_75_429 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_fill_2 FILLER_76_28 ();
 sg13g2_fill_1 FILLER_76_42 ();
 sg13g2_fill_1 FILLER_76_67 ();
 sg13g2_fill_2 FILLER_76_72 ();
 sg13g2_fill_1 FILLER_76_74 ();
 sg13g2_decap_8 FILLER_76_81 ();
 sg13g2_decap_4 FILLER_76_88 ();
 sg13g2_fill_1 FILLER_76_92 ();
 sg13g2_fill_2 FILLER_76_97 ();
 sg13g2_fill_2 FILLER_76_103 ();
 sg13g2_fill_1 FILLER_76_105 ();
 sg13g2_fill_2 FILLER_76_114 ();
 sg13g2_fill_1 FILLER_76_116 ();
 sg13g2_fill_2 FILLER_76_125 ();
 sg13g2_fill_1 FILLER_76_127 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_4 FILLER_76_189 ();
 sg13g2_fill_2 FILLER_76_193 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_fill_2 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_265 ();
 sg13g2_decap_8 FILLER_76_272 ();
 sg13g2_decap_8 FILLER_76_279 ();
 sg13g2_decap_4 FILLER_76_286 ();
 sg13g2_fill_2 FILLER_76_290 ();
 sg13g2_decap_8 FILLER_76_296 ();
 sg13g2_decap_8 FILLER_76_303 ();
 sg13g2_decap_8 FILLER_76_310 ();
 sg13g2_decap_8 FILLER_76_317 ();
 sg13g2_decap_8 FILLER_76_324 ();
 sg13g2_decap_8 FILLER_76_331 ();
 sg13g2_decap_8 FILLER_76_338 ();
 sg13g2_decap_8 FILLER_76_345 ();
 sg13g2_decap_8 FILLER_76_352 ();
 sg13g2_decap_8 FILLER_76_359 ();
 sg13g2_decap_8 FILLER_76_366 ();
 sg13g2_decap_8 FILLER_76_373 ();
 sg13g2_decap_8 FILLER_76_380 ();
 sg13g2_decap_8 FILLER_76_387 ();
 sg13g2_decap_8 FILLER_76_394 ();
 sg13g2_decap_8 FILLER_76_401 ();
 sg13g2_decap_8 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_76_415 ();
 sg13g2_decap_8 FILLER_76_422 ();
 sg13g2_fill_1 FILLER_76_429 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_4 FILLER_77_14 ();
 sg13g2_fill_2 FILLER_77_18 ();
 sg13g2_fill_1 FILLER_77_53 ();
 sg13g2_fill_2 FILLER_77_72 ();
 sg13g2_fill_1 FILLER_77_78 ();
 sg13g2_decap_4 FILLER_77_86 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_4 FILLER_77_105 ();
 sg13g2_fill_2 FILLER_77_109 ();
 sg13g2_fill_2 FILLER_77_132 ();
 sg13g2_decap_8 FILLER_77_138 ();
 sg13g2_decap_8 FILLER_77_145 ();
 sg13g2_decap_8 FILLER_77_152 ();
 sg13g2_decap_8 FILLER_77_159 ();
 sg13g2_decap_8 FILLER_77_166 ();
 sg13g2_decap_8 FILLER_77_173 ();
 sg13g2_decap_8 FILLER_77_180 ();
 sg13g2_decap_8 FILLER_77_187 ();
 sg13g2_decap_8 FILLER_77_194 ();
 sg13g2_fill_2 FILLER_77_201 ();
 sg13g2_fill_1 FILLER_77_203 ();
 sg13g2_decap_4 FILLER_77_208 ();
 sg13g2_fill_1 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_233 ();
 sg13g2_fill_2 FILLER_77_240 ();
 sg13g2_fill_1 FILLER_77_255 ();
 sg13g2_decap_8 FILLER_77_290 ();
 sg13g2_decap_8 FILLER_77_297 ();
 sg13g2_decap_8 FILLER_77_304 ();
 sg13g2_decap_8 FILLER_77_311 ();
 sg13g2_decap_8 FILLER_77_318 ();
 sg13g2_decap_8 FILLER_77_325 ();
 sg13g2_decap_8 FILLER_77_332 ();
 sg13g2_decap_8 FILLER_77_339 ();
 sg13g2_decap_8 FILLER_77_346 ();
 sg13g2_decap_8 FILLER_77_353 ();
 sg13g2_decap_8 FILLER_77_360 ();
 sg13g2_decap_8 FILLER_77_367 ();
 sg13g2_decap_8 FILLER_77_374 ();
 sg13g2_decap_8 FILLER_77_381 ();
 sg13g2_decap_8 FILLER_77_388 ();
 sg13g2_decap_8 FILLER_77_395 ();
 sg13g2_decap_8 FILLER_77_402 ();
 sg13g2_decap_8 FILLER_77_409 ();
 sg13g2_decap_8 FILLER_77_416 ();
 sg13g2_decap_8 FILLER_77_423 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_4 FILLER_78_21 ();
 sg13g2_fill_2 FILLER_78_25 ();
 sg13g2_fill_2 FILLER_78_39 ();
 sg13g2_fill_1 FILLER_78_41 ();
 sg13g2_fill_2 FILLER_78_46 ();
 sg13g2_decap_4 FILLER_78_56 ();
 sg13g2_fill_1 FILLER_78_60 ();
 sg13g2_fill_2 FILLER_78_70 ();
 sg13g2_decap_4 FILLER_78_80 ();
 sg13g2_fill_2 FILLER_78_84 ();
 sg13g2_decap_4 FILLER_78_90 ();
 sg13g2_decap_8 FILLER_78_102 ();
 sg13g2_decap_8 FILLER_78_113 ();
 sg13g2_decap_8 FILLER_78_120 ();
 sg13g2_decap_8 FILLER_78_127 ();
 sg13g2_fill_2 FILLER_78_134 ();
 sg13g2_fill_1 FILLER_78_136 ();
 sg13g2_decap_8 FILLER_78_141 ();
 sg13g2_decap_8 FILLER_78_148 ();
 sg13g2_decap_8 FILLER_78_155 ();
 sg13g2_decap_8 FILLER_78_162 ();
 sg13g2_decap_8 FILLER_78_169 ();
 sg13g2_decap_8 FILLER_78_176 ();
 sg13g2_decap_8 FILLER_78_183 ();
 sg13g2_decap_4 FILLER_78_190 ();
 sg13g2_fill_1 FILLER_78_194 ();
 sg13g2_fill_2 FILLER_78_229 ();
 sg13g2_decap_8 FILLER_78_290 ();
 sg13g2_decap_8 FILLER_78_297 ();
 sg13g2_decap_8 FILLER_78_304 ();
 sg13g2_decap_8 FILLER_78_311 ();
 sg13g2_decap_8 FILLER_78_318 ();
 sg13g2_decap_8 FILLER_78_325 ();
 sg13g2_decap_8 FILLER_78_332 ();
 sg13g2_decap_8 FILLER_78_339 ();
 sg13g2_decap_8 FILLER_78_346 ();
 sg13g2_decap_8 FILLER_78_353 ();
 sg13g2_decap_8 FILLER_78_360 ();
 sg13g2_decap_8 FILLER_78_367 ();
 sg13g2_decap_8 FILLER_78_374 ();
 sg13g2_decap_8 FILLER_78_381 ();
 sg13g2_decap_8 FILLER_78_388 ();
 sg13g2_decap_8 FILLER_78_395 ();
 sg13g2_decap_8 FILLER_78_402 ();
 sg13g2_decap_8 FILLER_78_409 ();
 sg13g2_decap_8 FILLER_78_416 ();
 sg13g2_decap_8 FILLER_78_423 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_fill_1 FILLER_79_35 ();
 sg13g2_fill_2 FILLER_79_62 ();
 sg13g2_fill_1 FILLER_79_64 ();
 sg13g2_decap_8 FILLER_79_125 ();
 sg13g2_decap_8 FILLER_79_132 ();
 sg13g2_decap_8 FILLER_79_139 ();
 sg13g2_decap_8 FILLER_79_146 ();
 sg13g2_decap_4 FILLER_79_153 ();
 sg13g2_fill_2 FILLER_79_157 ();
 sg13g2_decap_8 FILLER_79_167 ();
 sg13g2_decap_8 FILLER_79_174 ();
 sg13g2_decap_8 FILLER_79_181 ();
 sg13g2_decap_8 FILLER_79_188 ();
 sg13g2_decap_8 FILLER_79_195 ();
 sg13g2_fill_1 FILLER_79_202 ();
 sg13g2_decap_8 FILLER_79_233 ();
 sg13g2_fill_1 FILLER_79_240 ();
 sg13g2_fill_1 FILLER_79_245 ();
 sg13g2_fill_2 FILLER_79_267 ();
 sg13g2_fill_1 FILLER_79_269 ();
 sg13g2_fill_1 FILLER_79_274 ();
 sg13g2_decap_4 FILLER_79_279 ();
 sg13g2_fill_2 FILLER_79_283 ();
 sg13g2_decap_8 FILLER_79_289 ();
 sg13g2_decap_8 FILLER_79_296 ();
 sg13g2_decap_8 FILLER_79_303 ();
 sg13g2_decap_8 FILLER_79_310 ();
 sg13g2_decap_8 FILLER_79_317 ();
 sg13g2_decap_8 FILLER_79_324 ();
 sg13g2_decap_8 FILLER_79_331 ();
 sg13g2_decap_8 FILLER_79_338 ();
 sg13g2_decap_8 FILLER_79_345 ();
 sg13g2_decap_8 FILLER_79_352 ();
 sg13g2_decap_8 FILLER_79_359 ();
 sg13g2_decap_8 FILLER_79_366 ();
 sg13g2_decap_8 FILLER_79_373 ();
 sg13g2_decap_8 FILLER_79_380 ();
 sg13g2_decap_8 FILLER_79_387 ();
 sg13g2_decap_8 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_401 ();
 sg13g2_decap_8 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_79_415 ();
 sg13g2_decap_8 FILLER_79_422 ();
 sg13g2_fill_1 FILLER_79_429 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_46 ();
 sg13g2_decap_8 FILLER_80_53 ();
 sg13g2_decap_8 FILLER_80_60 ();
 sg13g2_fill_2 FILLER_80_67 ();
 sg13g2_fill_1 FILLER_80_69 ();
 sg13g2_decap_8 FILLER_80_78 ();
 sg13g2_fill_1 FILLER_80_85 ();
 sg13g2_decap_4 FILLER_80_90 ();
 sg13g2_fill_1 FILLER_80_94 ();
 sg13g2_fill_1 FILLER_80_99 ();
 sg13g2_fill_1 FILLER_80_104 ();
 sg13g2_fill_1 FILLER_80_109 ();
 sg13g2_fill_1 FILLER_80_118 ();
 sg13g2_decap_4 FILLER_80_135 ();
 sg13g2_fill_1 FILLER_80_139 ();
 sg13g2_decap_8 FILLER_80_160 ();
 sg13g2_fill_1 FILLER_80_175 ();
 sg13g2_decap_8 FILLER_80_200 ();
 sg13g2_decap_8 FILLER_80_207 ();
 sg13g2_decap_8 FILLER_80_218 ();
 sg13g2_fill_2 FILLER_80_225 ();
 sg13g2_fill_1 FILLER_80_227 ();
 sg13g2_fill_1 FILLER_80_236 ();
 sg13g2_fill_1 FILLER_80_241 ();
 sg13g2_fill_2 FILLER_80_250 ();
 sg13g2_decap_4 FILLER_80_256 ();
 sg13g2_decap_8 FILLER_80_268 ();
 sg13g2_decap_8 FILLER_80_275 ();
 sg13g2_decap_8 FILLER_80_282 ();
 sg13g2_decap_8 FILLER_80_289 ();
 sg13g2_decap_8 FILLER_80_296 ();
 sg13g2_decap_8 FILLER_80_307 ();
 sg13g2_decap_8 FILLER_80_314 ();
 sg13g2_decap_8 FILLER_80_321 ();
 sg13g2_decap_8 FILLER_80_328 ();
 sg13g2_decap_8 FILLER_80_335 ();
 sg13g2_decap_8 FILLER_80_342 ();
 sg13g2_decap_8 FILLER_80_349 ();
 sg13g2_decap_8 FILLER_80_356 ();
 sg13g2_decap_8 FILLER_80_363 ();
 sg13g2_decap_8 FILLER_80_370 ();
 sg13g2_decap_8 FILLER_80_377 ();
 sg13g2_decap_8 FILLER_80_384 ();
 sg13g2_decap_8 FILLER_80_391 ();
 sg13g2_decap_8 FILLER_80_398 ();
 sg13g2_decap_8 FILLER_80_405 ();
 sg13g2_decap_8 FILLER_80_412 ();
 sg13g2_decap_8 FILLER_80_419 ();
 sg13g2_decap_4 FILLER_80_426 ();
endmodule
