module tt_um_rebeccargb_universal_decoder (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;

 sg13g2_inv_1 _0688_ (.Y(_0170_),
    .A(net10));
 sg13g2_buf_1 _0689_ (.A(net8),
    .X(_0181_));
 sg13g2_buf_1 _0690_ (.A(uio_in[4]),
    .X(_0192_));
 sg13g2_inv_2 _0691_ (.Y(_0203_),
    .A(net95));
 sg13g2_buf_2 _0692_ (.A(net2),
    .X(_0213_));
 sg13g2_buf_8 _0693_ (.A(net94),
    .X(_0224_));
 sg13g2_buf_8 _0694_ (.A(net86),
    .X(_0235_));
 sg13g2_buf_1 _0695_ (.A(net71),
    .X(_0246_));
 sg13g2_buf_8 _0696_ (.A(net46),
    .X(_0257_));
 sg13g2_buf_8 _0697_ (.A(ui_in[2]),
    .X(_0268_));
 sg13g2_buf_8 _0698_ (.A(_0268_),
    .X(_0279_));
 sg13g2_buf_1 _0699_ (.A(net85),
    .X(_0290_));
 sg13g2_buf_1 _0700_ (.A(net70),
    .X(_0301_));
 sg13g2_buf_8 _0701_ (.A(ui_in[3]),
    .X(_0312_));
 sg13g2_inv_2 _0702_ (.Y(_0322_),
    .A(_0312_));
 sg13g2_buf_1 _0703_ (.A(_0322_),
    .X(_0333_));
 sg13g2_buf_8 _0704_ (.A(ui_in[6]),
    .X(_0344_));
 sg13g2_buf_8 _0705_ (.A(_0344_),
    .X(_0355_));
 sg13g2_buf_8 _0706_ (.A(net84),
    .X(_0366_));
 sg13g2_buf_1 _0707_ (.A(net68),
    .X(_0377_));
 sg13g2_buf_1 _0708_ (.A(net44),
    .X(_0388_));
 sg13g2_nor2_1 _0709_ (.A(net69),
    .B(net26),
    .Y(_0398_));
 sg13g2_buf_8 _0710_ (.A(net1),
    .X(_0409_));
 sg13g2_buf_8 _0711_ (.A(ui_in[0]),
    .X(_0420_));
 sg13g2_nand2_1 _0712_ (.Y(_0431_),
    .A(_0409_),
    .B(_0420_));
 sg13g2_buf_1 _0713_ (.A(_0431_),
    .X(_0442_));
 sg13g2_o21ai_1 _0714_ (.B1(net26),
    .Y(_0453_),
    .A1(net69),
    .A2(net67));
 sg13g2_o21ai_1 _0715_ (.B1(_0453_),
    .Y(_0464_),
    .A1(net45),
    .A2(_0398_));
 sg13g2_and2_1 _0716_ (.A(net93),
    .B(_0420_),
    .X(_0475_));
 sg13g2_buf_1 _0717_ (.A(_0475_),
    .X(_0485_));
 sg13g2_and2_1 _0718_ (.A(_0268_),
    .B(_0312_),
    .X(_0496_));
 sg13g2_buf_2 _0719_ (.A(_0496_),
    .X(_0507_));
 sg13g2_nand2_1 _0720_ (.Y(_0518_),
    .A(net66),
    .B(_0507_));
 sg13g2_inv_1 _0721_ (.Y(_0529_),
    .A(net7));
 sg13g2_buf_1 _0722_ (.A(_0529_),
    .X(_0540_));
 sg13g2_inv_1 _0723_ (.Y(_0550_),
    .A(net9));
 sg13g2_nor2_1 _0724_ (.A(net83),
    .B(net92),
    .Y(_0561_));
 sg13g2_o21ai_1 _0725_ (.B1(_0561_),
    .Y(_0572_),
    .A1(net27),
    .A2(_0518_));
 sg13g2_a21oi_1 _0726_ (.A1(net27),
    .A2(_0464_),
    .Y(_0583_),
    .B1(_0572_));
 sg13g2_buf_1 _0727_ (.A(net93),
    .X(_0593_));
 sg13g2_buf_1 _0728_ (.A(net82),
    .X(_0604_));
 sg13g2_buf_1 _0729_ (.A(net65),
    .X(_0615_));
 sg13g2_buf_8 _0730_ (.A(_0312_),
    .X(_0626_));
 sg13g2_buf_1 _0731_ (.A(net81),
    .X(_0637_));
 sg13g2_buf_8 _0732_ (.A(net64),
    .X(_0647_));
 sg13g2_buf_1 _0733_ (.A(net42),
    .X(_0658_));
 sg13g2_buf_8 _0734_ (.A(_0420_),
    .X(_0662_));
 sg13g2_buf_8 _0735_ (.A(net93),
    .X(_0663_));
 sg13g2_nand2b_2 _0736_ (.Y(_0664_),
    .B(net79),
    .A_N(net80));
 sg13g2_nand2_1 _0737_ (.Y(_0665_),
    .A(net92),
    .B(net6));
 sg13g2_a221oi_1 _0738_ (.B2(_0664_),
    .C1(_0665_),
    .B1(net25),
    .A1(net43),
    .Y(_0666_),
    .A2(net45));
 sg13g2_nor3_1 _0739_ (.A(_0203_),
    .B(_0583_),
    .C(_0666_),
    .Y(_0667_));
 sg13g2_xor2_1 _0740_ (.B(_0667_),
    .A(net96),
    .X(_0668_));
 sg13g2_nor2_1 _0741_ (.A(_0170_),
    .B(_0668_),
    .Y(net13));
 sg13g2_buf_1 _0742_ (.A(_0268_),
    .X(_0669_));
 sg13g2_buf_8 _0743_ (.A(net81),
    .X(_0670_));
 sg13g2_o21ai_1 _0744_ (.B1(net71),
    .Y(_0671_),
    .A1(net78),
    .A2(net63));
 sg13g2_or2_1 _0745_ (.X(_0672_),
    .B(_0671_),
    .A(net92));
 sg13g2_buf_1 _0746_ (.A(ui_in[5]),
    .X(_0673_));
 sg13g2_buf_1 _0747_ (.A(net91),
    .X(_0674_));
 sg13g2_buf_1 _0748_ (.A(net77),
    .X(_0675_));
 sg13g2_buf_1 _0749_ (.A(net62),
    .X(_0676_));
 sg13g2_nand2b_1 _0750_ (.Y(_0677_),
    .B(net91),
    .A_N(net2));
 sg13g2_buf_2 _0751_ (.A(_0677_),
    .X(_0678_));
 sg13g2_buf_1 _0752_ (.A(net3),
    .X(_0679_));
 sg13g2_buf_1 _0753_ (.A(_0679_),
    .X(_0680_));
 sg13g2_a221oi_1 _0754_ (.B2(net76),
    .C1(net83),
    .B1(_0678_),
    .A1(net26),
    .Y(_0681_),
    .A2(net41));
 sg13g2_nor2_1 _0755_ (.A(_0203_),
    .B(_0681_),
    .Y(_0682_));
 sg13g2_xnor2_1 _0756_ (.Y(_0683_),
    .A(net96),
    .B(_0682_));
 sg13g2_nand2_1 _0757_ (.Y(_0684_),
    .A(net92),
    .B(_0683_));
 sg13g2_a21oi_1 _0758_ (.A1(_0672_),
    .A2(_0684_),
    .Y(net14),
    .B1(net97));
 sg13g2_buf_1 _0759_ (.A(net7),
    .X(_0685_));
 sg13g2_buf_1 _0760_ (.A(net89),
    .X(_0686_));
 sg13g2_buf_1 _0761_ (.A(net75),
    .X(_0000_));
 sg13g2_nand3_1 _0762_ (.B(net94),
    .C(net91),
    .A(_0344_),
    .Y(_0001_));
 sg13g2_buf_1 _0763_ (.A(_0001_),
    .X(_0002_));
 sg13g2_nor2b_1 _0764_ (.A(net93),
    .B_N(_0420_),
    .Y(_0003_));
 sg13g2_buf_1 _0765_ (.A(_0003_),
    .X(_0004_));
 sg13g2_buf_8 _0766_ (.A(_0268_),
    .X(_0005_));
 sg13g2_nor2b_1 _0767_ (.A(net74),
    .B_N(_0312_),
    .Y(_0006_));
 sg13g2_a22oi_1 _0768_ (.Y(_0007_),
    .B1(_0006_),
    .B2(net66),
    .A2(net60),
    .A1(_0507_));
 sg13g2_nor2_1 _0769_ (.A(_0002_),
    .B(_0007_),
    .Y(_0008_));
 sg13g2_nand2b_1 _0770_ (.Y(_0009_),
    .B(net79),
    .A_N(net74));
 sg13g2_buf_8 _0771_ (.A(net80),
    .X(_0010_));
 sg13g2_buf_8 _0772_ (.A(net91),
    .X(_0011_));
 sg13g2_nor2b_2 _0773_ (.A(net73),
    .B_N(_0355_),
    .Y(_0012_));
 sg13g2_nor2b_2 _0774_ (.A(net68),
    .B_N(net73),
    .Y(_0013_));
 sg13g2_a21oi_1 _0775_ (.A1(net59),
    .A2(_0012_),
    .Y(_0014_),
    .B1(_0013_));
 sg13g2_nand3_1 _0776_ (.B(net60),
    .C(_0012_),
    .A(net70),
    .Y(_0015_));
 sg13g2_o21ai_1 _0777_ (.B1(_0015_),
    .Y(_0016_),
    .A1(_0009_),
    .A2(_0014_));
 sg13g2_inv_2 _0778_ (.Y(_0017_),
    .A(net71));
 sg13g2_nor2_1 _0779_ (.A(_0322_),
    .B(net40),
    .Y(_0018_));
 sg13g2_nor2b_2 _0780_ (.A(net82),
    .B_N(net85),
    .Y(_0019_));
 sg13g2_buf_1 _0781_ (.A(_0420_),
    .X(_0020_));
 sg13g2_nor2_2 _0782_ (.A(net72),
    .B(net86),
    .Y(_0021_));
 sg13g2_nand3_1 _0783_ (.B(_0019_),
    .C(_0021_),
    .A(_0529_),
    .Y(_0022_));
 sg13g2_nand2b_2 _0784_ (.Y(_0023_),
    .B(net80),
    .A_N(net79));
 sg13g2_nor2b_2 _0785_ (.A(_0268_),
    .B_N(net94),
    .Y(_0024_));
 sg13g2_and2_1 _0786_ (.A(net72),
    .B(net86),
    .X(_0025_));
 sg13g2_a22oi_1 _0787_ (.Y(_0026_),
    .B1(_0019_),
    .B2(_0025_),
    .A2(_0024_),
    .A1(_0023_));
 sg13g2_nand2_1 _0788_ (.Y(_0027_),
    .A(_0322_),
    .B(_0013_));
 sg13g2_a21oi_1 _0789_ (.A1(_0022_),
    .A2(_0026_),
    .Y(_0028_),
    .B1(_0027_));
 sg13g2_a221oi_1 _0790_ (.B2(_0018_),
    .C1(_0028_),
    .B1(_0016_),
    .A1(net61),
    .Y(_0029_),
    .A2(_0008_));
 sg13g2_nand3b_1 _0791_ (.B(net94),
    .C(net91),
    .Y(_0030_),
    .A_N(_0344_));
 sg13g2_buf_2 _0792_ (.A(_0030_),
    .X(_0031_));
 sg13g2_buf_1 _0793_ (.A(_0031_),
    .X(_0032_));
 sg13g2_inv_1 _0794_ (.Y(_0033_),
    .A(_0662_));
 sg13g2_inv_1 _0795_ (.Y(_0034_),
    .A(net4));
 sg13g2_nand3b_1 _0796_ (.B(net85),
    .C(net79),
    .Y(_0035_),
    .A_N(net81));
 sg13g2_a21oi_1 _0797_ (.A1(_0033_),
    .A2(_0034_),
    .Y(_0036_),
    .B1(_0035_));
 sg13g2_nand2b_1 _0798_ (.Y(_0037_),
    .B(_0670_),
    .A_N(net79));
 sg13g2_a21oi_1 _0799_ (.A1(net70),
    .A2(net83),
    .Y(_0038_),
    .B1(_0037_));
 sg13g2_nor2_1 _0800_ (.A(_0036_),
    .B(_0038_),
    .Y(_0039_));
 sg13g2_nor2_1 _0801_ (.A(net39),
    .B(_0039_),
    .Y(_0040_));
 sg13g2_nand2_1 _0802_ (.Y(_0041_),
    .A(_0268_),
    .B(net81));
 sg13g2_nor2_1 _0803_ (.A(net58),
    .B(_0023_),
    .Y(_0042_));
 sg13g2_nand2b_1 _0804_ (.Y(_0043_),
    .B(_0312_),
    .A_N(_0268_));
 sg13g2_buf_1 _0805_ (.A(_0043_),
    .X(_0044_));
 sg13g2_nor4_1 _0806_ (.A(net82),
    .B(net75),
    .C(net68),
    .D(_0044_),
    .Y(_0045_));
 sg13g2_a21oi_1 _0807_ (.A1(net44),
    .A2(_0042_),
    .Y(_0046_),
    .B1(_0045_));
 sg13g2_buf_8 _0808_ (.A(_0004_),
    .X(_0047_));
 sg13g2_buf_1 _0809_ (.A(_0006_),
    .X(_0048_));
 sg13g2_nand2_2 _0810_ (.Y(_0049_),
    .A(net90),
    .B(net77));
 sg13g2_nand2_1 _0811_ (.Y(_0050_),
    .A(_0540_),
    .B(_0049_));
 sg13g2_nor2b_1 _0812_ (.A(net94),
    .B_N(_0344_),
    .Y(_0051_));
 sg13g2_buf_8 _0813_ (.A(_0051_),
    .X(_0052_));
 sg13g2_nand4_1 _0814_ (.B(net37),
    .C(_0050_),
    .A(_0047_),
    .Y(_0053_),
    .D(net56));
 sg13g2_o21ai_1 _0815_ (.B1(_0053_),
    .Y(_0054_),
    .A1(_0678_),
    .A2(_0046_));
 sg13g2_nor2_1 _0816_ (.A(net59),
    .B(net75),
    .Y(_0055_));
 sg13g2_nand3_1 _0817_ (.B(net85),
    .C(net81),
    .A(_0663_),
    .Y(_0056_));
 sg13g2_nor3_1 _0818_ (.A(net39),
    .B(_0055_),
    .C(_0056_),
    .Y(_0057_));
 sg13g2_or3_1 _0819_ (.A(net93),
    .B(_0005_),
    .C(net81),
    .X(_0058_));
 sg13g2_inv_2 _0820_ (.Y(_0059_),
    .A(net73));
 sg13g2_nand2_1 _0821_ (.Y(_0060_),
    .A(_0059_),
    .B(net56));
 sg13g2_o21ai_1 _0822_ (.B1(net9),
    .Y(_0061_),
    .A1(_0058_),
    .A2(_0060_));
 sg13g2_nor2_1 _0823_ (.A(net74),
    .B(_0626_),
    .Y(_0062_));
 sg13g2_nor2b_2 _0824_ (.A(net94),
    .B_N(net91),
    .Y(_0063_));
 sg13g2_buf_8 _0825_ (.A(_0063_),
    .X(_0064_));
 sg13g2_nor2b_1 _0826_ (.A(net89),
    .B_N(net84),
    .Y(_0065_));
 sg13g2_nand4_1 _0827_ (.B(_0064_),
    .C(net60),
    .A(net55),
    .Y(_0066_),
    .D(_0065_));
 sg13g2_and3_1 _0828_ (.X(_0067_),
    .A(net84),
    .B(net86),
    .C(net73));
 sg13g2_nor2_2 _0829_ (.A(net93),
    .B(_0420_),
    .Y(_0068_));
 sg13g2_nor2b_1 _0830_ (.A(_0312_),
    .B_N(_0268_),
    .Y(_0069_));
 sg13g2_buf_8 _0831_ (.A(_0069_),
    .X(_0070_));
 sg13g2_nand3_1 _0832_ (.B(_0068_),
    .C(net53),
    .A(_0067_),
    .Y(_0071_));
 sg13g2_nand4_1 _0833_ (.B(net55),
    .C(net60),
    .A(net77),
    .Y(_0072_),
    .D(net56));
 sg13g2_a22oi_1 _0834_ (.Y(_0073_),
    .B1(_0071_),
    .B2(_0072_),
    .A2(_0066_),
    .A1(net76));
 sg13g2_or3_1 _0835_ (.A(_0057_),
    .B(_0061_),
    .C(_0073_),
    .X(_0074_));
 sg13g2_and2_1 _0836_ (.A(_0355_),
    .B(_0213_),
    .X(_0075_));
 sg13g2_buf_2 _0837_ (.A(_0075_),
    .X(_0076_));
 sg13g2_buf_1 _0838_ (.A(_0076_),
    .X(_0077_));
 sg13g2_or2_1 _0839_ (.X(_0078_),
    .B(_0420_),
    .A(net1));
 sg13g2_buf_1 _0840_ (.A(_0078_),
    .X(_0079_));
 sg13g2_xnor2_1 _0841_ (.Y(_0080_),
    .A(net74),
    .B(_0626_));
 sg13g2_buf_1 _0842_ (.A(_0059_),
    .X(_0081_));
 sg13g2_o21ai_1 _0843_ (.B1(_0081_),
    .Y(_0082_),
    .A1(net52),
    .A2(_0080_));
 sg13g2_nor2b_2 _0844_ (.A(net80),
    .B_N(net93),
    .Y(_0083_));
 sg13g2_nand2_1 _0845_ (.Y(_0084_),
    .A(_0507_),
    .B(_0083_));
 sg13g2_nand2_1 _0846_ (.Y(_0085_),
    .A(net41),
    .B(_0084_));
 sg13g2_and3_1 _0847_ (.X(_0086_),
    .A(_0077_),
    .B(_0082_),
    .C(_0085_));
 sg13g2_nor4_1 _0848_ (.A(_0040_),
    .B(_0054_),
    .C(_0074_),
    .D(_0086_),
    .Y(_0087_));
 sg13g2_nor2_1 _0849_ (.A(net68),
    .B(_0678_),
    .Y(_0088_));
 sg13g2_buf_1 _0850_ (.A(_0088_),
    .X(_0089_));
 sg13g2_nor2_1 _0851_ (.A(_0664_),
    .B(net57),
    .Y(_0090_));
 sg13g2_o21ai_1 _0852_ (.B1(_0058_),
    .Y(_0091_),
    .A1(_0675_),
    .A2(_0084_));
 sg13g2_a22oi_1 _0853_ (.Y(_0092_),
    .B1(_0091_),
    .B2(_0077_),
    .A2(_0090_),
    .A1(net23));
 sg13g2_nand2b_1 _0854_ (.Y(_0093_),
    .B(_0344_),
    .A_N(net2));
 sg13g2_buf_1 _0855_ (.A(_0093_),
    .X(_0094_));
 sg13g2_nor2_1 _0856_ (.A(_0011_),
    .B(net51),
    .Y(_0095_));
 sg13g2_nor2b_1 _0857_ (.A(net3),
    .B_N(net84),
    .Y(_0096_));
 sg13g2_nand2_1 _0858_ (.Y(_0097_),
    .A(_0063_),
    .B(_0096_));
 sg13g2_inv_1 _0859_ (.Y(_0098_),
    .A(_0097_));
 sg13g2_o21ai_1 _0860_ (.B1(_0507_),
    .Y(_0099_),
    .A1(_0083_),
    .A2(_0003_));
 sg13g2_o21ai_1 _0861_ (.B1(_0518_),
    .Y(_0100_),
    .A1(_0060_),
    .A2(_0099_));
 sg13g2_o21ai_1 _0862_ (.B1(_0100_),
    .Y(_0101_),
    .A1(_0095_),
    .A2(_0098_));
 sg13g2_nand3b_1 _0863_ (.B(net91),
    .C(_0344_),
    .Y(_0102_),
    .A_N(_0213_));
 sg13g2_buf_1 _0864_ (.A(_0102_),
    .X(_0103_));
 sg13g2_nand2b_2 _0865_ (.Y(_0104_),
    .B(net85),
    .A_N(net93));
 sg13g2_a21oi_1 _0866_ (.A1(_0009_),
    .A2(_0104_),
    .Y(_0105_),
    .B1(net90));
 sg13g2_nand2b_1 _0867_ (.Y(_0106_),
    .B(net72),
    .A_N(net7));
 sg13g2_nor2_1 _0868_ (.A(_0104_),
    .B(_0106_),
    .Y(_0107_));
 sg13g2_a221oi_1 _0869_ (.B2(net59),
    .C1(_0107_),
    .B1(_0105_),
    .A1(_0290_),
    .Y(_0108_),
    .A2(_0083_));
 sg13g2_or3_1 _0870_ (.A(net42),
    .B(net50),
    .C(_0108_),
    .X(_0109_));
 sg13g2_nand2_1 _0871_ (.Y(_0110_),
    .A(_0322_),
    .B(net84));
 sg13g2_a21oi_1 _0872_ (.A1(_0669_),
    .A2(_0063_),
    .Y(_0111_),
    .B1(_0024_));
 sg13g2_or3_1 _0873_ (.A(net67),
    .B(_0110_),
    .C(_0111_),
    .X(_0112_));
 sg13g2_buf_8 _0874_ (.A(_0083_),
    .X(_0113_));
 sg13g2_nand4_1 _0875_ (.B(net55),
    .C(_0076_),
    .A(net35),
    .Y(_0114_),
    .D(_0049_));
 sg13g2_and2_1 _0876_ (.A(_0112_),
    .B(_0114_),
    .X(_0115_));
 sg13g2_and4_1 _0877_ (.A(_0092_),
    .B(_0101_),
    .C(_0109_),
    .D(_0115_),
    .X(_0116_));
 sg13g2_nand2_2 _0878_ (.Y(_0117_),
    .A(net35),
    .B(net37));
 sg13g2_inv_2 _0879_ (.Y(_0118_),
    .A(net90));
 sg13g2_nand3_1 _0880_ (.B(net37),
    .C(_0068_),
    .A(_0118_),
    .Y(_0119_));
 sg13g2_a21oi_1 _0881_ (.A1(_0117_),
    .A2(_0119_),
    .Y(_0120_),
    .B1(net40));
 sg13g2_nor2b_1 _0882_ (.A(net73),
    .B_N(net80),
    .Y(_0121_));
 sg13g2_a22oi_1 _0883_ (.Y(_0122_),
    .B1(net53),
    .B2(_0121_),
    .A2(_0006_),
    .A1(_0485_));
 sg13g2_nor2b_2 _0884_ (.A(net74),
    .B_N(_0420_),
    .Y(_0123_));
 sg13g2_nor2b_1 _0885_ (.A(_0011_),
    .B_N(_0663_),
    .Y(_0124_));
 sg13g2_o21ai_1 _0886_ (.B1(_0124_),
    .Y(_0125_),
    .A1(net53),
    .A2(_0123_));
 sg13g2_a21oi_1 _0887_ (.A1(_0122_),
    .A2(_0125_),
    .Y(_0126_),
    .B1(net46));
 sg13g2_nor2_1 _0888_ (.A(_0120_),
    .B(_0126_),
    .Y(_0127_));
 sg13g2_nor2b_1 _0889_ (.A(net63),
    .B_N(net86),
    .Y(_0128_));
 sg13g2_nor2b_1 _0890_ (.A(net86),
    .B_N(net63),
    .Y(_0129_));
 sg13g2_mux2_1 _0891_ (.A0(_0128_),
    .A1(_0129_),
    .S(_0118_),
    .X(_0130_));
 sg13g2_nand4_1 _0892_ (.B(net41),
    .C(net35),
    .A(net45),
    .Y(_0131_),
    .D(_0130_));
 sg13g2_inv_2 _0893_ (.Y(_0132_),
    .A(net84));
 sg13g2_buf_1 _0894_ (.A(_0132_),
    .X(_0133_));
 sg13g2_a21o_1 _0895_ (.A2(_0131_),
    .A1(_0127_),
    .B1(net34),
    .X(_0134_));
 sg13g2_and4_1 _0896_ (.A(_0029_),
    .B(_0087_),
    .C(_0116_),
    .D(_0134_),
    .X(_0135_));
 sg13g2_buf_1 _0897_ (.A(_0033_),
    .X(_0136_));
 sg13g2_inv_1 _0898_ (.Y(_0137_),
    .A(_0279_));
 sg13g2_buf_1 _0899_ (.A(_0137_),
    .X(_0138_));
 sg13g2_nor4_1 _0900_ (.A(_0136_),
    .B(net32),
    .C(net69),
    .D(net39),
    .Y(_0139_));
 sg13g2_buf_1 _0901_ (.A(net53),
    .X(_0140_));
 sg13g2_or2_1 _0902_ (.X(_0141_),
    .B(net81),
    .A(net74));
 sg13g2_nor2_1 _0903_ (.A(net67),
    .B(_0141_),
    .Y(_0142_));
 sg13g2_a21o_1 _0904_ (.A2(_0140_),
    .A1(net38),
    .B1(_0142_),
    .X(_0143_));
 sg13g2_buf_1 _0905_ (.A(net72),
    .X(_0144_));
 sg13g2_nand3_1 _0906_ (.B(_0132_),
    .C(net54),
    .A(net49),
    .Y(_0145_));
 sg13g2_a21oi_1 _0907_ (.A1(net65),
    .A2(_0145_),
    .Y(_0146_),
    .B1(net57));
 sg13g2_nand2_2 _0908_ (.Y(_0147_),
    .A(net82),
    .B(net63));
 sg13g2_and2_1 _0909_ (.A(net78),
    .B(net86),
    .X(_0148_));
 sg13g2_nand2b_1 _0910_ (.Y(_0149_),
    .B(net72),
    .A_N(net73));
 sg13g2_a22oi_1 _0911_ (.Y(_0150_),
    .B1(_0148_),
    .B2(_0149_),
    .A2(_0123_),
    .A1(net54));
 sg13g2_nor3_1 _0912_ (.A(net34),
    .B(_0147_),
    .C(_0150_),
    .Y(_0151_));
 sg13g2_nor4_1 _0913_ (.A(_0139_),
    .B(_0143_),
    .C(_0146_),
    .D(_0151_),
    .Y(_0152_));
 sg13g2_buf_8 _0914_ (.A(_0507_),
    .X(_0153_));
 sg13g2_nand2_1 _0915_ (.Y(_0154_),
    .A(net30),
    .B(_0068_));
 sg13g2_nand3_1 _0916_ (.B(_0076_),
    .C(_0068_),
    .A(net30),
    .Y(_0155_));
 sg13g2_a22oi_1 _0917_ (.Y(_0156_),
    .B1(_0155_),
    .B2(net39),
    .A2(_0154_),
    .A1(_0117_));
 sg13g2_or4_1 _0918_ (.A(net79),
    .B(_0662_),
    .C(_0279_),
    .D(net81),
    .X(_0157_));
 sg13g2_nor2b_1 _0919_ (.A(net9),
    .B_N(net89),
    .Y(_0158_));
 sg13g2_o21ai_1 _0920_ (.B1(_0158_),
    .Y(_0159_),
    .A1(_0118_),
    .A2(_0157_));
 sg13g2_nand2_1 _0921_ (.Y(_0160_),
    .A(net35),
    .B(net55));
 sg13g2_nand2b_1 _0922_ (.Y(_0161_),
    .B(_0160_),
    .A_N(_0159_));
 sg13g2_nor2_1 _0923_ (.A(_0156_),
    .B(_0161_),
    .Y(_0162_));
 sg13g2_nor2_1 _0924_ (.A(_0013_),
    .B(_0012_),
    .Y(_0163_));
 sg13g2_nor3_1 _0925_ (.A(net27),
    .B(_0154_),
    .C(_0163_),
    .Y(_0164_));
 sg13g2_nand2b_1 _0926_ (.Y(_0165_),
    .B(net85),
    .A_N(net86));
 sg13g2_nand2b_1 _0927_ (.Y(_0166_),
    .B(_0165_),
    .A_N(_0024_));
 sg13g2_nor2_1 _0928_ (.A(_0322_),
    .B(_0132_),
    .Y(_0167_));
 sg13g2_and4_1 _0929_ (.A(net41),
    .B(net35),
    .C(_0166_),
    .D(_0167_),
    .X(_0168_));
 sg13g2_nor3_1 _0930_ (.A(_0036_),
    .B(_0164_),
    .C(_0168_),
    .Y(_0169_));
 sg13g2_nand3_1 _0931_ (.B(net30),
    .C(net38),
    .A(_0257_),
    .Y(_0171_));
 sg13g2_o21ai_1 _0932_ (.B1(_0171_),
    .Y(_0172_),
    .A1(net51),
    .A2(_0099_));
 sg13g2_nand2_1 _0933_ (.Y(_0173_),
    .A(net36),
    .B(_0172_));
 sg13g2_nand4_1 _0934_ (.B(_0162_),
    .C(_0169_),
    .A(_0152_),
    .Y(_0174_),
    .D(_0173_));
 sg13g2_nand3_1 _0935_ (.B(net97),
    .C(_0174_),
    .A(net95),
    .Y(_0175_));
 sg13g2_buf_1 _0936_ (.A(net82),
    .X(_0176_));
 sg13g2_nand2b_1 _0937_ (.Y(_0177_),
    .B(net72),
    .A_N(net85));
 sg13g2_o21ai_1 _0938_ (.B1(net26),
    .Y(_0178_),
    .A1(net48),
    .A2(_0177_));
 sg13g2_nand2_1 _0939_ (.Y(_0179_),
    .A(net27),
    .B(_0178_));
 sg13g2_and2_1 _0940_ (.A(net80),
    .B(net74),
    .X(_0180_));
 sg13g2_buf_2 _0941_ (.A(_0180_),
    .X(_0182_));
 sg13g2_buf_1 _0942_ (.A(net49),
    .X(_0183_));
 sg13g2_buf_1 _0943_ (.A(net70),
    .X(_0184_));
 sg13g2_nor3_1 _0944_ (.A(net29),
    .B(net28),
    .C(net46),
    .Y(_0185_));
 sg13g2_o21ai_1 _0945_ (.B1(net43),
    .Y(_0186_),
    .A1(_0182_),
    .A2(_0185_));
 sg13g2_nand2_1 _0946_ (.Y(_0187_),
    .A(net25),
    .B(_0561_));
 sg13g2_a21oi_1 _0947_ (.A1(_0179_),
    .A2(_0186_),
    .Y(_0188_),
    .B1(_0187_));
 sg13g2_o21ai_1 _0948_ (.B1(net42),
    .Y(_0189_),
    .A1(net48),
    .A2(net28));
 sg13g2_o21ai_1 _0949_ (.B1(_0141_),
    .Y(_0190_),
    .A1(_0136_),
    .A2(net58));
 sg13g2_a22oi_1 _0950_ (.Y(_0191_),
    .B1(_0190_),
    .B2(net43),
    .A2(_0189_),
    .A1(net33));
 sg13g2_nor2_1 _0951_ (.A(_0665_),
    .B(_0191_),
    .Y(_0193_));
 sg13g2_buf_1 _0952_ (.A(net9),
    .X(_0194_));
 sg13g2_nand2_1 _0953_ (.Y(_0195_),
    .A(net61),
    .B(net88));
 sg13g2_nor2b_1 _0954_ (.A(net68),
    .B_N(net71),
    .Y(_0196_));
 sg13g2_nor2_1 _0955_ (.A(net48),
    .B(net42),
    .Y(_0197_));
 sg13g2_or2_1 _0956_ (.X(_0198_),
    .B(_0165_),
    .A(net33));
 sg13g2_o21ai_1 _0957_ (.B1(_0198_),
    .Y(_0199_),
    .A1(net29),
    .A2(_0166_));
 sg13g2_a22oi_1 _0958_ (.Y(_0200_),
    .B1(_0197_),
    .B2(_0199_),
    .A2(_0196_),
    .A1(net45));
 sg13g2_o21ai_1 _0959_ (.B1(net95),
    .Y(_0201_),
    .A1(_0195_),
    .A2(_0200_));
 sg13g2_or4_1 _0960_ (.A(net97),
    .B(_0188_),
    .C(_0193_),
    .D(_0201_),
    .X(_0202_));
 sg13g2_o21ai_1 _0961_ (.B1(_0202_),
    .Y(_0204_),
    .A1(_0135_),
    .A2(_0175_));
 sg13g2_xnor2_1 _0962_ (.Y(net15),
    .A(net96),
    .B(_0204_));
 sg13g2_nor3_1 _0963_ (.A(_0431_),
    .B(_0002_),
    .C(net57),
    .Y(_0205_));
 sg13g2_nor3_1 _0964_ (.A(net58),
    .B(net52),
    .C(_0031_),
    .Y(_0206_));
 sg13g2_o21ai_1 _0965_ (.B1(_0540_),
    .Y(_0207_),
    .A1(_0205_),
    .A2(_0206_));
 sg13g2_nor2_1 _0966_ (.A(net65),
    .B(net70),
    .Y(_0208_));
 sg13g2_nand2b_1 _0967_ (.Y(_0209_),
    .B(_0005_),
    .A_N(_0312_));
 sg13g2_buf_2 _0968_ (.A(_0209_),
    .X(_0210_));
 sg13g2_nor2_1 _0969_ (.A(net67),
    .B(_0210_),
    .Y(_0211_));
 sg13g2_nand2b_1 _0970_ (.Y(_0212_),
    .B(net94),
    .A_N(net84));
 sg13g2_buf_2 _0971_ (.A(_0212_),
    .X(_0214_));
 sg13g2_nor2_2 _0972_ (.A(_0059_),
    .B(_0214_),
    .Y(_0215_));
 sg13g2_o21ai_1 _0973_ (.B1(_0215_),
    .Y(_0216_),
    .A1(_0208_),
    .A2(_0211_));
 sg13g2_nand2_1 _0974_ (.Y(_0217_),
    .A(net71),
    .B(_0059_));
 sg13g2_nor3_1 _0975_ (.A(net42),
    .B(_0104_),
    .C(_0217_),
    .Y(_0218_));
 sg13g2_nor2_1 _0976_ (.A(_0678_),
    .B(_0117_),
    .Y(_0219_));
 sg13g2_o21ai_1 _0977_ (.B1(net26),
    .Y(_0220_),
    .A1(_0218_),
    .A2(_0219_));
 sg13g2_nand3_1 _0978_ (.B(_0216_),
    .C(_0220_),
    .A(_0207_),
    .Y(_0221_));
 sg13g2_nor2b_2 _0979_ (.A(net63),
    .B_N(net59),
    .Y(_0222_));
 sg13g2_nor2b_1 _0980_ (.A(net59),
    .B_N(_0637_),
    .Y(_0223_));
 sg13g2_o21ai_1 _0981_ (.B1(net28),
    .Y(_0225_),
    .A1(_0222_),
    .A2(_0223_));
 sg13g2_nand3_1 _0982_ (.B(net37),
    .C(_0049_),
    .A(net29),
    .Y(_0226_));
 sg13g2_o21ai_1 _0983_ (.B1(_0226_),
    .Y(_0227_),
    .A1(_0049_),
    .A2(_0225_));
 sg13g2_nor2_1 _0984_ (.A(net43),
    .B(net51),
    .Y(_0228_));
 sg13g2_nand2_2 _0985_ (.Y(_0229_),
    .A(_0132_),
    .B(net54));
 sg13g2_nand3_1 _0986_ (.B(net36),
    .C(net24),
    .A(_0184_),
    .Y(_0230_));
 sg13g2_o21ai_1 _0987_ (.B1(_0230_),
    .Y(_0231_),
    .A1(net45),
    .A2(_0229_));
 sg13g2_nor2_1 _0988_ (.A(_0333_),
    .B(_0023_),
    .Y(_0232_));
 sg13g2_a22oi_1 _0989_ (.Y(_0233_),
    .B1(_0231_),
    .B2(_0232_),
    .A2(_0228_),
    .A1(_0227_));
 sg13g2_inv_1 _0990_ (.Y(_0234_),
    .A(_0409_));
 sg13g2_nor3_1 _0991_ (.A(_0234_),
    .B(_0141_),
    .C(_0229_),
    .Y(_0236_));
 sg13g2_nor2_1 _0992_ (.A(_0097_),
    .B(_0099_),
    .Y(_0237_));
 sg13g2_nor2_2 _0993_ (.A(_0044_),
    .B(_0079_),
    .Y(_0238_));
 sg13g2_and2_1 _0994_ (.A(_0095_),
    .B(_0238_),
    .X(_0239_));
 sg13g2_nand2_2 _0995_ (.Y(_0240_),
    .A(_0083_),
    .B(net53));
 sg13g2_nand3_1 _0996_ (.B(net60),
    .C(net53),
    .A(net77),
    .Y(_0241_));
 sg13g2_nand2_2 _0997_ (.Y(_0242_),
    .A(net84),
    .B(_0224_));
 sg13g2_a221oi_1 _0998_ (.B2(_0241_),
    .C1(_0242_),
    .B1(_0240_),
    .A1(net90),
    .Y(_0243_),
    .A2(_0675_));
 sg13g2_nor4_1 _0999_ (.A(_0236_),
    .B(_0237_),
    .C(_0239_),
    .D(_0243_),
    .Y(_0244_));
 sg13g2_o21ai_1 _1000_ (.B1(_0244_),
    .Y(_0245_),
    .A1(net61),
    .A2(_0233_));
 sg13g2_nor3_1 _1001_ (.A(_0074_),
    .B(_0221_),
    .C(_0245_),
    .Y(_0247_));
 sg13g2_nand2_1 _1002_ (.Y(_0248_),
    .A(_0092_),
    .B(_0101_));
 sg13g2_nand3_1 _1003_ (.B(_0678_),
    .C(_0090_),
    .A(net26),
    .Y(_0249_));
 sg13g2_nand2_1 _1004_ (.Y(_0250_),
    .A(_0062_),
    .B(_0004_));
 sg13g2_nand2_1 _1005_ (.Y(_0251_),
    .A(net34),
    .B(net40));
 sg13g2_nand4_1 _1006_ (.B(_0153_),
    .C(_0076_),
    .A(net61),
    .Y(_0252_),
    .D(net38));
 sg13g2_o21ai_1 _1007_ (.B1(_0252_),
    .Y(_0253_),
    .A1(_0250_),
    .A2(_0251_));
 sg13g2_nand2_1 _1008_ (.Y(_0254_),
    .A(net41),
    .B(_0253_));
 sg13g2_nor2_1 _1009_ (.A(net52),
    .B(_0210_),
    .Y(_0255_));
 sg13g2_a22oi_1 _1010_ (.Y(_0256_),
    .B1(_0238_),
    .B2(_0098_),
    .A2(_0255_),
    .A1(_0215_));
 sg13g2_nand3_1 _1011_ (.B(_0255_),
    .C(net23),
    .A(net61),
    .Y(_0258_));
 sg13g2_nand4_1 _1012_ (.B(_0254_),
    .C(_0256_),
    .A(_0249_),
    .Y(_0259_),
    .D(_0258_));
 sg13g2_nor2_1 _1013_ (.A(_0049_),
    .B(net51),
    .Y(_0260_));
 sg13g2_a21oi_1 _1014_ (.A1(_0089_),
    .A2(_0211_),
    .Y(_0261_),
    .B1(_0260_));
 sg13g2_nor2_1 _1015_ (.A(_0664_),
    .B(_0210_),
    .Y(_0262_));
 sg13g2_a21oi_1 _1016_ (.A1(_0000_),
    .A2(_0262_),
    .Y(_0263_),
    .B1(_0211_));
 sg13g2_nor2_1 _1017_ (.A(_0261_),
    .B(_0263_),
    .Y(_0264_));
 sg13g2_a22oi_1 _1018_ (.Y(_0265_),
    .B1(_0129_),
    .B2(net29),
    .A2(net55),
    .A1(net46));
 sg13g2_nand3b_1 _1019_ (.B(_0013_),
    .C(net48),
    .Y(_0266_),
    .A_N(_0265_));
 sg13g2_a22oi_1 _1020_ (.Y(_0267_),
    .B1(_0021_),
    .B2(net31),
    .A2(_0025_),
    .A1(net37));
 sg13g2_nor3_1 _1021_ (.A(net65),
    .B(net34),
    .C(_0267_),
    .Y(_0269_));
 sg13g2_a21oi_1 _1022_ (.A1(_0076_),
    .A2(_0211_),
    .Y(_0270_),
    .B1(net10));
 sg13g2_nor2b_1 _1023_ (.A(_0269_),
    .B_N(_0270_),
    .Y(_0271_));
 sg13g2_nand2_1 _1024_ (.Y(_0272_),
    .A(_0266_),
    .B(_0271_));
 sg13g2_nor4_1 _1025_ (.A(_0248_),
    .B(_0259_),
    .C(_0264_),
    .D(_0272_),
    .Y(_0273_));
 sg13g2_o21ai_1 _1026_ (.B1(_0184_),
    .Y(_0274_),
    .A1(net49),
    .A2(net50));
 sg13g2_nand2_1 _1027_ (.Y(_0275_),
    .A(net64),
    .B(_0067_));
 sg13g2_nand2_1 _1028_ (.Y(_0276_),
    .A(net28),
    .B(_0275_));
 sg13g2_a22oi_1 _1029_ (.Y(_0277_),
    .B1(_0276_),
    .B2(_0183_),
    .A2(_0274_),
    .A1(_0658_));
 sg13g2_nor3_1 _1030_ (.A(net28),
    .B(net39),
    .C(_0147_),
    .Y(_0278_));
 sg13g2_nor2_1 _1031_ (.A(_0159_),
    .B(_0278_),
    .Y(_0280_));
 sg13g2_o21ai_1 _1032_ (.B1(_0280_),
    .Y(_0281_),
    .A1(net43),
    .A2(_0277_));
 sg13g2_nand2b_1 _1033_ (.Y(_0282_),
    .B(net85),
    .A_N(net80));
 sg13g2_nand2_1 _1034_ (.Y(_0283_),
    .A(net64),
    .B(_0214_));
 sg13g2_buf_1 _1035_ (.A(_0234_),
    .X(_0284_));
 sg13g2_a22oi_1 _1036_ (.Y(_0285_),
    .B1(_0283_),
    .B2(net47),
    .A2(_0215_),
    .A1(net42));
 sg13g2_o21ai_1 _1037_ (.B1(_0160_),
    .Y(_0286_),
    .A1(_0282_),
    .A2(_0285_));
 sg13g2_nand2_1 _1038_ (.Y(_0287_),
    .A(net32),
    .B(net23));
 sg13g2_a21oi_1 _1039_ (.A1(net25),
    .A2(_0287_),
    .Y(_0288_),
    .B1(net67));
 sg13g2_nand2_1 _1040_ (.Y(_0289_),
    .A(net30),
    .B(net60));
 sg13g2_o21ai_1 _1041_ (.B1(net97),
    .Y(_0291_),
    .A1(_0289_),
    .A2(net39));
 sg13g2_or4_1 _1042_ (.A(_0168_),
    .B(_0286_),
    .C(_0288_),
    .D(_0291_),
    .X(_0292_));
 sg13g2_nor2b_1 _1043_ (.A(net80),
    .B_N(net74),
    .Y(_0293_));
 sg13g2_buf_2 _1044_ (.A(_0293_),
    .X(_0294_));
 sg13g2_buf_1 _1045_ (.A(net10),
    .X(_0295_));
 sg13g2_nand3_1 _1046_ (.B(net88),
    .C(net87),
    .A(net61),
    .Y(_0296_));
 sg13g2_a221oi_1 _1047_ (.B2(_0294_),
    .C1(_0296_),
    .B1(_0129_),
    .A1(_0123_),
    .Y(_0297_),
    .A2(_0128_));
 sg13g2_nand3_1 _1048_ (.B(net68),
    .C(net71),
    .A(net59),
    .Y(_0298_));
 sg13g2_a21oi_1 _1049_ (.A1(net64),
    .A2(_0298_),
    .Y(_0299_),
    .B1(net70));
 sg13g2_a221oi_1 _1050_ (.B2(_0214_),
    .C1(_0299_),
    .B1(_0222_),
    .A1(_0076_),
    .Y(_0300_),
    .A2(_0294_));
 sg13g2_o21ai_1 _1051_ (.B1(_0246_),
    .Y(_0302_),
    .A1(net32),
    .A2(_0132_));
 sg13g2_nand2_1 _1052_ (.Y(_0303_),
    .A(net64),
    .B(net68));
 sg13g2_nand2_1 _1053_ (.Y(_0304_),
    .A(_0165_),
    .B(_0303_));
 sg13g2_a221oi_1 _1054_ (.B2(net33),
    .C1(net48),
    .B1(_0304_),
    .A1(net42),
    .Y(_0305_),
    .A2(_0302_));
 sg13g2_a21o_1 _1055_ (.A2(_0300_),
    .A1(net43),
    .B1(_0305_),
    .X(_0306_));
 sg13g2_o21ai_1 _1056_ (.B1(net76),
    .Y(_0307_),
    .A1(_0013_),
    .A2(net56));
 sg13g2_nand2_1 _1057_ (.Y(_0308_),
    .A(_0118_),
    .B(net44));
 sg13g2_a21oi_1 _1058_ (.A1(net41),
    .A2(_0308_),
    .Y(_0309_),
    .B1(net40));
 sg13g2_nor4_1 _1059_ (.A(net83),
    .B(net88),
    .C(net97),
    .D(_0309_),
    .Y(_0310_));
 sg13g2_a221oi_1 _1060_ (.B2(_0310_),
    .C1(_0203_),
    .B1(_0307_),
    .A1(_0297_),
    .Y(_0311_),
    .A2(_0306_));
 sg13g2_o21ai_1 _1061_ (.B1(_0311_),
    .Y(_0313_),
    .A1(_0281_),
    .A2(_0292_));
 sg13g2_a21oi_1 _1062_ (.A1(_0247_),
    .A2(_0273_),
    .Y(_0314_),
    .B1(_0313_));
 sg13g2_xnor2_1 _1063_ (.Y(net16),
    .A(net96),
    .B(_0314_));
 sg13g2_nand3_1 _1064_ (.B(net31),
    .C(net56),
    .A(_0059_),
    .Y(_0315_));
 sg13g2_o21ai_1 _1065_ (.B1(_0315_),
    .Y(_0316_),
    .A1(net28),
    .A2(net39));
 sg13g2_a22oi_1 _1066_ (.Y(_0317_),
    .B1(_0316_),
    .B2(_0615_),
    .A2(_0095_),
    .A1(_0208_));
 sg13g2_mux2_1 _1067_ (.A0(_0031_),
    .A1(net51),
    .S(_0137_),
    .X(_0318_));
 sg13g2_nand2_1 _1068_ (.Y(_0319_),
    .A(_0322_),
    .B(net35));
 sg13g2_o21ai_1 _1069_ (.B1(_0194_),
    .Y(_0320_),
    .A1(_0318_),
    .A2(_0319_));
 sg13g2_nor2b_1 _1070_ (.A(net90),
    .B_N(_0685_),
    .Y(_0321_));
 sg13g2_nor4_1 _1071_ (.A(net67),
    .B(net58),
    .C(net50),
    .D(_0321_),
    .Y(_0323_));
 sg13g2_a21o_1 _1072_ (.A2(_0142_),
    .A1(net23),
    .B1(_0323_),
    .X(_0324_));
 sg13g2_o21ai_1 _1073_ (.B1(net59),
    .Y(_0325_),
    .A1(net89),
    .A2(net77));
 sg13g2_nand2_1 _1074_ (.Y(_0326_),
    .A(_0604_),
    .B(_0325_));
 sg13g2_nor2b_1 _1075_ (.A(net79),
    .B_N(net73),
    .Y(_0327_));
 sg13g2_nand3_1 _1076_ (.B(net49),
    .C(_0327_),
    .A(net76),
    .Y(_0328_));
 sg13g2_nand2_1 _1077_ (.Y(_0329_),
    .A(_0153_),
    .B(net56));
 sg13g2_a21oi_1 _1078_ (.A1(_0326_),
    .A2(_0328_),
    .Y(_0330_),
    .B1(_0329_));
 sg13g2_a21oi_1 _1079_ (.A1(net76),
    .A2(_0113_),
    .Y(_0331_),
    .B1(_0047_));
 sg13g2_nor3_1 _1080_ (.A(_0002_),
    .B(_0210_),
    .C(_0331_),
    .Y(_0332_));
 sg13g2_nor4_1 _1081_ (.A(_0320_),
    .B(_0324_),
    .C(_0330_),
    .D(_0332_),
    .Y(_0334_));
 sg13g2_o21ai_1 _1082_ (.B1(_0334_),
    .Y(_0335_),
    .A1(net33),
    .A2(_0317_));
 sg13g2_mux2_1 _1083_ (.A0(_0025_),
    .A1(_0021_),
    .S(net47),
    .X(_0336_));
 sg13g2_nor2b_1 _1084_ (.A(net62),
    .B_N(net63),
    .Y(_0337_));
 sg13g2_o21ai_1 _1085_ (.B1(_0025_),
    .Y(_0338_),
    .A1(net32),
    .A2(_0337_));
 sg13g2_o21ai_1 _1086_ (.B1(_0338_),
    .Y(_0339_),
    .A1(_0678_),
    .A2(net57));
 sg13g2_a22oi_1 _1087_ (.Y(_0340_),
    .B1(_0339_),
    .B2(net47),
    .A2(_0336_),
    .A1(net31));
 sg13g2_nand2_1 _1088_ (.Y(_0341_),
    .A(net66),
    .B(_0048_));
 sg13g2_o21ai_1 _1089_ (.B1(_0341_),
    .Y(_0342_),
    .A1(_0081_),
    .A2(_0250_));
 sg13g2_nor2_1 _1090_ (.A(_0676_),
    .B(_0242_),
    .Y(_0343_));
 sg13g2_nor2_1 _1091_ (.A(net58),
    .B(net52),
    .Y(_0345_));
 sg13g2_a22oi_1 _1092_ (.Y(_0346_),
    .B1(_0343_),
    .B2(_0345_),
    .A2(_0342_),
    .A1(_0052_));
 sg13g2_o21ai_1 _1093_ (.B1(_0346_),
    .Y(_0347_),
    .A1(net34),
    .A2(_0340_));
 sg13g2_a21oi_1 _1094_ (.A1(net47),
    .A2(net31),
    .Y(_0348_),
    .B1(net37));
 sg13g2_nand2b_1 _1095_ (.Y(_0349_),
    .B(net89),
    .A_N(net63));
 sg13g2_nand3_1 _1096_ (.B(_0294_),
    .C(_0349_),
    .A(_0284_),
    .Y(_0350_));
 sg13g2_o21ai_1 _1097_ (.B1(_0350_),
    .Y(_0351_),
    .A1(net33),
    .A2(_0348_));
 sg13g2_nand2_1 _1098_ (.Y(_0352_),
    .A(_0089_),
    .B(_0351_));
 sg13g2_nor2_1 _1099_ (.A(net49),
    .B(net57),
    .Y(_0353_));
 sg13g2_nor3_1 _1100_ (.A(_0176_),
    .B(_0032_),
    .C(_0210_),
    .Y(_0354_));
 sg13g2_a221oi_1 _1101_ (.B2(_0095_),
    .C1(_0354_),
    .B1(_0353_),
    .A1(_0345_),
    .Y(_0356_),
    .A2(_0260_));
 sg13g2_nand2b_1 _1102_ (.Y(_0357_),
    .B(_0118_),
    .A_N(_0071_));
 sg13g2_nand4_1 _1103_ (.B(_0352_),
    .C(_0356_),
    .A(_0112_),
    .Y(_0358_),
    .D(_0357_));
 sg13g2_nor4_1 _1104_ (.A(_0221_),
    .B(_0335_),
    .C(_0347_),
    .D(_0358_),
    .Y(_0359_));
 sg13g2_nor2_1 _1105_ (.A(_0234_),
    .B(net32),
    .Y(_0360_));
 sg13g2_nor3_1 _1106_ (.A(net62),
    .B(net67),
    .C(net57),
    .Y(_0361_));
 sg13g2_a21oi_1 _1107_ (.A1(net41),
    .A2(_0360_),
    .Y(_0362_),
    .B1(_0361_));
 sg13g2_a221oi_1 _1108_ (.B2(_0090_),
    .C1(net31),
    .B1(net23),
    .A1(_0215_),
    .Y(_0363_),
    .A2(_0182_));
 sg13g2_o21ai_1 _1109_ (.B1(_0363_),
    .Y(_0364_),
    .A1(_0214_),
    .A2(_0362_));
 sg13g2_nor2_1 _1110_ (.A(net45),
    .B(_0275_),
    .Y(_0365_));
 sg13g2_o21ai_1 _1111_ (.B1(net43),
    .Y(_0367_),
    .A1(_0222_),
    .A2(_0365_));
 sg13g2_nand2b_1 _1112_ (.Y(_0368_),
    .B(_0367_),
    .A_N(_0364_));
 sg13g2_o21ai_1 _1113_ (.B1(net97),
    .Y(_0369_),
    .A1(_0281_),
    .A2(_0368_));
 sg13g2_nor4_1 _1114_ (.A(_0203_),
    .B(net96),
    .C(_0359_),
    .D(_0369_),
    .Y(_0370_));
 sg13g2_nor2_1 _1115_ (.A(net72),
    .B(net78),
    .Y(_0371_));
 sg13g2_a21oi_1 _1116_ (.A1(net48),
    .A2(_0371_),
    .Y(_0372_),
    .B1(_0665_));
 sg13g2_o21ai_1 _1117_ (.B1(net25),
    .Y(_0373_),
    .A1(net47),
    .A2(_0182_));
 sg13g2_or2_1 _1118_ (.X(_0374_),
    .B(net78),
    .A(net90));
 sg13g2_a221oi_1 _1119_ (.B2(_0374_),
    .C1(net64),
    .B1(_0021_),
    .A1(net49),
    .Y(_0375_),
    .A2(_0024_));
 sg13g2_a21oi_1 _1120_ (.A1(net44),
    .A2(_0177_),
    .Y(_0376_),
    .B1(_0671_));
 sg13g2_nor3_1 _1121_ (.A(net48),
    .B(_0375_),
    .C(_0376_),
    .Y(_0378_));
 sg13g2_nor2_1 _1122_ (.A(_0195_),
    .B(_0378_),
    .Y(_0379_));
 sg13g2_nand3_1 _1123_ (.B(_0282_),
    .C(_0177_),
    .A(net64),
    .Y(_0380_));
 sg13g2_o21ai_1 _1124_ (.B1(_0380_),
    .Y(_0381_),
    .A1(net44),
    .A2(_0671_));
 sg13g2_nand2_1 _1125_ (.Y(_0382_),
    .A(_0033_),
    .B(net53));
 sg13g2_nand2_1 _1126_ (.Y(_0383_),
    .A(net59),
    .B(net64));
 sg13g2_a21oi_1 _1127_ (.A1(_0382_),
    .A2(_0383_),
    .Y(_0384_),
    .B1(net46));
 sg13g2_or3_1 _1128_ (.A(net47),
    .B(_0381_),
    .C(_0384_),
    .X(_0385_));
 sg13g2_a221oi_1 _1129_ (.B2(_0385_),
    .C1(net97),
    .B1(_0379_),
    .A1(_0372_),
    .Y(_0386_),
    .A2(_0373_));
 sg13g2_nor2b_1 _1130_ (.A(_0386_),
    .B_N(net8),
    .Y(_0387_));
 sg13g2_and2_1 _1131_ (.A(_0359_),
    .B(_0387_),
    .X(_0389_));
 sg13g2_nor2_1 _1132_ (.A(_0203_),
    .B(net8),
    .Y(_0390_));
 sg13g2_nor2b_1 _1133_ (.A(net95),
    .B_N(net8),
    .Y(_0391_));
 sg13g2_a21o_1 _1134_ (.A2(_0386_),
    .A1(_0390_),
    .B1(_0391_),
    .X(_0392_));
 sg13g2_a21o_1 _1135_ (.A2(_0387_),
    .A1(_0369_),
    .B1(_0392_),
    .X(_0393_));
 sg13g2_nor3_1 _1136_ (.A(_0370_),
    .B(_0389_),
    .C(_0393_),
    .Y(net17));
 sg13g2_nor2_1 _1137_ (.A(_0139_),
    .B(_0143_),
    .Y(_0394_));
 sg13g2_nand2_1 _1138_ (.Y(_0395_),
    .A(net49),
    .B(_0048_));
 sg13g2_o21ai_1 _1139_ (.B1(_0382_),
    .Y(_0396_),
    .A1(_0060_),
    .A2(_0395_));
 sg13g2_nor2b_1 _1140_ (.A(net77),
    .B_N(net71),
    .Y(_0397_));
 sg13g2_a21oi_1 _1141_ (.A1(net32),
    .A2(net54),
    .Y(_0399_),
    .B1(_0397_));
 sg13g2_nand2_1 _1142_ (.Y(_0400_),
    .A(net32),
    .B(_0397_));
 sg13g2_o21ai_1 _1143_ (.B1(_0400_),
    .Y(_0401_),
    .A1(net29),
    .A2(_0399_));
 sg13g2_nor2_1 _1144_ (.A(net44),
    .B(_0147_),
    .Y(_0402_));
 sg13g2_mux2_1 _1145_ (.A0(_0214_),
    .A1(net51),
    .S(_0033_),
    .X(_0403_));
 sg13g2_nor4_1 _1146_ (.A(net65),
    .B(_0676_),
    .C(net58),
    .D(_0403_),
    .Y(_0404_));
 sg13g2_a221oi_1 _1147_ (.B2(_0402_),
    .C1(_0404_),
    .B1(_0401_),
    .A1(_0615_),
    .Y(_0405_),
    .A2(_0396_));
 sg13g2_a22oi_1 _1148_ (.Y(_0406_),
    .B1(_0019_),
    .B2(net62),
    .A2(_0024_),
    .A1(net82));
 sg13g2_nor3_1 _1149_ (.A(net78),
    .B(_0235_),
    .C(net77),
    .Y(_0407_));
 sg13g2_o21ai_1 _1150_ (.B1(net35),
    .Y(_0408_),
    .A1(_0148_),
    .A2(_0407_));
 sg13g2_o21ai_1 _1151_ (.B1(_0408_),
    .Y(_0410_),
    .A1(net33),
    .A2(_0406_));
 sg13g2_and2_1 _1152_ (.A(_0167_),
    .B(_0410_),
    .X(_0411_));
 sg13g2_inv_1 _1153_ (.Y(_0412_),
    .A(net6));
 sg13g2_nand2_1 _1154_ (.Y(_0413_),
    .A(_0234_),
    .B(_0006_));
 sg13g2_a21oi_1 _1155_ (.A1(net49),
    .A2(_0412_),
    .Y(_0414_),
    .B1(_0413_));
 sg13g2_nor2_1 _1156_ (.A(net58),
    .B(_0664_),
    .Y(_0415_));
 sg13g2_nand2_1 _1157_ (.Y(_0416_),
    .A(_0415_),
    .B(net23));
 sg13g2_o21ai_1 _1158_ (.B1(_0416_),
    .Y(_0417_),
    .A1(_0341_),
    .A2(_0103_));
 sg13g2_nor4_1 _1159_ (.A(net87),
    .B(_0411_),
    .C(_0414_),
    .D(_0417_),
    .Y(_0418_));
 sg13g2_nand4_1 _1160_ (.B(_0162_),
    .C(_0405_),
    .A(_0394_),
    .Y(_0419_),
    .D(_0418_));
 sg13g2_a21oi_1 _1161_ (.A1(net70),
    .A2(_0242_),
    .Y(_0421_),
    .B1(net33));
 sg13g2_o21ai_1 _1162_ (.B1(net69),
    .Y(_0422_),
    .A1(_0024_),
    .A2(_0421_));
 sg13g2_nor3_1 _1163_ (.A(net69),
    .B(_0196_),
    .C(_0282_),
    .Y(_0423_));
 sg13g2_nor2_1 _1164_ (.A(net47),
    .B(_0423_),
    .Y(_0424_));
 sg13g2_nor3_1 _1165_ (.A(net34),
    .B(net40),
    .C(_0123_),
    .Y(_0425_));
 sg13g2_nor2_1 _1166_ (.A(net46),
    .B(_0294_),
    .Y(_0426_));
 sg13g2_o21ai_1 _1167_ (.B1(net25),
    .Y(_0427_),
    .A1(_0425_),
    .A2(_0426_));
 sg13g2_a21oi_1 _1168_ (.A1(_0021_),
    .A2(net31),
    .Y(_0428_),
    .B1(net48));
 sg13g2_a22oi_1 _1169_ (.Y(_0429_),
    .B1(_0427_),
    .B2(_0428_),
    .A2(_0424_),
    .A1(_0422_));
 sg13g2_o21ai_1 _1170_ (.B1(net76),
    .Y(_0430_),
    .A1(net36),
    .A2(net24));
 sg13g2_nand3_1 _1171_ (.B(_0229_),
    .C(_0430_),
    .A(_0550_),
    .Y(_0432_));
 sg13g2_o21ai_1 _1172_ (.B1(_0432_),
    .Y(_0433_),
    .A1(net92),
    .A2(_0429_));
 sg13g2_nand3_1 _1173_ (.B(_0295_),
    .C(_0433_),
    .A(net61),
    .Y(_0434_));
 sg13g2_nor2_2 _1174_ (.A(net94),
    .B(net91),
    .Y(_0435_));
 sg13g2_and2_1 _1175_ (.A(net2),
    .B(_0673_),
    .X(_0436_));
 sg13g2_buf_2 _1176_ (.A(_0436_),
    .X(_0437_));
 sg13g2_a22oi_1 _1177_ (.Y(_0438_),
    .B1(_0435_),
    .B2(_0144_),
    .A2(_0294_),
    .A1(_0437_));
 sg13g2_a221oi_1 _1178_ (.B2(_0435_),
    .C1(net82),
    .B1(_0371_),
    .A1(_0437_),
    .Y(_0439_),
    .A2(_0182_));
 sg13g2_a21oi_1 _1179_ (.A1(net65),
    .A2(_0438_),
    .Y(_0440_),
    .B1(_0439_));
 sg13g2_a21oi_1 _1180_ (.A1(_0182_),
    .A2(_0435_),
    .Y(_0441_),
    .B1(_0440_));
 sg13g2_nand2b_1 _1181_ (.Y(_0443_),
    .B(_0059_),
    .A_N(_0035_));
 sg13g2_nand3b_1 _1182_ (.B(net68),
    .C(_0224_),
    .Y(_0444_),
    .A_N(_0020_));
 sg13g2_a21oi_1 _1183_ (.A1(_0413_),
    .A2(_0443_),
    .Y(_0445_),
    .B1(_0444_));
 sg13g2_nor2_1 _1184_ (.A(_0320_),
    .B(_0445_),
    .Y(_0446_));
 sg13g2_o21ai_1 _1185_ (.B1(_0446_),
    .Y(_0447_),
    .A1(_0110_),
    .A2(_0441_));
 sg13g2_nand2b_1 _1186_ (.Y(_0448_),
    .B(net73),
    .A_N(net79));
 sg13g2_nor4_1 _1187_ (.A(_0118_),
    .B(net75),
    .C(_0110_),
    .D(_0448_),
    .Y(_0449_));
 sg13g2_a22oi_1 _1188_ (.Y(_0450_),
    .B1(_0449_),
    .B2(_0123_),
    .A2(_0345_),
    .A1(_0013_));
 sg13g2_mux2_1 _1189_ (.A0(_0042_),
    .A1(_0090_),
    .S(net62),
    .X(_0451_));
 sg13g2_a21oi_1 _1190_ (.A1(net56),
    .A2(_0451_),
    .Y(_0452_),
    .B1(net87));
 sg13g2_o21ai_1 _1191_ (.B1(_0452_),
    .Y(_0454_),
    .A1(_0257_),
    .A2(_0450_));
 sg13g2_a22oi_1 _1192_ (.Y(_0455_),
    .B1(_0415_),
    .B2(net23),
    .A2(_0215_),
    .A1(_0042_));
 sg13g2_o21ai_1 _1193_ (.B1(_0117_),
    .Y(_0456_),
    .A1(_0246_),
    .A2(_0154_));
 sg13g2_nand2_1 _1194_ (.Y(_0457_),
    .A(net53),
    .B(_0448_));
 sg13g2_a21oi_1 _1195_ (.A1(_0413_),
    .A2(_0457_),
    .Y(_0458_),
    .B1(_0298_));
 sg13g2_a221oi_1 _1196_ (.B2(_0012_),
    .C1(_0458_),
    .B1(_0456_),
    .A1(net23),
    .Y(_0459_),
    .A2(_0262_));
 sg13g2_o21ai_1 _1197_ (.B1(_0459_),
    .Y(_0460_),
    .A1(_0000_),
    .A2(_0455_));
 sg13g2_nor2b_1 _1198_ (.A(_0685_),
    .B_N(net3),
    .Y(_0461_));
 sg13g2_nor4_1 _1199_ (.A(net58),
    .B(net52),
    .C(net50),
    .D(_0461_),
    .Y(_0462_));
 sg13g2_a21oi_1 _1200_ (.A1(_0215_),
    .A2(_0414_),
    .Y(_0463_),
    .B1(_0462_));
 sg13g2_nor2_1 _1201_ (.A(net40),
    .B(_0282_),
    .Y(_0465_));
 sg13g2_nor2b_1 _1202_ (.A(net78),
    .B_N(net77),
    .Y(_0466_));
 sg13g2_a22oi_1 _1203_ (.Y(_0467_),
    .B1(_0466_),
    .B2(net66),
    .A2(_0149_),
    .A1(_0019_));
 sg13g2_nor3_1 _1204_ (.A(_0647_),
    .B(net51),
    .C(_0467_),
    .Y(_0468_));
 sg13g2_a21oi_1 _1205_ (.A1(_0449_),
    .A2(_0465_),
    .Y(_0469_),
    .B1(_0468_));
 sg13g2_nor3_1 _1206_ (.A(_0442_),
    .B(_0110_),
    .C(_0111_),
    .Y(_0470_));
 sg13g2_a21oi_1 _1207_ (.A1(_0413_),
    .A2(_0250_),
    .Y(_0471_),
    .B1(_0229_));
 sg13g2_a21oi_1 _1208_ (.A1(_0059_),
    .A2(_0182_),
    .Y(_0472_),
    .B1(_0371_));
 sg13g2_nor3_1 _1209_ (.A(_0242_),
    .B(_0147_),
    .C(_0472_),
    .Y(_0473_));
 sg13g2_and4_1 _1210_ (.A(_0593_),
    .B(_0020_),
    .C(_0669_),
    .D(_0670_),
    .X(_0474_));
 sg13g2_nand2_1 _1211_ (.Y(_0476_),
    .A(_0474_),
    .B(net56));
 sg13g2_o21ai_1 _1212_ (.B1(_0476_),
    .Y(_0477_),
    .A1(_0289_),
    .A2(_0097_));
 sg13g2_nor4_1 _1213_ (.A(_0470_),
    .B(_0471_),
    .C(_0473_),
    .D(_0477_),
    .Y(_0478_));
 sg13g2_nand4_1 _1214_ (.B(_0463_),
    .C(_0469_),
    .A(_0029_),
    .Y(_0479_),
    .D(_0478_));
 sg13g2_or4_1 _1215_ (.A(_0447_),
    .B(_0454_),
    .C(_0460_),
    .D(_0479_),
    .X(_0480_));
 sg13g2_nand4_1 _1216_ (.B(_0419_),
    .C(_0434_),
    .A(net95),
    .Y(_0481_),
    .D(_0480_));
 sg13g2_xor2_1 _1217_ (.B(_0481_),
    .A(net96),
    .X(net18));
 sg13g2_a21oi_1 _1218_ (.A1(net43),
    .A2(_0177_),
    .Y(_0482_),
    .B1(_0294_));
 sg13g2_nor2_1 _1219_ (.A(_0665_),
    .B(_0142_),
    .Y(_0483_));
 sg13g2_o21ai_1 _1220_ (.B1(_0483_),
    .Y(_0484_),
    .A1(net69),
    .A2(_0482_));
 sg13g2_a22oi_1 _1221_ (.Y(_0486_),
    .B1(_0019_),
    .B2(_0021_),
    .A2(_0024_),
    .A1(net66));
 sg13g2_nand3_1 _1222_ (.B(_0561_),
    .C(_0486_),
    .A(net69),
    .Y(_0487_));
 sg13g2_a22oi_1 _1223_ (.Y(_0488_),
    .B1(_0208_),
    .B2(net24),
    .A2(_0214_),
    .A1(_0360_));
 sg13g2_nor2_1 _1224_ (.A(net78),
    .B(net71),
    .Y(_0489_));
 sg13g2_a21o_1 _1225_ (.A2(net24),
    .A1(net28),
    .B1(_0489_),
    .X(_0490_));
 sg13g2_a21oi_1 _1226_ (.A1(net38),
    .A2(_0490_),
    .Y(_0491_),
    .B1(_0187_));
 sg13g2_o21ai_1 _1227_ (.B1(_0491_),
    .Y(_0492_),
    .A1(net29),
    .A2(_0488_));
 sg13g2_nand4_1 _1228_ (.B(_0484_),
    .C(_0487_),
    .A(net87),
    .Y(_0493_),
    .D(_0492_));
 sg13g2_nand3_1 _1229_ (.B(net37),
    .C(_0397_),
    .A(net66),
    .Y(_0494_));
 sg13g2_nand3_1 _1230_ (.B(_0128_),
    .C(_0448_),
    .A(_0182_),
    .Y(_0495_));
 sg13g2_nand2_1 _1231_ (.Y(_0497_),
    .A(net90),
    .B(net75));
 sg13g2_nand4_1 _1232_ (.B(net54),
    .C(net38),
    .A(net55),
    .Y(_0498_),
    .D(_0497_));
 sg13g2_nand3_1 _1233_ (.B(_0495_),
    .C(_0498_),
    .A(_0494_),
    .Y(_0499_));
 sg13g2_nor2_1 _1234_ (.A(net65),
    .B(net62),
    .Y(_0500_));
 sg13g2_a22oi_1 _1235_ (.Y(_0501_),
    .B1(_0129_),
    .B2(_0500_),
    .A2(net55),
    .A1(net46));
 sg13g2_nor2_1 _1236_ (.A(net29),
    .B(_0501_),
    .Y(_0502_));
 sg13g2_o21ai_1 _1237_ (.B1(net26),
    .Y(_0503_),
    .A1(_0499_),
    .A2(_0502_));
 sg13g2_a21oi_1 _1238_ (.A1(_0017_),
    .A2(_0474_),
    .Y(_0504_),
    .B1(_0238_));
 sg13g2_nor2_1 _1239_ (.A(_0133_),
    .B(_0238_),
    .Y(_0505_));
 sg13g2_or4_1 _1240_ (.A(net36),
    .B(net24),
    .C(_0504_),
    .D(_0505_),
    .X(_0506_));
 sg13g2_nor4_1 _1241_ (.A(net83),
    .B(net52),
    .C(_0210_),
    .D(_0229_),
    .Y(_0508_));
 sg13g2_nand3_1 _1242_ (.B(net54),
    .C(_0140_),
    .A(net66),
    .Y(_0509_));
 sg13g2_a221oi_1 _1243_ (.B2(_0509_),
    .C1(_0133_),
    .B1(_0117_),
    .A1(net76),
    .Y(_0510_),
    .A2(net54));
 sg13g2_nand4_1 _1244_ (.B(_0132_),
    .C(net30),
    .A(net75),
    .Y(_0511_),
    .D(_0113_));
 sg13g2_a21oi_1 _1245_ (.A1(_0240_),
    .A2(_0511_),
    .Y(_0512_),
    .B1(_0678_));
 sg13g2_nor4_1 _1246_ (.A(_0508_),
    .B(_0468_),
    .C(_0510_),
    .D(_0512_),
    .Y(_0513_));
 sg13g2_o21ai_1 _1247_ (.B1(_0160_),
    .Y(_0514_),
    .A1(_0388_),
    .A2(_0518_));
 sg13g2_nand2_1 _1248_ (.Y(_0515_),
    .A(_0437_),
    .B(_0514_));
 sg13g2_nand4_1 _1249_ (.B(_0506_),
    .C(_0513_),
    .A(_0503_),
    .Y(_0516_),
    .D(_0515_));
 sg13g2_o21ai_1 _1250_ (.B1(_0058_),
    .Y(_0517_),
    .A1(net89),
    .A2(_0056_));
 sg13g2_nor2_1 _1251_ (.A(_0010_),
    .B(_0031_),
    .Y(_0519_));
 sg13g2_a21oi_1 _1252_ (.A1(_0010_),
    .A2(net89),
    .Y(_0520_),
    .B1(_0104_));
 sg13g2_nor2_1 _1253_ (.A(_0322_),
    .B(_0002_),
    .Y(_0521_));
 sg13g2_a221oi_1 _1254_ (.B2(_0521_),
    .C1(_0462_),
    .B1(_0520_),
    .A1(_0517_),
    .Y(_0522_),
    .A2(_0519_));
 sg13g2_a21o_1 _1255_ (.A2(_0125_),
    .A1(_0122_),
    .B1(_0094_),
    .X(_0523_));
 sg13g2_nor2b_1 _1256_ (.A(_0058_),
    .B_N(_0435_),
    .Y(_0524_));
 sg13g2_and4_1 _1257_ (.A(_0679_),
    .B(_0068_),
    .C(_0437_),
    .D(_0069_),
    .X(_0525_));
 sg13g2_o21ai_1 _1258_ (.B1(net44),
    .Y(_0526_),
    .A1(_0524_),
    .A2(_0525_));
 sg13g2_and3_1 _1259_ (.X(_0527_),
    .A(_0522_),
    .B(_0523_),
    .C(_0526_));
 sg13g2_nand2_1 _1260_ (.Y(_0528_),
    .A(_0334_),
    .B(_0527_));
 sg13g2_nand4_1 _1261_ (.B(net62),
    .C(net30),
    .A(_0017_),
    .Y(_0530_),
    .D(net38));
 sg13g2_o21ai_1 _1262_ (.B1(_0530_),
    .Y(_0531_),
    .A1(_0007_),
    .A2(_0217_));
 sg13g2_nor3_1 _1263_ (.A(_0144_),
    .B(net32),
    .C(net50),
    .Y(_0532_));
 sg13g2_nor3_1 _1264_ (.A(_0234_),
    .B(_0290_),
    .C(_0002_),
    .Y(_0533_));
 sg13g2_or2_1 _1265_ (.X(_0534_),
    .B(_0533_),
    .A(_0532_));
 sg13g2_a221oi_1 _1266_ (.B2(net25),
    .C1(_0151_),
    .B1(_0534_),
    .A1(_0388_),
    .Y(_0535_),
    .A2(_0531_));
 sg13g2_a21oi_1 _1267_ (.A1(net36),
    .A2(_0196_),
    .Y(_0536_),
    .B1(_0147_));
 sg13g2_nor4_1 _1268_ (.A(net29),
    .B(net55),
    .C(_0019_),
    .D(_0536_),
    .Y(_0537_));
 sg13g2_nand4_1 _1269_ (.B(net46),
    .C(net30),
    .A(net44),
    .Y(_0538_),
    .D(net38));
 sg13g2_nand4_1 _1270_ (.B(net40),
    .C(net35),
    .A(net34),
    .Y(_0539_),
    .D(net37));
 sg13g2_a21oi_1 _1271_ (.A1(_0538_),
    .A2(_0539_),
    .Y(_0541_),
    .B1(net36));
 sg13g2_nor4_1 _1272_ (.A(_0156_),
    .B(_0161_),
    .C(_0537_),
    .D(_0541_),
    .Y(_0542_));
 sg13g2_a21oi_1 _1273_ (.A1(_0535_),
    .A2(_0542_),
    .Y(_0543_),
    .B1(_0295_));
 sg13g2_o21ai_1 _1274_ (.B1(_0543_),
    .Y(_0544_),
    .A1(_0516_),
    .A2(_0528_));
 sg13g2_a21oi_1 _1275_ (.A1(_0493_),
    .A2(_0544_),
    .Y(_0545_),
    .B1(_0203_));
 sg13g2_xnor2_1 _1276_ (.Y(net19),
    .A(net96),
    .B(_0545_));
 sg13g2_nor4_1 _1277_ (.A(_0366_),
    .B(_0678_),
    .C(net52),
    .D(_0080_),
    .Y(_0546_));
 sg13g2_nor4_1 _1278_ (.A(_0674_),
    .B(_0442_),
    .C(_0242_),
    .D(net57),
    .Y(_0547_));
 sg13g2_o21ai_1 _1279_ (.B1(_0529_),
    .Y(_0548_),
    .A1(_0546_),
    .A2(_0547_));
 sg13g2_nor3_1 _1280_ (.A(net72),
    .B(net78),
    .C(net50),
    .Y(_0549_));
 sg13g2_nor2_1 _1281_ (.A(_0031_),
    .B(_0080_),
    .Y(_0551_));
 sg13g2_o21ai_1 _1282_ (.B1(_0234_),
    .Y(_0552_),
    .A1(_0549_),
    .A2(_0551_));
 sg13g2_o21ai_1 _1283_ (.B1(_0686_),
    .Y(_0553_),
    .A1(_0205_),
    .A2(_0206_));
 sg13g2_nor3_1 _1284_ (.A(_0674_),
    .B(_0041_),
    .C(net52),
    .Y(_0554_));
 sg13g2_nor3_1 _1285_ (.A(_0235_),
    .B(_0664_),
    .C(_0141_),
    .Y(_0555_));
 sg13g2_o21ai_1 _1286_ (.B1(_0366_),
    .Y(_0556_),
    .A1(_0554_),
    .A2(_0555_));
 sg13g2_and4_1 _1287_ (.A(_0548_),
    .B(_0552_),
    .C(_0553_),
    .D(_0556_),
    .X(_0557_));
 sg13g2_nor2_1 _1288_ (.A(_0229_),
    .B(_0240_),
    .Y(_0558_));
 sg13g2_nand4_1 _1289_ (.B(_0064_),
    .C(net60),
    .A(_0132_),
    .Y(_0559_),
    .D(_0070_));
 sg13g2_o21ai_1 _1290_ (.B1(_0559_),
    .Y(_0560_),
    .A1(_0250_),
    .A2(_0097_));
 sg13g2_nor2_1 _1291_ (.A(_0033_),
    .B(net5),
    .Y(_0562_));
 sg13g2_or2_1 _1292_ (.X(_0563_),
    .B(_0035_),
    .A(_0031_));
 sg13g2_o21ai_1 _1293_ (.B1(_0194_),
    .Y(_0564_),
    .A1(_0562_),
    .A2(_0563_));
 sg13g2_nor4_1 _1294_ (.A(_0458_),
    .B(_0558_),
    .C(_0560_),
    .D(_0564_),
    .Y(_0565_));
 sg13g2_and4_1 _1295_ (.A(_0244_),
    .B(_0527_),
    .C(_0557_),
    .D(_0565_),
    .X(_0566_));
 sg13g2_o21ai_1 _1296_ (.B1(_0637_),
    .Y(_0567_),
    .A1(_0214_),
    .A2(_0327_));
 sg13g2_o21ai_1 _1297_ (.B1(_0593_),
    .Y(_0568_),
    .A1(_0322_),
    .A2(_0121_));
 sg13g2_nand3b_1 _1298_ (.B(net5),
    .C(net82),
    .Y(_0569_),
    .A_N(net63));
 sg13g2_o21ai_1 _1299_ (.B1(_0569_),
    .Y(_0570_),
    .A1(_0037_),
    .A2(_0444_));
 sg13g2_a21o_1 _1300_ (.A2(_0568_),
    .A1(_0567_),
    .B1(_0570_),
    .X(_0571_));
 sg13g2_o21ai_1 _1301_ (.B1(_0035_),
    .Y(_0573_),
    .A1(net57),
    .A2(_0032_));
 sg13g2_a221oi_1 _1302_ (.B2(net33),
    .C1(_0146_),
    .B1(_0573_),
    .A1(_0301_),
    .Y(_0574_),
    .A2(_0571_));
 sg13g2_nor2b_1 _1303_ (.A(_0159_),
    .B_N(_0574_),
    .Y(_0575_));
 sg13g2_a221oi_1 _1304_ (.B2(_0535_),
    .C1(net87),
    .B1(_0575_),
    .A1(_0116_),
    .Y(_0576_),
    .A2(_0566_));
 sg13g2_a21oi_1 _1305_ (.A1(net25),
    .A2(net67),
    .Y(_0577_),
    .B1(_0138_));
 sg13g2_o21ai_1 _1306_ (.B1(net27),
    .Y(_0578_),
    .A1(_0398_),
    .A2(_0577_));
 sg13g2_a21o_1 _1307_ (.A2(_0018_),
    .A1(_0138_),
    .B1(net31),
    .X(_0579_));
 sg13g2_nor3_1 _1308_ (.A(net28),
    .B(net42),
    .C(net27),
    .Y(_0580_));
 sg13g2_a21oi_1 _1309_ (.A1(_0068_),
    .A2(_0579_),
    .Y(_0581_),
    .B1(_0580_));
 sg13g2_nand3_1 _1310_ (.B(_0578_),
    .C(_0581_),
    .A(net88),
    .Y(_0582_));
 sg13g2_o21ai_1 _1311_ (.B1(net51),
    .Y(_0584_),
    .A1(net36),
    .A2(_0196_));
 sg13g2_mux2_1 _1312_ (.A0(_0215_),
    .A1(_0584_),
    .S(net76),
    .X(_0585_));
 sg13g2_a21oi_1 _1313_ (.A1(net92),
    .A2(_0585_),
    .Y(_0586_),
    .B1(net83));
 sg13g2_a21oi_1 _1314_ (.A1(_0582_),
    .A2(_0586_),
    .Y(_0587_),
    .B1(net97));
 sg13g2_o21ai_1 _1315_ (.B1(net95),
    .Y(_0588_),
    .A1(_0576_),
    .A2(_0587_));
 sg13g2_xor2_1 _1316_ (.B(_0588_),
    .A(_0181_),
    .X(net20));
 sg13g2_nand2_1 _1317_ (.Y(_0589_),
    .A(_0658_),
    .B(_0534_));
 sg13g2_nand3_1 _1318_ (.B(net30),
    .C(net38),
    .A(net62),
    .Y(_0590_));
 sg13g2_o21ai_1 _1319_ (.B1(_0590_),
    .Y(_0591_),
    .A1(net41),
    .A2(_0117_));
 sg13g2_o21ai_1 _1320_ (.B1(_0158_),
    .Y(_0592_),
    .A1(_0251_),
    .A2(_0590_));
 sg13g2_a21oi_1 _1321_ (.A1(net24),
    .A2(_0591_),
    .Y(_0594_),
    .B1(_0592_));
 sg13g2_nand3_1 _1322_ (.B(_0589_),
    .C(_0594_),
    .A(_0452_),
    .Y(_0595_));
 sg13g2_nand3b_1 _1323_ (.B(_0405_),
    .C(_0152_),
    .Y(_0596_),
    .A_N(_0286_));
 sg13g2_nor2_1 _1324_ (.A(_0595_),
    .B(_0596_),
    .Y(_0597_));
 sg13g2_nand2_1 _1325_ (.Y(_0598_),
    .A(net70),
    .B(net75));
 sg13g2_a22oi_1 _1326_ (.Y(_0599_),
    .B1(_0598_),
    .B2(_0222_),
    .A2(_0349_),
    .A1(_0294_));
 sg13g2_o21ai_1 _1327_ (.B1(_0289_),
    .Y(_0600_),
    .A1(_0284_),
    .A2(_0599_));
 sg13g2_nor2_1 _1328_ (.A(_0680_),
    .B(_0240_),
    .Y(_0601_));
 sg13g2_a21oi_1 _1329_ (.A1(_0680_),
    .A2(_0600_),
    .Y(_0602_),
    .B1(_0601_));
 sg13g2_nor2_1 _1330_ (.A(net50),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_nand4_1 _1331_ (.B(_0271_),
    .C(_0346_),
    .A(_0266_),
    .Y(_0605_),
    .D(_0446_));
 sg13g2_nand2b_1 _1332_ (.Y(_0606_),
    .B(net83),
    .A_N(_0147_));
 sg13g2_nand2b_1 _1333_ (.Y(_0607_),
    .B(_0333_),
    .A_N(_0049_));
 sg13g2_a21oi_1 _1334_ (.A1(_0606_),
    .A2(_0607_),
    .Y(_0608_),
    .B1(_0183_));
 sg13g2_a21oi_1 _1335_ (.A1(_0176_),
    .A2(_0106_),
    .Y(_0609_),
    .B1(_0647_));
 sg13g2_nor2_1 _1336_ (.A(_0301_),
    .B(_0242_),
    .Y(_0610_));
 sg13g2_o21ai_1 _1337_ (.B1(_0610_),
    .Y(_0611_),
    .A1(_0608_),
    .A2(_0609_));
 sg13g2_o21ai_1 _1338_ (.B1(_0604_),
    .Y(_0612_),
    .A1(net31),
    .A2(_0353_));
 sg13g2_a21o_1 _1339_ (.A2(_0612_),
    .A1(_0289_),
    .B1(_0229_),
    .X(_0613_));
 sg13g2_nand3_1 _1340_ (.B(_0611_),
    .C(_0613_),
    .A(_0552_),
    .Y(_0614_));
 sg13g2_a21oi_1 _1341_ (.A1(net75),
    .A2(_0489_),
    .Y(_0616_),
    .B1(_0148_));
 sg13g2_nor4_1 _1342_ (.A(_0377_),
    .B(net36),
    .C(_0037_),
    .D(_0616_),
    .Y(_0617_));
 sg13g2_nor2_1 _1343_ (.A(net90),
    .B(net89),
    .Y(_0618_));
 sg13g2_o21ai_1 _1344_ (.B1(net39),
    .Y(_0619_),
    .A1(net50),
    .A2(_0618_));
 sg13g2_and2_1 _1345_ (.A(_0474_),
    .B(_0619_),
    .X(_0620_));
 sg13g2_nor3_1 _1346_ (.A(_0008_),
    .B(_0617_),
    .C(_0620_),
    .Y(_0621_));
 sg13g2_nor2_1 _1347_ (.A(_0377_),
    .B(_0084_),
    .Y(_0622_));
 sg13g2_nor2_1 _1348_ (.A(_0308_),
    .B(_0240_),
    .Y(_0623_));
 sg13g2_o21ai_1 _1349_ (.B1(_0437_),
    .Y(_0624_),
    .A1(_0622_),
    .A2(_0623_));
 sg13g2_nor3_1 _1350_ (.A(_0686_),
    .B(_0023_),
    .C(_0210_),
    .Y(_0625_));
 sg13g2_a21o_1 _1351_ (.A2(_0238_),
    .A1(_0059_),
    .B1(_0625_),
    .X(_0627_));
 sg13g2_mux2_1 _1352_ (.A0(_0148_),
    .A1(_0166_),
    .S(net65),
    .X(_0628_));
 sg13g2_nor3_1 _1353_ (.A(net83),
    .B(_0149_),
    .C(_0303_),
    .Y(_0629_));
 sg13g2_nand4_1 _1354_ (.B(net60),
    .C(_0070_),
    .A(net54),
    .Y(_0630_),
    .D(_0096_));
 sg13g2_a221oi_1 _1355_ (.B2(_0630_),
    .C1(_0210_),
    .B1(_0060_),
    .A1(_0664_),
    .Y(_0631_),
    .A2(_0023_));
 sg13g2_a221oi_1 _1356_ (.B2(_0629_),
    .C1(_0631_),
    .B1(_0628_),
    .A1(_0052_),
    .Y(_0632_),
    .A2(_0627_));
 sg13g2_nand4_1 _1357_ (.B(_0621_),
    .C(_0624_),
    .A(_0526_),
    .Y(_0633_),
    .D(_0632_));
 sg13g2_nor4_1 _1358_ (.A(_0603_),
    .B(_0605_),
    .C(_0614_),
    .D(_0633_),
    .Y(_0634_));
 sg13g2_a21oi_1 _1359_ (.A1(net26),
    .A2(_0294_),
    .Y(_0635_),
    .B1(net40));
 sg13g2_o21ai_1 _1360_ (.B1(_0165_),
    .Y(_0636_),
    .A1(net47),
    .A2(_0635_));
 sg13g2_a21oi_1 _1361_ (.A1(net24),
    .A2(_0068_),
    .Y(_0638_),
    .B1(_0128_));
 sg13g2_a21oi_1 _1362_ (.A1(net69),
    .A2(net24),
    .Y(_0639_),
    .B1(_0296_));
 sg13g2_o21ai_1 _1363_ (.B1(_0639_),
    .Y(_0640_),
    .A1(net45),
    .A2(_0638_));
 sg13g2_a21oi_1 _1364_ (.A1(net25),
    .A2(_0636_),
    .Y(_0641_),
    .B1(_0640_));
 sg13g2_o21ai_1 _1365_ (.B1(_0147_),
    .Y(_0642_),
    .A1(_0104_),
    .A2(_0223_));
 sg13g2_nand3_1 _1366_ (.B(net6),
    .C(net87),
    .A(net92),
    .Y(_0643_));
 sg13g2_o21ai_1 _1367_ (.B1(net95),
    .Y(_0644_),
    .A1(_0642_),
    .A2(_0643_));
 sg13g2_nor4_1 _1368_ (.A(_0597_),
    .B(_0634_),
    .C(_0641_),
    .D(_0644_),
    .Y(_0645_));
 sg13g2_xnor2_1 _1369_ (.Y(net21),
    .A(_0181_),
    .B(_0645_));
 sg13g2_o21ai_1 _1370_ (.B1(_0012_),
    .Y(_0646_),
    .A1(_0118_),
    .A2(net27));
 sg13g2_nand3_1 _1371_ (.B(_0049_),
    .C(_0646_),
    .A(net61),
    .Y(_0648_));
 sg13g2_a21oi_1 _1372_ (.A1(net8),
    .A2(_0648_),
    .Y(_0649_),
    .B1(net88));
 sg13g2_nand2b_1 _1373_ (.Y(_0650_),
    .B(_0321_),
    .A_N(_0157_));
 sg13g2_nor3_1 _1374_ (.A(net27),
    .B(net92),
    .C(_0650_),
    .Y(_0651_));
 sg13g2_nor2_1 _1375_ (.A(_0649_),
    .B(_0651_),
    .Y(_0652_));
 sg13g2_nor2_1 _1376_ (.A(net88),
    .B(net96),
    .Y(_0653_));
 sg13g2_nand2_1 _1377_ (.Y(_0654_),
    .A(net95),
    .B(_0648_));
 sg13g2_a22oi_1 _1378_ (.Y(_0655_),
    .B1(_0653_),
    .B2(_0654_),
    .A2(_0652_),
    .A1(_0192_));
 sg13g2_o21ai_1 _1379_ (.B1(_0018_),
    .Y(_0656_),
    .A1(net45),
    .A2(net66));
 sg13g2_a21oi_1 _1380_ (.A1(_0068_),
    .A2(_0580_),
    .Y(_0657_),
    .B1(net34));
 sg13g2_nand2_1 _1381_ (.Y(_0659_),
    .A(_0656_),
    .B(_0657_));
 sg13g2_nor2_1 _1382_ (.A(_0203_),
    .B(net88),
    .Y(_0660_));
 sg13g2_a221oi_1 _1383_ (.B2(_0660_),
    .C1(net87),
    .B1(_0650_),
    .A1(net88),
    .Y(_0661_),
    .A2(_0659_));
 sg13g2_a21oi_1 _1384_ (.A1(net87),
    .A2(_0655_),
    .Y(net22),
    .B1(_0661_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_buf_1 _1386_ (.A(net10),
    .X(net11));
 sg13g2_buf_1 _1387_ (.A(net10),
    .X(net12));
 sg13g2_buf_1 _1388_ (.A(net98),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1389_ (.A(net99),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1390_ (.A(net100),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1391_ (.A(net101),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1392_ (.A(net102),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1393_ (.A(net103),
    .X(uio_oe[7]));
 sg13g2_buf_1 _1394_ (.A(net104),
    .X(uio_out[2]));
 sg13g2_buf_1 _1395_ (.A(net105),
    .X(uio_out[3]));
 sg13g2_buf_1 _1396_ (.A(net106),
    .X(uio_out[4]));
 sg13g2_buf_1 _1397_ (.A(net107),
    .X(uio_out[5]));
 sg13g2_buf_1 _1398_ (.A(net108),
    .X(uio_out[6]));
 sg13g2_buf_1 _1399_ (.A(net109),
    .X(uio_out[7]));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[4]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[7]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[0]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[1]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[2]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[3]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[5]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[6]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[7]),
    .X(net10));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_oe[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[0]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[1]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[0]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[1]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[2]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[3]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[4]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[5]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[6]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout23 (.A(_0089_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0077_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0658_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0388_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0257_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0184_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0183_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0153_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0140_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0138_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0136_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0133_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0113_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0081_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0048_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0047_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0032_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0017_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0676_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0647_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0615_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0377_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0301_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0246_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0284_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0176_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0144_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0103_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0094_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0079_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0070_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0064_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0062_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0052_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0044_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0041_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0010_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0004_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0000_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0675_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0670_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0637_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0604_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0485_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0442_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0366_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0333_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0290_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0235_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0020_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0011_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0005_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0686_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0680_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0674_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0669_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0663_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0662_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0626_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0593_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0540_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0355_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0279_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0224_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0295_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0194_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0685_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0679_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0673_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0550_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_0409_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_0213_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_0192_),
    .X(net95));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(_0181_));
 sg13g2_buf_2 fanout97 (.A(_0170_),
    .X(net97));
 sg13g2_tielo _1388__98 (.L_LO(net98));
 sg13g2_tielo _1389__99 (.L_LO(net99));
 sg13g2_tielo _1390__100 (.L_LO(net100));
 sg13g2_tielo _1391__101 (.L_LO(net101));
 sg13g2_tielo _1392__102 (.L_LO(net102));
 sg13g2_tielo _1393__103 (.L_LO(net103));
 sg13g2_tielo _1394__104 (.L_LO(net104));
 sg13g2_tielo _1395__105 (.L_LO(net105));
 sg13g2_tielo _1396__106 (.L_LO(net106));
 sg13g2_tielo _1397__107 (.L_LO(net107));
 sg13g2_tielo _1398__108 (.L_LO(net108));
 sg13g2_tielo _1399__109 (.L_LO(net109));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_17_427 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_fill_2 FILLER_18_427 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_4 FILLER_19_273 ();
 sg13g2_fill_2 FILLER_19_277 ();
 sg13g2_decap_8 FILLER_19_292 ();
 sg13g2_fill_2 FILLER_19_299 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_307 ();
 sg13g2_decap_8 FILLER_19_314 ();
 sg13g2_fill_2 FILLER_19_321 ();
 sg13g2_fill_1 FILLER_19_323 ();
 sg13g2_fill_1 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_19_370 ();
 sg13g2_decap_8 FILLER_19_377 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_8 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_19_412 ();
 sg13g2_decap_8 FILLER_19_419 ();
 sg13g2_decap_4 FILLER_19_426 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_fill_1 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_4 FILLER_20_189 ();
 sg13g2_fill_1 FILLER_20_193 ();
 sg13g2_decap_4 FILLER_20_199 ();
 sg13g2_fill_1 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_209 ();
 sg13g2_decap_8 FILLER_20_216 ();
 sg13g2_decap_8 FILLER_20_223 ();
 sg13g2_fill_2 FILLER_20_230 ();
 sg13g2_fill_1 FILLER_20_232 ();
 sg13g2_decap_4 FILLER_20_243 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_fill_1 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_268 ();
 sg13g2_fill_1 FILLER_20_275 ();
 sg13g2_fill_2 FILLER_20_284 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_fill_2 FILLER_20_291 ();
 sg13g2_fill_1 FILLER_20_313 ();
 sg13g2_fill_2 FILLER_20_322 ();
 sg13g2_decap_4 FILLER_20_328 ();
 sg13g2_fill_2 FILLER_20_337 ();
 sg13g2_fill_1 FILLER_20_339 ();
 sg13g2_decap_8 FILLER_20_353 ();
 sg13g2_fill_2 FILLER_20_360 ();
 sg13g2_fill_1 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_decap_8 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_20_415 ();
 sg13g2_decap_8 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_4 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_130 ();
 sg13g2_decap_4 FILLER_21_137 ();
 sg13g2_fill_1 FILLER_21_141 ();
 sg13g2_decap_4 FILLER_21_146 ();
 sg13g2_decap_8 FILLER_21_155 ();
 sg13g2_decap_8 FILLER_21_162 ();
 sg13g2_decap_8 FILLER_21_169 ();
 sg13g2_fill_1 FILLER_21_176 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_fill_1 FILLER_21_189 ();
 sg13g2_decap_4 FILLER_21_213 ();
 sg13g2_fill_2 FILLER_21_217 ();
 sg13g2_decap_4 FILLER_21_223 ();
 sg13g2_fill_1 FILLER_21_227 ();
 sg13g2_decap_8 FILLER_21_247 ();
 sg13g2_decap_8 FILLER_21_254 ();
 sg13g2_decap_8 FILLER_21_261 ();
 sg13g2_decap_4 FILLER_21_268 ();
 sg13g2_decap_8 FILLER_21_277 ();
 sg13g2_fill_2 FILLER_21_284 ();
 sg13g2_fill_1 FILLER_21_286 ();
 sg13g2_fill_1 FILLER_21_309 ();
 sg13g2_decap_4 FILLER_21_318 ();
 sg13g2_fill_2 FILLER_21_322 ();
 sg13g2_fill_2 FILLER_21_328 ();
 sg13g2_decap_4 FILLER_21_337 ();
 sg13g2_fill_2 FILLER_21_341 ();
 sg13g2_fill_1 FILLER_21_365 ();
 sg13g2_decap_4 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_decap_8 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_21_415 ();
 sg13g2_decap_8 FILLER_21_422 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_4 FILLER_22_105 ();
 sg13g2_decap_4 FILLER_22_122 ();
 sg13g2_fill_1 FILLER_22_136 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_154 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_fill_1 FILLER_22_175 ();
 sg13g2_fill_2 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_188 ();
 sg13g2_fill_2 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_219 ();
 sg13g2_decap_4 FILLER_22_225 ();
 sg13g2_fill_2 FILLER_22_253 ();
 sg13g2_decap_4 FILLER_22_263 ();
 sg13g2_fill_1 FILLER_22_272 ();
 sg13g2_fill_1 FILLER_22_278 ();
 sg13g2_fill_2 FILLER_22_311 ();
 sg13g2_fill_1 FILLER_22_313 ();
 sg13g2_fill_1 FILLER_22_325 ();
 sg13g2_decap_4 FILLER_22_337 ();
 sg13g2_fill_1 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_fill_1 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_22_414 ();
 sg13g2_decap_8 FILLER_22_421 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_4 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_102 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_fill_1 FILLER_23_110 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_fill_1 FILLER_23_122 ();
 sg13g2_fill_1 FILLER_23_154 ();
 sg13g2_fill_1 FILLER_23_164 ();
 sg13g2_decap_4 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_193 ();
 sg13g2_decap_4 FILLER_23_210 ();
 sg13g2_fill_2 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_221 ();
 sg13g2_fill_2 FILLER_23_248 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_decap_4 FILLER_23_284 ();
 sg13g2_fill_1 FILLER_23_288 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_decap_4 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_310 ();
 sg13g2_fill_1 FILLER_23_326 ();
 sg13g2_fill_2 FILLER_23_352 ();
 sg13g2_fill_1 FILLER_23_358 ();
 sg13g2_decap_4 FILLER_23_369 ();
 sg13g2_fill_2 FILLER_23_378 ();
 sg13g2_fill_1 FILLER_23_380 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_decap_8 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_23_414 ();
 sg13g2_decap_8 FILLER_23_421 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_91 ();
 sg13g2_fill_2 FILLER_24_97 ();
 sg13g2_fill_1 FILLER_24_99 ();
 sg13g2_fill_2 FILLER_24_115 ();
 sg13g2_fill_1 FILLER_24_130 ();
 sg13g2_fill_1 FILLER_24_135 ();
 sg13g2_decap_8 FILLER_24_145 ();
 sg13g2_fill_2 FILLER_24_152 ();
 sg13g2_fill_1 FILLER_24_165 ();
 sg13g2_decap_4 FILLER_24_184 ();
 sg13g2_decap_8 FILLER_24_211 ();
 sg13g2_fill_2 FILLER_24_218 ();
 sg13g2_fill_1 FILLER_24_220 ();
 sg13g2_decap_4 FILLER_24_227 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_fill_2 FILLER_24_257 ();
 sg13g2_fill_1 FILLER_24_274 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_fill_2 FILLER_24_293 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_fill_2 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_fill_2 FILLER_24_364 ();
 sg13g2_fill_1 FILLER_24_374 ();
 sg13g2_fill_2 FILLER_24_388 ();
 sg13g2_fill_1 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_8 FILLER_24_403 ();
 sg13g2_decap_8 FILLER_24_410 ();
 sg13g2_decap_8 FILLER_24_417 ();
 sg13g2_decap_4 FILLER_24_424 ();
 sg13g2_fill_2 FILLER_24_428 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_4 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_161 ();
 sg13g2_decap_4 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_190 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_4 FILLER_25_210 ();
 sg13g2_fill_1 FILLER_25_214 ();
 sg13g2_decap_4 FILLER_25_224 ();
 sg13g2_fill_2 FILLER_25_232 ();
 sg13g2_decap_4 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_267 ();
 sg13g2_fill_1 FILLER_25_280 ();
 sg13g2_fill_2 FILLER_25_298 ();
 sg13g2_fill_2 FILLER_25_305 ();
 sg13g2_fill_1 FILLER_25_335 ();
 sg13g2_fill_1 FILLER_25_341 ();
 sg13g2_decap_4 FILLER_25_370 ();
 sg13g2_decap_4 FILLER_25_379 ();
 sg13g2_decap_4 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_8 FILLER_25_404 ();
 sg13g2_decap_8 FILLER_25_411 ();
 sg13g2_decap_8 FILLER_25_418 ();
 sg13g2_decap_4 FILLER_25_425 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_fill_2 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_103 ();
 sg13g2_fill_1 FILLER_26_110 ();
 sg13g2_fill_1 FILLER_26_121 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_2 FILLER_26_139 ();
 sg13g2_fill_2 FILLER_26_146 ();
 sg13g2_fill_2 FILLER_26_199 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_decap_4 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_243 ();
 sg13g2_decap_4 FILLER_26_269 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_fill_2 FILLER_26_321 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_fill_1 FILLER_26_347 ();
 sg13g2_fill_1 FILLER_26_361 ();
 sg13g2_decap_4 FILLER_26_389 ();
 sg13g2_fill_1 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_26_414 ();
 sg13g2_decap_8 FILLER_26_421 ();
 sg13g2_fill_2 FILLER_26_428 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_4 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_88 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_4 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_124 ();
 sg13g2_fill_2 FILLER_27_146 ();
 sg13g2_fill_1 FILLER_27_148 ();
 sg13g2_decap_4 FILLER_27_187 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_decap_8 FILLER_27_197 ();
 sg13g2_decap_4 FILLER_27_204 ();
 sg13g2_fill_1 FILLER_27_208 ();
 sg13g2_decap_4 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_218 ();
 sg13g2_fill_1 FILLER_27_227 ();
 sg13g2_fill_2 FILLER_27_247 ();
 sg13g2_decap_8 FILLER_27_254 ();
 sg13g2_fill_2 FILLER_27_261 ();
 sg13g2_fill_2 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_282 ();
 sg13g2_fill_2 FILLER_27_289 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_fill_2 FILLER_27_320 ();
 sg13g2_fill_1 FILLER_27_322 ();
 sg13g2_fill_2 FILLER_27_360 ();
 sg13g2_fill_1 FILLER_27_362 ();
 sg13g2_fill_2 FILLER_27_376 ();
 sg13g2_fill_1 FILLER_27_378 ();
 sg13g2_fill_1 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_27_415 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_fill_2 FILLER_28_91 ();
 sg13g2_fill_1 FILLER_28_97 ();
 sg13g2_fill_2 FILLER_28_103 ();
 sg13g2_fill_1 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_fill_1 FILLER_28_148 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_4 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_fill_1 FILLER_28_211 ();
 sg13g2_decap_4 FILLER_28_217 ();
 sg13g2_fill_2 FILLER_28_221 ();
 sg13g2_fill_2 FILLER_28_240 ();
 sg13g2_decap_4 FILLER_28_248 ();
 sg13g2_decap_4 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_281 ();
 sg13g2_fill_2 FILLER_28_288 ();
 sg13g2_fill_1 FILLER_28_290 ();
 sg13g2_fill_1 FILLER_28_301 ();
 sg13g2_fill_2 FILLER_28_317 ();
 sg13g2_fill_1 FILLER_28_323 ();
 sg13g2_fill_2 FILLER_28_339 ();
 sg13g2_fill_1 FILLER_28_341 ();
 sg13g2_fill_2 FILLER_28_350 ();
 sg13g2_fill_1 FILLER_28_357 ();
 sg13g2_fill_1 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_410 ();
 sg13g2_decap_8 FILLER_28_417 ();
 sg13g2_decap_4 FILLER_28_424 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_fill_1 FILLER_29_84 ();
 sg13g2_fill_1 FILLER_29_89 ();
 sg13g2_fill_1 FILLER_29_115 ();
 sg13g2_fill_2 FILLER_29_121 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_decap_4 FILLER_29_132 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_fill_2 FILLER_29_148 ();
 sg13g2_fill_1 FILLER_29_150 ();
 sg13g2_fill_1 FILLER_29_161 ();
 sg13g2_fill_1 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_182 ();
 sg13g2_fill_2 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_decap_4 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_220 ();
 sg13g2_decap_4 FILLER_29_232 ();
 sg13g2_decap_8 FILLER_29_242 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_decap_4 FILLER_29_254 ();
 sg13g2_fill_1 FILLER_29_258 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_267 ();
 sg13g2_decap_4 FILLER_29_273 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_decap_4 FILLER_29_283 ();
 sg13g2_decap_8 FILLER_29_303 ();
 sg13g2_decap_4 FILLER_29_310 ();
 sg13g2_fill_2 FILLER_29_314 ();
 sg13g2_fill_1 FILLER_29_321 ();
 sg13g2_fill_2 FILLER_29_326 ();
 sg13g2_fill_1 FILLER_29_328 ();
 sg13g2_fill_2 FILLER_29_380 ();
 sg13g2_fill_2 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_414 ();
 sg13g2_decap_8 FILLER_29_421 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_fill_2 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_116 ();
 sg13g2_fill_1 FILLER_30_132 ();
 sg13g2_fill_2 FILLER_30_153 ();
 sg13g2_fill_1 FILLER_30_155 ();
 sg13g2_decap_4 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_218 ();
 sg13g2_decap_8 FILLER_30_225 ();
 sg13g2_fill_1 FILLER_30_272 ();
 sg13g2_fill_2 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_decap_8 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_318 ();
 sg13g2_fill_2 FILLER_30_324 ();
 sg13g2_fill_1 FILLER_30_347 ();
 sg13g2_fill_1 FILLER_30_358 ();
 sg13g2_fill_1 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_98 ();
 sg13g2_fill_1 FILLER_31_104 ();
 sg13g2_fill_2 FILLER_31_115 ();
 sg13g2_decap_8 FILLER_31_127 ();
 sg13g2_fill_1 FILLER_31_147 ();
 sg13g2_fill_1 FILLER_31_157 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_fill_1 FILLER_31_175 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_decap_4 FILLER_31_196 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_decap_8 FILLER_31_206 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_fill_2 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_241 ();
 sg13g2_decap_4 FILLER_31_252 ();
 sg13g2_fill_2 FILLER_31_256 ();
 sg13g2_decap_4 FILLER_31_263 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_fill_2 FILLER_31_287 ();
 sg13g2_fill_2 FILLER_31_308 ();
 sg13g2_fill_1 FILLER_31_310 ();
 sg13g2_fill_1 FILLER_31_316 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_339 ();
 sg13g2_decap_4 FILLER_31_354 ();
 sg13g2_fill_2 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_4 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_416 ();
 sg13g2_decap_8 FILLER_31_423 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_4 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_81 ();
 sg13g2_fill_1 FILLER_32_114 ();
 sg13g2_decap_4 FILLER_32_132 ();
 sg13g2_decap_4 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_144 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_fill_2 FILLER_32_216 ();
 sg13g2_decap_8 FILLER_32_230 ();
 sg13g2_fill_1 FILLER_32_241 ();
 sg13g2_decap_8 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_284 ();
 sg13g2_fill_2 FILLER_32_291 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_fill_2 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_319 ();
 sg13g2_decap_4 FILLER_32_326 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_decap_4 FILLER_32_359 ();
 sg13g2_fill_1 FILLER_32_363 ();
 sg13g2_decap_4 FILLER_32_369 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_fill_2 FILLER_32_385 ();
 sg13g2_fill_1 FILLER_32_387 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_decap_8 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_32_415 ();
 sg13g2_decap_8 FILLER_32_422 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_fill_2 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_90 ();
 sg13g2_decap_4 FILLER_33_100 ();
 sg13g2_fill_2 FILLER_33_104 ();
 sg13g2_decap_4 FILLER_33_110 ();
 sg13g2_decap_8 FILLER_33_123 ();
 sg13g2_decap_8 FILLER_33_130 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_fill_1 FILLER_33_153 ();
 sg13g2_decap_4 FILLER_33_159 ();
 sg13g2_fill_1 FILLER_33_163 ();
 sg13g2_fill_2 FILLER_33_174 ();
 sg13g2_fill_1 FILLER_33_176 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_fill_1 FILLER_33_198 ();
 sg13g2_decap_4 FILLER_33_212 ();
 sg13g2_decap_4 FILLER_33_222 ();
 sg13g2_fill_2 FILLER_33_226 ();
 sg13g2_decap_8 FILLER_33_236 ();
 sg13g2_decap_8 FILLER_33_243 ();
 sg13g2_decap_8 FILLER_33_250 ();
 sg13g2_fill_2 FILLER_33_257 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_265 ();
 sg13g2_decap_8 FILLER_33_272 ();
 sg13g2_decap_4 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_fill_2 FILLER_33_288 ();
 sg13g2_fill_1 FILLER_33_290 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_fill_2 FILLER_33_318 ();
 sg13g2_fill_2 FILLER_33_351 ();
 sg13g2_fill_1 FILLER_33_373 ();
 sg13g2_fill_1 FILLER_33_379 ();
 sg13g2_decap_4 FILLER_33_384 ();
 sg13g2_decap_8 FILLER_33_395 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_33_409 ();
 sg13g2_decap_8 FILLER_33_416 ();
 sg13g2_decap_8 FILLER_33_423 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_4 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_81 ();
 sg13g2_decap_8 FILLER_34_100 ();
 sg13g2_fill_2 FILLER_34_107 ();
 sg13g2_decap_4 FILLER_34_117 ();
 sg13g2_fill_1 FILLER_34_121 ();
 sg13g2_fill_2 FILLER_34_132 ();
 sg13g2_decap_4 FILLER_34_143 ();
 sg13g2_fill_2 FILLER_34_175 ();
 sg13g2_fill_2 FILLER_34_191 ();
 sg13g2_decap_4 FILLER_34_207 ();
 sg13g2_fill_2 FILLER_34_211 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_decap_4 FILLER_34_223 ();
 sg13g2_fill_1 FILLER_34_227 ();
 sg13g2_fill_1 FILLER_34_233 ();
 sg13g2_fill_1 FILLER_34_248 ();
 sg13g2_fill_2 FILLER_34_254 ();
 sg13g2_fill_1 FILLER_34_261 ();
 sg13g2_fill_2 FILLER_34_287 ();
 sg13g2_fill_2 FILLER_34_299 ();
 sg13g2_fill_1 FILLER_34_301 ();
 sg13g2_fill_2 FILLER_34_306 ();
 sg13g2_fill_1 FILLER_34_368 ();
 sg13g2_fill_1 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_403 ();
 sg13g2_fill_1 FILLER_34_410 ();
 sg13g2_decap_4 FILLER_34_424 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_fill_2 FILLER_35_77 ();
 sg13g2_decap_4 FILLER_35_92 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_fill_2 FILLER_35_106 ();
 sg13g2_fill_1 FILLER_35_108 ();
 sg13g2_fill_2 FILLER_35_119 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_132 ();
 sg13g2_decap_8 FILLER_35_139 ();
 sg13g2_decap_8 FILLER_35_146 ();
 sg13g2_fill_2 FILLER_35_170 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_decap_8 FILLER_35_183 ();
 sg13g2_decap_4 FILLER_35_190 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_decap_8 FILLER_35_221 ();
 sg13g2_fill_1 FILLER_35_238 ();
 sg13g2_fill_1 FILLER_35_244 ();
 sg13g2_fill_1 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_decap_8 FILLER_35_262 ();
 sg13g2_fill_2 FILLER_35_269 ();
 sg13g2_fill_1 FILLER_35_271 ();
 sg13g2_fill_2 FILLER_35_289 ();
 sg13g2_decap_4 FILLER_35_295 ();
 sg13g2_fill_2 FILLER_35_304 ();
 sg13g2_fill_1 FILLER_35_317 ();
 sg13g2_fill_1 FILLER_35_322 ();
 sg13g2_fill_1 FILLER_35_328 ();
 sg13g2_decap_4 FILLER_35_334 ();
 sg13g2_fill_2 FILLER_35_338 ();
 sg13g2_fill_2 FILLER_35_348 ();
 sg13g2_fill_2 FILLER_35_364 ();
 sg13g2_decap_4 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_8 FILLER_35_404 ();
 sg13g2_decap_8 FILLER_35_411 ();
 sg13g2_decap_8 FILLER_35_418 ();
 sg13g2_decap_4 FILLER_35_425 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_fill_2 FILLER_36_105 ();
 sg13g2_decap_4 FILLER_36_117 ();
 sg13g2_fill_2 FILLER_36_146 ();
 sg13g2_fill_1 FILLER_36_148 ();
 sg13g2_decap_8 FILLER_36_153 ();
 sg13g2_fill_1 FILLER_36_160 ();
 sg13g2_fill_2 FILLER_36_166 ();
 sg13g2_fill_1 FILLER_36_168 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_fill_2 FILLER_36_192 ();
 sg13g2_fill_1 FILLER_36_194 ();
 sg13g2_fill_1 FILLER_36_200 ();
 sg13g2_decap_4 FILLER_36_211 ();
 sg13g2_fill_2 FILLER_36_215 ();
 sg13g2_decap_8 FILLER_36_222 ();
 sg13g2_fill_2 FILLER_36_229 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_255 ();
 sg13g2_decap_8 FILLER_36_262 ();
 sg13g2_decap_8 FILLER_36_269 ();
 sg13g2_fill_1 FILLER_36_276 ();
 sg13g2_fill_1 FILLER_36_291 ();
 sg13g2_fill_2 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_297 ();
 sg13g2_decap_8 FILLER_36_307 ();
 sg13g2_fill_1 FILLER_36_314 ();
 sg13g2_decap_4 FILLER_36_318 ();
 sg13g2_fill_1 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_327 ();
 sg13g2_fill_1 FILLER_36_334 ();
 sg13g2_decap_4 FILLER_36_349 ();
 sg13g2_fill_1 FILLER_36_358 ();
 sg13g2_fill_1 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_36_409 ();
 sg13g2_decap_8 FILLER_36_416 ();
 sg13g2_decap_8 FILLER_36_423 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_84 ();
 sg13g2_fill_1 FILLER_37_86 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_4 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_124 ();
 sg13g2_decap_4 FILLER_37_131 ();
 sg13g2_fill_2 FILLER_37_147 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_decap_4 FILLER_37_154 ();
 sg13g2_fill_1 FILLER_37_158 ();
 sg13g2_fill_1 FILLER_37_163 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_202 ();
 sg13g2_decap_4 FILLER_37_219 ();
 sg13g2_fill_1 FILLER_37_231 ();
 sg13g2_decap_4 FILLER_37_240 ();
 sg13g2_fill_1 FILLER_37_244 ();
 sg13g2_fill_1 FILLER_37_265 ();
 sg13g2_fill_2 FILLER_37_288 ();
 sg13g2_decap_4 FILLER_37_299 ();
 sg13g2_fill_1 FILLER_37_303 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_4 FILLER_37_315 ();
 sg13g2_fill_1 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_324 ();
 sg13g2_decap_4 FILLER_37_331 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_fill_2 FILLER_37_341 ();
 sg13g2_fill_2 FILLER_37_356 ();
 sg13g2_fill_1 FILLER_37_358 ();
 sg13g2_fill_2 FILLER_37_363 ();
 sg13g2_fill_1 FILLER_37_365 ();
 sg13g2_fill_2 FILLER_37_379 ();
 sg13g2_fill_1 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_decap_8 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_37_414 ();
 sg13g2_decap_8 FILLER_37_421 ();
 sg13g2_fill_2 FILLER_37_428 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_4 FILLER_38_70 ();
 sg13g2_fill_2 FILLER_38_134 ();
 sg13g2_fill_1 FILLER_38_144 ();
 sg13g2_fill_1 FILLER_38_181 ();
 sg13g2_decap_8 FILLER_38_186 ();
 sg13g2_fill_2 FILLER_38_213 ();
 sg13g2_fill_2 FILLER_38_227 ();
 sg13g2_fill_2 FILLER_38_241 ();
 sg13g2_fill_2 FILLER_38_255 ();
 sg13g2_fill_1 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_262 ();
 sg13g2_fill_2 FILLER_38_267 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_323 ();
 sg13g2_decap_8 FILLER_38_330 ();
 sg13g2_decap_8 FILLER_38_337 ();
 sg13g2_fill_2 FILLER_38_344 ();
 sg13g2_fill_1 FILLER_38_346 ();
 sg13g2_decap_8 FILLER_38_351 ();
 sg13g2_fill_2 FILLER_38_358 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_fill_2 FILLER_38_371 ();
 sg13g2_fill_1 FILLER_38_373 ();
 sg13g2_fill_2 FILLER_38_387 ();
 sg13g2_fill_1 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_403 ();
 sg13g2_decap_8 FILLER_38_410 ();
 sg13g2_decap_8 FILLER_38_417 ();
 sg13g2_decap_4 FILLER_38_424 ();
 sg13g2_fill_2 FILLER_38_428 ();
endmodule
