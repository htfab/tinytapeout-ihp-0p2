module tt_um_NicklausThompson_SkyKing (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire BNC_trig;
 wire \BNC_x[0] ;
 wire \BNC_x[1] ;
 wire \BNC_x[2] ;
 wire \BNC_x[3] ;
 wire \BNC_x[4] ;
 wire \BNC_x[5] ;
 wire \BNC_x[6] ;
 wire \BNC_x[7] ;
 wire \BNC_y[0] ;
 wire \BNC_y[1] ;
 wire \BNC_y[2] ;
 wire \BNC_y[3] ;
 wire \BNC_y[4] ;
 wire \BNC_y[5] ;
 wire \BNC_y[6] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire clknet_0_clk;
 wire \bnc_image_generator.counter[0] ;
 wire \bnc_image_generator.counter[1] ;
 wire \bnc_image_generator.counter[2] ;
 wire \bnc_image_generator.counter[4] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \vga_image_generator.character_hold[0] ;
 wire \vga_image_generator.character_hold[10] ;
 wire \vga_image_generator.character_hold[11] ;
 wire \vga_image_generator.character_hold[12] ;
 wire \vga_image_generator.character_hold[13] ;
 wire \vga_image_generator.character_hold[14] ;
 wire \vga_image_generator.character_hold[15] ;
 wire \vga_image_generator.character_hold[16] ;
 wire \vga_image_generator.character_hold[17] ;
 wire \vga_image_generator.character_hold[1] ;
 wire \vga_image_generator.character_hold[2] ;
 wire \vga_image_generator.character_hold[3] ;
 wire \vga_image_generator.character_hold[4] ;
 wire \vga_image_generator.character_hold[5] ;
 wire \vga_image_generator.character_hold[6] ;
 wire \vga_image_generator.character_hold[7] ;
 wire \vga_image_generator.character_hold[8] ;
 wire \vga_image_generator.character_hold[9] ;
 wire \vga_image_generator.counter[0] ;
 wire \vga_image_generator.counter[10] ;
 wire \vga_image_generator.counter[11] ;
 wire \vga_image_generator.counter[12] ;
 wire \vga_image_generator.counter[13] ;
 wire \vga_image_generator.counter[14] ;
 wire \vga_image_generator.counter[15] ;
 wire \vga_image_generator.counter[16] ;
 wire \vga_image_generator.counter[17] ;
 wire \vga_image_generator.counter[18] ;
 wire \vga_image_generator.counter[19] ;
 wire \vga_image_generator.counter[1] ;
 wire \vga_image_generator.counter[20] ;
 wire \vga_image_generator.counter[21] ;
 wire \vga_image_generator.counter[22] ;
 wire \vga_image_generator.counter[23] ;
 wire \vga_image_generator.counter[24] ;
 wire \vga_image_generator.counter[2] ;
 wire \vga_image_generator.counter[3] ;
 wire \vga_image_generator.counter[4] ;
 wire \vga_image_generator.counter[5] ;
 wire \vga_image_generator.counter[6] ;
 wire \vga_image_generator.counter[7] ;
 wire \vga_image_generator.counter[8] ;
 wire \vga_image_generator.counter[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_inv_1 _0874_ (.Y(_0107_),
    .A(\hvsync_gen.vpos[1] ));
 sg13g2_buf_1 _0875_ (.A(\hvsync_gen.vpos[2] ),
    .X(_0108_));
 sg13g2_buf_8 _0876_ (.A(\hvsync_gen.vpos[3] ),
    .X(_0109_));
 sg13g2_inv_2 _0877_ (.Y(_0110_),
    .A(_0109_));
 sg13g2_nor2_1 _0878_ (.A(net68),
    .B(_0110_),
    .Y(_0111_));
 sg13g2_buf_1 _0879_ (.A(\hvsync_gen.vpos[8] ),
    .X(_0112_));
 sg13g2_inv_2 _0880_ (.Y(_0113_),
    .A(net67));
 sg13g2_nor2_1 _0881_ (.A(_0113_),
    .B(\hvsync_gen.vpos[9] ),
    .Y(_0114_));
 sg13g2_nand2b_1 _0882_ (.Y(_0115_),
    .B(\hvsync_gen.vpos[5] ),
    .A_N(\hvsync_gen.vpos[4] ));
 sg13g2_buf_2 _0883_ (.A(_0115_),
    .X(_0116_));
 sg13g2_a21oi_1 _0884_ (.A1(\hvsync_gen.vpos[0] ),
    .A2(_0021_),
    .Y(_0117_),
    .B1(_0116_));
 sg13g2_nand3_1 _0885_ (.B(_0114_),
    .C(_0117_),
    .A(_0111_),
    .Y(_0118_));
 sg13g2_buf_1 _0886_ (.A(\hvsync_gen.vpos[7] ),
    .X(_0119_));
 sg13g2_buf_1 _0887_ (.A(\hvsync_gen.vpos[6] ),
    .X(_0120_));
 sg13g2_nand2_1 _0888_ (.Y(_0121_),
    .A(net66),
    .B(net65));
 sg13g2_nor3_1 _0889_ (.A(_0107_),
    .B(_0118_),
    .C(_0121_),
    .Y(_0016_));
 sg13g2_buf_1 _0890_ (.A(\hvsync_gen.hpos[9] ),
    .X(_0122_));
 sg13g2_inv_2 _0891_ (.Y(_0123_),
    .A(_0122_));
 sg13g2_buf_2 _0892_ (.A(_0022_),
    .X(_0124_));
 sg13g2_buf_2 _0893_ (.A(\hvsync_gen.hpos[6] ),
    .X(_0125_));
 sg13g2_buf_8 _0894_ (.A(_0125_),
    .X(_0126_));
 sg13g2_buf_1 _0895_ (.A(\hvsync_gen.hpos[5] ),
    .X(_0127_));
 sg13g2_buf_1 _0896_ (.A(\hvsync_gen.hpos[4] ),
    .X(_0128_));
 sg13g2_and2_1 _0897_ (.A(net64),
    .B(_0128_),
    .X(_0129_));
 sg13g2_buf_1 _0898_ (.A(_0129_),
    .X(_0130_));
 sg13g2_buf_1 _0899_ (.A(\hvsync_gen.hpos[8] ),
    .X(_0131_));
 sg13g2_buf_1 _0900_ (.A(net62),
    .X(_0132_));
 sg13g2_a21oi_1 _0901_ (.A1(net51),
    .A2(net28),
    .Y(_0133_),
    .B1(net50));
 sg13g2_nor2_1 _0902_ (.A(_0124_),
    .B(_0133_),
    .Y(_0134_));
 sg13g2_buf_2 _0903_ (.A(\hvsync_gen.hpos[7] ),
    .X(_0135_));
 sg13g2_buf_1 _0904_ (.A(_0135_),
    .X(_0136_));
 sg13g2_or3_1 _0905_ (.A(net64),
    .B(net63),
    .C(net51),
    .X(_0137_));
 sg13g2_a21oi_1 _0906_ (.A1(net49),
    .A2(_0137_),
    .Y(_0138_),
    .B1(net50));
 sg13g2_nor3_1 _0907_ (.A(_0123_),
    .B(_0134_),
    .C(_0138_),
    .Y(_0015_));
 sg13g2_buf_1 _0908_ (.A(BNC_trig),
    .X(_0139_));
 sg13g2_buf_1 _0909_ (.A(net61),
    .X(_0140_));
 sg13g2_buf_1 _0910_ (.A(\bnc_image_generator.counter[0] ),
    .X(_0141_));
 sg13g2_buf_1 _0911_ (.A(net60),
    .X(_0142_));
 sg13g2_inv_1 _0912_ (.Y(_0143_),
    .A(\bnc_image_generator.counter[2] ));
 sg13g2_buf_2 _0913_ (.A(\bnc_image_generator.counter[4] ),
    .X(_0144_));
 sg13g2_buf_1 _0914_ (.A(_0144_),
    .X(_0145_));
 sg13g2_nand2_2 _0915_ (.Y(_0146_),
    .A(net59),
    .B(net46));
 sg13g2_buf_1 _0916_ (.A(\bnc_image_generator.counter[2] ),
    .X(_0147_));
 sg13g2_nand2b_1 _0917_ (.Y(_0148_),
    .B(net58),
    .A_N(_0144_));
 sg13g2_nand3_1 _0918_ (.B(_0146_),
    .C(_0148_),
    .A(net47),
    .Y(_0149_));
 sg13g2_o21ai_1 _0919_ (.B1(_0149_),
    .Y(_0150_),
    .A1(net47),
    .A2(_0146_));
 sg13g2_buf_1 _0920_ (.A(\bnc_image_generator.counter[1] ),
    .X(_0151_));
 sg13g2_buf_1 _0921_ (.A(net57),
    .X(_0152_));
 sg13g2_buf_1 _0922_ (.A(net61),
    .X(_0153_));
 sg13g2_nand2b_1 _0923_ (.Y(_0154_),
    .B(net58),
    .A_N(net60));
 sg13g2_nand2_1 _0924_ (.Y(_0155_),
    .A(net60),
    .B(net59));
 sg13g2_a22oi_1 _0925_ (.Y(_0156_),
    .B1(_0154_),
    .B2(_0155_),
    .A2(net46),
    .A1(net44));
 sg13g2_inv_2 _0926_ (.Y(_0157_),
    .A(net57));
 sg13g2_or2_1 _0927_ (.X(_0158_),
    .B(_0154_),
    .A(_0157_));
 sg13g2_inv_1 _0928_ (.Y(_0159_),
    .A(BNC_trig));
 sg13g2_buf_1 _0929_ (.A(_0159_),
    .X(_0160_));
 sg13g2_nand2b_1 _0930_ (.Y(_0161_),
    .B(net43),
    .A_N(_0158_));
 sg13g2_o21ai_1 _0931_ (.B1(_0161_),
    .Y(_0162_),
    .A1(net45),
    .A2(_0156_));
 sg13g2_a21oi_1 _0932_ (.A1(net48),
    .A2(_0150_),
    .Y(_0000_),
    .B1(_0162_));
 sg13g2_a21oi_1 _0933_ (.A1(_0146_),
    .A2(_0148_),
    .Y(_0163_),
    .B1(_0157_));
 sg13g2_nand2_1 _0934_ (.Y(_0164_),
    .A(net58),
    .B(_0144_));
 sg13g2_nor2_1 _0935_ (.A(net45),
    .B(_0164_),
    .Y(_0165_));
 sg13g2_nor2_1 _0936_ (.A(_0163_),
    .B(_0165_),
    .Y(_0166_));
 sg13g2_nor2_1 _0937_ (.A(net59),
    .B(_0144_),
    .Y(_0167_));
 sg13g2_a22oi_1 _0938_ (.Y(_0168_),
    .B1(_0167_),
    .B2(net45),
    .A2(_0145_),
    .A1(net61));
 sg13g2_nor2_1 _0939_ (.A(net47),
    .B(_0168_),
    .Y(_0169_));
 sg13g2_buf_1 _0940_ (.A(net58),
    .X(_0170_));
 sg13g2_nand2_2 _0941_ (.Y(_0171_),
    .A(_0157_),
    .B(net60));
 sg13g2_nor3_1 _0942_ (.A(net42),
    .B(net46),
    .C(_0171_),
    .Y(_0172_));
 sg13g2_nor2_1 _0943_ (.A(net57),
    .B(_0144_),
    .Y(_0173_));
 sg13g2_nand2_1 _0944_ (.Y(_0174_),
    .A(_0154_),
    .B(_0173_));
 sg13g2_a21oi_1 _0945_ (.A1(_0155_),
    .A2(_0174_),
    .Y(_0175_),
    .B1(net44));
 sg13g2_nor3_1 _0946_ (.A(_0169_),
    .B(_0172_),
    .C(_0175_),
    .Y(_0176_));
 sg13g2_o21ai_1 _0947_ (.B1(_0176_),
    .Y(_0001_),
    .A1(net43),
    .A2(_0166_));
 sg13g2_buf_1 _0948_ (.A(net46),
    .X(_0177_));
 sg13g2_and2_1 _0949_ (.A(net57),
    .B(net60),
    .X(_0178_));
 sg13g2_buf_1 _0950_ (.A(_0178_),
    .X(_0179_));
 sg13g2_xnor2_1 _0951_ (.Y(_0180_),
    .A(net42),
    .B(_0179_));
 sg13g2_nand2b_2 _0952_ (.Y(_0181_),
    .B(net57),
    .A_N(net60));
 sg13g2_a21oi_1 _0953_ (.A1(_0171_),
    .A2(_0181_),
    .Y(_0182_),
    .B1(_0018_));
 sg13g2_nor2_1 _0954_ (.A(net44),
    .B(_0182_),
    .Y(_0183_));
 sg13g2_a21oi_1 _0955_ (.A1(net48),
    .A2(_0180_),
    .Y(_0184_),
    .B1(_0183_));
 sg13g2_nand2_1 _0956_ (.Y(_0185_),
    .A(net58),
    .B(_0019_));
 sg13g2_nand2_1 _0957_ (.Y(_0186_),
    .A(net44),
    .B(_0185_));
 sg13g2_nand3_1 _0958_ (.B(_0158_),
    .C(_0171_),
    .A(net43),
    .Y(_0187_));
 sg13g2_buf_1 _0959_ (.A(net46),
    .X(_0188_));
 sg13g2_a221oi_1 _0960_ (.B2(_0187_),
    .C1(net26),
    .B1(_0186_),
    .A1(net59),
    .Y(_0189_),
    .A2(_0179_));
 sg13g2_a21oi_1 _0961_ (.A1(net27),
    .A2(_0184_),
    .Y(_0002_),
    .B1(_0189_));
 sg13g2_inv_1 _0962_ (.Y(_0190_),
    .A(_0030_));
 sg13g2_nand2_1 _0963_ (.Y(_0191_),
    .A(_0151_),
    .B(net47));
 sg13g2_nor2_1 _0964_ (.A(net58),
    .B(_0191_),
    .Y(_0192_));
 sg13g2_nor2_1 _0965_ (.A(net57),
    .B(net60),
    .Y(_0193_));
 sg13g2_nor2_1 _0966_ (.A(_0147_),
    .B(_0193_),
    .Y(_0194_));
 sg13g2_nor2_1 _0967_ (.A(net61),
    .B(_0194_),
    .Y(_0195_));
 sg13g2_a221oi_1 _0968_ (.B2(net44),
    .C1(_0195_),
    .B1(_0192_),
    .A1(net42),
    .Y(_0196_),
    .A2(_0190_));
 sg13g2_o21ai_1 _0969_ (.B1(_0142_),
    .Y(_0197_),
    .A1(_0152_),
    .A2(_0170_));
 sg13g2_nor2_1 _0970_ (.A(_0141_),
    .B(\bnc_image_generator.counter[2] ),
    .Y(_0198_));
 sg13g2_a221oi_1 _0971_ (.B2(_0152_),
    .C1(_0188_),
    .B1(_0198_),
    .A1(_0153_),
    .Y(_0199_),
    .A2(_0197_));
 sg13g2_a21o_1 _0972_ (.A2(_0196_),
    .A1(_0177_),
    .B1(_0199_),
    .X(_0003_));
 sg13g2_nor2_1 _0973_ (.A(net43),
    .B(net26),
    .Y(_0200_));
 sg13g2_nor3_1 _0974_ (.A(net44),
    .B(net47),
    .C(_0146_),
    .Y(_0201_));
 sg13g2_o21ai_1 _0975_ (.B1(net45),
    .Y(_0202_),
    .A1(_0200_),
    .A2(_0201_));
 sg13g2_nand3_1 _0976_ (.B(_0142_),
    .C(net59),
    .A(_0157_),
    .Y(_0203_));
 sg13g2_nand2_1 _0977_ (.Y(_0204_),
    .A(_0185_),
    .B(_0203_));
 sg13g2_nand3_1 _0978_ (.B(net26),
    .C(_0204_),
    .A(net48),
    .Y(_0205_));
 sg13g2_a21oi_1 _0979_ (.A1(net61),
    .A2(_0198_),
    .Y(_0206_),
    .B1(_0195_));
 sg13g2_or2_1 _0980_ (.X(_0207_),
    .B(_0206_),
    .A(net26));
 sg13g2_nand3_1 _0981_ (.B(_0205_),
    .C(_0207_),
    .A(_0202_),
    .Y(_0004_));
 sg13g2_inv_1 _0982_ (.Y(_0208_),
    .A(_0198_));
 sg13g2_nand2_1 _0983_ (.Y(_0209_),
    .A(net47),
    .B(_0147_));
 sg13g2_o21ai_1 _0984_ (.B1(_0209_),
    .Y(_0210_),
    .A1(_0157_),
    .A2(_0208_));
 sg13g2_nor2_1 _0985_ (.A(net61),
    .B(_0203_),
    .Y(_0211_));
 sg13g2_a21oi_1 _0986_ (.A1(_0140_),
    .A2(_0210_),
    .Y(_0212_),
    .B1(_0211_));
 sg13g2_xor2_1 _0987_ (.B(_0212_),
    .A(net27),
    .X(_0005_));
 sg13g2_nor2b_1 _0988_ (.A(net61),
    .B_N(_0144_),
    .Y(_0213_));
 sg13g2_a21o_1 _0989_ (.A2(_0179_),
    .A1(_0145_),
    .B1(_0173_),
    .X(_0214_));
 sg13g2_a22oi_1 _0990_ (.Y(_0215_),
    .B1(_0214_),
    .B2(net48),
    .A2(_0213_),
    .A1(_0193_));
 sg13g2_a22oi_1 _0991_ (.Y(_0216_),
    .B1(_0208_),
    .B2(_0159_),
    .A2(_0155_),
    .A1(net45));
 sg13g2_nand4_1 _0992_ (.B(net42),
    .C(net46),
    .A(net44),
    .Y(_0217_),
    .D(_0019_));
 sg13g2_o21ai_1 _0993_ (.B1(_0217_),
    .Y(_0218_),
    .A1(_0188_),
    .A2(_0216_));
 sg13g2_inv_1 _0994_ (.Y(_0219_),
    .A(_0218_));
 sg13g2_o21ai_1 _0995_ (.B1(_0219_),
    .Y(_0006_),
    .A1(net42),
    .A2(_0215_));
 sg13g2_nand3_1 _0996_ (.B(net45),
    .C(_0170_),
    .A(_0153_),
    .Y(_0220_));
 sg13g2_nand2_1 _0997_ (.Y(_0221_),
    .A(net57),
    .B(net58));
 sg13g2_o21ai_1 _0998_ (.B1(net26),
    .Y(_0222_),
    .A1(_0017_),
    .A2(_0221_));
 sg13g2_o21ai_1 _0999_ (.B1(_0222_),
    .Y(_0223_),
    .A1(net27),
    .A2(_0220_));
 sg13g2_inv_1 _1000_ (.Y(_0007_),
    .A(_0223_));
 sg13g2_nor2b_2 _1001_ (.A(_0141_),
    .B_N(_0144_),
    .Y(_0224_));
 sg13g2_nor2_1 _1002_ (.A(net42),
    .B(_0224_),
    .Y(_0225_));
 sg13g2_a22oi_1 _1003_ (.Y(_0226_),
    .B1(_0225_),
    .B2(net48),
    .A2(_0213_),
    .A1(_0208_));
 sg13g2_nand2b_1 _1004_ (.Y(_0227_),
    .B(net61),
    .A_N(net47));
 sg13g2_o21ai_1 _1005_ (.B1(_0146_),
    .Y(_0228_),
    .A1(_0148_),
    .A2(_0227_));
 sg13g2_o21ai_1 _1006_ (.B1(_0203_),
    .Y(_0229_),
    .A1(net46),
    .A2(_0185_));
 sg13g2_a22oi_1 _1007_ (.Y(_0230_),
    .B1(_0229_),
    .B2(net43),
    .A2(_0228_),
    .A1(_0157_));
 sg13g2_o21ai_1 _1008_ (.B1(_0230_),
    .Y(_0008_),
    .A1(_0157_),
    .A2(_0226_));
 sg13g2_xnor2_1 _1009_ (.Y(_0231_),
    .A(net58),
    .B(_0224_));
 sg13g2_nor2b_1 _1010_ (.A(_0144_),
    .B_N(net60),
    .Y(_0232_));
 sg13g2_nor3_1 _1011_ (.A(net57),
    .B(_0224_),
    .C(_0232_),
    .Y(_0233_));
 sg13g2_a21oi_1 _1012_ (.A1(net45),
    .A2(_0231_),
    .Y(_0234_),
    .B1(_0233_));
 sg13g2_a21oi_1 _1013_ (.A1(_0018_),
    .A2(_0224_),
    .Y(_0235_),
    .B1(_0167_));
 sg13g2_mux2_1 _1014_ (.A0(_0234_),
    .A1(_0235_),
    .S(net43),
    .X(_0236_));
 sg13g2_o21ai_1 _1015_ (.B1(_0236_),
    .Y(_0009_),
    .A1(net27),
    .A2(_0191_));
 sg13g2_o21ai_1 _1016_ (.B1(_0148_),
    .Y(_0237_),
    .A1(_0146_),
    .A2(_0181_));
 sg13g2_a21oi_1 _1017_ (.A1(_0179_),
    .A2(_0213_),
    .Y(_0238_),
    .B1(_0173_));
 sg13g2_nor2_1 _1018_ (.A(_0030_),
    .B(_0164_),
    .Y(_0239_));
 sg13g2_nor2_1 _1019_ (.A(net47),
    .B(net46),
    .Y(_0240_));
 sg13g2_o21ai_1 _1020_ (.B1(net43),
    .Y(_0241_),
    .A1(_0239_),
    .A2(_0240_));
 sg13g2_o21ai_1 _1021_ (.B1(_0241_),
    .Y(_0242_),
    .A1(net42),
    .A2(_0238_));
 sg13g2_a21oi_1 _1022_ (.A1(net48),
    .A2(_0237_),
    .Y(_0010_),
    .B1(_0242_));
 sg13g2_o21ai_1 _1023_ (.B1(_0185_),
    .Y(_0243_),
    .A1(net43),
    .A2(_0194_));
 sg13g2_nor2_1 _1024_ (.A(_0211_),
    .B(_0243_),
    .Y(_0244_));
 sg13g2_o21ai_1 _1025_ (.B1(_0181_),
    .Y(_0245_),
    .A1(_0159_),
    .A2(_0171_));
 sg13g2_nand2_1 _1026_ (.Y(_0246_),
    .A(_0157_),
    .B(_0208_));
 sg13g2_a221oi_1 _1027_ (.B2(_0160_),
    .C1(net26),
    .B1(_0246_),
    .A1(net59),
    .Y(_0247_),
    .A2(_0245_));
 sg13g2_a21oi_1 _1028_ (.A1(net27),
    .A2(_0244_),
    .Y(_0011_),
    .B1(_0247_));
 sg13g2_a21oi_1 _1029_ (.A1(net48),
    .A2(_0171_),
    .Y(_0248_),
    .B1(_0210_));
 sg13g2_nor2_1 _1030_ (.A(_0139_),
    .B(net59),
    .Y(_0249_));
 sg13g2_nand2_1 _1031_ (.Y(_0250_),
    .A(_0159_),
    .B(_0181_));
 sg13g2_nand2_1 _1032_ (.Y(_0251_),
    .A(_0171_),
    .B(_0250_));
 sg13g2_a221oi_1 _1033_ (.B2(net59),
    .C1(net26),
    .B1(_0251_),
    .A1(_0030_),
    .Y(_0252_),
    .A2(_0249_));
 sg13g2_a21oi_1 _1034_ (.A1(net27),
    .A2(_0248_),
    .Y(_0012_),
    .B1(_0252_));
 sg13g2_nor2_1 _1035_ (.A(_0159_),
    .B(_0193_),
    .Y(_0253_));
 sg13g2_nor2_1 _1036_ (.A(_0192_),
    .B(_0253_),
    .Y(_0254_));
 sg13g2_o21ai_1 _1037_ (.B1(_0254_),
    .Y(_0255_),
    .A1(net45),
    .A2(_0143_));
 sg13g2_nand2b_1 _1038_ (.Y(_0256_),
    .B(_0249_),
    .A_N(_0019_));
 sg13g2_nor2_1 _1039_ (.A(_0139_),
    .B(_0179_),
    .Y(_0257_));
 sg13g2_o21ai_1 _1040_ (.B1(_0143_),
    .Y(_0258_),
    .A1(_0193_),
    .A2(_0257_));
 sg13g2_nand3_1 _1041_ (.B(_0256_),
    .C(_0258_),
    .A(net27),
    .Y(_0259_));
 sg13g2_o21ai_1 _1042_ (.B1(_0259_),
    .Y(_0013_),
    .A1(_0177_),
    .A2(_0255_));
 sg13g2_a21oi_1 _1043_ (.A1(_0017_),
    .A2(_0221_),
    .Y(_0260_),
    .B1(net27));
 sg13g2_a21oi_1 _1044_ (.A1(_0213_),
    .A2(_0221_),
    .Y(_0014_),
    .B1(_0260_));
 sg13g2_buf_1 _1045_ (.A(rst_n),
    .X(_0261_));
 sg13g2_buf_2 _1046_ (.A(\hvsync_gen.hpos[2] ),
    .X(_0262_));
 sg13g2_buf_8 _1047_ (.A(\hvsync_gen.hpos[3] ),
    .X(_0263_));
 sg13g2_nand2_1 _1048_ (.Y(_0264_),
    .A(_0262_),
    .B(_0263_));
 sg13g2_buf_1 _1049_ (.A(\hvsync_gen.hpos[1] ),
    .X(_0265_));
 sg13g2_buf_2 _1050_ (.A(\hvsync_gen.hpos[0] ),
    .X(_0266_));
 sg13g2_nand2_2 _1051_ (.Y(_0267_),
    .A(net55),
    .B(_0266_));
 sg13g2_nor2_2 _1052_ (.A(_0264_),
    .B(_0267_),
    .Y(_0268_));
 sg13g2_or2_1 _1053_ (.X(_0269_),
    .B(_0135_),
    .A(_0125_));
 sg13g2_buf_2 _1054_ (.A(_0269_),
    .X(_0270_));
 sg13g2_nand2b_1 _1055_ (.Y(_0271_),
    .B(net63),
    .A_N(net64));
 sg13g2_nor2_1 _1056_ (.A(_0270_),
    .B(_0271_),
    .Y(_0272_));
 sg13g2_nand3_1 _1057_ (.B(_0268_),
    .C(_0272_),
    .A(net62),
    .Y(_0273_));
 sg13g2_or2_1 _1058_ (.X(_0274_),
    .B(_0273_),
    .A(_0123_));
 sg13g2_and2_1 _1059_ (.A(_0261_),
    .B(_0274_),
    .X(_0275_));
 sg13g2_buf_1 _1060_ (.A(_0275_),
    .X(_0276_));
 sg13g2_buf_1 _1061_ (.A(\hvsync_gen.vpos[5] ),
    .X(_0277_));
 sg13g2_buf_1 _1062_ (.A(\hvsync_gen.vpos[4] ),
    .X(_0278_));
 sg13g2_inv_1 _1063_ (.Y(_0279_),
    .A(\hvsync_gen.vpos[9] ));
 sg13g2_nor4_1 _1064_ (.A(net54),
    .B(net53),
    .C(net67),
    .D(_0279_),
    .Y(_0280_));
 sg13g2_or2_1 _1065_ (.X(_0281_),
    .B(\hvsync_gen.vpos[0] ),
    .A(\hvsync_gen.vpos[1] ));
 sg13g2_buf_1 _1066_ (.A(_0281_),
    .X(_0282_));
 sg13g2_nand2_1 _1067_ (.Y(_0283_),
    .A(net68),
    .B(_0109_));
 sg13g2_nor4_1 _1068_ (.A(net66),
    .B(net65),
    .C(_0282_),
    .D(_0283_),
    .Y(_0284_));
 sg13g2_inv_1 _1069_ (.Y(_0285_),
    .A(_0261_));
 sg13g2_a21o_1 _1070_ (.A2(_0284_),
    .A1(_0280_),
    .B1(_0285_),
    .X(_0286_));
 sg13g2_buf_1 _1071_ (.A(_0286_),
    .X(_0287_));
 sg13g2_or2_1 _1072_ (.X(_0288_),
    .B(net21),
    .A(_0274_));
 sg13g2_buf_2 _1073_ (.A(_0288_),
    .X(_0289_));
 sg13g2_inv_1 _1074_ (.Y(_0290_),
    .A(_0289_));
 sg13g2_a22oi_1 _1075_ (.Y(_0291_),
    .B1(_0290_),
    .B2(_0029_),
    .A2(net19),
    .A1(\hvsync_gen.vpos[0] ));
 sg13g2_inv_1 _1076_ (.Y(_0047_),
    .A(_0291_));
 sg13g2_nand2_1 _1077_ (.Y(_0292_),
    .A(_0107_),
    .B(\hvsync_gen.vpos[0] ));
 sg13g2_nand2_2 _1078_ (.Y(_0293_),
    .A(_0261_),
    .B(_0274_));
 sg13g2_o21ai_1 _1079_ (.B1(_0293_),
    .Y(_0294_),
    .A1(\hvsync_gen.vpos[0] ),
    .A2(_0289_));
 sg13g2_nand2_1 _1080_ (.Y(_0295_),
    .A(\hvsync_gen.vpos[1] ),
    .B(_0294_));
 sg13g2_o21ai_1 _1081_ (.B1(_0295_),
    .Y(_0048_),
    .A1(_0289_),
    .A2(_0292_));
 sg13g2_buf_1 _1082_ (.A(net68),
    .X(_0296_));
 sg13g2_and2_1 _1083_ (.A(\hvsync_gen.vpos[1] ),
    .B(\hvsync_gen.vpos[0] ),
    .X(_0297_));
 sg13g2_buf_2 _1084_ (.A(_0297_),
    .X(_0298_));
 sg13g2_nor2_1 _1085_ (.A(net19),
    .B(net21),
    .Y(_0299_));
 sg13g2_nand2_1 _1086_ (.Y(_0300_),
    .A(_0298_),
    .B(_0299_));
 sg13g2_nor2_1 _1087_ (.A(net21),
    .B(_0298_),
    .Y(_0301_));
 sg13g2_o21ai_1 _1088_ (.B1(net41),
    .Y(_0302_),
    .A1(net19),
    .A2(_0301_));
 sg13g2_o21ai_1 _1089_ (.B1(_0302_),
    .Y(_0049_),
    .A1(net41),
    .A2(_0300_));
 sg13g2_nand3_1 _1090_ (.B(_0110_),
    .C(_0298_),
    .A(net41),
    .Y(_0303_));
 sg13g2_a21oi_1 _1091_ (.A1(net41),
    .A2(_0298_),
    .Y(_0304_),
    .B1(net21));
 sg13g2_buf_1 _1092_ (.A(_0109_),
    .X(_0305_));
 sg13g2_o21ai_1 _1093_ (.B1(net40),
    .Y(_0306_),
    .A1(net19),
    .A2(_0304_));
 sg13g2_o21ai_1 _1094_ (.B1(_0306_),
    .Y(_0050_),
    .A1(_0289_),
    .A2(_0303_));
 sg13g2_inv_1 _1095_ (.Y(_0307_),
    .A(net53));
 sg13g2_nor2b_2 _1096_ (.A(_0283_),
    .B_N(_0298_),
    .Y(_0308_));
 sg13g2_nand2_1 _1097_ (.Y(_0309_),
    .A(_0307_),
    .B(_0308_));
 sg13g2_nor2_1 _1098_ (.A(net21),
    .B(_0308_),
    .Y(_0310_));
 sg13g2_buf_1 _1099_ (.A(net53),
    .X(_0311_));
 sg13g2_o21ai_1 _1100_ (.B1(net39),
    .Y(_0312_),
    .A1(net19),
    .A2(_0310_));
 sg13g2_o21ai_1 _1101_ (.B1(_0312_),
    .Y(_0051_),
    .A1(_0289_),
    .A2(_0309_));
 sg13g2_inv_2 _1102_ (.Y(_0313_),
    .A(net54));
 sg13g2_nand3_1 _1103_ (.B(net39),
    .C(_0308_),
    .A(_0313_),
    .Y(_0314_));
 sg13g2_a21oi_1 _1104_ (.A1(net39),
    .A2(_0308_),
    .Y(_0315_),
    .B1(net21));
 sg13g2_o21ai_1 _1105_ (.B1(_0277_),
    .Y(_0316_),
    .A1(net19),
    .A2(_0315_));
 sg13g2_o21ai_1 _1106_ (.B1(_0316_),
    .Y(_0052_),
    .A1(_0289_),
    .A2(_0314_));
 sg13g2_and3_1 _1107_ (.X(_0317_),
    .A(_0277_),
    .B(_0311_),
    .C(_0308_));
 sg13g2_buf_1 _1108_ (.A(_0317_),
    .X(_0318_));
 sg13g2_nand2_1 _1109_ (.Y(_0319_),
    .A(_0299_),
    .B(_0318_));
 sg13g2_nor2_1 _1110_ (.A(net21),
    .B(_0318_),
    .Y(_0320_));
 sg13g2_o21ai_1 _1111_ (.B1(net65),
    .Y(_0321_),
    .A1(net19),
    .A2(_0320_));
 sg13g2_o21ai_1 _1112_ (.B1(_0321_),
    .Y(_0053_),
    .A1(net65),
    .A2(_0319_));
 sg13g2_nand3_1 _1113_ (.B(_0299_),
    .C(_0318_),
    .A(_0120_),
    .Y(_0322_));
 sg13g2_a21oi_1 _1114_ (.A1(_0120_),
    .A2(_0318_),
    .Y(_0323_),
    .B1(net21));
 sg13g2_o21ai_1 _1115_ (.B1(net66),
    .Y(_0324_),
    .A1(_0276_),
    .A2(_0323_));
 sg13g2_o21ai_1 _1116_ (.B1(_0324_),
    .Y(_0054_),
    .A1(net66),
    .A2(_0322_));
 sg13g2_nor2b_1 _1117_ (.A(_0121_),
    .B_N(_0318_),
    .Y(_0325_));
 sg13g2_nand2_1 _1118_ (.Y(_0326_),
    .A(_0299_),
    .B(_0325_));
 sg13g2_o21ai_1 _1119_ (.B1(_0293_),
    .Y(_0327_),
    .A1(_0287_),
    .A2(_0325_));
 sg13g2_nand2_1 _1120_ (.Y(_0328_),
    .A(net67),
    .B(_0327_));
 sg13g2_o21ai_1 _1121_ (.B1(_0328_),
    .Y(_0055_),
    .A1(net67),
    .A2(_0326_));
 sg13g2_nand2_1 _1122_ (.Y(_0329_),
    .A(_0114_),
    .B(_0325_));
 sg13g2_a21oi_1 _1123_ (.A1(net67),
    .A2(_0325_),
    .Y(_0330_),
    .B1(_0289_));
 sg13g2_o21ai_1 _1124_ (.B1(\hvsync_gen.vpos[9] ),
    .Y(_0331_),
    .A1(net19),
    .A2(_0330_));
 sg13g2_o21ai_1 _1125_ (.B1(_0331_),
    .Y(_0056_),
    .A1(_0289_),
    .A2(_0329_));
 sg13g2_and2_1 _1126_ (.A(_0028_),
    .B(_0276_),
    .X(_0037_));
 sg13g2_buf_1 _1127_ (.A(_0285_),
    .X(_0332_));
 sg13g2_buf_1 _1128_ (.A(_0332_),
    .X(_0333_));
 sg13g2_xnor2_1 _1129_ (.Y(_0334_),
    .A(net55),
    .B(_0266_));
 sg13g2_nor2_1 _1130_ (.A(net25),
    .B(_0334_),
    .Y(_0038_));
 sg13g2_buf_1 _1131_ (.A(_0262_),
    .X(_0335_));
 sg13g2_and2_1 _1132_ (.A(net55),
    .B(_0266_),
    .X(_0336_));
 sg13g2_buf_1 _1133_ (.A(_0336_),
    .X(_0337_));
 sg13g2_xnor2_1 _1134_ (.Y(_0338_),
    .A(net37),
    .B(_0337_));
 sg13g2_nor2_1 _1135_ (.A(net25),
    .B(_0338_),
    .Y(_0039_));
 sg13g2_inv_2 _1136_ (.Y(_0339_),
    .A(net56));
 sg13g2_nand2_1 _1137_ (.Y(_0340_),
    .A(net37),
    .B(_0337_));
 sg13g2_xnor2_1 _1138_ (.Y(_0341_),
    .A(_0339_),
    .B(_0340_));
 sg13g2_nor2_1 _1139_ (.A(net25),
    .B(_0341_),
    .Y(_0040_));
 sg13g2_buf_1 _1140_ (.A(net63),
    .X(_0342_));
 sg13g2_xnor2_1 _1141_ (.Y(_0343_),
    .A(net36),
    .B(_0268_));
 sg13g2_nor2_1 _1142_ (.A(_0293_),
    .B(_0343_),
    .Y(_0041_));
 sg13g2_inv_1 _1143_ (.Y(_0344_),
    .A(_0127_));
 sg13g2_nand2_1 _1144_ (.Y(_0345_),
    .A(_0342_),
    .B(_0268_));
 sg13g2_xnor2_1 _1145_ (.Y(_0346_),
    .A(_0344_),
    .B(_0345_));
 sg13g2_nor2_1 _1146_ (.A(_0293_),
    .B(_0346_),
    .Y(_0042_));
 sg13g2_inv_1 _1147_ (.Y(_0347_),
    .A(net51));
 sg13g2_buf_1 _1148_ (.A(net64),
    .X(_0348_));
 sg13g2_nand3_1 _1149_ (.B(_0342_),
    .C(_0268_),
    .A(net35),
    .Y(_0349_));
 sg13g2_xnor2_1 _1150_ (.Y(_0350_),
    .A(_0347_),
    .B(_0349_));
 sg13g2_nor2_1 _1151_ (.A(_0293_),
    .B(_0350_),
    .Y(_0043_));
 sg13g2_nor3_2 _1152_ (.A(_0344_),
    .B(_0347_),
    .C(_0345_),
    .Y(_0351_));
 sg13g2_xnor2_1 _1153_ (.Y(_0352_),
    .A(net49),
    .B(_0351_));
 sg13g2_nor2_1 _1154_ (.A(_0293_),
    .B(_0352_),
    .Y(_0044_));
 sg13g2_nand2_1 _1155_ (.Y(_0353_),
    .A(net49),
    .B(_0351_));
 sg13g2_xor2_1 _1156_ (.B(_0353_),
    .A(net50),
    .X(_0354_));
 sg13g2_nor2_1 _1157_ (.A(_0293_),
    .B(_0354_),
    .Y(_0045_));
 sg13g2_nand3_1 _1158_ (.B(net50),
    .C(_0351_),
    .A(net49),
    .Y(_0355_));
 sg13g2_xnor2_1 _1159_ (.Y(_0356_),
    .A(_0123_),
    .B(_0355_));
 sg13g2_nor2_1 _1160_ (.A(_0293_),
    .B(_0356_),
    .Y(_0046_));
 sg13g2_nor2_1 _1161_ (.A(net25),
    .B(_0190_),
    .Y(_0032_));
 sg13g2_a21oi_1 _1162_ (.A1(_0171_),
    .A2(_0181_),
    .Y(_0033_),
    .B1(_0332_));
 sg13g2_nor2_1 _1163_ (.A(net25),
    .B(_0180_),
    .Y(_0034_));
 sg13g2_nor2_1 _1164_ (.A(_0030_),
    .B(_0221_),
    .Y(_0357_));
 sg13g2_xnor2_1 _1165_ (.Y(_0358_),
    .A(net48),
    .B(_0357_));
 sg13g2_nor2_1 _1166_ (.A(net25),
    .B(_0358_),
    .Y(_0035_));
 sg13g2_nand3_1 _1167_ (.B(net42),
    .C(_0179_),
    .A(net44),
    .Y(_0359_));
 sg13g2_xor2_1 _1168_ (.B(_0359_),
    .A(net26),
    .X(_0360_));
 sg13g2_nor2_1 _1169_ (.A(net25),
    .B(_0360_),
    .Y(_0036_));
 sg13g2_buf_2 _1170_ (.A(\vga_image_generator.counter[22] ),
    .X(_0361_));
 sg13g2_buf_1 _1171_ (.A(\vga_image_generator.counter[23] ),
    .X(_0362_));
 sg13g2_nor2_1 _1172_ (.A(_0361_),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_buf_2 _1173_ (.A(\vga_image_generator.counter[20] ),
    .X(_0364_));
 sg13g2_buf_2 _1174_ (.A(\vga_image_generator.counter[24] ),
    .X(_0365_));
 sg13g2_nor3_2 _1175_ (.A(\vga_image_generator.counter[21] ),
    .B(_0364_),
    .C(_0365_),
    .Y(_0366_));
 sg13g2_a21oi_1 _1176_ (.A1(_0363_),
    .A2(_0366_),
    .Y(_0367_),
    .B1(\vga_image_generator.character_hold[0] ));
 sg13g2_nor2_1 _1177_ (.A(net25),
    .B(_0367_),
    .Y(_0057_));
 sg13g2_nor2b_1 _1178_ (.A(_0361_),
    .B_N(_0362_),
    .Y(_0368_));
 sg13g2_nor2b_1 _1179_ (.A(_0365_),
    .B_N(_0368_),
    .Y(_0369_));
 sg13g2_nor2b_1 _1180_ (.A(_0364_),
    .B_N(\vga_image_generator.counter[21] ),
    .Y(_0370_));
 sg13g2_a21oi_1 _1181_ (.A1(_0369_),
    .A2(_0370_),
    .Y(_0371_),
    .B1(\vga_image_generator.character_hold[10] ));
 sg13g2_nor2_1 _1182_ (.A(_0333_),
    .B(_0371_),
    .Y(_0058_));
 sg13g2_and2_1 _1183_ (.A(\vga_image_generator.counter[21] ),
    .B(_0364_),
    .X(_0372_));
 sg13g2_a21oi_1 _1184_ (.A1(_0369_),
    .A2(_0372_),
    .Y(_0373_),
    .B1(\vga_image_generator.character_hold[11] ));
 sg13g2_nor2_1 _1185_ (.A(_0333_),
    .B(_0373_),
    .Y(_0059_));
 sg13g2_buf_1 _1186_ (.A(_0285_),
    .X(_0374_));
 sg13g2_and2_1 _1187_ (.A(_0361_),
    .B(_0362_),
    .X(_0375_));
 sg13g2_buf_1 _1188_ (.A(_0375_),
    .X(_0376_));
 sg13g2_a21oi_1 _1189_ (.A1(_0366_),
    .A2(_0376_),
    .Y(_0377_),
    .B1(\vga_image_generator.character_hold[12] ));
 sg13g2_nor2_1 _1190_ (.A(net34),
    .B(_0377_),
    .Y(_0060_));
 sg13g2_nor2b_1 _1191_ (.A(\vga_image_generator.counter[21] ),
    .B_N(_0364_),
    .Y(_0378_));
 sg13g2_nor2b_1 _1192_ (.A(_0365_),
    .B_N(_0378_),
    .Y(_0379_));
 sg13g2_a21oi_1 _1193_ (.A1(_0376_),
    .A2(_0379_),
    .Y(_0380_),
    .B1(\vga_image_generator.character_hold[13] ));
 sg13g2_nor2_1 _1194_ (.A(_0374_),
    .B(_0380_),
    .Y(_0061_));
 sg13g2_nor2b_1 _1195_ (.A(_0365_),
    .B_N(_0370_),
    .Y(_0381_));
 sg13g2_a21oi_1 _1196_ (.A1(_0376_),
    .A2(_0381_),
    .Y(_0382_),
    .B1(\vga_image_generator.character_hold[14] ));
 sg13g2_nor2_1 _1197_ (.A(_0374_),
    .B(_0382_),
    .Y(_0062_));
 sg13g2_nor2b_1 _1198_ (.A(_0365_),
    .B_N(_0372_),
    .Y(_0383_));
 sg13g2_a21oi_1 _1199_ (.A1(_0376_),
    .A2(_0383_),
    .Y(_0384_),
    .B1(\vga_image_generator.character_hold[15] ));
 sg13g2_nor2_1 _1200_ (.A(net34),
    .B(_0384_),
    .Y(_0063_));
 sg13g2_nor3_1 _1201_ (.A(_0361_),
    .B(_0362_),
    .C(_0020_),
    .Y(_0385_));
 sg13g2_a21oi_1 _1202_ (.A1(_0378_),
    .A2(_0385_),
    .Y(_0386_),
    .B1(\vga_image_generator.character_hold[16] ));
 sg13g2_nor2_1 _1203_ (.A(net34),
    .B(_0386_),
    .Y(_0064_));
 sg13g2_a21oi_1 _1204_ (.A1(_0370_),
    .A2(_0385_),
    .Y(_0387_),
    .B1(\vga_image_generator.character_hold[17] ));
 sg13g2_nor2_1 _1205_ (.A(net34),
    .B(_0387_),
    .Y(_0065_));
 sg13g2_a21oi_1 _1206_ (.A1(_0363_),
    .A2(_0379_),
    .Y(_0388_),
    .B1(\vga_image_generator.character_hold[1] ));
 sg13g2_nor2_1 _1207_ (.A(net34),
    .B(_0388_),
    .Y(_0066_));
 sg13g2_a21oi_1 _1208_ (.A1(_0363_),
    .A2(_0381_),
    .Y(_0389_),
    .B1(\vga_image_generator.character_hold[2] ));
 sg13g2_nor2_1 _1209_ (.A(net34),
    .B(_0389_),
    .Y(_0067_));
 sg13g2_a21oi_1 _1210_ (.A1(_0363_),
    .A2(_0383_),
    .Y(_0390_),
    .B1(\vga_image_generator.character_hold[3] ));
 sg13g2_nor2_1 _1211_ (.A(net34),
    .B(_0390_),
    .Y(_0068_));
 sg13g2_nor2b_1 _1212_ (.A(_0362_),
    .B_N(_0361_),
    .Y(_0391_));
 sg13g2_a21oi_1 _1213_ (.A1(_0366_),
    .A2(_0391_),
    .Y(_0392_),
    .B1(\vga_image_generator.character_hold[4] ));
 sg13g2_nor2_1 _1214_ (.A(net34),
    .B(_0392_),
    .Y(_0069_));
 sg13g2_buf_1 _1215_ (.A(_0285_),
    .X(_0393_));
 sg13g2_a21oi_1 _1216_ (.A1(_0379_),
    .A2(_0391_),
    .Y(_0394_),
    .B1(\vga_image_generator.character_hold[5] ));
 sg13g2_nor2_1 _1217_ (.A(net33),
    .B(_0394_),
    .Y(_0070_));
 sg13g2_a21oi_1 _1218_ (.A1(_0381_),
    .A2(_0391_),
    .Y(_0395_),
    .B1(\vga_image_generator.character_hold[6] ));
 sg13g2_nor2_1 _1219_ (.A(net33),
    .B(_0395_),
    .Y(_0071_));
 sg13g2_a21oi_1 _1220_ (.A1(_0383_),
    .A2(_0391_),
    .Y(_0396_),
    .B1(\vga_image_generator.character_hold[7] ));
 sg13g2_nor2_1 _1221_ (.A(net33),
    .B(_0396_),
    .Y(_0072_));
 sg13g2_a21oi_1 _1222_ (.A1(_0366_),
    .A2(_0368_),
    .Y(_0397_),
    .B1(\vga_image_generator.character_hold[8] ));
 sg13g2_nor2_1 _1223_ (.A(_0393_),
    .B(_0397_),
    .Y(_0073_));
 sg13g2_a21oi_1 _1224_ (.A1(_0369_),
    .A2(_0378_),
    .Y(_0398_),
    .B1(\vga_image_generator.character_hold[9] ));
 sg13g2_nor2_1 _1225_ (.A(_0393_),
    .B(_0398_),
    .Y(_0074_));
 sg13g2_and2_1 _1226_ (.A(_0261_),
    .B(_0031_),
    .X(_0075_));
 sg13g2_inv_1 _1227_ (.Y(_0399_),
    .A(\vga_image_generator.counter[8] ));
 sg13g2_and4_1 _1228_ (.A(\vga_image_generator.counter[1] ),
    .B(\vga_image_generator.counter[0] ),
    .C(\vga_image_generator.counter[2] ),
    .D(\vga_image_generator.counter[3] ),
    .X(_0400_));
 sg13g2_buf_8 _1229_ (.A(_0400_),
    .X(_0401_));
 sg13g2_and2_1 _1230_ (.A(\vga_image_generator.counter[6] ),
    .B(\vga_image_generator.counter[7] ),
    .X(_0402_));
 sg13g2_nand4_1 _1231_ (.B(\vga_image_generator.counter[5] ),
    .C(_0401_),
    .A(\vga_image_generator.counter[4] ),
    .Y(_0403_),
    .D(_0402_));
 sg13g2_buf_2 _1232_ (.A(_0403_),
    .X(_0404_));
 sg13g2_nor2_1 _1233_ (.A(_0399_),
    .B(_0404_),
    .Y(_0405_));
 sg13g2_nand2_1 _1234_ (.Y(_0406_),
    .A(\vga_image_generator.counter[9] ),
    .B(_0405_));
 sg13g2_xor2_1 _1235_ (.B(_0406_),
    .A(\vga_image_generator.counter[10] ),
    .X(_0407_));
 sg13g2_nor2_1 _1236_ (.A(net33),
    .B(_0407_),
    .Y(_0076_));
 sg13g2_nand2_1 _1237_ (.Y(_0408_),
    .A(\vga_image_generator.counter[9] ),
    .B(\vga_image_generator.counter[10] ));
 sg13g2_nor3_1 _1238_ (.A(_0399_),
    .B(_0404_),
    .C(_0408_),
    .Y(_0409_));
 sg13g2_xnor2_1 _1239_ (.Y(_0410_),
    .A(\vga_image_generator.counter[11] ),
    .B(_0409_));
 sg13g2_nor2_1 _1240_ (.A(net33),
    .B(_0410_),
    .Y(_0077_));
 sg13g2_inv_1 _1241_ (.Y(_0411_),
    .A(\vga_image_generator.counter[12] ));
 sg13g2_nand4_1 _1242_ (.B(\vga_image_generator.counter[10] ),
    .C(\vga_image_generator.counter[11] ),
    .A(\vga_image_generator.counter[9] ),
    .Y(_0412_),
    .D(_0405_));
 sg13g2_xnor2_1 _1243_ (.Y(_0413_),
    .A(_0411_),
    .B(_0412_));
 sg13g2_nor2_1 _1244_ (.A(net33),
    .B(_0413_),
    .Y(_0078_));
 sg13g2_nand4_1 _1245_ (.B(\vga_image_generator.counter[9] ),
    .C(\vga_image_generator.counter[10] ),
    .A(\vga_image_generator.counter[8] ),
    .Y(_0414_),
    .D(\vga_image_generator.counter[11] ));
 sg13g2_nor3_1 _1246_ (.A(_0411_),
    .B(_0404_),
    .C(_0414_),
    .Y(_0415_));
 sg13g2_xnor2_1 _1247_ (.Y(_0416_),
    .A(\vga_image_generator.counter[13] ),
    .B(_0415_));
 sg13g2_nor2_1 _1248_ (.A(net33),
    .B(_0416_),
    .Y(_0079_));
 sg13g2_nand2_1 _1249_ (.Y(_0417_),
    .A(\vga_image_generator.counter[13] ),
    .B(_0415_));
 sg13g2_xor2_1 _1250_ (.B(_0417_),
    .A(\vga_image_generator.counter[14] ),
    .X(_0418_));
 sg13g2_nor2_1 _1251_ (.A(net33),
    .B(_0418_),
    .Y(_0080_));
 sg13g2_buf_1 _1252_ (.A(_0285_),
    .X(_0419_));
 sg13g2_nand2_1 _1253_ (.Y(_0420_),
    .A(\vga_image_generator.counter[13] ),
    .B(\vga_image_generator.counter[14] ));
 sg13g2_nor4_2 _1254_ (.A(_0411_),
    .B(_0404_),
    .C(_0414_),
    .Y(_0421_),
    .D(_0420_));
 sg13g2_xnor2_1 _1255_ (.Y(_0422_),
    .A(\vga_image_generator.counter[15] ),
    .B(_0421_));
 sg13g2_nor2_1 _1256_ (.A(net32),
    .B(_0422_),
    .Y(_0081_));
 sg13g2_inv_1 _1257_ (.Y(_0423_),
    .A(\vga_image_generator.counter[16] ));
 sg13g2_nand2_1 _1258_ (.Y(_0424_),
    .A(\vga_image_generator.counter[11] ),
    .B(\vga_image_generator.counter[12] ));
 sg13g2_nor4_1 _1259_ (.A(_0399_),
    .B(_0404_),
    .C(_0408_),
    .D(_0424_),
    .Y(_0425_));
 sg13g2_nand4_1 _1260_ (.B(\vga_image_generator.counter[14] ),
    .C(\vga_image_generator.counter[15] ),
    .A(\vga_image_generator.counter[13] ),
    .Y(_0426_),
    .D(_0425_));
 sg13g2_xnor2_1 _1261_ (.Y(_0427_),
    .A(_0423_),
    .B(_0426_));
 sg13g2_nor2_1 _1262_ (.A(net32),
    .B(_0427_),
    .Y(_0082_));
 sg13g2_nor2_1 _1263_ (.A(_0423_),
    .B(_0426_),
    .Y(_0428_));
 sg13g2_xnor2_1 _1264_ (.Y(_0429_),
    .A(\vga_image_generator.counter[17] ),
    .B(_0428_));
 sg13g2_nor2_1 _1265_ (.A(net32),
    .B(_0429_),
    .Y(_0083_));
 sg13g2_nand2_1 _1266_ (.Y(_0430_),
    .A(\vga_image_generator.counter[17] ),
    .B(_0428_));
 sg13g2_xor2_1 _1267_ (.B(_0430_),
    .A(\vga_image_generator.counter[18] ),
    .X(_0431_));
 sg13g2_nor2_1 _1268_ (.A(net32),
    .B(_0431_),
    .Y(_0084_));
 sg13g2_inv_1 _1269_ (.Y(_0432_),
    .A(\vga_image_generator.counter[19] ));
 sg13g2_nand3_1 _1270_ (.B(\vga_image_generator.counter[18] ),
    .C(_0428_),
    .A(\vga_image_generator.counter[17] ),
    .Y(_0433_));
 sg13g2_xnor2_1 _1271_ (.Y(_0434_),
    .A(_0432_),
    .B(_0433_));
 sg13g2_nor2_1 _1272_ (.A(net32),
    .B(_0434_),
    .Y(_0085_));
 sg13g2_xnor2_1 _1273_ (.Y(_0435_),
    .A(\vga_image_generator.counter[1] ),
    .B(\vga_image_generator.counter[0] ));
 sg13g2_nor2_1 _1274_ (.A(net32),
    .B(_0435_),
    .Y(_0086_));
 sg13g2_nand4_1 _1275_ (.B(\vga_image_generator.counter[16] ),
    .C(\vga_image_generator.counter[17] ),
    .A(\vga_image_generator.counter[15] ),
    .Y(_0436_),
    .D(\vga_image_generator.counter[18] ));
 sg13g2_nor2_1 _1276_ (.A(_0432_),
    .B(_0436_),
    .Y(_0437_));
 sg13g2_nand2_1 _1277_ (.Y(_0438_),
    .A(_0421_),
    .B(_0437_));
 sg13g2_xor2_1 _1278_ (.B(_0438_),
    .A(_0364_),
    .X(_0439_));
 sg13g2_nor2_1 _1279_ (.A(_0419_),
    .B(_0439_),
    .Y(_0087_));
 sg13g2_nand3_1 _1280_ (.B(_0421_),
    .C(_0437_),
    .A(_0364_),
    .Y(_0440_));
 sg13g2_xor2_1 _1281_ (.B(_0440_),
    .A(\vga_image_generator.counter[21] ),
    .X(_0441_));
 sg13g2_nor2_1 _1282_ (.A(net32),
    .B(_0441_),
    .Y(_0088_));
 sg13g2_nand3_1 _1283_ (.B(_0421_),
    .C(_0437_),
    .A(_0372_),
    .Y(_0442_));
 sg13g2_xor2_1 _1284_ (.B(_0442_),
    .A(_0361_),
    .X(_0443_));
 sg13g2_nor2_1 _1285_ (.A(net32),
    .B(_0443_),
    .Y(_0089_));
 sg13g2_inv_2 _1286_ (.Y(_0444_),
    .A(_0442_));
 sg13g2_nand2_1 _1287_ (.Y(_0445_),
    .A(_0361_),
    .B(_0444_));
 sg13g2_xnor2_1 _1288_ (.Y(_0446_),
    .A(_0362_),
    .B(_0445_));
 sg13g2_and2_1 _1289_ (.A(_0261_),
    .B(_0446_),
    .X(_0090_));
 sg13g2_and2_1 _1290_ (.A(_0376_),
    .B(_0444_),
    .X(_0447_));
 sg13g2_xnor2_1 _1291_ (.Y(_0448_),
    .A(_0365_),
    .B(_0447_));
 sg13g2_nor2_1 _1292_ (.A(_0419_),
    .B(_0448_),
    .Y(_0091_));
 sg13g2_nand2_1 _1293_ (.Y(_0449_),
    .A(\vga_image_generator.counter[1] ),
    .B(\vga_image_generator.counter[0] ));
 sg13g2_xor2_1 _1294_ (.B(_0449_),
    .A(\vga_image_generator.counter[2] ),
    .X(_0450_));
 sg13g2_nor2_1 _1295_ (.A(net38),
    .B(_0450_),
    .Y(_0092_));
 sg13g2_nand3_1 _1296_ (.B(\vga_image_generator.counter[0] ),
    .C(\vga_image_generator.counter[2] ),
    .A(\vga_image_generator.counter[1] ),
    .Y(_0451_));
 sg13g2_xor2_1 _1297_ (.B(_0451_),
    .A(\vga_image_generator.counter[3] ),
    .X(_0452_));
 sg13g2_nor2_1 _1298_ (.A(net38),
    .B(_0452_),
    .Y(_0093_));
 sg13g2_xnor2_1 _1299_ (.Y(_0453_),
    .A(\vga_image_generator.counter[4] ),
    .B(_0401_));
 sg13g2_nor2_1 _1300_ (.A(net38),
    .B(_0453_),
    .Y(_0094_));
 sg13g2_nand2_1 _1301_ (.Y(_0454_),
    .A(\vga_image_generator.counter[4] ),
    .B(_0401_));
 sg13g2_xor2_1 _1302_ (.B(_0454_),
    .A(\vga_image_generator.counter[5] ),
    .X(_0455_));
 sg13g2_nor2_1 _1303_ (.A(net38),
    .B(_0455_),
    .Y(_0095_));
 sg13g2_nand3_1 _1304_ (.B(\vga_image_generator.counter[5] ),
    .C(_0401_),
    .A(\vga_image_generator.counter[4] ),
    .Y(_0456_));
 sg13g2_xor2_1 _1305_ (.B(_0456_),
    .A(\vga_image_generator.counter[6] ),
    .X(_0457_));
 sg13g2_nor2_1 _1306_ (.A(net38),
    .B(_0457_),
    .Y(_0096_));
 sg13g2_nand4_1 _1307_ (.B(\vga_image_generator.counter[5] ),
    .C(\vga_image_generator.counter[6] ),
    .A(\vga_image_generator.counter[4] ),
    .Y(_0458_),
    .D(_0401_));
 sg13g2_xor2_1 _1308_ (.B(_0458_),
    .A(\vga_image_generator.counter[7] ),
    .X(_0459_));
 sg13g2_nor2_1 _1309_ (.A(net38),
    .B(_0459_),
    .Y(_0097_));
 sg13g2_xnor2_1 _1310_ (.Y(_0460_),
    .A(_0399_),
    .B(_0404_));
 sg13g2_nor2_1 _1311_ (.A(net38),
    .B(_0460_),
    .Y(_0098_));
 sg13g2_xnor2_1 _1312_ (.Y(_0461_),
    .A(\vga_image_generator.counter[9] ),
    .B(_0405_));
 sg13g2_nor2_1 _1313_ (.A(net38),
    .B(_0461_),
    .Y(_0099_));
 sg13g2_buf_1 _1314_ (.A(ui_in[1]),
    .X(_0462_));
 sg13g2_buf_1 _1315_ (.A(net71),
    .X(_0463_));
 sg13g2_and2_1 _1316_ (.A(_0463_),
    .B(\BNC_x[0] ),
    .X(net3));
 sg13g2_and2_1 _1317_ (.A(net52),
    .B(\BNC_x[2] ),
    .X(net4));
 sg13g2_and2_1 _1318_ (.A(net52),
    .B(\BNC_x[4] ),
    .X(net5));
 sg13g2_and2_1 _1319_ (.A(_0463_),
    .B(\BNC_x[6] ),
    .X(net6));
 sg13g2_and2_1 _1320_ (.A(net52),
    .B(\BNC_x[1] ),
    .X(net7));
 sg13g2_and2_1 _1321_ (.A(net52),
    .B(\BNC_x[3] ),
    .X(net8));
 sg13g2_and2_1 _1322_ (.A(net52),
    .B(\BNC_x[5] ),
    .X(net9));
 sg13g2_and2_1 _1323_ (.A(net52),
    .B(\BNC_x[7] ),
    .X(net10));
 sg13g2_inv_1 _1324_ (.Y(_0464_),
    .A(net1));
 sg13g2_nor2_1 _1325_ (.A(_0160_),
    .B(_0462_),
    .Y(_0465_));
 sg13g2_a21oi_1 _1326_ (.A1(\BNC_y[0] ),
    .A2(_0462_),
    .Y(_0466_),
    .B1(_0465_));
 sg13g2_nor2_1 _1327_ (.A(_0125_),
    .B(_0135_),
    .Y(_0467_));
 sg13g2_nand2_1 _1328_ (.Y(_0468_),
    .A(_0344_),
    .B(_0467_));
 sg13g2_buf_1 _1329_ (.A(_0122_),
    .X(_0469_));
 sg13g2_a21oi_1 _1330_ (.A1(net50),
    .A2(_0468_),
    .Y(_0470_),
    .B1(net31));
 sg13g2_nand2b_1 _1331_ (.Y(_0471_),
    .B(net37),
    .A_N(_0024_));
 sg13g2_buf_1 _1332_ (.A(net56),
    .X(_0472_));
 sg13g2_nand2b_1 _1333_ (.Y(_0473_),
    .B(net35),
    .A_N(net63));
 sg13g2_nor2_1 _1334_ (.A(net30),
    .B(_0473_),
    .Y(_0474_));
 sg13g2_a21o_1 _1335_ (.A2(_0474_),
    .A1(_0471_),
    .B1(_0023_),
    .X(_0475_));
 sg13g2_nand3_1 _1336_ (.B(_0467_),
    .C(_0475_),
    .A(_0123_),
    .Y(_0476_));
 sg13g2_nor2b_1 _1337_ (.A(net55),
    .B_N(_0266_),
    .Y(_0477_));
 sg13g2_nor2b_2 _1338_ (.A(net56),
    .B_N(_0262_),
    .Y(_0478_));
 sg13g2_nor2b_1 _1339_ (.A(_0122_),
    .B_N(net62),
    .Y(_0479_));
 sg13g2_and3_1 _1340_ (.X(_0480_),
    .A(_0477_),
    .B(_0478_),
    .C(_0479_));
 sg13g2_nor2_1 _1341_ (.A(_0270_),
    .B(_0473_),
    .Y(_0481_));
 sg13g2_buf_1 _1342_ (.A(net62),
    .X(_0482_));
 sg13g2_nor2_1 _1343_ (.A(net29),
    .B(net31),
    .Y(_0483_));
 sg13g2_a21oi_1 _1344_ (.A1(_0480_),
    .A2(_0481_),
    .Y(_0484_),
    .B1(_0483_));
 sg13g2_a22oi_1 _1345_ (.Y(_0485_),
    .B1(_0476_),
    .B2(_0484_),
    .A2(_0470_),
    .A1(_0273_));
 sg13g2_a21oi_2 _1346_ (.B1(net31),
    .Y(_0486_),
    .A2(_0270_),
    .A1(net62));
 sg13g2_nand2b_2 _1347_ (.Y(_0487_),
    .B(\hvsync_gen.hpos[8] ),
    .A_N(_0135_));
 sg13g2_nand2b_1 _1348_ (.Y(_0488_),
    .B(_0125_),
    .A_N(net64));
 sg13g2_nor3_1 _1349_ (.A(_0122_),
    .B(_0487_),
    .C(_0488_),
    .Y(_0489_));
 sg13g2_nor2_1 _1350_ (.A(_0024_),
    .B(_0477_),
    .Y(_0490_));
 sg13g2_nor2b_1 _1351_ (.A(_0135_),
    .B_N(_0125_),
    .Y(_0491_));
 sg13g2_buf_1 _1352_ (.A(_0491_),
    .X(_0492_));
 sg13g2_nand2_1 _1353_ (.Y(_0493_),
    .A(_0479_),
    .B(net24));
 sg13g2_nor2b_1 _1354_ (.A(\hvsync_gen.hpos[4] ),
    .B_N(net64),
    .Y(_0494_));
 sg13g2_buf_2 _1355_ (.A(_0494_),
    .X(_0495_));
 sg13g2_nor2_2 _1356_ (.A(_0262_),
    .B(net56),
    .Y(_0496_));
 sg13g2_nand2_1 _1357_ (.Y(_0497_),
    .A(_0495_),
    .B(_0496_));
 sg13g2_nor3_1 _1358_ (.A(_0490_),
    .B(_0493_),
    .C(_0497_),
    .Y(_0498_));
 sg13g2_nor3_1 _1359_ (.A(_0486_),
    .B(_0489_),
    .C(_0498_),
    .Y(_0499_));
 sg13g2_nor2b_1 _1360_ (.A(net64),
    .B_N(\hvsync_gen.hpos[4] ),
    .Y(_0500_));
 sg13g2_buf_1 _1361_ (.A(_0500_),
    .X(_0501_));
 sg13g2_nand2_1 _1362_ (.Y(_0502_),
    .A(net23),
    .B(net24));
 sg13g2_nor2b_1 _1363_ (.A(_0262_),
    .B_N(net56),
    .Y(_0503_));
 sg13g2_buf_2 _1364_ (.A(_0503_),
    .X(_0504_));
 sg13g2_nand2_1 _1365_ (.Y(_0505_),
    .A(_0337_),
    .B(_0504_));
 sg13g2_and2_1 _1366_ (.A(_0262_),
    .B(net56),
    .X(_0506_));
 sg13g2_buf_1 _1367_ (.A(_0506_),
    .X(_0507_));
 sg13g2_and2_1 _1368_ (.A(net63),
    .B(net51),
    .X(_0508_));
 sg13g2_a221oi_1 _1369_ (.B2(_0508_),
    .C1(net49),
    .B1(net22),
    .A1(net35),
    .Y(_0509_),
    .A2(net51));
 sg13g2_o21ai_1 _1370_ (.B1(_0509_),
    .Y(_0510_),
    .A1(_0502_),
    .A2(_0505_));
 sg13g2_a21oi_1 _1371_ (.A1(net50),
    .A2(_0510_),
    .Y(_0511_),
    .B1(net31));
 sg13g2_nor2_1 _1372_ (.A(_0499_),
    .B(_0511_),
    .Y(_0512_));
 sg13g2_or2_1 _1373_ (.X(_0513_),
    .B(_0109_),
    .A(net68));
 sg13g2_buf_2 _1374_ (.A(_0513_),
    .X(_0514_));
 sg13g2_o21ai_1 _1375_ (.B1(net39),
    .Y(_0515_),
    .A1(\hvsync_gen.vpos[1] ),
    .A2(_0514_));
 sg13g2_nor2_2 _1376_ (.A(net67),
    .B(\hvsync_gen.vpos[9] ),
    .Y(_0516_));
 sg13g2_nand2b_1 _1377_ (.Y(_0517_),
    .B(_0516_),
    .A_N(_0121_));
 sg13g2_a21oi_1 _1378_ (.A1(_0313_),
    .A2(_0515_),
    .Y(_0518_),
    .B1(_0517_));
 sg13g2_o21ai_1 _1379_ (.B1(_0518_),
    .Y(_0519_),
    .A1(_0485_),
    .A2(_0512_));
 sg13g2_or2_1 _1380_ (.X(_0520_),
    .B(net56),
    .A(_0262_));
 sg13g2_buf_1 _1381_ (.A(_0520_),
    .X(_0521_));
 sg13g2_or2_1 _1382_ (.X(_0522_),
    .B(net36),
    .A(net55));
 sg13g2_o21ai_1 _1383_ (.B1(net35),
    .Y(_0523_),
    .A1(_0521_),
    .A2(_0522_));
 sg13g2_nand2_1 _1384_ (.Y(_0524_),
    .A(_0113_),
    .B(_0279_));
 sg13g2_nor2_1 _1385_ (.A(_0109_),
    .B(net53),
    .Y(_0525_));
 sg13g2_and2_1 _1386_ (.A(net54),
    .B(_0525_),
    .X(_0526_));
 sg13g2_nor4_2 _1387_ (.A(net66),
    .B(net65),
    .C(_0113_),
    .Y(_0527_),
    .D(\hvsync_gen.vpos[9] ));
 sg13g2_o21ai_1 _1388_ (.B1(_0527_),
    .Y(_0528_),
    .A1(_0021_),
    .A2(_0526_));
 sg13g2_nand2_1 _1389_ (.Y(_0529_),
    .A(_0524_),
    .B(_0528_));
 sg13g2_nand4_1 _1390_ (.B(_0298_),
    .C(_0527_),
    .A(_0296_),
    .Y(_0530_),
    .D(_0526_));
 sg13g2_nor3_1 _1391_ (.A(_0264_),
    .B(_0337_),
    .C(_0502_),
    .Y(_0531_));
 sg13g2_o21ai_1 _1392_ (.B1(_0479_),
    .Y(_0532_),
    .A1(_0509_),
    .A2(_0531_));
 sg13g2_a221oi_1 _1393_ (.B2(_0530_),
    .C1(_0532_),
    .B1(_0529_),
    .A1(_0467_),
    .Y(_0533_),
    .A2(_0523_));
 sg13g2_nand2_1 _1394_ (.Y(_0534_),
    .A(\hvsync_gen.vpos[5] ),
    .B(net53));
 sg13g2_nor2_1 _1395_ (.A(_0108_),
    .B(_0109_),
    .Y(_0535_));
 sg13g2_nor2_1 _1396_ (.A(_0534_),
    .B(_0535_),
    .Y(_0536_));
 sg13g2_o21ai_1 _1397_ (.B1(_0119_),
    .Y(_0537_),
    .A1(net65),
    .A2(_0536_));
 sg13g2_nor2_1 _1398_ (.A(_0348_),
    .B(_0128_),
    .Y(_0538_));
 sg13g2_and2_1 _1399_ (.A(_0538_),
    .B(_0504_),
    .X(_0539_));
 sg13g2_nand4_1 _1400_ (.B(_0479_),
    .C(net24),
    .A(_0267_),
    .Y(_0540_),
    .D(_0539_));
 sg13g2_nand2_1 _1401_ (.Y(_0541_),
    .A(net29),
    .B(_0123_));
 sg13g2_a21oi_1 _1402_ (.A1(net55),
    .A2(net37),
    .Y(_0542_),
    .B1(net30));
 sg13g2_nor3_1 _1403_ (.A(_0270_),
    .B(_0541_),
    .C(_0542_),
    .Y(_0543_));
 sg13g2_or2_1 _1404_ (.X(_0544_),
    .B(net63),
    .A(net56));
 sg13g2_nor2b_1 _1405_ (.A(_0544_),
    .B_N(_0489_),
    .Y(_0545_));
 sg13g2_a21oi_1 _1406_ (.A1(net28),
    .A2(_0543_),
    .Y(_0546_),
    .B1(_0545_));
 sg13g2_a22oi_1 _1407_ (.Y(_0547_),
    .B1(_0540_),
    .B2(_0546_),
    .A2(_0537_),
    .A1(_0516_));
 sg13g2_inv_1 _1408_ (.Y(_0548_),
    .A(net68));
 sg13g2_nor2_1 _1409_ (.A(_0548_),
    .B(_0110_),
    .Y(_0549_));
 sg13g2_a21oi_1 _1410_ (.A1(_0282_),
    .A2(_0549_),
    .Y(_0550_),
    .B1(_0116_));
 sg13g2_o21ai_1 _1411_ (.B1(_0527_),
    .Y(_0551_),
    .A1(_0021_),
    .A2(_0550_));
 sg13g2_nand2_1 _1412_ (.Y(_0552_),
    .A(_0524_),
    .B(_0551_));
 sg13g2_o21ai_1 _1413_ (.B1(_0552_),
    .Y(_0553_),
    .A1(_0533_),
    .A2(_0547_));
 sg13g2_o21ai_1 _1414_ (.B1(_0525_),
    .Y(_0554_),
    .A1(_0107_),
    .A2(_0548_));
 sg13g2_nand2_1 _1415_ (.Y(_0555_),
    .A(net54),
    .B(_0554_));
 sg13g2_nand2b_1 _1416_ (.Y(_0556_),
    .B(_0496_),
    .A_N(_0137_));
 sg13g2_o21ai_1 _1417_ (.B1(_0311_),
    .Y(_0557_),
    .A1(_0282_),
    .A2(_0514_));
 sg13g2_or2_1 _1418_ (.X(_0558_),
    .B(_0266_),
    .A(net55));
 sg13g2_buf_1 _1419_ (.A(_0558_),
    .X(_0559_));
 sg13g2_nand4_1 _1420_ (.B(net28),
    .C(net22),
    .A(net51),
    .Y(_0560_),
    .D(_0559_));
 sg13g2_nor3_1 _1421_ (.A(net31),
    .B(_0517_),
    .C(_0487_),
    .Y(_0561_));
 sg13g2_nand4_1 _1422_ (.B(_0557_),
    .C(_0560_),
    .A(_0556_),
    .Y(_0562_),
    .D(_0561_));
 sg13g2_o21ai_1 _1423_ (.B1(net31),
    .Y(_0563_),
    .A1(net49),
    .A2(_0482_));
 sg13g2_and3_1 _1424_ (.X(_0564_),
    .A(_0279_),
    .B(_0464_),
    .C(_0563_));
 sg13g2_o21ai_1 _1425_ (.B1(_0564_),
    .Y(_0565_),
    .A1(_0555_),
    .A2(_0562_));
 sg13g2_nand2b_1 _1426_ (.Y(_0566_),
    .B(net53),
    .A_N(_0109_));
 sg13g2_a21o_1 _1427_ (.A2(_0282_),
    .A1(_0296_),
    .B1(_0566_),
    .X(_0567_));
 sg13g2_nand2b_1 _1428_ (.Y(_0568_),
    .B(_0267_),
    .A_N(net37));
 sg13g2_and2_1 _1429_ (.A(net30),
    .B(net29),
    .X(_0569_));
 sg13g2_nand4_1 _1430_ (.B(_0486_),
    .C(_0568_),
    .A(net28),
    .Y(_0570_),
    .D(_0569_));
 sg13g2_and2_1 _1431_ (.A(_0538_),
    .B(net24),
    .X(_0571_));
 sg13g2_a22oi_1 _1432_ (.Y(_0572_),
    .B1(_0571_),
    .B2(_0480_),
    .A2(_0545_),
    .A1(_0471_));
 sg13g2_nor2b_1 _1433_ (.A(net65),
    .B_N(_0119_),
    .Y(_0573_));
 sg13g2_nand3_1 _1434_ (.B(_0516_),
    .C(_0573_),
    .A(net54),
    .Y(_0574_));
 sg13g2_a221oi_1 _1435_ (.B2(_0572_),
    .C1(_0574_),
    .B1(_0570_),
    .A1(_0309_),
    .Y(_0575_),
    .A2(_0567_));
 sg13g2_nand3_1 _1436_ (.B(net65),
    .C(net67),
    .A(net66),
    .Y(_0576_));
 sg13g2_a21oi_1 _1437_ (.A1(net41),
    .A2(_0282_),
    .Y(_0577_),
    .B1(_0566_));
 sg13g2_a21o_1 _1438_ (.A2(_0507_),
    .A1(_0265_),
    .B1(_0137_),
    .X(_0578_));
 sg13g2_nand2_1 _1439_ (.Y(_0579_),
    .A(_0267_),
    .B(_0496_));
 sg13g2_nand3_1 _1440_ (.B(net28),
    .C(_0579_),
    .A(net51),
    .Y(_0580_));
 sg13g2_nand4_1 _1441_ (.B(_0577_),
    .C(_0578_),
    .A(_0561_),
    .Y(_0581_),
    .D(_0580_));
 sg13g2_a21oi_1 _1442_ (.A1(_0576_),
    .A2(_0581_),
    .Y(_0582_),
    .B1(_0313_));
 sg13g2_a21oi_1 _1443_ (.A1(net37),
    .A2(_0559_),
    .Y(_0583_),
    .B1(net30));
 sg13g2_nand2b_1 _1444_ (.Y(_0584_),
    .B(net36),
    .A_N(_0583_));
 sg13g2_a21oi_1 _1445_ (.A1(_0489_),
    .A2(_0584_),
    .Y(_0585_),
    .B1(_0486_));
 sg13g2_o21ai_1 _1446_ (.B1(net50),
    .Y(_0586_),
    .A1(net28),
    .A2(_0270_));
 sg13g2_nor2_1 _1447_ (.A(net55),
    .B(_0266_),
    .Y(_0587_));
 sg13g2_o21ai_1 _1448_ (.B1(_0587_),
    .Y(_0588_),
    .A1(net36),
    .A2(_0270_));
 sg13g2_nand4_1 _1449_ (.B(net22),
    .C(_0468_),
    .A(net29),
    .Y(_0589_),
    .D(_0588_));
 sg13g2_and3_1 _1450_ (.X(_0590_),
    .A(_0123_),
    .B(_0586_),
    .C(_0589_));
 sg13g2_nor2_1 _1451_ (.A(_0548_),
    .B(_0292_),
    .Y(_0591_));
 sg13g2_nor2_1 _1452_ (.A(_0313_),
    .B(_0516_),
    .Y(_0592_));
 sg13g2_a22oi_1 _1453_ (.Y(_0593_),
    .B1(_0592_),
    .B2(_0554_),
    .A2(_0591_),
    .A1(_0526_));
 sg13g2_nor4_1 _1454_ (.A(_0528_),
    .B(_0585_),
    .C(_0590_),
    .D(_0593_),
    .Y(_0594_));
 sg13g2_nor4_1 _1455_ (.A(_0565_),
    .B(_0575_),
    .C(_0582_),
    .D(_0594_),
    .Y(_0595_));
 sg13g2_nand2b_1 _1456_ (.Y(_0596_),
    .B(net30),
    .A_N(net37));
 sg13g2_o21ai_1 _1457_ (.B1(_0025_),
    .Y(_0597_),
    .A1(_0596_),
    .A2(_0559_));
 sg13g2_nand2_1 _1458_ (.Y(_0598_),
    .A(net29),
    .B(_0495_));
 sg13g2_a21oi_1 _1459_ (.A1(net22),
    .A2(_0559_),
    .Y(_0599_),
    .B1(_0598_));
 sg13g2_a21oi_1 _1460_ (.A1(net23),
    .A2(_0597_),
    .Y(_0600_),
    .B1(_0599_));
 sg13g2_nor3_1 _1461_ (.A(_0270_),
    .B(_0541_),
    .C(_0600_),
    .Y(_0601_));
 sg13g2_a21o_1 _1462_ (.A2(_0587_),
    .A1(_0504_),
    .B1(_0025_),
    .X(_0602_));
 sg13g2_a22oi_1 _1463_ (.Y(_0603_),
    .B1(_0602_),
    .B2(_0495_),
    .A2(_0486_),
    .A1(net35));
 sg13g2_nand2_1 _1464_ (.Y(_0604_),
    .A(net23),
    .B(_0521_));
 sg13g2_a21oi_1 _1465_ (.A1(_0603_),
    .A2(_0604_),
    .Y(_0605_),
    .B1(_0493_));
 sg13g2_nand3b_1 _1466_ (.B(_0548_),
    .C(net40),
    .Y(_0606_),
    .A_N(_0282_));
 sg13g2_a21oi_1 _1467_ (.A1(net40),
    .A2(net53),
    .Y(_0607_),
    .B1(net54));
 sg13g2_o21ai_1 _1468_ (.B1(_0516_),
    .Y(_0608_),
    .A1(_0121_),
    .A2(_0607_));
 sg13g2_mux2_1 _1469_ (.A0(_0303_),
    .A1(_0606_),
    .S(_0608_),
    .X(_0609_));
 sg13g2_nor4_1 _1470_ (.A(net54),
    .B(_0307_),
    .C(_0517_),
    .D(_0609_),
    .Y(_0610_));
 sg13g2_o21ai_1 _1471_ (.B1(_0610_),
    .Y(_0611_),
    .A1(_0601_),
    .A2(_0605_));
 sg13g2_nand4_1 _1472_ (.B(_0553_),
    .C(_0595_),
    .A(_0519_),
    .Y(_0612_),
    .D(_0611_));
 sg13g2_buf_2 _1473_ (.A(_0612_),
    .X(_0613_));
 sg13g2_o21ai_1 _1474_ (.B1(_0613_),
    .Y(net11),
    .A1(_0464_),
    .A2(_0466_));
 sg13g2_buf_1 _1475_ (.A(net1),
    .X(_0614_));
 sg13g2_mux2_1 _1476_ (.A0(\BNC_y[5] ),
    .A1(\BNC_y[2] ),
    .S(net71),
    .X(_0615_));
 sg13g2_nand2_1 _1477_ (.Y(_0616_),
    .A(net70),
    .B(_0615_));
 sg13g2_nand2_1 _1478_ (.Y(_0617_),
    .A(net64),
    .B(net63));
 sg13g2_nor2_1 _1479_ (.A(net62),
    .B(_0617_),
    .Y(_0618_));
 sg13g2_nand4_1 _1480_ (.B(\vga_image_generator.character_hold[4] ),
    .C(net24),
    .A(_0124_),
    .Y(_0619_),
    .D(_0618_));
 sg13g2_buf_2 _1481_ (.A(_0026_),
    .X(_0620_));
 sg13g2_nand2b_1 _1482_ (.Y(_0621_),
    .B(\hvsync_gen.vpos[7] ),
    .A_N(\hvsync_gen.vpos[6] ));
 sg13g2_buf_2 _1483_ (.A(_0621_),
    .X(_0622_));
 sg13g2_nor4_2 _1484_ (.A(net68),
    .B(_0313_),
    .C(_0620_),
    .Y(_0623_),
    .D(_0622_));
 sg13g2_buf_1 _1485_ (.A(net2),
    .X(_0624_));
 sg13g2_nand2b_1 _1486_ (.Y(_0625_),
    .B(_0109_),
    .A_N(_0278_));
 sg13g2_nand2b_1 _1487_ (.Y(_0626_),
    .B(net69),
    .A_N(net40));
 sg13g2_o21ai_1 _1488_ (.B1(_0626_),
    .Y(_0627_),
    .A1(net69),
    .A2(_0625_));
 sg13g2_nor4_1 _1489_ (.A(_0620_),
    .B(_0534_),
    .C(_0514_),
    .D(_0622_),
    .Y(_0628_));
 sg13g2_buf_1 _1490_ (.A(_0628_),
    .X(_0629_));
 sg13g2_xor2_1 _1491_ (.B(_0263_),
    .A(_0262_),
    .X(_0630_));
 sg13g2_nor2_1 _1492_ (.A(net69),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_a22oi_1 _1493_ (.Y(_0632_),
    .B1(net20),
    .B2(_0631_),
    .A2(_0627_),
    .A1(_0623_));
 sg13g2_or2_1 _1494_ (.X(_0633_),
    .B(_0632_),
    .A(_0619_));
 sg13g2_inv_1 _1495_ (.Y(_0634_),
    .A(_0124_));
 sg13g2_nor3_2 _1496_ (.A(_0113_),
    .B(_0116_),
    .C(_0622_),
    .Y(_0635_));
 sg13g2_nor4_2 _1497_ (.A(net68),
    .B(_0620_),
    .C(_0116_),
    .Y(_0636_),
    .D(_0622_));
 sg13g2_a21oi_1 _1498_ (.A1(net22),
    .A2(_0635_),
    .Y(_0637_),
    .B1(_0636_));
 sg13g2_nor3_2 _1499_ (.A(_0125_),
    .B(_0135_),
    .C(_0131_),
    .Y(_0638_));
 sg13g2_nand3_1 _1500_ (.B(_0538_),
    .C(_0638_),
    .A(\vga_image_generator.character_hold[0] ),
    .Y(_0639_));
 sg13g2_or4_1 _1501_ (.A(_0110_),
    .B(_0634_),
    .C(_0637_),
    .D(_0639_),
    .X(_0640_));
 sg13g2_nor3_2 _1502_ (.A(_0620_),
    .B(_0116_),
    .C(_0622_),
    .Y(_0641_));
 sg13g2_nor4_2 _1503_ (.A(_0110_),
    .B(_0113_),
    .C(_0116_),
    .Y(_0642_),
    .D(_0622_));
 sg13g2_a22oi_1 _1504_ (.Y(_0643_),
    .B1(_0642_),
    .B2(_0335_),
    .A2(_0641_),
    .A1(_0111_));
 sg13g2_nand2_1 _1505_ (.Y(_0644_),
    .A(_0136_),
    .B(\vga_image_generator.character_hold[5] ));
 sg13g2_nor4_2 _1506_ (.A(net35),
    .B(net51),
    .C(_0131_),
    .Y(_0645_),
    .D(_0644_));
 sg13g2_nor2b_1 _1507_ (.A(net30),
    .B_N(net36),
    .Y(_0646_));
 sg13g2_nor2_1 _1508_ (.A(_0634_),
    .B(_0624_),
    .Y(_0647_));
 sg13g2_and2_1 _1509_ (.A(_0646_),
    .B(_0647_),
    .X(_0648_));
 sg13g2_nand3b_1 _1510_ (.B(_0645_),
    .C(_0648_),
    .Y(_0649_),
    .A_N(_0643_));
 sg13g2_a22oi_1 _1511_ (.Y(_0650_),
    .B1(_0504_),
    .B2(net23),
    .A2(_0495_),
    .A1(_0478_));
 sg13g2_inv_1 _1512_ (.Y(_0651_),
    .A(_0027_));
 sg13g2_nor2b_1 _1513_ (.A(_0125_),
    .B_N(_0135_),
    .Y(_0652_));
 sg13g2_and2_1 _1514_ (.A(_0651_),
    .B(_0652_),
    .X(_0653_));
 sg13g2_nand3b_1 _1515_ (.B(_0653_),
    .C(\vga_image_generator.character_hold[15] ),
    .Y(_0654_),
    .A_N(_0650_));
 sg13g2_nand2_1 _1516_ (.Y(_0655_),
    .A(_0126_),
    .B(net49));
 sg13g2_nor3_1 _1517_ (.A(net62),
    .B(_0617_),
    .C(_0655_),
    .Y(_0656_));
 sg13g2_nand3_1 _1518_ (.B(_0504_),
    .C(_0656_),
    .A(\vga_image_generator.character_hold[9] ),
    .Y(_0657_));
 sg13g2_nor2b_1 _1519_ (.A(_0278_),
    .B_N(\hvsync_gen.vpos[5] ),
    .Y(_0658_));
 sg13g2_nand3b_1 _1520_ (.B(_0658_),
    .C(_0573_),
    .Y(_0659_),
    .A_N(_0620_));
 sg13g2_buf_2 _1521_ (.A(_0659_),
    .X(_0660_));
 sg13g2_a21o_1 _1522_ (.A2(_0657_),
    .A1(_0654_),
    .B1(_0660_),
    .X(_0661_));
 sg13g2_and4_1 _1523_ (.A(_0633_),
    .B(_0640_),
    .C(_0649_),
    .D(_0661_),
    .X(_0662_));
 sg13g2_nand4_1 _1524_ (.B(\vga_image_generator.character_hold[12] ),
    .C(_0501_),
    .A(_0651_),
    .Y(_0663_),
    .D(net24));
 sg13g2_inv_1 _1525_ (.Y(_0664_),
    .A(\vga_image_generator.character_hold[11] ));
 sg13g2_nor3_1 _1526_ (.A(_0027_),
    .B(_0664_),
    .C(_0617_),
    .Y(_0665_));
 sg13g2_nand3_1 _1527_ (.B(_0504_),
    .C(_0665_),
    .A(_0467_),
    .Y(_0666_));
 sg13g2_o21ai_1 _1528_ (.B1(_0666_),
    .Y(_0667_),
    .A1(_0630_),
    .A2(_0663_));
 sg13g2_nand2_1 _1529_ (.Y(_0668_),
    .A(net41),
    .B(_0521_));
 sg13g2_a21oi_1 _1530_ (.A1(_0641_),
    .A2(_0668_),
    .Y(_0669_),
    .B1(net20));
 sg13g2_nand3_1 _1531_ (.B(\vga_image_generator.character_hold[10] ),
    .C(_0272_),
    .A(_0651_),
    .Y(_0670_));
 sg13g2_nor2_1 _1532_ (.A(_0669_),
    .B(_0670_),
    .Y(_0671_));
 sg13g2_a21oi_1 _1533_ (.A1(_0641_),
    .A2(_0667_),
    .Y(_0672_),
    .B1(_0671_));
 sg13g2_a22oi_1 _1534_ (.Y(_0673_),
    .B1(_0635_),
    .B2(_0496_),
    .A2(_0623_),
    .A1(net39));
 sg13g2_nor4_1 _1535_ (.A(net40),
    .B(_0634_),
    .C(_0639_),
    .D(_0673_),
    .Y(_0674_));
 sg13g2_nor2_1 _1536_ (.A(_0339_),
    .B(_0271_),
    .Y(_0675_));
 sg13g2_nor3_1 _1537_ (.A(_0344_),
    .B(net31),
    .C(_0544_),
    .Y(_0676_));
 sg13g2_a21oi_1 _1538_ (.A1(_0124_),
    .A2(_0675_),
    .Y(_0677_),
    .B1(_0676_));
 sg13g2_nand3_1 _1539_ (.B(_0638_),
    .C(_0641_),
    .A(\vga_image_generator.character_hold[1] ),
    .Y(_0678_));
 sg13g2_nor3_1 _1540_ (.A(_0514_),
    .B(_0677_),
    .C(_0678_),
    .Y(_0679_));
 sg13g2_nor2_1 _1541_ (.A(_0674_),
    .B(_0679_),
    .Y(_0680_));
 sg13g2_nor4_1 _1542_ (.A(_0339_),
    .B(net29),
    .C(_0617_),
    .D(_0655_),
    .Y(_0681_));
 sg13g2_nor3_1 _1543_ (.A(net30),
    .B(_0137_),
    .C(_0487_),
    .Y(_0682_));
 sg13g2_o21ai_1 _1544_ (.B1(\vga_image_generator.character_hold[9] ),
    .Y(_0683_),
    .A1(_0681_),
    .A2(_0682_));
 sg13g2_nor3_2 _1545_ (.A(_0313_),
    .B(_0620_),
    .C(_0622_),
    .Y(_0684_));
 sg13g2_nand2_1 _1546_ (.Y(_0685_),
    .A(_0535_),
    .B(_0684_));
 sg13g2_a21oi_1 _1547_ (.A1(_0663_),
    .A2(_0683_),
    .Y(_0686_),
    .B1(_0685_));
 sg13g2_xnor2_1 _1548_ (.Y(_0687_),
    .A(_0472_),
    .B(net63));
 sg13g2_nand4_1 _1549_ (.B(net49),
    .C(net62),
    .A(_0361_),
    .Y(_0688_),
    .D(\vga_image_generator.character_hold[17] ));
 sg13g2_nor2_1 _1550_ (.A(_0488_),
    .B(_0688_),
    .Y(_0689_));
 sg13g2_nand3_1 _1551_ (.B(_0126_),
    .C(\vga_image_generator.character_hold[13] ),
    .A(net35),
    .Y(_0690_));
 sg13g2_nor2_1 _1552_ (.A(_0487_),
    .B(_0690_),
    .Y(_0691_));
 sg13g2_a22oi_1 _1553_ (.Y(_0692_),
    .B1(_0691_),
    .B2(_0642_),
    .A2(_0689_),
    .A1(net20));
 sg13g2_nor2_1 _1554_ (.A(_0687_),
    .B(_0692_),
    .Y(_0693_));
 sg13g2_xor2_1 _1555_ (.B(_0472_),
    .A(net40),
    .X(_0694_));
 sg13g2_nor3_1 _1556_ (.A(_0548_),
    .B(net69),
    .C(_0694_),
    .Y(_0695_));
 sg13g2_o21ai_1 _1557_ (.B1(_0641_),
    .Y(_0696_),
    .A1(net22),
    .A2(_0695_));
 sg13g2_nor2_1 _1558_ (.A(_0619_),
    .B(_0696_),
    .Y(_0697_));
 sg13g2_nand2_1 _1559_ (.Y(_0698_),
    .A(_0684_),
    .B(_0645_));
 sg13g2_and2_1 _1560_ (.A(net36),
    .B(net69),
    .X(_0699_));
 sg13g2_nor3_1 _1561_ (.A(_0335_),
    .B(_0339_),
    .C(net36),
    .Y(_0700_));
 sg13g2_inv_1 _1562_ (.Y(_0701_),
    .A(net2));
 sg13g2_nand2_1 _1563_ (.Y(_0702_),
    .A(net31),
    .B(_0701_));
 sg13g2_a22oi_1 _1564_ (.Y(_0703_),
    .B1(_0700_),
    .B2(_0702_),
    .A2(_0699_),
    .A1(_0478_));
 sg13g2_nor3_1 _1565_ (.A(net39),
    .B(_0698_),
    .C(_0703_),
    .Y(_0704_));
 sg13g2_nor4_1 _1566_ (.A(_0686_),
    .B(_0693_),
    .C(_0697_),
    .D(_0704_),
    .Y(_0705_));
 sg13g2_nand4_1 _1567_ (.B(_0672_),
    .C(_0680_),
    .A(_0662_),
    .Y(_0706_),
    .D(_0705_));
 sg13g2_nand3_1 _1568_ (.B(net28),
    .C(_0653_),
    .A(\vga_image_generator.character_hold[16] ),
    .Y(_0707_));
 sg13g2_xnor2_1 _1569_ (.Y(_0708_),
    .A(_0305_),
    .B(_0630_));
 sg13g2_a22oi_1 _1570_ (.Y(_0709_),
    .B1(_0635_),
    .B2(_0708_),
    .A2(_0630_),
    .A1(net20));
 sg13g2_nor2_1 _1571_ (.A(_0707_),
    .B(_0709_),
    .Y(_0710_));
 sg13g2_nand4_1 _1572_ (.B(\vga_image_generator.character_hold[16] ),
    .C(_0130_),
    .A(_0132_),
    .Y(_0711_),
    .D(_0652_));
 sg13g2_nor4_1 _1573_ (.A(net41),
    .B(_0110_),
    .C(_0660_),
    .D(_0711_),
    .Y(_0712_));
 sg13g2_nor2_1 _1574_ (.A(net20),
    .B(_0641_),
    .Y(_0713_));
 sg13g2_and2_1 _1575_ (.A(net37),
    .B(_0646_),
    .X(_0714_));
 sg13g2_nor3_1 _1576_ (.A(_0136_),
    .B(_0027_),
    .C(_0690_),
    .Y(_0715_));
 sg13g2_o21ai_1 _1577_ (.B1(_0715_),
    .Y(_0716_),
    .A1(_0700_),
    .A2(_0714_));
 sg13g2_nor2_1 _1578_ (.A(_0713_),
    .B(_0716_),
    .Y(_0717_));
 sg13g2_nand4_1 _1579_ (.B(\vga_image_generator.character_hold[2] ),
    .C(net28),
    .A(_0624_),
    .Y(_0718_),
    .D(_0638_));
 sg13g2_nand2_1 _1580_ (.Y(_0719_),
    .A(net54),
    .B(_0124_));
 sg13g2_nor4_1 _1581_ (.A(_0620_),
    .B(_0622_),
    .C(_0718_),
    .D(_0719_),
    .Y(_0720_));
 sg13g2_a21oi_1 _1582_ (.A1(_0625_),
    .A2(_0566_),
    .Y(_0721_),
    .B1(net68));
 sg13g2_a21o_1 _1583_ (.A2(_0496_),
    .A1(_0307_),
    .B1(_0721_),
    .X(_0722_));
 sg13g2_nor2_1 _1584_ (.A(_0122_),
    .B(_0620_),
    .Y(_0723_));
 sg13g2_nand4_1 _1585_ (.B(_0535_),
    .C(_0573_),
    .A(_0658_),
    .Y(_0724_),
    .D(_0723_));
 sg13g2_a21oi_1 _1586_ (.A1(_0639_),
    .A2(_0718_),
    .Y(_0725_),
    .B1(_0724_));
 sg13g2_a21o_1 _1587_ (.A2(_0722_),
    .A1(_0720_),
    .B1(_0725_),
    .X(_0726_));
 sg13g2_nor4_1 _1588_ (.A(_0710_),
    .B(_0712_),
    .C(_0717_),
    .D(_0726_),
    .Y(_0727_));
 sg13g2_nor2_1 _1589_ (.A(_0514_),
    .B(_0687_),
    .Y(_0728_));
 sg13g2_mux2_1 _1590_ (.A0(_0647_),
    .A1(_0702_),
    .S(net39),
    .X(_0729_));
 sg13g2_nand4_1 _1591_ (.B(_0645_),
    .C(_0728_),
    .A(_0684_),
    .Y(_0730_),
    .D(_0729_));
 sg13g2_o21ai_1 _1592_ (.B1(net41),
    .Y(_0731_),
    .A1(net39),
    .A2(_0630_));
 sg13g2_nand2_1 _1593_ (.Y(_0732_),
    .A(_0305_),
    .B(net53));
 sg13g2_and3_1 _1594_ (.X(_0733_),
    .A(\vga_image_generator.character_hold[14] ),
    .B(_0538_),
    .C(_0732_));
 sg13g2_nand4_1 _1595_ (.B(_0653_),
    .C(_0731_),
    .A(_0684_),
    .Y(_0734_),
    .D(_0733_));
 sg13g2_nor2_1 _1596_ (.A(net29),
    .B(_0655_),
    .Y(_0735_));
 sg13g2_nand4_1 _1597_ (.B(_0495_),
    .C(_0636_),
    .A(\vga_image_generator.character_hold[8] ),
    .Y(_0736_),
    .D(_0735_));
 sg13g2_nand4_1 _1598_ (.B(net35),
    .C(net36),
    .A(net30),
    .Y(_0737_),
    .D(_0347_));
 sg13g2_o21ai_1 _1599_ (.B1(_0737_),
    .Y(_0738_),
    .A1(_0544_),
    .A2(_0488_));
 sg13g2_nor2_1 _1600_ (.A(_0664_),
    .B(_0487_),
    .Y(_0739_));
 sg13g2_nand4_1 _1601_ (.B(_0684_),
    .C(_0738_),
    .A(_0535_),
    .Y(_0740_),
    .D(_0739_));
 sg13g2_and4_1 _1602_ (.A(_0730_),
    .B(_0734_),
    .C(_0736_),
    .D(_0740_),
    .X(_0741_));
 sg13g2_nand3_1 _1603_ (.B(_0495_),
    .C(_0735_),
    .A(\vga_image_generator.character_hold[8] ),
    .Y(_0742_));
 sg13g2_nor3_1 _1604_ (.A(_0630_),
    .B(_0713_),
    .C(_0742_),
    .Y(_0743_));
 sg13g2_nand3_1 _1605_ (.B(_0492_),
    .C(_0618_),
    .A(\vga_image_generator.character_hold[4] ),
    .Y(_0744_));
 sg13g2_nor4_1 _1606_ (.A(_0469_),
    .B(_0521_),
    .C(_0744_),
    .D(_0660_),
    .Y(_0745_));
 sg13g2_nand3_1 _1607_ (.B(_0658_),
    .C(_0573_),
    .A(_0112_),
    .Y(_0746_));
 sg13g2_nand2_1 _1608_ (.Y(_0747_),
    .A(net23),
    .B(_0478_));
 sg13g2_nand2_1 _1609_ (.Y(_0748_),
    .A(\vga_image_generator.character_hold[7] ),
    .B(_0735_));
 sg13g2_nor4_1 _1610_ (.A(net40),
    .B(_0746_),
    .C(_0747_),
    .D(_0748_),
    .Y(_0749_));
 sg13g2_mux2_1 _1611_ (.A0(net23),
    .A1(_0495_),
    .S(_0339_),
    .X(_0750_));
 sg13g2_nand4_1 _1612_ (.B(\vga_image_generator.character_hold[15] ),
    .C(_0652_),
    .A(_0132_),
    .Y(_0751_),
    .D(_0750_));
 sg13g2_nor2_1 _1613_ (.A(_0685_),
    .B(_0751_),
    .Y(_0752_));
 sg13g2_nor4_1 _1614_ (.A(_0743_),
    .B(_0745_),
    .C(_0749_),
    .D(_0752_),
    .Y(_0753_));
 sg13g2_or4_1 _1615_ (.A(_0482_),
    .B(_0469_),
    .C(_0521_),
    .D(_0660_),
    .X(_0754_));
 sg13g2_nand3_1 _1616_ (.B(_0027_),
    .C(net20),
    .A(_0124_),
    .Y(_0755_));
 sg13g2_nand3_1 _1617_ (.B(\vga_image_generator.character_hold[2] ),
    .C(_0571_),
    .A(_0701_),
    .Y(_0756_));
 sg13g2_a21oi_1 _1618_ (.A1(_0754_),
    .A2(_0755_),
    .Y(_0757_),
    .B1(_0756_));
 sg13g2_mux2_1 _1619_ (.A0(net22),
    .A1(_0496_),
    .S(_0110_),
    .X(_0758_));
 sg13g2_a221oi_1 _1620_ (.B2(_0758_),
    .C1(_0629_),
    .B1(_0635_),
    .A1(_0307_),
    .Y(_0759_),
    .A2(_0623_));
 sg13g2_nand3_1 _1621_ (.B(_0618_),
    .C(_0652_),
    .A(\vga_image_generator.character_hold[6] ),
    .Y(_0760_));
 sg13g2_nor2_1 _1622_ (.A(_0759_),
    .B(_0760_),
    .Y(_0761_));
 sg13g2_nor2_1 _1623_ (.A(_0348_),
    .B(_0687_),
    .Y(_0762_));
 sg13g2_a21oi_1 _1624_ (.A1(_0636_),
    .A2(_0762_),
    .Y(_0763_),
    .B1(_0539_));
 sg13g2_nor3_1 _1625_ (.A(_0713_),
    .B(_0748_),
    .C(_0763_),
    .Y(_0764_));
 sg13g2_o21ai_1 _1626_ (.B1(_0566_),
    .Y(_0765_),
    .A1(_0701_),
    .A2(_0625_));
 sg13g2_nand3_1 _1627_ (.B(_0750_),
    .C(_0765_),
    .A(_0623_),
    .Y(_0766_));
 sg13g2_o21ai_1 _1628_ (.B1(net69),
    .Y(_0767_),
    .A1(_0271_),
    .A2(_0596_));
 sg13g2_nand3b_1 _1629_ (.B(_0767_),
    .C(_0641_),
    .Y(_0768_),
    .A_N(_0650_));
 sg13g2_nand3_1 _1630_ (.B(\vga_image_generator.character_hold[1] ),
    .C(_0638_),
    .A(_0124_),
    .Y(_0769_));
 sg13g2_a21oi_1 _1631_ (.A1(_0766_),
    .A2(_0768_),
    .Y(_0770_),
    .B1(_0769_));
 sg13g2_nor4_1 _1632_ (.A(_0757_),
    .B(_0761_),
    .C(_0764_),
    .D(_0770_),
    .Y(_0771_));
 sg13g2_nand4_1 _1633_ (.B(_0741_),
    .C(_0753_),
    .A(_0727_),
    .Y(_0772_),
    .D(_0771_));
 sg13g2_inv_1 _1634_ (.Y(_0773_),
    .A(\vga_image_generator.character_hold[3] ));
 sg13g2_nand2_1 _1635_ (.Y(_0774_),
    .A(_0478_),
    .B(_0495_));
 sg13g2_nand3b_1 _1636_ (.B(_0124_),
    .C(net24),
    .Y(_0775_),
    .A_N(net29));
 sg13g2_buf_1 _1637_ (.A(_0775_),
    .X(_0776_));
 sg13g2_nand4_1 _1638_ (.B(_0483_),
    .C(net24),
    .A(net23),
    .Y(_0777_),
    .D(_0504_));
 sg13g2_o21ai_1 _1639_ (.B1(_0777_),
    .Y(_0778_),
    .A1(_0774_),
    .A2(_0776_));
 sg13g2_nor2_1 _1640_ (.A(net40),
    .B(_0746_),
    .Y(_0779_));
 sg13g2_or2_1 _1641_ (.X(_0780_),
    .B(_0642_),
    .A(net20));
 sg13g2_nand2_1 _1642_ (.Y(_0781_),
    .A(net22),
    .B(net23));
 sg13g2_a21oi_1 _1643_ (.A1(_0497_),
    .A2(_0781_),
    .Y(_0782_),
    .B1(_0776_));
 sg13g2_nand3_1 _1644_ (.B(_0641_),
    .C(_0750_),
    .A(_0111_),
    .Y(_0783_));
 sg13g2_o21ai_1 _1645_ (.B1(net69),
    .Y(_0784_),
    .A1(_0776_),
    .A2(_0783_));
 sg13g2_a221oi_1 _1646_ (.B2(_0782_),
    .C1(_0784_),
    .B1(_0780_),
    .A1(_0778_),
    .Y(_0785_),
    .A2(_0779_));
 sg13g2_a21oi_1 _1647_ (.A1(net20),
    .A2(_0675_),
    .Y(_0786_),
    .B1(_0474_));
 sg13g2_nor3_1 _1648_ (.A(_0685_),
    .B(_0776_),
    .C(_0786_),
    .Y(_0787_));
 sg13g2_nor3_1 _1649_ (.A(_0660_),
    .B(_0650_),
    .C(_0776_),
    .Y(_0788_));
 sg13g2_nor4_1 _1650_ (.A(_0339_),
    .B(net50),
    .C(_0502_),
    .D(_0724_),
    .Y(_0789_));
 sg13g2_nor4_1 _1651_ (.A(net69),
    .B(_0787_),
    .C(_0788_),
    .D(_0789_),
    .Y(_0790_));
 sg13g2_nor3_1 _1652_ (.A(_0773_),
    .B(_0785_),
    .C(_0790_),
    .Y(_0791_));
 sg13g2_nor3_2 _1653_ (.A(_0706_),
    .B(_0772_),
    .C(_0791_),
    .Y(_0792_));
 sg13g2_a21oi_1 _1654_ (.A1(net70),
    .A2(_0615_),
    .Y(_0793_),
    .B1(_0113_));
 sg13g2_a22oi_1 _1655_ (.Y(net12),
    .B1(_0792_),
    .B2(_0793_),
    .A2(_0616_),
    .A1(_0613_));
 sg13g2_mux2_1 _1656_ (.A0(\BNC_x[7] ),
    .A1(\BNC_y[4] ),
    .S(net71),
    .X(_0794_));
 sg13g2_nand2_1 _1657_ (.Y(_0795_),
    .A(net70),
    .B(_0794_));
 sg13g2_o21ai_1 _1658_ (.B1(_0795_),
    .Y(net13),
    .A1(_0613_),
    .A2(_0792_));
 sg13g2_nor2b_1 _1659_ (.A(net71),
    .B_N(\BNC_x[5] ),
    .Y(_0796_));
 sg13g2_a21oi_1 _1660_ (.A1(net52),
    .A2(\BNC_y[6] ),
    .Y(_0797_),
    .B1(_0796_));
 sg13g2_nor2_1 _1661_ (.A(_0614_),
    .B(\hvsync_gen.vsync ),
    .Y(_0798_));
 sg13g2_a21oi_1 _1662_ (.A1(_0614_),
    .A2(_0797_),
    .Y(net14),
    .B1(_0798_));
 sg13g2_mux2_1 _1663_ (.A0(\BNC_y[6] ),
    .A1(\BNC_y[1] ),
    .S(net71),
    .X(_0799_));
 sg13g2_nand2_1 _1664_ (.Y(_0800_),
    .A(net70),
    .B(_0799_));
 sg13g2_and3_1 _1665_ (.X(_0801_),
    .A(net66),
    .B(net67),
    .C(_0800_));
 sg13g2_a22oi_1 _1666_ (.Y(net15),
    .B1(_0801_),
    .B2(_0792_),
    .A2(_0800_),
    .A1(_0613_));
 sg13g2_mux2_1 _1667_ (.A0(\BNC_y[4] ),
    .A1(\BNC_y[3] ),
    .S(net71),
    .X(_0802_));
 sg13g2_nand2_1 _1668_ (.Y(_0100_),
    .A(net70),
    .B(_0802_));
 sg13g2_and2_1 _1669_ (.A(net66),
    .B(_0100_),
    .X(_0101_));
 sg13g2_a22oi_1 _1670_ (.Y(net16),
    .B1(_0101_),
    .B2(_0792_),
    .A2(_0100_),
    .A1(_0613_));
 sg13g2_mux2_1 _1671_ (.A0(\BNC_x[6] ),
    .A1(\BNC_y[5] ),
    .S(net71),
    .X(_0102_));
 sg13g2_nand2_1 _1672_ (.Y(_0103_),
    .A(net70),
    .B(_0102_));
 sg13g2_o21ai_1 _1673_ (.B1(_0103_),
    .Y(net17),
    .A1(_0613_),
    .A2(_0792_));
 sg13g2_nor2b_1 _1674_ (.A(net71),
    .B_N(\BNC_x[4] ),
    .Y(_0104_));
 sg13g2_a21oi_1 _1675_ (.A1(_0140_),
    .A2(net52),
    .Y(_0105_),
    .B1(_0104_));
 sg13g2_nor2_1 _1676_ (.A(net70),
    .B(hsync),
    .Y(_0106_));
 sg13g2_a21oi_1 _1677_ (.A1(net70),
    .A2(_0105_),
    .Y(net18),
    .B1(_0106_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _1679_ (.A(net72),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1680_ (.A(net73),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1681_ (.A(net74),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1682_ (.A(net75),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1683_ (.A(net76),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1684_ (.A(net77),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1685_ (.A(net78),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1686_ (.A(net79),
    .X(uio_oe[7]));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[0]$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net80),
    .D(_0000_),
    .Q_N(_0858_),
    .Q(\BNC_x[0] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[1]$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net81),
    .D(_0001_),
    .Q_N(_0859_),
    .Q(\BNC_x[1] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[2]$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net82),
    .D(_0002_),
    .Q_N(_0860_),
    .Q(\BNC_x[2] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[3]$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net83),
    .D(_0003_),
    .Q_N(_0861_),
    .Q(\BNC_x[3] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[4]$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net84),
    .D(_0004_),
    .Q_N(_0862_),
    .Q(\BNC_x[4] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[5]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net85),
    .D(_0005_),
    .Q_N(_0863_),
    .Q(\BNC_x[5] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[6]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net86),
    .D(_0006_),
    .Q_N(_0864_),
    .Q(\BNC_x[6] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_x[7]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net87),
    .D(_0007_),
    .Q_N(_0865_),
    .Q(\BNC_x[7] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[0]$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net88),
    .D(_0008_),
    .Q_N(_0866_),
    .Q(\BNC_y[0] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[1]$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net89),
    .D(_0009_),
    .Q_N(_0867_),
    .Q(\BNC_y[1] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[2]$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net90),
    .D(_0010_),
    .Q_N(_0868_),
    .Q(\BNC_y[2] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[3]$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net91),
    .D(_0011_),
    .Q_N(_0869_),
    .Q(\BNC_y[3] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[4]$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net92),
    .D(_0012_),
    .Q_N(_0870_),
    .Q(\BNC_y[4] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[5]$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net93),
    .D(_0013_),
    .Q_N(_0871_),
    .Q(\BNC_y[5] ));
 sg13g2_dfrbp_1 \bnc_image_generator.BNC_y[6]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net94),
    .D(_0014_),
    .Q_N(_0857_),
    .Q(\BNC_y[6] ));
 sg13g2_dfrbp_1 \bnc_image_generator.counter[0]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net95),
    .D(_0032_),
    .Q_N(_0030_),
    .Q(\bnc_image_generator.counter[0] ));
 sg13g2_dfrbp_1 \bnc_image_generator.counter[1]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net96),
    .D(_0033_),
    .Q_N(_0019_),
    .Q(\bnc_image_generator.counter[1] ));
 sg13g2_dfrbp_1 \bnc_image_generator.counter[2]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net97),
    .D(_0034_),
    .Q_N(_0018_),
    .Q(\bnc_image_generator.counter[2] ));
 sg13g2_dfrbp_1 \bnc_image_generator.counter[3]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net98),
    .D(_0035_),
    .Q_N(_0017_),
    .Q(BNC_trig));
 sg13g2_dfrbp_1 \bnc_image_generator.counter[4]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net99),
    .D(_0036_),
    .Q_N(_0856_),
    .Q(\bnc_image_generator.counter[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[0]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net100),
    .D(_0037_),
    .Q_N(_0028_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[1]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net101),
    .D(_0038_),
    .Q_N(_0024_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[2]$_SDFF_PP0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net102),
    .D(_0039_),
    .Q_N(_0855_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[3]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net103),
    .D(_0040_),
    .Q_N(_0025_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[4]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net104),
    .D(_0041_),
    .Q_N(_0854_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[5]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net105),
    .D(_0042_),
    .Q_N(_0023_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[6]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net106),
    .D(_0043_),
    .Q_N(_0853_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[7]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net107),
    .D(_0044_),
    .Q_N(_0852_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[8]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net108),
    .D(_0045_),
    .Q_N(_0027_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[9]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net109),
    .D(_0046_),
    .Q_N(_0022_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.hsync$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net110),
    .D(_0015_),
    .Q_N(_0851_),
    .Q(hsync));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[0]$_SDFFCE_PP0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net111),
    .D(_0047_),
    .Q_N(_0029_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[1]$_SDFFCE_PP0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net112),
    .D(_0048_),
    .Q_N(_0850_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[2]$_SDFFCE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net113),
    .D(_0049_),
    .Q_N(_0849_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[3]$_SDFFCE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net114),
    .D(_0050_),
    .Q_N(_0848_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[4]$_SDFFCE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net115),
    .D(_0051_),
    .Q_N(_0847_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[5]$_SDFFCE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net116),
    .D(_0052_),
    .Q_N(_0021_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[6]$_SDFFCE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net117),
    .D(_0053_),
    .Q_N(_0846_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[7]$_SDFFCE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net118),
    .D(_0054_),
    .Q_N(_0845_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[8]$_SDFFCE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net119),
    .D(_0055_),
    .Q_N(_0026_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[9]$_SDFFCE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net120),
    .D(_0056_),
    .Q_N(_0872_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.vsync$_DFF_P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net121),
    .D(_0016_),
    .Q_N(_0844_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[0]$_SDFFE_PN0N_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net122),
    .D(_0057_),
    .Q_N(_0843_),
    .Q(\vga_image_generator.character_hold[0] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[10]$_SDFFE_PN0N_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net123),
    .D(_0058_),
    .Q_N(_0842_),
    .Q(\vga_image_generator.character_hold[10] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[11]$_SDFFE_PN0N_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net124),
    .D(_0059_),
    .Q_N(_0841_),
    .Q(\vga_image_generator.character_hold[11] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[12]$_SDFFE_PN0N_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net125),
    .D(_0060_),
    .Q_N(_0840_),
    .Q(\vga_image_generator.character_hold[12] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[13]$_SDFFE_PN0N_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net126),
    .D(_0061_),
    .Q_N(_0839_),
    .Q(\vga_image_generator.character_hold[13] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[14]$_SDFFE_PN0N_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net127),
    .D(_0062_),
    .Q_N(_0838_),
    .Q(\vga_image_generator.character_hold[14] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[15]$_SDFFE_PN0N_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net128),
    .D(_0063_),
    .Q_N(_0837_),
    .Q(\vga_image_generator.character_hold[15] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[16]$_SDFFE_PN0N_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net129),
    .D(_0064_),
    .Q_N(_0836_),
    .Q(\vga_image_generator.character_hold[16] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[17]$_SDFFE_PN0N_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net130),
    .D(_0065_),
    .Q_N(_0835_),
    .Q(\vga_image_generator.character_hold[17] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[1]$_SDFFE_PN0N_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net131),
    .D(_0066_),
    .Q_N(_0834_),
    .Q(\vga_image_generator.character_hold[1] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[2]$_SDFFE_PN0N_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net132),
    .D(_0067_),
    .Q_N(_0833_),
    .Q(\vga_image_generator.character_hold[2] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[3]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net133),
    .D(_0068_),
    .Q_N(_0832_),
    .Q(\vga_image_generator.character_hold[3] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[4]$_SDFFE_PN0N_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net134),
    .D(_0069_),
    .Q_N(_0831_),
    .Q(\vga_image_generator.character_hold[4] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[5]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net135),
    .D(_0070_),
    .Q_N(_0830_),
    .Q(\vga_image_generator.character_hold[5] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[6]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net136),
    .D(_0071_),
    .Q_N(_0829_),
    .Q(\vga_image_generator.character_hold[6] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[7]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net137),
    .D(_0072_),
    .Q_N(_0828_),
    .Q(\vga_image_generator.character_hold[7] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[8]$_SDFFE_PN0N_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net138),
    .D(_0073_),
    .Q_N(_0827_),
    .Q(\vga_image_generator.character_hold[8] ));
 sg13g2_dfrbp_1 \vga_image_generator.character_hold[9]$_SDFFE_PN0N_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net139),
    .D(_0074_),
    .Q_N(_0826_),
    .Q(\vga_image_generator.character_hold[9] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[0]$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net140),
    .D(_0075_),
    .Q_N(_0031_),
    .Q(\vga_image_generator.counter[0] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[10]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net141),
    .D(_0076_),
    .Q_N(_0825_),
    .Q(\vga_image_generator.counter[10] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[11]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net142),
    .D(_0077_),
    .Q_N(_0824_),
    .Q(\vga_image_generator.counter[11] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[12]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net143),
    .D(_0078_),
    .Q_N(_0823_),
    .Q(\vga_image_generator.counter[12] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[13]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net144),
    .D(_0079_),
    .Q_N(_0822_),
    .Q(\vga_image_generator.counter[13] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[14]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net145),
    .D(_0080_),
    .Q_N(_0821_),
    .Q(\vga_image_generator.counter[14] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[15]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net146),
    .D(_0081_),
    .Q_N(_0820_),
    .Q(\vga_image_generator.counter[15] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[16]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net147),
    .D(_0082_),
    .Q_N(_0819_),
    .Q(\vga_image_generator.counter[16] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[17]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net148),
    .D(_0083_),
    .Q_N(_0818_),
    .Q(\vga_image_generator.counter[17] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[18]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net149),
    .D(_0084_),
    .Q_N(_0817_),
    .Q(\vga_image_generator.counter[18] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[19]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net150),
    .D(_0085_),
    .Q_N(_0816_),
    .Q(\vga_image_generator.counter[19] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[1]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net151),
    .D(_0086_),
    .Q_N(_0815_),
    .Q(\vga_image_generator.counter[1] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[20]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net152),
    .D(_0087_),
    .Q_N(_0814_),
    .Q(\vga_image_generator.counter[20] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[21]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net153),
    .D(_0088_),
    .Q_N(_0813_),
    .Q(\vga_image_generator.counter[21] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[22]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net154),
    .D(_0089_),
    .Q_N(_0812_),
    .Q(\vga_image_generator.counter[22] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[23]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net155),
    .D(_0090_),
    .Q_N(_0811_),
    .Q(\vga_image_generator.counter[23] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[24]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net156),
    .D(_0091_),
    .Q_N(_0020_),
    .Q(\vga_image_generator.counter[24] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[2]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net157),
    .D(_0092_),
    .Q_N(_0810_),
    .Q(\vga_image_generator.counter[2] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[3]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net158),
    .D(_0093_),
    .Q_N(_0809_),
    .Q(\vga_image_generator.counter[3] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[4]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net159),
    .D(_0094_),
    .Q_N(_0808_),
    .Q(\vga_image_generator.counter[4] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[5]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net160),
    .D(_0095_),
    .Q_N(_0807_),
    .Q(\vga_image_generator.counter[5] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[6]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net161),
    .D(_0096_),
    .Q_N(_0806_),
    .Q(\vga_image_generator.counter[6] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[7]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net162),
    .D(_0097_),
    .Q_N(_0805_),
    .Q(\vga_image_generator.counter[7] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[8]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net163),
    .D(_0098_),
    .Q_N(_0804_),
    .Q(\vga_image_generator.counter[8] ));
 sg13g2_dfrbp_1 \vga_image_generator.counter[9]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net164),
    .D(_0099_),
    .Q_N(_0803_),
    .Q(\vga_image_generator.counter[9] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_out[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_out[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout19 (.A(_0276_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0629_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0287_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0507_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0501_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0492_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0333_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0188_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0177_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0130_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0482_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0472_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0469_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0419_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0393_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0374_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0348_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0342_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0335_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0332_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0311_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0305_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0296_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0170_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0160_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0153_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0152_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0145_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0142_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0140_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0136_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0132_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0126_),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(_0463_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0278_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0277_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0265_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0263_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0151_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0147_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0143_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0141_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0139_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0131_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0128_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0127_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0120_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0119_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0112_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0108_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0624_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0614_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0462_),
    .X(net71));
 sg13g2_tiehi _1679__72 (.L_HI(net72));
 sg13g2_tiehi _1680__73 (.L_HI(net73));
 sg13g2_tiehi _1681__74 (.L_HI(net74));
 sg13g2_tiehi _1682__75 (.L_HI(net75));
 sg13g2_tiehi _1683__76 (.L_HI(net76));
 sg13g2_tiehi _1684__77 (.L_HI(net77));
 sg13g2_tiehi _1685__78 (.L_HI(net78));
 sg13g2_tiehi _1686__79 (.L_HI(net79));
 sg13g2_tiehi \bnc_image_generator.BNC_x[0]$_DFF_P__80  (.L_HI(net80));
 sg13g2_tiehi \bnc_image_generator.BNC_x[1]$_DFF_P__81  (.L_HI(net81));
 sg13g2_tiehi \bnc_image_generator.BNC_x[2]$_DFF_P__82  (.L_HI(net82));
 sg13g2_tiehi \bnc_image_generator.BNC_x[3]$_DFF_P__83  (.L_HI(net83));
 sg13g2_tiehi \bnc_image_generator.BNC_x[4]$_DFF_P__84  (.L_HI(net84));
 sg13g2_tiehi \bnc_image_generator.BNC_x[5]$_DFF_P__85  (.L_HI(net85));
 sg13g2_tiehi \bnc_image_generator.BNC_x[6]$_DFF_P__86  (.L_HI(net86));
 sg13g2_tiehi \bnc_image_generator.BNC_x[7]$_DFF_P__87  (.L_HI(net87));
 sg13g2_tiehi \bnc_image_generator.BNC_y[0]$_DFF_P__88  (.L_HI(net88));
 sg13g2_tiehi \bnc_image_generator.BNC_y[1]$_DFF_P__89  (.L_HI(net89));
 sg13g2_tiehi \bnc_image_generator.BNC_y[2]$_DFF_P__90  (.L_HI(net90));
 sg13g2_tiehi \bnc_image_generator.BNC_y[3]$_DFF_P__91  (.L_HI(net91));
 sg13g2_tiehi \bnc_image_generator.BNC_y[4]$_DFF_P__92  (.L_HI(net92));
 sg13g2_tiehi \bnc_image_generator.BNC_y[5]$_DFF_P__93  (.L_HI(net93));
 sg13g2_tiehi \bnc_image_generator.BNC_y[6]$_DFF_P__94  (.L_HI(net94));
 sg13g2_tiehi \bnc_image_generator.counter[0]$_SDFF_PN0__95  (.L_HI(net95));
 sg13g2_tiehi \bnc_image_generator.counter[1]$_SDFF_PN0__96  (.L_HI(net96));
 sg13g2_tiehi \bnc_image_generator.counter[2]$_SDFF_PN0__97  (.L_HI(net97));
 sg13g2_tiehi \bnc_image_generator.counter[3]$_SDFF_PN0__98  (.L_HI(net98));
 sg13g2_tiehi \bnc_image_generator.counter[4]$_SDFF_PN0__99  (.L_HI(net99));
 sg13g2_tiehi \hvsync_gen.hpos[0]$_SDFF_PP0__100  (.L_HI(net100));
 sg13g2_tiehi \hvsync_gen.hpos[1]$_SDFF_PP0__101  (.L_HI(net101));
 sg13g2_tiehi \hvsync_gen.hpos[2]$_SDFF_PP0__102  (.L_HI(net102));
 sg13g2_tiehi \hvsync_gen.hpos[3]$_SDFF_PP0__103  (.L_HI(net103));
 sg13g2_tiehi \hvsync_gen.hpos[4]$_SDFF_PP0__104  (.L_HI(net104));
 sg13g2_tiehi \hvsync_gen.hpos[5]$_SDFF_PP0__105  (.L_HI(net105));
 sg13g2_tiehi \hvsync_gen.hpos[6]$_SDFF_PP0__106  (.L_HI(net106));
 sg13g2_tiehi \hvsync_gen.hpos[7]$_SDFF_PP0__107  (.L_HI(net107));
 sg13g2_tiehi \hvsync_gen.hpos[8]$_SDFF_PP0__108  (.L_HI(net108));
 sg13g2_tiehi \hvsync_gen.hpos[9]$_SDFF_PP0__109  (.L_HI(net109));
 sg13g2_tiehi \hvsync_gen.hsync$_DFF_P__110  (.L_HI(net110));
 sg13g2_tiehi \hvsync_gen.vpos[0]$_SDFFCE_PP0P__111  (.L_HI(net111));
 sg13g2_tiehi \hvsync_gen.vpos[1]$_SDFFCE_PP0P__112  (.L_HI(net112));
 sg13g2_tiehi \hvsync_gen.vpos[2]$_SDFFCE_PP0P__113  (.L_HI(net113));
 sg13g2_tiehi \hvsync_gen.vpos[3]$_SDFFCE_PP0P__114  (.L_HI(net114));
 sg13g2_tiehi \hvsync_gen.vpos[4]$_SDFFCE_PP0P__115  (.L_HI(net115));
 sg13g2_tiehi \hvsync_gen.vpos[5]$_SDFFCE_PP0P__116  (.L_HI(net116));
 sg13g2_tiehi \hvsync_gen.vpos[6]$_SDFFCE_PP0P__117  (.L_HI(net117));
 sg13g2_tiehi \hvsync_gen.vpos[7]$_SDFFCE_PP0P__118  (.L_HI(net118));
 sg13g2_tiehi \hvsync_gen.vpos[8]$_SDFFCE_PP0P__119  (.L_HI(net119));
 sg13g2_tiehi \hvsync_gen.vpos[9]$_SDFFCE_PP0P__120  (.L_HI(net120));
 sg13g2_tiehi \hvsync_gen.vsync$_DFF_P__121  (.L_HI(net121));
 sg13g2_tiehi \vga_image_generator.character_hold[0]$_SDFFE_PN0N__122  (.L_HI(net122));
 sg13g2_tiehi \vga_image_generator.character_hold[10]$_SDFFE_PN0N__123  (.L_HI(net123));
 sg13g2_tiehi \vga_image_generator.character_hold[11]$_SDFFE_PN0N__124  (.L_HI(net124));
 sg13g2_tiehi \vga_image_generator.character_hold[12]$_SDFFE_PN0N__125  (.L_HI(net125));
 sg13g2_tiehi \vga_image_generator.character_hold[13]$_SDFFE_PN0N__126  (.L_HI(net126));
 sg13g2_tiehi \vga_image_generator.character_hold[14]$_SDFFE_PN0N__127  (.L_HI(net127));
 sg13g2_tiehi \vga_image_generator.character_hold[15]$_SDFFE_PN0N__128  (.L_HI(net128));
 sg13g2_tiehi \vga_image_generator.character_hold[16]$_SDFFE_PN0N__129  (.L_HI(net129));
 sg13g2_tiehi \vga_image_generator.character_hold[17]$_SDFFE_PN0N__130  (.L_HI(net130));
 sg13g2_tiehi \vga_image_generator.character_hold[1]$_SDFFE_PN0N__131  (.L_HI(net131));
 sg13g2_tiehi \vga_image_generator.character_hold[2]$_SDFFE_PN0N__132  (.L_HI(net132));
 sg13g2_tiehi \vga_image_generator.character_hold[3]$_SDFFE_PN0N__133  (.L_HI(net133));
 sg13g2_tiehi \vga_image_generator.character_hold[4]$_SDFFE_PN0N__134  (.L_HI(net134));
 sg13g2_tiehi \vga_image_generator.character_hold[5]$_SDFFE_PN0N__135  (.L_HI(net135));
 sg13g2_tiehi \vga_image_generator.character_hold[6]$_SDFFE_PN0N__136  (.L_HI(net136));
 sg13g2_tiehi \vga_image_generator.character_hold[7]$_SDFFE_PN0N__137  (.L_HI(net137));
 sg13g2_tiehi \vga_image_generator.character_hold[8]$_SDFFE_PN0N__138  (.L_HI(net138));
 sg13g2_tiehi \vga_image_generator.character_hold[9]$_SDFFE_PN0N__139  (.L_HI(net139));
 sg13g2_tiehi \vga_image_generator.counter[0]$_SDFF_PN0__140  (.L_HI(net140));
 sg13g2_tiehi \vga_image_generator.counter[10]$_SDFF_PN0__141  (.L_HI(net141));
 sg13g2_tiehi \vga_image_generator.counter[11]$_SDFF_PN0__142  (.L_HI(net142));
 sg13g2_tiehi \vga_image_generator.counter[12]$_SDFF_PN0__143  (.L_HI(net143));
 sg13g2_tiehi \vga_image_generator.counter[13]$_SDFF_PN0__144  (.L_HI(net144));
 sg13g2_tiehi \vga_image_generator.counter[14]$_SDFF_PN0__145  (.L_HI(net145));
 sg13g2_tiehi \vga_image_generator.counter[15]$_SDFF_PN0__146  (.L_HI(net146));
 sg13g2_tiehi \vga_image_generator.counter[16]$_SDFF_PN0__147  (.L_HI(net147));
 sg13g2_tiehi \vga_image_generator.counter[17]$_SDFF_PN0__148  (.L_HI(net148));
 sg13g2_tiehi \vga_image_generator.counter[18]$_SDFF_PN0__149  (.L_HI(net149));
 sg13g2_tiehi \vga_image_generator.counter[19]$_SDFF_PN0__150  (.L_HI(net150));
 sg13g2_tiehi \vga_image_generator.counter[1]$_SDFF_PN0__151  (.L_HI(net151));
 sg13g2_tiehi \vga_image_generator.counter[20]$_SDFF_PN0__152  (.L_HI(net152));
 sg13g2_tiehi \vga_image_generator.counter[21]$_SDFF_PN0__153  (.L_HI(net153));
 sg13g2_tiehi \vga_image_generator.counter[22]$_SDFF_PN0__154  (.L_HI(net154));
 sg13g2_tiehi \vga_image_generator.counter[23]$_SDFF_PN0__155  (.L_HI(net155));
 sg13g2_tiehi \vga_image_generator.counter[24]$_SDFF_PN0__156  (.L_HI(net156));
 sg13g2_tiehi \vga_image_generator.counter[2]$_SDFF_PN0__157  (.L_HI(net157));
 sg13g2_tiehi \vga_image_generator.counter[3]$_SDFF_PN0__158  (.L_HI(net158));
 sg13g2_tiehi \vga_image_generator.counter[4]$_SDFF_PN0__159  (.L_HI(net159));
 sg13g2_tiehi \vga_image_generator.counter[5]$_SDFF_PN0__160  (.L_HI(net160));
 sg13g2_tiehi \vga_image_generator.counter[6]$_SDFF_PN0__161  (.L_HI(net161));
 sg13g2_tiehi \vga_image_generator.counter[7]$_SDFF_PN0__162  (.L_HI(net162));
 sg13g2_tiehi \vga_image_generator.counter[8]$_SDFF_PN0__163  (.L_HI(net163));
 sg13g2_tiehi \vga_image_generator.counter[9]$_SDFF_PN0__164  (.L_HI(net164));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_fill_2 FILLER_9_112 ();
 sg13g2_fill_1 FILLER_9_114 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_140 ();
 sg13g2_fill_1 FILLER_9_146 ();
 sg13g2_decap_8 FILLER_9_159 ();
 sg13g2_decap_8 FILLER_9_166 ();
 sg13g2_decap_8 FILLER_9_173 ();
 sg13g2_decap_8 FILLER_9_180 ();
 sg13g2_decap_8 FILLER_9_190 ();
 sg13g2_decap_8 FILLER_9_197 ();
 sg13g2_decap_8 FILLER_9_204 ();
 sg13g2_decap_8 FILLER_9_211 ();
 sg13g2_decap_8 FILLER_9_218 ();
 sg13g2_decap_8 FILLER_9_225 ();
 sg13g2_decap_4 FILLER_9_232 ();
 sg13g2_fill_2 FILLER_9_236 ();
 sg13g2_decap_8 FILLER_9_242 ();
 sg13g2_decap_8 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_256 ();
 sg13g2_decap_8 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_decap_8 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_284 ();
 sg13g2_decap_8 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_decap_8 FILLER_9_312 ();
 sg13g2_decap_8 FILLER_9_319 ();
 sg13g2_decap_8 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_340 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_9_410 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_decap_4 FILLER_9_424 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_fill_2 FILLER_10_105 ();
 sg13g2_fill_1 FILLER_10_107 ();
 sg13g2_fill_2 FILLER_10_134 ();
 sg13g2_fill_1 FILLER_10_136 ();
 sg13g2_fill_2 FILLER_10_141 ();
 sg13g2_fill_2 FILLER_10_229 ();
 sg13g2_decap_8 FILLER_10_262 ();
 sg13g2_decap_8 FILLER_10_269 ();
 sg13g2_decap_8 FILLER_10_276 ();
 sg13g2_decap_8 FILLER_10_283 ();
 sg13g2_decap_8 FILLER_10_290 ();
 sg13g2_decap_8 FILLER_10_297 ();
 sg13g2_fill_2 FILLER_10_304 ();
 sg13g2_decap_8 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_324 ();
 sg13g2_decap_8 FILLER_10_331 ();
 sg13g2_decap_8 FILLER_10_338 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_decap_8 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_10_415 ();
 sg13g2_decap_8 FILLER_10_422 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_fill_2 FILLER_11_84 ();
 sg13g2_fill_1 FILLER_11_86 ();
 sg13g2_fill_2 FILLER_11_91 ();
 sg13g2_fill_1 FILLER_11_93 ();
 sg13g2_decap_8 FILLER_11_120 ();
 sg13g2_fill_2 FILLER_11_127 ();
 sg13g2_decap_4 FILLER_11_137 ();
 sg13g2_fill_1 FILLER_11_153 ();
 sg13g2_decap_4 FILLER_11_159 ();
 sg13g2_decap_8 FILLER_11_171 ();
 sg13g2_decap_4 FILLER_11_178 ();
 sg13g2_decap_4 FILLER_11_186 ();
 sg13g2_fill_1 FILLER_11_190 ();
 sg13g2_fill_2 FILLER_11_208 ();
 sg13g2_fill_1 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_232 ();
 sg13g2_fill_2 FILLER_11_239 ();
 sg13g2_decap_8 FILLER_11_267 ();
 sg13g2_fill_1 FILLER_11_274 ();
 sg13g2_fill_2 FILLER_11_331 ();
 sg13g2_fill_1 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_decap_4 FILLER_11_345 ();
 sg13g2_fill_1 FILLER_11_349 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_4 FILLER_11_424 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_4 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_60 ();
 sg13g2_fill_2 FILLER_12_92 ();
 sg13g2_fill_1 FILLER_12_94 ();
 sg13g2_decap_8 FILLER_12_107 ();
 sg13g2_decap_8 FILLER_12_114 ();
 sg13g2_decap_8 FILLER_12_121 ();
 sg13g2_fill_1 FILLER_12_171 ();
 sg13g2_decap_8 FILLER_12_176 ();
 sg13g2_decap_8 FILLER_12_183 ();
 sg13g2_fill_2 FILLER_12_190 ();
 sg13g2_fill_1 FILLER_12_192 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_decap_4 FILLER_12_214 ();
 sg13g2_fill_2 FILLER_12_222 ();
 sg13g2_fill_1 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_233 ();
 sg13g2_decap_4 FILLER_12_240 ();
 sg13g2_fill_2 FILLER_12_244 ();
 sg13g2_decap_8 FILLER_12_250 ();
 sg13g2_fill_2 FILLER_12_257 ();
 sg13g2_fill_1 FILLER_12_259 ();
 sg13g2_fill_1 FILLER_12_265 ();
 sg13g2_fill_2 FILLER_12_271 ();
 sg13g2_fill_1 FILLER_12_273 ();
 sg13g2_decap_4 FILLER_12_278 ();
 sg13g2_fill_1 FILLER_12_282 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_4 FILLER_12_294 ();
 sg13g2_fill_1 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_303 ();
 sg13g2_fill_2 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_8 FILLER_12_403 ();
 sg13g2_decap_8 FILLER_12_410 ();
 sg13g2_decap_8 FILLER_12_417 ();
 sg13g2_decap_4 FILLER_12_424 ();
 sg13g2_fill_2 FILLER_12_428 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_4 FILLER_13_63 ();
 sg13g2_fill_2 FILLER_13_67 ();
 sg13g2_decap_8 FILLER_13_73 ();
 sg13g2_fill_2 FILLER_13_95 ();
 sg13g2_decap_8 FILLER_13_101 ();
 sg13g2_fill_2 FILLER_13_108 ();
 sg13g2_fill_1 FILLER_13_110 ();
 sg13g2_fill_1 FILLER_13_115 ();
 sg13g2_decap_4 FILLER_13_122 ();
 sg13g2_decap_4 FILLER_13_138 ();
 sg13g2_fill_1 FILLER_13_142 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_fill_1 FILLER_13_161 ();
 sg13g2_fill_2 FILLER_13_200 ();
 sg13g2_decap_4 FILLER_13_210 ();
 sg13g2_fill_1 FILLER_13_214 ();
 sg13g2_fill_2 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_285 ();
 sg13g2_fill_2 FILLER_13_297 ();
 sg13g2_fill_1 FILLER_13_299 ();
 sg13g2_decap_8 FILLER_13_305 ();
 sg13g2_fill_2 FILLER_13_312 ();
 sg13g2_fill_1 FILLER_13_314 ();
 sg13g2_decap_4 FILLER_13_320 ();
 sg13g2_decap_8 FILLER_13_338 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_8 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_13_412 ();
 sg13g2_decap_8 FILLER_13_419 ();
 sg13g2_decap_4 FILLER_13_426 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_89 ();
 sg13g2_fill_1 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_104 ();
 sg13g2_decap_8 FILLER_14_117 ();
 sg13g2_decap_8 FILLER_14_124 ();
 sg13g2_fill_1 FILLER_14_131 ();
 sg13g2_decap_4 FILLER_14_162 ();
 sg13g2_fill_2 FILLER_14_171 ();
 sg13g2_decap_8 FILLER_14_177 ();
 sg13g2_decap_8 FILLER_14_184 ();
 sg13g2_fill_2 FILLER_14_191 ();
 sg13g2_fill_1 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_199 ();
 sg13g2_fill_1 FILLER_14_206 ();
 sg13g2_fill_2 FILLER_14_212 ();
 sg13g2_decap_4 FILLER_14_232 ();
 sg13g2_decap_4 FILLER_14_241 ();
 sg13g2_fill_1 FILLER_14_245 ();
 sg13g2_decap_4 FILLER_14_250 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_fill_1 FILLER_14_260 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_fill_2 FILLER_14_273 ();
 sg13g2_fill_1 FILLER_14_275 ();
 sg13g2_fill_1 FILLER_14_280 ();
 sg13g2_decap_4 FILLER_14_286 ();
 sg13g2_fill_2 FILLER_14_334 ();
 sg13g2_fill_1 FILLER_14_336 ();
 sg13g2_fill_1 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_8 FILLER_14_404 ();
 sg13g2_decap_8 FILLER_14_411 ();
 sg13g2_decap_8 FILLER_14_418 ();
 sg13g2_decap_4 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_fill_2 FILLER_15_56 ();
 sg13g2_decap_4 FILLER_15_62 ();
 sg13g2_fill_1 FILLER_15_66 ();
 sg13g2_decap_8 FILLER_15_71 ();
 sg13g2_decap_4 FILLER_15_78 ();
 sg13g2_fill_2 FILLER_15_82 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_fill_2 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_139 ();
 sg13g2_decap_8 FILLER_15_146 ();
 sg13g2_decap_8 FILLER_15_153 ();
 sg13g2_fill_1 FILLER_15_160 ();
 sg13g2_fill_2 FILLER_15_169 ();
 sg13g2_fill_1 FILLER_15_201 ();
 sg13g2_decap_8 FILLER_15_206 ();
 sg13g2_fill_1 FILLER_15_218 ();
 sg13g2_fill_1 FILLER_15_224 ();
 sg13g2_fill_2 FILLER_15_230 ();
 sg13g2_fill_2 FILLER_15_258 ();
 sg13g2_fill_2 FILLER_15_295 ();
 sg13g2_fill_2 FILLER_15_302 ();
 sg13g2_fill_1 FILLER_15_308 ();
 sg13g2_fill_2 FILLER_15_313 ();
 sg13g2_fill_2 FILLER_15_319 ();
 sg13g2_fill_1 FILLER_15_321 ();
 sg13g2_fill_1 FILLER_15_326 ();
 sg13g2_fill_2 FILLER_15_367 ();
 sg13g2_fill_1 FILLER_15_369 ();
 sg13g2_decap_4 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_404 ();
 sg13g2_decap_8 FILLER_15_411 ();
 sg13g2_decap_8 FILLER_15_418 ();
 sg13g2_decap_4 FILLER_15_425 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_fill_2 FILLER_16_49 ();
 sg13g2_fill_2 FILLER_16_77 ();
 sg13g2_fill_1 FILLER_16_79 ();
 sg13g2_fill_2 FILLER_16_84 ();
 sg13g2_fill_1 FILLER_16_86 ();
 sg13g2_fill_2 FILLER_16_117 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_161 ();
 sg13g2_fill_1 FILLER_16_163 ();
 sg13g2_decap_8 FILLER_16_169 ();
 sg13g2_decap_4 FILLER_16_176 ();
 sg13g2_fill_2 FILLER_16_180 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_fill_1 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_243 ();
 sg13g2_fill_1 FILLER_16_255 ();
 sg13g2_fill_1 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_272 ();
 sg13g2_fill_2 FILLER_16_279 ();
 sg13g2_fill_1 FILLER_16_281 ();
 sg13g2_fill_2 FILLER_16_312 ();
 sg13g2_fill_1 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_decap_8 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_4 FILLER_16_372 ();
 sg13g2_fill_1 FILLER_16_376 ();
 sg13g2_fill_2 FILLER_16_381 ();
 sg13g2_fill_1 FILLER_16_383 ();
 sg13g2_fill_2 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_4 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_16_410 ();
 sg13g2_decap_8 FILLER_16_417 ();
 sg13g2_decap_4 FILLER_16_424 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_fill_2 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_76 ();
 sg13g2_decap_4 FILLER_17_83 ();
 sg13g2_fill_2 FILLER_17_87 ();
 sg13g2_fill_2 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_111 ();
 sg13g2_decap_8 FILLER_17_118 ();
 sg13g2_fill_1 FILLER_17_125 ();
 sg13g2_decap_4 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_134 ();
 sg13g2_decap_8 FILLER_17_166 ();
 sg13g2_decap_8 FILLER_17_173 ();
 sg13g2_fill_1 FILLER_17_180 ();
 sg13g2_decap_8 FILLER_17_185 ();
 sg13g2_fill_2 FILLER_17_192 ();
 sg13g2_decap_8 FILLER_17_198 ();
 sg13g2_decap_4 FILLER_17_205 ();
 sg13g2_fill_2 FILLER_17_209 ();
 sg13g2_fill_1 FILLER_17_215 ();
 sg13g2_fill_2 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_254 ();
 sg13g2_decap_8 FILLER_17_281 ();
 sg13g2_fill_2 FILLER_17_288 ();
 sg13g2_fill_1 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_295 ();
 sg13g2_decap_8 FILLER_17_302 ();
 sg13g2_fill_2 FILLER_17_309 ();
 sg13g2_fill_1 FILLER_17_311 ();
 sg13g2_fill_1 FILLER_17_320 ();
 sg13g2_decap_4 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_4 FILLER_17_395 ();
 sg13g2_decap_4 FILLER_17_425 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_fill_2 FILLER_18_63 ();
 sg13g2_fill_2 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_93 ();
 sg13g2_fill_1 FILLER_18_99 ();
 sg13g2_fill_2 FILLER_18_126 ();
 sg13g2_decap_4 FILLER_18_132 ();
 sg13g2_decap_8 FILLER_18_160 ();
 sg13g2_fill_2 FILLER_18_167 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_fill_2 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_fill_1 FILLER_18_217 ();
 sg13g2_fill_1 FILLER_18_223 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_fill_1 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_fill_1 FILLER_18_262 ();
 sg13g2_decap_8 FILLER_18_271 ();
 sg13g2_decap_4 FILLER_18_278 ();
 sg13g2_decap_8 FILLER_18_295 ();
 sg13g2_fill_2 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_309 ();
 sg13g2_fill_2 FILLER_18_314 ();
 sg13g2_fill_1 FILLER_18_316 ();
 sg13g2_decap_4 FILLER_18_322 ();
 sg13g2_fill_2 FILLER_18_350 ();
 sg13g2_fill_2 FILLER_18_361 ();
 sg13g2_fill_1 FILLER_18_363 ();
 sg13g2_fill_2 FILLER_18_372 ();
 sg13g2_fill_1 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_379 ();
 sg13g2_decap_4 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_4 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_405 ();
 sg13g2_fill_2 FILLER_18_410 ();
 sg13g2_fill_1 FILLER_18_412 ();
 sg13g2_decap_8 FILLER_18_418 ();
 sg13g2_decap_4 FILLER_18_425 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_fill_1 FILLER_19_84 ();
 sg13g2_fill_1 FILLER_19_102 ();
 sg13g2_decap_4 FILLER_19_111 ();
 sg13g2_fill_2 FILLER_19_115 ();
 sg13g2_fill_2 FILLER_19_160 ();
 sg13g2_fill_1 FILLER_19_188 ();
 sg13g2_decap_4 FILLER_19_193 ();
 sg13g2_fill_2 FILLER_19_197 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_4 FILLER_19_231 ();
 sg13g2_fill_1 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_241 ();
 sg13g2_fill_2 FILLER_19_247 ();
 sg13g2_fill_2 FILLER_19_258 ();
 sg13g2_fill_2 FILLER_19_279 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_fill_2 FILLER_19_317 ();
 sg13g2_decap_4 FILLER_19_337 ();
 sg13g2_fill_1 FILLER_19_341 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_356 ();
 sg13g2_fill_1 FILLER_19_361 ();
 sg13g2_fill_1 FILLER_19_372 ();
 sg13g2_fill_2 FILLER_19_393 ();
 sg13g2_decap_4 FILLER_19_425 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_110 ();
 sg13g2_decap_8 FILLER_20_117 ();
 sg13g2_decap_4 FILLER_20_124 ();
 sg13g2_fill_1 FILLER_20_128 ();
 sg13g2_decap_4 FILLER_20_150 ();
 sg13g2_decap_8 FILLER_20_162 ();
 sg13g2_decap_8 FILLER_20_173 ();
 sg13g2_decap_4 FILLER_20_185 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_216 ();
 sg13g2_decap_8 FILLER_20_223 ();
 sg13g2_decap_8 FILLER_20_230 ();
 sg13g2_decap_4 FILLER_20_237 ();
 sg13g2_fill_1 FILLER_20_241 ();
 sg13g2_fill_2 FILLER_20_251 ();
 sg13g2_fill_2 FILLER_20_257 ();
 sg13g2_fill_1 FILLER_20_259 ();
 sg13g2_fill_2 FILLER_20_299 ();
 sg13g2_decap_4 FILLER_20_307 ();
 sg13g2_fill_2 FILLER_20_315 ();
 sg13g2_fill_1 FILLER_20_317 ();
 sg13g2_fill_1 FILLER_20_323 ();
 sg13g2_decap_8 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_fill_2 FILLER_20_372 ();
 sg13g2_fill_1 FILLER_20_374 ();
 sg13g2_fill_2 FILLER_20_393 ();
 sg13g2_fill_1 FILLER_20_395 ();
 sg13g2_fill_2 FILLER_20_401 ();
 sg13g2_decap_4 FILLER_20_408 ();
 sg13g2_fill_1 FILLER_20_412 ();
 sg13g2_decap_8 FILLER_20_417 ();
 sg13g2_decap_4 FILLER_20_424 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_4 FILLER_21_77 ();
 sg13g2_fill_2 FILLER_21_81 ();
 sg13g2_decap_8 FILLER_21_95 ();
 sg13g2_decap_4 FILLER_21_102 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_fill_1 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_155 ();
 sg13g2_decap_8 FILLER_21_162 ();
 sg13g2_decap_8 FILLER_21_169 ();
 sg13g2_decap_8 FILLER_21_176 ();
 sg13g2_decap_8 FILLER_21_183 ();
 sg13g2_decap_8 FILLER_21_190 ();
 sg13g2_decap_4 FILLER_21_197 ();
 sg13g2_fill_2 FILLER_21_201 ();
 sg13g2_fill_2 FILLER_21_208 ();
 sg13g2_decap_8 FILLER_21_219 ();
 sg13g2_decap_8 FILLER_21_226 ();
 sg13g2_fill_1 FILLER_21_242 ();
 sg13g2_fill_1 FILLER_21_258 ();
 sg13g2_decap_4 FILLER_21_264 ();
 sg13g2_decap_4 FILLER_21_278 ();
 sg13g2_fill_1 FILLER_21_282 ();
 sg13g2_decap_4 FILLER_21_293 ();
 sg13g2_fill_1 FILLER_21_347 ();
 sg13g2_fill_2 FILLER_21_352 ();
 sg13g2_fill_1 FILLER_21_354 ();
 sg13g2_fill_1 FILLER_21_361 ();
 sg13g2_fill_1 FILLER_21_367 ();
 sg13g2_fill_1 FILLER_21_379 ();
 sg13g2_decap_4 FILLER_21_384 ();
 sg13g2_fill_2 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_fill_1 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_21_411 ();
 sg13g2_decap_8 FILLER_21_418 ();
 sg13g2_decap_4 FILLER_21_425 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_4 FILLER_22_56 ();
 sg13g2_fill_1 FILLER_22_86 ();
 sg13g2_fill_1 FILLER_22_91 ();
 sg13g2_fill_1 FILLER_22_96 ();
 sg13g2_fill_2 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_115 ();
 sg13g2_fill_2 FILLER_22_122 ();
 sg13g2_fill_1 FILLER_22_124 ();
 sg13g2_decap_8 FILLER_22_129 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_4 FILLER_22_147 ();
 sg13g2_fill_1 FILLER_22_155 ();
 sg13g2_fill_1 FILLER_22_182 ();
 sg13g2_fill_2 FILLER_22_196 ();
 sg13g2_fill_2 FILLER_22_203 ();
 sg13g2_fill_1 FILLER_22_205 ();
 sg13g2_fill_2 FILLER_22_223 ();
 sg13g2_fill_1 FILLER_22_225 ();
 sg13g2_fill_1 FILLER_22_230 ();
 sg13g2_fill_2 FILLER_22_236 ();
 sg13g2_fill_1 FILLER_22_238 ();
 sg13g2_fill_2 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_decap_8 FILLER_22_255 ();
 sg13g2_fill_2 FILLER_22_262 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_269 ();
 sg13g2_fill_1 FILLER_22_276 ();
 sg13g2_fill_1 FILLER_22_282 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_307 ();
 sg13g2_decap_8 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_321 ();
 sg13g2_fill_1 FILLER_22_332 ();
 sg13g2_fill_1 FILLER_22_343 ();
 sg13g2_decap_4 FILLER_22_357 ();
 sg13g2_decap_4 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_2 FILLER_22_413 ();
 sg13g2_fill_1 FILLER_22_415 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_fill_2 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_65 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_4 FILLER_23_84 ();
 sg13g2_fill_2 FILLER_23_88 ();
 sg13g2_decap_4 FILLER_23_94 ();
 sg13g2_decap_8 FILLER_23_144 ();
 sg13g2_decap_8 FILLER_23_151 ();
 sg13g2_decap_8 FILLER_23_158 ();
 sg13g2_fill_1 FILLER_23_165 ();
 sg13g2_decap_8 FILLER_23_178 ();
 sg13g2_decap_8 FILLER_23_185 ();
 sg13g2_decap_4 FILLER_23_192 ();
 sg13g2_fill_1 FILLER_23_196 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_fill_1 FILLER_23_236 ();
 sg13g2_fill_1 FILLER_23_247 ();
 sg13g2_fill_2 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_278 ();
 sg13g2_decap_4 FILLER_23_284 ();
 sg13g2_fill_2 FILLER_23_288 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_304 ();
 sg13g2_fill_2 FILLER_23_311 ();
 sg13g2_fill_1 FILLER_23_313 ();
 sg13g2_fill_1 FILLER_23_334 ();
 sg13g2_fill_2 FILLER_23_346 ();
 sg13g2_fill_1 FILLER_23_352 ();
 sg13g2_fill_2 FILLER_23_359 ();
 sg13g2_fill_1 FILLER_23_366 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_fill_1 FILLER_23_401 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_4 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_88 ();
 sg13g2_decap_8 FILLER_24_115 ();
 sg13g2_fill_2 FILLER_24_122 ();
 sg13g2_fill_1 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_160 ();
 sg13g2_fill_2 FILLER_24_167 ();
 sg13g2_fill_1 FILLER_24_169 ();
 sg13g2_decap_4 FILLER_24_179 ();
 sg13g2_fill_2 FILLER_24_183 ();
 sg13g2_fill_1 FILLER_24_194 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_213 ();
 sg13g2_fill_2 FILLER_24_218 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_fill_2 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_254 ();
 sg13g2_fill_1 FILLER_24_266 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_decap_4 FILLER_24_309 ();
 sg13g2_fill_1 FILLER_24_313 ();
 sg13g2_fill_1 FILLER_24_320 ();
 sg13g2_fill_1 FILLER_24_326 ();
 sg13g2_fill_1 FILLER_24_332 ();
 sg13g2_fill_2 FILLER_24_343 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_350 ();
 sg13g2_fill_1 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_363 ();
 sg13g2_fill_2 FILLER_24_369 ();
 sg13g2_fill_2 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_fill_1 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_412 ();
 sg13g2_decap_8 FILLER_24_419 ();
 sg13g2_decap_4 FILLER_24_426 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_48 ();
 sg13g2_decap_8 FILLER_25_55 ();
 sg13g2_decap_8 FILLER_25_62 ();
 sg13g2_decap_8 FILLER_25_69 ();
 sg13g2_decap_8 FILLER_25_76 ();
 sg13g2_decap_8 FILLER_25_83 ();
 sg13g2_decap_4 FILLER_25_90 ();
 sg13g2_fill_1 FILLER_25_94 ();
 sg13g2_decap_8 FILLER_25_99 ();
 sg13g2_decap_8 FILLER_25_106 ();
 sg13g2_decap_8 FILLER_25_113 ();
 sg13g2_decap_8 FILLER_25_120 ();
 sg13g2_decap_8 FILLER_25_127 ();
 sg13g2_decap_4 FILLER_25_134 ();
 sg13g2_fill_1 FILLER_25_138 ();
 sg13g2_decap_8 FILLER_25_143 ();
 sg13g2_decap_8 FILLER_25_150 ();
 sg13g2_decap_4 FILLER_25_157 ();
 sg13g2_fill_1 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_193 ();
 sg13g2_fill_2 FILLER_25_210 ();
 sg13g2_fill_1 FILLER_25_212 ();
 sg13g2_fill_1 FILLER_25_229 ();
 sg13g2_fill_2 FILLER_25_243 ();
 sg13g2_fill_1 FILLER_25_245 ();
 sg13g2_fill_2 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_264 ();
 sg13g2_fill_2 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_281 ();
 sg13g2_decap_4 FILLER_25_288 ();
 sg13g2_fill_1 FILLER_25_292 ();
 sg13g2_fill_1 FILLER_25_298 ();
 sg13g2_decap_4 FILLER_25_310 ();
 sg13g2_fill_2 FILLER_25_322 ();
 sg13g2_decap_4 FILLER_25_330 ();
 sg13g2_fill_2 FILLER_25_334 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_4 FILLER_25_377 ();
 sg13g2_fill_1 FILLER_25_381 ();
 sg13g2_fill_1 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_fill_2 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_427 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_68 ();
 sg13g2_decap_4 FILLER_26_75 ();
 sg13g2_fill_2 FILLER_26_79 ();
 sg13g2_decap_8 FILLER_26_111 ();
 sg13g2_fill_1 FILLER_26_118 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_128 ();
 sg13g2_decap_8 FILLER_26_135 ();
 sg13g2_decap_8 FILLER_26_142 ();
 sg13g2_fill_2 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_decap_8 FILLER_26_156 ();
 sg13g2_decap_8 FILLER_26_163 ();
 sg13g2_fill_2 FILLER_26_170 ();
 sg13g2_decap_4 FILLER_26_180 ();
 sg13g2_fill_1 FILLER_26_192 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_fill_1 FILLER_26_206 ();
 sg13g2_fill_2 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_265 ();
 sg13g2_decap_8 FILLER_26_272 ();
 sg13g2_decap_4 FILLER_26_279 ();
 sg13g2_decap_4 FILLER_26_310 ();
 sg13g2_fill_2 FILLER_26_314 ();
 sg13g2_fill_2 FILLER_26_372 ();
 sg13g2_fill_2 FILLER_26_379 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_fill_1 FILLER_26_401 ();
 sg13g2_decap_8 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_26_414 ();
 sg13g2_decap_8 FILLER_26_419 ();
 sg13g2_decap_4 FILLER_26_426 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_37 ();
 sg13g2_decap_8 FILLER_27_68 ();
 sg13g2_fill_2 FILLER_27_75 ();
 sg13g2_fill_2 FILLER_27_82 ();
 sg13g2_fill_1 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_97 ();
 sg13g2_decap_4 FILLER_27_108 ();
 sg13g2_decap_8 FILLER_27_138 ();
 sg13g2_decap_4 FILLER_27_145 ();
 sg13g2_fill_1 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_185 ();
 sg13g2_decap_4 FILLER_27_192 ();
 sg13g2_fill_1 FILLER_27_196 ();
 sg13g2_fill_2 FILLER_27_201 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_2 FILLER_27_225 ();
 sg13g2_fill_2 FILLER_27_237 ();
 sg13g2_fill_1 FILLER_27_239 ();
 sg13g2_fill_2 FILLER_27_251 ();
 sg13g2_fill_2 FILLER_27_268 ();
 sg13g2_fill_1 FILLER_27_274 ();
 sg13g2_decap_4 FILLER_27_280 ();
 sg13g2_fill_1 FILLER_27_294 ();
 sg13g2_fill_2 FILLER_27_317 ();
 sg13g2_fill_1 FILLER_27_319 ();
 sg13g2_decap_4 FILLER_27_325 ();
 sg13g2_fill_1 FILLER_27_329 ();
 sg13g2_fill_2 FILLER_27_335 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_fill_2 FILLER_27_347 ();
 sg13g2_fill_1 FILLER_27_354 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_fill_2 FILLER_27_378 ();
 sg13g2_fill_1 FILLER_27_384 ();
 sg13g2_fill_1 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_414 ();
 sg13g2_decap_8 FILLER_27_421 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_4 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_32 ();
 sg13g2_fill_2 FILLER_28_46 ();
 sg13g2_fill_1 FILLER_28_48 ();
 sg13g2_fill_2 FILLER_28_53 ();
 sg13g2_fill_1 FILLER_28_55 ();
 sg13g2_fill_1 FILLER_28_60 ();
 sg13g2_fill_1 FILLER_28_66 ();
 sg13g2_fill_2 FILLER_28_75 ();
 sg13g2_fill_1 FILLER_28_82 ();
 sg13g2_fill_1 FILLER_28_107 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_decap_4 FILLER_28_118 ();
 sg13g2_fill_1 FILLER_28_122 ();
 sg13g2_fill_2 FILLER_28_128 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_fill_1 FILLER_28_139 ();
 sg13g2_decap_8 FILLER_28_166 ();
 sg13g2_decap_8 FILLER_28_173 ();
 sg13g2_decap_8 FILLER_28_180 ();
 sg13g2_fill_2 FILLER_28_187 ();
 sg13g2_fill_1 FILLER_28_189 ();
 sg13g2_decap_4 FILLER_28_199 ();
 sg13g2_fill_2 FILLER_28_203 ();
 sg13g2_fill_2 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_224 ();
 sg13g2_fill_1 FILLER_28_240 ();
 sg13g2_decap_4 FILLER_28_255 ();
 sg13g2_fill_2 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_4 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_4 FILLER_28_301 ();
 sg13g2_fill_2 FILLER_28_318 ();
 sg13g2_fill_1 FILLER_28_320 ();
 sg13g2_fill_2 FILLER_28_379 ();
 sg13g2_decap_4 FILLER_28_390 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_420 ();
 sg13g2_fill_2 FILLER_28_427 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_30 ();
 sg13g2_fill_1 FILLER_29_36 ();
 sg13g2_fill_2 FILLER_29_54 ();
 sg13g2_fill_2 FILLER_29_61 ();
 sg13g2_fill_1 FILLER_29_72 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_fill_1 FILLER_29_99 ();
 sg13g2_fill_1 FILLER_29_104 ();
 sg13g2_fill_2 FILLER_29_110 ();
 sg13g2_fill_2 FILLER_29_125 ();
 sg13g2_fill_1 FILLER_29_127 ();
 sg13g2_fill_1 FILLER_29_132 ();
 sg13g2_fill_2 FILLER_29_146 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_fill_1 FILLER_29_156 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_fill_2 FILLER_29_168 ();
 sg13g2_fill_1 FILLER_29_170 ();
 sg13g2_fill_2 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_178 ();
 sg13g2_fill_2 FILLER_29_183 ();
 sg13g2_fill_1 FILLER_29_221 ();
 sg13g2_decap_4 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_232 ();
 sg13g2_decap_8 FILLER_29_243 ();
 sg13g2_fill_1 FILLER_29_255 ();
 sg13g2_decap_8 FILLER_29_260 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_decap_8 FILLER_29_292 ();
 sg13g2_fill_1 FILLER_29_299 ();
 sg13g2_decap_8 FILLER_29_305 ();
 sg13g2_decap_8 FILLER_29_312 ();
 sg13g2_decap_4 FILLER_29_319 ();
 sg13g2_fill_1 FILLER_29_343 ();
 sg13g2_fill_1 FILLER_29_351 ();
 sg13g2_fill_2 FILLER_29_378 ();
 sg13g2_fill_1 FILLER_29_380 ();
 sg13g2_fill_1 FILLER_29_387 ();
 sg13g2_fill_1 FILLER_29_392 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_fill_2 FILLER_29_427 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_41 ();
 sg13g2_fill_1 FILLER_30_46 ();
 sg13g2_fill_2 FILLER_30_52 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_fill_1 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_139 ();
 sg13g2_fill_2 FILLER_30_149 ();
 sg13g2_fill_1 FILLER_30_155 ();
 sg13g2_decap_8 FILLER_30_185 ();
 sg13g2_decap_8 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_199 ();
 sg13g2_decap_8 FILLER_30_206 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_decap_8 FILLER_30_220 ();
 sg13g2_decap_8 FILLER_30_227 ();
 sg13g2_decap_8 FILLER_30_244 ();
 sg13g2_decap_4 FILLER_30_251 ();
 sg13g2_decap_4 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_273 ();
 sg13g2_fill_2 FILLER_30_279 ();
 sg13g2_decap_4 FILLER_30_288 ();
 sg13g2_fill_2 FILLER_30_297 ();
 sg13g2_fill_2 FILLER_30_304 ();
 sg13g2_fill_2 FILLER_30_311 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_fill_2 FILLER_30_320 ();
 sg13g2_fill_1 FILLER_30_322 ();
 sg13g2_fill_2 FILLER_30_326 ();
 sg13g2_fill_1 FILLER_30_340 ();
 sg13g2_fill_1 FILLER_30_351 ();
 sg13g2_fill_2 FILLER_30_368 ();
 sg13g2_fill_1 FILLER_30_370 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_fill_1 FILLER_30_390 ();
 sg13g2_fill_1 FILLER_30_396 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_decap_4 FILLER_30_408 ();
 sg13g2_fill_1 FILLER_30_412 ();
 sg13g2_decap_8 FILLER_30_417 ();
 sg13g2_decap_4 FILLER_30_424 ();
 sg13g2_fill_2 FILLER_30_428 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_28 ();
 sg13g2_fill_1 FILLER_31_30 ();
 sg13g2_fill_1 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_64 ();
 sg13g2_fill_1 FILLER_31_77 ();
 sg13g2_fill_2 FILLER_31_87 ();
 sg13g2_fill_1 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_108 ();
 sg13g2_fill_1 FILLER_31_110 ();
 sg13g2_fill_1 FILLER_31_120 ();
 sg13g2_fill_1 FILLER_31_134 ();
 sg13g2_fill_2 FILLER_31_139 ();
 sg13g2_decap_8 FILLER_31_151 ();
 sg13g2_decap_8 FILLER_31_158 ();
 sg13g2_decap_8 FILLER_31_165 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_251 ();
 sg13g2_decap_8 FILLER_31_258 ();
 sg13g2_decap_8 FILLER_31_265 ();
 sg13g2_fill_2 FILLER_31_272 ();
 sg13g2_fill_1 FILLER_31_274 ();
 sg13g2_fill_2 FILLER_31_280 ();
 sg13g2_fill_2 FILLER_31_287 ();
 sg13g2_fill_1 FILLER_31_328 ();
 sg13g2_decap_4 FILLER_31_333 ();
 sg13g2_fill_2 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_decap_4 FILLER_31_357 ();
 sg13g2_fill_1 FILLER_31_361 ();
 sg13g2_fill_2 FILLER_31_367 ();
 sg13g2_decap_8 FILLER_31_373 ();
 sg13g2_decap_4 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_fill_2 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_403 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_fill_2 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_30 ();
 sg13g2_fill_1 FILLER_32_51 ();
 sg13g2_fill_2 FILLER_32_57 ();
 sg13g2_fill_1 FILLER_32_63 ();
 sg13g2_fill_1 FILLER_32_87 ();
 sg13g2_fill_1 FILLER_32_103 ();
 sg13g2_fill_1 FILLER_32_110 ();
 sg13g2_fill_1 FILLER_32_115 ();
 sg13g2_fill_2 FILLER_32_120 ();
 sg13g2_fill_2 FILLER_32_127 ();
 sg13g2_fill_2 FILLER_32_134 ();
 sg13g2_decap_4 FILLER_32_146 ();
 sg13g2_fill_2 FILLER_32_150 ();
 sg13g2_decap_8 FILLER_32_156 ();
 sg13g2_decap_8 FILLER_32_167 ();
 sg13g2_fill_2 FILLER_32_174 ();
 sg13g2_fill_1 FILLER_32_176 ();
 sg13g2_decap_8 FILLER_32_181 ();
 sg13g2_decap_8 FILLER_32_188 ();
 sg13g2_decap_8 FILLER_32_195 ();
 sg13g2_fill_2 FILLER_32_202 ();
 sg13g2_fill_1 FILLER_32_204 ();
 sg13g2_decap_4 FILLER_32_209 ();
 sg13g2_fill_2 FILLER_32_213 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_238 ();
 sg13g2_fill_1 FILLER_32_240 ();
 sg13g2_fill_1 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_254 ();
 sg13g2_decap_8 FILLER_32_261 ();
 sg13g2_decap_4 FILLER_32_268 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_fill_1 FILLER_32_277 ();
 sg13g2_fill_2 FILLER_32_289 ();
 sg13g2_fill_1 FILLER_32_291 ();
 sg13g2_decap_8 FILLER_32_297 ();
 sg13g2_fill_1 FILLER_32_304 ();
 sg13g2_decap_8 FILLER_32_311 ();
 sg13g2_fill_1 FILLER_32_318 ();
 sg13g2_decap_4 FILLER_32_346 ();
 sg13g2_decap_4 FILLER_32_383 ();
 sg13g2_fill_1 FILLER_32_387 ();
 sg13g2_fill_2 FILLER_32_427 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_4 FILLER_33_21 ();
 sg13g2_fill_2 FILLER_33_25 ();
 sg13g2_decap_4 FILLER_33_52 ();
 sg13g2_fill_1 FILLER_33_60 ();
 sg13g2_decap_8 FILLER_33_71 ();
 sg13g2_decap_8 FILLER_33_78 ();
 sg13g2_fill_2 FILLER_33_85 ();
 sg13g2_fill_2 FILLER_33_91 ();
 sg13g2_fill_1 FILLER_33_93 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_fill_2 FILLER_33_119 ();
 sg13g2_decap_4 FILLER_33_125 ();
 sg13g2_fill_1 FILLER_33_142 ();
 sg13g2_decap_8 FILLER_33_234 ();
 sg13g2_fill_2 FILLER_33_241 ();
 sg13g2_fill_1 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_256 ();
 sg13g2_fill_1 FILLER_33_279 ();
 sg13g2_decap_4 FILLER_33_285 ();
 sg13g2_fill_1 FILLER_33_289 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_303 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_fill_1 FILLER_33_318 ();
 sg13g2_fill_2 FILLER_33_329 ();
 sg13g2_fill_1 FILLER_33_342 ();
 sg13g2_fill_2 FILLER_33_350 ();
 sg13g2_fill_2 FILLER_33_357 ();
 sg13g2_fill_1 FILLER_33_359 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_fill_1 FILLER_33_367 ();
 sg13g2_fill_1 FILLER_33_399 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_decap_8 FILLER_33_412 ();
 sg13g2_decap_8 FILLER_33_419 ();
 sg13g2_decap_4 FILLER_33_426 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_25 ();
 sg13g2_fill_1 FILLER_34_41 ();
 sg13g2_fill_1 FILLER_34_47 ();
 sg13g2_fill_2 FILLER_34_53 ();
 sg13g2_fill_2 FILLER_34_61 ();
 sg13g2_fill_2 FILLER_34_68 ();
 sg13g2_fill_1 FILLER_34_76 ();
 sg13g2_fill_1 FILLER_34_82 ();
 sg13g2_fill_1 FILLER_34_88 ();
 sg13g2_fill_1 FILLER_34_99 ();
 sg13g2_fill_1 FILLER_34_112 ();
 sg13g2_fill_2 FILLER_34_127 ();
 sg13g2_fill_1 FILLER_34_129 ();
 sg13g2_decap_8 FILLER_34_144 ();
 sg13g2_fill_1 FILLER_34_154 ();
 sg13g2_fill_2 FILLER_34_181 ();
 sg13g2_decap_8 FILLER_34_209 ();
 sg13g2_decap_4 FILLER_34_242 ();
 sg13g2_fill_1 FILLER_34_246 ();
 sg13g2_decap_8 FILLER_34_256 ();
 sg13g2_decap_8 FILLER_34_263 ();
 sg13g2_decap_4 FILLER_34_270 ();
 sg13g2_fill_1 FILLER_34_274 ();
 sg13g2_decap_8 FILLER_34_279 ();
 sg13g2_fill_1 FILLER_34_286 ();
 sg13g2_decap_4 FILLER_34_306 ();
 sg13g2_fill_1 FILLER_34_310 ();
 sg13g2_decap_8 FILLER_34_328 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_fill_1 FILLER_34_341 ();
 sg13g2_fill_1 FILLER_34_346 ();
 sg13g2_decap_4 FILLER_34_351 ();
 sg13g2_fill_2 FILLER_34_355 ();
 sg13g2_decap_4 FILLER_34_375 ();
 sg13g2_fill_1 FILLER_34_379 ();
 sg13g2_decap_8 FILLER_34_410 ();
 sg13g2_decap_8 FILLER_34_417 ();
 sg13g2_decap_4 FILLER_34_424 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_37 ();
 sg13g2_decap_4 FILLER_35_48 ();
 sg13g2_fill_1 FILLER_35_52 ();
 sg13g2_decap_4 FILLER_35_72 ();
 sg13g2_fill_1 FILLER_35_85 ();
 sg13g2_fill_1 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_100 ();
 sg13g2_fill_2 FILLER_35_106 ();
 sg13g2_decap_8 FILLER_35_115 ();
 sg13g2_decap_4 FILLER_35_122 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_135 ();
 sg13g2_fill_2 FILLER_35_142 ();
 sg13g2_fill_2 FILLER_35_170 ();
 sg13g2_fill_2 FILLER_35_176 ();
 sg13g2_fill_1 FILLER_35_178 ();
 sg13g2_fill_1 FILLER_35_189 ();
 sg13g2_fill_2 FILLER_35_194 ();
 sg13g2_fill_1 FILLER_35_196 ();
 sg13g2_decap_4 FILLER_35_201 ();
 sg13g2_fill_2 FILLER_35_205 ();
 sg13g2_decap_4 FILLER_35_217 ();
 sg13g2_fill_2 FILLER_35_221 ();
 sg13g2_fill_1 FILLER_35_227 ();
 sg13g2_fill_2 FILLER_35_238 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_fill_2 FILLER_35_286 ();
 sg13g2_fill_1 FILLER_35_304 ();
 sg13g2_fill_1 FILLER_35_326 ();
 sg13g2_decap_8 FILLER_35_332 ();
 sg13g2_decap_8 FILLER_35_339 ();
 sg13g2_fill_2 FILLER_35_346 ();
 sg13g2_fill_1 FILLER_35_348 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_8 FILLER_35_404 ();
 sg13g2_decap_8 FILLER_35_411 ();
 sg13g2_decap_8 FILLER_35_418 ();
 sg13g2_decap_4 FILLER_35_425 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_fill_2 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_fill_1 FILLER_36_77 ();
 sg13g2_decap_4 FILLER_36_83 ();
 sg13g2_fill_1 FILLER_36_87 ();
 sg13g2_decap_8 FILLER_36_97 ();
 sg13g2_decap_8 FILLER_36_104 ();
 sg13g2_fill_2 FILLER_36_111 ();
 sg13g2_fill_1 FILLER_36_113 ();
 sg13g2_decap_8 FILLER_36_118 ();
 sg13g2_decap_8 FILLER_36_125 ();
 sg13g2_decap_8 FILLER_36_132 ();
 sg13g2_decap_8 FILLER_36_143 ();
 sg13g2_fill_2 FILLER_36_150 ();
 sg13g2_decap_8 FILLER_36_156 ();
 sg13g2_decap_4 FILLER_36_163 ();
 sg13g2_fill_2 FILLER_36_167 ();
 sg13g2_fill_1 FILLER_36_178 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_decap_4 FILLER_36_190 ();
 sg13g2_decap_8 FILLER_36_226 ();
 sg13g2_decap_8 FILLER_36_233 ();
 sg13g2_decap_8 FILLER_36_240 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_fill_2 FILLER_36_252 ();
 sg13g2_fill_2 FILLER_36_259 ();
 sg13g2_decap_4 FILLER_36_264 ();
 sg13g2_fill_2 FILLER_36_268 ();
 sg13g2_decap_8 FILLER_36_274 ();
 sg13g2_decap_8 FILLER_36_281 ();
 sg13g2_decap_8 FILLER_36_288 ();
 sg13g2_fill_2 FILLER_36_295 ();
 sg13g2_fill_2 FILLER_36_302 ();
 sg13g2_fill_1 FILLER_36_304 ();
 sg13g2_fill_2 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_321 ();
 sg13g2_fill_1 FILLER_36_336 ();
 sg13g2_decap_4 FILLER_36_342 ();
 sg13g2_fill_2 FILLER_36_350 ();
 sg13g2_fill_2 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_4 FILLER_36_384 ();
 sg13g2_fill_1 FILLER_36_388 ();
 sg13g2_fill_1 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_36_414 ();
 sg13g2_decap_8 FILLER_36_421 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_fill_1 FILLER_37_46 ();
 sg13g2_decap_4 FILLER_37_51 ();
 sg13g2_fill_1 FILLER_37_164 ();
 sg13g2_decap_8 FILLER_37_188 ();
 sg13g2_decap_4 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_199 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_fill_2 FILLER_37_217 ();
 sg13g2_fill_1 FILLER_37_219 ();
 sg13g2_fill_1 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_248 ();
 sg13g2_fill_2 FILLER_37_255 ();
 sg13g2_decap_4 FILLER_37_262 ();
 sg13g2_fill_2 FILLER_37_266 ();
 sg13g2_fill_2 FILLER_37_320 ();
 sg13g2_fill_2 FILLER_37_332 ();
 sg13g2_fill_2 FILLER_37_338 ();
 sg13g2_fill_2 FILLER_37_344 ();
 sg13g2_fill_1 FILLER_37_346 ();
 sg13g2_decap_4 FILLER_37_352 ();
 sg13g2_fill_2 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_4 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_423 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_61 ();
 sg13g2_decap_4 FILLER_38_67 ();
 sg13g2_fill_2 FILLER_38_176 ();
 sg13g2_fill_1 FILLER_38_178 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_4 FILLER_38_198 ();
 sg13g2_fill_2 FILLER_38_202 ();
 sg13g2_decap_4 FILLER_38_208 ();
 sg13g2_fill_1 FILLER_38_212 ();
 sg13g2_fill_2 FILLER_38_249 ();
 sg13g2_fill_1 FILLER_38_255 ();
 sg13g2_fill_2 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_279 ();
 sg13g2_decap_8 FILLER_38_286 ();
 sg13g2_decap_4 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_304 ();
 sg13g2_decap_4 FILLER_38_315 ();
 sg13g2_fill_2 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_328 ();
 sg13g2_decap_4 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_fill_1 FILLER_38_404 ();
 sg13g2_decap_8 FILLER_38_409 ();
 sg13g2_decap_8 FILLER_38_416 ();
 sg13g2_decap_8 FILLER_38_423 ();
endmodule
