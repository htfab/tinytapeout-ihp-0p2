module tt_um_cfib_demo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire clknet_0_clk;
 wire net83;
 wire hsync;
 wire pwm;
 wire \top_inst.pwm_inst.cntr[0] ;
 wire \top_inst.pwm_inst.cntr[1] ;
 wire \top_inst.pwm_inst.cntr[2] ;
 wire \top_inst.pwm_inst.cntr[3] ;
 wire \top_inst.sample_ena ;
 wire \top_inst.sndgen_inst.bar_counter[0] ;
 wire \top_inst.sndgen_inst.bar_counter[1] ;
 wire \top_inst.sndgen_inst.bar_counter[2] ;
 wire \top_inst.sndgen_inst.bar_counter[3] ;
 wire \top_inst.sndgen_inst.c1[0] ;
 wire \top_inst.sndgen_inst.c1[1] ;
 wire \top_inst.sndgen_inst.c2[0] ;
 wire \top_inst.sndgen_inst.c2[1] ;
 wire \top_inst.sndgen_inst.c2[2] ;
 wire \top_inst.sndgen_inst.c3[0] ;
 wire \top_inst.sndgen_inst.c3[1] ;
 wire \top_inst.sndgen_inst.c3[2] ;
 wire \top_inst.sndgen_inst.c4[2] ;
 wire \top_inst.sndgen_inst.lfsr[0] ;
 wire \top_inst.sndgen_inst.lfsr[1] ;
 wire \top_inst.sndgen_inst.lfsr[2] ;
 wire \top_inst.sndgen_inst.lfsr[3] ;
 wire \top_inst.sndgen_inst.lfsr[4] ;
 wire \top_inst.sndgen_inst.lfsr[5] ;
 wire \top_inst.sndgen_inst.lfsr[6] ;
 wire \top_inst.sndgen_inst.lfsr[7] ;
 wire \top_inst.sndgen_inst.mask_1[0] ;
 wire \top_inst.sndgen_inst.mask_1[1] ;
 wire \top_inst.sndgen_inst.mask_1[2] ;
 wire \top_inst.sndgen_inst.mask_1[3] ;
 wire \top_inst.sndgen_inst.mask_2 ;
 wire \top_inst.sndgen_inst.p_c2[0] ;
 wire \top_inst.sndgen_inst.p_c2[10] ;
 wire \top_inst.sndgen_inst.p_c2[1] ;
 wire \top_inst.sndgen_inst.p_c2[2] ;
 wire \top_inst.sndgen_inst.p_c2[3] ;
 wire \top_inst.sndgen_inst.p_c2[4] ;
 wire \top_inst.sndgen_inst.p_c2[5] ;
 wire \top_inst.sndgen_inst.p_c2[6] ;
 wire \top_inst.sndgen_inst.p_c2[7] ;
 wire \top_inst.sndgen_inst.p_c3[0] ;
 wire \top_inst.sndgen_inst.p_c3[10] ;
 wire \top_inst.sndgen_inst.p_c3[1] ;
 wire \top_inst.sndgen_inst.p_c3[2] ;
 wire \top_inst.sndgen_inst.p_c3[3] ;
 wire \top_inst.sndgen_inst.p_c3[4] ;
 wire \top_inst.sndgen_inst.p_c3[5] ;
 wire \top_inst.sndgen_inst.p_c3[6] ;
 wire \top_inst.sndgen_inst.p_c3[7] ;
 wire \top_inst.sndgen_inst.p_c4[0] ;
 wire \top_inst.sndgen_inst.p_c4[10] ;
 wire \top_inst.sndgen_inst.p_c4[1] ;
 wire \top_inst.sndgen_inst.p_c4[2] ;
 wire \top_inst.sndgen_inst.p_c4[3] ;
 wire \top_inst.sndgen_inst.p_c4[4] ;
 wire \top_inst.sndgen_inst.p_c4[5] ;
 wire \top_inst.sndgen_inst.p_c4[6] ;
 wire \top_inst.sndgen_inst.p_c4[7] ;
 wire \top_inst.sndgen_inst.phacc2[0] ;
 wire \top_inst.sndgen_inst.phacc2[10] ;
 wire \top_inst.sndgen_inst.phacc2[11] ;
 wire \top_inst.sndgen_inst.phacc2[12] ;
 wire \top_inst.sndgen_inst.phacc2[13] ;
 wire \top_inst.sndgen_inst.phacc2[1] ;
 wire \top_inst.sndgen_inst.phacc2[2] ;
 wire \top_inst.sndgen_inst.phacc2[3] ;
 wire \top_inst.sndgen_inst.phacc2[4] ;
 wire \top_inst.sndgen_inst.phacc2[5] ;
 wire \top_inst.sndgen_inst.phacc2[6] ;
 wire \top_inst.sndgen_inst.phacc2[7] ;
 wire \top_inst.sndgen_inst.phacc2[8] ;
 wire \top_inst.sndgen_inst.phacc2[9] ;
 wire \top_inst.sndgen_inst.phacc3[0] ;
 wire \top_inst.sndgen_inst.phacc3[10] ;
 wire \top_inst.sndgen_inst.phacc3[11] ;
 wire \top_inst.sndgen_inst.phacc3[12] ;
 wire \top_inst.sndgen_inst.phacc3[13] ;
 wire \top_inst.sndgen_inst.phacc3[1] ;
 wire \top_inst.sndgen_inst.phacc3[2] ;
 wire \top_inst.sndgen_inst.phacc3[3] ;
 wire \top_inst.sndgen_inst.phacc3[4] ;
 wire \top_inst.sndgen_inst.phacc3[5] ;
 wire \top_inst.sndgen_inst.phacc3[6] ;
 wire \top_inst.sndgen_inst.phacc3[7] ;
 wire \top_inst.sndgen_inst.phacc3[8] ;
 wire \top_inst.sndgen_inst.phacc3[9] ;
 wire \top_inst.sndgen_inst.phacc4[0] ;
 wire \top_inst.sndgen_inst.phacc4[10] ;
 wire \top_inst.sndgen_inst.phacc4[11] ;
 wire \top_inst.sndgen_inst.phacc4[12] ;
 wire \top_inst.sndgen_inst.phacc4[13] ;
 wire \top_inst.sndgen_inst.phacc4[1] ;
 wire \top_inst.sndgen_inst.phacc4[2] ;
 wire \top_inst.sndgen_inst.phacc4[3] ;
 wire \top_inst.sndgen_inst.phacc4[4] ;
 wire \top_inst.sndgen_inst.phacc4[5] ;
 wire \top_inst.sndgen_inst.phacc4[6] ;
 wire \top_inst.sndgen_inst.phacc4[7] ;
 wire \top_inst.sndgen_inst.phacc4[8] ;
 wire \top_inst.sndgen_inst.phacc4[9] ;
 wire \top_inst.sndgen_inst.rom_addr[0] ;
 wire \top_inst.sndgen_inst.rom_addr[1] ;
 wire \top_inst.sndgen_inst.rom_addr[2] ;
 wire \top_inst.sndgen_inst.rom_addr[3] ;
 wire \top_inst.sndgen_inst.sample_ena_delay[0] ;
 wire \top_inst.sndgen_inst.sample_ena_delay[1] ;
 wire \top_inst.sndgen_inst.sample_ena_delay[2] ;
 wire \top_inst.sndgen_inst.slot_counter[0] ;
 wire \top_inst.sndgen_inst.slot_counter[10] ;
 wire \top_inst.sndgen_inst.slot_counter[1] ;
 wire \top_inst.sndgen_inst.slot_counter[2] ;
 wire \top_inst.sndgen_inst.slot_counter[3] ;
 wire \top_inst.sndgen_inst.slot_counter[4] ;
 wire \top_inst.sndgen_inst.slot_counter[5] ;
 wire \top_inst.sndgen_inst.slot_counter[6] ;
 wire \top_inst.sndgen_inst.slot_counter[7] ;
 wire \top_inst.sndgen_inst.slot_counter[8] ;
 wire \top_inst.sndgen_inst.slot_counter[9] ;
 wire \top_inst.sys_presc[0] ;
 wire \top_inst.sys_presc[1] ;
 wire \top_inst.sys_presc[2] ;
 wire \top_inst.sys_presc[3] ;
 wire \top_inst.sys_presc[4] ;
 wire \top_inst.vga_inst.bg[0] ;
 wire \top_inst.vga_inst.bg[1] ;
 wire \top_inst.vga_inst.bg[4] ;
 wire \top_inst.vga_inst.bg[5] ;
 wire \top_inst.vga_inst.sr1[0] ;
 wire \top_inst.vga_inst.sr1[1] ;
 wire \top_inst.vga_inst.sr1[2] ;
 wire \top_inst.vga_inst.sr1[3] ;
 wire \top_inst.vga_inst.sx1[0] ;
 wire \top_inst.vga_inst.sx1[1] ;
 wire \top_inst.vga_inst.sx1[2] ;
 wire \top_inst.vga_inst.sx1[3] ;
 wire \top_inst.vga_inst.vsync ;
 wire \top_inst.vga_inst.x1[0] ;
 wire \top_inst.vga_inst.x1[1] ;
 wire \top_inst.vga_inst.x1[2] ;
 wire \top_inst.vga_inst.x1[3] ;
 wire \top_inst.vga_inst.x1[4] ;
 wire \top_inst.vga_inst.x1[5] ;
 wire \top_inst.vga_inst.x1[6] ;
 wire \top_inst.vga_inst.x1[7] ;
 wire \top_inst.vga_inst.x[0] ;
 wire \top_inst.vga_inst.x[1] ;
 wire \top_inst.vga_inst.x[2] ;
 wire \top_inst.vga_inst.x[3] ;
 wire \top_inst.vga_inst.x[4] ;
 wire \top_inst.vga_inst.x[5] ;
 wire \top_inst.vga_inst.x[6] ;
 wire \top_inst.vga_inst.x[7] ;
 wire \top_inst.vga_inst.x[8] ;
 wire \top_inst.vga_inst.x[9] ;
 wire \top_inst.vga_inst.xmax[0] ;
 wire \top_inst.vga_inst.xmax[1] ;
 wire \top_inst.vga_inst.xmax[2] ;
 wire \top_inst.vga_inst.xmax[3] ;
 wire \top_inst.vga_inst.xmin[0] ;
 wire \top_inst.vga_inst.xmin[1] ;
 wire \top_inst.vga_inst.xmin[2] ;
 wire \top_inst.vga_inst.xmin[3] ;
 wire \top_inst.vga_inst.y[0] ;
 wire \top_inst.vga_inst.y[1] ;
 wire \top_inst.vga_inst.y[2] ;
 wire \top_inst.vga_inst.y[7] ;
 wire \top_inst.vga_inst.y[8] ;
 wire \top_inst.vga_inst.y[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_2 _1055_ (.A(\top_inst.vga_inst.x[6] ),
    .X(_0387_));
 sg13g2_buf_2 _1056_ (.A(\top_inst.vga_inst.x[0] ),
    .X(_0388_));
 sg13g2_nor4_2 _1057_ (.A(\top_inst.vga_inst.x[3] ),
    .B(\top_inst.vga_inst.x[2] ),
    .C(\top_inst.vga_inst.x[1] ),
    .Y(_0389_),
    .D(_0388_));
 sg13g2_buf_2 _1058_ (.A(\top_inst.vga_inst.x[4] ),
    .X(_0390_));
 sg13g2_buf_1 _1059_ (.A(\top_inst.vga_inst.x[5] ),
    .X(_0391_));
 sg13g2_nor2_1 _1060_ (.A(_0390_),
    .B(net38),
    .Y(_0392_));
 sg13g2_nand2_1 _1061_ (.Y(_0393_),
    .A(_0389_),
    .B(_0392_));
 sg13g2_buf_1 _1062_ (.A(\top_inst.vga_inst.x[9] ),
    .X(_0394_));
 sg13g2_buf_2 _1063_ (.A(\top_inst.vga_inst.x[7] ),
    .X(_0395_));
 sg13g2_nand3b_1 _1064_ (.B(net37),
    .C(_0395_),
    .Y(_0396_),
    .A_N(\top_inst.vga_inst.x[8] ));
 sg13g2_buf_1 _1065_ (.A(\top_inst.vga_inst.y[0] ),
    .X(_0397_));
 sg13g2_buf_2 _1066_ (.A(\top_inst.sys_presc[0] ),
    .X(_0398_));
 sg13g2_nand2_1 _1067_ (.Y(_0399_),
    .A(net36),
    .B(_0398_));
 sg13g2_nor4_2 _1068_ (.A(_0387_),
    .B(_0393_),
    .C(_0396_),
    .Y(_0400_),
    .D(_0399_));
 sg13g2_buf_1 _1069_ (.A(_0400_),
    .X(\top_inst.sample_ena ));
 sg13g2_buf_1 _1070_ (.A(_0398_),
    .X(_0401_));
 sg13g2_xor2_1 _1071_ (.B(\top_inst.sys_presc[1] ),
    .A(net27),
    .X(_0014_));
 sg13g2_nand2_1 _1072_ (.Y(_0402_),
    .A(net27),
    .B(\top_inst.sys_presc[1] ));
 sg13g2_xnor2_1 _1073_ (.Y(_0015_),
    .A(\top_inst.sys_presc[2] ),
    .B(_0402_));
 sg13g2_nand3_1 _1074_ (.B(\top_inst.sys_presc[1] ),
    .C(\top_inst.sys_presc[2] ),
    .A(net27),
    .Y(_0403_));
 sg13g2_xnor2_1 _1075_ (.Y(_0016_),
    .A(\top_inst.sys_presc[3] ),
    .B(_0403_));
 sg13g2_nand4_1 _1076_ (.B(\top_inst.sys_presc[1] ),
    .C(\top_inst.sys_presc[3] ),
    .A(net27),
    .Y(_0404_),
    .D(\top_inst.sys_presc[2] ));
 sg13g2_xnor2_1 _1077_ (.Y(_0017_),
    .A(\top_inst.sys_presc[4] ),
    .B(_0404_));
 sg13g2_and3_1 _1078_ (.X(_0405_),
    .A(\top_inst.sndgen_inst.slot_counter[5] ),
    .B(\top_inst.sndgen_inst.slot_counter[4] ),
    .C(\top_inst.sndgen_inst.slot_counter[6] ));
 sg13g2_nand3_1 _1079_ (.B(\top_inst.sndgen_inst.slot_counter[7] ),
    .C(_0405_),
    .A(\top_inst.sndgen_inst.slot_counter[8] ),
    .Y(_0406_));
 sg13g2_nand2_1 _1080_ (.Y(_0407_),
    .A(\top_inst.sndgen_inst.slot_counter[9] ),
    .B(\top_inst.sndgen_inst.slot_counter[10] ));
 sg13g2_inv_1 _1081_ (.Y(_0408_),
    .A(_0407_));
 sg13g2_buf_1 _1082_ (.A(\top_inst.sndgen_inst.slot_counter[1] ),
    .X(_0409_));
 sg13g2_and3_1 _1083_ (.X(_0410_),
    .A(net35),
    .B(\top_inst.sndgen_inst.slot_counter[3] ),
    .C(\top_inst.sndgen_inst.slot_counter[2] ));
 sg13g2_buf_1 _1084_ (.A(_0410_),
    .X(_0411_));
 sg13g2_nand3b_1 _1085_ (.B(_0408_),
    .C(_0411_),
    .Y(_0412_),
    .A_N(_0406_));
 sg13g2_nor2b_1 _1086_ (.A(_0019_),
    .B_N(_0400_),
    .Y(_0413_));
 sg13g2_nand2b_1 _1087_ (.Y(_0414_),
    .B(_0413_),
    .A_N(_0412_));
 sg13g2_buf_1 _1088_ (.A(_0414_),
    .X(_0415_));
 sg13g2_buf_2 _1089_ (.A(\top_inst.sndgen_inst.bar_counter[0] ),
    .X(_0416_));
 sg13g2_buf_2 _1090_ (.A(\top_inst.sndgen_inst.bar_counter[2] ),
    .X(_0417_));
 sg13g2_nand2_1 _1091_ (.Y(_0418_),
    .A(_0416_),
    .B(_0417_));
 sg13g2_buf_2 _1092_ (.A(\top_inst.sndgen_inst.bar_counter[1] ),
    .X(_0419_));
 sg13g2_mux2_1 _1093_ (.A0(_0418_),
    .A1(_0416_),
    .S(_0419_),
    .X(_0420_));
 sg13g2_nand2_1 _1094_ (.Y(_0421_),
    .A(\top_inst.sndgen_inst.c1[0] ),
    .B(net12));
 sg13g2_o21ai_1 _1095_ (.B1(_0421_),
    .Y(_0027_),
    .A1(net12),
    .A2(_0420_));
 sg13g2_inv_1 _1096_ (.Y(_0422_),
    .A(_0020_));
 sg13g2_nor2_1 _1097_ (.A(_0417_),
    .B(_0010_),
    .Y(_0423_));
 sg13g2_nor4_1 _1098_ (.A(_0419_),
    .B(_0416_),
    .C(_0414_),
    .D(_0423_),
    .Y(_0424_));
 sg13g2_a21oi_1 _1099_ (.A1(_0422_),
    .A2(net12),
    .Y(_0028_),
    .B1(_0424_));
 sg13g2_nand2_1 _1100_ (.Y(_0425_),
    .A(_0419_),
    .B(_0416_));
 sg13g2_buf_2 _1101_ (.A(\top_inst.sndgen_inst.slot_counter[0] ),
    .X(_0426_));
 sg13g2_nand3_1 _1102_ (.B(_0400_),
    .C(_0411_),
    .A(_0426_),
    .Y(_0427_));
 sg13g2_nor2_1 _1103_ (.A(_0406_),
    .B(_0427_),
    .Y(_0428_));
 sg13g2_nand2_1 _1104_ (.Y(_0429_),
    .A(\top_inst.sndgen_inst.slot_counter[9] ),
    .B(_0428_));
 sg13g2_or3_1 _1105_ (.A(_0002_),
    .B(_0425_),
    .C(_0429_),
    .X(_0430_));
 sg13g2_buf_1 _1106_ (.A(_0430_),
    .X(_0431_));
 sg13g2_nand2b_1 _1107_ (.Y(_0029_),
    .B(_0431_),
    .A_N(\top_inst.sndgen_inst.c2[0] ));
 sg13g2_xnor2_1 _1108_ (.Y(_0432_),
    .A(_0417_),
    .B(\top_inst.sndgen_inst.bar_counter[3] ));
 sg13g2_nand2_1 _1109_ (.Y(_0433_),
    .A(\top_inst.sndgen_inst.c2[1] ),
    .B(_0431_));
 sg13g2_o21ai_1 _1110_ (.B1(_0433_),
    .Y(_0030_),
    .A1(_0431_),
    .A2(_0432_));
 sg13g2_mux2_1 _1111_ (.A0(\top_inst.sndgen_inst.bar_counter[3] ),
    .A1(\top_inst.sndgen_inst.c2[2] ),
    .S(_0431_),
    .X(_0031_));
 sg13g2_buf_8 _1112_ (.A(\top_inst.sndgen_inst.lfsr[7] ),
    .X(_0434_));
 sg13g2_mux2_1 _1113_ (.A0(net34),
    .A1(\top_inst.sndgen_inst.c3[0] ),
    .S(net12),
    .X(_0032_));
 sg13g2_buf_2 _1114_ (.A(\top_inst.sndgen_inst.lfsr[5] ),
    .X(_0435_));
 sg13g2_nand2_1 _1115_ (.Y(_0436_),
    .A(_0435_),
    .B(_0009_));
 sg13g2_nand3_1 _1116_ (.B(net34),
    .C(_0436_),
    .A(\top_inst.sndgen_inst.lfsr[3] ),
    .Y(_0437_));
 sg13g2_nand2_1 _1117_ (.Y(_0438_),
    .A(\top_inst.sndgen_inst.c3[1] ),
    .B(net12));
 sg13g2_o21ai_1 _1118_ (.B1(_0438_),
    .Y(_0033_),
    .A1(net12),
    .A2(_0437_));
 sg13g2_nand2b_1 _1119_ (.Y(_0439_),
    .B(net34),
    .A_N(_0435_));
 sg13g2_nand2_1 _1120_ (.Y(_0440_),
    .A(\top_inst.sndgen_inst.c4[2] ),
    .B(net12));
 sg13g2_o21ai_1 _1121_ (.B1(_0440_),
    .Y(_0034_),
    .A1(net12),
    .A2(_0439_));
 sg13g2_nand2_1 _1122_ (.Y(_0441_),
    .A(net34),
    .B(_0435_));
 sg13g2_nand2_1 _1123_ (.Y(_0442_),
    .A(\top_inst.sndgen_inst.c3[2] ),
    .B(_0415_));
 sg13g2_o21ai_1 _1124_ (.B1(_0442_),
    .Y(_0035_),
    .A1(_0415_),
    .A2(_0441_));
 sg13g2_inv_1 _1125_ (.Y(_0443_),
    .A(_0396_));
 sg13g2_inv_2 _1126_ (.Y(_0444_),
    .A(_0390_));
 sg13g2_nor2_1 _1127_ (.A(net38),
    .B(_0387_),
    .Y(_0445_));
 sg13g2_and3_1 _1128_ (.X(_0446_),
    .A(_0444_),
    .B(net36),
    .C(_0445_));
 sg13g2_nand4_1 _1129_ (.B(_0389_),
    .C(_0443_),
    .A(_0398_),
    .Y(_0447_),
    .D(_0446_));
 sg13g2_buf_1 _1130_ (.A(_0447_),
    .X(_0448_));
 sg13g2_buf_1 _1131_ (.A(net21),
    .X(_0449_));
 sg13g2_mux2_1 _1132_ (.A0(_0009_),
    .A1(_0021_),
    .S(_0449_),
    .X(_0036_));
 sg13g2_and4_1 _1133_ (.A(_0398_),
    .B(_0389_),
    .C(_0443_),
    .D(_0446_),
    .X(_0450_));
 sg13g2_buf_2 _1134_ (.A(_0450_),
    .X(_0451_));
 sg13g2_buf_1 _1135_ (.A(_0451_),
    .X(_0452_));
 sg13g2_mux2_1 _1136_ (.A0(\top_inst.sndgen_inst.lfsr[1] ),
    .A1(\top_inst.sndgen_inst.lfsr[0] ),
    .S(net16),
    .X(_0037_));
 sg13g2_mux2_1 _1137_ (.A0(\top_inst.sndgen_inst.lfsr[2] ),
    .A1(\top_inst.sndgen_inst.lfsr[1] ),
    .S(net16),
    .X(_0038_));
 sg13g2_mux2_1 _1138_ (.A0(\top_inst.sndgen_inst.lfsr[3] ),
    .A1(\top_inst.sndgen_inst.lfsr[2] ),
    .S(net16),
    .X(_0039_));
 sg13g2_buf_1 _1139_ (.A(net21),
    .X(_0453_));
 sg13g2_xnor2_1 _1140_ (.Y(_0454_),
    .A(\top_inst.sndgen_inst.lfsr[3] ),
    .B(net34));
 sg13g2_nand2_1 _1141_ (.Y(_0455_),
    .A(\top_inst.sndgen_inst.lfsr[4] ),
    .B(net15));
 sg13g2_o21ai_1 _1142_ (.B1(_0455_),
    .Y(_0040_),
    .A1(net15),
    .A2(_0454_));
 sg13g2_xnor2_1 _1143_ (.Y(_0456_),
    .A(net34),
    .B(\top_inst.sndgen_inst.lfsr[4] ));
 sg13g2_nand2_1 _1144_ (.Y(_0457_),
    .A(_0435_),
    .B(net15));
 sg13g2_o21ai_1 _1145_ (.B1(_0457_),
    .Y(_0041_),
    .A1(net15),
    .A2(_0456_));
 sg13g2_xnor2_1 _1146_ (.Y(_0458_),
    .A(_0434_),
    .B(_0435_));
 sg13g2_nor2_1 _1147_ (.A(\top_inst.sndgen_inst.lfsr[6] ),
    .B(net16),
    .Y(_0459_));
 sg13g2_a21oi_1 _1148_ (.A1(net16),
    .A2(_0458_),
    .Y(_0042_),
    .B1(_0459_));
 sg13g2_mux2_1 _1149_ (.A0(_0434_),
    .A1(\top_inst.sndgen_inst.lfsr[6] ),
    .S(net16),
    .X(_0043_));
 sg13g2_nand4_1 _1150_ (.B(_0416_),
    .C(_0417_),
    .A(_0419_),
    .Y(_0460_),
    .D(\top_inst.sndgen_inst.bar_counter[3] ));
 sg13g2_nor4_1 _1151_ (.A(_0019_),
    .B(_0412_),
    .C(net21),
    .D(_0460_),
    .Y(_0461_));
 sg13g2_buf_2 _1152_ (.A(_0461_),
    .X(_0462_));
 sg13g2_mux2_1 _1153_ (.A0(\top_inst.sndgen_inst.mask_1[0] ),
    .A1(\top_inst.sndgen_inst.lfsr[1] ),
    .S(_0462_),
    .X(_0044_));
 sg13g2_mux2_1 _1154_ (.A0(\top_inst.sndgen_inst.mask_1[1] ),
    .A1(\top_inst.sndgen_inst.lfsr[2] ),
    .S(_0462_),
    .X(_0045_));
 sg13g2_buf_1 _1155_ (.A(\top_inst.sndgen_inst.mask_1[2] ),
    .X(_0463_));
 sg13g2_inv_2 _1156_ (.Y(_0464_),
    .A(_0463_));
 sg13g2_nand2_1 _1157_ (.Y(_0465_),
    .A(\top_inst.sndgen_inst.lfsr[3] ),
    .B(_0462_));
 sg13g2_o21ai_1 _1158_ (.B1(_0465_),
    .Y(_0046_),
    .A1(_0464_),
    .A2(_0462_));
 sg13g2_buf_1 _1159_ (.A(\top_inst.sndgen_inst.mask_1[3] ),
    .X(_0466_));
 sg13g2_inv_1 _1160_ (.Y(_0467_),
    .A(_0466_));
 sg13g2_nand2_1 _1161_ (.Y(_0468_),
    .A(\top_inst.sndgen_inst.lfsr[4] ),
    .B(_0462_));
 sg13g2_o21ai_1 _1162_ (.B1(_0468_),
    .Y(_0047_),
    .A1(_0467_),
    .A2(_0462_));
 sg13g2_nor3_1 _1163_ (.A(\top_inst.sndgen_inst.lfsr[3] ),
    .B(\top_inst.sndgen_inst.lfsr[2] ),
    .C(\top_inst.sndgen_inst.lfsr[1] ),
    .Y(_0469_));
 sg13g2_nor2_1 _1164_ (.A(_0022_),
    .B(_0462_),
    .Y(_0470_));
 sg13g2_a21oi_1 _1165_ (.A1(_0462_),
    .A2(_0469_),
    .Y(_0048_),
    .B1(_0470_));
 sg13g2_buf_2 _1166_ (.A(\top_inst.sndgen_inst.rom_addr[3] ),
    .X(_0471_));
 sg13g2_buf_1 _1167_ (.A(\top_inst.sndgen_inst.rom_addr[1] ),
    .X(_0472_));
 sg13g2_nand2_1 _1168_ (.Y(_0473_),
    .A(net32),
    .B(_0004_));
 sg13g2_buf_2 _1169_ (.A(\top_inst.sndgen_inst.rom_addr[0] ),
    .X(_0474_));
 sg13g2_inv_1 _1170_ (.Y(_0475_),
    .A(_0474_));
 sg13g2_a21oi_2 _1171_ (.B1(_0475_),
    .Y(_0476_),
    .A2(_0473_),
    .A1(_0471_));
 sg13g2_buf_1 _1172_ (.A(\top_inst.sndgen_inst.sample_ena_delay[0] ),
    .X(_0477_));
 sg13g2_buf_1 _1173_ (.A(net31),
    .X(_0478_));
 sg13g2_mux2_1 _1174_ (.A0(\top_inst.sndgen_inst.p_c2[0] ),
    .A1(_0476_),
    .S(net26),
    .X(_0049_));
 sg13g2_buf_2 _1175_ (.A(\top_inst.sndgen_inst.rom_addr[2] ),
    .X(_0479_));
 sg13g2_nor2_2 _1176_ (.A(_0475_),
    .B(_0479_),
    .Y(_0480_));
 sg13g2_a21oi_1 _1177_ (.A1(_0479_),
    .A2(_0003_),
    .Y(_0481_),
    .B1(_0480_));
 sg13g2_nor2_1 _1178_ (.A(net31),
    .B(\top_inst.sndgen_inst.p_c2[10] ),
    .Y(_0482_));
 sg13g2_a21oi_1 _1179_ (.A1(net26),
    .A2(_0481_),
    .Y(_0050_),
    .B1(_0482_));
 sg13g2_inv_1 _1180_ (.Y(_0483_),
    .A(\top_inst.sndgen_inst.p_c2[1] ));
 sg13g2_inv_1 _1181_ (.Y(_0484_),
    .A(_0471_));
 sg13g2_inv_1 _1182_ (.Y(_0485_),
    .A(_0480_));
 sg13g2_nand2_2 _1183_ (.Y(_0486_),
    .A(_0479_),
    .B(_0484_));
 sg13g2_a22oi_1 _1184_ (.Y(_0487_),
    .B1(_0485_),
    .B2(_0486_),
    .A2(_0484_),
    .A1(_0472_));
 sg13g2_nand2_1 _1185_ (.Y(_0488_),
    .A(net26),
    .B(_0487_));
 sg13g2_o21ai_1 _1186_ (.B1(_0488_),
    .Y(_0051_),
    .A1(net26),
    .A2(_0483_));
 sg13g2_buf_2 _1187_ (.A(\top_inst.sndgen_inst.p_c2[2] ),
    .X(_0489_));
 sg13g2_nand2_1 _1188_ (.Y(_0490_),
    .A(_0471_),
    .B(_0480_));
 sg13g2_a21oi_2 _1189_ (.B1(net32),
    .Y(_0491_),
    .A2(_0490_),
    .A1(_0486_));
 sg13g2_mux2_1 _1190_ (.A0(_0489_),
    .A1(_0491_),
    .S(_0478_),
    .X(_0052_));
 sg13g2_nor2_1 _1191_ (.A(_0474_),
    .B(_0486_),
    .Y(_0492_));
 sg13g2_o21ai_1 _1192_ (.B1(_0479_),
    .Y(_0493_),
    .A1(net32),
    .A2(_0471_));
 sg13g2_a22oi_1 _1193_ (.Y(_0494_),
    .B1(_0493_),
    .B2(_0474_),
    .A2(_0492_),
    .A1(_0472_));
 sg13g2_nor2_1 _1194_ (.A(_0477_),
    .B(\top_inst.sndgen_inst.p_c2[3] ),
    .Y(_0495_));
 sg13g2_a21oi_1 _1195_ (.A1(_0478_),
    .A2(_0494_),
    .Y(_0053_),
    .B1(_0495_));
 sg13g2_nand3_1 _1196_ (.B(_0004_),
    .C(_0471_),
    .A(net32),
    .Y(_0496_));
 sg13g2_mux2_1 _1197_ (.A0(_0486_),
    .A1(_0496_),
    .S(_0474_),
    .X(_0497_));
 sg13g2_nor2_1 _1198_ (.A(net31),
    .B(\top_inst.sndgen_inst.p_c2[4] ),
    .Y(_0498_));
 sg13g2_a21oi_1 _1199_ (.A1(net26),
    .A2(_0497_),
    .Y(_0054_),
    .B1(_0498_));
 sg13g2_nand2_1 _1200_ (.Y(_0499_),
    .A(net32),
    .B(_0484_));
 sg13g2_inv_1 _1201_ (.Y(_0500_),
    .A(net32));
 sg13g2_a21oi_1 _1202_ (.A1(_0500_),
    .A2(_0474_),
    .Y(_0501_),
    .B1(_0471_));
 sg13g2_a22oi_1 _1203_ (.Y(_0502_),
    .B1(_0501_),
    .B2(_0479_),
    .A2(_0499_),
    .A1(_0480_));
 sg13g2_buf_2 _1204_ (.A(\top_inst.sndgen_inst.p_c2[5] ),
    .X(_0503_));
 sg13g2_nor2_1 _1205_ (.A(net31),
    .B(_0503_),
    .Y(_0504_));
 sg13g2_a21oi_1 _1206_ (.A1(net26),
    .A2(_0502_),
    .Y(_0055_),
    .B1(_0504_));
 sg13g2_inv_1 _1207_ (.Y(_0505_),
    .A(_0004_));
 sg13g2_o21ai_1 _1208_ (.B1(_0486_),
    .Y(_0506_),
    .A1(_0475_),
    .A2(_0505_));
 sg13g2_a22oi_1 _1209_ (.Y(_0507_),
    .B1(_0506_),
    .B2(net32),
    .A2(_0480_),
    .A1(_0484_));
 sg13g2_nor2_1 _1210_ (.A(net31),
    .B(\top_inst.sndgen_inst.p_c2[6] ),
    .Y(_0508_));
 sg13g2_a21oi_1 _1211_ (.A1(net26),
    .A2(_0507_),
    .Y(_0056_),
    .B1(_0508_));
 sg13g2_o21ai_1 _1212_ (.B1(_0496_),
    .Y(_0509_),
    .A1(_0479_),
    .A2(_0471_));
 sg13g2_nor2_1 _1213_ (.A(net32),
    .B(_0486_),
    .Y(_0510_));
 sg13g2_a21oi_1 _1214_ (.A1(_0474_),
    .A2(_0509_),
    .Y(_0511_),
    .B1(_0510_));
 sg13g2_nor2_1 _1215_ (.A(net31),
    .B(\top_inst.sndgen_inst.p_c2[7] ),
    .Y(_0512_));
 sg13g2_a21oi_1 _1216_ (.A1(net26),
    .A2(_0511_),
    .Y(_0057_),
    .B1(_0512_));
 sg13g2_buf_1 _1217_ (.A(\top_inst.sndgen_inst.sample_ena_delay[1] ),
    .X(_0513_));
 sg13g2_buf_1 _1218_ (.A(_0513_),
    .X(_0514_));
 sg13g2_mux2_1 _1219_ (.A0(\top_inst.sndgen_inst.p_c3[0] ),
    .A1(_0476_),
    .S(net25),
    .X(_0058_));
 sg13g2_nor2_1 _1220_ (.A(net30),
    .B(\top_inst.sndgen_inst.p_c3[10] ),
    .Y(_0515_));
 sg13g2_a21oi_1 _1221_ (.A1(_0514_),
    .A2(_0481_),
    .Y(_0059_),
    .B1(_0515_));
 sg13g2_mux2_1 _1222_ (.A0(\top_inst.sndgen_inst.p_c3[1] ),
    .A1(_0487_),
    .S(net30),
    .X(_0060_));
 sg13g2_mux2_1 _1223_ (.A0(\top_inst.sndgen_inst.p_c3[2] ),
    .A1(_0491_),
    .S(net30),
    .X(_0061_));
 sg13g2_nor2_1 _1224_ (.A(net30),
    .B(\top_inst.sndgen_inst.p_c3[3] ),
    .Y(_0516_));
 sg13g2_a21oi_1 _1225_ (.A1(net25),
    .A2(_0494_),
    .Y(_0062_),
    .B1(_0516_));
 sg13g2_buf_1 _1226_ (.A(\top_inst.sndgen_inst.p_c3[4] ),
    .X(_0517_));
 sg13g2_nor2_1 _1227_ (.A(net30),
    .B(_0517_),
    .Y(_0518_));
 sg13g2_a21oi_1 _1228_ (.A1(net25),
    .A2(_0497_),
    .Y(_0063_),
    .B1(_0518_));
 sg13g2_buf_2 _1229_ (.A(\top_inst.sndgen_inst.p_c3[5] ),
    .X(_0519_));
 sg13g2_nor2_1 _1230_ (.A(net30),
    .B(_0519_),
    .Y(_0520_));
 sg13g2_a21oi_1 _1231_ (.A1(net25),
    .A2(_0502_),
    .Y(_0064_),
    .B1(_0520_));
 sg13g2_nor2_1 _1232_ (.A(net30),
    .B(\top_inst.sndgen_inst.p_c3[6] ),
    .Y(_0521_));
 sg13g2_a21oi_1 _1233_ (.A1(net25),
    .A2(_0507_),
    .Y(_0065_),
    .B1(_0521_));
 sg13g2_buf_1 _1234_ (.A(\top_inst.sndgen_inst.p_c3[7] ),
    .X(_0522_));
 sg13g2_nor2_1 _1235_ (.A(net30),
    .B(_0522_),
    .Y(_0523_));
 sg13g2_a21oi_1 _1236_ (.A1(_0514_),
    .A2(_0511_),
    .Y(_0066_),
    .B1(_0523_));
 sg13g2_buf_2 _1237_ (.A(\top_inst.sndgen_inst.sample_ena_delay[2] ),
    .X(_0524_));
 sg13g2_mux2_1 _1238_ (.A0(\top_inst.sndgen_inst.p_c4[0] ),
    .A1(_0476_),
    .S(_0524_),
    .X(_0067_));
 sg13g2_buf_1 _1239_ (.A(_0524_),
    .X(_0525_));
 sg13g2_nor2_1 _1240_ (.A(\top_inst.sndgen_inst.p_c4[10] ),
    .B(net24),
    .Y(_0526_));
 sg13g2_a21oi_1 _1241_ (.A1(net24),
    .A2(_0481_),
    .Y(_0068_),
    .B1(_0526_));
 sg13g2_inv_1 _1242_ (.Y(_0527_),
    .A(\top_inst.sndgen_inst.p_c4[1] ));
 sg13g2_nand2_1 _1243_ (.Y(_0528_),
    .A(net24),
    .B(_0487_));
 sg13g2_o21ai_1 _1244_ (.B1(_0528_),
    .Y(_0069_),
    .A1(_0527_),
    .A2(net24));
 sg13g2_mux2_1 _1245_ (.A0(\top_inst.sndgen_inst.p_c4[2] ),
    .A1(_0491_),
    .S(_0524_),
    .X(_0070_));
 sg13g2_nor2_1 _1246_ (.A(\top_inst.sndgen_inst.p_c4[3] ),
    .B(net24),
    .Y(_0529_));
 sg13g2_a21oi_1 _1247_ (.A1(net24),
    .A2(_0494_),
    .Y(_0071_),
    .B1(_0529_));
 sg13g2_nor2_1 _1248_ (.A(\top_inst.sndgen_inst.p_c4[4] ),
    .B(_0524_),
    .Y(_0530_));
 sg13g2_a21oi_1 _1249_ (.A1(net24),
    .A2(_0497_),
    .Y(_0072_),
    .B1(_0530_));
 sg13g2_nor2_1 _1250_ (.A(\top_inst.sndgen_inst.p_c4[5] ),
    .B(_0524_),
    .Y(_0531_));
 sg13g2_a21oi_1 _1251_ (.A1(_0525_),
    .A2(_0502_),
    .Y(_0073_),
    .B1(_0531_));
 sg13g2_buf_2 _1252_ (.A(\top_inst.sndgen_inst.p_c4[6] ),
    .X(_0532_));
 sg13g2_nor2_1 _1253_ (.A(_0532_),
    .B(_0524_),
    .Y(_0533_));
 sg13g2_a21oi_1 _1254_ (.A1(_0525_),
    .A2(_0507_),
    .Y(_0074_),
    .B1(_0533_));
 sg13g2_nor2_1 _1255_ (.A(\top_inst.sndgen_inst.p_c4[7] ),
    .B(_0524_),
    .Y(_0534_));
 sg13g2_a21oi_1 _1256_ (.A1(net24),
    .A2(_0511_),
    .Y(_0075_),
    .B1(_0534_));
 sg13g2_and2_1 _1257_ (.A(net35),
    .B(_0413_),
    .X(_0535_));
 sg13g2_buf_8 _1258_ (.A(_0535_),
    .X(_0536_));
 sg13g2_nand2_1 _1259_ (.Y(_0537_),
    .A(\top_inst.sndgen_inst.p_c2[0] ),
    .B(_0536_));
 sg13g2_xnor2_1 _1260_ (.Y(_0076_),
    .A(\top_inst.sndgen_inst.phacc2[0] ),
    .B(_0537_));
 sg13g2_inv_1 _1261_ (.Y(_0538_),
    .A(\top_inst.sndgen_inst.phacc2[4] ));
 sg13g2_nand3_1 _1262_ (.B(\top_inst.sndgen_inst.p_c2[0] ),
    .C(\top_inst.sndgen_inst.phacc2[0] ),
    .A(\top_inst.sndgen_inst.phacc2[1] ),
    .Y(_0539_));
 sg13g2_buf_2 _1263_ (.A(\top_inst.sndgen_inst.phacc2[2] ),
    .X(_0540_));
 sg13g2_o21ai_1 _1264_ (.B1(\top_inst.sndgen_inst.phacc2[3] ),
    .Y(_0541_),
    .A1(_0489_),
    .A2(_0540_));
 sg13g2_o21ai_1 _1265_ (.B1(\top_inst.sndgen_inst.p_c2[3] ),
    .Y(_0542_),
    .A1(_0489_),
    .A2(_0540_));
 sg13g2_a21oi_1 _1266_ (.A1(\top_inst.sndgen_inst.p_c2[0] ),
    .A2(\top_inst.sndgen_inst.phacc2[0] ),
    .Y(_0543_),
    .B1(\top_inst.sndgen_inst.phacc2[1] ));
 sg13g2_a221oi_1 _1267_ (.B2(_0542_),
    .C1(_0543_),
    .B1(_0541_),
    .A1(_0483_),
    .Y(_0544_),
    .A2(_0539_));
 sg13g2_nand2_1 _1268_ (.Y(_0545_),
    .A(\top_inst.sndgen_inst.p_c2[3] ),
    .B(\top_inst.sndgen_inst.phacc2[3] ));
 sg13g2_nand3_1 _1269_ (.B(_0540_),
    .C(\top_inst.sndgen_inst.phacc2[3] ),
    .A(_0489_),
    .Y(_0546_));
 sg13g2_nand3_1 _1270_ (.B(_0540_),
    .C(\top_inst.sndgen_inst.p_c2[3] ),
    .A(_0489_),
    .Y(_0547_));
 sg13g2_nand3_1 _1271_ (.B(_0546_),
    .C(_0547_),
    .A(_0545_),
    .Y(_0548_));
 sg13g2_nor2_1 _1272_ (.A(_0544_),
    .B(_0548_),
    .Y(_0549_));
 sg13g2_buf_1 _1273_ (.A(\top_inst.sndgen_inst.phacc2[5] ),
    .X(_0550_));
 sg13g2_o21ai_1 _1274_ (.B1(_0550_),
    .Y(_0551_),
    .A1(\top_inst.sndgen_inst.p_c2[6] ),
    .A2(\top_inst.sndgen_inst.phacc2[6] ));
 sg13g2_o21ai_1 _1275_ (.B1(_0503_),
    .Y(_0552_),
    .A1(\top_inst.sndgen_inst.p_c2[6] ),
    .A2(\top_inst.sndgen_inst.phacc2[6] ));
 sg13g2_inv_1 _1276_ (.Y(_0553_),
    .A(\top_inst.sndgen_inst.p_c2[4] ));
 sg13g2_a221oi_1 _1277_ (.B2(_0552_),
    .C1(_0553_),
    .B1(_0551_),
    .A1(_0538_),
    .Y(_0554_),
    .A2(_0549_));
 sg13g2_inv_1 _1278_ (.Y(_0555_),
    .A(\top_inst.sndgen_inst.p_c2[6] ));
 sg13g2_inv_1 _1279_ (.Y(_0556_),
    .A(\top_inst.sndgen_inst.phacc2[6] ));
 sg13g2_nand2_1 _1280_ (.Y(_0557_),
    .A(\top_inst.sndgen_inst.phacc2[4] ),
    .B(_0550_));
 sg13g2_nand2_1 _1281_ (.Y(_0558_),
    .A(\top_inst.sndgen_inst.phacc2[4] ),
    .B(_0503_));
 sg13g2_a221oi_1 _1282_ (.B2(_0558_),
    .C1(_0549_),
    .B1(_0557_),
    .A1(_0555_),
    .Y(_0559_),
    .A2(_0556_));
 sg13g2_nand2_1 _1283_ (.Y(_0560_),
    .A(_0503_),
    .B(_0550_));
 sg13g2_a21oi_1 _1284_ (.A1(_0555_),
    .A2(_0556_),
    .Y(_0561_),
    .B1(_0560_));
 sg13g2_nor2_1 _1285_ (.A(_0555_),
    .B(_0556_),
    .Y(_0562_));
 sg13g2_or4_1 _1286_ (.A(_0554_),
    .B(_0559_),
    .C(_0561_),
    .D(_0562_),
    .X(_0563_));
 sg13g2_buf_1 _1287_ (.A(_0563_),
    .X(_0564_));
 sg13g2_o21ai_1 _1288_ (.B1(\top_inst.sndgen_inst.p_c2[7] ),
    .Y(_0565_),
    .A1(\top_inst.sndgen_inst.phacc2[7] ),
    .A2(_0564_));
 sg13g2_nand2_1 _1289_ (.Y(_0566_),
    .A(\top_inst.sndgen_inst.phacc2[7] ),
    .B(_0564_));
 sg13g2_a21oi_1 _1290_ (.A1(_0565_),
    .A2(_0566_),
    .Y(_0567_),
    .B1(_0001_));
 sg13g2_nand2b_1 _1291_ (.Y(_0568_),
    .B(\top_inst.sndgen_inst.p_c2[10] ),
    .A_N(\top_inst.sndgen_inst.phacc2[9] ));
 sg13g2_nor2_1 _1292_ (.A(_0567_),
    .B(_0568_),
    .Y(_0569_));
 sg13g2_nor2b_1 _1293_ (.A(\top_inst.sndgen_inst.p_c2[10] ),
    .B_N(\top_inst.sndgen_inst.phacc2[9] ),
    .Y(_0570_));
 sg13g2_and2_1 _1294_ (.A(_0567_),
    .B(_0570_),
    .X(_0571_));
 sg13g2_o21ai_1 _1295_ (.B1(_0536_),
    .Y(_0572_),
    .A1(_0569_),
    .A2(_0571_));
 sg13g2_xnor2_1 _1296_ (.Y(_0077_),
    .A(\top_inst.sndgen_inst.phacc2[10] ),
    .B(_0572_));
 sg13g2_nor2_1 _1297_ (.A(_0019_),
    .B(net21),
    .Y(_0573_));
 sg13g2_nand4_1 _1298_ (.B(\top_inst.sndgen_inst.phacc2[10] ),
    .C(_0573_),
    .A(_0409_),
    .Y(_0574_),
    .D(_0570_));
 sg13g2_nand2_1 _1299_ (.Y(_0575_),
    .A(net35),
    .B(_0573_));
 sg13g2_or3_1 _1300_ (.A(\top_inst.sndgen_inst.phacc2[10] ),
    .B(net11),
    .C(_0568_),
    .X(_0576_));
 sg13g2_nand2b_1 _1301_ (.Y(_0577_),
    .B(_0564_),
    .A_N(_0001_));
 sg13g2_nand2_1 _1302_ (.Y(_0578_),
    .A(\top_inst.sndgen_inst.phacc2[7] ),
    .B(\top_inst.sndgen_inst.phacc2[8] ));
 sg13g2_o21ai_1 _1303_ (.B1(_0578_),
    .Y(_0579_),
    .A1(\top_inst.sndgen_inst.phacc2[7] ),
    .A2(_0577_));
 sg13g2_nor3_1 _1304_ (.A(\top_inst.sndgen_inst.p_c2[7] ),
    .B(_0001_),
    .C(_0566_),
    .Y(_0580_));
 sg13g2_a21oi_2 _1305_ (.B1(_0580_),
    .Y(_0581_),
    .A2(_0579_),
    .A1(\top_inst.sndgen_inst.p_c2[7] ));
 sg13g2_mux2_1 _1306_ (.A0(_0574_),
    .A1(_0576_),
    .S(_0581_),
    .X(_0582_));
 sg13g2_xnor2_1 _1307_ (.Y(_0078_),
    .A(\top_inst.sndgen_inst.phacc2[11] ),
    .B(_0582_));
 sg13g2_nor3_1 _1308_ (.A(\top_inst.sndgen_inst.phacc2[10] ),
    .B(\top_inst.sndgen_inst.phacc2[11] ),
    .C(_0568_),
    .Y(_0583_));
 sg13g2_nand2_1 _1309_ (.Y(_0584_),
    .A(_0536_),
    .B(_0583_));
 sg13g2_nand4_1 _1310_ (.B(\top_inst.sndgen_inst.phacc2[11] ),
    .C(_0536_),
    .A(\top_inst.sndgen_inst.phacc2[10] ),
    .Y(_0585_),
    .D(_0570_));
 sg13g2_mux2_1 _1311_ (.A0(_0584_),
    .A1(_0585_),
    .S(_0567_),
    .X(_0586_));
 sg13g2_xnor2_1 _1312_ (.Y(_0079_),
    .A(\top_inst.sndgen_inst.phacc2[12] ),
    .B(_0586_));
 sg13g2_inv_1 _1313_ (.Y(_0587_),
    .A(\top_inst.sndgen_inst.phacc2[12] ));
 sg13g2_or2_1 _1314_ (.X(_0588_),
    .B(_0585_),
    .A(_0587_));
 sg13g2_nand3_1 _1315_ (.B(_0536_),
    .C(_0583_),
    .A(_0587_),
    .Y(_0589_));
 sg13g2_mux2_1 _1316_ (.A0(_0588_),
    .A1(_0589_),
    .S(_0581_),
    .X(_0590_));
 sg13g2_xnor2_1 _1317_ (.Y(_0080_),
    .A(\top_inst.sndgen_inst.phacc2[13] ),
    .B(_0590_));
 sg13g2_nand2_1 _1318_ (.Y(_0591_),
    .A(\top_inst.sndgen_inst.p_c2[0] ),
    .B(\top_inst.sndgen_inst.phacc2[0] ));
 sg13g2_xnor2_1 _1319_ (.Y(_0592_),
    .A(_0483_),
    .B(_0591_));
 sg13g2_nor2_1 _1320_ (.A(net11),
    .B(_0592_),
    .Y(_0593_));
 sg13g2_xor2_1 _1321_ (.B(_0593_),
    .A(\top_inst.sndgen_inst.phacc2[1] ),
    .X(_0081_));
 sg13g2_o21ai_1 _1322_ (.B1(_0539_),
    .Y(_0594_),
    .A1(_0483_),
    .A2(_0543_));
 sg13g2_xnor2_1 _1323_ (.Y(_0595_),
    .A(_0489_),
    .B(_0594_));
 sg13g2_nor2_1 _1324_ (.A(net11),
    .B(_0595_),
    .Y(_0596_));
 sg13g2_xor2_1 _1325_ (.B(_0596_),
    .A(_0540_),
    .X(_0082_));
 sg13g2_a21o_1 _1326_ (.A2(_0540_),
    .A1(_0489_),
    .B1(_0594_),
    .X(_0597_));
 sg13g2_o21ai_1 _1327_ (.B1(_0597_),
    .Y(_0598_),
    .A1(_0489_),
    .A2(_0540_));
 sg13g2_xor2_1 _1328_ (.B(_0598_),
    .A(\top_inst.sndgen_inst.p_c2[3] ),
    .X(_0599_));
 sg13g2_nor2_1 _1329_ (.A(net11),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_xor2_1 _1330_ (.B(_0600_),
    .A(\top_inst.sndgen_inst.phacc2[3] ),
    .X(_0083_));
 sg13g2_or2_1 _1331_ (.X(_0601_),
    .B(_0548_),
    .A(_0544_));
 sg13g2_xnor2_1 _1332_ (.Y(_0602_),
    .A(\top_inst.sndgen_inst.p_c2[4] ),
    .B(_0601_));
 sg13g2_nor2_1 _1333_ (.A(_0575_),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_xnor2_1 _1334_ (.Y(_0084_),
    .A(_0538_),
    .B(_0603_));
 sg13g2_o21ai_1 _1335_ (.B1(\top_inst.sndgen_inst.p_c2[4] ),
    .Y(_0604_),
    .A1(\top_inst.sndgen_inst.phacc2[4] ),
    .A2(_0601_));
 sg13g2_nand2_1 _1336_ (.Y(_0605_),
    .A(\top_inst.sndgen_inst.phacc2[4] ),
    .B(_0601_));
 sg13g2_and2_1 _1337_ (.A(_0604_),
    .B(_0605_),
    .X(_0606_));
 sg13g2_xor2_1 _1338_ (.B(_0606_),
    .A(_0503_),
    .X(_0607_));
 sg13g2_nor2_1 _1339_ (.A(net11),
    .B(_0607_),
    .Y(_0608_));
 sg13g2_xor2_1 _1340_ (.B(_0608_),
    .A(_0550_),
    .X(_0085_));
 sg13g2_nand2b_1 _1341_ (.Y(_0609_),
    .B(_0606_),
    .A_N(_0550_));
 sg13g2_nor2b_1 _1342_ (.A(_0606_),
    .B_N(_0550_),
    .Y(_0610_));
 sg13g2_a21oi_1 _1343_ (.A1(_0503_),
    .A2(_0609_),
    .Y(_0611_),
    .B1(_0610_));
 sg13g2_xnor2_1 _1344_ (.Y(_0612_),
    .A(_0555_),
    .B(_0611_));
 sg13g2_nor2_1 _1345_ (.A(net11),
    .B(_0612_),
    .Y(_0613_));
 sg13g2_xnor2_1 _1346_ (.Y(_0086_),
    .A(_0556_),
    .B(_0613_));
 sg13g2_xnor2_1 _1347_ (.Y(_0614_),
    .A(\top_inst.sndgen_inst.p_c2[7] ),
    .B(_0564_));
 sg13g2_nor2_1 _1348_ (.A(net11),
    .B(_0614_),
    .Y(_0615_));
 sg13g2_xor2_1 _1349_ (.B(_0615_),
    .A(\top_inst.sndgen_inst.phacc2[7] ),
    .X(_0087_));
 sg13g2_nand2_1 _1350_ (.Y(_0616_),
    .A(_0565_),
    .B(_0566_));
 sg13g2_xor2_1 _1351_ (.B(_0616_),
    .A(_0001_),
    .X(_0617_));
 sg13g2_nor2_1 _1352_ (.A(\top_inst.sndgen_inst.phacc2[8] ),
    .B(_0536_),
    .Y(_0618_));
 sg13g2_a21oi_1 _1353_ (.A1(_0536_),
    .A2(_0617_),
    .Y(_0088_),
    .B1(_0618_));
 sg13g2_or2_1 _1354_ (.X(_0619_),
    .B(net11),
    .A(\top_inst.sndgen_inst.p_c2[10] ));
 sg13g2_nand3_1 _1355_ (.B(\top_inst.sndgen_inst.p_c2[10] ),
    .C(_0573_),
    .A(net35),
    .Y(_0620_));
 sg13g2_mux2_1 _1356_ (.A0(_0619_),
    .A1(_0620_),
    .S(_0581_),
    .X(_0621_));
 sg13g2_xnor2_1 _1357_ (.Y(_0089_),
    .A(\top_inst.sndgen_inst.phacc2[9] ),
    .B(_0621_));
 sg13g2_buf_1 _1358_ (.A(_0451_),
    .X(_0622_));
 sg13g2_nand2_1 _1359_ (.Y(_0623_),
    .A(\top_inst.sndgen_inst.p_c3[0] ),
    .B(net14));
 sg13g2_xnor2_1 _1360_ (.Y(_0090_),
    .A(\top_inst.sndgen_inst.phacc3[0] ),
    .B(_0623_));
 sg13g2_nor2b_1 _1361_ (.A(\top_inst.sndgen_inst.p_c3[10] ),
    .B_N(\top_inst.sndgen_inst.phacc3[9] ),
    .Y(_0624_));
 sg13g2_nand2_1 _1362_ (.Y(_0625_),
    .A(net22),
    .B(_0624_));
 sg13g2_nor2b_1 _1363_ (.A(\top_inst.sndgen_inst.phacc3[9] ),
    .B_N(\top_inst.sndgen_inst.p_c3[10] ),
    .Y(_0626_));
 sg13g2_nand2_1 _1364_ (.Y(_0627_),
    .A(net22),
    .B(_0626_));
 sg13g2_buf_1 _1365_ (.A(\top_inst.sndgen_inst.phacc3[7] ),
    .X(_0628_));
 sg13g2_nor2_2 _1366_ (.A(\top_inst.sndgen_inst.p_c3[6] ),
    .B(\top_inst.sndgen_inst.phacc3[6] ),
    .Y(_0629_));
 sg13g2_buf_2 _1367_ (.A(\top_inst.sndgen_inst.phacc3[4] ),
    .X(_0630_));
 sg13g2_buf_2 _1368_ (.A(\top_inst.sndgen_inst.phacc3[5] ),
    .X(_0631_));
 sg13g2_nand2_1 _1369_ (.Y(_0632_),
    .A(_0630_),
    .B(_0631_));
 sg13g2_nor2_1 _1370_ (.A(_0629_),
    .B(_0632_),
    .Y(_0633_));
 sg13g2_nand2_1 _1371_ (.Y(_0634_),
    .A(_0517_),
    .B(_0631_));
 sg13g2_nor2_1 _1372_ (.A(_0629_),
    .B(_0634_),
    .Y(_0635_));
 sg13g2_and2_1 _1373_ (.A(\top_inst.sndgen_inst.p_c3[0] ),
    .B(\top_inst.sndgen_inst.phacc3[0] ),
    .X(_0636_));
 sg13g2_o21ai_1 _1374_ (.B1(\top_inst.sndgen_inst.p_c3[1] ),
    .Y(_0637_),
    .A1(\top_inst.sndgen_inst.phacc3[1] ),
    .A2(_0636_));
 sg13g2_nand3_1 _1375_ (.B(\top_inst.sndgen_inst.p_c3[0] ),
    .C(\top_inst.sndgen_inst.phacc3[0] ),
    .A(\top_inst.sndgen_inst.phacc3[1] ),
    .Y(_0638_));
 sg13g2_a22oi_1 _1376_ (.Y(_0639_),
    .B1(\top_inst.sndgen_inst.p_c3[3] ),
    .B2(\top_inst.sndgen_inst.phacc3[3] ),
    .A2(\top_inst.sndgen_inst.phacc3[2] ),
    .A1(\top_inst.sndgen_inst.p_c3[2] ));
 sg13g2_and2_1 _1377_ (.A(_0638_),
    .B(_0639_),
    .X(_0640_));
 sg13g2_nor2_1 _1378_ (.A(\top_inst.sndgen_inst.p_c3[2] ),
    .B(\top_inst.sndgen_inst.phacc3[2] ),
    .Y(_0641_));
 sg13g2_nor2_1 _1379_ (.A(\top_inst.sndgen_inst.p_c3[3] ),
    .B(\top_inst.sndgen_inst.phacc3[3] ),
    .Y(_0642_));
 sg13g2_a221oi_1 _1380_ (.B2(_0639_),
    .C1(_0642_),
    .B1(_0641_),
    .A1(_0637_),
    .Y(_0643_),
    .A2(_0640_));
 sg13g2_buf_1 _1381_ (.A(_0643_),
    .X(_0644_));
 sg13g2_o21ai_1 _1382_ (.B1(_0644_),
    .Y(_0645_),
    .A1(_0633_),
    .A2(_0635_));
 sg13g2_nand2_1 _1383_ (.Y(_0646_),
    .A(_0630_),
    .B(_0519_));
 sg13g2_nor2_1 _1384_ (.A(_0629_),
    .B(_0646_),
    .Y(_0647_));
 sg13g2_nand2_1 _1385_ (.Y(_0648_),
    .A(_0517_),
    .B(_0519_));
 sg13g2_nor2_1 _1386_ (.A(_0629_),
    .B(_0648_),
    .Y(_0649_));
 sg13g2_o21ai_1 _1387_ (.B1(_0644_),
    .Y(_0650_),
    .A1(_0647_),
    .A2(_0649_));
 sg13g2_nand2_1 _1388_ (.Y(_0651_),
    .A(_0519_),
    .B(_0631_));
 sg13g2_nor2_1 _1389_ (.A(_0629_),
    .B(_0651_),
    .Y(_0652_));
 sg13g2_nand2_1 _1390_ (.Y(_0653_),
    .A(_0517_),
    .B(_0630_));
 sg13g2_nor2_1 _1391_ (.A(_0629_),
    .B(_0653_),
    .Y(_0654_));
 sg13g2_o21ai_1 _1392_ (.B1(_0654_),
    .Y(_0655_),
    .A1(_0519_),
    .A2(_0631_));
 sg13g2_nor2b_1 _1393_ (.A(_0652_),
    .B_N(_0655_),
    .Y(_0656_));
 sg13g2_nand2_1 _1394_ (.Y(_0657_),
    .A(\top_inst.sndgen_inst.p_c3[6] ),
    .B(\top_inst.sndgen_inst.phacc3[6] ));
 sg13g2_nand4_1 _1395_ (.B(_0650_),
    .C(_0656_),
    .A(_0645_),
    .Y(_0658_),
    .D(_0657_));
 sg13g2_buf_1 _1396_ (.A(_0658_),
    .X(_0659_));
 sg13g2_nor2_1 _1397_ (.A(_0628_),
    .B(_0659_),
    .Y(_0660_));
 sg13g2_a21oi_1 _1398_ (.A1(_0628_),
    .A2(_0659_),
    .Y(_0661_),
    .B1(_0522_));
 sg13g2_nor2_1 _1399_ (.A(_0660_),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_nand2b_1 _1400_ (.Y(_0663_),
    .B(_0662_),
    .A_N(_0013_));
 sg13g2_mux2_1 _1401_ (.A0(_0625_),
    .A1(_0627_),
    .S(_0663_),
    .X(_0664_));
 sg13g2_xnor2_1 _1402_ (.Y(_0091_),
    .A(\top_inst.sndgen_inst.phacc3[10] ),
    .B(_0664_));
 sg13g2_inv_1 _1403_ (.Y(_0665_),
    .A(\top_inst.sndgen_inst.phacc3[11] ));
 sg13g2_nand2b_1 _1404_ (.Y(_0666_),
    .B(_0626_),
    .A_N(\top_inst.sndgen_inst.phacc3[10] ));
 sg13g2_nand2_1 _1405_ (.Y(_0667_),
    .A(\top_inst.sndgen_inst.phacc3[10] ),
    .B(_0624_));
 sg13g2_nand3_1 _1406_ (.B(_0628_),
    .C(\top_inst.sndgen_inst.phacc3[8] ),
    .A(_0522_),
    .Y(_0668_));
 sg13g2_nor2b_1 _1407_ (.A(_0522_),
    .B_N(_0628_),
    .Y(_0669_));
 sg13g2_nand3b_1 _1408_ (.B(_0659_),
    .C(_0669_),
    .Y(_0670_),
    .A_N(_0013_));
 sg13g2_nor2b_1 _1409_ (.A(_0628_),
    .B_N(_0522_),
    .Y(_0671_));
 sg13g2_nand3b_1 _1410_ (.B(_0659_),
    .C(_0671_),
    .Y(_0672_),
    .A_N(_0013_));
 sg13g2_nand3_1 _1411_ (.B(_0670_),
    .C(_0672_),
    .A(_0668_),
    .Y(_0673_));
 sg13g2_mux2_1 _1412_ (.A0(_0666_),
    .A1(_0667_),
    .S(_0673_),
    .X(_0674_));
 sg13g2_nor2_1 _1413_ (.A(net17),
    .B(_0674_),
    .Y(_0675_));
 sg13g2_xnor2_1 _1414_ (.Y(_0092_),
    .A(_0665_),
    .B(_0675_));
 sg13g2_nor3_1 _1415_ (.A(_0665_),
    .B(net21),
    .C(_0667_),
    .Y(_0676_));
 sg13g2_nor3_1 _1416_ (.A(\top_inst.sndgen_inst.phacc3[11] ),
    .B(net21),
    .C(_0666_),
    .Y(_0677_));
 sg13g2_mux2_1 _1417_ (.A0(_0676_),
    .A1(_0677_),
    .S(_0663_),
    .X(_0678_));
 sg13g2_xor2_1 _1418_ (.B(_0678_),
    .A(\top_inst.sndgen_inst.phacc3[12] ),
    .X(_0093_));
 sg13g2_inv_1 _1419_ (.Y(_0679_),
    .A(\top_inst.sndgen_inst.phacc3[13] ));
 sg13g2_or4_1 _1420_ (.A(\top_inst.sndgen_inst.phacc3[11] ),
    .B(\top_inst.sndgen_inst.phacc3[12] ),
    .C(_0673_),
    .D(_0666_),
    .X(_0680_));
 sg13g2_nand4_1 _1421_ (.B(\top_inst.sndgen_inst.phacc3[11] ),
    .C(\top_inst.sndgen_inst.phacc3[12] ),
    .A(\top_inst.sndgen_inst.phacc3[10] ),
    .Y(_0681_),
    .D(_0624_));
 sg13g2_nand2b_1 _1422_ (.Y(_0682_),
    .B(_0673_),
    .A_N(_0681_));
 sg13g2_a21oi_1 _1423_ (.A1(_0680_),
    .A2(_0682_),
    .Y(_0683_),
    .B1(net17));
 sg13g2_xnor2_1 _1424_ (.Y(_0094_),
    .A(_0679_),
    .B(_0683_));
 sg13g2_xor2_1 _1425_ (.B(_0636_),
    .A(\top_inst.sndgen_inst.p_c3[1] ),
    .X(_0684_));
 sg13g2_nand2_1 _1426_ (.Y(_0685_),
    .A(net22),
    .B(_0684_));
 sg13g2_xnor2_1 _1427_ (.Y(_0095_),
    .A(\top_inst.sndgen_inst.phacc3[1] ),
    .B(_0685_));
 sg13g2_inv_1 _1428_ (.Y(_0686_),
    .A(\top_inst.sndgen_inst.phacc3[2] ));
 sg13g2_and2_1 _1429_ (.A(_0638_),
    .B(_0637_),
    .X(_0687_));
 sg13g2_xor2_1 _1430_ (.B(_0687_),
    .A(\top_inst.sndgen_inst.p_c3[2] ),
    .X(_0688_));
 sg13g2_nor2_1 _1431_ (.A(net17),
    .B(_0688_),
    .Y(_0689_));
 sg13g2_xnor2_1 _1432_ (.Y(_0096_),
    .A(_0686_),
    .B(_0689_));
 sg13g2_nand2_1 _1433_ (.Y(_0690_),
    .A(_0686_),
    .B(_0687_));
 sg13g2_nor2_1 _1434_ (.A(_0686_),
    .B(_0687_),
    .Y(_0691_));
 sg13g2_a21oi_1 _1435_ (.A1(\top_inst.sndgen_inst.p_c3[2] ),
    .A2(_0690_),
    .Y(_0692_),
    .B1(_0691_));
 sg13g2_xor2_1 _1436_ (.B(_0692_),
    .A(\top_inst.sndgen_inst.p_c3[3] ),
    .X(_0693_));
 sg13g2_nor2_1 _1437_ (.A(net17),
    .B(_0693_),
    .Y(_0694_));
 sg13g2_xor2_1 _1438_ (.B(_0694_),
    .A(\top_inst.sndgen_inst.phacc3[3] ),
    .X(_0097_));
 sg13g2_buf_1 _1439_ (.A(net21),
    .X(_0695_));
 sg13g2_xnor2_1 _1440_ (.Y(_0696_),
    .A(_0517_),
    .B(_0644_));
 sg13g2_nor2_1 _1441_ (.A(net13),
    .B(_0696_),
    .Y(_0697_));
 sg13g2_xor2_1 _1442_ (.B(_0697_),
    .A(_0630_),
    .X(_0098_));
 sg13g2_nand2_1 _1443_ (.Y(_0698_),
    .A(_0630_),
    .B(_0644_));
 sg13g2_o21ai_1 _1444_ (.B1(_0517_),
    .Y(_0699_),
    .A1(_0630_),
    .A2(_0644_));
 sg13g2_nand2_1 _1445_ (.Y(_0700_),
    .A(_0698_),
    .B(_0699_));
 sg13g2_xnor2_1 _1446_ (.Y(_0701_),
    .A(_0519_),
    .B(_0700_));
 sg13g2_nor2_1 _1447_ (.A(net13),
    .B(_0701_),
    .Y(_0702_));
 sg13g2_xor2_1 _1448_ (.B(_0702_),
    .A(_0631_),
    .X(_0099_));
 sg13g2_o21ai_1 _1449_ (.B1(_0700_),
    .Y(_0703_),
    .A1(_0519_),
    .A2(_0631_));
 sg13g2_nand2_1 _1450_ (.Y(_0704_),
    .A(_0651_),
    .B(_0703_));
 sg13g2_xnor2_1 _1451_ (.Y(_0705_),
    .A(\top_inst.sndgen_inst.p_c3[6] ),
    .B(_0704_));
 sg13g2_nor2_1 _1452_ (.A(net13),
    .B(_0705_),
    .Y(_0706_));
 sg13g2_xor2_1 _1453_ (.B(_0706_),
    .A(\top_inst.sndgen_inst.phacc3[6] ),
    .X(_0100_));
 sg13g2_xnor2_1 _1454_ (.Y(_0707_),
    .A(_0522_),
    .B(_0659_));
 sg13g2_nor2_1 _1455_ (.A(net13),
    .B(_0707_),
    .Y(_0708_));
 sg13g2_xor2_1 _1456_ (.B(_0708_),
    .A(_0628_),
    .X(_0101_));
 sg13g2_xor2_1 _1457_ (.B(_0662_),
    .A(_0013_),
    .X(_0709_));
 sg13g2_nor2_1 _1458_ (.A(\top_inst.sndgen_inst.phacc3[8] ),
    .B(net22),
    .Y(_0710_));
 sg13g2_a21oi_1 _1459_ (.A1(\top_inst.sample_ena ),
    .A2(_0709_),
    .Y(_0102_),
    .B1(_0710_));
 sg13g2_xnor2_1 _1460_ (.Y(_0711_),
    .A(\top_inst.sndgen_inst.p_c3[10] ),
    .B(_0673_));
 sg13g2_nor2_1 _1461_ (.A(net13),
    .B(_0711_),
    .Y(_0712_));
 sg13g2_xor2_1 _1462_ (.B(_0712_),
    .A(\top_inst.sndgen_inst.phacc3[9] ),
    .X(_0103_));
 sg13g2_nand2_1 _1463_ (.Y(_0713_),
    .A(\top_inst.sndgen_inst.p_c4[0] ),
    .B(_0622_));
 sg13g2_xnor2_1 _1464_ (.Y(_0104_),
    .A(\top_inst.sndgen_inst.phacc4[0] ),
    .B(_0713_));
 sg13g2_inv_1 _1465_ (.Y(_0714_),
    .A(\top_inst.sndgen_inst.p_c4[10] ));
 sg13g2_nor3_1 _1466_ (.A(_0714_),
    .B(\top_inst.sndgen_inst.phacc4[9] ),
    .C(_0448_),
    .Y(_0715_));
 sg13g2_nor2b_1 _1467_ (.A(\top_inst.sndgen_inst.p_c4[10] ),
    .B_N(\top_inst.sndgen_inst.phacc4[9] ),
    .Y(_0716_));
 sg13g2_and2_1 _1468_ (.A(_0451_),
    .B(_0716_),
    .X(_0717_));
 sg13g2_buf_1 _1469_ (.A(\top_inst.sndgen_inst.phacc4[6] ),
    .X(_0718_));
 sg13g2_nor2_1 _1470_ (.A(_0532_),
    .B(_0718_),
    .Y(_0719_));
 sg13g2_a21oi_1 _1471_ (.A1(\top_inst.sndgen_inst.p_c4[0] ),
    .A2(\top_inst.sndgen_inst.phacc4[0] ),
    .Y(_0720_),
    .B1(\top_inst.sndgen_inst.phacc4[1] ));
 sg13g2_nand3_1 _1472_ (.B(\top_inst.sndgen_inst.p_c4[0] ),
    .C(\top_inst.sndgen_inst.phacc4[0] ),
    .A(\top_inst.sndgen_inst.phacc4[1] ),
    .Y(_0721_));
 sg13g2_o21ai_1 _1473_ (.B1(_0721_),
    .Y(_0722_),
    .A1(_0527_),
    .A2(_0720_));
 sg13g2_or2_1 _1474_ (.X(_0723_),
    .B(\top_inst.sndgen_inst.phacc4[2] ),
    .A(\top_inst.sndgen_inst.p_c4[2] ));
 sg13g2_a22oi_1 _1475_ (.Y(_0724_),
    .B1(\top_inst.sndgen_inst.p_c4[4] ),
    .B2(\top_inst.sndgen_inst.phacc4[4] ),
    .A2(\top_inst.sndgen_inst.phacc4[2] ),
    .A1(\top_inst.sndgen_inst.p_c4[2] ));
 sg13g2_inv_1 _1476_ (.Y(_0725_),
    .A(_0724_));
 sg13g2_a221oi_1 _1477_ (.B2(_0723_),
    .C1(_0725_),
    .B1(_0722_),
    .A1(\top_inst.sndgen_inst.p_c4[3] ),
    .Y(_0726_),
    .A2(\top_inst.sndgen_inst.phacc4[3] ));
 sg13g2_and2_1 _1478_ (.A(\top_inst.sndgen_inst.p_c4[4] ),
    .B(\top_inst.sndgen_inst.phacc4[4] ),
    .X(_0727_));
 sg13g2_or3_1 _1479_ (.A(\top_inst.sndgen_inst.p_c4[3] ),
    .B(\top_inst.sndgen_inst.phacc4[3] ),
    .C(_0727_),
    .X(_0728_));
 sg13g2_o21ai_1 _1480_ (.B1(_0728_),
    .Y(_0729_),
    .A1(\top_inst.sndgen_inst.p_c4[4] ),
    .A2(\top_inst.sndgen_inst.phacc4[4] ));
 sg13g2_inv_1 _1481_ (.Y(_0730_),
    .A(\top_inst.sndgen_inst.phacc4[5] ));
 sg13g2_o21ai_1 _1482_ (.B1(_0730_),
    .Y(_0731_),
    .A1(_0726_),
    .A2(_0729_));
 sg13g2_nor3_1 _1483_ (.A(_0730_),
    .B(_0726_),
    .C(_0729_),
    .Y(_0732_));
 sg13g2_a21oi_2 _1484_ (.B1(_0732_),
    .Y(_0733_),
    .A2(_0731_),
    .A1(\top_inst.sndgen_inst.p_c4[5] ));
 sg13g2_buf_1 _1485_ (.A(\top_inst.sndgen_inst.phacc4[7] ),
    .X(_0734_));
 sg13g2_a21oi_1 _1486_ (.A1(_0532_),
    .A2(_0718_),
    .Y(_0735_),
    .B1(net29));
 sg13g2_o21ai_1 _1487_ (.B1(_0735_),
    .Y(_0736_),
    .A1(_0719_),
    .A2(_0733_));
 sg13g2_nor2_1 _1488_ (.A(_0726_),
    .B(_0729_),
    .Y(_0737_));
 sg13g2_inv_1 _1489_ (.Y(_0738_),
    .A(_0719_));
 sg13g2_nand4_1 _1490_ (.B(net29),
    .C(_0737_),
    .A(\top_inst.sndgen_inst.phacc4[5] ),
    .Y(_0739_),
    .D(_0738_));
 sg13g2_nand4_1 _1491_ (.B(net29),
    .C(_0737_),
    .A(\top_inst.sndgen_inst.p_c4[5] ),
    .Y(_0740_),
    .D(_0738_));
 sg13g2_nand3_1 _1492_ (.B(_0718_),
    .C(net29),
    .A(_0532_),
    .Y(_0741_));
 sg13g2_nand4_1 _1493_ (.B(\top_inst.sndgen_inst.phacc4[5] ),
    .C(net29),
    .A(\top_inst.sndgen_inst.p_c4[5] ),
    .Y(_0742_),
    .D(_0738_));
 sg13g2_nand4_1 _1494_ (.B(_0740_),
    .C(_0741_),
    .A(_0739_),
    .Y(_0743_),
    .D(_0742_));
 sg13g2_a21oi_1 _1495_ (.A1(\top_inst.sndgen_inst.p_c4[7] ),
    .A2(_0736_),
    .Y(_0744_),
    .B1(_0743_));
 sg13g2_nor2_1 _1496_ (.A(_0000_),
    .B(_0744_),
    .Y(_0745_));
 sg13g2_mux2_1 _1497_ (.A0(_0715_),
    .A1(_0717_),
    .S(_0745_),
    .X(_0746_));
 sg13g2_xor2_1 _1498_ (.B(_0746_),
    .A(\top_inst.sndgen_inst.phacc4[10] ),
    .X(_0105_));
 sg13g2_nand3_1 _1499_ (.B(net22),
    .C(_0716_),
    .A(\top_inst.sndgen_inst.phacc4[10] ),
    .Y(_0747_));
 sg13g2_nor3_1 _1500_ (.A(_0714_),
    .B(\top_inst.sndgen_inst.phacc4[9] ),
    .C(\top_inst.sndgen_inst.phacc4[10] ),
    .Y(_0748_));
 sg13g2_nand2_1 _1501_ (.Y(_0749_),
    .A(_0400_),
    .B(_0748_));
 sg13g2_nor2_1 _1502_ (.A(_0719_),
    .B(_0733_),
    .Y(_0750_));
 sg13g2_inv_1 _1503_ (.Y(_0751_),
    .A(\top_inst.sndgen_inst.p_c4[7] ));
 sg13g2_nor3_1 _1504_ (.A(_0751_),
    .B(net29),
    .C(_0000_),
    .Y(_0752_));
 sg13g2_nor2_1 _1505_ (.A(\top_inst.sndgen_inst.p_c4[7] ),
    .B(_0000_),
    .Y(_0753_));
 sg13g2_nand2_1 _1506_ (.Y(_0754_),
    .A(_0532_),
    .B(_0718_));
 sg13g2_nor3_1 _1507_ (.A(net29),
    .B(_0000_),
    .C(_0754_),
    .Y(_0755_));
 sg13g2_a21oi_1 _1508_ (.A1(net29),
    .A2(\top_inst.sndgen_inst.phacc4[8] ),
    .Y(_0756_),
    .B1(_0755_));
 sg13g2_nor2_1 _1509_ (.A(_0751_),
    .B(_0756_),
    .Y(_0757_));
 sg13g2_a221oi_1 _1510_ (.B2(_0743_),
    .C1(_0757_),
    .B1(_0753_),
    .A1(_0750_),
    .Y(_0758_),
    .A2(_0752_));
 sg13g2_buf_1 _1511_ (.A(_0758_),
    .X(_0759_));
 sg13g2_mux2_1 _1512_ (.A0(_0747_),
    .A1(_0749_),
    .S(_0759_),
    .X(_0760_));
 sg13g2_xnor2_1 _1513_ (.Y(_0106_),
    .A(\top_inst.sndgen_inst.phacc4[11] ),
    .B(_0760_));
 sg13g2_or2_1 _1514_ (.X(_0761_),
    .B(_0749_),
    .A(\top_inst.sndgen_inst.phacc4[11] ));
 sg13g2_nand4_1 _1515_ (.B(\top_inst.sndgen_inst.phacc4[11] ),
    .C(net22),
    .A(\top_inst.sndgen_inst.phacc4[10] ),
    .Y(_0762_),
    .D(_0716_));
 sg13g2_mux2_1 _1516_ (.A0(_0761_),
    .A1(_0762_),
    .S(_0745_),
    .X(_0763_));
 sg13g2_xnor2_1 _1517_ (.Y(_0107_),
    .A(\top_inst.sndgen_inst.phacc4[12] ),
    .B(_0763_));
 sg13g2_buf_2 _1518_ (.A(\top_inst.sndgen_inst.phacc4[13] ),
    .X(_0764_));
 sg13g2_nor3_1 _1519_ (.A(\top_inst.sndgen_inst.phacc4[11] ),
    .B(\top_inst.sndgen_inst.phacc4[12] ),
    .C(_0749_),
    .Y(_0765_));
 sg13g2_nand2_1 _1520_ (.Y(_0766_),
    .A(\top_inst.sndgen_inst.phacc4[11] ),
    .B(\top_inst.sndgen_inst.phacc4[12] ));
 sg13g2_nor3_1 _1521_ (.A(_0759_),
    .B(_0747_),
    .C(_0766_),
    .Y(_0767_));
 sg13g2_a21o_1 _1522_ (.A2(_0765_),
    .A1(_0759_),
    .B1(_0767_),
    .X(_0768_));
 sg13g2_xor2_1 _1523_ (.B(_0768_),
    .A(_0764_),
    .X(_0108_));
 sg13g2_nand2_1 _1524_ (.Y(_0769_),
    .A(\top_inst.sndgen_inst.p_c4[0] ),
    .B(\top_inst.sndgen_inst.phacc4[0] ));
 sg13g2_xnor2_1 _1525_ (.Y(_0770_),
    .A(_0527_),
    .B(_0769_));
 sg13g2_nor2_1 _1526_ (.A(net13),
    .B(_0770_),
    .Y(_0771_));
 sg13g2_xor2_1 _1527_ (.B(_0771_),
    .A(\top_inst.sndgen_inst.phacc4[1] ),
    .X(_0109_));
 sg13g2_xnor2_1 _1528_ (.Y(_0772_),
    .A(\top_inst.sndgen_inst.p_c4[2] ),
    .B(_0722_));
 sg13g2_nor2_1 _1529_ (.A(net13),
    .B(_0772_),
    .Y(_0773_));
 sg13g2_xor2_1 _1530_ (.B(_0773_),
    .A(\top_inst.sndgen_inst.phacc4[2] ),
    .X(_0110_));
 sg13g2_and2_1 _1531_ (.A(\top_inst.sndgen_inst.p_c4[2] ),
    .B(\top_inst.sndgen_inst.phacc4[2] ),
    .X(_0774_));
 sg13g2_a21o_1 _1532_ (.A2(_0723_),
    .A1(_0722_),
    .B1(_0774_),
    .X(_0775_));
 sg13g2_xnor2_1 _1533_ (.Y(_0776_),
    .A(\top_inst.sndgen_inst.p_c4[3] ),
    .B(_0775_));
 sg13g2_nor2_1 _1534_ (.A(_0695_),
    .B(_0776_),
    .Y(_0777_));
 sg13g2_xor2_1 _1535_ (.B(_0777_),
    .A(\top_inst.sndgen_inst.phacc4[3] ),
    .X(_0111_));
 sg13g2_nor2_1 _1536_ (.A(\top_inst.sndgen_inst.phacc4[3] ),
    .B(_0775_),
    .Y(_0778_));
 sg13g2_a21oi_1 _1537_ (.A1(\top_inst.sndgen_inst.phacc4[3] ),
    .A2(_0775_),
    .Y(_0779_),
    .B1(\top_inst.sndgen_inst.p_c4[3] ));
 sg13g2_nor2_1 _1538_ (.A(_0778_),
    .B(_0779_),
    .Y(_0780_));
 sg13g2_xnor2_1 _1539_ (.Y(_0781_),
    .A(\top_inst.sndgen_inst.p_c4[4] ),
    .B(_0780_));
 sg13g2_nor2_1 _1540_ (.A(_0695_),
    .B(_0781_),
    .Y(_0782_));
 sg13g2_xor2_1 _1541_ (.B(_0782_),
    .A(\top_inst.sndgen_inst.phacc4[4] ),
    .X(_0112_));
 sg13g2_xnor2_1 _1542_ (.Y(_0783_),
    .A(\top_inst.sndgen_inst.p_c4[5] ),
    .B(_0737_));
 sg13g2_nor2_1 _1543_ (.A(net17),
    .B(_0783_),
    .Y(_0784_));
 sg13g2_xnor2_1 _1544_ (.Y(_0113_),
    .A(_0730_),
    .B(_0784_));
 sg13g2_xnor2_1 _1545_ (.Y(_0785_),
    .A(_0532_),
    .B(_0733_));
 sg13g2_nand2_1 _1546_ (.Y(_0786_),
    .A(_0622_),
    .B(_0785_));
 sg13g2_xnor2_1 _1547_ (.Y(_0114_),
    .A(_0718_),
    .B(_0786_));
 sg13g2_a21oi_1 _1548_ (.A1(_0532_),
    .A2(_0718_),
    .Y(_0787_),
    .B1(_0750_));
 sg13g2_xnor2_1 _1549_ (.Y(_0788_),
    .A(_0751_),
    .B(_0787_));
 sg13g2_nor2_1 _1550_ (.A(net13),
    .B(_0788_),
    .Y(_0789_));
 sg13g2_xor2_1 _1551_ (.B(_0789_),
    .A(_0734_),
    .X(_0115_));
 sg13g2_xnor2_1 _1552_ (.Y(_0790_),
    .A(_0000_),
    .B(_0744_));
 sg13g2_nand2_1 _1553_ (.Y(_0791_),
    .A(\top_inst.sndgen_inst.phacc4[8] ),
    .B(net15));
 sg13g2_o21ai_1 _1554_ (.B1(_0791_),
    .Y(_0116_),
    .A1(net15),
    .A2(_0790_));
 sg13g2_xnor2_1 _1555_ (.Y(_0792_),
    .A(\top_inst.sndgen_inst.p_c4[10] ),
    .B(_0759_));
 sg13g2_nand2_1 _1556_ (.Y(_0793_),
    .A(net22),
    .B(_0792_));
 sg13g2_xnor2_1 _1557_ (.Y(_0117_),
    .A(\top_inst.sndgen_inst.phacc4[9] ),
    .B(_0793_));
 sg13g2_nor2_2 _1558_ (.A(_0477_),
    .B(_0513_),
    .Y(_0794_));
 sg13g2_nor2_1 _1559_ (.A(_0475_),
    .B(_0451_),
    .Y(_0795_));
 sg13g2_a21oi_1 _1560_ (.A1(\top_inst.sndgen_inst.c2[0] ),
    .A2(net14),
    .Y(_0796_),
    .B1(_0795_));
 sg13g2_nor2_1 _1561_ (.A(\top_inst.sndgen_inst.c3[0] ),
    .B(_0794_),
    .Y(_0797_));
 sg13g2_a21oi_1 _1562_ (.A1(_0794_),
    .A2(_0796_),
    .Y(_0118_),
    .B1(_0797_));
 sg13g2_nor2_1 _1563_ (.A(_0500_),
    .B(_0451_),
    .Y(_0798_));
 sg13g2_a21oi_1 _1564_ (.A1(\top_inst.sndgen_inst.c2[1] ),
    .A2(net14),
    .Y(_0799_),
    .B1(_0798_));
 sg13g2_nor2_1 _1565_ (.A(\top_inst.sndgen_inst.c3[1] ),
    .B(_0794_),
    .Y(_0800_));
 sg13g2_a21oi_1 _1566_ (.A1(_0794_),
    .A2(_0799_),
    .Y(_0119_),
    .B1(_0800_));
 sg13g2_nand2_1 _1567_ (.Y(_0801_),
    .A(_0479_),
    .B(net21));
 sg13g2_nand2_1 _1568_ (.Y(_0802_),
    .A(\top_inst.sndgen_inst.c2[2] ),
    .B(_0451_));
 sg13g2_a21oi_1 _1569_ (.A1(_0801_),
    .A2(_0802_),
    .Y(_0803_),
    .B1(net31));
 sg13g2_a21oi_1 _1570_ (.A1(net31),
    .A2(\top_inst.sndgen_inst.c3[2] ),
    .Y(_0804_),
    .B1(_0803_));
 sg13g2_nand2_1 _1571_ (.Y(_0805_),
    .A(net25),
    .B(\top_inst.sndgen_inst.c4[2] ));
 sg13g2_o21ai_1 _1572_ (.B1(_0805_),
    .Y(_0120_),
    .A1(net25),
    .A2(_0804_));
 sg13g2_nand2_1 _1573_ (.Y(_0806_),
    .A(_0471_),
    .B(_0794_));
 sg13g2_nand2_1 _1574_ (.Y(_0807_),
    .A(net25),
    .B(\top_inst.sndgen_inst.c3[2] ));
 sg13g2_o21ai_1 _1575_ (.B1(_0807_),
    .Y(_0121_),
    .A1(net16),
    .A2(_0806_));
 sg13g2_mux2_1 _1576_ (.A0(_0426_),
    .A1(_0019_),
    .S(net14),
    .X(_0122_));
 sg13g2_xnor2_1 _1577_ (.Y(_0123_),
    .A(\top_inst.sndgen_inst.slot_counter[10] ),
    .B(_0429_));
 sg13g2_nand3_1 _1578_ (.B(_0411_),
    .C(_0451_),
    .A(_0426_),
    .Y(_0808_));
 sg13g2_nor3_2 _1579_ (.A(_0406_),
    .B(_0407_),
    .C(_0808_),
    .Y(_0809_));
 sg13g2_xor2_1 _1580_ (.B(_0809_),
    .A(_0416_),
    .X(_0124_));
 sg13g2_nand2_1 _1581_ (.Y(_0810_),
    .A(_0416_),
    .B(_0809_));
 sg13g2_xnor2_1 _1582_ (.Y(_0125_),
    .A(_0419_),
    .B(_0810_));
 sg13g2_nand2b_1 _1583_ (.Y(_0811_),
    .B(_0809_),
    .A_N(_0425_));
 sg13g2_xnor2_1 _1584_ (.Y(_0126_),
    .A(_0417_),
    .B(_0811_));
 sg13g2_nand4_1 _1585_ (.B(_0416_),
    .C(_0417_),
    .A(_0419_),
    .Y(_0812_),
    .D(_0809_));
 sg13g2_xnor2_1 _1586_ (.Y(_0127_),
    .A(\top_inst.sndgen_inst.bar_counter[3] ),
    .B(_0812_));
 sg13g2_nand2_1 _1587_ (.Y(_0813_),
    .A(_0426_),
    .B(\top_inst.sample_ena ));
 sg13g2_xnor2_1 _1588_ (.Y(_0128_),
    .A(net35),
    .B(_0813_));
 sg13g2_nand3_1 _1589_ (.B(_0426_),
    .C(net14),
    .A(net35),
    .Y(_0814_));
 sg13g2_xnor2_1 _1590_ (.Y(_0129_),
    .A(\top_inst.sndgen_inst.slot_counter[2] ),
    .B(_0814_));
 sg13g2_nand4_1 _1591_ (.B(_0426_),
    .C(\top_inst.sndgen_inst.slot_counter[2] ),
    .A(net35),
    .Y(_0815_),
    .D(net14));
 sg13g2_xnor2_1 _1592_ (.Y(_0130_),
    .A(\top_inst.sndgen_inst.slot_counter[3] ),
    .B(_0815_));
 sg13g2_xnor2_1 _1593_ (.Y(_0131_),
    .A(\top_inst.sndgen_inst.slot_counter[4] ),
    .B(_0808_));
 sg13g2_and3_1 _1594_ (.X(_0816_),
    .A(_0426_),
    .B(_0411_),
    .C(_0451_));
 sg13g2_buf_1 _1595_ (.A(_0816_),
    .X(_0817_));
 sg13g2_nand2_1 _1596_ (.Y(_0818_),
    .A(\top_inst.sndgen_inst.slot_counter[4] ),
    .B(_0817_));
 sg13g2_xnor2_1 _1597_ (.Y(_0132_),
    .A(\top_inst.sndgen_inst.slot_counter[5] ),
    .B(_0818_));
 sg13g2_nand3_1 _1598_ (.B(\top_inst.sndgen_inst.slot_counter[4] ),
    .C(_0817_),
    .A(\top_inst.sndgen_inst.slot_counter[5] ),
    .Y(_0819_));
 sg13g2_xnor2_1 _1599_ (.Y(_0133_),
    .A(\top_inst.sndgen_inst.slot_counter[6] ),
    .B(_0819_));
 sg13g2_nand2_1 _1600_ (.Y(_0820_),
    .A(_0405_),
    .B(_0817_));
 sg13g2_xnor2_1 _1601_ (.Y(_0134_),
    .A(\top_inst.sndgen_inst.slot_counter[7] ),
    .B(_0820_));
 sg13g2_nand3_1 _1602_ (.B(_0405_),
    .C(_0817_),
    .A(\top_inst.sndgen_inst.slot_counter[7] ),
    .Y(_0821_));
 sg13g2_xnor2_1 _1603_ (.Y(_0135_),
    .A(\top_inst.sndgen_inst.slot_counter[8] ),
    .B(_0821_));
 sg13g2_xor2_1 _1604_ (.B(_0428_),
    .A(\top_inst.sndgen_inst.slot_counter[9] ),
    .X(_0136_));
 sg13g2_inv_1 _1605_ (.Y(_0822_),
    .A(\top_inst.vga_inst.sx1[0] ));
 sg13g2_nand2_1 _1606_ (.Y(_0823_),
    .A(\top_inst.vga_inst.sr1[0] ),
    .B(net15));
 sg13g2_o21ai_1 _1607_ (.B1(_0823_),
    .Y(_0137_),
    .A1(_0822_),
    .A2(_0453_));
 sg13g2_mux2_1 _1608_ (.A0(\top_inst.vga_inst.sx1[1] ),
    .A1(\top_inst.vga_inst.sr1[1] ),
    .S(net17),
    .X(_0138_));
 sg13g2_mux2_1 _1609_ (.A0(\top_inst.vga_inst.sx1[2] ),
    .A1(\top_inst.vga_inst.sr1[2] ),
    .S(net17),
    .X(_0139_));
 sg13g2_inv_1 _1610_ (.Y(_0824_),
    .A(\top_inst.vga_inst.sx1[3] ));
 sg13g2_nand2_1 _1611_ (.Y(_0825_),
    .A(\top_inst.vga_inst.sr1[3] ),
    .B(net17));
 sg13g2_o21ai_1 _1612_ (.B1(_0825_),
    .Y(_0140_),
    .A1(_0824_),
    .A2(_0453_));
 sg13g2_nor2_1 _1613_ (.A(\top_inst.sndgen_inst.slot_counter[6] ),
    .B(_0002_),
    .Y(_0826_));
 sg13g2_nor4_1 _1614_ (.A(\top_inst.sndgen_inst.slot_counter[3] ),
    .B(\top_inst.sndgen_inst.slot_counter[2] ),
    .C(\top_inst.sndgen_inst.slot_counter[8] ),
    .D(\top_inst.sndgen_inst.slot_counter[7] ),
    .Y(_0827_));
 sg13g2_nor4_1 _1615_ (.A(net35),
    .B(_0426_),
    .C(\top_inst.sndgen_inst.slot_counter[5] ),
    .D(\top_inst.sndgen_inst.slot_counter[4] ),
    .Y(_0828_));
 sg13g2_nand3_1 _1616_ (.B(_0827_),
    .C(_0828_),
    .A(_0826_),
    .Y(_0829_));
 sg13g2_nand2_2 _1617_ (.Y(_0830_),
    .A(_0408_),
    .B(_0829_));
 sg13g2_buf_2 _1618_ (.A(_0012_),
    .X(_0831_));
 sg13g2_nand2_1 _1619_ (.Y(_0832_),
    .A(_0435_),
    .B(\top_inst.sndgen_inst.c1[1] ));
 sg13g2_nand3b_1 _1620_ (.B(\top_inst.sndgen_inst.c1[0] ),
    .C(net34),
    .Y(_0833_),
    .A_N(\top_inst.sndgen_inst.c1[1] ));
 sg13g2_nor2_1 _1621_ (.A(\top_inst.sndgen_inst.mask_1[0] ),
    .B(\top_inst.sndgen_inst.mask_2 ),
    .Y(_0834_));
 sg13g2_a21oi_2 _1622_ (.B1(_0834_),
    .Y(_0835_),
    .A2(_0833_),
    .A1(_0832_));
 sg13g2_xnor2_1 _1623_ (.Y(_0836_),
    .A(_0831_),
    .B(_0835_));
 sg13g2_nand2_1 _1624_ (.Y(_0837_),
    .A(_0830_),
    .B(_0836_));
 sg13g2_xnor2_1 _1625_ (.Y(_0838_),
    .A(_0464_),
    .B(_0837_));
 sg13g2_nand2_1 _1626_ (.Y(_0839_),
    .A(_0467_),
    .B(_0838_));
 sg13g2_xnor2_1 _1627_ (.Y(_0840_),
    .A(_0463_),
    .B(_0837_));
 sg13g2_nand2_1 _1628_ (.Y(_0841_),
    .A(net33),
    .B(_0840_));
 sg13g2_nand3_1 _1629_ (.B(_0839_),
    .C(_0841_),
    .A(net14),
    .Y(_0842_));
 sg13g2_o21ai_1 _1630_ (.B1(_0842_),
    .Y(_0141_),
    .A1(_0822_),
    .A2(_0452_));
 sg13g2_nand2_1 _1631_ (.Y(_0843_),
    .A(_0831_),
    .B(_0464_));
 sg13g2_inv_1 _1632_ (.Y(_0844_),
    .A(_0831_));
 sg13g2_nor2_1 _1633_ (.A(_0844_),
    .B(_0679_),
    .Y(_0845_));
 sg13g2_a21o_1 _1634_ (.A2(_0833_),
    .A1(_0832_),
    .B1(_0834_),
    .X(_0846_));
 sg13g2_o21ai_1 _1635_ (.B1(_0846_),
    .Y(_0847_),
    .A1(_0464_),
    .A2(_0845_));
 sg13g2_nand2b_1 _1636_ (.Y(_0848_),
    .B(\top_inst.sndgen_inst.c1[1] ),
    .A_N(net34));
 sg13g2_nand2b_1 _1637_ (.Y(_0849_),
    .B(\top_inst.sndgen_inst.c1[0] ),
    .A_N(\top_inst.sndgen_inst.c1[1] ));
 sg13g2_a21oi_1 _1638_ (.A1(_0848_),
    .A2(_0849_),
    .Y(_0850_),
    .B1(_0834_));
 sg13g2_buf_1 _1639_ (.A(_0850_),
    .X(_0851_));
 sg13g2_nor2_2 _1640_ (.A(_0831_),
    .B(\top_inst.sndgen_inst.phacc2[13] ),
    .Y(_0852_));
 sg13g2_xnor2_1 _1641_ (.Y(_0853_),
    .A(net23),
    .B(_0852_));
 sg13g2_a221oi_1 _1642_ (.B2(_0847_),
    .C1(_0853_),
    .B1(_0843_),
    .A1(_0408_),
    .Y(_0854_),
    .A2(_0829_));
 sg13g2_nand2_1 _1643_ (.Y(_0855_),
    .A(_0463_),
    .B(_0679_));
 sg13g2_nor2_1 _1644_ (.A(_0830_),
    .B(_0855_),
    .Y(_0856_));
 sg13g2_nor2_1 _1645_ (.A(_0464_),
    .B(\top_inst.sndgen_inst.phacc3[13] ),
    .Y(_0857_));
 sg13g2_o21ai_1 _1646_ (.B1(_0857_),
    .Y(_0858_),
    .A1(_0844_),
    .A2(_0835_));
 sg13g2_or4_1 _1647_ (.A(_0844_),
    .B(_0835_),
    .C(net23),
    .D(_0855_),
    .X(_0859_));
 sg13g2_o21ai_1 _1648_ (.B1(_0859_),
    .Y(_0860_),
    .A1(_0853_),
    .A2(_0858_));
 sg13g2_nor2_1 _1649_ (.A(_0464_),
    .B(_0679_),
    .Y(_0861_));
 sg13g2_nand2_1 _1650_ (.Y(_0862_),
    .A(_0844_),
    .B(_0861_));
 sg13g2_nor2_1 _1651_ (.A(_0831_),
    .B(_0463_),
    .Y(_0863_));
 sg13g2_o21ai_1 _1652_ (.B1(_0835_),
    .Y(_0864_),
    .A1(_0863_),
    .A2(_0861_));
 sg13g2_xor2_1 _1653_ (.B(_0852_),
    .A(net23),
    .X(_0865_));
 sg13g2_a221oi_1 _1654_ (.B2(_0864_),
    .C1(_0865_),
    .B1(_0862_),
    .A1(_0408_),
    .Y(_0866_),
    .A2(_0829_));
 sg13g2_or4_1 _1655_ (.A(_0854_),
    .B(_0856_),
    .C(_0860_),
    .D(_0866_),
    .X(_0867_));
 sg13g2_buf_2 _1656_ (.A(_0867_),
    .X(_0868_));
 sg13g2_xnor2_1 _1657_ (.Y(_0869_),
    .A(_0764_),
    .B(_0838_));
 sg13g2_nor2_1 _1658_ (.A(_0467_),
    .B(_0869_),
    .Y(_0870_));
 sg13g2_xnor2_1 _1659_ (.Y(_0871_),
    .A(_0868_),
    .B(_0870_));
 sg13g2_nand2_1 _1660_ (.Y(_0872_),
    .A(\top_inst.vga_inst.sx1[1] ),
    .B(_0449_));
 sg13g2_o21ai_1 _1661_ (.B1(_0872_),
    .Y(_0142_),
    .A1(net15),
    .A2(_0871_));
 sg13g2_o21ai_1 _1662_ (.B1(_0852_),
    .Y(_0873_),
    .A1(_0851_),
    .A2(_0857_));
 sg13g2_nand2_1 _1663_ (.Y(_0874_),
    .A(net23),
    .B(_0857_));
 sg13g2_a22oi_1 _1664_ (.Y(_0875_),
    .B1(_0873_),
    .B2(_0874_),
    .A2(_0829_),
    .A1(_0408_));
 sg13g2_buf_1 _1665_ (.A(_0875_),
    .X(_0876_));
 sg13g2_nor3_1 _1666_ (.A(_0679_),
    .B(net23),
    .C(_0852_),
    .Y(_0877_));
 sg13g2_nor2_1 _1667_ (.A(\top_inst.sndgen_inst.phacc3[13] ),
    .B(_0852_),
    .Y(_0878_));
 sg13g2_and2_1 _1668_ (.A(net23),
    .B(_0878_),
    .X(_0879_));
 sg13g2_nor4_1 _1669_ (.A(_0831_),
    .B(\top_inst.sndgen_inst.phacc2[13] ),
    .C(\top_inst.sndgen_inst.phacc3[13] ),
    .D(net23),
    .Y(_0880_));
 sg13g2_and3_1 _1670_ (.X(_0881_),
    .A(\top_inst.sndgen_inst.phacc3[13] ),
    .B(net23),
    .C(_0852_));
 sg13g2_nor4_1 _1671_ (.A(_0877_),
    .B(_0879_),
    .C(_0880_),
    .D(_0881_),
    .Y(_0882_));
 sg13g2_a21oi_1 _1672_ (.A1(_0831_),
    .A2(_0846_),
    .Y(_0883_),
    .B1(_0464_));
 sg13g2_nand2_1 _1673_ (.Y(_0884_),
    .A(_0830_),
    .B(_0883_));
 sg13g2_nand4_1 _1674_ (.B(_0835_),
    .C(_0853_),
    .A(_0830_),
    .Y(_0885_),
    .D(_0863_));
 sg13g2_o21ai_1 _1675_ (.B1(_0885_),
    .Y(_0886_),
    .A1(_0882_),
    .A2(_0884_));
 sg13g2_nand2b_1 _1676_ (.Y(_0887_),
    .B(net33),
    .A_N(_0764_));
 sg13g2_o21ai_1 _1677_ (.B1(_0859_),
    .Y(_0888_),
    .A1(_0830_),
    .A2(_0855_));
 sg13g2_nor2_1 _1678_ (.A(_0854_),
    .B(_0888_),
    .Y(_0889_));
 sg13g2_o21ai_1 _1679_ (.B1(_0889_),
    .Y(_0890_),
    .A1(_0886_),
    .A2(_0887_));
 sg13g2_and2_1 _1680_ (.A(net33),
    .B(_0764_),
    .X(_0891_));
 sg13g2_xnor2_1 _1681_ (.Y(_0892_),
    .A(_0464_),
    .B(_0836_));
 sg13g2_and2_1 _1682_ (.A(_0891_),
    .B(_0892_),
    .X(_0893_));
 sg13g2_nor2_1 _1683_ (.A(_0889_),
    .B(_0887_),
    .Y(_0894_));
 sg13g2_a221oi_1 _1684_ (.B2(_0886_),
    .C1(_0894_),
    .B1(_0893_),
    .A1(_0841_),
    .Y(_0895_),
    .A2(_0890_));
 sg13g2_xnor2_1 _1685_ (.Y(_0896_),
    .A(_0876_),
    .B(_0895_));
 sg13g2_mux2_1 _1686_ (.A0(\top_inst.vga_inst.sx1[2] ),
    .A1(_0896_),
    .S(net14),
    .X(_0143_));
 sg13g2_nor2b_1 _1687_ (.A(_0886_),
    .B_N(_0876_),
    .Y(_0897_));
 sg13g2_nand2b_1 _1688_ (.Y(_0898_),
    .B(_0889_),
    .A_N(_0876_));
 sg13g2_o21ai_1 _1689_ (.B1(_0898_),
    .Y(_0899_),
    .A1(_0841_),
    .A2(_0897_));
 sg13g2_inv_1 _1690_ (.Y(_0900_),
    .A(_0886_));
 sg13g2_o21ai_1 _1691_ (.B1(_0889_),
    .Y(_0901_),
    .A1(_0467_),
    .A2(_0840_));
 sg13g2_a21oi_1 _1692_ (.A1(_0900_),
    .A2(_0901_),
    .Y(_0902_),
    .B1(_0876_));
 sg13g2_a21o_1 _1693_ (.A2(_0899_),
    .A1(_0764_),
    .B1(_0902_),
    .X(_0903_));
 sg13g2_nand2_1 _1694_ (.Y(_0904_),
    .A(net16),
    .B(_0903_));
 sg13g2_o21ai_1 _1695_ (.B1(_0904_),
    .Y(_0144_),
    .A1(_0824_),
    .A2(_0452_));
 sg13g2_buf_1 _1696_ (.A(\top_inst.vga_inst.x[8] ),
    .X(_0905_));
 sg13g2_inv_1 _1697_ (.Y(_0181_),
    .A(_0398_));
 sg13g2_nand2_1 _1698_ (.Y(_0182_),
    .A(_0395_),
    .B(_0387_));
 sg13g2_nor2_1 _1699_ (.A(_0392_),
    .B(_0182_),
    .Y(_0183_));
 sg13g2_nor4_1 _1700_ (.A(net37),
    .B(net28),
    .C(_0181_),
    .D(_0183_),
    .Y(_0184_));
 sg13g2_buf_1 _1701_ (.A(_0184_),
    .X(_0185_));
 sg13g2_xnor2_1 _1702_ (.Y(_0186_),
    .A(_0401_),
    .B(\top_inst.vga_inst.x1[0] ));
 sg13g2_nor2_1 _1703_ (.A(net20),
    .B(_0186_),
    .Y(_0145_));
 sg13g2_nand2_1 _1704_ (.Y(_0187_),
    .A(_0398_),
    .B(\top_inst.vga_inst.x1[0] ));
 sg13g2_xor2_1 _1705_ (.B(_0187_),
    .A(\top_inst.vga_inst.x1[1] ),
    .X(_0188_));
 sg13g2_nor2_1 _1706_ (.A(net20),
    .B(_0188_),
    .Y(_0146_));
 sg13g2_inv_1 _1707_ (.Y(_0189_),
    .A(\top_inst.vga_inst.x1[2] ));
 sg13g2_nand3_1 _1708_ (.B(\top_inst.vga_inst.x1[0] ),
    .C(\top_inst.vga_inst.x1[1] ),
    .A(_0398_),
    .Y(_0190_));
 sg13g2_xnor2_1 _1709_ (.Y(_0191_),
    .A(_0189_),
    .B(_0190_));
 sg13g2_nor2_1 _1710_ (.A(net20),
    .B(_0191_),
    .Y(_0147_));
 sg13g2_nor2_2 _1711_ (.A(_0189_),
    .B(_0190_),
    .Y(_0192_));
 sg13g2_xnor2_1 _1712_ (.Y(_0193_),
    .A(\top_inst.vga_inst.x1[3] ),
    .B(_0192_));
 sg13g2_nor2_1 _1713_ (.A(net20),
    .B(_0193_),
    .Y(_0148_));
 sg13g2_buf_1 _1714_ (.A(\top_inst.vga_inst.x1[4] ),
    .X(_0194_));
 sg13g2_nand2_1 _1715_ (.Y(_0195_),
    .A(\top_inst.vga_inst.x1[3] ),
    .B(_0192_));
 sg13g2_xor2_1 _1716_ (.B(_0195_),
    .A(_0194_),
    .X(_0196_));
 sg13g2_nor2_1 _1717_ (.A(net20),
    .B(_0196_),
    .Y(_0149_));
 sg13g2_buf_2 _1718_ (.A(\top_inst.vga_inst.x1[5] ),
    .X(_0197_));
 sg13g2_nand3_1 _1719_ (.B(_0194_),
    .C(_0192_),
    .A(\top_inst.vga_inst.x1[3] ),
    .Y(_0198_));
 sg13g2_xor2_1 _1720_ (.B(_0198_),
    .A(_0197_),
    .X(_0199_));
 sg13g2_nor2_1 _1721_ (.A(_0185_),
    .B(_0199_),
    .Y(_0150_));
 sg13g2_inv_1 _1722_ (.Y(_0200_),
    .A(\top_inst.vga_inst.x1[6] ));
 sg13g2_nand4_1 _1723_ (.B(_0194_),
    .C(_0197_),
    .A(\top_inst.vga_inst.x1[3] ),
    .Y(_0201_),
    .D(_0192_));
 sg13g2_xnor2_1 _1724_ (.Y(_0202_),
    .A(_0200_),
    .B(_0201_));
 sg13g2_nor2_1 _1725_ (.A(_0185_),
    .B(_0202_),
    .Y(_0151_));
 sg13g2_nor2_1 _1726_ (.A(_0200_),
    .B(_0201_),
    .Y(_0203_));
 sg13g2_xnor2_1 _1727_ (.Y(_0204_),
    .A(\top_inst.vga_inst.x1[7] ),
    .B(_0203_));
 sg13g2_nor2_1 _1728_ (.A(net20),
    .B(_0204_),
    .Y(_0152_));
 sg13g2_xor2_1 _1729_ (.B(net27),
    .A(_0388_),
    .X(_0153_));
 sg13g2_nand2_1 _1730_ (.Y(_0205_),
    .A(_0388_),
    .B(net27));
 sg13g2_xnor2_1 _1731_ (.Y(_0154_),
    .A(\top_inst.vga_inst.x[1] ),
    .B(_0205_));
 sg13g2_nand3_1 _1732_ (.B(_0388_),
    .C(net27),
    .A(\top_inst.vga_inst.x[1] ),
    .Y(_0206_));
 sg13g2_xnor2_1 _1733_ (.Y(_0155_),
    .A(\top_inst.vga_inst.x[2] ),
    .B(_0206_));
 sg13g2_nand4_1 _1734_ (.B(\top_inst.vga_inst.x[1] ),
    .C(_0388_),
    .A(\top_inst.vga_inst.x[2] ),
    .Y(_0207_),
    .D(net27));
 sg13g2_xnor2_1 _1735_ (.Y(_0156_),
    .A(\top_inst.vga_inst.x[3] ),
    .B(_0207_));
 sg13g2_and4_1 _1736_ (.A(\top_inst.vga_inst.x[3] ),
    .B(\top_inst.vga_inst.x[2] ),
    .C(\top_inst.vga_inst.x[1] ),
    .D(_0388_),
    .X(_0208_));
 sg13g2_and2_1 _1737_ (.A(_0398_),
    .B(_0208_),
    .X(_0209_));
 sg13g2_buf_2 _1738_ (.A(_0209_),
    .X(_0210_));
 sg13g2_xnor2_1 _1739_ (.Y(_0157_),
    .A(_0444_),
    .B(_0210_));
 sg13g2_nand2_1 _1740_ (.Y(_0211_),
    .A(_0390_),
    .B(_0210_));
 sg13g2_nand3_1 _1741_ (.B(\top_inst.vga_inst.x[8] ),
    .C(_0445_),
    .A(net37),
    .Y(_0212_));
 sg13g2_nor3_2 _1742_ (.A(_0444_),
    .B(_0395_),
    .C(_0212_),
    .Y(_0213_));
 sg13g2_nor3_1 _1743_ (.A(net38),
    .B(_0211_),
    .C(_0213_),
    .Y(_0214_));
 sg13g2_a21o_1 _1744_ (.A2(_0211_),
    .A1(net38),
    .B1(_0214_),
    .X(_0158_));
 sg13g2_nand3_1 _1745_ (.B(_0391_),
    .C(_0210_),
    .A(_0390_),
    .Y(_0215_));
 sg13g2_xnor2_1 _1746_ (.Y(_0159_),
    .A(_0387_),
    .B(_0215_));
 sg13g2_and3_1 _1747_ (.X(_0216_),
    .A(_0390_),
    .B(_0391_),
    .C(_0387_));
 sg13g2_buf_1 _1748_ (.A(_0216_),
    .X(_0217_));
 sg13g2_nand3_1 _1749_ (.B(_0208_),
    .C(_0217_),
    .A(_0005_),
    .Y(_0218_));
 sg13g2_o21ai_1 _1750_ (.B1(_0218_),
    .Y(_0219_),
    .A1(_0005_),
    .A2(_0217_));
 sg13g2_nand2b_1 _1751_ (.Y(_0220_),
    .B(_0219_),
    .A_N(_0213_));
 sg13g2_o21ai_1 _1752_ (.B1(_0220_),
    .Y(_0221_),
    .A1(_0005_),
    .A2(_0208_));
 sg13g2_mux2_1 _1753_ (.A0(_0395_),
    .A1(_0221_),
    .S(_0401_),
    .X(_0160_));
 sg13g2_and2_1 _1754_ (.A(_0395_),
    .B(_0387_),
    .X(_0222_));
 sg13g2_buf_1 _1755_ (.A(_0222_),
    .X(_0223_));
 sg13g2_and3_1 _1756_ (.X(_0224_),
    .A(_0390_),
    .B(net38),
    .C(_0223_));
 sg13g2_o21ai_1 _1757_ (.B1(_0210_),
    .Y(_0225_),
    .A1(_0213_),
    .A2(_0224_));
 sg13g2_nor3_1 _1758_ (.A(net28),
    .B(_0182_),
    .C(_0215_),
    .Y(_0226_));
 sg13g2_a21o_1 _1759_ (.A2(_0225_),
    .A1(net28),
    .B1(_0226_),
    .X(_0161_));
 sg13g2_and3_1 _1760_ (.X(_0227_),
    .A(_0395_),
    .B(net28),
    .C(_0217_));
 sg13g2_nand2_1 _1761_ (.Y(_0228_),
    .A(_0210_),
    .B(_0227_));
 sg13g2_o21ai_1 _1762_ (.B1(_0210_),
    .Y(_0229_),
    .A1(_0213_),
    .A2(_0227_));
 sg13g2_nand2_1 _1763_ (.Y(_0230_),
    .A(net37),
    .B(_0229_));
 sg13g2_o21ai_1 _1764_ (.B1(_0230_),
    .Y(_0162_),
    .A1(_0394_),
    .A2(_0228_));
 sg13g2_inv_1 _1765_ (.Y(_0231_),
    .A(\top_inst.vga_inst.sr1[3] ));
 sg13g2_nor2b_1 _1766_ (.A(\top_inst.vga_inst.sx1[0] ),
    .B_N(\top_inst.vga_inst.sr1[0] ),
    .Y(_0232_));
 sg13g2_nor2_1 _1767_ (.A(\top_inst.vga_inst.sr1[1] ),
    .B(_0232_),
    .Y(_0233_));
 sg13g2_nand2_1 _1768_ (.Y(_0234_),
    .A(\top_inst.vga_inst.sr1[1] ),
    .B(_0232_));
 sg13g2_o21ai_1 _1769_ (.B1(_0234_),
    .Y(_0235_),
    .A1(\top_inst.vga_inst.sx1[1] ),
    .A2(_0233_));
 sg13g2_nand2_1 _1770_ (.Y(_0236_),
    .A(\top_inst.vga_inst.sr1[2] ),
    .B(_0235_));
 sg13g2_nor2_1 _1771_ (.A(\top_inst.vga_inst.sr1[2] ),
    .B(_0235_),
    .Y(_0237_));
 sg13g2_a221oi_1 _1772_ (.B2(_0236_),
    .C1(_0237_),
    .B1(\top_inst.vga_inst.sx1[2] ),
    .A1(_0231_),
    .Y(_0238_),
    .A2(\top_inst.vga_inst.sx1[3] ));
 sg13g2_a21oi_2 _1773_ (.B1(_0238_),
    .Y(_0239_),
    .A2(_0824_),
    .A1(\top_inst.vga_inst.sr1[3] ));
 sg13g2_mux2_1 _1774_ (.A0(\top_inst.vga_inst.sr1[0] ),
    .A1(\top_inst.vga_inst.sx1[0] ),
    .S(_0239_),
    .X(_0240_));
 sg13g2_buf_1 _1775_ (.A(_0184_),
    .X(_0241_));
 sg13g2_mux2_1 _1776_ (.A0(\top_inst.vga_inst.xmax[0] ),
    .A1(_0240_),
    .S(net19),
    .X(_0163_));
 sg13g2_mux2_1 _1777_ (.A0(\top_inst.vga_inst.sr1[1] ),
    .A1(\top_inst.vga_inst.sx1[1] ),
    .S(_0239_),
    .X(_0242_));
 sg13g2_mux2_1 _1778_ (.A0(\top_inst.vga_inst.xmax[1] ),
    .A1(_0242_),
    .S(net19),
    .X(_0164_));
 sg13g2_inv_1 _1779_ (.Y(_0243_),
    .A(\top_inst.vga_inst.xmax[2] ));
 sg13g2_mux2_1 _1780_ (.A0(\top_inst.vga_inst.sr1[2] ),
    .A1(\top_inst.vga_inst.sx1[2] ),
    .S(_0239_),
    .X(_0244_));
 sg13g2_nand2_1 _1781_ (.Y(_0245_),
    .A(net19),
    .B(_0244_));
 sg13g2_o21ai_1 _1782_ (.B1(_0245_),
    .Y(_0165_),
    .A1(_0243_),
    .A2(net20));
 sg13g2_inv_1 _1783_ (.Y(_0246_),
    .A(\top_inst.vga_inst.xmax[3] ));
 sg13g2_o21ai_1 _1784_ (.B1(net19),
    .Y(_0247_),
    .A1(\top_inst.vga_inst.sr1[3] ),
    .A2(\top_inst.vga_inst.sx1[3] ));
 sg13g2_o21ai_1 _1785_ (.B1(_0247_),
    .Y(_0166_),
    .A1(_0246_),
    .A2(net20));
 sg13g2_mux2_1 _1786_ (.A0(\top_inst.vga_inst.sx1[0] ),
    .A1(\top_inst.vga_inst.sr1[0] ),
    .S(_0239_),
    .X(_0248_));
 sg13g2_mux2_1 _1787_ (.A0(\top_inst.vga_inst.xmin[0] ),
    .A1(_0248_),
    .S(_0241_),
    .X(_0167_));
 sg13g2_mux2_1 _1788_ (.A0(\top_inst.vga_inst.sx1[1] ),
    .A1(\top_inst.vga_inst.sr1[1] ),
    .S(_0239_),
    .X(_0249_));
 sg13g2_mux2_1 _1789_ (.A0(\top_inst.vga_inst.xmin[1] ),
    .A1(_0249_),
    .S(_0241_),
    .X(_0168_));
 sg13g2_inv_1 _1790_ (.Y(_0250_),
    .A(\top_inst.vga_inst.xmin[2] ));
 sg13g2_mux2_1 _1791_ (.A0(\top_inst.vga_inst.sx1[2] ),
    .A1(\top_inst.vga_inst.sr1[2] ),
    .S(_0239_),
    .X(_0251_));
 sg13g2_nand2_1 _1792_ (.Y(_0252_),
    .A(net19),
    .B(_0251_));
 sg13g2_o21ai_1 _1793_ (.B1(_0252_),
    .Y(_0169_),
    .A1(_0250_),
    .A2(net19));
 sg13g2_inv_1 _1794_ (.Y(_0253_),
    .A(\top_inst.vga_inst.xmin[3] ));
 sg13g2_nand3_1 _1795_ (.B(\top_inst.vga_inst.sx1[3] ),
    .C(net19),
    .A(\top_inst.vga_inst.sr1[3] ),
    .Y(_0254_));
 sg13g2_o21ai_1 _1796_ (.B1(_0254_),
    .Y(_0170_),
    .A1(_0253_),
    .A2(net19));
 sg13g2_buf_2 _1797_ (.A(\top_inst.vga_inst.y[2] ),
    .X(_0255_));
 sg13g2_buf_2 _1798_ (.A(\top_inst.vga_inst.y[9] ),
    .X(_0256_));
 sg13g2_buf_1 _1799_ (.A(\top_inst.vga_inst.y[7] ),
    .X(_0257_));
 sg13g2_buf_1 _1800_ (.A(\top_inst.vga_inst.bg[4] ),
    .X(_0258_));
 sg13g2_nor4_1 _1801_ (.A(_0257_),
    .B(\top_inst.vga_inst.bg[5] ),
    .C(_0258_),
    .D(\top_inst.vga_inst.y[8] ),
    .Y(_0259_));
 sg13g2_buf_2 _1802_ (.A(\top_inst.vga_inst.y[1] ),
    .X(_0260_));
 sg13g2_buf_2 _1803_ (.A(\top_inst.vga_inst.bg[0] ),
    .X(_0261_));
 sg13g2_buf_2 _1804_ (.A(\top_inst.vga_inst.bg[1] ),
    .X(_0262_));
 sg13g2_inv_1 _1805_ (.Y(_0263_),
    .A(_0262_));
 sg13g2_nand2_1 _1806_ (.Y(_0264_),
    .A(_0261_),
    .B(_0263_));
 sg13g2_nor3_1 _1807_ (.A(net36),
    .B(_0260_),
    .C(_0264_),
    .Y(_0265_));
 sg13g2_and4_1 _1808_ (.A(_0255_),
    .B(_0256_),
    .C(_0259_),
    .D(_0265_),
    .X(_0266_));
 sg13g2_buf_1 _1809_ (.A(_0266_),
    .X(_0267_));
 sg13g2_and2_1 _1810_ (.A(_0210_),
    .B(_0213_),
    .X(_0268_));
 sg13g2_nand2b_2 _1811_ (.Y(_0269_),
    .B(_0268_),
    .A_N(_0267_));
 sg13g2_nand2_1 _1812_ (.Y(_0270_),
    .A(_0210_),
    .B(_0213_));
 sg13g2_nand2_1 _1813_ (.Y(_0271_),
    .A(net36),
    .B(net18));
 sg13g2_o21ai_1 _1814_ (.B1(_0271_),
    .Y(_0171_),
    .A1(net36),
    .A2(_0269_));
 sg13g2_nand2_1 _1815_ (.Y(_0272_),
    .A(net36),
    .B(_0268_));
 sg13g2_xnor2_1 _1816_ (.Y(_0172_),
    .A(_0260_),
    .B(_0272_));
 sg13g2_nand2_1 _1817_ (.Y(_0273_),
    .A(net36),
    .B(_0260_));
 sg13g2_nor3_1 _1818_ (.A(_0255_),
    .B(net18),
    .C(_0273_),
    .Y(_0274_));
 sg13g2_a21oi_1 _1819_ (.A1(_0255_),
    .A2(_0273_),
    .Y(_0275_),
    .B1(_0274_));
 sg13g2_nand2_1 _1820_ (.Y(_0276_),
    .A(_0255_),
    .B(net18));
 sg13g2_o21ai_1 _1821_ (.B1(_0276_),
    .Y(_0173_),
    .A1(_0267_),
    .A2(_0275_));
 sg13g2_nand3_1 _1822_ (.B(_0260_),
    .C(_0255_),
    .A(net36),
    .Y(_0277_));
 sg13g2_or2_1 _1823_ (.X(_0278_),
    .B(_0277_),
    .A(net18));
 sg13g2_nor2b_1 _1824_ (.A(_0267_),
    .B_N(_0277_),
    .Y(_0279_));
 sg13g2_o21ai_1 _1825_ (.B1(_0261_),
    .Y(_0280_),
    .A1(net18),
    .A2(_0279_));
 sg13g2_o21ai_1 _1826_ (.B1(_0280_),
    .Y(_0174_),
    .A1(_0261_),
    .A2(_0278_));
 sg13g2_inv_1 _1827_ (.Y(_0281_),
    .A(_0261_));
 sg13g2_nor2_1 _1828_ (.A(_0281_),
    .B(_0277_),
    .Y(_0282_));
 sg13g2_xor2_1 _1829_ (.B(_0282_),
    .A(_0006_),
    .X(_0283_));
 sg13g2_nand2_1 _1830_ (.Y(_0284_),
    .A(_0262_),
    .B(net18));
 sg13g2_o21ai_1 _1831_ (.B1(_0284_),
    .Y(_0175_),
    .A1(_0269_),
    .A2(_0283_));
 sg13g2_nand2_1 _1832_ (.Y(_0285_),
    .A(_0262_),
    .B(_0282_));
 sg13g2_xnor2_1 _1833_ (.Y(_0286_),
    .A(_0008_),
    .B(_0285_));
 sg13g2_nand2_1 _1834_ (.Y(_0287_),
    .A(_0258_),
    .B(net18));
 sg13g2_o21ai_1 _1835_ (.B1(_0287_),
    .Y(_0176_),
    .A1(_0269_),
    .A2(_0286_));
 sg13g2_nand3_1 _1836_ (.B(_0262_),
    .C(_0282_),
    .A(_0258_),
    .Y(_0288_));
 sg13g2_xnor2_1 _1837_ (.Y(_0289_),
    .A(_0007_),
    .B(_0288_));
 sg13g2_nand2_1 _1838_ (.Y(_0290_),
    .A(\top_inst.vga_inst.bg[5] ),
    .B(net18));
 sg13g2_o21ai_1 _1839_ (.B1(_0290_),
    .Y(_0177_),
    .A1(_0269_),
    .A2(_0289_));
 sg13g2_nand2_1 _1840_ (.Y(_0291_),
    .A(\top_inst.vga_inst.bg[5] ),
    .B(_0258_));
 sg13g2_nor3_2 _1841_ (.A(_0270_),
    .B(_0285_),
    .C(_0291_),
    .Y(_0292_));
 sg13g2_xor2_1 _1842_ (.B(_0292_),
    .A(_0257_),
    .X(_0178_));
 sg13g2_nand2_1 _1843_ (.Y(_0293_),
    .A(_0257_),
    .B(_0292_));
 sg13g2_xnor2_1 _1844_ (.Y(_0179_),
    .A(\top_inst.vga_inst.y[8] ),
    .B(_0293_));
 sg13g2_nand3_1 _1845_ (.B(\top_inst.vga_inst.y[8] ),
    .C(_0292_),
    .A(_0257_),
    .Y(_0294_));
 sg13g2_xor2_1 _1846_ (.B(_0294_),
    .A(_0256_),
    .X(_0295_));
 sg13g2_a21oi_1 _1847_ (.A1(_0268_),
    .A2(_0267_),
    .Y(_0180_),
    .B1(_0295_));
 sg13g2_nor4_1 _1848_ (.A(\top_inst.sys_presc[1] ),
    .B(\top_inst.sys_presc[3] ),
    .C(\top_inst.sys_presc[2] ),
    .D(\top_inst.sys_presc[4] ),
    .Y(_0296_));
 sg13g2_and2_1 _1849_ (.A(_0181_),
    .B(_0296_),
    .X(_0297_));
 sg13g2_buf_1 _1850_ (.A(_0297_),
    .X(_0298_));
 sg13g2_mux2_1 _1851_ (.A0(\top_inst.pwm_inst.cntr[0] ),
    .A1(_0018_),
    .S(_0298_),
    .X(_0023_));
 sg13g2_nand2_1 _1852_ (.Y(_0299_),
    .A(\top_inst.pwm_inst.cntr[0] ),
    .B(_0298_));
 sg13g2_xnor2_1 _1853_ (.Y(_0024_),
    .A(\top_inst.pwm_inst.cntr[1] ),
    .B(_0299_));
 sg13g2_nand3_1 _1854_ (.B(\top_inst.pwm_inst.cntr[0] ),
    .C(_0298_),
    .A(\top_inst.pwm_inst.cntr[1] ),
    .Y(_0300_));
 sg13g2_xnor2_1 _1855_ (.Y(_0025_),
    .A(\top_inst.pwm_inst.cntr[2] ),
    .B(_0300_));
 sg13g2_nand4_1 _1856_ (.B(\top_inst.pwm_inst.cntr[1] ),
    .C(\top_inst.pwm_inst.cntr[0] ),
    .A(\top_inst.pwm_inst.cntr[2] ),
    .Y(_0301_),
    .D(_0298_));
 sg13g2_xnor2_1 _1857_ (.Y(_0026_),
    .A(\top_inst.pwm_inst.cntr[3] ),
    .B(_0301_));
 sg13g2_nor3_1 _1858_ (.A(_0390_),
    .B(net38),
    .C(_0387_),
    .Y(_0302_));
 sg13g2_or3_1 _1859_ (.A(_0396_),
    .B(_0217_),
    .C(_0302_),
    .X(hsync));
 sg13g2_nand2_1 _1860_ (.Y(_0303_),
    .A(net33),
    .B(_0838_));
 sg13g2_xor2_1 _1861_ (.B(_0868_),
    .A(_0764_),
    .X(_0304_));
 sg13g2_nand3b_1 _1862_ (.B(_0840_),
    .C(_0868_),
    .Y(_0305_),
    .A_N(net33));
 sg13g2_o21ai_1 _1863_ (.B1(_0305_),
    .Y(_0306_),
    .A1(_0303_),
    .A2(_0304_));
 sg13g2_nor3_1 _1864_ (.A(net33),
    .B(_0018_),
    .C(_0868_),
    .Y(_0307_));
 sg13g2_nor3_1 _1865_ (.A(net33),
    .B(_0840_),
    .C(_0868_),
    .Y(_0308_));
 sg13g2_nor2_1 _1866_ (.A(_0467_),
    .B(_0764_),
    .Y(_0309_));
 sg13g2_nor2b_1 _1867_ (.A(_0018_),
    .B_N(_0764_),
    .Y(_0310_));
 sg13g2_nor2_1 _1868_ (.A(_0018_),
    .B(_0887_),
    .Y(_0311_));
 sg13g2_mux4_1 _1869_ (.S0(_0868_),
    .A0(_0309_),
    .A1(_0891_),
    .A2(_0310_),
    .A3(_0311_),
    .S1(_0838_),
    .X(_0312_));
 sg13g2_nor4_1 _1870_ (.A(\top_inst.pwm_inst.cntr[1] ),
    .B(_0307_),
    .C(_0308_),
    .D(_0312_),
    .Y(_0313_));
 sg13g2_a21o_1 _1871_ (.A2(_0306_),
    .A1(_0018_),
    .B1(_0313_),
    .X(_0314_));
 sg13g2_nand3_1 _1872_ (.B(_0896_),
    .C(_0314_),
    .A(_0011_),
    .Y(_0315_));
 sg13g2_nor2b_1 _1873_ (.A(\top_inst.pwm_inst.cntr[2] ),
    .B_N(_0011_),
    .Y(_0316_));
 sg13g2_nand2_1 _1874_ (.Y(_0317_),
    .A(_0314_),
    .B(_0316_));
 sg13g2_nand3b_1 _1875_ (.B(_0903_),
    .C(_0314_),
    .Y(_0318_),
    .A_N(\top_inst.pwm_inst.cntr[2] ));
 sg13g2_nand2_1 _1876_ (.Y(_0319_),
    .A(_0886_),
    .B(_0893_));
 sg13g2_nor3_1 _1877_ (.A(\top_inst.pwm_inst.cntr[2] ),
    .B(_0876_),
    .C(_0319_),
    .Y(_0320_));
 sg13g2_a221oi_1 _1878_ (.B2(_0896_),
    .C1(_0320_),
    .B1(_0316_),
    .A1(_0011_),
    .Y(_0321_),
    .A2(_0903_));
 sg13g2_nand4_1 _1879_ (.B(_0317_),
    .C(_0318_),
    .A(_0315_),
    .Y(pwm),
    .D(_0321_));
 sg13g2_nand4_1 _1880_ (.B(\top_inst.vga_inst.bg[5] ),
    .C(_0258_),
    .A(_0257_),
    .Y(_0322_),
    .D(\top_inst.vga_inst.y[8] ));
 sg13g2_nor4_1 _1881_ (.A(_0255_),
    .B(_0256_),
    .C(_0264_),
    .D(_0322_),
    .Y(_0323_));
 sg13g2_nand2_1 _1882_ (.Y(\top_inst.vga_inst.vsync ),
    .A(_0260_),
    .B(_0323_));
 sg13g2_nor4_2 _1883_ (.A(_0397_),
    .B(_0260_),
    .C(_0255_),
    .Y(_0324_),
    .D(_0261_));
 sg13g2_inv_1 _1884_ (.Y(_0325_),
    .A(_0258_));
 sg13g2_o21ai_1 _1885_ (.B1(_0325_),
    .Y(_0326_),
    .A1(_0263_),
    .A2(_0324_));
 sg13g2_nand4_1 _1886_ (.B(\top_inst.vga_inst.bg[5] ),
    .C(\top_inst.vga_inst.y[8] ),
    .A(_0257_),
    .Y(_0327_),
    .D(_0326_));
 sg13g2_nand3_1 _1887_ (.B(_0393_),
    .C(_0223_),
    .A(net28),
    .Y(_0328_));
 sg13g2_nor2b_2 _1888_ (.A(_0256_),
    .B_N(_0259_),
    .Y(_0329_));
 sg13g2_nor2_1 _1889_ (.A(net37),
    .B(_0256_),
    .Y(_0330_));
 sg13g2_o21ai_1 _1890_ (.B1(_0330_),
    .Y(_0331_),
    .A1(net28),
    .A2(_0223_));
 sg13g2_a21oi_1 _1891_ (.A1(_0263_),
    .A2(_0329_),
    .Y(_0332_),
    .B1(_0331_));
 sg13g2_nand3_1 _1892_ (.B(_0328_),
    .C(_0332_),
    .A(_0327_),
    .Y(_0333_));
 sg13g2_inv_1 _1893_ (.Y(_0334_),
    .A(_0005_));
 sg13g2_o21ai_1 _1894_ (.B1(_0394_),
    .Y(_0335_),
    .A1(net28),
    .A2(_0334_));
 sg13g2_nand2_1 _1895_ (.Y(_0336_),
    .A(_0322_),
    .B(_0335_));
 sg13g2_xnor2_1 _1896_ (.Y(_0337_),
    .A(_0905_),
    .B(_0183_));
 sg13g2_nor3_1 _1897_ (.A(net37),
    .B(_0329_),
    .C(_0337_),
    .Y(_0338_));
 sg13g2_nor3_1 _1898_ (.A(_0256_),
    .B(_0336_),
    .C(_0338_),
    .Y(_0339_));
 sg13g2_nand2_1 _1899_ (.Y(_0340_),
    .A(_0333_),
    .B(_0339_));
 sg13g2_nor2_1 _1900_ (.A(_0007_),
    .B(_0340_),
    .Y(net3));
 sg13g2_nor4_1 _1901_ (.A(net37),
    .B(net28),
    .C(_0389_),
    .D(_0182_),
    .Y(_0341_));
 sg13g2_nand2b_1 _1902_ (.Y(_0342_),
    .B(_0197_),
    .A_N(\top_inst.vga_inst.xmin[1] ));
 sg13g2_nor2b_1 _1903_ (.A(_0194_),
    .B_N(\top_inst.vga_inst.xmin[0] ),
    .Y(_0343_));
 sg13g2_nor2b_1 _1904_ (.A(_0197_),
    .B_N(\top_inst.vga_inst.xmin[1] ),
    .Y(_0344_));
 sg13g2_a221oi_1 _1905_ (.B2(_0343_),
    .C1(_0344_),
    .B1(_0342_),
    .A1(_0200_),
    .Y(_0345_),
    .A2(\top_inst.vga_inst.xmin[2] ));
 sg13g2_a21oi_1 _1906_ (.A1(\top_inst.vga_inst.x1[6] ),
    .A2(_0250_),
    .Y(_0346_),
    .B1(_0345_));
 sg13g2_nor3_1 _1907_ (.A(\top_inst.vga_inst.x1[7] ),
    .B(\top_inst.vga_inst.xmin[3] ),
    .C(_0346_),
    .Y(_0347_));
 sg13g2_nand2b_1 _1908_ (.Y(_0348_),
    .B(_0197_),
    .A_N(\top_inst.vga_inst.xmax[1] ));
 sg13g2_nor2b_1 _1909_ (.A(\top_inst.vga_inst.xmax[0] ),
    .B_N(_0194_),
    .Y(_0349_));
 sg13g2_or2_1 _1910_ (.X(_0350_),
    .B(\top_inst.vga_inst.x1[3] ),
    .A(\top_inst.vga_inst.x1[2] ));
 sg13g2_nand2b_1 _1911_ (.Y(_0351_),
    .B(\top_inst.vga_inst.xmax[0] ),
    .A_N(_0194_));
 sg13g2_o21ai_1 _1912_ (.B1(_0351_),
    .Y(_0352_),
    .A1(_0349_),
    .A2(_0350_));
 sg13g2_nor2b_1 _1913_ (.A(_0197_),
    .B_N(\top_inst.vga_inst.xmax[1] ),
    .Y(_0353_));
 sg13g2_a221oi_1 _1914_ (.B2(_0352_),
    .C1(_0353_),
    .B1(_0348_),
    .A1(_0200_),
    .Y(_0354_),
    .A2(\top_inst.vga_inst.xmax[2] ));
 sg13g2_a21oi_1 _1915_ (.A1(\top_inst.vga_inst.x1[6] ),
    .A2(_0243_),
    .Y(_0355_),
    .B1(_0354_));
 sg13g2_inv_1 _1916_ (.Y(_0356_),
    .A(\top_inst.vga_inst.x1[7] ));
 sg13g2_a21oi_1 _1917_ (.A1(\top_inst.vga_inst.xmin[3] ),
    .A2(_0346_),
    .Y(_0357_),
    .B1(_0356_));
 sg13g2_a21o_1 _1918_ (.A2(_0357_),
    .A1(_0355_),
    .B1(_0347_),
    .X(_0358_));
 sg13g2_a22oi_1 _1919_ (.Y(_0359_),
    .B1(_0358_),
    .B2(\top_inst.vga_inst.xmax[3] ),
    .A2(_0355_),
    .A1(_0347_));
 sg13g2_nor2_1 _1920_ (.A(_0389_),
    .B(_0324_),
    .Y(_0360_));
 sg13g2_nand2_1 _1921_ (.Y(_0361_),
    .A(_0359_),
    .B(_0360_));
 sg13g2_nor3_1 _1922_ (.A(\top_inst.sndgen_inst.c2[0] ),
    .B(\top_inst.sndgen_inst.c2[1] ),
    .C(\top_inst.sndgen_inst.c2[2] ),
    .Y(_0362_));
 sg13g2_or2_1 _1923_ (.X(_0363_),
    .B(_0362_),
    .A(_0831_));
 sg13g2_nor2_1 _1924_ (.A(\top_inst.sndgen_inst.c1[1] ),
    .B(\top_inst.sndgen_inst.c1[0] ),
    .Y(_0364_));
 sg13g2_or2_1 _1925_ (.X(_0365_),
    .B(_0364_),
    .A(_0834_));
 sg13g2_nor3_1 _1926_ (.A(\top_inst.sndgen_inst.c3[0] ),
    .B(\top_inst.sndgen_inst.c3[1] ),
    .C(\top_inst.sndgen_inst.c3[2] ),
    .Y(_0366_));
 sg13g2_nor2b_1 _1927_ (.A(\top_inst.sndgen_inst.c4[2] ),
    .B_N(_0366_),
    .Y(_0367_));
 sg13g2_nand2b_1 _1928_ (.Y(_0368_),
    .B(net33),
    .A_N(_0367_));
 sg13g2_nand2b_1 _1929_ (.Y(_0369_),
    .B(_0463_),
    .A_N(_0366_));
 sg13g2_mux4_1 _1930_ (.S0(_0444_),
    .A0(_0363_),
    .A1(_0365_),
    .A2(_0368_),
    .A3(_0369_),
    .S1(net38),
    .X(_0370_));
 sg13g2_nand4_1 _1931_ (.B(_0329_),
    .C(_0341_),
    .A(_0262_),
    .Y(_0371_),
    .D(_0370_));
 sg13g2_o21ai_1 _1932_ (.B1(_0371_),
    .Y(_0372_),
    .A1(_0341_),
    .A2(_0361_));
 sg13g2_nor2b_1 _1933_ (.A(_0324_),
    .B_N(_0372_),
    .Y(_0373_));
 sg13g2_a21oi_1 _1934_ (.A1(_0262_),
    .A2(_0329_),
    .Y(_0374_),
    .B1(_0361_));
 sg13g2_nor3_1 _1935_ (.A(_0333_),
    .B(_0373_),
    .C(_0374_),
    .Y(net4));
 sg13g2_nor2_1 _1936_ (.A(_0006_),
    .B(_0340_),
    .Y(net5));
 sg13g2_inv_1 _1937_ (.Y(_0375_),
    .A(_0333_));
 sg13g2_inv_1 _1938_ (.Y(_0376_),
    .A(_0007_));
 sg13g2_a21oi_1 _1939_ (.A1(net37),
    .A2(_0389_),
    .Y(_0377_),
    .B1(_0444_));
 sg13g2_o21ai_1 _1940_ (.B1(_0223_),
    .Y(_0378_),
    .A1(net38),
    .A2(_0377_));
 sg13g2_nor3_1 _1941_ (.A(\top_inst.vga_inst.x[8] ),
    .B(_0392_),
    .C(_0182_),
    .Y(_0379_));
 sg13g2_a21oi_1 _1942_ (.A1(_0905_),
    .A2(_0378_),
    .Y(_0380_),
    .B1(_0379_));
 sg13g2_nand2_1 _1943_ (.Y(_0381_),
    .A(_0322_),
    .B(_0330_));
 sg13g2_nor3_1 _1944_ (.A(_0329_),
    .B(_0380_),
    .C(_0381_),
    .Y(_0382_));
 sg13g2_nor4_1 _1945_ (.A(_0256_),
    .B(_0008_),
    .C(_0336_),
    .D(_0382_),
    .Y(_0383_));
 sg13g2_a21oi_1 _1946_ (.A1(_0376_),
    .A2(_0382_),
    .Y(_0384_),
    .B1(_0383_));
 sg13g2_nor2_1 _1947_ (.A(_0375_),
    .B(_0384_),
    .Y(net7));
 sg13g2_inv_1 _1948_ (.Y(_0385_),
    .A(_0360_));
 sg13g2_a21oi_1 _1949_ (.A1(_0359_),
    .A2(_0385_),
    .Y(net8),
    .B1(_0333_));
 sg13g2_a22oi_1 _1950_ (.Y(_0386_),
    .B1(_0382_),
    .B2(_0262_),
    .A2(_0339_),
    .A1(_0261_));
 sg13g2_nor2_1 _1951_ (.A(_0375_),
    .B(_0386_),
    .Y(net9));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _1961__83 (.L_HI(net83));
 sg13g2_buf_1 _1954_ (.A(net69),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1955_ (.A(net70),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1956_ (.A(net71),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1957_ (.A(net72),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1958_ (.A(net73),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1959_ (.A(net74),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1960_ (.A(net75),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1961_ (.A(net83),
    .X(uio_oe[7]));
 sg13g2_buf_1 _1962_ (.A(net76),
    .X(uio_out[0]));
 sg13g2_buf_1 _1963_ (.A(net77),
    .X(uio_out[1]));
 sg13g2_buf_1 _1964_ (.A(net78),
    .X(uio_out[2]));
 sg13g2_buf_1 _1965_ (.A(net79),
    .X(uio_out[3]));
 sg13g2_buf_1 _1966_ (.A(net80),
    .X(uio_out[4]));
 sg13g2_buf_1 _1967_ (.A(net81),
    .X(uio_out[5]));
 sg13g2_buf_1 _1968_ (.A(net82),
    .X(uio_out[6]));
 sg13g2_buf_1 _1969_ (.A(pwm),
    .X(net2));
 sg13g2_buf_1 _1970_ (.A(\top_inst.vga_inst.vsync ),
    .X(net6));
 sg13g2_buf_1 _1971_ (.A(hsync),
    .X(net10));
 sg13g2_dfrbp_1 \top_inst.pwm_inst.cntr[0]$_DFFE_PN0N_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net46),
    .D(_0023_),
    .Q_N(_0018_),
    .Q(\top_inst.pwm_inst.cntr[0] ));
 sg13g2_dfrbp_1 \top_inst.pwm_inst.cntr[1]$_DFFE_PN0N_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net46),
    .D(_0024_),
    .Q_N(_1046_),
    .Q(\top_inst.pwm_inst.cntr[1] ));
 sg13g2_dfrbp_1 \top_inst.pwm_inst.cntr[2]$_DFFE_PN0N_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net46),
    .D(_0025_),
    .Q_N(_1045_),
    .Q(\top_inst.pwm_inst.cntr[2] ));
 sg13g2_dfrbp_1 \top_inst.pwm_inst.cntr[3]$_DFFE_PN0N_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net46),
    .D(_0026_),
    .Q_N(_0011_),
    .Q(\top_inst.pwm_inst.cntr[3] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.c1[0]$_DFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net40),
    .D(_0027_),
    .Q_N(_1044_),
    .Q(\top_inst.sndgen_inst.c1[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.c1[1]$_DFFE_PN1P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net40),
    .D(_0028_),
    .Q_N(\top_inst.sndgen_inst.c1[1] ),
    .Q(_0020_));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.c2[0]$_DFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net43),
    .D(_0029_),
    .Q_N(_1043_),
    .Q(\top_inst.sndgen_inst.c2[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.c2[1]$_DFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net43),
    .D(_0030_),
    .Q_N(_1042_),
    .Q(\top_inst.sndgen_inst.c2[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.c2[2]$_DFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net43),
    .D(_0031_),
    .Q_N(_1041_),
    .Q(\top_inst.sndgen_inst.c2[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.c3[0]$_DFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net43),
    .D(_0032_),
    .Q_N(_1040_),
    .Q(\top_inst.sndgen_inst.c3[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.c3[1]$_DFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net43),
    .D(_0033_),
    .Q_N(_1039_),
    .Q(\top_inst.sndgen_inst.c3[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.c4[2]$_DFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net43),
    .D(_0034_),
    .Q_N(_1038_),
    .Q(\top_inst.sndgen_inst.c4[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.c4[3]$_DFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net43),
    .D(_0035_),
    .Q_N(_1037_),
    .Q(\top_inst.sndgen_inst.c3[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.lfsr[0]$_DFFE_PN1P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net49),
    .D(_0036_),
    .Q_N(\top_inst.sndgen_inst.lfsr[0] ),
    .Q(_0021_));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.lfsr[1]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net49),
    .D(_0037_),
    .Q_N(_1036_),
    .Q(\top_inst.sndgen_inst.lfsr[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.lfsr[2]$_DFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net49),
    .D(_0038_),
    .Q_N(_1035_),
    .Q(\top_inst.sndgen_inst.lfsr[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.lfsr[3]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net49),
    .D(_0039_),
    .Q_N(_1034_),
    .Q(\top_inst.sndgen_inst.lfsr[3] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.lfsr[4]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net50),
    .D(_0040_),
    .Q_N(_1033_),
    .Q(\top_inst.sndgen_inst.lfsr[4] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.lfsr[5]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net50),
    .D(_0041_),
    .Q_N(_1032_),
    .Q(\top_inst.sndgen_inst.lfsr[5] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.lfsr[6]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net50),
    .D(_0042_),
    .Q_N(_1031_),
    .Q(\top_inst.sndgen_inst.lfsr[6] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.lfsr[7]$_DFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net49),
    .D(_0043_),
    .Q_N(_0009_),
    .Q(\top_inst.sndgen_inst.lfsr[7] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.mask_1[0]$_DFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net49),
    .D(_0044_),
    .Q_N(_1030_),
    .Q(\top_inst.sndgen_inst.mask_1[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.mask_1[1]$_DFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net49),
    .D(_0045_),
    .Q_N(_0012_),
    .Q(\top_inst.sndgen_inst.mask_1[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.mask_1[2]$_DFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net48),
    .D(_0046_),
    .Q_N(_1029_),
    .Q(\top_inst.sndgen_inst.mask_1[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.mask_1[3]$_DFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net48),
    .D(_0047_),
    .Q_N(_1028_),
    .Q(\top_inst.sndgen_inst.mask_1[3] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.mask_2$_DFFE_PN1P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net49),
    .D(_0048_),
    .Q_N(\top_inst.sndgen_inst.mask_2 ),
    .Q(_0022_));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c2[0]$_DFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net53),
    .D(_0049_),
    .Q_N(_1027_),
    .Q(\top_inst.sndgen_inst.p_c2[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c2[12]$_DFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net42),
    .D(_0050_),
    .Q_N(_1026_),
    .Q(\top_inst.sndgen_inst.p_c2[10] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c2[1]$_DFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net53),
    .D(_0051_),
    .Q_N(_1025_),
    .Q(\top_inst.sndgen_inst.p_c2[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c2[2]$_DFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net53),
    .D(_0052_),
    .Q_N(_1024_),
    .Q(\top_inst.sndgen_inst.p_c2[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c2[3]$_DFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net53),
    .D(_0053_),
    .Q_N(_1023_),
    .Q(\top_inst.sndgen_inst.p_c2[3] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c2[4]$_DFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net42),
    .D(_0054_),
    .Q_N(_1022_),
    .Q(\top_inst.sndgen_inst.p_c2[4] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c2[5]$_DFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net42),
    .D(_0055_),
    .Q_N(_1021_),
    .Q(\top_inst.sndgen_inst.p_c2[5] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c2[6]$_DFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net42),
    .D(_0056_),
    .Q_N(_1020_),
    .Q(\top_inst.sndgen_inst.p_c2[6] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c2[7]$_DFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net44),
    .D(_0057_),
    .Q_N(_1019_),
    .Q(\top_inst.sndgen_inst.p_c2[7] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c3[0]$_DFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net53),
    .D(_0058_),
    .Q_N(_1018_),
    .Q(\top_inst.sndgen_inst.p_c3[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c3[12]$_DFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net55),
    .D(_0059_),
    .Q_N(_1017_),
    .Q(\top_inst.sndgen_inst.p_c3[10] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c3[1]$_DFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net53),
    .D(_0060_),
    .Q_N(_1016_),
    .Q(\top_inst.sndgen_inst.p_c3[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c3[2]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net58),
    .D(_0061_),
    .Q_N(_1015_),
    .Q(\top_inst.sndgen_inst.p_c3[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c3[3]$_DFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net56),
    .D(_0062_),
    .Q_N(_1014_),
    .Q(\top_inst.sndgen_inst.p_c3[3] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c3[4]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net60),
    .D(_0063_),
    .Q_N(_1013_),
    .Q(\top_inst.sndgen_inst.p_c3[4] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c3[5]$_DFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net54),
    .D(_0064_),
    .Q_N(_1012_),
    .Q(\top_inst.sndgen_inst.p_c3[5] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c3[6]$_DFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net54),
    .D(_0065_),
    .Q_N(_1011_),
    .Q(\top_inst.sndgen_inst.p_c3[6] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c3[7]$_DFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net56),
    .D(_0066_),
    .Q_N(_1010_),
    .Q(\top_inst.sndgen_inst.p_c3[7] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c4[0]$_DFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net60),
    .D(_0067_),
    .Q_N(_1009_),
    .Q(\top_inst.sndgen_inst.p_c4[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c4[12]$_DFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net55),
    .D(_0068_),
    .Q_N(_1008_),
    .Q(\top_inst.sndgen_inst.p_c4[10] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c4[1]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net60),
    .D(_0069_),
    .Q_N(_1007_),
    .Q(\top_inst.sndgen_inst.p_c4[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c4[2]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net58),
    .D(_0070_),
    .Q_N(_1006_),
    .Q(\top_inst.sndgen_inst.p_c4[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c4[3]$_DFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net58),
    .D(_0071_),
    .Q_N(_1005_),
    .Q(\top_inst.sndgen_inst.p_c4[3] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c4[4]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net58),
    .D(_0072_),
    .Q_N(_1004_),
    .Q(\top_inst.sndgen_inst.p_c4[4] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c4[5]$_DFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net58),
    .D(_0073_),
    .Q_N(_1003_),
    .Q(\top_inst.sndgen_inst.p_c4[5] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c4[6]$_DFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net58),
    .D(_0074_),
    .Q_N(_1002_),
    .Q(\top_inst.sndgen_inst.p_c4[6] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.p_c4[7]$_DFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net58),
    .D(_0075_),
    .Q_N(_1001_),
    .Q(\top_inst.sndgen_inst.p_c4[7] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[0]$_DFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net53),
    .D(_0076_),
    .Q_N(_1000_),
    .Q(\top_inst.sndgen_inst.phacc2[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[10]$_DFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net42),
    .D(_0077_),
    .Q_N(_0999_),
    .Q(\top_inst.sndgen_inst.phacc2[10] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[11]$_DFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net41),
    .D(_0078_),
    .Q_N(_0998_),
    .Q(\top_inst.sndgen_inst.phacc2[11] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[12]$_DFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net41),
    .D(_0079_),
    .Q_N(_0997_),
    .Q(\top_inst.sndgen_inst.phacc2[12] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[13]$_DFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net48),
    .D(_0080_),
    .Q_N(_0996_),
    .Q(\top_inst.sndgen_inst.phacc2[13] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[1]$_DFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net53),
    .D(_0081_),
    .Q_N(_0995_),
    .Q(\top_inst.sndgen_inst.phacc2[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[2]$_DFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net54),
    .D(_0082_),
    .Q_N(_0994_),
    .Q(\top_inst.sndgen_inst.phacc2[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[3]$_DFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net54),
    .D(_0083_),
    .Q_N(_0993_),
    .Q(\top_inst.sndgen_inst.phacc2[3] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[4]$_DFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net44),
    .D(_0084_),
    .Q_N(_0992_),
    .Q(\top_inst.sndgen_inst.phacc2[4] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[5]$_DFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net42),
    .D(_0085_),
    .Q_N(_0991_),
    .Q(\top_inst.sndgen_inst.phacc2[5] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[6]$_DFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net42),
    .D(_0086_),
    .Q_N(_0990_),
    .Q(\top_inst.sndgen_inst.phacc2[6] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[7]$_DFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net41),
    .D(_0087_),
    .Q_N(_0989_),
    .Q(\top_inst.sndgen_inst.phacc2[7] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[8]$_DFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net41),
    .D(_0088_),
    .Q_N(_0001_),
    .Q(\top_inst.sndgen_inst.phacc2[8] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc2[9]$_DFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net42),
    .D(_0089_),
    .Q_N(_0988_),
    .Q(\top_inst.sndgen_inst.phacc2[9] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[0]$_DFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net55),
    .D(_0090_),
    .Q_N(_0987_),
    .Q(\top_inst.sndgen_inst.phacc3[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[10]$_DFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net63),
    .D(_0091_),
    .Q_N(_0986_),
    .Q(\top_inst.sndgen_inst.phacc3[10] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[11]$_DFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net61),
    .D(_0092_),
    .Q_N(_0985_),
    .Q(\top_inst.sndgen_inst.phacc3[11] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[12]$_DFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net63),
    .D(_0093_),
    .Q_N(_0984_),
    .Q(\top_inst.sndgen_inst.phacc3[12] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[13]$_DFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net48),
    .D(_0094_),
    .Q_N(_0983_),
    .Q(\top_inst.sndgen_inst.phacc3[13] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[1]$_DFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net55),
    .D(_0095_),
    .Q_N(_0982_),
    .Q(\top_inst.sndgen_inst.phacc3[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[2]$_DFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net56),
    .D(_0096_),
    .Q_N(_0981_),
    .Q(\top_inst.sndgen_inst.phacc3[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[3]$_DFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net58),
    .D(_0097_),
    .Q_N(_0980_),
    .Q(\top_inst.sndgen_inst.phacc3[3] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[4]$_DFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net60),
    .D(_0098_),
    .Q_N(_0979_),
    .Q(\top_inst.sndgen_inst.phacc3[4] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[5]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net60),
    .D(_0099_),
    .Q_N(_0978_),
    .Q(\top_inst.sndgen_inst.phacc3[5] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[6]$_DFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net54),
    .D(_0100_),
    .Q_N(_0977_),
    .Q(\top_inst.sndgen_inst.phacc3[6] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[7]$_DFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net63),
    .D(_0101_),
    .Q_N(_0976_),
    .Q(\top_inst.sndgen_inst.phacc3[7] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[8]$_DFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net56),
    .D(_0102_),
    .Q_N(_0013_),
    .Q(\top_inst.sndgen_inst.phacc3[8] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc3[9]$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net61),
    .D(_0103_),
    .Q_N(_0975_),
    .Q(\top_inst.sndgen_inst.phacc3[9] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[0]$_DFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net60),
    .D(_0104_),
    .Q_N(_0974_),
    .Q(\top_inst.sndgen_inst.phacc4[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[10]$_DFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net61),
    .D(_0105_),
    .Q_N(_0973_),
    .Q(\top_inst.sndgen_inst.phacc4[10] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[11]$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net61),
    .D(_0106_),
    .Q_N(_0972_),
    .Q(\top_inst.sndgen_inst.phacc4[11] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[12]$_DFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net61),
    .D(_0107_),
    .Q_N(_0971_),
    .Q(\top_inst.sndgen_inst.phacc4[12] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[13]$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net61),
    .D(_0108_),
    .Q_N(_0970_),
    .Q(\top_inst.sndgen_inst.phacc4[13] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[1]$_DFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net60),
    .D(_0109_),
    .Q_N(_0969_),
    .Q(\top_inst.sndgen_inst.phacc4[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[2]$_DFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net59),
    .D(_0110_),
    .Q_N(_0968_),
    .Q(\top_inst.sndgen_inst.phacc4[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[3]$_DFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net59),
    .D(_0111_),
    .Q_N(_0967_),
    .Q(\top_inst.sndgen_inst.phacc4[3] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[4]$_DFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net59),
    .D(_0112_),
    .Q_N(_0966_),
    .Q(\top_inst.sndgen_inst.phacc4[4] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[5]$_DFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net59),
    .D(_0113_),
    .Q_N(_0965_),
    .Q(\top_inst.sndgen_inst.phacc4[5] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[6]$_DFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net63),
    .D(_0114_),
    .Q_N(_0964_),
    .Q(\top_inst.sndgen_inst.phacc4[6] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[7]$_DFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net63),
    .D(_0115_),
    .Q_N(_0963_),
    .Q(\top_inst.sndgen_inst.phacc4[7] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[8]$_DFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net63),
    .D(_0116_),
    .Q_N(_0000_),
    .Q(\top_inst.sndgen_inst.phacc4[8] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.phacc4[9]$_DFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net55),
    .D(_0117_),
    .Q_N(_0962_),
    .Q(\top_inst.sndgen_inst.phacc4[9] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.rom_addr[0]$_DFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net44),
    .D(_0118_),
    .Q_N(_0961_),
    .Q(\top_inst.sndgen_inst.rom_addr[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.rom_addr[1]$_DFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net44),
    .D(_0119_),
    .Q_N(_0960_),
    .Q(\top_inst.sndgen_inst.rom_addr[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.rom_addr[2]$_DFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net44),
    .D(_0120_),
    .Q_N(_0004_),
    .Q(\top_inst.sndgen_inst.rom_addr[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.rom_addr[3]$_DFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net55),
    .D(_0121_),
    .Q_N(_0003_),
    .Q(\top_inst.sndgen_inst.rom_addr[3] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.sample_ena_delay[0]$_DFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net55),
    .D(net22),
    .Q_N(_1047_),
    .Q(\top_inst.sndgen_inst.sample_ena_delay[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.sample_ena_delay[1]$_DFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net55),
    .D(\top_inst.sndgen_inst.sample_ena_delay[0] ),
    .Q_N(_1048_),
    .Q(\top_inst.sndgen_inst.sample_ena_delay[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.sample_ena_delay[2]$_DFF_PN0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net59),
    .D(\top_inst.sndgen_inst.sample_ena_delay[1] ),
    .Q_N(_0959_),
    .Q(\top_inst.sndgen_inst.sample_ena_delay[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[0]$_DFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net40),
    .D(_0122_),
    .Q_N(_0019_),
    .Q(\top_inst.sndgen_inst.slot_counter[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[10]$_DFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net39),
    .D(_0123_),
    .Q_N(_0002_),
    .Q(\top_inst.sndgen_inst.slot_counter[10] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[11]$_DFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net39),
    .D(_0124_),
    .Q_N(_0958_),
    .Q(\top_inst.sndgen_inst.bar_counter[0] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[12]$_DFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net39),
    .D(_0125_),
    .Q_N(_0957_),
    .Q(\top_inst.sndgen_inst.bar_counter[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[13]$_DFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net39),
    .D(_0126_),
    .Q_N(_0010_),
    .Q(\top_inst.sndgen_inst.bar_counter[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[14]$_DFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net39),
    .D(_0127_),
    .Q_N(_0956_),
    .Q(\top_inst.sndgen_inst.bar_counter[3] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[1]$_DFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net43),
    .D(_0128_),
    .Q_N(_0955_),
    .Q(\top_inst.sndgen_inst.slot_counter[1] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[2]$_DFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net40),
    .D(_0129_),
    .Q_N(_0954_),
    .Q(\top_inst.sndgen_inst.slot_counter[2] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[3]$_DFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net41),
    .D(_0130_),
    .Q_N(_0953_),
    .Q(\top_inst.sndgen_inst.slot_counter[3] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[4]$_DFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net39),
    .D(_0131_),
    .Q_N(_0952_),
    .Q(\top_inst.sndgen_inst.slot_counter[4] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[5]$_DFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net41),
    .D(_0132_),
    .Q_N(_0951_),
    .Q(\top_inst.sndgen_inst.slot_counter[5] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[6]$_DFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net39),
    .D(_0133_),
    .Q_N(_0950_),
    .Q(\top_inst.sndgen_inst.slot_counter[6] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[7]$_DFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net41),
    .D(_0134_),
    .Q_N(_0949_),
    .Q(\top_inst.sndgen_inst.slot_counter[7] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[8]$_DFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net41),
    .D(_0135_),
    .Q_N(_0948_),
    .Q(\top_inst.sndgen_inst.slot_counter[8] ));
 sg13g2_dfrbp_1 \top_inst.sndgen_inst.slot_counter[9]$_DFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net39),
    .D(_0136_),
    .Q_N(_1049_),
    .Q(\top_inst.sndgen_inst.slot_counter[9] ));
 sg13g2_dfrbp_1 \top_inst.sys_presc[0]$_DFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net50),
    .D(_0906_),
    .Q_N(_0906_),
    .Q(\top_inst.sys_presc[0] ));
 sg13g2_dfrbp_1 \top_inst.sys_presc[1]$_DFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net46),
    .D(_0014_),
    .Q_N(_1050_),
    .Q(\top_inst.sys_presc[1] ));
 sg13g2_dfrbp_1 \top_inst.sys_presc[2]$_DFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net46),
    .D(_0015_),
    .Q_N(_1051_),
    .Q(\top_inst.sys_presc[2] ));
 sg13g2_dfrbp_1 \top_inst.sys_presc[3]$_DFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net46),
    .D(_0016_),
    .Q_N(_1052_),
    .Q(\top_inst.sys_presc[3] ));
 sg13g2_dfrbp_1 \top_inst.sys_presc[4]$_DFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net46),
    .D(_0017_),
    .Q_N(_0947_),
    .Q(\top_inst.sys_presc[4] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.sr1[0]$_DFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net63),
    .D(_0137_),
    .Q_N(_0946_),
    .Q(\top_inst.vga_inst.sr1[0] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.sr1[1]$_DFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net66),
    .D(_0138_),
    .Q_N(_0945_),
    .Q(\top_inst.vga_inst.sr1[1] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.sr1[2]$_DFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net63),
    .D(_0139_),
    .Q_N(_0944_),
    .Q(\top_inst.vga_inst.sr1[2] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.sr1[3]$_DFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net61),
    .D(_0140_),
    .Q_N(_0943_),
    .Q(\top_inst.vga_inst.sr1[3] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.sx1[0]$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net61),
    .D(_0141_),
    .Q_N(_0942_),
    .Q(\top_inst.vga_inst.sx1[0] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.sx1[1]$_DFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net66),
    .D(_0142_),
    .Q_N(_0941_),
    .Q(\top_inst.vga_inst.sx1[1] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.sx1[2]$_DFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net47),
    .D(_0143_),
    .Q_N(_0940_),
    .Q(\top_inst.vga_inst.sx1[2] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.sx1[3]$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net62),
    .D(_0144_),
    .Q_N(_0939_),
    .Q(\top_inst.vga_inst.sx1[3] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x1[0]$_DFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net62),
    .D(_0145_),
    .Q_N(_0938_),
    .Q(\top_inst.vga_inst.x1[0] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x1[1]$_DFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net64),
    .D(_0146_),
    .Q_N(_0937_),
    .Q(\top_inst.vga_inst.x1[1] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x1[2]$_DFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net64),
    .D(_0147_),
    .Q_N(_0936_),
    .Q(\top_inst.vga_inst.x1[2] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x1[3]$_DFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net65),
    .D(_0148_),
    .Q_N(_0935_),
    .Q(\top_inst.vga_inst.x1[3] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x1[4]$_DFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net65),
    .D(_0149_),
    .Q_N(_0934_),
    .Q(\top_inst.vga_inst.x1[4] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x1[5]$_DFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net65),
    .D(_0150_),
    .Q_N(_0933_),
    .Q(\top_inst.vga_inst.x1[5] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x1[6]$_DFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net64),
    .D(_0151_),
    .Q_N(_0932_),
    .Q(\top_inst.vga_inst.x1[6] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x1[7]$_DFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net64),
    .D(_0152_),
    .Q_N(_0931_),
    .Q(\top_inst.vga_inst.x1[7] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x[0]$_DFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net47),
    .D(_0153_),
    .Q_N(_0930_),
    .Q(\top_inst.vga_inst.x[0] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x[1]$_DFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net47),
    .D(_0154_),
    .Q_N(_0929_),
    .Q(\top_inst.vga_inst.x[1] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x[2]$_DFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net47),
    .D(_0155_),
    .Q_N(_0928_),
    .Q(\top_inst.vga_inst.x[2] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x[3]$_DFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net47),
    .D(_0156_),
    .Q_N(_0927_),
    .Q(\top_inst.vga_inst.x[3] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x[4]$_DFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net50),
    .D(_0157_),
    .Q_N(_0926_),
    .Q(\top_inst.vga_inst.x[4] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x[5]$_DFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net47),
    .D(_0158_),
    .Q_N(_0925_),
    .Q(\top_inst.vga_inst.x[5] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x[6]$_DFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net50),
    .D(_0159_),
    .Q_N(_0924_),
    .Q(\top_inst.vga_inst.x[6] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x[7]$_DFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net50),
    .D(_0160_),
    .Q_N(_0005_),
    .Q(\top_inst.vga_inst.x[7] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x[8]$_DFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net47),
    .D(_0161_),
    .Q_N(_0923_),
    .Q(\top_inst.vga_inst.x[8] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.x[9]$_DFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net51),
    .D(_0162_),
    .Q_N(_0922_),
    .Q(\top_inst.vga_inst.x[9] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.xmax[0]$_DFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net65),
    .D(_0163_),
    .Q_N(_0921_),
    .Q(\top_inst.vga_inst.xmax[0] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.xmax[1]$_DFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net65),
    .D(_0164_),
    .Q_N(_0920_),
    .Q(\top_inst.vga_inst.xmax[1] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.xmax[2]$_DFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net64),
    .D(_0165_),
    .Q_N(_0919_),
    .Q(\top_inst.vga_inst.xmax[2] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.xmax[3]$_DFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net64),
    .D(_0166_),
    .Q_N(_0918_),
    .Q(\top_inst.vga_inst.xmax[3] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.xmin[0]$_DFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net65),
    .D(_0167_),
    .Q_N(_0917_),
    .Q(\top_inst.vga_inst.xmin[0] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.xmin[1]$_DFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net66),
    .D(_0168_),
    .Q_N(_0916_),
    .Q(\top_inst.vga_inst.xmin[1] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.xmin[2]$_DFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net64),
    .D(_0169_),
    .Q_N(_0915_),
    .Q(\top_inst.vga_inst.xmin[2] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.xmin[3]$_DFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net64),
    .D(_0170_),
    .Q_N(_0914_),
    .Q(\top_inst.vga_inst.xmin[3] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.y[0]$_DFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net51),
    .D(_0171_),
    .Q_N(_0913_),
    .Q(\top_inst.vga_inst.y[0] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.y[1]$_DFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net51),
    .D(_0172_),
    .Q_N(_0912_),
    .Q(\top_inst.vga_inst.y[1] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.y[2]$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net62),
    .D(_0173_),
    .Q_N(_0911_),
    .Q(\top_inst.vga_inst.y[2] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.y[3]$_DFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net62),
    .D(_0174_),
    .Q_N(_0910_),
    .Q(\top_inst.vga_inst.bg[0] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.y[4]$_DFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net51),
    .D(_0175_),
    .Q_N(_0006_),
    .Q(\top_inst.vga_inst.bg[1] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.y[5]$_DFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net62),
    .D(_0176_),
    .Q_N(_0008_),
    .Q(\top_inst.vga_inst.bg[4] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.y[6]$_DFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net62),
    .D(_0177_),
    .Q_N(_0007_),
    .Q(\top_inst.vga_inst.bg[5] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.y[7]$_DFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net62),
    .D(_0178_),
    .Q_N(_0909_),
    .Q(\top_inst.vga_inst.y[7] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.y[8]$_DFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net67),
    .D(_0179_),
    .Q_N(_0908_),
    .Q(\top_inst.vga_inst.y[8] ));
 sg13g2_dfrbp_1 \top_inst.vga_inst.y[9]$_DFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net67),
    .D(_0180_),
    .Q_N(_0907_),
    .Q(\top_inst.vga_inst.y[9] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uio_out[7]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout11 (.A(_0575_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_0415_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0695_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_0622_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_0453_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0452_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0449_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0270_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0241_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0185_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0448_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(\top_inst.sample_ena ),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0851_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0525_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0514_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0478_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0401_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0905_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0734_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0513_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0477_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0472_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0466_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0434_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0409_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0397_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0394_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0391_),
    .X(net38));
 sg13g2_buf_4 fanout39 (.X(net39),
    .A(net45));
 sg13g2_buf_2 fanout40 (.A(net45),
    .X(net40));
 sg13g2_buf_4 fanout41 (.X(net41),
    .A(net45));
 sg13g2_buf_4 fanout42 (.X(net42),
    .A(net44));
 sg13g2_buf_4 fanout43 (.X(net43),
    .A(net44));
 sg13g2_buf_4 fanout44 (.X(net44),
    .A(net45));
 sg13g2_buf_1 fanout45 (.A(net52),
    .X(net45));
 sg13g2_buf_4 fanout46 (.X(net46),
    .A(net47));
 sg13g2_buf_4 fanout47 (.X(net47),
    .A(net48));
 sg13g2_buf_2 fanout48 (.A(net52),
    .X(net48));
 sg13g2_buf_4 fanout49 (.X(net49),
    .A(net50));
 sg13g2_buf_4 fanout50 (.X(net50),
    .A(net52));
 sg13g2_buf_2 fanout51 (.A(net52),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(net68),
    .X(net52));
 sg13g2_buf_4 fanout53 (.X(net53),
    .A(net57));
 sg13g2_buf_2 fanout54 (.A(net57),
    .X(net54));
 sg13g2_buf_4 fanout55 (.X(net55),
    .A(net57));
 sg13g2_buf_2 fanout56 (.A(net57),
    .X(net56));
 sg13g2_buf_1 fanout57 (.A(net68),
    .X(net57));
 sg13g2_buf_4 fanout58 (.X(net58),
    .A(net59));
 sg13g2_buf_2 fanout59 (.A(net60),
    .X(net59));
 sg13g2_buf_4 fanout60 (.X(net60),
    .A(net68));
 sg13g2_buf_4 fanout61 (.X(net61),
    .A(net62));
 sg13g2_buf_4 fanout62 (.X(net62),
    .A(net67));
 sg13g2_buf_4 fanout63 (.X(net63),
    .A(net66));
 sg13g2_buf_4 fanout64 (.X(net64),
    .A(net66));
 sg13g2_buf_2 fanout65 (.A(net66),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(net67),
    .X(net66));
 sg13g2_buf_1 fanout67 (.A(net68),
    .X(net67));
 sg13g2_buf_1 fanout68 (.A(net1),
    .X(net68));
 sg13g2_tielo _1954__69 (.L_LO(net69));
 sg13g2_tielo _1955__70 (.L_LO(net70));
 sg13g2_tielo _1956__71 (.L_LO(net71));
 sg13g2_tielo _1957__72 (.L_LO(net72));
 sg13g2_tielo _1958__73 (.L_LO(net73));
 sg13g2_tielo _1959__74 (.L_LO(net74));
 sg13g2_tielo _1960__75 (.L_LO(net75));
 sg13g2_tielo _1962__76 (.L_LO(net76));
 sg13g2_tielo _1963__77 (.L_LO(net77));
 sg13g2_tielo _1964__78 (.L_LO(net78));
 sg13g2_tielo _1965__79 (.L_LO(net79));
 sg13g2_tielo _1966__80 (.L_LO(net80));
 sg13g2_tielo _1967__81 (.L_LO(net81));
 sg13g2_tielo _1968__82 (.L_LO(net82));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_25__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_fill_2 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_215 ();
 sg13g2_decap_8 FILLER_0_222 ();
 sg13g2_decap_8 FILLER_0_229 ();
 sg13g2_decap_8 FILLER_0_236 ();
 sg13g2_decap_8 FILLER_0_243 ();
 sg13g2_decap_8 FILLER_0_250 ();
 sg13g2_decap_8 FILLER_0_257 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_313 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_decap_8 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_0_334 ();
 sg13g2_decap_8 FILLER_0_341 ();
 sg13g2_decap_8 FILLER_0_348 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_8 FILLER_0_404 ();
 sg13g2_decap_8 FILLER_0_411 ();
 sg13g2_decap_8 FILLER_0_418 ();
 sg13g2_decap_4 FILLER_0_425 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_fill_2 FILLER_1_125 ();
 sg13g2_decap_8 FILLER_1_131 ();
 sg13g2_decap_4 FILLER_1_138 ();
 sg13g2_decap_8 FILLER_1_159 ();
 sg13g2_decap_4 FILLER_1_166 ();
 sg13g2_fill_2 FILLER_1_170 ();
 sg13g2_fill_1 FILLER_1_180 ();
 sg13g2_decap_4 FILLER_1_193 ();
 sg13g2_fill_2 FILLER_1_205 ();
 sg13g2_decap_8 FILLER_1_212 ();
 sg13g2_decap_4 FILLER_1_219 ();
 sg13g2_fill_2 FILLER_1_223 ();
 sg13g2_fill_2 FILLER_1_237 ();
 sg13g2_fill_1 FILLER_1_239 ();
 sg13g2_fill_1 FILLER_1_282 ();
 sg13g2_decap_8 FILLER_1_309 ();
 sg13g2_decap_8 FILLER_1_316 ();
 sg13g2_decap_8 FILLER_1_323 ();
 sg13g2_decap_8 FILLER_1_330 ();
 sg13g2_decap_8 FILLER_1_337 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_decap_8 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_4 FILLER_2_91 ();
 sg13g2_fill_1 FILLER_2_95 ();
 sg13g2_fill_2 FILLER_2_104 ();
 sg13g2_decap_8 FILLER_2_110 ();
 sg13g2_fill_2 FILLER_2_117 ();
 sg13g2_fill_1 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_132 ();
 sg13g2_decap_4 FILLER_2_139 ();
 sg13g2_fill_1 FILLER_2_161 ();
 sg13g2_decap_4 FILLER_2_183 ();
 sg13g2_fill_1 FILLER_2_187 ();
 sg13g2_decap_8 FILLER_2_191 ();
 sg13g2_decap_8 FILLER_2_198 ();
 sg13g2_decap_4 FILLER_2_214 ();
 sg13g2_fill_1 FILLER_2_218 ();
 sg13g2_fill_1 FILLER_2_231 ();
 sg13g2_fill_2 FILLER_2_242 ();
 sg13g2_decap_4 FILLER_2_249 ();
 sg13g2_fill_1 FILLER_2_253 ();
 sg13g2_fill_1 FILLER_2_268 ();
 sg13g2_decap_8 FILLER_2_324 ();
 sg13g2_decap_8 FILLER_2_331 ();
 sg13g2_decap_4 FILLER_2_338 ();
 sg13g2_fill_1 FILLER_2_342 ();
 sg13g2_decap_8 FILLER_2_351 ();
 sg13g2_decap_8 FILLER_2_358 ();
 sg13g2_decap_8 FILLER_2_365 ();
 sg13g2_decap_8 FILLER_2_372 ();
 sg13g2_decap_8 FILLER_2_379 ();
 sg13g2_decap_8 FILLER_2_386 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_decap_8 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_2_414 ();
 sg13g2_decap_8 FILLER_2_421 ();
 sg13g2_fill_2 FILLER_2_428 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_fill_1 FILLER_3_70 ();
 sg13g2_fill_1 FILLER_3_115 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_4 FILLER_3_133 ();
 sg13g2_decap_4 FILLER_3_149 ();
 sg13g2_decap_4 FILLER_3_157 ();
 sg13g2_fill_1 FILLER_3_161 ();
 sg13g2_fill_1 FILLER_3_182 ();
 sg13g2_decap_4 FILLER_3_191 ();
 sg13g2_fill_2 FILLER_3_198 ();
 sg13g2_decap_4 FILLER_3_212 ();
 sg13g2_fill_1 FILLER_3_220 ();
 sg13g2_decap_8 FILLER_3_226 ();
 sg13g2_decap_4 FILLER_3_233 ();
 sg13g2_fill_2 FILLER_3_237 ();
 sg13g2_decap_4 FILLER_3_247 ();
 sg13g2_fill_1 FILLER_3_251 ();
 sg13g2_decap_8 FILLER_3_267 ();
 sg13g2_decap_8 FILLER_3_286 ();
 sg13g2_decap_8 FILLER_3_293 ();
 sg13g2_decap_8 FILLER_3_300 ();
 sg13g2_fill_2 FILLER_3_307 ();
 sg13g2_fill_1 FILLER_3_309 ();
 sg13g2_fill_1 FILLER_3_322 ();
 sg13g2_decap_4 FILLER_3_348 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_fill_2 FILLER_4_63 ();
 sg13g2_fill_1 FILLER_4_65 ();
 sg13g2_decap_8 FILLER_4_95 ();
 sg13g2_decap_4 FILLER_4_102 ();
 sg13g2_fill_1 FILLER_4_106 ();
 sg13g2_decap_8 FILLER_4_125 ();
 sg13g2_decap_8 FILLER_4_132 ();
 sg13g2_decap_4 FILLER_4_176 ();
 sg13g2_decap_8 FILLER_4_185 ();
 sg13g2_fill_2 FILLER_4_192 ();
 sg13g2_fill_1 FILLER_4_194 ();
 sg13g2_decap_8 FILLER_4_198 ();
 sg13g2_fill_2 FILLER_4_205 ();
 sg13g2_decap_8 FILLER_4_233 ();
 sg13g2_decap_8 FILLER_4_240 ();
 sg13g2_decap_8 FILLER_4_247 ();
 sg13g2_decap_8 FILLER_4_254 ();
 sg13g2_decap_8 FILLER_4_261 ();
 sg13g2_decap_8 FILLER_4_268 ();
 sg13g2_decap_8 FILLER_4_275 ();
 sg13g2_decap_8 FILLER_4_282 ();
 sg13g2_decap_4 FILLER_4_289 ();
 sg13g2_fill_1 FILLER_4_293 ();
 sg13g2_decap_8 FILLER_4_297 ();
 sg13g2_decap_4 FILLER_4_304 ();
 sg13g2_fill_1 FILLER_4_316 ();
 sg13g2_decap_8 FILLER_4_323 ();
 sg13g2_fill_1 FILLER_4_330 ();
 sg13g2_fill_2 FILLER_4_335 ();
 sg13g2_fill_1 FILLER_4_337 ();
 sg13g2_fill_1 FILLER_4_346 ();
 sg13g2_fill_2 FILLER_4_351 ();
 sg13g2_fill_1 FILLER_4_353 ();
 sg13g2_decap_4 FILLER_4_367 ();
 sg13g2_fill_1 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_377 ();
 sg13g2_decap_4 FILLER_4_384 ();
 sg13g2_fill_2 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_8 FILLER_4_416 ();
 sg13g2_decap_8 FILLER_4_423 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_fill_1 FILLER_5_89 ();
 sg13g2_fill_2 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_125 ();
 sg13g2_decap_8 FILLER_5_132 ();
 sg13g2_fill_2 FILLER_5_139 ();
 sg13g2_decap_8 FILLER_5_145 ();
 sg13g2_decap_8 FILLER_5_152 ();
 sg13g2_decap_8 FILLER_5_159 ();
 sg13g2_decap_4 FILLER_5_166 ();
 sg13g2_decap_8 FILLER_5_208 ();
 sg13g2_decap_4 FILLER_5_215 ();
 sg13g2_fill_1 FILLER_5_219 ();
 sg13g2_decap_8 FILLER_5_249 ();
 sg13g2_fill_2 FILLER_5_317 ();
 sg13g2_fill_1 FILLER_5_319 ();
 sg13g2_fill_2 FILLER_5_324 ();
 sg13g2_fill_1 FILLER_5_348 ();
 sg13g2_fill_2 FILLER_5_353 ();
 sg13g2_fill_1 FILLER_5_355 ();
 sg13g2_fill_2 FILLER_5_364 ();
 sg13g2_fill_2 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_fill_2 FILLER_6_70 ();
 sg13g2_fill_1 FILLER_6_104 ();
 sg13g2_decap_4 FILLER_6_110 ();
 sg13g2_fill_1 FILLER_6_114 ();
 sg13g2_decap_8 FILLER_6_214 ();
 sg13g2_decap_8 FILLER_6_226 ();
 sg13g2_decap_8 FILLER_6_233 ();
 sg13g2_decap_4 FILLER_6_240 ();
 sg13g2_decap_8 FILLER_6_258 ();
 sg13g2_decap_8 FILLER_6_265 ();
 sg13g2_decap_4 FILLER_6_272 ();
 sg13g2_decap_4 FILLER_6_302 ();
 sg13g2_fill_2 FILLER_6_306 ();
 sg13g2_decap_4 FILLER_6_312 ();
 sg13g2_fill_1 FILLER_6_320 ();
 sg13g2_decap_4 FILLER_6_336 ();
 sg13g2_fill_1 FILLER_6_340 ();
 sg13g2_decap_4 FILLER_6_350 ();
 sg13g2_fill_2 FILLER_6_383 ();
 sg13g2_fill_1 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_4 FILLER_7_21 ();
 sg13g2_fill_2 FILLER_7_25 ();
 sg13g2_decap_4 FILLER_7_95 ();
 sg13g2_fill_1 FILLER_7_99 ();
 sg13g2_fill_1 FILLER_7_107 ();
 sg13g2_fill_1 FILLER_7_114 ();
 sg13g2_fill_1 FILLER_7_120 ();
 sg13g2_fill_1 FILLER_7_126 ();
 sg13g2_fill_1 FILLER_7_132 ();
 sg13g2_decap_8 FILLER_7_141 ();
 sg13g2_decap_8 FILLER_7_148 ();
 sg13g2_fill_2 FILLER_7_191 ();
 sg13g2_fill_1 FILLER_7_193 ();
 sg13g2_decap_4 FILLER_7_203 ();
 sg13g2_fill_2 FILLER_7_207 ();
 sg13g2_decap_8 FILLER_7_213 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_fill_2 FILLER_7_280 ();
 sg13g2_fill_1 FILLER_7_282 ();
 sg13g2_decap_4 FILLER_7_288 ();
 sg13g2_fill_1 FILLER_7_292 ();
 sg13g2_fill_2 FILLER_7_306 ();
 sg13g2_fill_1 FILLER_7_308 ();
 sg13g2_fill_2 FILLER_7_313 ();
 sg13g2_fill_2 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_356 ();
 sg13g2_decap_8 FILLER_7_363 ();
 sg13g2_decap_8 FILLER_7_370 ();
 sg13g2_decap_8 FILLER_7_377 ();
 sg13g2_decap_4 FILLER_7_384 ();
 sg13g2_fill_2 FILLER_7_402 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_2 ();
 sg13g2_fill_1 FILLER_8_41 ();
 sg13g2_decap_8 FILLER_8_47 ();
 sg13g2_decap_8 FILLER_8_54 ();
 sg13g2_decap_8 FILLER_8_61 ();
 sg13g2_decap_8 FILLER_8_68 ();
 sg13g2_decap_8 FILLER_8_75 ();
 sg13g2_decap_4 FILLER_8_82 ();
 sg13g2_fill_2 FILLER_8_99 ();
 sg13g2_decap_4 FILLER_8_120 ();
 sg13g2_decap_4 FILLER_8_134 ();
 sg13g2_decap_4 FILLER_8_164 ();
 sg13g2_fill_2 FILLER_8_168 ();
 sg13g2_fill_2 FILLER_8_178 ();
 sg13g2_decap_8 FILLER_8_185 ();
 sg13g2_decap_8 FILLER_8_192 ();
 sg13g2_decap_8 FILLER_8_199 ();
 sg13g2_decap_4 FILLER_8_206 ();
 sg13g2_fill_1 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_decap_4 FILLER_8_256 ();
 sg13g2_fill_1 FILLER_8_260 ();
 sg13g2_decap_4 FILLER_8_271 ();
 sg13g2_fill_2 FILLER_8_275 ();
 sg13g2_decap_8 FILLER_8_290 ();
 sg13g2_decap_4 FILLER_8_297 ();
 sg13g2_fill_1 FILLER_8_301 ();
 sg13g2_decap_4 FILLER_8_333 ();
 sg13g2_fill_2 FILLER_8_337 ();
 sg13g2_fill_2 FILLER_8_343 ();
 sg13g2_fill_1 FILLER_8_345 ();
 sg13g2_decap_8 FILLER_8_351 ();
 sg13g2_decap_8 FILLER_8_358 ();
 sg13g2_decap_8 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_4 FILLER_8_386 ();
 sg13g2_fill_1 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_4 FILLER_8_424 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_71 ();
 sg13g2_decap_8 FILLER_9_78 ();
 sg13g2_decap_8 FILLER_9_85 ();
 sg13g2_decap_8 FILLER_9_92 ();
 sg13g2_decap_8 FILLER_9_99 ();
 sg13g2_decap_8 FILLER_9_106 ();
 sg13g2_fill_1 FILLER_9_113 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_140 ();
 sg13g2_fill_1 FILLER_9_142 ();
 sg13g2_fill_2 FILLER_9_179 ();
 sg13g2_decap_8 FILLER_9_186 ();
 sg13g2_fill_2 FILLER_9_193 ();
 sg13g2_fill_1 FILLER_9_195 ();
 sg13g2_fill_2 FILLER_9_199 ();
 sg13g2_fill_1 FILLER_9_206 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_4 FILLER_9_224 ();
 sg13g2_fill_2 FILLER_9_228 ();
 sg13g2_decap_8 FILLER_9_292 ();
 sg13g2_decap_8 FILLER_9_299 ();
 sg13g2_decap_8 FILLER_9_316 ();
 sg13g2_decap_8 FILLER_9_323 ();
 sg13g2_decap_8 FILLER_9_330 ();
 sg13g2_fill_2 FILLER_9_337 ();
 sg13g2_fill_1 FILLER_9_339 ();
 sg13g2_fill_2 FILLER_9_350 ();
 sg13g2_fill_1 FILLER_9_352 ();
 sg13g2_fill_1 FILLER_9_363 ();
 sg13g2_fill_1 FILLER_9_390 ();
 sg13g2_fill_1 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_fill_2 FILLER_10_40 ();
 sg13g2_fill_1 FILLER_10_42 ();
 sg13g2_fill_2 FILLER_10_54 ();
 sg13g2_fill_1 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_102 ();
 sg13g2_decap_8 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_116 ();
 sg13g2_decap_4 FILLER_10_123 ();
 sg13g2_fill_2 FILLER_10_127 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_fill_1 FILLER_10_204 ();
 sg13g2_fill_2 FILLER_10_211 ();
 sg13g2_fill_1 FILLER_10_234 ();
 sg13g2_decap_8 FILLER_10_239 ();
 sg13g2_decap_8 FILLER_10_246 ();
 sg13g2_decap_4 FILLER_10_253 ();
 sg13g2_fill_2 FILLER_10_257 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_fill_1 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_276 ();
 sg13g2_fill_1 FILLER_10_283 ();
 sg13g2_fill_2 FILLER_10_310 ();
 sg13g2_fill_1 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_339 ();
 sg13g2_fill_2 FILLER_10_346 ();
 sg13g2_decap_8 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_fill_1 FILLER_10_388 ();
 sg13g2_fill_2 FILLER_10_397 ();
 sg13g2_decap_8 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_10_414 ();
 sg13g2_decap_8 FILLER_10_421 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_45 ();
 sg13g2_decap_4 FILLER_11_53 ();
 sg13g2_decap_8 FILLER_11_141 ();
 sg13g2_decap_8 FILLER_11_148 ();
 sg13g2_decap_8 FILLER_11_155 ();
 sg13g2_decap_8 FILLER_11_162 ();
 sg13g2_decap_8 FILLER_11_169 ();
 sg13g2_fill_2 FILLER_11_176 ();
 sg13g2_fill_1 FILLER_11_178 ();
 sg13g2_fill_1 FILLER_11_206 ();
 sg13g2_decap_4 FILLER_11_213 ();
 sg13g2_fill_2 FILLER_11_222 ();
 sg13g2_decap_4 FILLER_11_228 ();
 sg13g2_fill_2 FILLER_11_286 ();
 sg13g2_fill_1 FILLER_11_288 ();
 sg13g2_decap_4 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_4 FILLER_11_319 ();
 sg13g2_decap_4 FILLER_11_328 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_4 FILLER_11_374 ();
 sg13g2_fill_1 FILLER_11_378 ();
 sg13g2_fill_2 FILLER_11_385 ();
 sg13g2_fill_2 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_403 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_fill_2 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_80 ();
 sg13g2_decap_8 FILLER_12_87 ();
 sg13g2_decap_8 FILLER_12_94 ();
 sg13g2_decap_4 FILLER_12_101 ();
 sg13g2_fill_2 FILLER_12_105 ();
 sg13g2_fill_1 FILLER_12_111 ();
 sg13g2_decap_8 FILLER_12_117 ();
 sg13g2_decap_8 FILLER_12_124 ();
 sg13g2_decap_8 FILLER_12_131 ();
 sg13g2_decap_8 FILLER_12_138 ();
 sg13g2_decap_8 FILLER_12_145 ();
 sg13g2_fill_2 FILLER_12_152 ();
 sg13g2_fill_1 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_160 ();
 sg13g2_decap_4 FILLER_12_167 ();
 sg13g2_fill_2 FILLER_12_171 ();
 sg13g2_fill_2 FILLER_12_185 ();
 sg13g2_fill_2 FILLER_12_190 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_fill_1 FILLER_12_214 ();
 sg13g2_decap_8 FILLER_12_226 ();
 sg13g2_decap_8 FILLER_12_233 ();
 sg13g2_decap_8 FILLER_12_240 ();
 sg13g2_decap_8 FILLER_12_247 ();
 sg13g2_decap_8 FILLER_12_254 ();
 sg13g2_decap_4 FILLER_12_261 ();
 sg13g2_fill_2 FILLER_12_265 ();
 sg13g2_fill_2 FILLER_12_280 ();
 sg13g2_fill_1 FILLER_12_282 ();
 sg13g2_fill_1 FILLER_12_288 ();
 sg13g2_fill_2 FILLER_12_293 ();
 sg13g2_fill_1 FILLER_12_295 ();
 sg13g2_decap_8 FILLER_12_313 ();
 sg13g2_decap_4 FILLER_12_320 ();
 sg13g2_fill_1 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_4 FILLER_12_379 ();
 sg13g2_fill_1 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_12_409 ();
 sg13g2_decap_8 FILLER_12_416 ();
 sg13g2_decap_8 FILLER_12_423 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_fill_2 FILLER_13_25 ();
 sg13g2_fill_2 FILLER_13_65 ();
 sg13g2_fill_1 FILLER_13_67 ();
 sg13g2_fill_1 FILLER_13_119 ();
 sg13g2_fill_1 FILLER_13_151 ();
 sg13g2_fill_2 FILLER_13_183 ();
 sg13g2_fill_1 FILLER_13_185 ();
 sg13g2_fill_1 FILLER_13_190 ();
 sg13g2_fill_2 FILLER_13_202 ();
 sg13g2_fill_1 FILLER_13_204 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_fill_1 FILLER_13_266 ();
 sg13g2_fill_2 FILLER_13_275 ();
 sg13g2_fill_1 FILLER_13_277 ();
 sg13g2_fill_1 FILLER_13_290 ();
 sg13g2_fill_1 FILLER_13_295 ();
 sg13g2_decap_8 FILLER_13_309 ();
 sg13g2_decap_8 FILLER_13_316 ();
 sg13g2_decap_8 FILLER_13_323 ();
 sg13g2_decap_8 FILLER_13_330 ();
 sg13g2_decap_8 FILLER_13_337 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_4 FILLER_13_372 ();
 sg13g2_fill_2 FILLER_13_376 ();
 sg13g2_decap_4 FILLER_13_400 ();
 sg13g2_decap_8 FILLER_13_412 ();
 sg13g2_decap_8 FILLER_13_419 ();
 sg13g2_decap_4 FILLER_13_426 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_18 ();
 sg13g2_fill_2 FILLER_14_48 ();
 sg13g2_decap_8 FILLER_14_53 ();
 sg13g2_decap_4 FILLER_14_60 ();
 sg13g2_fill_1 FILLER_14_64 ();
 sg13g2_decap_8 FILLER_14_72 ();
 sg13g2_fill_2 FILLER_14_79 ();
 sg13g2_fill_1 FILLER_14_86 ();
 sg13g2_decap_4 FILLER_14_93 ();
 sg13g2_fill_1 FILLER_14_106 ();
 sg13g2_fill_1 FILLER_14_111 ();
 sg13g2_decap_4 FILLER_14_120 ();
 sg13g2_decap_8 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_141 ();
 sg13g2_fill_2 FILLER_14_148 ();
 sg13g2_fill_1 FILLER_14_150 ();
 sg13g2_decap_4 FILLER_14_156 ();
 sg13g2_fill_1 FILLER_14_160 ();
 sg13g2_decap_8 FILLER_14_174 ();
 sg13g2_decap_4 FILLER_14_181 ();
 sg13g2_fill_1 FILLER_14_185 ();
 sg13g2_fill_1 FILLER_14_199 ();
 sg13g2_decap_4 FILLER_14_205 ();
 sg13g2_decap_8 FILLER_14_214 ();
 sg13g2_fill_2 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_239 ();
 sg13g2_fill_2 FILLER_14_276 ();
 sg13g2_decap_8 FILLER_14_290 ();
 sg13g2_fill_2 FILLER_14_297 ();
 sg13g2_fill_1 FILLER_14_299 ();
 sg13g2_fill_2 FILLER_14_341 ();
 sg13g2_decap_4 FILLER_14_373 ();
 sg13g2_fill_1 FILLER_14_384 ();
 sg13g2_fill_2 FILLER_14_389 ();
 sg13g2_fill_1 FILLER_14_391 ();
 sg13g2_decap_4 FILLER_14_400 ();
 sg13g2_decap_4 FILLER_15_26 ();
 sg13g2_fill_2 FILLER_15_30 ();
 sg13g2_decap_8 FILLER_15_76 ();
 sg13g2_fill_1 FILLER_15_83 ();
 sg13g2_fill_1 FILLER_15_90 ();
 sg13g2_decap_4 FILLER_15_99 ();
 sg13g2_decap_4 FILLER_15_170 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_179 ();
 sg13g2_fill_2 FILLER_15_186 ();
 sg13g2_fill_2 FILLER_15_214 ();
 sg13g2_fill_2 FILLER_15_220 ();
 sg13g2_fill_1 FILLER_15_222 ();
 sg13g2_fill_1 FILLER_15_249 ();
 sg13g2_fill_2 FILLER_15_276 ();
 sg13g2_fill_1 FILLER_15_278 ();
 sg13g2_decap_8 FILLER_15_305 ();
 sg13g2_fill_2 FILLER_15_312 ();
 sg13g2_fill_1 FILLER_15_314 ();
 sg13g2_fill_2 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_fill_1 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_fill_2 FILLER_16_21 ();
 sg13g2_fill_1 FILLER_16_23 ();
 sg13g2_decap_4 FILLER_16_29 ();
 sg13g2_fill_2 FILLER_16_33 ();
 sg13g2_fill_1 FILLER_16_40 ();
 sg13g2_decap_8 FILLER_16_45 ();
 sg13g2_decap_8 FILLER_16_52 ();
 sg13g2_decap_8 FILLER_16_72 ();
 sg13g2_fill_1 FILLER_16_79 ();
 sg13g2_decap_4 FILLER_16_90 ();
 sg13g2_fill_2 FILLER_16_94 ();
 sg13g2_decap_8 FILLER_16_122 ();
 sg13g2_decap_4 FILLER_16_129 ();
 sg13g2_fill_1 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_138 ();
 sg13g2_decap_4 FILLER_16_145 ();
 sg13g2_fill_1 FILLER_16_149 ();
 sg13g2_fill_1 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_163 ();
 sg13g2_decap_8 FILLER_16_170 ();
 sg13g2_decap_4 FILLER_16_177 ();
 sg13g2_fill_2 FILLER_16_181 ();
 sg13g2_decap_8 FILLER_16_191 ();
 sg13g2_decap_4 FILLER_16_198 ();
 sg13g2_decap_8 FILLER_16_206 ();
 sg13g2_decap_8 FILLER_16_213 ();
 sg13g2_decap_8 FILLER_16_220 ();
 sg13g2_decap_4 FILLER_16_227 ();
 sg13g2_fill_1 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_242 ();
 sg13g2_fill_2 FILLER_16_249 ();
 sg13g2_fill_1 FILLER_16_251 ();
 sg13g2_fill_2 FILLER_16_274 ();
 sg13g2_decap_4 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_288 ();
 sg13g2_decap_4 FILLER_16_332 ();
 sg13g2_fill_2 FILLER_16_336 ();
 sg13g2_fill_2 FILLER_16_346 ();
 sg13g2_fill_1 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_fill_1 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_16_412 ();
 sg13g2_decap_8 FILLER_16_419 ();
 sg13g2_decap_4 FILLER_16_426 ();
 sg13g2_fill_2 FILLER_17_46 ();
 sg13g2_decap_4 FILLER_17_78 ();
 sg13g2_fill_2 FILLER_17_82 ();
 sg13g2_decap_8 FILLER_17_103 ();
 sg13g2_fill_2 FILLER_17_110 ();
 sg13g2_decap_8 FILLER_17_116 ();
 sg13g2_decap_4 FILLER_17_123 ();
 sg13g2_fill_1 FILLER_17_127 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_161 ();
 sg13g2_fill_1 FILLER_17_163 ();
 sg13g2_decap_8 FILLER_17_190 ();
 sg13g2_decap_8 FILLER_17_197 ();
 sg13g2_fill_2 FILLER_17_204 ();
 sg13g2_decap_8 FILLER_17_236 ();
 sg13g2_fill_2 FILLER_17_243 ();
 sg13g2_fill_1 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_272 ();
 sg13g2_fill_2 FILLER_17_284 ();
 sg13g2_fill_1 FILLER_17_295 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_fill_2 FILLER_17_307 ();
 sg13g2_fill_1 FILLER_17_309 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_332 ();
 sg13g2_fill_2 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_4 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_fill_2 FILLER_17_380 ();
 sg13g2_fill_1 FILLER_17_394 ();
 sg13g2_fill_1 FILLER_17_403 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_4 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_64 ();
 sg13g2_decap_8 FILLER_18_71 ();
 sg13g2_decap_8 FILLER_18_78 ();
 sg13g2_decap_8 FILLER_18_93 ();
 sg13g2_decap_4 FILLER_18_100 ();
 sg13g2_decap_8 FILLER_18_109 ();
 sg13g2_fill_1 FILLER_18_116 ();
 sg13g2_decap_8 FILLER_18_122 ();
 sg13g2_fill_2 FILLER_18_129 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_decap_4 FILLER_18_146 ();
 sg13g2_fill_2 FILLER_18_150 ();
 sg13g2_fill_1 FILLER_18_157 ();
 sg13g2_decap_4 FILLER_18_167 ();
 sg13g2_fill_2 FILLER_18_180 ();
 sg13g2_decap_8 FILLER_18_208 ();
 sg13g2_decap_8 FILLER_18_215 ();
 sg13g2_decap_4 FILLER_18_222 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_4 FILLER_18_259 ();
 sg13g2_fill_1 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_313 ();
 sg13g2_decap_8 FILLER_18_331 ();
 sg13g2_fill_1 FILLER_18_338 ();
 sg13g2_decap_8 FILLER_18_365 ();
 sg13g2_fill_2 FILLER_18_372 ();
 sg13g2_fill_1 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_fill_2 FILLER_18_427 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_decap_4 FILLER_19_29 ();
 sg13g2_decap_8 FILLER_19_41 ();
 sg13g2_decap_4 FILLER_19_48 ();
 sg13g2_decap_8 FILLER_19_62 ();
 sg13g2_decap_8 FILLER_19_69 ();
 sg13g2_decap_4 FILLER_19_107 ();
 sg13g2_fill_2 FILLER_19_116 ();
 sg13g2_fill_2 FILLER_19_123 ();
 sg13g2_fill_2 FILLER_19_130 ();
 sg13g2_decap_4 FILLER_19_158 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_decap_8 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_188 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_4 FILLER_19_211 ();
 sg13g2_decap_8 FILLER_19_239 ();
 sg13g2_decap_8 FILLER_19_246 ();
 sg13g2_decap_8 FILLER_19_253 ();
 sg13g2_decap_4 FILLER_19_260 ();
 sg13g2_decap_8 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_275 ();
 sg13g2_decap_8 FILLER_19_282 ();
 sg13g2_decap_4 FILLER_19_289 ();
 sg13g2_fill_1 FILLER_19_293 ();
 sg13g2_fill_2 FILLER_19_313 ();
 sg13g2_decap_4 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_327 ();
 sg13g2_decap_8 FILLER_19_334 ();
 sg13g2_fill_2 FILLER_19_341 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_fill_1 FILLER_19_361 ();
 sg13g2_fill_2 FILLER_19_369 ();
 sg13g2_fill_1 FILLER_19_390 ();
 sg13g2_fill_1 FILLER_19_404 ();
 sg13g2_decap_8 FILLER_19_409 ();
 sg13g2_decap_8 FILLER_19_416 ();
 sg13g2_decap_8 FILLER_19_423 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_11 ();
 sg13g2_fill_1 FILLER_20_16 ();
 sg13g2_fill_1 FILLER_20_29 ();
 sg13g2_fill_1 FILLER_20_36 ();
 sg13g2_fill_2 FILLER_20_45 ();
 sg13g2_decap_4 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_69 ();
 sg13g2_decap_8 FILLER_20_80 ();
 sg13g2_decap_8 FILLER_20_87 ();
 sg13g2_decap_4 FILLER_20_94 ();
 sg13g2_fill_2 FILLER_20_114 ();
 sg13g2_fill_1 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_121 ();
 sg13g2_fill_2 FILLER_20_128 ();
 sg13g2_fill_1 FILLER_20_130 ();
 sg13g2_decap_8 FILLER_20_136 ();
 sg13g2_decap_8 FILLER_20_143 ();
 sg13g2_decap_8 FILLER_20_150 ();
 sg13g2_decap_8 FILLER_20_157 ();
 sg13g2_decap_4 FILLER_20_164 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_fill_2 FILLER_20_218 ();
 sg13g2_decap_8 FILLER_20_233 ();
 sg13g2_fill_2 FILLER_20_240 ();
 sg13g2_fill_1 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_269 ();
 sg13g2_decap_8 FILLER_20_276 ();
 sg13g2_fill_1 FILLER_20_283 ();
 sg13g2_fill_2 FILLER_20_296 ();
 sg13g2_fill_1 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_304 ();
 sg13g2_fill_1 FILLER_20_311 ();
 sg13g2_fill_1 FILLER_20_317 ();
 sg13g2_fill_2 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_19 ();
 sg13g2_fill_1 FILLER_21_25 ();
 sg13g2_fill_1 FILLER_21_38 ();
 sg13g2_fill_1 FILLER_21_43 ();
 sg13g2_fill_1 FILLER_21_47 ();
 sg13g2_fill_2 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_85 ();
 sg13g2_fill_2 FILLER_21_92 ();
 sg13g2_decap_8 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_116 ();
 sg13g2_decap_8 FILLER_21_128 ();
 sg13g2_decap_8 FILLER_21_135 ();
 sg13g2_decap_8 FILLER_21_142 ();
 sg13g2_fill_1 FILLER_21_149 ();
 sg13g2_fill_2 FILLER_21_194 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_fill_2 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_227 ();
 sg13g2_decap_8 FILLER_21_246 ();
 sg13g2_decap_4 FILLER_21_253 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_decap_4 FILLER_21_297 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_4 FILLER_21_350 ();
 sg13g2_fill_1 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_359 ();
 sg13g2_fill_2 FILLER_21_366 ();
 sg13g2_fill_2 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_423 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_11 ();
 sg13g2_fill_2 FILLER_22_79 ();
 sg13g2_fill_1 FILLER_22_86 ();
 sg13g2_decap_8 FILLER_22_92 ();
 sg13g2_decap_8 FILLER_22_99 ();
 sg13g2_fill_2 FILLER_22_106 ();
 sg13g2_fill_1 FILLER_22_108 ();
 sg13g2_fill_1 FILLER_22_143 ();
 sg13g2_decap_4 FILLER_22_174 ();
 sg13g2_fill_1 FILLER_22_183 ();
 sg13g2_decap_8 FILLER_22_214 ();
 sg13g2_fill_1 FILLER_22_221 ();
 sg13g2_fill_1 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_248 ();
 sg13g2_decap_8 FILLER_22_255 ();
 sg13g2_decap_8 FILLER_22_262 ();
 sg13g2_decap_8 FILLER_22_269 ();
 sg13g2_decap_8 FILLER_22_276 ();
 sg13g2_decap_4 FILLER_22_283 ();
 sg13g2_fill_2 FILLER_22_287 ();
 sg13g2_decap_4 FILLER_22_294 ();
 sg13g2_decap_4 FILLER_22_307 ();
 sg13g2_decap_8 FILLER_22_345 ();
 sg13g2_fill_1 FILLER_22_352 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_4 FILLER_22_375 ();
 sg13g2_fill_2 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_409 ();
 sg13g2_decap_8 FILLER_22_416 ();
 sg13g2_decap_8 FILLER_22_423 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_31 ();
 sg13g2_decap_8 FILLER_23_38 ();
 sg13g2_fill_2 FILLER_23_45 ();
 sg13g2_fill_2 FILLER_23_51 ();
 sg13g2_fill_1 FILLER_23_53 ();
 sg13g2_fill_2 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_78 ();
 sg13g2_decap_4 FILLER_23_85 ();
 sg13g2_decap_8 FILLER_23_94 ();
 sg13g2_decap_8 FILLER_23_101 ();
 sg13g2_decap_8 FILLER_23_108 ();
 sg13g2_decap_4 FILLER_23_115 ();
 sg13g2_fill_1 FILLER_23_119 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_decap_8 FILLER_23_149 ();
 sg13g2_decap_8 FILLER_23_156 ();
 sg13g2_decap_8 FILLER_23_163 ();
 sg13g2_fill_2 FILLER_23_170 ();
 sg13g2_decap_8 FILLER_23_198 ();
 sg13g2_decap_8 FILLER_23_205 ();
 sg13g2_decap_8 FILLER_23_212 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_234 ();
 sg13g2_decap_4 FILLER_23_240 ();
 sg13g2_decap_4 FILLER_23_278 ();
 sg13g2_fill_1 FILLER_23_282 ();
 sg13g2_fill_2 FILLER_23_288 ();
 sg13g2_fill_1 FILLER_23_290 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_fill_2 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_325 ();
 sg13g2_decap_8 FILLER_23_332 ();
 sg13g2_decap_4 FILLER_23_339 ();
 sg13g2_fill_1 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_decap_8 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_23_409 ();
 sg13g2_decap_8 FILLER_23_416 ();
 sg13g2_decap_8 FILLER_23_423 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_fill_1 FILLER_24_59 ();
 sg13g2_decap_8 FILLER_24_72 ();
 sg13g2_decap_4 FILLER_24_79 ();
 sg13g2_fill_1 FILLER_24_83 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_1 FILLER_24_125 ();
 sg13g2_decap_4 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_140 ();
 sg13g2_decap_4 FILLER_24_146 ();
 sg13g2_fill_1 FILLER_24_150 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_4 FILLER_24_175 ();
 sg13g2_fill_2 FILLER_24_179 ();
 sg13g2_fill_2 FILLER_24_216 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_decap_8 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_256 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_decap_4 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_293 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_decap_4 FILLER_24_347 ();
 sg13g2_fill_2 FILLER_24_351 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_8 FILLER_24_404 ();
 sg13g2_decap_8 FILLER_24_411 ();
 sg13g2_decap_8 FILLER_24_418 ();
 sg13g2_decap_4 FILLER_24_425 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_1 FILLER_25_37 ();
 sg13g2_decap_8 FILLER_25_62 ();
 sg13g2_fill_1 FILLER_25_69 ();
 sg13g2_decap_8 FILLER_25_75 ();
 sg13g2_decap_8 FILLER_25_82 ();
 sg13g2_decap_8 FILLER_25_89 ();
 sg13g2_decap_8 FILLER_25_96 ();
 sg13g2_decap_4 FILLER_25_108 ();
 sg13g2_fill_1 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_149 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_decap_4 FILLER_25_191 ();
 sg13g2_decap_8 FILLER_25_199 ();
 sg13g2_decap_8 FILLER_25_206 ();
 sg13g2_fill_2 FILLER_25_221 ();
 sg13g2_fill_2 FILLER_25_228 ();
 sg13g2_fill_1 FILLER_25_230 ();
 sg13g2_decap_4 FILLER_25_295 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_324 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_8 FILLER_25_338 ();
 sg13g2_decap_8 FILLER_25_345 ();
 sg13g2_fill_2 FILLER_25_352 ();
 sg13g2_fill_1 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_404 ();
 sg13g2_decap_8 FILLER_25_411 ();
 sg13g2_decap_8 FILLER_25_418 ();
 sg13g2_decap_4 FILLER_25_425 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_11 ();
 sg13g2_fill_2 FILLER_26_17 ();
 sg13g2_fill_1 FILLER_26_19 ();
 sg13g2_decap_8 FILLER_26_41 ();
 sg13g2_decap_8 FILLER_26_48 ();
 sg13g2_decap_4 FILLER_26_55 ();
 sg13g2_fill_2 FILLER_26_59 ();
 sg13g2_decap_8 FILLER_26_85 ();
 sg13g2_decap_4 FILLER_26_92 ();
 sg13g2_decap_8 FILLER_26_122 ();
 sg13g2_decap_8 FILLER_26_129 ();
 sg13g2_fill_2 FILLER_26_136 ();
 sg13g2_fill_1 FILLER_26_138 ();
 sg13g2_fill_2 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_decap_8 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_202 ();
 sg13g2_decap_4 FILLER_26_208 ();
 sg13g2_decap_8 FILLER_26_247 ();
 sg13g2_decap_4 FILLER_26_254 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_fill_2 FILLER_26_304 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_fill_2 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_414 ();
 sg13g2_decap_8 FILLER_26_421 ();
 sg13g2_fill_2 FILLER_26_428 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_41 ();
 sg13g2_fill_2 FILLER_27_52 ();
 sg13g2_fill_2 FILLER_27_58 ();
 sg13g2_fill_2 FILLER_27_83 ();
 sg13g2_fill_2 FILLER_27_90 ();
 sg13g2_fill_1 FILLER_27_92 ();
 sg13g2_decap_8 FILLER_27_97 ();
 sg13g2_fill_2 FILLER_27_104 ();
 sg13g2_fill_1 FILLER_27_106 ();
 sg13g2_decap_4 FILLER_27_110 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_fill_1 FILLER_27_120 ();
 sg13g2_decap_4 FILLER_27_125 ();
 sg13g2_fill_1 FILLER_27_129 ();
 sg13g2_fill_1 FILLER_27_139 ();
 sg13g2_fill_2 FILLER_27_166 ();
 sg13g2_decap_8 FILLER_27_204 ();
 sg13g2_decap_8 FILLER_27_211 ();
 sg13g2_decap_8 FILLER_27_218 ();
 sg13g2_decap_8 FILLER_27_225 ();
 sg13g2_fill_2 FILLER_27_232 ();
 sg13g2_fill_1 FILLER_27_234 ();
 sg13g2_decap_8 FILLER_27_239 ();
 sg13g2_fill_2 FILLER_27_308 ();
 sg13g2_fill_2 FILLER_27_315 ();
 sg13g2_fill_1 FILLER_27_317 ();
 sg13g2_decap_4 FILLER_27_322 ();
 sg13g2_fill_2 FILLER_27_352 ();
 sg13g2_fill_1 FILLER_27_354 ();
 sg13g2_fill_1 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_decap_8 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_27_414 ();
 sg13g2_decap_8 FILLER_27_421 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_33 ();
 sg13g2_decap_8 FILLER_28_40 ();
 sg13g2_decap_8 FILLER_28_47 ();
 sg13g2_fill_1 FILLER_28_54 ();
 sg13g2_decap_8 FILLER_28_81 ();
 sg13g2_fill_1 FILLER_28_124 ();
 sg13g2_decap_8 FILLER_28_146 ();
 sg13g2_decap_4 FILLER_28_153 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_decap_4 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_172 ();
 sg13g2_fill_2 FILLER_28_178 ();
 sg13g2_decap_8 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_201 ();
 sg13g2_decap_8 FILLER_28_206 ();
 sg13g2_decap_8 FILLER_28_213 ();
 sg13g2_decap_8 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_227 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_fill_2 FILLER_28_292 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_319 ();
 sg13g2_decap_4 FILLER_28_324 ();
 sg13g2_fill_2 FILLER_28_328 ();
 sg13g2_decap_4 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_fill_2 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_fill_2 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_23 ();
 sg13g2_fill_2 FILLER_29_70 ();
 sg13g2_fill_2 FILLER_29_90 ();
 sg13g2_fill_1 FILLER_29_92 ();
 sg13g2_decap_8 FILLER_29_96 ();
 sg13g2_decap_8 FILLER_29_103 ();
 sg13g2_decap_8 FILLER_29_110 ();
 sg13g2_decap_8 FILLER_29_117 ();
 sg13g2_fill_2 FILLER_29_124 ();
 sg13g2_fill_1 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_132 ();
 sg13g2_fill_1 FILLER_29_165 ();
 sg13g2_decap_4 FILLER_29_190 ();
 sg13g2_decap_8 FILLER_29_220 ();
 sg13g2_decap_4 FILLER_29_227 ();
 sg13g2_decap_8 FILLER_29_240 ();
 sg13g2_fill_2 FILLER_29_247 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_decap_8 FILLER_29_260 ();
 sg13g2_decap_8 FILLER_29_267 ();
 sg13g2_decap_8 FILLER_29_279 ();
 sg13g2_decap_8 FILLER_29_286 ();
 sg13g2_decap_4 FILLER_29_293 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_309 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_decap_8 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_29_327 ();
 sg13g2_fill_2 FILLER_29_334 ();
 sg13g2_fill_2 FILLER_29_340 ();
 sg13g2_fill_1 FILLER_29_342 ();
 sg13g2_decap_4 FILLER_29_352 ();
 sg13g2_fill_2 FILLER_29_356 ();
 sg13g2_fill_1 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_86 ();
 sg13g2_decap_8 FILLER_30_93 ();
 sg13g2_decap_4 FILLER_30_100 ();
 sg13g2_fill_2 FILLER_30_104 ();
 sg13g2_decap_4 FILLER_30_132 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_decap_8 FILLER_30_145 ();
 sg13g2_decap_4 FILLER_30_152 ();
 sg13g2_fill_2 FILLER_30_156 ();
 sg13g2_fill_1 FILLER_30_163 ();
 sg13g2_decap_8 FILLER_30_184 ();
 sg13g2_decap_8 FILLER_30_191 ();
 sg13g2_decap_8 FILLER_30_198 ();
 sg13g2_decap_8 FILLER_30_205 ();
 sg13g2_decap_4 FILLER_30_212 ();
 sg13g2_fill_2 FILLER_30_216 ();
 sg13g2_decap_4 FILLER_30_222 ();
 sg13g2_fill_1 FILLER_30_226 ();
 sg13g2_fill_2 FILLER_30_246 ();
 sg13g2_fill_1 FILLER_30_248 ();
 sg13g2_decap_8 FILLER_30_290 ();
 sg13g2_decap_4 FILLER_30_297 ();
 sg13g2_fill_1 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_370 ();
 sg13g2_fill_2 FILLER_30_377 ();
 sg13g2_fill_1 FILLER_30_379 ();
 sg13g2_decap_4 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_33 ();
 sg13g2_decap_8 FILLER_31_48 ();
 sg13g2_decap_8 FILLER_31_55 ();
 sg13g2_decap_8 FILLER_31_62 ();
 sg13g2_decap_4 FILLER_31_69 ();
 sg13g2_fill_2 FILLER_31_73 ();
 sg13g2_decap_4 FILLER_31_101 ();
 sg13g2_fill_1 FILLER_31_105 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_129 ();
 sg13g2_fill_1 FILLER_31_136 ();
 sg13g2_decap_4 FILLER_31_142 ();
 sg13g2_fill_2 FILLER_31_146 ();
 sg13g2_decap_4 FILLER_31_161 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_fill_1 FILLER_31_182 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_decap_8 FILLER_31_205 ();
 sg13g2_fill_2 FILLER_31_212 ();
 sg13g2_fill_1 FILLER_31_236 ();
 sg13g2_decap_4 FILLER_31_249 ();
 sg13g2_decap_8 FILLER_31_261 ();
 sg13g2_decap_8 FILLER_31_268 ();
 sg13g2_decap_4 FILLER_31_275 ();
 sg13g2_decap_8 FILLER_31_284 ();
 sg13g2_decap_8 FILLER_31_291 ();
 sg13g2_fill_1 FILLER_31_298 ();
 sg13g2_decap_8 FILLER_31_309 ();
 sg13g2_decap_4 FILLER_31_320 ();
 sg13g2_fill_1 FILLER_31_324 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_fill_2 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_345 ();
 sg13g2_decap_8 FILLER_31_351 ();
 sg13g2_decap_4 FILLER_31_358 ();
 sg13g2_decap_8 FILLER_31_367 ();
 sg13g2_fill_2 FILLER_31_374 ();
 sg13g2_fill_1 FILLER_31_376 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_406 ();
 sg13g2_decap_8 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_fill_2 FILLER_31_427 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_4 FILLER_32_26 ();
 sg13g2_fill_1 FILLER_32_30 ();
 sg13g2_decap_8 FILLER_32_44 ();
 sg13g2_decap_8 FILLER_32_51 ();
 sg13g2_decap_8 FILLER_32_58 ();
 sg13g2_decap_8 FILLER_32_65 ();
 sg13g2_decap_8 FILLER_32_72 ();
 sg13g2_decap_8 FILLER_32_79 ();
 sg13g2_decap_8 FILLER_32_86 ();
 sg13g2_decap_4 FILLER_32_93 ();
 sg13g2_fill_2 FILLER_32_97 ();
 sg13g2_decap_4 FILLER_32_111 ();
 sg13g2_decap_4 FILLER_32_119 ();
 sg13g2_fill_2 FILLER_32_130 ();
 sg13g2_decap_8 FILLER_32_146 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_fill_2 FILLER_32_161 ();
 sg13g2_fill_2 FILLER_32_173 ();
 sg13g2_fill_1 FILLER_32_175 ();
 sg13g2_fill_1 FILLER_32_180 ();
 sg13g2_fill_2 FILLER_32_187 ();
 sg13g2_decap_4 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_fill_2 FILLER_32_226 ();
 sg13g2_fill_1 FILLER_32_228 ();
 sg13g2_decap_4 FILLER_32_234 ();
 sg13g2_fill_2 FILLER_32_244 ();
 sg13g2_fill_1 FILLER_32_246 ();
 sg13g2_fill_2 FILLER_32_259 ();
 sg13g2_fill_1 FILLER_32_261 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_fill_2 FILLER_32_299 ();
 sg13g2_fill_1 FILLER_32_335 ();
 sg13g2_fill_2 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_346 ();
 sg13g2_fill_1 FILLER_32_389 ();
 sg13g2_decap_8 FILLER_32_416 ();
 sg13g2_decap_8 FILLER_32_423 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_58 ();
 sg13g2_decap_8 FILLER_33_65 ();
 sg13g2_fill_2 FILLER_33_72 ();
 sg13g2_decap_8 FILLER_33_82 ();
 sg13g2_fill_2 FILLER_33_89 ();
 sg13g2_fill_1 FILLER_33_117 ();
 sg13g2_fill_2 FILLER_33_154 ();
 sg13g2_fill_1 FILLER_33_156 ();
 sg13g2_fill_2 FILLER_33_162 ();
 sg13g2_fill_1 FILLER_33_164 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_200 ();
 sg13g2_fill_1 FILLER_33_216 ();
 sg13g2_fill_1 FILLER_33_222 ();
 sg13g2_fill_1 FILLER_33_228 ();
 sg13g2_fill_2 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_239 ();
 sg13g2_fill_1 FILLER_33_248 ();
 sg13g2_decap_4 FILLER_33_256 ();
 sg13g2_decap_8 FILLER_33_268 ();
 sg13g2_decap_8 FILLER_33_275 ();
 sg13g2_decap_8 FILLER_33_282 ();
 sg13g2_decap_8 FILLER_33_289 ();
 sg13g2_decap_8 FILLER_33_296 ();
 sg13g2_decap_8 FILLER_33_303 ();
 sg13g2_decap_8 FILLER_33_310 ();
 sg13g2_decap_8 FILLER_33_321 ();
 sg13g2_fill_1 FILLER_33_328 ();
 sg13g2_decap_8 FILLER_33_342 ();
 sg13g2_decap_8 FILLER_33_349 ();
 sg13g2_decap_8 FILLER_33_356 ();
 sg13g2_fill_2 FILLER_33_363 ();
 sg13g2_decap_4 FILLER_33_370 ();
 sg13g2_fill_2 FILLER_33_374 ();
 sg13g2_fill_1 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_395 ();
 sg13g2_fill_2 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_33_409 ();
 sg13g2_decap_8 FILLER_33_416 ();
 sg13g2_decap_8 FILLER_33_423 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_11 ();
 sg13g2_decap_4 FILLER_34_20 ();
 sg13g2_fill_2 FILLER_34_24 ();
 sg13g2_decap_8 FILLER_34_40 ();
 sg13g2_decap_8 FILLER_34_47 ();
 sg13g2_decap_4 FILLER_34_54 ();
 sg13g2_decap_8 FILLER_34_96 ();
 sg13g2_decap_8 FILLER_34_103 ();
 sg13g2_decap_4 FILLER_34_110 ();
 sg13g2_fill_2 FILLER_34_114 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_fill_1 FILLER_34_140 ();
 sg13g2_decap_4 FILLER_34_145 ();
 sg13g2_fill_2 FILLER_34_149 ();
 sg13g2_fill_1 FILLER_34_159 ();
 sg13g2_decap_8 FILLER_34_167 ();
 sg13g2_decap_8 FILLER_34_174 ();
 sg13g2_decap_8 FILLER_34_181 ();
 sg13g2_fill_2 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_190 ();
 sg13g2_decap_8 FILLER_34_205 ();
 sg13g2_fill_2 FILLER_34_212 ();
 sg13g2_fill_1 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_220 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_fill_1 FILLER_34_230 ();
 sg13g2_decap_4 FILLER_34_236 ();
 sg13g2_fill_2 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_263 ();
 sg13g2_fill_1 FILLER_34_270 ();
 sg13g2_fill_2 FILLER_34_276 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_decap_8 FILLER_34_317 ();
 sg13g2_decap_8 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_331 ();
 sg13g2_decap_4 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_decap_8 FILLER_34_370 ();
 sg13g2_fill_2 FILLER_34_377 ();
 sg13g2_fill_1 FILLER_34_379 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_34_409 ();
 sg13g2_decap_8 FILLER_34_416 ();
 sg13g2_decap_8 FILLER_34_423 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_17 ();
 sg13g2_decap_4 FILLER_35_24 ();
 sg13g2_fill_2 FILLER_35_28 ();
 sg13g2_decap_4 FILLER_35_36 ();
 sg13g2_fill_1 FILLER_35_40 ();
 sg13g2_decap_8 FILLER_35_53 ();
 sg13g2_decap_8 FILLER_35_60 ();
 sg13g2_decap_4 FILLER_35_67 ();
 sg13g2_decap_8 FILLER_35_94 ();
 sg13g2_decap_8 FILLER_35_101 ();
 sg13g2_fill_1 FILLER_35_108 ();
 sg13g2_decap_8 FILLER_35_129 ();
 sg13g2_decap_8 FILLER_35_136 ();
 sg13g2_fill_2 FILLER_35_143 ();
 sg13g2_fill_1 FILLER_35_145 ();
 sg13g2_decap_4 FILLER_35_151 ();
 sg13g2_fill_2 FILLER_35_180 ();
 sg13g2_decap_8 FILLER_35_190 ();
 sg13g2_decap_8 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_208 ();
 sg13g2_fill_2 FILLER_35_215 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_4 FILLER_35_238 ();
 sg13g2_fill_1 FILLER_35_242 ();
 sg13g2_decap_8 FILLER_35_247 ();
 sg13g2_decap_8 FILLER_35_258 ();
 sg13g2_decap_8 FILLER_35_278 ();
 sg13g2_fill_1 FILLER_35_293 ();
 sg13g2_fill_2 FILLER_35_320 ();
 sg13g2_fill_1 FILLER_35_348 ();
 sg13g2_decap_4 FILLER_35_379 ();
 sg13g2_fill_1 FILLER_35_383 ();
 sg13g2_fill_1 FILLER_35_392 ();
 sg13g2_fill_2 FILLER_35_398 ();
 sg13g2_decap_8 FILLER_35_404 ();
 sg13g2_decap_8 FILLER_35_411 ();
 sg13g2_decap_8 FILLER_35_418 ();
 sg13g2_decap_4 FILLER_35_425 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_4 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_46 ();
 sg13g2_decap_8 FILLER_36_73 ();
 sg13g2_decap_8 FILLER_36_88 ();
 sg13g2_decap_8 FILLER_36_95 ();
 sg13g2_fill_1 FILLER_36_102 ();
 sg13g2_fill_2 FILLER_36_156 ();
 sg13g2_decap_8 FILLER_36_162 ();
 sg13g2_decap_8 FILLER_36_174 ();
 sg13g2_decap_8 FILLER_36_181 ();
 sg13g2_decap_8 FILLER_36_192 ();
 sg13g2_decap_8 FILLER_36_199 ();
 sg13g2_fill_1 FILLER_36_206 ();
 sg13g2_fill_1 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_294 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_decap_8 FILLER_36_313 ();
 sg13g2_fill_2 FILLER_36_320 ();
 sg13g2_fill_1 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_328 ();
 sg13g2_decap_8 FILLER_36_335 ();
 sg13g2_decap_8 FILLER_36_342 ();
 sg13g2_decap_8 FILLER_36_349 ();
 sg13g2_fill_1 FILLER_36_356 ();
 sg13g2_fill_1 FILLER_36_365 ();
 sg13g2_fill_2 FILLER_36_375 ();
 sg13g2_fill_1 FILLER_36_377 ();
 sg13g2_fill_2 FILLER_36_383 ();
 sg13g2_fill_1 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_416 ();
 sg13g2_decap_8 FILLER_36_423 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_17 ();
 sg13g2_decap_8 FILLER_37_24 ();
 sg13g2_fill_2 FILLER_37_31 ();
 sg13g2_fill_1 FILLER_37_33 ();
 sg13g2_fill_2 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_52 ();
 sg13g2_decap_8 FILLER_37_59 ();
 sg13g2_fill_1 FILLER_37_71 ();
 sg13g2_fill_1 FILLER_37_76 ();
 sg13g2_fill_1 FILLER_37_103 ();
 sg13g2_fill_1 FILLER_37_117 ();
 sg13g2_fill_2 FILLER_37_122 ();
 sg13g2_fill_1 FILLER_37_124 ();
 sg13g2_fill_2 FILLER_37_129 ();
 sg13g2_fill_1 FILLER_37_135 ();
 sg13g2_fill_1 FILLER_37_144 ();
 sg13g2_fill_1 FILLER_37_150 ();
 sg13g2_fill_2 FILLER_37_155 ();
 sg13g2_fill_2 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_193 ();
 sg13g2_fill_1 FILLER_37_200 ();
 sg13g2_fill_1 FILLER_37_206 ();
 sg13g2_fill_1 FILLER_37_211 ();
 sg13g2_fill_2 FILLER_37_216 ();
 sg13g2_fill_2 FILLER_37_223 ();
 sg13g2_fill_2 FILLER_37_229 ();
 sg13g2_fill_1 FILLER_37_231 ();
 sg13g2_fill_2 FILLER_37_244 ();
 sg13g2_fill_1 FILLER_37_246 ();
 sg13g2_decap_4 FILLER_37_290 ();
 sg13g2_fill_2 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_304 ();
 sg13g2_decap_8 FILLER_37_309 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_fill_1 FILLER_37_365 ();
 sg13g2_fill_2 FILLER_37_374 ();
 sg13g2_fill_1 FILLER_37_376 ();
 sg13g2_fill_2 FILLER_37_382 ();
 sg13g2_fill_1 FILLER_37_384 ();
 sg13g2_decap_8 FILLER_37_416 ();
 sg13g2_decap_8 FILLER_37_423 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_14 ();
 sg13g2_decap_4 FILLER_38_41 ();
 sg13g2_fill_2 FILLER_38_45 ();
 sg13g2_fill_1 FILLER_38_85 ();
 sg13g2_fill_1 FILLER_38_106 ();
 sg13g2_fill_2 FILLER_38_111 ();
 sg13g2_fill_2 FILLER_38_121 ();
 sg13g2_fill_1 FILLER_38_153 ();
 sg13g2_decap_4 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_260 ();
 sg13g2_decap_8 FILLER_38_267 ();
 sg13g2_decap_8 FILLER_38_274 ();
 sg13g2_decap_8 FILLER_38_281 ();
 sg13g2_decap_8 FILLER_38_288 ();
 sg13g2_decap_4 FILLER_38_295 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_4 FILLER_38_350 ();
 sg13g2_fill_1 FILLER_38_354 ();
 sg13g2_fill_2 FILLER_38_381 ();
 sg13g2_fill_1 FILLER_38_395 ();
 sg13g2_fill_1 FILLER_38_400 ();
 sg13g2_fill_1 FILLER_38_405 ();
 sg13g2_decap_8 FILLER_38_410 ();
 sg13g2_decap_8 FILLER_38_417 ();
 sg13g2_decap_4 FILLER_38_424 ();
 sg13g2_fill_2 FILLER_38_428 ();
endmodule
