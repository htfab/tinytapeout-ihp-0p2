module tt_um_frequency_counter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire clknet_0_clk;
 wire \frequency_counter.clk_counter[0] ;
 wire \frequency_counter.clk_counter[10] ;
 wire \frequency_counter.clk_counter[11] ;
 wire \frequency_counter.clk_counter[1] ;
 wire \frequency_counter.clk_counter[2] ;
 wire \frequency_counter.clk_counter[3] ;
 wire \frequency_counter.clk_counter[4] ;
 wire \frequency_counter.clk_counter[5] ;
 wire \frequency_counter.clk_counter[6] ;
 wire \frequency_counter.clk_counter[7] ;
 wire \frequency_counter.clk_counter[8] ;
 wire \frequency_counter.clk_counter[9] ;
 wire \frequency_counter.digit ;
 wire \frequency_counter.edge_counter[0] ;
 wire \frequency_counter.edge_counter[1] ;
 wire \frequency_counter.edge_counter[2] ;
 wire \frequency_counter.edge_counter[3] ;
 wire \frequency_counter.edge_counter[4] ;
 wire \frequency_counter.edge_counter[5] ;
 wire \frequency_counter.edge_counter[6] ;
 wire \frequency_counter.edge_detect0.q0 ;
 wire \frequency_counter.edge_detect0.q1 ;
 wire \frequency_counter.edge_detect0.q2 ;
 wire \frequency_counter.seven_segment0.load ;
 wire \frequency_counter.seven_segment0.ten_count[0] ;
 wire \frequency_counter.seven_segment0.ten_count[1] ;
 wire \frequency_counter.seven_segment0.ten_count[2] ;
 wire \frequency_counter.seven_segment0.ten_count[3] ;
 wire \frequency_counter.seven_segment0.ten_count_reg[0] ;
 wire \frequency_counter.seven_segment0.ten_count_reg[1] ;
 wire \frequency_counter.seven_segment0.ten_count_reg[2] ;
 wire \frequency_counter.seven_segment0.ten_count_reg[3] ;
 wire \frequency_counter.seven_segment0.unit_count[0] ;
 wire \frequency_counter.seven_segment0.unit_count[1] ;
 wire \frequency_counter.seven_segment0.unit_count[2] ;
 wire \frequency_counter.seven_segment0.unit_count[3] ;
 wire \frequency_counter.seven_segment0.unit_count_reg[0] ;
 wire \frequency_counter.seven_segment0.unit_count_reg[1] ;
 wire \frequency_counter.seven_segment0.unit_count_reg[2] ;
 wire \frequency_counter.seven_segment0.unit_count_reg[3] ;
 wire \frequency_counter.update_period[0] ;
 wire \frequency_counter.update_period[10] ;
 wire \frequency_counter.update_period[11] ;
 wire \frequency_counter.update_period[1] ;
 wire \frequency_counter.update_period[2] ;
 wire \frequency_counter.update_period[3] ;
 wire \frequency_counter.update_period[4] ;
 wire \frequency_counter.update_period[5] ;
 wire \frequency_counter.update_period[6] ;
 wire \frequency_counter.update_period[7] ;
 wire \frequency_counter.update_period[8] ;
 wire \frequency_counter.update_period[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net107;

 sg13g2_inv_1 _354_ (.Y(_054_),
    .A(\frequency_counter.clk_counter[11] ));
 sg13g2_inv_1 _355_ (.Y(_055_),
    .A(\frequency_counter.clk_counter[10] ));
 sg13g2_inv_1 _356_ (.Y(_056_),
    .A(\frequency_counter.update_period[10] ));
 sg13g2_nand2b_1 _357_ (.Y(_057_),
    .B(\frequency_counter.clk_counter[8] ),
    .A_N(\frequency_counter.update_period[8] ));
 sg13g2_nand2_1 _358_ (.Y(_058_),
    .A(\frequency_counter.update_period[9] ),
    .B(_057_));
 sg13g2_nor2_1 _359_ (.A(\frequency_counter.update_period[9] ),
    .B(_057_),
    .Y(_059_));
 sg13g2_a221oi_1 _360_ (.B2(_058_),
    .C1(_059_),
    .B1(\frequency_counter.clk_counter[9] ),
    .A1(\frequency_counter.clk_counter[10] ),
    .Y(_060_),
    .A2(_056_));
 sg13g2_a221oi_1 _361_ (.B2(\frequency_counter.update_period[10] ),
    .C1(_060_),
    .B1(_055_),
    .A1(_054_),
    .Y(_061_),
    .A2(\frequency_counter.update_period[11] ));
 sg13g2_inv_1 _362_ (.Y(_062_),
    .A(\frequency_counter.clk_counter[1] ));
 sg13g2_nor2b_1 _363_ (.A(\frequency_counter.clk_counter[0] ),
    .B_N(\frequency_counter.update_period[0] ),
    .Y(_063_));
 sg13g2_a21oi_1 _364_ (.A1(_062_),
    .A2(_063_),
    .Y(_064_),
    .B1(\frequency_counter.update_period[1] ));
 sg13g2_nor2_1 _365_ (.A(_062_),
    .B(_063_),
    .Y(_065_));
 sg13g2_nand2b_1 _366_ (.Y(_066_),
    .B(\frequency_counter.update_period[2] ),
    .A_N(\frequency_counter.clk_counter[2] ));
 sg13g2_o21ai_1 _367_ (.B1(_066_),
    .Y(_067_),
    .A1(_064_),
    .A2(_065_));
 sg13g2_inv_1 _368_ (.Y(_068_),
    .A(\frequency_counter.update_period[3] ));
 sg13g2_inv_1 _369_ (.Y(_069_),
    .A(\frequency_counter.update_period[2] ));
 sg13g2_a22oi_1 _370_ (.Y(_070_),
    .B1(\frequency_counter.clk_counter[2] ),
    .B2(_069_),
    .A2(_068_),
    .A1(\frequency_counter.clk_counter[3] ));
 sg13g2_xor2_1 _371_ (.B(\frequency_counter.update_period[7] ),
    .A(\frequency_counter.clk_counter[7] ),
    .X(_071_));
 sg13g2_xor2_1 _372_ (.B(\frequency_counter.update_period[6] ),
    .A(\frequency_counter.clk_counter[6] ),
    .X(_072_));
 sg13g2_nor2b_1 _373_ (.A(\frequency_counter.clk_counter[5] ),
    .B_N(\frequency_counter.update_period[5] ),
    .Y(_073_));
 sg13g2_nor3_1 _374_ (.A(_071_),
    .B(_072_),
    .C(_073_),
    .Y(_074_));
 sg13g2_xor2_1 _375_ (.B(\frequency_counter.update_period[8] ),
    .A(\frequency_counter.clk_counter[8] ),
    .X(_075_));
 sg13g2_xor2_1 _376_ (.B(\frequency_counter.update_period[11] ),
    .A(\frequency_counter.clk_counter[11] ),
    .X(_076_));
 sg13g2_xor2_1 _377_ (.B(\frequency_counter.update_period[9] ),
    .A(\frequency_counter.clk_counter[9] ),
    .X(_077_));
 sg13g2_xor2_1 _378_ (.B(\frequency_counter.update_period[10] ),
    .A(\frequency_counter.clk_counter[10] ),
    .X(_078_));
 sg13g2_nor4_1 _379_ (.A(_075_),
    .B(_076_),
    .C(_077_),
    .D(_078_),
    .Y(_079_));
 sg13g2_inv_1 _380_ (.Y(_080_),
    .A(\frequency_counter.update_period[5] ));
 sg13g2_inv_1 _381_ (.Y(_081_),
    .A(\frequency_counter.clk_counter[3] ));
 sg13g2_a22oi_1 _382_ (.Y(_082_),
    .B1(_081_),
    .B2(\frequency_counter.update_period[3] ),
    .A2(_080_),
    .A1(\frequency_counter.clk_counter[5] ));
 sg13g2_xnor2_1 _383_ (.Y(_083_),
    .A(\frequency_counter.clk_counter[4] ),
    .B(\frequency_counter.update_period[4] ));
 sg13g2_nand4_1 _384_ (.B(_079_),
    .C(_082_),
    .A(_074_),
    .Y(_084_),
    .D(_083_));
 sg13g2_a21oi_1 _385_ (.A1(_067_),
    .A2(_070_),
    .Y(_085_),
    .B1(_084_));
 sg13g2_inv_1 _386_ (.Y(_086_),
    .A(\frequency_counter.update_period[11] ));
 sg13g2_a21oi_1 _387_ (.A1(\frequency_counter.clk_counter[11] ),
    .A2(_086_),
    .Y(_087_),
    .B1(_079_));
 sg13g2_inv_1 _388_ (.Y(_088_),
    .A(\frequency_counter.clk_counter[4] ));
 sg13g2_nand2b_1 _389_ (.Y(_089_),
    .B(\frequency_counter.clk_counter[5] ),
    .A_N(\frequency_counter.update_period[5] ));
 sg13g2_o21ai_1 _390_ (.B1(_089_),
    .Y(_090_),
    .A1(_088_),
    .A2(\frequency_counter.update_period[4] ));
 sg13g2_nand2b_1 _391_ (.Y(_091_),
    .B(\frequency_counter.clk_counter[6] ),
    .A_N(\frequency_counter.update_period[6] ));
 sg13g2_nand2_1 _392_ (.Y(_092_),
    .A(\frequency_counter.update_period[7] ),
    .B(_091_));
 sg13g2_nand2b_1 _393_ (.Y(_093_),
    .B(\frequency_counter.clk_counter[11] ),
    .A_N(\frequency_counter.update_period[11] ));
 sg13g2_o21ai_1 _394_ (.B1(_093_),
    .Y(_094_),
    .A1(\frequency_counter.update_period[7] ),
    .A2(_091_));
 sg13g2_a221oi_1 _395_ (.B2(\frequency_counter.clk_counter[7] ),
    .C1(_094_),
    .B1(_092_),
    .A1(_074_),
    .Y(_095_),
    .A2(_090_));
 sg13g2_nor2_1 _396_ (.A(_087_),
    .B(_095_),
    .Y(_096_));
 sg13g2_nor3_2 _397_ (.A(_061_),
    .B(_085_),
    .C(_096_),
    .Y(_097_));
 sg13g2_buf_8 _398_ (.A(net23),
    .X(_098_));
 sg13g2_nor2_2 _399_ (.A(_098_),
    .B(net24),
    .Y(_099_));
 sg13g2_nand3b_1 _400_ (.B(_097_),
    .C(_099_),
    .Y(_100_),
    .A_N(\frequency_counter.clk_counter[0] ));
 sg13g2_inv_2 _401_ (.Y(_101_),
    .A(_098_));
 sg13g2_inv_2 _402_ (.Y(_102_),
    .A(net24));
 sg13g2_nand2_2 _403_ (.Y(_103_),
    .A(_101_),
    .B(net51));
 sg13g2_nand2_1 _404_ (.Y(_104_),
    .A(\frequency_counter.clk_counter[0] ),
    .B(_103_));
 sg13g2_buf_2 _405_ (.A(rst_n),
    .X(_105_));
 sg13g2_inv_1 _406_ (.Y(_106_),
    .A(_105_));
 sg13g2_buf_1 _407_ (.A(_106_),
    .X(_107_));
 sg13g2_a21oi_1 _408_ (.A1(_100_),
    .A2(_104_),
    .Y(_003_),
    .B1(net44));
 sg13g2_o21ai_1 _409_ (.B1(_105_),
    .Y(_108_),
    .A1(_097_),
    .A2(_103_));
 sg13g2_buf_8 _410_ (.A(_108_),
    .X(_109_));
 sg13g2_nand3_1 _411_ (.B(\frequency_counter.clk_counter[3] ),
    .C(\frequency_counter.clk_counter[2] ),
    .A(\frequency_counter.clk_counter[4] ),
    .Y(_110_));
 sg13g2_nand2_1 _412_ (.Y(_111_),
    .A(\frequency_counter.clk_counter[6] ),
    .B(\frequency_counter.clk_counter[5] ));
 sg13g2_nand3_1 _413_ (.B(\frequency_counter.clk_counter[1] ),
    .C(\frequency_counter.clk_counter[0] ),
    .A(\frequency_counter.clk_counter[7] ),
    .Y(_112_));
 sg13g2_nor3_2 _414_ (.A(_110_),
    .B(_111_),
    .C(_112_),
    .Y(_113_));
 sg13g2_nand4_1 _415_ (.B(\frequency_counter.clk_counter[8] ),
    .C(_099_),
    .A(\frequency_counter.clk_counter[9] ),
    .Y(_114_),
    .D(_113_));
 sg13g2_xnor2_1 _416_ (.Y(_115_),
    .A(_055_),
    .B(_114_));
 sg13g2_nor2_1 _417_ (.A(net39),
    .B(_115_),
    .Y(_004_));
 sg13g2_or2_1 _418_ (.X(_116_),
    .B(_114_),
    .A(_055_));
 sg13g2_xnor2_1 _419_ (.Y(_117_),
    .A(_054_),
    .B(_116_));
 sg13g2_nor2_1 _420_ (.A(net39),
    .B(_117_),
    .Y(_005_));
 sg13g2_nand2_1 _421_ (.Y(_118_),
    .A(\frequency_counter.clk_counter[0] ),
    .B(_099_));
 sg13g2_xnor2_1 _422_ (.Y(_119_),
    .A(_062_),
    .B(_118_));
 sg13g2_nor2_1 _423_ (.A(net39),
    .B(_119_),
    .Y(_006_));
 sg13g2_nor2_1 _424_ (.A(_062_),
    .B(_118_),
    .Y(_120_));
 sg13g2_xnor2_1 _425_ (.Y(_121_),
    .A(\frequency_counter.clk_counter[2] ),
    .B(_120_));
 sg13g2_nor2_1 _426_ (.A(net39),
    .B(_121_),
    .Y(_007_));
 sg13g2_nand2_1 _427_ (.Y(_122_),
    .A(\frequency_counter.clk_counter[2] ),
    .B(_120_));
 sg13g2_xnor2_1 _428_ (.Y(_123_),
    .A(_081_),
    .B(_122_));
 sg13g2_nor2_1 _429_ (.A(net39),
    .B(_123_),
    .Y(_008_));
 sg13g2_nand3_1 _430_ (.B(\frequency_counter.clk_counter[2] ),
    .C(_120_),
    .A(\frequency_counter.clk_counter[3] ),
    .Y(_124_));
 sg13g2_xnor2_1 _431_ (.Y(_125_),
    .A(_088_),
    .B(_124_));
 sg13g2_nor2_1 _432_ (.A(net39),
    .B(_125_),
    .Y(_009_));
 sg13g2_nor3_2 _433_ (.A(_062_),
    .B(_110_),
    .C(_118_),
    .Y(_126_));
 sg13g2_xnor2_1 _434_ (.Y(_127_),
    .A(\frequency_counter.clk_counter[5] ),
    .B(_126_));
 sg13g2_nor2_1 _435_ (.A(net39),
    .B(_127_),
    .Y(_010_));
 sg13g2_nand2_1 _436_ (.Y(_128_),
    .A(\frequency_counter.clk_counter[5] ),
    .B(_126_));
 sg13g2_xor2_1 _437_ (.B(_128_),
    .A(\frequency_counter.clk_counter[6] ),
    .X(_129_));
 sg13g2_nor2_1 _438_ (.A(_109_),
    .B(_129_),
    .Y(_011_));
 sg13g2_nand2b_1 _439_ (.Y(_130_),
    .B(_126_),
    .A_N(_111_));
 sg13g2_xor2_1 _440_ (.B(_130_),
    .A(\frequency_counter.clk_counter[7] ),
    .X(_131_));
 sg13g2_nor2_1 _441_ (.A(_109_),
    .B(_131_),
    .Y(_012_));
 sg13g2_nand2_1 _442_ (.Y(_132_),
    .A(\frequency_counter.clk_counter[8] ),
    .B(_103_));
 sg13g2_nand2b_1 _443_ (.Y(_133_),
    .B(\frequency_counter.clk_counter[8] ),
    .A_N(_113_));
 sg13g2_nand3b_1 _444_ (.B(_099_),
    .C(_113_),
    .Y(_134_),
    .A_N(\frequency_counter.clk_counter[8] ));
 sg13g2_or3_1 _445_ (.A(_061_),
    .B(_085_),
    .C(_096_),
    .X(_135_));
 sg13g2_a21o_1 _446_ (.A2(_134_),
    .A1(_133_),
    .B1(_135_),
    .X(_136_));
 sg13g2_a21oi_1 _447_ (.A1(_132_),
    .A2(_136_),
    .Y(_013_),
    .B1(_107_));
 sg13g2_nand2_1 _448_ (.Y(_137_),
    .A(\frequency_counter.clk_counter[9] ),
    .B(_103_));
 sg13g2_nand2_1 _449_ (.Y(_138_),
    .A(\frequency_counter.clk_counter[8] ),
    .B(_113_));
 sg13g2_and2_1 _450_ (.A(\frequency_counter.clk_counter[9] ),
    .B(_138_),
    .X(_139_));
 sg13g2_nor3_1 _451_ (.A(\frequency_counter.clk_counter[9] ),
    .B(_103_),
    .C(_138_),
    .Y(_140_));
 sg13g2_o21ai_1 _452_ (.B1(_097_),
    .Y(_141_),
    .A1(_139_),
    .A2(_140_));
 sg13g2_a21oi_1 _453_ (.A1(_137_),
    .A2(_141_),
    .Y(_014_),
    .B1(net44));
 sg13g2_buf_1 _454_ (.A(_098_),
    .X(_142_));
 sg13g2_buf_1 _455_ (.A(\frequency_counter.edge_counter[0] ),
    .X(_143_));
 sg13g2_nand2b_2 _456_ (.Y(_144_),
    .B(\frequency_counter.edge_detect0.q1 ),
    .A_N(\frequency_counter.edge_detect0.q2 ));
 sg13g2_nor3_1 _457_ (.A(_098_),
    .B(net50),
    .C(_144_),
    .Y(_145_));
 sg13g2_a21o_1 _458_ (.A2(_144_),
    .A1(net50),
    .B1(_145_),
    .X(_146_));
 sg13g2_a22oi_1 _459_ (.Y(_147_),
    .B1(_146_),
    .B2(net51),
    .A2(net50),
    .A1(net43));
 sg13g2_nor2_1 _460_ (.A(net44),
    .B(_147_),
    .Y(_015_));
 sg13g2_buf_1 _461_ (.A(\frequency_counter.edge_counter[1] ),
    .X(_148_));
 sg13g2_o21ai_1 _462_ (.B1(net51),
    .Y(_149_),
    .A1(net49),
    .A2(net50));
 sg13g2_a21oi_1 _463_ (.A1(net51),
    .A2(_144_),
    .Y(_150_),
    .B1(_098_));
 sg13g2_buf_2 _464_ (.A(\frequency_counter.edge_counter[2] ),
    .X(_151_));
 sg13g2_nand2b_1 _465_ (.Y(_152_),
    .B(_002_),
    .A_N(net50));
 sg13g2_inv_1 _466_ (.Y(_153_),
    .A(\frequency_counter.edge_counter[1] ));
 sg13g2_a21oi_1 _467_ (.A1(_001_),
    .A2(_152_),
    .Y(_154_),
    .B1(_153_));
 sg13g2_o21ai_1 _468_ (.B1(\frequency_counter.edge_counter[3] ),
    .Y(_155_),
    .A1(net48),
    .A2(_154_));
 sg13g2_nor3_1 _469_ (.A(\frequency_counter.edge_counter[5] ),
    .B(\frequency_counter.edge_counter[6] ),
    .C(\frequency_counter.edge_counter[4] ),
    .Y(_156_));
 sg13g2_nor2_1 _470_ (.A(_101_),
    .B(net24),
    .Y(_157_));
 sg13g2_inv_1 _471_ (.Y(_158_),
    .A(_157_));
 sg13g2_a21oi_2 _472_ (.B1(_158_),
    .Y(_159_),
    .A2(_156_),
    .A1(_155_));
 sg13g2_nor2_1 _473_ (.A(_150_),
    .B(_159_),
    .Y(_160_));
 sg13g2_nor2_1 _474_ (.A(net51),
    .B(_143_),
    .Y(_161_));
 sg13g2_or3_1 _475_ (.A(net49),
    .B(net40),
    .C(_161_),
    .X(_162_));
 sg13g2_nor2_1 _476_ (.A(net50),
    .B(net41),
    .Y(_163_));
 sg13g2_o21ai_1 _477_ (.B1(net49),
    .Y(_164_),
    .A1(net40),
    .A2(_163_));
 sg13g2_a221oi_1 _478_ (.B2(_164_),
    .C1(_106_),
    .B1(_162_),
    .A1(_101_),
    .Y(_016_),
    .A2(_149_));
 sg13g2_buf_1 _479_ (.A(net24),
    .X(_165_));
 sg13g2_and2_1 _480_ (.A(_155_),
    .B(_156_),
    .X(_166_));
 sg13g2_nor3_1 _481_ (.A(_165_),
    .B(net49),
    .C(_166_),
    .Y(_167_));
 sg13g2_xnor2_1 _482_ (.Y(_168_),
    .A(_151_),
    .B(_167_));
 sg13g2_buf_1 _483_ (.A(_105_),
    .X(_169_));
 sg13g2_nand2_1 _484_ (.Y(_170_),
    .A(net49),
    .B(_143_));
 sg13g2_nor2_1 _485_ (.A(_144_),
    .B(_170_),
    .Y(_171_));
 sg13g2_xnor2_1 _486_ (.Y(_172_),
    .A(_151_),
    .B(_171_));
 sg13g2_o21ai_1 _487_ (.B1(_101_),
    .Y(_173_),
    .A1(net47),
    .A2(_172_));
 sg13g2_nand2_1 _488_ (.Y(_174_),
    .A(net46),
    .B(_173_));
 sg13g2_a21oi_1 _489_ (.A1(net43),
    .A2(_168_),
    .Y(_017_),
    .B1(_174_));
 sg13g2_and2_1 _490_ (.A(net49),
    .B(net50),
    .X(_175_));
 sg13g2_or2_1 _491_ (.X(_176_),
    .B(net49),
    .A(net48));
 sg13g2_nor2_2 _492_ (.A(_098_),
    .B(net51),
    .Y(_177_));
 sg13g2_a221oi_1 _493_ (.B2(net41),
    .C1(_177_),
    .B1(_176_),
    .A1(net48),
    .Y(_178_),
    .A2(_175_));
 sg13g2_o21ai_1 _494_ (.B1(\frequency_counter.edge_counter[3] ),
    .Y(_179_),
    .A1(net40),
    .A2(_178_));
 sg13g2_a21oi_1 _495_ (.A1(net47),
    .A2(_170_),
    .Y(_180_),
    .B1(_101_));
 sg13g2_a21o_1 _496_ (.A2(_175_),
    .A1(net51),
    .B1(_180_),
    .X(_181_));
 sg13g2_a22oi_1 _497_ (.Y(_182_),
    .B1(_181_),
    .B2(net48),
    .A2(net41),
    .A1(net49));
 sg13g2_or3_1 _498_ (.A(\frequency_counter.edge_counter[3] ),
    .B(net40),
    .C(_182_),
    .X(_183_));
 sg13g2_a21oi_1 _499_ (.A1(_179_),
    .A2(_183_),
    .Y(_018_),
    .B1(net44));
 sg13g2_o21ai_1 _500_ (.B1(\frequency_counter.edge_counter[3] ),
    .Y(_184_),
    .A1(net48),
    .A2(\frequency_counter.edge_counter[1] ));
 sg13g2_and4_1 _501_ (.A(\frequency_counter.edge_counter[3] ),
    .B(net48),
    .C(\frequency_counter.edge_counter[1] ),
    .D(net50),
    .X(_185_));
 sg13g2_a22oi_1 _502_ (.Y(_186_),
    .B1(_185_),
    .B2(net47),
    .A2(_184_),
    .A1(net41));
 sg13g2_o21ai_1 _503_ (.B1(_101_),
    .Y(_187_),
    .A1(net47),
    .A2(_185_));
 sg13g2_and2_1 _504_ (.A(_186_),
    .B(_187_),
    .X(_188_));
 sg13g2_o21ai_1 _505_ (.B1(\frequency_counter.edge_counter[4] ),
    .Y(_189_),
    .A1(net40),
    .A2(_188_));
 sg13g2_nor2b_1 _506_ (.A(\frequency_counter.edge_counter[4] ),
    .B_N(_184_),
    .Y(_190_));
 sg13g2_nor3_1 _507_ (.A(\frequency_counter.edge_counter[4] ),
    .B(_103_),
    .C(_144_),
    .Y(_191_));
 sg13g2_a22oi_1 _508_ (.Y(_192_),
    .B1(_185_),
    .B2(_191_),
    .A2(_190_),
    .A1(_159_));
 sg13g2_a21oi_1 _509_ (.A1(_189_),
    .A2(_192_),
    .Y(_019_),
    .B1(net44));
 sg13g2_and2_1 _510_ (.A(\frequency_counter.edge_counter[4] ),
    .B(_185_),
    .X(_193_));
 sg13g2_mux2_1 _511_ (.A0(_190_),
    .A1(_193_),
    .S(net47),
    .X(_194_));
 sg13g2_nor2_1 _512_ (.A(net47),
    .B(_193_),
    .Y(_195_));
 sg13g2_nor2_1 _513_ (.A(_098_),
    .B(_195_),
    .Y(_196_));
 sg13g2_a21oi_1 _514_ (.A1(net43),
    .A2(_194_),
    .Y(_197_),
    .B1(_196_));
 sg13g2_o21ai_1 _515_ (.B1(\frequency_counter.edge_counter[5] ),
    .Y(_198_),
    .A1(net40),
    .A2(_197_));
 sg13g2_a22oi_1 _516_ (.Y(_199_),
    .B1(_194_),
    .B2(net43),
    .A2(_193_),
    .A1(_099_));
 sg13g2_or3_1 _517_ (.A(\frequency_counter.edge_counter[5] ),
    .B(_160_),
    .C(_199_),
    .X(_200_));
 sg13g2_a21oi_1 _518_ (.A1(_198_),
    .A2(_200_),
    .Y(_020_),
    .B1(net44));
 sg13g2_nor2b_1 _519_ (.A(\frequency_counter.edge_counter[5] ),
    .B_N(_190_),
    .Y(_201_));
 sg13g2_xnor2_1 _520_ (.Y(_202_),
    .A(_002_),
    .B(_201_));
 sg13g2_nand2_1 _521_ (.Y(_203_),
    .A(net41),
    .B(_202_));
 sg13g2_nand2_1 _522_ (.Y(_204_),
    .A(\frequency_counter.edge_counter[5] ),
    .B(_193_));
 sg13g2_or4_1 _523_ (.A(\frequency_counter.edge_counter[6] ),
    .B(net41),
    .C(_177_),
    .D(_204_),
    .X(_205_));
 sg13g2_a21o_1 _524_ (.A2(_205_),
    .A1(_203_),
    .B1(net40),
    .X(_206_));
 sg13g2_inv_1 _525_ (.Y(_207_),
    .A(\frequency_counter.edge_counter[6] ));
 sg13g2_nor3_1 _526_ (.A(_207_),
    .B(net41),
    .C(_177_),
    .Y(_208_));
 sg13g2_a22oi_1 _527_ (.Y(_209_),
    .B1(_204_),
    .B2(_208_),
    .A2(net40),
    .A1(\frequency_counter.edge_counter[6] ));
 sg13g2_a21oi_1 _528_ (.A1(_206_),
    .A2(_209_),
    .Y(_021_),
    .B1(net44));
 sg13g2_and2_1 _529_ (.A(net46),
    .B(_000_),
    .X(_022_));
 sg13g2_buf_1 _530_ (.A(\frequency_counter.seven_segment0.load ),
    .X(_210_));
 sg13g2_nand2_1 _531_ (.Y(_211_),
    .A(\frequency_counter.seven_segment0.ten_count[0] ),
    .B(_210_));
 sg13g2_nand2b_1 _532_ (.Y(_212_),
    .B(\frequency_counter.seven_segment0.ten_count_reg[0] ),
    .A_N(net45));
 sg13g2_buf_1 _533_ (.A(_106_),
    .X(_213_));
 sg13g2_a21oi_1 _534_ (.A1(_211_),
    .A2(_212_),
    .Y(_023_),
    .B1(net42));
 sg13g2_nand2_1 _535_ (.Y(_214_),
    .A(\frequency_counter.seven_segment0.ten_count[1] ),
    .B(net45));
 sg13g2_nand2b_1 _536_ (.Y(_215_),
    .B(\frequency_counter.seven_segment0.ten_count_reg[1] ),
    .A_N(\frequency_counter.seven_segment0.load ));
 sg13g2_a21oi_1 _537_ (.A1(_214_),
    .A2(_215_),
    .Y(_024_),
    .B1(net42));
 sg13g2_nand2_1 _538_ (.Y(_216_),
    .A(\frequency_counter.seven_segment0.ten_count[2] ),
    .B(net45));
 sg13g2_nand2b_1 _539_ (.Y(_217_),
    .B(\frequency_counter.seven_segment0.ten_count_reg[2] ),
    .A_N(\frequency_counter.seven_segment0.load ));
 sg13g2_a21oi_1 _540_ (.A1(_216_),
    .A2(_217_),
    .Y(_025_),
    .B1(net42));
 sg13g2_nand2_1 _541_ (.Y(_218_),
    .A(\frequency_counter.seven_segment0.ten_count[3] ),
    .B(_210_));
 sg13g2_nand2b_1 _542_ (.Y(_219_),
    .B(\frequency_counter.seven_segment0.ten_count_reg[3] ),
    .A_N(\frequency_counter.seven_segment0.load ));
 sg13g2_a21oi_1 _543_ (.A1(_218_),
    .A2(_219_),
    .Y(_026_),
    .B1(net42));
 sg13g2_nand2_1 _544_ (.Y(_220_),
    .A(net45),
    .B(\frequency_counter.seven_segment0.unit_count[0] ));
 sg13g2_nand2b_1 _545_ (.Y(_221_),
    .B(\frequency_counter.seven_segment0.unit_count_reg[0] ),
    .A_N(\frequency_counter.seven_segment0.load ));
 sg13g2_a21oi_1 _546_ (.A1(_220_),
    .A2(_221_),
    .Y(_027_),
    .B1(net42));
 sg13g2_nand2_1 _547_ (.Y(_222_),
    .A(net45),
    .B(\frequency_counter.seven_segment0.unit_count[1] ));
 sg13g2_nand2b_1 _548_ (.Y(_223_),
    .B(\frequency_counter.seven_segment0.unit_count_reg[1] ),
    .A_N(\frequency_counter.seven_segment0.load ));
 sg13g2_a21oi_1 _549_ (.A1(_222_),
    .A2(_223_),
    .Y(_028_),
    .B1(net42));
 sg13g2_nand2_1 _550_ (.Y(_224_),
    .A(net45),
    .B(\frequency_counter.seven_segment0.unit_count[2] ));
 sg13g2_nand2b_1 _551_ (.Y(_225_),
    .B(\frequency_counter.seven_segment0.unit_count_reg[2] ),
    .A_N(\frequency_counter.seven_segment0.load ));
 sg13g2_a21oi_1 _552_ (.A1(_224_),
    .A2(_225_),
    .Y(_029_),
    .B1(net42));
 sg13g2_nand2_1 _553_ (.Y(_226_),
    .A(net45),
    .B(\frequency_counter.seven_segment0.unit_count[3] ));
 sg13g2_nand2b_1 _554_ (.Y(_227_),
    .B(\frequency_counter.seven_segment0.unit_count_reg[3] ),
    .A_N(\frequency_counter.seven_segment0.load ));
 sg13g2_a21oi_1 _555_ (.A1(_226_),
    .A2(_227_),
    .Y(_030_),
    .B1(net42));
 sg13g2_a21oi_1 _556_ (.A1(_135_),
    .A2(_099_),
    .Y(_228_),
    .B1(_159_));
 sg13g2_nor2_1 _557_ (.A(_107_),
    .B(_228_),
    .Y(_031_));
 sg13g2_and3_1 _558_ (.X(_032_),
    .A(net46),
    .B(_157_),
    .C(_166_));
 sg13g2_xnor2_1 _559_ (.Y(_229_),
    .A(\frequency_counter.seven_segment0.ten_count[0] ),
    .B(_159_));
 sg13g2_nor2_1 _560_ (.A(net39),
    .B(_229_),
    .Y(_033_));
 sg13g2_nand2_1 _561_ (.Y(_230_),
    .A(\frequency_counter.seven_segment0.ten_count[0] ),
    .B(_159_));
 sg13g2_xor2_1 _562_ (.B(_230_),
    .A(\frequency_counter.seven_segment0.ten_count[1] ),
    .X(_231_));
 sg13g2_nor2_1 _563_ (.A(_108_),
    .B(_231_),
    .Y(_034_));
 sg13g2_nand2b_1 _564_ (.Y(_232_),
    .B(\frequency_counter.seven_segment0.ten_count[2] ),
    .A_N(_159_));
 sg13g2_nand2_1 _565_ (.Y(_233_),
    .A(\frequency_counter.seven_segment0.ten_count[0] ),
    .B(\frequency_counter.seven_segment0.ten_count[1] ));
 sg13g2_or2_1 _566_ (.X(_234_),
    .B(_233_),
    .A(\frequency_counter.seven_segment0.ten_count[2] ));
 sg13g2_nand2_1 _567_ (.Y(_235_),
    .A(\frequency_counter.seven_segment0.ten_count[2] ),
    .B(_233_));
 sg13g2_o21ai_1 _568_ (.B1(_235_),
    .Y(_236_),
    .A1(_166_),
    .A2(_234_));
 sg13g2_nand3_1 _569_ (.B(net41),
    .C(_236_),
    .A(_105_),
    .Y(_237_));
 sg13g2_o21ai_1 _570_ (.B1(_237_),
    .Y(_035_),
    .A1(_108_),
    .A2(_232_));
 sg13g2_nand4_1 _571_ (.B(\frequency_counter.seven_segment0.ten_count[1] ),
    .C(\frequency_counter.seven_segment0.ten_count[2] ),
    .A(\frequency_counter.seven_segment0.ten_count[0] ),
    .Y(_238_),
    .D(_159_));
 sg13g2_xor2_1 _572_ (.B(_238_),
    .A(\frequency_counter.seven_segment0.ten_count[3] ),
    .X(_239_));
 sg13g2_nor2_1 _573_ (.A(_108_),
    .B(_239_),
    .Y(_036_));
 sg13g2_nand2_1 _574_ (.Y(_240_),
    .A(_102_),
    .B(_097_));
 sg13g2_nor3_1 _575_ (.A(net43),
    .B(net51),
    .C(_001_),
    .Y(_241_));
 sg13g2_nor2_1 _576_ (.A(net43),
    .B(_241_),
    .Y(_242_));
 sg13g2_o21ai_1 _577_ (.B1(_105_),
    .Y(_243_),
    .A1(\frequency_counter.seven_segment0.unit_count[0] ),
    .A2(_241_));
 sg13g2_a21oi_1 _578_ (.A1(_240_),
    .A2(_242_),
    .Y(_037_),
    .B1(_243_));
 sg13g2_a21oi_1 _579_ (.A1(net47),
    .A2(_148_),
    .Y(_244_),
    .B1(_142_));
 sg13g2_a21oi_1 _580_ (.A1(_148_),
    .A2(_177_),
    .Y(_245_),
    .B1(\frequency_counter.seven_segment0.unit_count[1] ));
 sg13g2_nand2b_1 _581_ (.Y(_246_),
    .B(_105_),
    .A_N(_245_));
 sg13g2_a21oi_1 _582_ (.A1(_240_),
    .A2(_244_),
    .Y(_038_),
    .B1(_246_));
 sg13g2_a21oi_1 _583_ (.A1(_165_),
    .A2(net48),
    .Y(_247_),
    .B1(net43));
 sg13g2_a21oi_1 _584_ (.A1(net48),
    .A2(_177_),
    .Y(_248_),
    .B1(\frequency_counter.seven_segment0.unit_count[2] ));
 sg13g2_nand2b_1 _585_ (.Y(_249_),
    .B(_105_),
    .A_N(_248_));
 sg13g2_a21oi_1 _586_ (.A1(_240_),
    .A2(_247_),
    .Y(_039_),
    .B1(_249_));
 sg13g2_a21oi_1 _587_ (.A1(net47),
    .A2(\frequency_counter.edge_counter[3] ),
    .Y(_250_),
    .B1(net43));
 sg13g2_a21oi_1 _588_ (.A1(\frequency_counter.edge_counter[3] ),
    .A2(_177_),
    .Y(_251_),
    .B1(\frequency_counter.seven_segment0.unit_count[3] ));
 sg13g2_nand2b_1 _589_ (.Y(_252_),
    .B(_105_),
    .A_N(_251_));
 sg13g2_a21oi_1 _590_ (.A1(_240_),
    .A2(_250_),
    .Y(_040_),
    .B1(_252_));
 sg13g2_a21oi_1 _591_ (.A1(_142_),
    .A2(net45),
    .Y(_253_),
    .B1(_177_));
 sg13g2_nor2_1 _592_ (.A(net44),
    .B(_253_),
    .Y(_041_));
 sg13g2_buf_1 _593_ (.A(net2),
    .X(_254_));
 sg13g2_nand2b_1 _594_ (.Y(_255_),
    .B(\frequency_counter.update_period[0] ),
    .A_N(net52));
 sg13g2_nand2_1 _595_ (.Y(_256_),
    .A(net7),
    .B(_254_));
 sg13g2_nand3_1 _596_ (.B(_255_),
    .C(_256_),
    .A(net46),
    .Y(_042_));
 sg13g2_nand2b_1 _597_ (.Y(_257_),
    .B(\frequency_counter.update_period[10] ),
    .A_N(net52));
 sg13g2_buf_2 _598_ (.A(net2),
    .X(_258_));
 sg13g2_nand2_1 _599_ (.Y(_259_),
    .A(net107),
    .B(net5));
 sg13g2_nand3_1 _600_ (.B(_257_),
    .C(_259_),
    .A(net46),
    .Y(_043_));
 sg13g2_nand2_1 _601_ (.Y(_260_),
    .A(_258_),
    .B(net6));
 sg13g2_nand2b_1 _602_ (.Y(_261_),
    .B(\frequency_counter.update_period[11] ),
    .A_N(net52));
 sg13g2_a21oi_1 _603_ (.A1(_260_),
    .A2(_261_),
    .Y(_044_),
    .B1(_213_));
 sg13g2_nand2b_1 _604_ (.Y(_262_),
    .B(\frequency_counter.update_period[1] ),
    .A_N(net52));
 sg13g2_nand2_1 _605_ (.Y(_263_),
    .A(net107),
    .B(net8));
 sg13g2_nand3_1 _606_ (.B(_262_),
    .C(_263_),
    .A(net46),
    .Y(_045_));
 sg13g2_nand2b_1 _607_ (.Y(_264_),
    .B(\frequency_counter.update_period[2] ),
    .A_N(net52));
 sg13g2_nand2_1 _608_ (.Y(_265_),
    .A(net107),
    .B(net9));
 sg13g2_nand3_1 _609_ (.B(_264_),
    .C(_265_),
    .A(net46),
    .Y(_046_));
 sg13g2_nand2b_1 _610_ (.Y(_266_),
    .B(\frequency_counter.update_period[3] ),
    .A_N(net52));
 sg13g2_nand2_1 _611_ (.Y(_267_),
    .A(net107),
    .B(net10));
 sg13g2_nand3_1 _612_ (.B(_266_),
    .C(_267_),
    .A(net46),
    .Y(_047_));
 sg13g2_nand2_1 _613_ (.Y(_268_),
    .A(_258_),
    .B(net11));
 sg13g2_nand2b_1 _614_ (.Y(_269_),
    .B(\frequency_counter.update_period[4] ),
    .A_N(net2));
 sg13g2_a21oi_1 _615_ (.A1(_268_),
    .A2(_269_),
    .Y(_048_),
    .B1(_213_));
 sg13g2_nand2b_1 _616_ (.Y(_270_),
    .B(\frequency_counter.update_period[5] ),
    .A_N(net52));
 sg13g2_nand2_1 _617_ (.Y(_271_),
    .A(net107),
    .B(net12));
 sg13g2_nand3_1 _618_ (.B(_270_),
    .C(_271_),
    .A(_169_),
    .Y(_049_));
 sg13g2_nand2_1 _619_ (.Y(_272_),
    .A(net107),
    .B(net13));
 sg13g2_nand2b_1 _620_ (.Y(_273_),
    .B(\frequency_counter.update_period[6] ),
    .A_N(net2));
 sg13g2_a21oi_1 _621_ (.A1(_272_),
    .A2(_273_),
    .Y(_050_),
    .B1(_106_));
 sg13g2_nand2b_1 _622_ (.Y(_274_),
    .B(\frequency_counter.update_period[7] ),
    .A_N(net52));
 sg13g2_nand2_1 _623_ (.Y(_275_),
    .A(net107),
    .B(net14));
 sg13g2_nand3_1 _624_ (.B(_274_),
    .C(_275_),
    .A(_169_),
    .Y(_051_));
 sg13g2_nand2_1 _625_ (.Y(_276_),
    .A(net107),
    .B(net3));
 sg13g2_nand2b_1 _626_ (.Y(_277_),
    .B(\frequency_counter.update_period[8] ),
    .A_N(net2));
 sg13g2_a21oi_1 _627_ (.A1(_276_),
    .A2(_277_),
    .Y(_052_),
    .B1(_106_));
 sg13g2_nand2_1 _628_ (.Y(_278_),
    .A(_254_),
    .B(net4));
 sg13g2_nand2b_1 _629_ (.Y(_279_),
    .B(\frequency_counter.update_period[9] ),
    .A_N(net2));
 sg13g2_a21oi_1 _630_ (.A1(_278_),
    .A2(_279_),
    .Y(_053_),
    .B1(_106_));
 sg13g2_mux2_2 _631_ (.A0(\frequency_counter.seven_segment0.unit_count_reg[2] ),
    .A1(\frequency_counter.seven_segment0.ten_count_reg[2] ),
    .S(\frequency_counter.digit ),
    .X(_280_));
 sg13g2_mux2_2 _632_ (.A0(\frequency_counter.seven_segment0.unit_count_reg[1] ),
    .A1(\frequency_counter.seven_segment0.ten_count_reg[1] ),
    .S(\frequency_counter.digit ),
    .X(_281_));
 sg13g2_or2_1 _633_ (.X(_282_),
    .B(_281_),
    .A(_280_));
 sg13g2_mux2_1 _634_ (.A0(\frequency_counter.seven_segment0.unit_count_reg[3] ),
    .A1(\frequency_counter.seven_segment0.ten_count_reg[3] ),
    .S(\frequency_counter.digit ),
    .X(_283_));
 sg13g2_buf_2 _635_ (.A(_283_),
    .X(_284_));
 sg13g2_and2_1 _636_ (.A(_282_),
    .B(_284_),
    .X(_285_));
 sg13g2_nor2b_1 _637_ (.A(\frequency_counter.digit ),
    .B_N(\frequency_counter.seven_segment0.unit_count_reg[0] ),
    .Y(_286_));
 sg13g2_a21o_1 _638_ (.A2(\frequency_counter.digit ),
    .A1(\frequency_counter.seven_segment0.ten_count_reg[0] ),
    .B1(_286_),
    .X(_287_));
 sg13g2_nand2b_1 _639_ (.Y(_288_),
    .B(_287_),
    .A_N(_284_));
 sg13g2_a21oi_2 _640_ (.B1(_286_),
    .Y(_289_),
    .A2(\frequency_counter.digit ),
    .A1(\frequency_counter.seven_segment0.ten_count_reg[0] ));
 sg13g2_nand2_1 _641_ (.Y(_290_),
    .A(_280_),
    .B(_289_));
 sg13g2_o21ai_1 _642_ (.B1(_290_),
    .Y(_291_),
    .A1(_282_),
    .A2(_288_));
 sg13g2_nor2_1 _643_ (.A(_285_),
    .B(_291_),
    .Y(net31));
 sg13g2_xnor2_1 _644_ (.Y(_292_),
    .A(_289_),
    .B(_281_));
 sg13g2_a21oi_1 _645_ (.A1(_280_),
    .A2(_292_),
    .Y(net32),
    .B1(_285_));
 sg13g2_nor2_1 _646_ (.A(_280_),
    .B(_287_),
    .Y(_293_));
 sg13g2_o21ai_1 _647_ (.B1(_282_),
    .Y(net33),
    .A1(_284_),
    .A2(_293_));
 sg13g2_nand2_1 _648_ (.Y(_294_),
    .A(_280_),
    .B(_287_));
 sg13g2_nor2_1 _649_ (.A(_284_),
    .B(_294_),
    .Y(_295_));
 sg13g2_nor2_1 _650_ (.A(_293_),
    .B(_295_),
    .Y(_296_));
 sg13g2_nand2b_1 _651_ (.Y(_297_),
    .B(_281_),
    .A_N(_284_));
 sg13g2_nand2b_1 _652_ (.Y(_298_),
    .B(_294_),
    .A_N(_297_));
 sg13g2_o21ai_1 _653_ (.B1(_298_),
    .Y(net34),
    .A1(_281_),
    .A2(_296_));
 sg13g2_a21oi_1 _654_ (.A1(_282_),
    .A2(_297_),
    .Y(net35),
    .B1(_287_));
 sg13g2_nor3_1 _655_ (.A(_280_),
    .B(_289_),
    .C(_284_),
    .Y(_299_));
 sg13g2_a221oi_1 _656_ (.B2(_280_),
    .C1(_299_),
    .B1(_284_),
    .A1(_290_),
    .Y(net36),
    .A2(_281_));
 sg13g2_nor2b_1 _657_ (.A(_294_),
    .B_N(_281_),
    .Y(_300_));
 sg13g2_nor2_1 _658_ (.A(_282_),
    .B(_284_),
    .Y(_301_));
 sg13g2_nor3_1 _659_ (.A(_285_),
    .B(_300_),
    .C(_301_),
    .Y(net37));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _661_ (.A(ui_in[1]),
    .X(net15));
 sg13g2_buf_1 _662_ (.A(ui_in[1]),
    .X(net16));
 sg13g2_buf_1 _663_ (.A(ui_in[1]),
    .X(net17));
 sg13g2_buf_1 _664_ (.A(ui_in[1]),
    .X(net18));
 sg13g2_buf_1 _665_ (.A(ui_in[1]),
    .X(net19));
 sg13g2_buf_1 _666_ (.A(ui_in[1]),
    .X(net20));
 sg13g2_buf_1 _667_ (.A(ui_in[1]),
    .X(net21));
 sg13g2_buf_1 _668_ (.A(ui_in[1]),
    .X(net22));
 sg13g2_buf_1 _669_ (.A(\frequency_counter.clk_counter[9] ),
    .X(net25));
 sg13g2_buf_1 _670_ (.A(\frequency_counter.clk_counter[10] ),
    .X(net26));
 sg13g2_buf_1 _671_ (.A(\frequency_counter.clk_counter[11] ),
    .X(net27));
 sg13g2_buf_1 _672_ (.A(\frequency_counter.edge_counter[4] ),
    .X(net28));
 sg13g2_buf_1 _673_ (.A(\frequency_counter.edge_counter[5] ),
    .X(net29));
 sg13g2_buf_1 _674_ (.A(\frequency_counter.edge_counter[6] ),
    .X(net30));
 sg13g2_buf_1 _675_ (.A(\frequency_counter.digit ),
    .X(net38));
 sg13g2_dfrbp_1 \frequency_counter.clk_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net53),
    .D(_003_),
    .Q_N(_350_),
    .Q(\frequency_counter.clk_counter[0] ));
 sg13g2_dfrbp_1 \frequency_counter.clk_counter[10]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net54),
    .D(_004_),
    .Q_N(_349_),
    .Q(\frequency_counter.clk_counter[10] ));
 sg13g2_dfrbp_1 \frequency_counter.clk_counter[11]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net55),
    .D(_005_),
    .Q_N(_348_),
    .Q(\frequency_counter.clk_counter[11] ));
 sg13g2_dfrbp_1 \frequency_counter.clk_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net56),
    .D(_006_),
    .Q_N(_347_),
    .Q(\frequency_counter.clk_counter[1] ));
 sg13g2_dfrbp_1 \frequency_counter.clk_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net57),
    .D(_007_),
    .Q_N(_346_),
    .Q(\frequency_counter.clk_counter[2] ));
 sg13g2_dfrbp_1 \frequency_counter.clk_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net58),
    .D(_008_),
    .Q_N(_345_),
    .Q(\frequency_counter.clk_counter[3] ));
 sg13g2_dfrbp_1 \frequency_counter.clk_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net59),
    .D(_009_),
    .Q_N(_344_),
    .Q(\frequency_counter.clk_counter[4] ));
 sg13g2_dfrbp_1 \frequency_counter.clk_counter[5]$_SDFFE_PN0P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net60),
    .D(_010_),
    .Q_N(_343_),
    .Q(\frequency_counter.clk_counter[5] ));
 sg13g2_dfrbp_1 \frequency_counter.clk_counter[6]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net61),
    .D(_011_),
    .Q_N(_342_),
    .Q(\frequency_counter.clk_counter[6] ));
 sg13g2_dfrbp_1 \frequency_counter.clk_counter[7]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net62),
    .D(_012_),
    .Q_N(_341_),
    .Q(\frequency_counter.clk_counter[7] ));
 sg13g2_dfrbp_1 \frequency_counter.clk_counter[8]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net63),
    .D(_013_),
    .Q_N(_340_),
    .Q(\frequency_counter.clk_counter[8] ));
 sg13g2_dfrbp_1 \frequency_counter.clk_counter[9]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net64),
    .D(_014_),
    .Q_N(_339_),
    .Q(\frequency_counter.clk_counter[9] ));
 sg13g2_dfrbp_1 \frequency_counter.edge_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net65),
    .D(_015_),
    .Q_N(_001_),
    .Q(\frequency_counter.edge_counter[0] ));
 sg13g2_dfrbp_1 \frequency_counter.edge_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net66),
    .D(_016_),
    .Q_N(_338_),
    .Q(\frequency_counter.edge_counter[1] ));
 sg13g2_dfrbp_1 \frequency_counter.edge_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net67),
    .D(_017_),
    .Q_N(_337_),
    .Q(\frequency_counter.edge_counter[2] ));
 sg13g2_dfrbp_1 \frequency_counter.edge_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net68),
    .D(_018_),
    .Q_N(_336_),
    .Q(\frequency_counter.edge_counter[3] ));
 sg13g2_dfrbp_1 \frequency_counter.edge_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net69),
    .D(_019_),
    .Q_N(_335_),
    .Q(\frequency_counter.edge_counter[4] ));
 sg13g2_dfrbp_1 \frequency_counter.edge_counter[5]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net70),
    .D(_020_),
    .Q_N(_334_),
    .Q(\frequency_counter.edge_counter[5] ));
 sg13g2_dfrbp_1 \frequency_counter.edge_counter[6]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net71),
    .D(_021_),
    .Q_N(_002_),
    .Q(\frequency_counter.edge_counter[6] ));
 sg13g2_dfrbp_1 \frequency_counter.edge_detect0.q0$_DFF_P_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net72),
    .D(net1),
    .Q_N(_351_),
    .Q(\frequency_counter.edge_detect0.q0 ));
 sg13g2_dfrbp_1 \frequency_counter.edge_detect0.q1$_DFF_P_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net73),
    .D(\frequency_counter.edge_detect0.q0 ),
    .Q_N(_352_),
    .Q(\frequency_counter.edge_detect0.q1 ));
 sg13g2_dfrbp_1 \frequency_counter.edge_detect0.q2$_DFF_P_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net74),
    .D(\frequency_counter.edge_detect0.q1 ),
    .Q_N(_333_),
    .Q(\frequency_counter.edge_detect0.q2 ));
 sg13g2_dfrbp_1 \frequency_counter.seven_segment0.digit$_SDFF_PN0_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net75),
    .D(_022_),
    .Q_N(_000_),
    .Q(\frequency_counter.digit ));
 sg13g2_dfrbp_1 \frequency_counter.seven_segment0.ten_count_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net76),
    .D(_023_),
    .Q_N(_332_),
    .Q(\frequency_counter.seven_segment0.ten_count_reg[0] ));
 sg13g2_dfrbp_1 \frequency_counter.seven_segment0.ten_count_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net77),
    .D(_024_),
    .Q_N(_331_),
    .Q(\frequency_counter.seven_segment0.ten_count_reg[1] ));
 sg13g2_dfrbp_1 \frequency_counter.seven_segment0.ten_count_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net78),
    .D(_025_),
    .Q_N(_330_),
    .Q(\frequency_counter.seven_segment0.ten_count_reg[2] ));
 sg13g2_dfrbp_1 \frequency_counter.seven_segment0.ten_count_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net79),
    .D(_026_),
    .Q_N(_329_),
    .Q(\frequency_counter.seven_segment0.ten_count_reg[3] ));
 sg13g2_dfrbp_1 \frequency_counter.seven_segment0.unit_count_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net80),
    .D(_027_),
    .Q_N(_328_),
    .Q(\frequency_counter.seven_segment0.unit_count_reg[0] ));
 sg13g2_dfrbp_1 \frequency_counter.seven_segment0.unit_count_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net81),
    .D(_028_),
    .Q_N(_327_),
    .Q(\frequency_counter.seven_segment0.unit_count_reg[1] ));
 sg13g2_dfrbp_1 \frequency_counter.seven_segment0.unit_count_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net82),
    .D(_029_),
    .Q_N(_326_),
    .Q(\frequency_counter.seven_segment0.unit_count_reg[2] ));
 sg13g2_dfrbp_1 \frequency_counter.seven_segment0.unit_count_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net83),
    .D(_030_),
    .Q_N(_325_),
    .Q(\frequency_counter.seven_segment0.unit_count_reg[3] ));
 sg13g2_dfrbp_1 \frequency_counter.state[0]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net84),
    .D(_031_),
    .Q_N(_324_),
    .Q(net23));
 sg13g2_dfrbp_1 \frequency_counter.state[1]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net85),
    .D(_032_),
    .Q_N(_323_),
    .Q(net24));
 sg13g2_dfrbp_1 \frequency_counter.ten_count[0]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net86),
    .D(_033_),
    .Q_N(_322_),
    .Q(\frequency_counter.seven_segment0.ten_count[0] ));
 sg13g2_dfrbp_1 \frequency_counter.ten_count[1]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net87),
    .D(_034_),
    .Q_N(_321_),
    .Q(\frequency_counter.seven_segment0.ten_count[1] ));
 sg13g2_dfrbp_1 \frequency_counter.ten_count[2]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net88),
    .D(_035_),
    .Q_N(_320_),
    .Q(\frequency_counter.seven_segment0.ten_count[2] ));
 sg13g2_dfrbp_1 \frequency_counter.ten_count[3]$_SDFFE_PN0P_  (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net89),
    .D(_036_),
    .Q_N(_319_),
    .Q(\frequency_counter.seven_segment0.ten_count[3] ));
 sg13g2_dfrbp_1 \frequency_counter.unit_count[0]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net90),
    .D(_037_),
    .Q_N(_318_),
    .Q(\frequency_counter.seven_segment0.unit_count[0] ));
 sg13g2_dfrbp_1 \frequency_counter.unit_count[1]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net91),
    .D(_038_),
    .Q_N(_317_),
    .Q(\frequency_counter.seven_segment0.unit_count[1] ));
 sg13g2_dfrbp_1 \frequency_counter.unit_count[2]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net92),
    .D(_039_),
    .Q_N(_316_),
    .Q(\frequency_counter.seven_segment0.unit_count[2] ));
 sg13g2_dfrbp_1 \frequency_counter.unit_count[3]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net93),
    .D(_040_),
    .Q_N(_315_),
    .Q(\frequency_counter.seven_segment0.unit_count[3] ));
 sg13g2_dfrbp_1 \frequency_counter.update_digits$_SDFFE_PN0N_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net94),
    .D(_041_),
    .Q_N(_314_),
    .Q(\frequency_counter.seven_segment0.load ));
 sg13g2_dfrbp_1 \frequency_counter.update_period[0]$_SDFFE_PN1P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net95),
    .D(_042_),
    .Q_N(_313_),
    .Q(\frequency_counter.update_period[0] ));
 sg13g2_dfrbp_1 \frequency_counter.update_period[10]$_SDFFE_PN1P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net96),
    .D(_043_),
    .Q_N(_312_),
    .Q(\frequency_counter.update_period[10] ));
 sg13g2_dfrbp_1 \frequency_counter.update_period[11]$_SDFFE_PN0P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net97),
    .D(_044_),
    .Q_N(_311_),
    .Q(\frequency_counter.update_period[11] ));
 sg13g2_dfrbp_1 \frequency_counter.update_period[1]$_SDFFE_PN1P_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net98),
    .D(_045_),
    .Q_N(_310_),
    .Q(\frequency_counter.update_period[1] ));
 sg13g2_dfrbp_1 \frequency_counter.update_period[2]$_SDFFE_PN1P_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net99),
    .D(_046_),
    .Q_N(_309_),
    .Q(\frequency_counter.update_period[2] ));
 sg13g2_dfrbp_1 \frequency_counter.update_period[3]$_SDFFE_PN1P_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net100),
    .D(_047_),
    .Q_N(_308_),
    .Q(\frequency_counter.update_period[3] ));
 sg13g2_dfrbp_1 \frequency_counter.update_period[4]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net101),
    .D(_048_),
    .Q_N(_307_),
    .Q(\frequency_counter.update_period[4] ));
 sg13g2_dfrbp_1 \frequency_counter.update_period[5]$_SDFFE_PN1P_  (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net102),
    .D(_049_),
    .Q_N(_306_),
    .Q(\frequency_counter.update_period[5] ));
 sg13g2_dfrbp_1 \frequency_counter.update_period[6]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net103),
    .D(_050_),
    .Q_N(_305_),
    .Q(\frequency_counter.update_period[6] ));
 sg13g2_dfrbp_1 \frequency_counter.update_period[7]$_SDFFE_PN1P_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net104),
    .D(_051_),
    .Q_N(_304_),
    .Q(\frequency_counter.update_period[7] ));
 sg13g2_dfrbp_1 \frequency_counter.update_period[8]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net105),
    .D(_052_),
    .Q_N(_303_),
    .Q(\frequency_counter.update_period[8] ));
 sg13g2_dfrbp_1 \frequency_counter.update_period[9]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net106),
    .D(_053_),
    .Q_N(_302_),
    .Q(\frequency_counter.update_period[9] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[0]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[6]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[7]),
    .X(net14));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[0]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_oe[1]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_oe[2]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_oe[3]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_oe[4]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_oe[5]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_oe[6]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_oe[7]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[0]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[1]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uio_out[2]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uio_out[3]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uio_out[4]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uio_out[5]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uio_out[6]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uio_out[7]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[0]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uo_out[1]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(uo_out[2]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(uo_out[3]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(uo_out[4]));
 sg13g2_buf_1 output36 (.A(net36),
    .X(uo_out[5]));
 sg13g2_buf_1 output37 (.A(net37),
    .X(uo_out[6]));
 sg13g2_buf_1 output38 (.A(net38),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout39 (.A(_109_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_160_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_157_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_213_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_142_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_107_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_210_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_169_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_165_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_151_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_148_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_143_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_102_),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(_254_),
    .X(net52));
 sg13g2_tiehi \frequency_counter.clk_counter[0]$_SDFFE_PN0P__53  (.L_HI(net53));
 sg13g2_tiehi \frequency_counter.clk_counter[10]$_SDFFE_PN0P__54  (.L_HI(net54));
 sg13g2_tiehi \frequency_counter.clk_counter[11]$_SDFFE_PN0P__55  (.L_HI(net55));
 sg13g2_tiehi \frequency_counter.clk_counter[1]$_SDFFE_PN0P__56  (.L_HI(net56));
 sg13g2_tiehi \frequency_counter.clk_counter[2]$_SDFFE_PN0P__57  (.L_HI(net57));
 sg13g2_tiehi \frequency_counter.clk_counter[3]$_SDFFE_PN0P__58  (.L_HI(net58));
 sg13g2_tiehi \frequency_counter.clk_counter[4]$_SDFFE_PN0P__59  (.L_HI(net59));
 sg13g2_tiehi \frequency_counter.clk_counter[5]$_SDFFE_PN0P__60  (.L_HI(net60));
 sg13g2_tiehi \frequency_counter.clk_counter[6]$_SDFFE_PN0P__61  (.L_HI(net61));
 sg13g2_tiehi \frequency_counter.clk_counter[7]$_SDFFE_PN0P__62  (.L_HI(net62));
 sg13g2_tiehi \frequency_counter.clk_counter[8]$_SDFFE_PN0P__63  (.L_HI(net63));
 sg13g2_tiehi \frequency_counter.clk_counter[9]$_SDFFE_PN0P__64  (.L_HI(net64));
 sg13g2_tiehi \frequency_counter.edge_counter[0]$_SDFFE_PN0P__65  (.L_HI(net65));
 sg13g2_tiehi \frequency_counter.edge_counter[1]$_SDFFE_PN0P__66  (.L_HI(net66));
 sg13g2_tiehi \frequency_counter.edge_counter[2]$_SDFFE_PN0P__67  (.L_HI(net67));
 sg13g2_tiehi \frequency_counter.edge_counter[3]$_SDFFE_PN0P__68  (.L_HI(net68));
 sg13g2_tiehi \frequency_counter.edge_counter[4]$_SDFFE_PN0P__69  (.L_HI(net69));
 sg13g2_tiehi \frequency_counter.edge_counter[5]$_SDFFE_PN0P__70  (.L_HI(net70));
 sg13g2_tiehi \frequency_counter.edge_counter[6]$_SDFFE_PN0P__71  (.L_HI(net71));
 sg13g2_tiehi \frequency_counter.edge_detect0.q0$_DFF_P__72  (.L_HI(net72));
 sg13g2_tiehi \frequency_counter.edge_detect0.q1$_DFF_P__73  (.L_HI(net73));
 sg13g2_tiehi \frequency_counter.edge_detect0.q2$_DFF_P__74  (.L_HI(net74));
 sg13g2_tiehi \frequency_counter.seven_segment0.digit$_SDFF_PN0__75  (.L_HI(net75));
 sg13g2_tiehi \frequency_counter.seven_segment0.ten_count_reg[0]$_SDFFE_PN0P__76  (.L_HI(net76));
 sg13g2_tiehi \frequency_counter.seven_segment0.ten_count_reg[1]$_SDFFE_PN0P__77  (.L_HI(net77));
 sg13g2_tiehi \frequency_counter.seven_segment0.ten_count_reg[2]$_SDFFE_PN0P__78  (.L_HI(net78));
 sg13g2_tiehi \frequency_counter.seven_segment0.ten_count_reg[3]$_SDFFE_PN0P__79  (.L_HI(net79));
 sg13g2_tiehi \frequency_counter.seven_segment0.unit_count_reg[0]$_SDFFE_PN0P__80  (.L_HI(net80));
 sg13g2_tiehi \frequency_counter.seven_segment0.unit_count_reg[1]$_SDFFE_PN0P__81  (.L_HI(net81));
 sg13g2_tiehi \frequency_counter.seven_segment0.unit_count_reg[2]$_SDFFE_PN0P__82  (.L_HI(net82));
 sg13g2_tiehi \frequency_counter.seven_segment0.unit_count_reg[3]$_SDFFE_PN0P__83  (.L_HI(net83));
 sg13g2_tiehi \frequency_counter.state[0]$_SDFFE_PN0P__84  (.L_HI(net84));
 sg13g2_tiehi \frequency_counter.state[1]$_SDFFE_PN0P__85  (.L_HI(net85));
 sg13g2_tiehi \frequency_counter.ten_count[0]$_SDFFE_PN0P__86  (.L_HI(net86));
 sg13g2_tiehi \frequency_counter.ten_count[1]$_SDFFE_PN0P__87  (.L_HI(net87));
 sg13g2_tiehi \frequency_counter.ten_count[2]$_SDFFE_PN0P__88  (.L_HI(net88));
 sg13g2_tiehi \frequency_counter.ten_count[3]$_SDFFE_PN0P__89  (.L_HI(net89));
 sg13g2_tiehi \frequency_counter.unit_count[0]$_SDFFE_PN0P__90  (.L_HI(net90));
 sg13g2_tiehi \frequency_counter.unit_count[1]$_SDFFE_PN0P__91  (.L_HI(net91));
 sg13g2_tiehi \frequency_counter.unit_count[2]$_SDFFE_PN0P__92  (.L_HI(net92));
 sg13g2_tiehi \frequency_counter.unit_count[3]$_SDFFE_PN0P__93  (.L_HI(net93));
 sg13g2_tiehi \frequency_counter.update_digits$_SDFFE_PN0N__94  (.L_HI(net94));
 sg13g2_tiehi \frequency_counter.update_period[0]$_SDFFE_PN1P__95  (.L_HI(net95));
 sg13g2_tiehi \frequency_counter.update_period[10]$_SDFFE_PN1P__96  (.L_HI(net96));
 sg13g2_tiehi \frequency_counter.update_period[11]$_SDFFE_PN0P__97  (.L_HI(net97));
 sg13g2_tiehi \frequency_counter.update_period[1]$_SDFFE_PN1P__98  (.L_HI(net98));
 sg13g2_tiehi \frequency_counter.update_period[2]$_SDFFE_PN1P__99  (.L_HI(net99));
 sg13g2_tiehi \frequency_counter.update_period[3]$_SDFFE_PN1P__100  (.L_HI(net100));
 sg13g2_tiehi \frequency_counter.update_period[4]$_SDFFE_PN0P__101  (.L_HI(net101));
 sg13g2_tiehi \frequency_counter.update_period[5]$_SDFFE_PN1P__102  (.L_HI(net102));
 sg13g2_tiehi \frequency_counter.update_period[6]$_SDFFE_PN0P__103  (.L_HI(net103));
 sg13g2_tiehi \frequency_counter.update_period[7]$_SDFFE_PN1P__104  (.L_HI(net104));
 sg13g2_tiehi \frequency_counter.update_period[8]$_SDFFE_PN0P__105  (.L_HI(net105));
 sg13g2_tiehi \frequency_counter.update_period[9]$_SDFFE_PN0P__106  (.L_HI(net106));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_7__leaf_clk));
 sg13g2_buf_1 fanout1 (.A(_258_),
    .X(net107));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_17_427 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_fill_2 FILLER_18_427 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_fill_2 FILLER_20_427 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_fill_2 FILLER_21_427 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_fill_2 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_125 ();
 sg13g2_decap_8 FILLER_24_132 ();
 sg13g2_decap_8 FILLER_24_139 ();
 sg13g2_decap_8 FILLER_24_146 ();
 sg13g2_fill_2 FILLER_24_153 ();
 sg13g2_decap_8 FILLER_24_185 ();
 sg13g2_decap_4 FILLER_24_192 ();
 sg13g2_fill_1 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_201 ();
 sg13g2_decap_8 FILLER_24_208 ();
 sg13g2_decap_8 FILLER_24_215 ();
 sg13g2_decap_8 FILLER_24_222 ();
 sg13g2_decap_8 FILLER_24_229 ();
 sg13g2_decap_8 FILLER_24_236 ();
 sg13g2_decap_8 FILLER_24_243 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_257 ();
 sg13g2_decap_8 FILLER_24_264 ();
 sg13g2_decap_8 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_decap_8 FILLER_24_299 ();
 sg13g2_decap_8 FILLER_24_306 ();
 sg13g2_decap_8 FILLER_24_313 ();
 sg13g2_decap_8 FILLER_24_320 ();
 sg13g2_decap_8 FILLER_24_327 ();
 sg13g2_decap_8 FILLER_24_334 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_8 FILLER_24_404 ();
 sg13g2_decap_8 FILLER_24_411 ();
 sg13g2_decap_8 FILLER_24_418 ();
 sg13g2_decap_4 FILLER_24_425 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_112 ();
 sg13g2_fill_1 FILLER_25_144 ();
 sg13g2_fill_1 FILLER_25_153 ();
 sg13g2_decap_4 FILLER_25_158 ();
 sg13g2_fill_2 FILLER_25_174 ();
 sg13g2_fill_1 FILLER_25_176 ();
 sg13g2_fill_1 FILLER_25_185 ();
 sg13g2_decap_8 FILLER_25_247 ();
 sg13g2_decap_8 FILLER_25_254 ();
 sg13g2_decap_8 FILLER_25_261 ();
 sg13g2_decap_8 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_275 ();
 sg13g2_decap_8 FILLER_25_282 ();
 sg13g2_decap_8 FILLER_25_289 ();
 sg13g2_decap_8 FILLER_25_296 ();
 sg13g2_decap_4 FILLER_25_303 ();
 sg13g2_fill_1 FILLER_25_307 ();
 sg13g2_decap_8 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_319 ();
 sg13g2_decap_8 FILLER_25_326 ();
 sg13g2_decap_4 FILLER_25_333 ();
 sg13g2_fill_1 FILLER_25_337 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_8 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_4 FILLER_25_424 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_4 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_116 ();
 sg13g2_decap_8 FILLER_26_143 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_fill_2 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_163 ();
 sg13g2_fill_2 FILLER_26_170 ();
 sg13g2_decap_4 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_180 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_256 ();
 sg13g2_decap_8 FILLER_26_263 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_284 ();
 sg13g2_decap_4 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_295 ();
 sg13g2_fill_1 FILLER_26_335 ();
 sg13g2_decap_4 FILLER_26_340 ();
 sg13g2_fill_2 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_fill_2 FILLER_26_427 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_4 FILLER_27_84 ();
 sg13g2_decap_4 FILLER_27_118 ();
 sg13g2_fill_2 FILLER_27_122 ();
 sg13g2_decap_8 FILLER_27_128 ();
 sg13g2_decap_4 FILLER_27_135 ();
 sg13g2_decap_4 FILLER_27_158 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_4 FILLER_27_190 ();
 sg13g2_fill_1 FILLER_27_194 ();
 sg13g2_fill_1 FILLER_27_199 ();
 sg13g2_fill_1 FILLER_27_205 ();
 sg13g2_fill_2 FILLER_27_216 ();
 sg13g2_fill_1 FILLER_27_218 ();
 sg13g2_fill_1 FILLER_27_224 ();
 sg13g2_fill_2 FILLER_27_230 ();
 sg13g2_fill_1 FILLER_27_232 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_fill_2 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_279 ();
 sg13g2_decap_8 FILLER_27_286 ();
 sg13g2_decap_4 FILLER_27_293 ();
 sg13g2_decap_4 FILLER_27_301 ();
 sg13g2_fill_1 FILLER_27_305 ();
 sg13g2_decap_8 FILLER_27_310 ();
 sg13g2_decap_8 FILLER_27_317 ();
 sg13g2_decap_8 FILLER_27_324 ();
 sg13g2_fill_2 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_27_412 ();
 sg13g2_decap_8 FILLER_27_419 ();
 sg13g2_decap_4 FILLER_27_426 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_51 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_fill_1 FILLER_28_70 ();
 sg13g2_decap_4 FILLER_28_102 ();
 sg13g2_fill_1 FILLER_28_106 ();
 sg13g2_decap_8 FILLER_28_111 ();
 sg13g2_fill_2 FILLER_28_118 ();
 sg13g2_decap_8 FILLER_28_129 ();
 sg13g2_decap_8 FILLER_28_136 ();
 sg13g2_decap_4 FILLER_28_143 ();
 sg13g2_fill_1 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_153 ();
 sg13g2_decap_4 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_162 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_200 ();
 sg13g2_decap_4 FILLER_28_232 ();
 sg13g2_fill_2 FILLER_28_236 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_decap_8 FILLER_28_254 ();
 sg13g2_fill_2 FILLER_28_261 ();
 sg13g2_fill_1 FILLER_28_263 ();
 sg13g2_fill_2 FILLER_28_294 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_fill_2 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_342 ();
 sg13g2_decap_4 FILLER_28_351 ();
 sg13g2_decap_8 FILLER_28_363 ();
 sg13g2_decap_4 FILLER_28_370 ();
 sg13g2_fill_1 FILLER_28_374 ();
 sg13g2_fill_2 FILLER_28_387 ();
 sg13g2_fill_1 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_4 FILLER_28_401 ();
 sg13g2_fill_2 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_28_411 ();
 sg13g2_decap_8 FILLER_28_418 ();
 sg13g2_decap_4 FILLER_28_425 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_fill_2 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_44 ();
 sg13g2_decap_4 FILLER_29_71 ();
 sg13g2_fill_2 FILLER_29_75 ();
 sg13g2_decap_8 FILLER_29_81 ();
 sg13g2_decap_4 FILLER_29_88 ();
 sg13g2_fill_1 FILLER_29_92 ();
 sg13g2_fill_2 FILLER_29_103 ();
 sg13g2_fill_2 FILLER_29_110 ();
 sg13g2_fill_1 FILLER_29_112 ();
 sg13g2_fill_1 FILLER_29_118 ();
 sg13g2_fill_2 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_153 ();
 sg13g2_fill_2 FILLER_29_164 ();
 sg13g2_fill_1 FILLER_29_166 ();
 sg13g2_decap_4 FILLER_29_218 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_decap_8 FILLER_29_234 ();
 sg13g2_fill_2 FILLER_29_241 ();
 sg13g2_fill_2 FILLER_29_269 ();
 sg13g2_fill_1 FILLER_29_271 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_fill_1 FILLER_29_329 ();
 sg13g2_decap_4 FILLER_29_361 ();
 sg13g2_fill_2 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_370 ();
 sg13g2_fill_2 FILLER_29_377 ();
 sg13g2_decap_4 FILLER_29_426 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_fill_2 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_30 ();
 sg13g2_decap_8 FILLER_30_78 ();
 sg13g2_decap_4 FILLER_30_85 ();
 sg13g2_fill_2 FILLER_30_89 ();
 sg13g2_decap_4 FILLER_30_100 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_decap_4 FILLER_30_110 ();
 sg13g2_fill_2 FILLER_30_114 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_4 FILLER_30_147 ();
 sg13g2_fill_2 FILLER_30_151 ();
 sg13g2_decap_8 FILLER_30_162 ();
 sg13g2_decap_8 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_188 ();
 sg13g2_decap_8 FILLER_30_195 ();
 sg13g2_fill_1 FILLER_30_202 ();
 sg13g2_decap_8 FILLER_30_223 ();
 sg13g2_decap_4 FILLER_30_230 ();
 sg13g2_decap_8 FILLER_30_250 ();
 sg13g2_decap_8 FILLER_30_257 ();
 sg13g2_fill_1 FILLER_30_271 ();
 sg13g2_fill_1 FILLER_30_281 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_4 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_305 ();
 sg13g2_decap_4 FILLER_30_313 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_decap_4 FILLER_30_349 ();
 sg13g2_fill_1 FILLER_30_368 ();
 sg13g2_fill_2 FILLER_30_377 ();
 sg13g2_fill_1 FILLER_30_379 ();
 sg13g2_fill_1 FILLER_30_399 ();
 sg13g2_decap_4 FILLER_30_426 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_65 ();
 sg13g2_fill_1 FILLER_31_72 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_decap_4 FILLER_31_105 ();
 sg13g2_decap_4 FILLER_31_114 ();
 sg13g2_fill_2 FILLER_31_146 ();
 sg13g2_fill_2 FILLER_31_178 ();
 sg13g2_fill_1 FILLER_31_180 ();
 sg13g2_decap_4 FILLER_31_212 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_fill_2 FILLER_31_222 ();
 sg13g2_fill_1 FILLER_31_224 ();
 sg13g2_fill_1 FILLER_31_233 ();
 sg13g2_fill_2 FILLER_31_249 ();
 sg13g2_fill_1 FILLER_31_255 ();
 sg13g2_fill_2 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_262 ();
 sg13g2_decap_8 FILLER_31_275 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_303 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_fill_1 FILLER_31_328 ();
 sg13g2_decap_8 FILLER_31_337 ();
 sg13g2_decap_8 FILLER_31_344 ();
 sg13g2_decap_8 FILLER_31_351 ();
 sg13g2_decap_4 FILLER_31_358 ();
 sg13g2_fill_1 FILLER_31_362 ();
 sg13g2_fill_2 FILLER_31_369 ();
 sg13g2_fill_1 FILLER_31_371 ();
 sg13g2_fill_2 FILLER_31_377 ();
 sg13g2_fill_1 FILLER_31_379 ();
 sg13g2_fill_2 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_1 FILLER_31_406 ();
 sg13g2_decap_8 FILLER_31_411 ();
 sg13g2_decap_8 FILLER_31_418 ();
 sg13g2_decap_4 FILLER_31_425 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_32 ();
 sg13g2_decap_4 FILLER_32_59 ();
 sg13g2_decap_4 FILLER_32_67 ();
 sg13g2_fill_2 FILLER_32_71 ();
 sg13g2_decap_4 FILLER_32_87 ();
 sg13g2_fill_1 FILLER_32_95 ();
 sg13g2_decap_8 FILLER_32_102 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_fill_2 FILLER_32_148 ();
 sg13g2_decap_8 FILLER_32_155 ();
 sg13g2_decap_8 FILLER_32_162 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_fill_2 FILLER_32_174 ();
 sg13g2_decap_8 FILLER_32_180 ();
 sg13g2_fill_2 FILLER_32_187 ();
 sg13g2_fill_1 FILLER_32_189 ();
 sg13g2_fill_1 FILLER_32_194 ();
 sg13g2_decap_8 FILLER_32_199 ();
 sg13g2_decap_8 FILLER_32_206 ();
 sg13g2_decap_8 FILLER_32_213 ();
 sg13g2_decap_4 FILLER_32_220 ();
 sg13g2_fill_2 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_4 FILLER_32_245 ();
 sg13g2_fill_2 FILLER_32_249 ();
 sg13g2_fill_2 FILLER_32_256 ();
 sg13g2_decap_8 FILLER_32_262 ();
 sg13g2_decap_8 FILLER_32_269 ();
 sg13g2_decap_4 FILLER_32_276 ();
 sg13g2_decap_8 FILLER_32_299 ();
 sg13g2_decap_8 FILLER_32_306 ();
 sg13g2_decap_8 FILLER_32_317 ();
 sg13g2_decap_8 FILLER_32_324 ();
 sg13g2_decap_8 FILLER_32_331 ();
 sg13g2_decap_4 FILLER_32_338 ();
 sg13g2_fill_2 FILLER_32_342 ();
 sg13g2_decap_8 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_decap_4 FILLER_32_362 ();
 sg13g2_fill_1 FILLER_32_380 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_404 ();
 sg13g2_decap_8 FILLER_32_411 ();
 sg13g2_decap_8 FILLER_32_418 ();
 sg13g2_decap_4 FILLER_32_425 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_4 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_43 ();
 sg13g2_decap_4 FILLER_33_50 ();
 sg13g2_fill_1 FILLER_33_54 ();
 sg13g2_decap_4 FILLER_33_63 ();
 sg13g2_fill_2 FILLER_33_93 ();
 sg13g2_fill_1 FILLER_33_95 ();
 sg13g2_fill_1 FILLER_33_100 ();
 sg13g2_decap_4 FILLER_33_113 ();
 sg13g2_fill_1 FILLER_33_117 ();
 sg13g2_decap_8 FILLER_33_146 ();
 sg13g2_decap_4 FILLER_33_153 ();
 sg13g2_fill_1 FILLER_33_157 ();
 sg13g2_fill_1 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_189 ();
 sg13g2_fill_1 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_201 ();
 sg13g2_fill_2 FILLER_33_208 ();
 sg13g2_fill_1 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_decap_4 FILLER_33_373 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_383 ();
 sg13g2_fill_2 FILLER_33_390 ();
 sg13g2_fill_1 FILLER_33_392 ();
 sg13g2_fill_2 FILLER_33_427 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_30 ();
 sg13g2_fill_1 FILLER_34_57 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_4 FILLER_34_79 ();
 sg13g2_fill_1 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_110 ();
 sg13g2_decap_4 FILLER_34_123 ();
 sg13g2_decap_8 FILLER_34_164 ();
 sg13g2_fill_2 FILLER_34_171 ();
 sg13g2_fill_2 FILLER_34_177 ();
 sg13g2_fill_1 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_222 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_fill_2 FILLER_34_273 ();
 sg13g2_fill_1 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_299 ();
 sg13g2_decap_8 FILLER_34_306 ();
 sg13g2_fill_2 FILLER_34_313 ();
 sg13g2_fill_2 FILLER_34_334 ();
 sg13g2_fill_1 FILLER_34_336 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_decap_4 FILLER_34_349 ();
 sg13g2_fill_2 FILLER_34_353 ();
 sg13g2_decap_4 FILLER_34_362 ();
 sg13g2_fill_1 FILLER_34_366 ();
 sg13g2_decap_4 FILLER_34_398 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_41 ();
 sg13g2_decap_8 FILLER_35_48 ();
 sg13g2_fill_1 FILLER_35_55 ();
 sg13g2_fill_2 FILLER_35_64 ();
 sg13g2_fill_2 FILLER_35_74 ();
 sg13g2_fill_1 FILLER_35_76 ();
 sg13g2_fill_1 FILLER_35_85 ();
 sg13g2_fill_2 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_93 ();
 sg13g2_fill_1 FILLER_35_107 ();
 sg13g2_fill_1 FILLER_35_113 ();
 sg13g2_fill_1 FILLER_35_123 ();
 sg13g2_fill_1 FILLER_35_130 ();
 sg13g2_fill_1 FILLER_35_136 ();
 sg13g2_fill_2 FILLER_35_142 ();
 sg13g2_decap_8 FILLER_35_149 ();
 sg13g2_fill_2 FILLER_35_156 ();
 sg13g2_fill_2 FILLER_35_187 ();
 sg13g2_decap_8 FILLER_35_193 ();
 sg13g2_decap_8 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_fill_2 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_236 ();
 sg13g2_fill_2 FILLER_35_278 ();
 sg13g2_decap_8 FILLER_35_285 ();
 sg13g2_fill_2 FILLER_35_292 ();
 sg13g2_decap_8 FILLER_35_302 ();
 sg13g2_decap_4 FILLER_35_309 ();
 sg13g2_fill_2 FILLER_35_313 ();
 sg13g2_fill_2 FILLER_35_346 ();
 sg13g2_fill_1 FILLER_35_378 ();
 sg13g2_fill_2 FILLER_35_384 ();
 sg13g2_decap_8 FILLER_35_390 ();
 sg13g2_fill_2 FILLER_35_397 ();
 sg13g2_fill_1 FILLER_35_399 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_28 ();
 sg13g2_fill_1 FILLER_36_32 ();
 sg13g2_fill_2 FILLER_36_75 ();
 sg13g2_fill_1 FILLER_36_77 ();
 sg13g2_decap_4 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_127 ();
 sg13g2_fill_1 FILLER_36_134 ();
 sg13g2_decap_8 FILLER_36_139 ();
 sg13g2_decap_8 FILLER_36_146 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_fill_2 FILLER_36_177 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_decap_4 FILLER_36_211 ();
 sg13g2_fill_2 FILLER_36_215 ();
 sg13g2_fill_2 FILLER_36_222 ();
 sg13g2_decap_8 FILLER_36_250 ();
 sg13g2_decap_4 FILLER_36_257 ();
 sg13g2_fill_1 FILLER_36_261 ();
 sg13g2_decap_4 FILLER_36_266 ();
 sg13g2_fill_2 FILLER_36_270 ();
 sg13g2_decap_4 FILLER_36_276 ();
 sg13g2_decap_8 FILLER_36_285 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_decap_8 FILLER_36_319 ();
 sg13g2_fill_1 FILLER_36_326 ();
 sg13g2_decap_8 FILLER_36_341 ();
 sg13g2_fill_2 FILLER_36_352 ();
 sg13g2_fill_1 FILLER_36_354 ();
 sg13g2_fill_2 FILLER_36_359 ();
 sg13g2_fill_1 FILLER_36_361 ();
 sg13g2_fill_2 FILLER_36_376 ();
 sg13g2_fill_1 FILLER_36_378 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_36_413 ();
 sg13g2_decap_8 FILLER_36_420 ();
 sg13g2_fill_2 FILLER_36_427 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_fill_2 FILLER_37_35 ();
 sg13g2_fill_1 FILLER_37_37 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_fill_1 FILLER_37_70 ();
 sg13g2_fill_1 FILLER_37_75 ();
 sg13g2_fill_1 FILLER_37_92 ();
 sg13g2_decap_8 FILLER_37_115 ();
 sg13g2_fill_2 FILLER_37_122 ();
 sg13g2_fill_1 FILLER_37_124 ();
 sg13g2_decap_8 FILLER_37_159 ();
 sg13g2_decap_8 FILLER_37_166 ();
 sg13g2_decap_4 FILLER_37_173 ();
 sg13g2_fill_2 FILLER_37_177 ();
 sg13g2_decap_4 FILLER_37_183 ();
 sg13g2_fill_1 FILLER_37_187 ();
 sg13g2_fill_1 FILLER_37_192 ();
 sg13g2_decap_8 FILLER_37_197 ();
 sg13g2_fill_1 FILLER_37_212 ();
 sg13g2_fill_1 FILLER_37_222 ();
 sg13g2_fill_1 FILLER_37_251 ();
 sg13g2_fill_2 FILLER_37_257 ();
 sg13g2_fill_2 FILLER_37_290 ();
 sg13g2_fill_1 FILLER_37_301 ();
 sg13g2_fill_2 FILLER_37_315 ();
 sg13g2_fill_1 FILLER_37_334 ();
 sg13g2_fill_1 FILLER_37_361 ();
 sg13g2_fill_1 FILLER_37_371 ();
 sg13g2_fill_2 FILLER_37_402 ();
 sg13g2_fill_1 FILLER_37_404 ();
 sg13g2_decap_8 FILLER_37_409 ();
 sg13g2_decap_8 FILLER_37_416 ();
 sg13g2_decap_8 FILLER_37_423 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_56 ();
 sg13g2_fill_2 FILLER_38_90 ();
 sg13g2_fill_2 FILLER_38_148 ();
 sg13g2_fill_2 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_160 ();
 sg13g2_fill_1 FILLER_38_167 ();
 sg13g2_fill_1 FILLER_38_198 ();
 sg13g2_fill_1 FILLER_38_203 ();
 sg13g2_fill_1 FILLER_38_208 ();
 sg13g2_fill_1 FILLER_38_213 ();
 sg13g2_fill_1 FILLER_38_218 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_fill_2 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_238 ();
 sg13g2_fill_1 FILLER_38_265 ();
 sg13g2_fill_2 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_313 ();
 sg13g2_fill_1 FILLER_38_318 ();
 sg13g2_fill_1 FILLER_38_323 ();
 sg13g2_fill_1 FILLER_38_387 ();
 sg13g2_fill_1 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_424 ();
 sg13g2_fill_2 FILLER_38_428 ();
endmodule
