module tt_um_z2a_rgb_mixer (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire clknet_0_clk;
 wire net53;
 wire \enc0[0] ;
 wire \enc0[1] ;
 wire \enc0[2] ;
 wire \enc0[3] ;
 wire \enc0[4] ;
 wire \enc0[5] ;
 wire \enc0[6] ;
 wire \enc0[7] ;
 wire \enc1[0] ;
 wire \enc1[1] ;
 wire \enc1[2] ;
 wire \enc1[3] ;
 wire \enc1[4] ;
 wire \enc1[5] ;
 wire \enc1[6] ;
 wire \enc1[7] ;
 wire \enc2[0] ;
 wire \enc2[1] ;
 wire \enc2[2] ;
 wire \enc2[3] ;
 wire \enc2[4] ;
 wire \enc2[5] ;
 wire \enc2[6] ;
 wire \enc2[7] ;
 wire \rgb_mixer.debounce0_a.button_hist[0] ;
 wire \rgb_mixer.debounce0_a.button_hist[1] ;
 wire \rgb_mixer.debounce0_a.button_hist[2] ;
 wire \rgb_mixer.debounce0_a.button_hist[3] ;
 wire \rgb_mixer.debounce0_a.button_hist[4] ;
 wire \rgb_mixer.debounce0_a.button_hist[5] ;
 wire \rgb_mixer.debounce0_a.button_hist[6] ;
 wire \rgb_mixer.debounce0_a.button_hist[7] ;
 wire \rgb_mixer.debounce0_a.debounced ;
 wire \rgb_mixer.debounce0_b.button_hist[0] ;
 wire \rgb_mixer.debounce0_b.button_hist[1] ;
 wire \rgb_mixer.debounce0_b.button_hist[2] ;
 wire \rgb_mixer.debounce0_b.button_hist[3] ;
 wire \rgb_mixer.debounce0_b.button_hist[4] ;
 wire \rgb_mixer.debounce0_b.button_hist[5] ;
 wire \rgb_mixer.debounce0_b.button_hist[6] ;
 wire \rgb_mixer.debounce0_b.button_hist[7] ;
 wire \rgb_mixer.debounce0_b.debounced ;
 wire \rgb_mixer.debounce1_a.button_hist[0] ;
 wire \rgb_mixer.debounce1_a.button_hist[1] ;
 wire \rgb_mixer.debounce1_a.button_hist[2] ;
 wire \rgb_mixer.debounce1_a.button_hist[3] ;
 wire \rgb_mixer.debounce1_a.button_hist[4] ;
 wire \rgb_mixer.debounce1_a.button_hist[5] ;
 wire \rgb_mixer.debounce1_a.button_hist[6] ;
 wire \rgb_mixer.debounce1_a.button_hist[7] ;
 wire \rgb_mixer.debounce1_a.debounced ;
 wire \rgb_mixer.debounce1_b.button_hist[0] ;
 wire \rgb_mixer.debounce1_b.button_hist[1] ;
 wire \rgb_mixer.debounce1_b.button_hist[2] ;
 wire \rgb_mixer.debounce1_b.button_hist[3] ;
 wire \rgb_mixer.debounce1_b.button_hist[4] ;
 wire \rgb_mixer.debounce1_b.button_hist[5] ;
 wire \rgb_mixer.debounce1_b.button_hist[6] ;
 wire \rgb_mixer.debounce1_b.button_hist[7] ;
 wire \rgb_mixer.debounce1_b.debounced ;
 wire \rgb_mixer.debounce2_a.button_hist[0] ;
 wire \rgb_mixer.debounce2_a.button_hist[1] ;
 wire \rgb_mixer.debounce2_a.button_hist[2] ;
 wire \rgb_mixer.debounce2_a.button_hist[3] ;
 wire \rgb_mixer.debounce2_a.button_hist[4] ;
 wire \rgb_mixer.debounce2_a.button_hist[5] ;
 wire \rgb_mixer.debounce2_a.button_hist[6] ;
 wire \rgb_mixer.debounce2_a.button_hist[7] ;
 wire \rgb_mixer.debounce2_a.debounced ;
 wire \rgb_mixer.debounce2_b.button_hist[0] ;
 wire \rgb_mixer.debounce2_b.button_hist[1] ;
 wire \rgb_mixer.debounce2_b.button_hist[2] ;
 wire \rgb_mixer.debounce2_b.button_hist[3] ;
 wire \rgb_mixer.debounce2_b.button_hist[4] ;
 wire \rgb_mixer.debounce2_b.button_hist[5] ;
 wire \rgb_mixer.debounce2_b.button_hist[6] ;
 wire \rgb_mixer.debounce2_b.button_hist[7] ;
 wire \rgb_mixer.debounce2_b.debounced ;
 wire \rgb_mixer.encoder0.old_a ;
 wire \rgb_mixer.encoder0.old_b ;
 wire \rgb_mixer.encoder1.old_a ;
 wire \rgb_mixer.encoder1.old_b ;
 wire \rgb_mixer.encoder2.old_a ;
 wire \rgb_mixer.encoder2.old_b ;
 wire \rgb_mixer.pwm0.count[0] ;
 wire \rgb_mixer.pwm0.count[1] ;
 wire \rgb_mixer.pwm0.count[2] ;
 wire \rgb_mixer.pwm0.count[3] ;
 wire \rgb_mixer.pwm0.count[4] ;
 wire \rgb_mixer.pwm0.count[5] ;
 wire \rgb_mixer.pwm0.count[6] ;
 wire \rgb_mixer.pwm0.count[7] ;
 wire \rgb_mixer.pwm0.out ;
 wire \rgb_mixer.pwm1.count[0] ;
 wire \rgb_mixer.pwm1.count[1] ;
 wire \rgb_mixer.pwm1.count[2] ;
 wire \rgb_mixer.pwm1.count[3] ;
 wire \rgb_mixer.pwm1.count[4] ;
 wire \rgb_mixer.pwm1.count[5] ;
 wire \rgb_mixer.pwm1.count[6] ;
 wire \rgb_mixer.pwm1.count[7] ;
 wire \rgb_mixer.pwm1.out ;
 wire \rgb_mixer.pwm2.count[0] ;
 wire \rgb_mixer.pwm2.count[1] ;
 wire \rgb_mixer.pwm2.count[2] ;
 wire \rgb_mixer.pwm2.count[3] ;
 wire \rgb_mixer.pwm2.count[4] ;
 wire \rgb_mixer.pwm2.count[5] ;
 wire \rgb_mixer.pwm2.count[6] ;
 wire \rgb_mixer.pwm2.count[7] ;
 wire \rgb_mixer.pwm2.out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_1 _0699_ (.A(rst_n),
    .X(_0123_));
 sg13g2_buf_1 _0700_ (.A(_0123_),
    .X(_0124_));
 sg13g2_buf_1 _0701_ (.A(net46),
    .X(_0125_));
 sg13g2_buf_1 _0702_ (.A(net29),
    .X(_0126_));
 sg13g2_and2_1 _0703_ (.A(net1),
    .B(net27),
    .X(_0012_));
 sg13g2_and2_1 _0704_ (.A(\rgb_mixer.debounce0_a.button_hist[0] ),
    .B(_0124_),
    .X(_0013_));
 sg13g2_and2_1 _0705_ (.A(\rgb_mixer.debounce0_a.button_hist[1] ),
    .B(net27),
    .X(_0014_));
 sg13g2_and2_1 _0706_ (.A(\rgb_mixer.debounce0_a.button_hist[2] ),
    .B(net27),
    .X(_0015_));
 sg13g2_and2_1 _0707_ (.A(\rgb_mixer.debounce0_a.button_hist[3] ),
    .B(net27),
    .X(_0016_));
 sg13g2_and2_1 _0708_ (.A(\rgb_mixer.debounce0_a.button_hist[4] ),
    .B(net27),
    .X(_0017_));
 sg13g2_and2_1 _0709_ (.A(\rgb_mixer.debounce0_a.button_hist[5] ),
    .B(net27),
    .X(_0018_));
 sg13g2_and2_1 _0710_ (.A(\rgb_mixer.debounce0_a.button_hist[6] ),
    .B(_0126_),
    .X(_0019_));
 sg13g2_nand4_1 _0711_ (.B(\rgb_mixer.debounce0_a.button_hist[2] ),
    .C(\rgb_mixer.debounce0_a.button_hist[4] ),
    .A(\rgb_mixer.debounce0_a.button_hist[3] ),
    .Y(_0127_),
    .D(\rgb_mixer.debounce0_a.button_hist[7] ));
 sg13g2_nand3_1 _0712_ (.B(\rgb_mixer.debounce0_a.button_hist[6] ),
    .C(_0013_),
    .A(\rgb_mixer.debounce0_a.button_hist[1] ),
    .Y(_0128_));
 sg13g2_nand2_1 _0713_ (.Y(_0129_),
    .A(\rgb_mixer.debounce0_a.debounced ),
    .B(_0124_));
 sg13g2_o21ai_1 _0714_ (.B1(_0129_),
    .Y(_0130_),
    .A1(_0127_),
    .A2(_0128_));
 sg13g2_nor4_1 _0715_ (.A(\rgb_mixer.debounce0_a.button_hist[2] ),
    .B(\rgb_mixer.debounce0_a.button_hist[4] ),
    .C(\rgb_mixer.debounce0_a.button_hist[7] ),
    .D(\rgb_mixer.debounce0_a.button_hist[6] ),
    .Y(_0131_));
 sg13g2_nor3_1 _0716_ (.A(\rgb_mixer.debounce0_a.button_hist[1] ),
    .B(\rgb_mixer.debounce0_a.button_hist[0] ),
    .C(\rgb_mixer.debounce0_a.button_hist[3] ),
    .Y(_0132_));
 sg13g2_a21oi_1 _0717_ (.A1(_0131_),
    .A2(_0132_),
    .Y(_0133_),
    .B1(_0129_));
 sg13g2_a21o_1 _0718_ (.A2(_0130_),
    .A1(\rgb_mixer.debounce0_a.button_hist[5] ),
    .B1(_0133_),
    .X(_0020_));
 sg13g2_buf_1 _0719_ (.A(net29),
    .X(_0134_));
 sg13g2_and2_1 _0720_ (.A(net26),
    .B(net2),
    .X(_0021_));
 sg13g2_and2_1 _0721_ (.A(\rgb_mixer.debounce0_b.button_hist[0] ),
    .B(_0126_),
    .X(_0022_));
 sg13g2_buf_1 _0722_ (.A(_0125_),
    .X(_0135_));
 sg13g2_and2_1 _0723_ (.A(\rgb_mixer.debounce0_b.button_hist[1] ),
    .B(net25),
    .X(_0023_));
 sg13g2_and2_1 _0724_ (.A(\rgb_mixer.debounce0_b.button_hist[2] ),
    .B(_0123_),
    .X(_0024_));
 sg13g2_and2_1 _0725_ (.A(\rgb_mixer.debounce0_b.button_hist[3] ),
    .B(net25),
    .X(_0025_));
 sg13g2_and2_1 _0726_ (.A(\rgb_mixer.debounce0_b.button_hist[4] ),
    .B(net25),
    .X(_0026_));
 sg13g2_and2_1 _0727_ (.A(\rgb_mixer.debounce0_b.button_hist[5] ),
    .B(_0135_),
    .X(_0027_));
 sg13g2_and2_1 _0728_ (.A(\rgb_mixer.debounce0_b.button_hist[6] ),
    .B(_0135_),
    .X(_0028_));
 sg13g2_nand4_1 _0729_ (.B(\rgb_mixer.debounce0_b.button_hist[3] ),
    .C(\rgb_mixer.debounce0_b.button_hist[4] ),
    .A(\rgb_mixer.debounce0_b.button_hist[0] ),
    .Y(_0136_),
    .D(\rgb_mixer.debounce0_b.button_hist[7] ));
 sg13g2_nand3_1 _0730_ (.B(\rgb_mixer.debounce0_b.button_hist[6] ),
    .C(_0024_),
    .A(\rgb_mixer.debounce0_b.button_hist[1] ),
    .Y(_0137_));
 sg13g2_buf_1 _0731_ (.A(\rgb_mixer.debounce0_b.debounced ),
    .X(_0138_));
 sg13g2_nand2_1 _0732_ (.Y(_0139_),
    .A(net45),
    .B(net46));
 sg13g2_o21ai_1 _0733_ (.B1(_0139_),
    .Y(_0140_),
    .A1(_0136_),
    .A2(_0137_));
 sg13g2_nor4_1 _0734_ (.A(\rgb_mixer.debounce0_b.button_hist[2] ),
    .B(\rgb_mixer.debounce0_b.button_hist[4] ),
    .C(\rgb_mixer.debounce0_b.button_hist[7] ),
    .D(\rgb_mixer.debounce0_b.button_hist[6] ),
    .Y(_0141_));
 sg13g2_nor3_1 _0735_ (.A(\rgb_mixer.debounce0_b.button_hist[1] ),
    .B(\rgb_mixer.debounce0_b.button_hist[0] ),
    .C(\rgb_mixer.debounce0_b.button_hist[3] ),
    .Y(_0142_));
 sg13g2_a21oi_1 _0736_ (.A1(_0141_),
    .A2(_0142_),
    .Y(_0143_),
    .B1(_0139_));
 sg13g2_a21o_1 _0737_ (.A2(_0140_),
    .A1(\rgb_mixer.debounce0_b.button_hist[5] ),
    .B1(_0143_),
    .X(_0029_));
 sg13g2_and2_1 _0738_ (.A(net26),
    .B(net3),
    .X(_0030_));
 sg13g2_and2_1 _0739_ (.A(\rgb_mixer.debounce1_a.button_hist[0] ),
    .B(net25),
    .X(_0031_));
 sg13g2_and2_1 _0740_ (.A(\rgb_mixer.debounce1_a.button_hist[1] ),
    .B(net25),
    .X(_0032_));
 sg13g2_and2_1 _0741_ (.A(\rgb_mixer.debounce1_a.button_hist[2] ),
    .B(net25),
    .X(_0033_));
 sg13g2_and2_1 _0742_ (.A(\rgb_mixer.debounce1_a.button_hist[3] ),
    .B(net25),
    .X(_0034_));
 sg13g2_and2_1 _0743_ (.A(\rgb_mixer.debounce1_a.button_hist[4] ),
    .B(net25),
    .X(_0035_));
 sg13g2_buf_1 _0744_ (.A(_0125_),
    .X(_0144_));
 sg13g2_and2_1 _0745_ (.A(\rgb_mixer.debounce1_a.button_hist[5] ),
    .B(net24),
    .X(_0036_));
 sg13g2_and2_1 _0746_ (.A(\rgb_mixer.debounce1_a.button_hist[6] ),
    .B(_0123_),
    .X(_0037_));
 sg13g2_nand4_1 _0747_ (.B(\rgb_mixer.debounce1_a.button_hist[3] ),
    .C(\rgb_mixer.debounce1_a.button_hist[2] ),
    .A(\rgb_mixer.debounce1_a.button_hist[0] ),
    .Y(_0145_),
    .D(\rgb_mixer.debounce1_a.button_hist[4] ));
 sg13g2_nand3_1 _0748_ (.B(\rgb_mixer.debounce1_a.button_hist[7] ),
    .C(_0037_),
    .A(\rgb_mixer.debounce1_a.button_hist[1] ),
    .Y(_0146_));
 sg13g2_nand2_1 _0749_ (.Y(_0147_),
    .A(\rgb_mixer.debounce1_a.debounced ),
    .B(net46));
 sg13g2_o21ai_1 _0750_ (.B1(_0147_),
    .Y(_0148_),
    .A1(_0145_),
    .A2(_0146_));
 sg13g2_nor4_1 _0751_ (.A(\rgb_mixer.debounce1_a.button_hist[2] ),
    .B(\rgb_mixer.debounce1_a.button_hist[4] ),
    .C(\rgb_mixer.debounce1_a.button_hist[7] ),
    .D(\rgb_mixer.debounce1_a.button_hist[6] ),
    .Y(_0149_));
 sg13g2_nor3_1 _0752_ (.A(\rgb_mixer.debounce1_a.button_hist[1] ),
    .B(\rgb_mixer.debounce1_a.button_hist[0] ),
    .C(\rgb_mixer.debounce1_a.button_hist[3] ),
    .Y(_0150_));
 sg13g2_a21oi_1 _0753_ (.A1(_0149_),
    .A2(_0150_),
    .Y(_0151_),
    .B1(_0147_));
 sg13g2_a21o_1 _0754_ (.A2(_0148_),
    .A1(\rgb_mixer.debounce1_a.button_hist[5] ),
    .B1(_0151_),
    .X(_0038_));
 sg13g2_and2_1 _0755_ (.A(net26),
    .B(net4),
    .X(_0039_));
 sg13g2_and2_1 _0756_ (.A(\rgb_mixer.debounce1_b.button_hist[0] ),
    .B(net24),
    .X(_0040_));
 sg13g2_and2_1 _0757_ (.A(\rgb_mixer.debounce1_b.button_hist[1] ),
    .B(_0123_),
    .X(_0041_));
 sg13g2_and2_1 _0758_ (.A(\rgb_mixer.debounce1_b.button_hist[2] ),
    .B(net24),
    .X(_0042_));
 sg13g2_and2_1 _0759_ (.A(\rgb_mixer.debounce1_b.button_hist[3] ),
    .B(net24),
    .X(_0043_));
 sg13g2_and2_1 _0760_ (.A(\rgb_mixer.debounce1_b.button_hist[4] ),
    .B(net24),
    .X(_0044_));
 sg13g2_and2_1 _0761_ (.A(\rgb_mixer.debounce1_b.button_hist[5] ),
    .B(_0144_),
    .X(_0045_));
 sg13g2_and2_1 _0762_ (.A(\rgb_mixer.debounce1_b.button_hist[6] ),
    .B(_0144_),
    .X(_0046_));
 sg13g2_nand4_1 _0763_ (.B(\rgb_mixer.debounce1_b.button_hist[2] ),
    .C(\rgb_mixer.debounce1_b.button_hist[4] ),
    .A(\rgb_mixer.debounce1_b.button_hist[3] ),
    .Y(_0152_),
    .D(\rgb_mixer.debounce1_b.button_hist[7] ));
 sg13g2_nand3_1 _0764_ (.B(\rgb_mixer.debounce1_b.button_hist[6] ),
    .C(_0041_),
    .A(\rgb_mixer.debounce1_b.button_hist[0] ),
    .Y(_0153_));
 sg13g2_nand2_1 _0765_ (.Y(_0154_),
    .A(\rgb_mixer.debounce1_b.debounced ),
    .B(net46));
 sg13g2_o21ai_1 _0766_ (.B1(_0154_),
    .Y(_0155_),
    .A1(_0152_),
    .A2(_0153_));
 sg13g2_nor4_1 _0767_ (.A(\rgb_mixer.debounce1_b.button_hist[2] ),
    .B(\rgb_mixer.debounce1_b.button_hist[4] ),
    .C(\rgb_mixer.debounce1_b.button_hist[7] ),
    .D(\rgb_mixer.debounce1_b.button_hist[6] ),
    .Y(_0156_));
 sg13g2_nor3_1 _0768_ (.A(\rgb_mixer.debounce1_b.button_hist[1] ),
    .B(\rgb_mixer.debounce1_b.button_hist[0] ),
    .C(\rgb_mixer.debounce1_b.button_hist[3] ),
    .Y(_0157_));
 sg13g2_a21oi_1 _0769_ (.A1(_0156_),
    .A2(_0157_),
    .Y(_0158_),
    .B1(_0154_));
 sg13g2_a21o_1 _0770_ (.A2(_0155_),
    .A1(\rgb_mixer.debounce1_b.button_hist[5] ),
    .B1(_0158_),
    .X(_0047_));
 sg13g2_and2_1 _0771_ (.A(_0134_),
    .B(net5),
    .X(_0048_));
 sg13g2_and2_1 _0772_ (.A(\rgb_mixer.debounce2_a.button_hist[0] ),
    .B(net24),
    .X(_0049_));
 sg13g2_and2_1 _0773_ (.A(\rgb_mixer.debounce2_a.button_hist[1] ),
    .B(_0123_),
    .X(_0050_));
 sg13g2_and2_1 _0774_ (.A(\rgb_mixer.debounce2_a.button_hist[2] ),
    .B(net24),
    .X(_0051_));
 sg13g2_and2_1 _0775_ (.A(\rgb_mixer.debounce2_a.button_hist[3] ),
    .B(net24),
    .X(_0052_));
 sg13g2_buf_1 _0776_ (.A(net46),
    .X(_0159_));
 sg13g2_and2_1 _0777_ (.A(\rgb_mixer.debounce2_a.button_hist[4] ),
    .B(_0159_),
    .X(_0053_));
 sg13g2_and2_1 _0778_ (.A(\rgb_mixer.debounce2_a.button_hist[5] ),
    .B(net28),
    .X(_0054_));
 sg13g2_and2_1 _0779_ (.A(\rgb_mixer.debounce2_a.button_hist[6] ),
    .B(net28),
    .X(_0055_));
 sg13g2_nand4_1 _0780_ (.B(\rgb_mixer.debounce2_a.button_hist[2] ),
    .C(\rgb_mixer.debounce2_a.button_hist[4] ),
    .A(\rgb_mixer.debounce2_a.button_hist[3] ),
    .Y(_0160_),
    .D(\rgb_mixer.debounce2_a.button_hist[7] ));
 sg13g2_nand3_1 _0781_ (.B(\rgb_mixer.debounce2_a.button_hist[6] ),
    .C(_0050_),
    .A(\rgb_mixer.debounce2_a.button_hist[0] ),
    .Y(_0161_));
 sg13g2_buf_2 _0782_ (.A(\rgb_mixer.debounce2_a.debounced ),
    .X(_0162_));
 sg13g2_nand2_1 _0783_ (.Y(_0163_),
    .A(_0162_),
    .B(net46));
 sg13g2_o21ai_1 _0784_ (.B1(_0163_),
    .Y(_0164_),
    .A1(_0160_),
    .A2(_0161_));
 sg13g2_nor4_1 _0785_ (.A(\rgb_mixer.debounce2_a.button_hist[2] ),
    .B(\rgb_mixer.debounce2_a.button_hist[4] ),
    .C(\rgb_mixer.debounce2_a.button_hist[7] ),
    .D(\rgb_mixer.debounce2_a.button_hist[6] ),
    .Y(_0165_));
 sg13g2_nor3_1 _0786_ (.A(\rgb_mixer.debounce2_a.button_hist[1] ),
    .B(\rgb_mixer.debounce2_a.button_hist[0] ),
    .C(\rgb_mixer.debounce2_a.button_hist[3] ),
    .Y(_0166_));
 sg13g2_a21oi_1 _0787_ (.A1(_0165_),
    .A2(_0166_),
    .Y(_0167_),
    .B1(_0163_));
 sg13g2_a21o_1 _0788_ (.A2(_0164_),
    .A1(\rgb_mixer.debounce2_a.button_hist[5] ),
    .B1(_0167_),
    .X(_0056_));
 sg13g2_and2_1 _0789_ (.A(_0134_),
    .B(net6),
    .X(_0057_));
 sg13g2_and2_1 _0790_ (.A(\rgb_mixer.debounce2_b.button_hist[0] ),
    .B(net28),
    .X(_0058_));
 sg13g2_and2_1 _0791_ (.A(\rgb_mixer.debounce2_b.button_hist[1] ),
    .B(_0123_),
    .X(_0059_));
 sg13g2_and2_1 _0792_ (.A(\rgb_mixer.debounce2_b.button_hist[2] ),
    .B(net28),
    .X(_0060_));
 sg13g2_and2_1 _0793_ (.A(\rgb_mixer.debounce2_b.button_hist[3] ),
    .B(net28),
    .X(_0061_));
 sg13g2_and2_1 _0794_ (.A(\rgb_mixer.debounce2_b.button_hist[4] ),
    .B(net28),
    .X(_0062_));
 sg13g2_and2_1 _0795_ (.A(\rgb_mixer.debounce2_b.button_hist[5] ),
    .B(net28),
    .X(_0063_));
 sg13g2_and2_1 _0796_ (.A(\rgb_mixer.debounce2_b.button_hist[6] ),
    .B(_0159_),
    .X(_0064_));
 sg13g2_nand4_1 _0797_ (.B(\rgb_mixer.debounce2_b.button_hist[3] ),
    .C(\rgb_mixer.debounce2_b.button_hist[5] ),
    .A(\rgb_mixer.debounce2_b.button_hist[2] ),
    .Y(_0168_),
    .D(\rgb_mixer.debounce2_b.button_hist[7] ));
 sg13g2_nand3_1 _0798_ (.B(\rgb_mixer.debounce2_b.button_hist[6] ),
    .C(_0059_),
    .A(\rgb_mixer.debounce2_b.button_hist[0] ),
    .Y(_0169_));
 sg13g2_buf_1 _0799_ (.A(\rgb_mixer.debounce2_b.debounced ),
    .X(_0170_));
 sg13g2_nand2_1 _0800_ (.Y(_0171_),
    .A(_0170_),
    .B(net46));
 sg13g2_o21ai_1 _0801_ (.B1(_0171_),
    .Y(_0172_),
    .A1(_0168_),
    .A2(_0169_));
 sg13g2_nor4_1 _0802_ (.A(\rgb_mixer.debounce2_b.button_hist[3] ),
    .B(\rgb_mixer.debounce2_b.button_hist[5] ),
    .C(\rgb_mixer.debounce2_b.button_hist[7] ),
    .D(\rgb_mixer.debounce2_b.button_hist[6] ),
    .Y(_0173_));
 sg13g2_nor3_1 _0803_ (.A(\rgb_mixer.debounce2_b.button_hist[0] ),
    .B(\rgb_mixer.debounce2_b.button_hist[1] ),
    .C(\rgb_mixer.debounce2_b.button_hist[2] ),
    .Y(_0174_));
 sg13g2_a21oi_1 _0804_ (.A1(_0173_),
    .A2(_0174_),
    .Y(_0175_),
    .B1(_0171_));
 sg13g2_a21o_1 _0805_ (.A2(_0172_),
    .A1(\rgb_mixer.debounce2_b.button_hist[4] ),
    .B1(_0175_),
    .X(_0065_));
 sg13g2_inv_1 _0806_ (.Y(_0066_),
    .A(_0129_));
 sg13g2_inv_1 _0807_ (.Y(_0067_),
    .A(_0139_));
 sg13g2_buf_1 _0808_ (.A(\rgb_mixer.encoder0.old_b ),
    .X(_0176_));
 sg13g2_buf_2 _0809_ (.A(\rgb_mixer.encoder0.old_a ),
    .X(_0177_));
 sg13g2_and2_1 _0810_ (.A(net43),
    .B(_0177_),
    .X(_0178_));
 sg13g2_nor2_1 _0811_ (.A(net43),
    .B(_0177_),
    .Y(_0179_));
 sg13g2_or2_1 _0812_ (.X(_0180_),
    .B(_0179_),
    .A(_0178_));
 sg13g2_nor2b_1 _0813_ (.A(net45),
    .B_N(\rgb_mixer.debounce0_a.debounced ),
    .Y(_0181_));
 sg13g2_nand2b_2 _0814_ (.Y(_0182_),
    .B(net45),
    .A_N(\rgb_mixer.debounce0_a.debounced ));
 sg13g2_nand2b_1 _0815_ (.Y(_0183_),
    .B(_0182_),
    .A_N(_0181_));
 sg13g2_and2_1 _0816_ (.A(_0180_),
    .B(_0183_),
    .X(_0184_));
 sg13g2_buf_1 _0817_ (.A(_0184_),
    .X(_0185_));
 sg13g2_nand2_1 _0818_ (.Y(_0186_),
    .A(_0009_),
    .B(_0185_));
 sg13g2_buf_2 _0819_ (.A(\enc0[0] ),
    .X(_0187_));
 sg13g2_nand2_2 _0820_ (.Y(_0188_),
    .A(_0180_),
    .B(_0183_));
 sg13g2_nand2_1 _0821_ (.Y(_0189_),
    .A(_0187_),
    .B(_0188_));
 sg13g2_inv_2 _0822_ (.Y(_0190_),
    .A(net46));
 sg13g2_buf_1 _0823_ (.A(_0190_),
    .X(_0191_));
 sg13g2_a21oi_1 _0824_ (.A1(_0186_),
    .A2(_0189_),
    .Y(_0068_),
    .B1(_0191_));
 sg13g2_buf_1 _0825_ (.A(_0190_),
    .X(_0192_));
 sg13g2_buf_1 _0826_ (.A(\enc0[1] ),
    .X(_0193_));
 sg13g2_nor2b_1 _0827_ (.A(\rgb_mixer.debounce0_a.debounced ),
    .B_N(net45),
    .Y(_0194_));
 sg13g2_a22oi_1 _0828_ (.Y(_0195_),
    .B1(_0194_),
    .B2(_0179_),
    .A2(_0181_),
    .A1(_0178_));
 sg13g2_buf_2 _0829_ (.A(_0195_),
    .X(_0196_));
 sg13g2_xnor2_1 _0830_ (.Y(_0197_),
    .A(_0009_),
    .B(_0196_));
 sg13g2_nor2_1 _0831_ (.A(_0188_),
    .B(_0197_),
    .Y(_0198_));
 sg13g2_xnor2_1 _0832_ (.Y(_0199_),
    .A(net42),
    .B(_0198_));
 sg13g2_nor2_1 _0833_ (.A(_0192_),
    .B(_0199_),
    .Y(_0069_));
 sg13g2_buf_1 _0834_ (.A(_0190_),
    .X(_0200_));
 sg13g2_buf_1 _0835_ (.A(\enc0[2] ),
    .X(_0201_));
 sg13g2_nor2_1 _0836_ (.A(net41),
    .B(_0185_),
    .Y(_0202_));
 sg13g2_nand3_1 _0837_ (.B(_0187_),
    .C(_0196_),
    .A(net42),
    .Y(_0203_));
 sg13g2_nor2_1 _0838_ (.A(net42),
    .B(_0187_),
    .Y(_0204_));
 sg13g2_nand2b_1 _0839_ (.Y(_0205_),
    .B(_0204_),
    .A_N(_0196_));
 sg13g2_nand2_1 _0840_ (.Y(_0206_),
    .A(_0203_),
    .B(_0205_));
 sg13g2_xnor2_1 _0841_ (.Y(_0207_),
    .A(_0004_),
    .B(_0206_));
 sg13g2_nor2_1 _0842_ (.A(_0188_),
    .B(_0207_),
    .Y(_0208_));
 sg13g2_nor3_1 _0843_ (.A(net21),
    .B(_0202_),
    .C(_0208_),
    .Y(_0070_));
 sg13g2_inv_1 _0844_ (.Y(_0209_),
    .A(_0004_));
 sg13g2_nor2_1 _0845_ (.A(_0209_),
    .B(_0196_),
    .Y(_0210_));
 sg13g2_nand2b_1 _0846_ (.Y(_0211_),
    .B(_0004_),
    .A_N(_0196_));
 sg13g2_o21ai_1 _0847_ (.B1(_0203_),
    .Y(_0212_),
    .A1(net42),
    .A2(_0211_));
 sg13g2_a22oi_1 _0848_ (.Y(_0213_),
    .B1(_0212_),
    .B2(net41),
    .A2(_0210_),
    .A1(_0204_));
 sg13g2_xnor2_1 _0849_ (.Y(_0214_),
    .A(_0005_),
    .B(_0213_));
 sg13g2_buf_1 _0850_ (.A(\enc0[3] ),
    .X(_0215_));
 sg13g2_o21ai_1 _0851_ (.B1(net28),
    .Y(_0216_),
    .A1(net40),
    .A2(_0185_));
 sg13g2_a21oi_1 _0852_ (.A1(_0185_),
    .A2(_0214_),
    .Y(_0071_),
    .B1(_0216_));
 sg13g2_buf_1 _0853_ (.A(\enc0[4] ),
    .X(_0217_));
 sg13g2_nor2_1 _0854_ (.A(net39),
    .B(net21),
    .Y(_0218_));
 sg13g2_and2_1 _0855_ (.A(net39),
    .B(net29),
    .X(_0219_));
 sg13g2_nand3_1 _0856_ (.B(net40),
    .C(net41),
    .A(net45),
    .Y(_0220_));
 sg13g2_nand3b_1 _0857_ (.B(\rgb_mixer.debounce0_a.debounced ),
    .C(_0177_),
    .Y(_0221_),
    .A_N(\rgb_mixer.debounce0_b.debounced ));
 sg13g2_or3_1 _0858_ (.A(net40),
    .B(net41),
    .C(_0221_),
    .X(_0222_));
 sg13g2_nand3_1 _0859_ (.B(_0220_),
    .C(_0222_),
    .A(net43),
    .Y(_0223_));
 sg13g2_nor4_1 _0860_ (.A(_0177_),
    .B(net40),
    .C(_0201_),
    .D(_0182_),
    .Y(_0224_));
 sg13g2_nand2_1 _0861_ (.Y(_0225_),
    .A(net40),
    .B(\enc0[2] ));
 sg13g2_nor2_1 _0862_ (.A(net45),
    .B(_0225_),
    .Y(_0226_));
 sg13g2_or3_1 _0863_ (.A(net43),
    .B(_0224_),
    .C(_0226_),
    .X(_0227_));
 sg13g2_o21ai_1 _0864_ (.B1(_0221_),
    .Y(_0228_),
    .A1(_0177_),
    .A2(_0182_));
 sg13g2_nor2_1 _0865_ (.A(_0225_),
    .B(_0228_),
    .Y(_0229_));
 sg13g2_a21oi_1 _0866_ (.A1(_0223_),
    .A2(_0227_),
    .Y(_0230_),
    .B1(_0229_));
 sg13g2_or2_1 _0867_ (.X(_0231_),
    .B(_0230_),
    .A(_0204_));
 sg13g2_and2_1 _0868_ (.A(_0005_),
    .B(_0210_),
    .X(_0232_));
 sg13g2_nor3_1 _0869_ (.A(_0188_),
    .B(_0203_),
    .C(_0230_),
    .Y(_0233_));
 sg13g2_a21oi_1 _0870_ (.A1(_0231_),
    .A2(_0232_),
    .Y(_0234_),
    .B1(_0233_));
 sg13g2_mux2_1 _0871_ (.A0(_0218_),
    .A1(_0219_),
    .S(_0234_),
    .X(_0072_));
 sg13g2_buf_1 _0872_ (.A(\enc0[5] ),
    .X(_0235_));
 sg13g2_nand2_1 _0873_ (.Y(_0236_),
    .A(net39),
    .B(net40));
 sg13g2_or2_1 _0874_ (.X(_0237_),
    .B(_0236_),
    .A(_0228_));
 sg13g2_or2_1 _0875_ (.X(_0238_),
    .B(net40),
    .A(net39));
 sg13g2_nand3_1 _0876_ (.B(net39),
    .C(_0215_),
    .A(net45),
    .Y(_0239_));
 sg13g2_o21ai_1 _0877_ (.B1(_0239_),
    .Y(_0240_),
    .A1(_0221_),
    .A2(_0238_));
 sg13g2_nor2_1 _0878_ (.A(net43),
    .B(_0238_),
    .Y(_0241_));
 sg13g2_nor2_1 _0879_ (.A(_0177_),
    .B(_0182_),
    .Y(_0242_));
 sg13g2_nor3_1 _0880_ (.A(net45),
    .B(net43),
    .C(_0236_),
    .Y(_0243_));
 sg13g2_a221oi_1 _0881_ (.B2(_0242_),
    .C1(_0243_),
    .B1(_0241_),
    .A1(net43),
    .Y(_0244_),
    .A2(_0240_));
 sg13g2_nand2_1 _0882_ (.Y(_0245_),
    .A(_0237_),
    .B(_0244_));
 sg13g2_nand2b_1 _0883_ (.Y(_0246_),
    .B(_0187_),
    .A_N(net41));
 sg13g2_nand3b_1 _0884_ (.B(_0004_),
    .C(_0246_),
    .Y(_0247_),
    .A_N(net42));
 sg13g2_nor2b_1 _0885_ (.A(_0217_),
    .B_N(_0005_),
    .Y(_0248_));
 sg13g2_nand2b_1 _0886_ (.Y(_0249_),
    .B(_0248_),
    .A_N(_0196_));
 sg13g2_a21o_1 _0887_ (.A2(_0247_),
    .A1(_0245_),
    .B1(_0249_),
    .X(_0250_));
 sg13g2_nand4_1 _0888_ (.B(net42),
    .C(_0187_),
    .A(_0201_),
    .Y(_0251_),
    .D(_0196_));
 sg13g2_a21oi_1 _0889_ (.A1(_0237_),
    .A2(_0244_),
    .Y(_0252_),
    .B1(_0251_));
 sg13g2_nand2_1 _0890_ (.Y(_0253_),
    .A(_0185_),
    .B(_0252_));
 sg13g2_nand3_1 _0891_ (.B(_0250_),
    .C(_0253_),
    .A(net38),
    .Y(_0254_));
 sg13g2_a21o_1 _0892_ (.A2(_0253_),
    .A1(_0250_),
    .B1(net38),
    .X(_0255_));
 sg13g2_a21oi_1 _0893_ (.A1(_0254_),
    .A2(_0255_),
    .Y(_0073_),
    .B1(_0191_));
 sg13g2_buf_1 _0894_ (.A(\enc0[6] ),
    .X(_0256_));
 sg13g2_nor2_1 _0895_ (.A(net37),
    .B(net21),
    .Y(_0257_));
 sg13g2_and2_1 _0896_ (.A(net37),
    .B(net29),
    .X(_0258_));
 sg13g2_nor3_1 _0897_ (.A(net38),
    .B(_0209_),
    .C(_0249_),
    .Y(_0259_));
 sg13g2_and2_1 _0898_ (.A(net38),
    .B(_0217_),
    .X(_0260_));
 sg13g2_a22oi_1 _0899_ (.Y(_0261_),
    .B1(_0260_),
    .B2(_0233_),
    .A2(_0259_),
    .A1(_0231_));
 sg13g2_mux2_1 _0900_ (.A0(_0257_),
    .A1(_0258_),
    .S(_0261_),
    .X(_0074_));
 sg13g2_and2_1 _0901_ (.A(_0237_),
    .B(_0244_),
    .X(_0262_));
 sg13g2_or2_1 _0902_ (.X(_0263_),
    .B(net38),
    .A(net37));
 sg13g2_buf_1 _0903_ (.A(_0263_),
    .X(_0264_));
 sg13g2_nor2_1 _0904_ (.A(_0249_),
    .B(_0264_),
    .Y(_0265_));
 sg13g2_inv_1 _0905_ (.Y(_0266_),
    .A(_0176_));
 sg13g2_nand3_1 _0906_ (.B(net37),
    .C(_0235_),
    .A(_0138_),
    .Y(_0267_));
 sg13g2_o21ai_1 _0907_ (.B1(_0267_),
    .Y(_0268_),
    .A1(_0221_),
    .A2(_0264_));
 sg13g2_nor2_1 _0908_ (.A(_0266_),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_nand2_1 _0909_ (.Y(_0270_),
    .A(_0256_),
    .B(_0235_));
 sg13g2_nor2_1 _0910_ (.A(_0138_),
    .B(_0270_),
    .Y(_0271_));
 sg13g2_nor3_1 _0911_ (.A(_0177_),
    .B(_0182_),
    .C(_0264_),
    .Y(_0272_));
 sg13g2_nor3_1 _0912_ (.A(net43),
    .B(_0271_),
    .C(_0272_),
    .Y(_0273_));
 sg13g2_or2_1 _0913_ (.X(_0274_),
    .B(_0270_),
    .A(_0228_));
 sg13g2_o21ai_1 _0914_ (.B1(_0274_),
    .Y(_0275_),
    .A1(_0269_),
    .A2(_0273_));
 sg13g2_nor3_1 _0915_ (.A(_0249_),
    .B(_0247_),
    .C(_0264_),
    .Y(_0276_));
 sg13g2_a221oi_1 _0916_ (.B2(_0252_),
    .C1(_0276_),
    .B1(_0275_),
    .A1(_0262_),
    .Y(_0277_),
    .A2(_0265_));
 sg13g2_o21ai_1 _0917_ (.B1(\enc0[7] ),
    .Y(_0278_),
    .A1(_0188_),
    .A2(_0277_));
 sg13g2_or3_1 _0918_ (.A(\enc0[7] ),
    .B(_0188_),
    .C(_0277_),
    .X(_0279_));
 sg13g2_a21oi_1 _0919_ (.A1(_0278_),
    .A2(_0279_),
    .Y(_0075_),
    .B1(_0200_));
 sg13g2_inv_1 _0920_ (.Y(_0076_),
    .A(_0147_));
 sg13g2_inv_1 _0921_ (.Y(_0077_),
    .A(_0154_));
 sg13g2_buf_2 _0922_ (.A(\enc1[0] ),
    .X(_0280_));
 sg13g2_buf_2 _0923_ (.A(\rgb_mixer.encoder1.old_b ),
    .X(_0281_));
 sg13g2_nand2_1 _0924_ (.Y(_0282_),
    .A(_0281_),
    .B(\rgb_mixer.encoder1.old_a ));
 sg13g2_nor2_2 _0925_ (.A(_0281_),
    .B(\rgb_mixer.encoder1.old_a ),
    .Y(_0283_));
 sg13g2_inv_1 _0926_ (.Y(_0284_),
    .A(_0283_));
 sg13g2_nor2b_2 _0927_ (.A(\rgb_mixer.debounce1_b.debounced ),
    .B_N(\rgb_mixer.debounce1_a.debounced ),
    .Y(_0285_));
 sg13g2_nor2b_2 _0928_ (.A(\rgb_mixer.debounce1_a.debounced ),
    .B_N(\rgb_mixer.debounce1_b.debounced ),
    .Y(_0286_));
 sg13g2_nor2_1 _0929_ (.A(_0285_),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_a21oi_2 _0930_ (.B1(_0287_),
    .Y(_0288_),
    .A2(_0284_),
    .A1(_0282_));
 sg13g2_mux2_1 _0931_ (.A0(_0280_),
    .A1(_0010_),
    .S(_0288_),
    .X(_0289_));
 sg13g2_and2_1 _0932_ (.A(net26),
    .B(_0289_),
    .X(_0078_));
 sg13g2_buf_2 _0933_ (.A(\enc1[1] ),
    .X(_0290_));
 sg13g2_inv_1 _0934_ (.Y(_0291_),
    .A(_0290_));
 sg13g2_and2_1 _0935_ (.A(_0281_),
    .B(\rgb_mixer.encoder1.old_a ),
    .X(_0292_));
 sg13g2_a22oi_1 _0936_ (.Y(_0293_),
    .B1(_0286_),
    .B2(_0283_),
    .A2(_0285_),
    .A1(_0292_));
 sg13g2_buf_1 _0937_ (.A(_0293_),
    .X(_0294_));
 sg13g2_xor2_1 _0938_ (.B(net19),
    .A(_0010_),
    .X(_0295_));
 sg13g2_nand2_1 _0939_ (.Y(_0296_),
    .A(_0288_),
    .B(_0295_));
 sg13g2_xnor2_1 _0940_ (.Y(_0297_),
    .A(_0291_),
    .B(_0296_));
 sg13g2_nor2_1 _0941_ (.A(net22),
    .B(_0297_),
    .Y(_0079_));
 sg13g2_buf_2 _0942_ (.A(\enc1[2] ),
    .X(_0298_));
 sg13g2_or2_1 _0943_ (.X(_0299_),
    .B(net19),
    .A(_0290_));
 sg13g2_nand3_1 _0944_ (.B(_0290_),
    .C(net19),
    .A(_0280_),
    .Y(_0300_));
 sg13g2_o21ai_1 _0945_ (.B1(_0300_),
    .Y(_0301_),
    .A1(_0280_),
    .A2(_0299_));
 sg13g2_xnor2_1 _0946_ (.Y(_0302_),
    .A(_0002_),
    .B(_0301_));
 sg13g2_mux2_1 _0947_ (.A0(_0298_),
    .A1(_0302_),
    .S(_0288_),
    .X(_0303_));
 sg13g2_and2_1 _0948_ (.A(net26),
    .B(_0303_),
    .X(_0080_));
 sg13g2_buf_2 _0949_ (.A(\enc1[3] ),
    .X(_0304_));
 sg13g2_nor2_1 _0950_ (.A(_0304_),
    .B(_0288_),
    .Y(_0305_));
 sg13g2_a221oi_1 _0951_ (.B2(_0283_),
    .C1(_0298_),
    .B1(_0286_),
    .A1(_0292_),
    .Y(_0306_),
    .A2(_0285_));
 sg13g2_nand2_1 _0952_ (.Y(_0307_),
    .A(_0291_),
    .B(_0298_));
 sg13g2_nand3b_1 _0953_ (.B(_0307_),
    .C(_0280_),
    .Y(_0308_),
    .A_N(_0306_));
 sg13g2_a21o_1 _0954_ (.A2(_0002_),
    .A1(_0291_),
    .B1(net19),
    .X(_0309_));
 sg13g2_and2_1 _0955_ (.A(_0308_),
    .B(_0309_),
    .X(_0310_));
 sg13g2_xnor2_1 _0956_ (.Y(_0311_),
    .A(_0003_),
    .B(net19));
 sg13g2_xnor2_1 _0957_ (.Y(_0312_),
    .A(_0310_),
    .B(_0311_));
 sg13g2_and2_1 _0958_ (.A(_0288_),
    .B(_0312_),
    .X(_0313_));
 sg13g2_nor3_1 _0959_ (.A(net21),
    .B(_0305_),
    .C(_0313_),
    .Y(_0081_));
 sg13g2_buf_1 _0960_ (.A(\enc1[4] ),
    .X(_0314_));
 sg13g2_a22oi_1 _0961_ (.Y(_0315_),
    .B1(_0286_),
    .B2(_0292_),
    .A2(_0285_),
    .A1(_0283_));
 sg13g2_nor2b_1 _0962_ (.A(_0294_),
    .B_N(_0003_),
    .Y(_0316_));
 sg13g2_nand2_1 _0963_ (.Y(_0317_),
    .A(_0002_),
    .B(_0316_));
 sg13g2_nor2_1 _0964_ (.A(_0298_),
    .B(_0304_),
    .Y(_0318_));
 sg13g2_nor2b_1 _0965_ (.A(net19),
    .B_N(_0318_),
    .Y(_0319_));
 sg13g2_and3_1 _0966_ (.X(_0320_),
    .A(_0290_),
    .B(_0298_),
    .C(_0304_));
 sg13g2_mux2_1 _0967_ (.A0(_0318_),
    .A1(_0320_),
    .S(net19),
    .X(_0321_));
 sg13g2_a22oi_1 _0968_ (.Y(_0322_),
    .B1(_0321_),
    .B2(_0280_),
    .A2(_0319_),
    .A1(_0290_));
 sg13g2_mux2_1 _0969_ (.A0(_0315_),
    .A1(_0317_),
    .S(_0322_),
    .X(_0323_));
 sg13g2_xor2_1 _0970_ (.B(_0323_),
    .A(_0314_),
    .X(_0324_));
 sg13g2_nor2_1 _0971_ (.A(net22),
    .B(_0324_),
    .Y(_0082_));
 sg13g2_buf_2 _0972_ (.A(\enc1[5] ),
    .X(_0325_));
 sg13g2_nor2_1 _0973_ (.A(_0325_),
    .B(_0200_),
    .Y(_0326_));
 sg13g2_and2_1 _0974_ (.A(_0325_),
    .B(net29),
    .X(_0327_));
 sg13g2_nor2b_1 _0975_ (.A(net36),
    .B_N(_0003_),
    .Y(_0328_));
 sg13g2_a22oi_1 _0976_ (.Y(_0329_),
    .B1(_0328_),
    .B2(_0285_),
    .A2(_0286_),
    .A1(net36));
 sg13g2_nor2_1 _0977_ (.A(_0282_),
    .B(_0329_),
    .Y(_0330_));
 sg13g2_a22oi_1 _0978_ (.Y(_0331_),
    .B1(_0286_),
    .B2(_0328_),
    .A2(_0285_),
    .A1(net36));
 sg13g2_nor2_1 _0979_ (.A(_0284_),
    .B(_0331_),
    .Y(_0332_));
 sg13g2_nor2b_1 _0980_ (.A(_0294_),
    .B_N(_0328_),
    .Y(_0333_));
 sg13g2_mux2_1 _0981_ (.A0(_0304_),
    .A1(_0333_),
    .S(_0310_),
    .X(_0334_));
 sg13g2_o21ai_1 _0982_ (.B1(_0334_),
    .Y(_0335_),
    .A1(_0330_),
    .A2(_0332_));
 sg13g2_mux2_1 _0983_ (.A0(_0326_),
    .A1(_0327_),
    .S(_0335_),
    .X(_0083_));
 sg13g2_buf_2 _0984_ (.A(\enc1[6] ),
    .X(_0336_));
 sg13g2_nor2_1 _0985_ (.A(_0336_),
    .B(net21),
    .Y(_0337_));
 sg13g2_inv_1 _0986_ (.Y(_0338_),
    .A(_0336_));
 sg13g2_nor2_1 _0987_ (.A(_0338_),
    .B(_0190_),
    .Y(_0339_));
 sg13g2_nor2_2 _0988_ (.A(net36),
    .B(_0325_),
    .Y(_0340_));
 sg13g2_nand4_1 _0989_ (.B(_0288_),
    .C(_0316_),
    .A(_0002_),
    .Y(_0341_),
    .D(_0340_));
 sg13g2_and2_1 _0990_ (.A(net36),
    .B(_0325_),
    .X(_0342_));
 sg13g2_nor3_1 _0991_ (.A(_0281_),
    .B(\rgb_mixer.debounce1_a.debounced ),
    .C(\rgb_mixer.encoder1.old_a ),
    .Y(_0343_));
 sg13g2_and3_1 _0992_ (.X(_0344_),
    .A(_0281_),
    .B(\rgb_mixer.debounce1_a.debounced ),
    .C(\rgb_mixer.encoder1.old_a ));
 sg13g2_nor2_1 _0993_ (.A(_0343_),
    .B(_0344_),
    .Y(_0345_));
 sg13g2_nand2_1 _0994_ (.Y(_0346_),
    .A(_0342_),
    .B(_0345_));
 sg13g2_a22oi_1 _0995_ (.Y(_0347_),
    .B1(_0343_),
    .B2(_0340_),
    .A2(_0342_),
    .A1(_0281_));
 sg13g2_inv_1 _0996_ (.Y(_0348_),
    .A(_0281_));
 sg13g2_a221oi_1 _0997_ (.B2(_0340_),
    .C1(\rgb_mixer.debounce1_b.debounced ),
    .B1(_0344_),
    .A1(_0348_),
    .Y(_0349_),
    .A2(_0342_));
 sg13g2_a21o_1 _0998_ (.A2(_0347_),
    .A1(\rgb_mixer.debounce1_b.debounced ),
    .B1(_0349_),
    .X(_0350_));
 sg13g2_a21oi_1 _0999_ (.A1(_0346_),
    .A2(_0350_),
    .Y(_0351_),
    .B1(_0322_));
 sg13g2_mux2_1 _1000_ (.A0(_0341_),
    .A1(_0315_),
    .S(_0351_),
    .X(_0352_));
 sg13g2_mux2_1 _1001_ (.A0(_0337_),
    .A1(_0339_),
    .S(_0352_),
    .X(_0084_));
 sg13g2_nand3_1 _1002_ (.B(_0316_),
    .C(_0340_),
    .A(_0338_),
    .Y(_0353_));
 sg13g2_nand2b_1 _1003_ (.Y(_0354_),
    .B(_0336_),
    .A_N(_0315_));
 sg13g2_xor2_1 _1004_ (.B(net19),
    .A(_0304_),
    .X(_0355_));
 sg13g2_a221oi_1 _1005_ (.B2(_0350_),
    .C1(_0355_),
    .B1(_0346_),
    .A1(_0308_),
    .Y(_0356_),
    .A2(_0309_));
 sg13g2_mux2_1 _1006_ (.A0(_0353_),
    .A1(_0354_),
    .S(_0356_),
    .X(_0357_));
 sg13g2_xnor2_1 _1007_ (.Y(_0358_),
    .A(\enc1[7] ),
    .B(_0357_));
 sg13g2_and2_1 _1008_ (.A(net26),
    .B(_0358_),
    .X(_0085_));
 sg13g2_inv_1 _1009_ (.Y(_0086_),
    .A(_0163_));
 sg13g2_inv_1 _1010_ (.Y(_0087_),
    .A(_0171_));
 sg13g2_buf_2 _1011_ (.A(\enc2[0] ),
    .X(_0359_));
 sg13g2_nand2b_1 _1012_ (.Y(_0360_),
    .B(net44),
    .A_N(_0162_));
 sg13g2_nand2b_1 _1013_ (.Y(_0361_),
    .B(_0162_),
    .A_N(net44));
 sg13g2_buf_1 _1014_ (.A(\rgb_mixer.encoder2.old_b ),
    .X(_0362_));
 sg13g2_buf_2 _1015_ (.A(\rgb_mixer.encoder2.old_a ),
    .X(_0363_));
 sg13g2_xor2_1 _1016_ (.B(_0363_),
    .A(_0362_),
    .X(_0364_));
 sg13g2_a21oi_2 _1017_ (.B1(_0364_),
    .Y(_0365_),
    .A2(_0361_),
    .A1(_0360_));
 sg13g2_mux2_1 _1018_ (.A0(_0359_),
    .A1(_0011_),
    .S(_0365_),
    .X(_0366_));
 sg13g2_and2_1 _1019_ (.A(net26),
    .B(_0366_),
    .X(_0088_));
 sg13g2_buf_1 _1020_ (.A(\enc2[1] ),
    .X(_0367_));
 sg13g2_nor2_1 _1021_ (.A(_0362_),
    .B(_0363_),
    .Y(_0368_));
 sg13g2_nor2b_1 _1022_ (.A(_0162_),
    .B_N(\rgb_mixer.debounce2_b.debounced ),
    .Y(_0369_));
 sg13g2_and2_1 _1023_ (.A(_0162_),
    .B(_0363_),
    .X(_0370_));
 sg13g2_nor2b_1 _1024_ (.A(_0170_),
    .B_N(\rgb_mixer.encoder2.old_b ),
    .Y(_0371_));
 sg13g2_a22oi_1 _1025_ (.Y(_0372_),
    .B1(_0370_),
    .B2(_0371_),
    .A2(_0369_),
    .A1(_0368_));
 sg13g2_buf_1 _1026_ (.A(_0372_),
    .X(_0373_));
 sg13g2_xor2_1 _1027_ (.B(net18),
    .A(_0011_),
    .X(_0374_));
 sg13g2_nand2_1 _1028_ (.Y(_0375_),
    .A(_0365_),
    .B(_0374_));
 sg13g2_xor2_1 _1029_ (.B(_0375_),
    .A(net34),
    .X(_0376_));
 sg13g2_nor2_1 _1030_ (.A(net22),
    .B(_0376_),
    .Y(_0089_));
 sg13g2_or2_1 _1031_ (.X(_0377_),
    .B(net34),
    .A(_0359_));
 sg13g2_nand2_1 _1032_ (.Y(_0378_),
    .A(_0359_),
    .B(net34));
 sg13g2_mux2_1 _1033_ (.A0(_0377_),
    .A1(_0378_),
    .S(net18),
    .X(_0379_));
 sg13g2_xor2_1 _1034_ (.B(_0379_),
    .A(_0000_),
    .X(_0380_));
 sg13g2_buf_2 _1035_ (.A(\enc2[2] ),
    .X(_0381_));
 sg13g2_inv_1 _1036_ (.Y(_0382_),
    .A(_0381_));
 sg13g2_nor2_1 _1037_ (.A(_0382_),
    .B(_0365_),
    .Y(_0383_));
 sg13g2_a21oi_1 _1038_ (.A1(_0365_),
    .A2(_0380_),
    .Y(_0384_),
    .B1(_0383_));
 sg13g2_nor2_1 _1039_ (.A(net22),
    .B(_0384_),
    .Y(_0090_));
 sg13g2_nor2b_1 _1040_ (.A(net18),
    .B_N(_0000_),
    .Y(_0385_));
 sg13g2_a21oi_1 _1041_ (.A1(_0359_),
    .A2(_0382_),
    .Y(_0386_),
    .B1(net34));
 sg13g2_nor2_1 _1042_ (.A(_0382_),
    .B(_0378_),
    .Y(_0387_));
 sg13g2_a22oi_1 _1043_ (.Y(_0388_),
    .B1(_0387_),
    .B2(net18),
    .A2(_0386_),
    .A1(_0385_));
 sg13g2_xor2_1 _1044_ (.B(_0388_),
    .A(_0001_),
    .X(_0389_));
 sg13g2_buf_1 _1045_ (.A(\enc2[3] ),
    .X(_0390_));
 sg13g2_nor2b_1 _1046_ (.A(_0365_),
    .B_N(net33),
    .Y(_0391_));
 sg13g2_a21oi_1 _1047_ (.A1(_0365_),
    .A2(_0389_),
    .Y(_0392_),
    .B1(_0391_));
 sg13g2_nor2_1 _1048_ (.A(net22),
    .B(_0392_),
    .Y(_0091_));
 sg13g2_buf_1 _1049_ (.A(\enc2[4] ),
    .X(_0393_));
 sg13g2_nand3b_1 _1050_ (.B(_0162_),
    .C(_0363_),
    .Y(_0394_),
    .A_N(net44));
 sg13g2_inv_1 _1051_ (.Y(_0395_),
    .A(_0363_));
 sg13g2_nand2_1 _1052_ (.Y(_0396_),
    .A(_0395_),
    .B(_0369_));
 sg13g2_and4_1 _1053_ (.A(_0381_),
    .B(net33),
    .C(_0394_),
    .D(_0396_),
    .X(_0397_));
 sg13g2_and3_1 _1054_ (.X(_0398_),
    .A(net44),
    .B(_0381_),
    .C(net33));
 sg13g2_nor3_1 _1055_ (.A(_0381_),
    .B(net33),
    .C(_0394_),
    .Y(_0399_));
 sg13g2_o21ai_1 _1056_ (.B1(net35),
    .Y(_0400_),
    .A1(_0398_),
    .A2(_0399_));
 sg13g2_inv_1 _1057_ (.Y(_0401_),
    .A(net44));
 sg13g2_and3_1 _1058_ (.X(_0402_),
    .A(_0401_),
    .B(_0381_),
    .C(\enc2[3] ));
 sg13g2_nor4_1 _1059_ (.A(_0363_),
    .B(_0381_),
    .C(net33),
    .D(_0360_),
    .Y(_0403_));
 sg13g2_inv_1 _1060_ (.Y(_0404_),
    .A(net35));
 sg13g2_o21ai_1 _1061_ (.B1(_0404_),
    .Y(_0405_),
    .A1(_0402_),
    .A2(_0403_));
 sg13g2_nand3b_1 _1062_ (.B(_0400_),
    .C(_0405_),
    .Y(_0406_),
    .A_N(_0397_));
 sg13g2_nand2_1 _1063_ (.Y(_0407_),
    .A(_0365_),
    .B(net18));
 sg13g2_nor2_1 _1064_ (.A(_0378_),
    .B(_0407_),
    .Y(_0408_));
 sg13g2_and3_1 _1065_ (.X(_0409_),
    .A(_0001_),
    .B(_0385_),
    .C(_0400_));
 sg13g2_nor2b_1 _1066_ (.A(_0397_),
    .B_N(_0405_),
    .Y(_0410_));
 sg13g2_nor2_1 _1067_ (.A(_0359_),
    .B(net34),
    .Y(_0411_));
 sg13g2_and3_1 _1068_ (.X(_0412_),
    .A(_0001_),
    .B(_0411_),
    .C(_0385_));
 sg13g2_a221oi_1 _1069_ (.B2(_0410_),
    .C1(_0412_),
    .B1(_0409_),
    .A1(_0406_),
    .Y(_0413_),
    .A2(_0408_));
 sg13g2_xor2_1 _1070_ (.B(_0413_),
    .A(net32),
    .X(_0414_));
 sg13g2_nor2_1 _1071_ (.A(net22),
    .B(_0414_),
    .Y(_0092_));
 sg13g2_buf_1 _1072_ (.A(\enc2[5] ),
    .X(_0415_));
 sg13g2_nor2_1 _1073_ (.A(net31),
    .B(net21),
    .Y(_0416_));
 sg13g2_and2_1 _1074_ (.A(net31),
    .B(net29),
    .X(_0417_));
 sg13g2_nand2b_1 _1075_ (.Y(_0418_),
    .B(_0001_),
    .A_N(net32));
 sg13g2_nor2_1 _1076_ (.A(net18),
    .B(_0418_),
    .Y(_0419_));
 sg13g2_or4_1 _1077_ (.A(net35),
    .B(net33),
    .C(net32),
    .D(_0396_),
    .X(_0420_));
 sg13g2_nand2_1 _1078_ (.Y(_0421_),
    .A(\enc2[3] ),
    .B(net32));
 sg13g2_a221oi_1 _1079_ (.B2(_0401_),
    .C1(_0421_),
    .B1(_0370_),
    .A1(_0395_),
    .Y(_0422_),
    .A2(_0369_));
 sg13g2_nand2_1 _1080_ (.Y(_0423_),
    .A(net44),
    .B(net35));
 sg13g2_or2_1 _1081_ (.X(_0424_),
    .B(net35),
    .A(net44));
 sg13g2_a21oi_1 _1082_ (.A1(_0423_),
    .A2(_0424_),
    .Y(_0425_),
    .B1(_0421_));
 sg13g2_nor4_1 _1083_ (.A(_0404_),
    .B(net33),
    .C(net32),
    .D(_0394_),
    .Y(_0426_));
 sg13g2_nor3_1 _1084_ (.A(_0422_),
    .B(_0425_),
    .C(_0426_),
    .Y(_0427_));
 sg13g2_o21ai_1 _1085_ (.B1(_0359_),
    .Y(_0428_),
    .A1(_0367_),
    .A2(_0382_));
 sg13g2_a21o_1 _1086_ (.A2(_0372_),
    .A1(_0382_),
    .B1(_0428_),
    .X(_0429_));
 sg13g2_nand2b_1 _1087_ (.Y(_0430_),
    .B(_0000_),
    .A_N(net34));
 sg13g2_nand2b_1 _1088_ (.Y(_0431_),
    .B(_0430_),
    .A_N(_0373_));
 sg13g2_a22oi_1 _1089_ (.Y(_0432_),
    .B1(_0429_),
    .B2(_0431_),
    .A2(_0427_),
    .A1(_0420_));
 sg13g2_mux2_1 _1090_ (.A0(_0419_),
    .A1(_0373_),
    .S(_0432_),
    .X(_0433_));
 sg13g2_nand2_1 _1091_ (.Y(_0434_),
    .A(_0365_),
    .B(_0433_));
 sg13g2_mux2_1 _1092_ (.A0(_0416_),
    .A1(_0417_),
    .S(_0434_),
    .X(_0093_));
 sg13g2_buf_2 _1093_ (.A(\enc2[6] ),
    .X(_0435_));
 sg13g2_inv_1 _1094_ (.Y(_0436_),
    .A(_0435_));
 sg13g2_nor2_1 _1095_ (.A(_0436_),
    .B(_0190_),
    .Y(_0437_));
 sg13g2_nor2_1 _1096_ (.A(_0435_),
    .B(_0190_),
    .Y(_0438_));
 sg13g2_and2_1 _1097_ (.A(_0377_),
    .B(_0406_),
    .X(_0439_));
 sg13g2_nor2_1 _1098_ (.A(net31),
    .B(_0418_),
    .Y(_0440_));
 sg13g2_nand2_1 _1099_ (.Y(_0441_),
    .A(_0385_),
    .B(_0440_));
 sg13g2_nand4_1 _1100_ (.B(net31),
    .C(_0406_),
    .A(net32),
    .Y(_0442_),
    .D(_0408_));
 sg13g2_o21ai_1 _1101_ (.B1(_0442_),
    .Y(_0443_),
    .A1(_0439_),
    .A2(_0441_));
 sg13g2_mux2_1 _1102_ (.A0(_0437_),
    .A1(_0438_),
    .S(_0443_),
    .X(_0094_));
 sg13g2_nor2_1 _1103_ (.A(\enc2[7] ),
    .B(_0190_),
    .Y(_0444_));
 sg13g2_and2_1 _1104_ (.A(\enc2[7] ),
    .B(net29),
    .X(_0445_));
 sg13g2_and2_1 _1105_ (.A(net31),
    .B(_0435_),
    .X(_0446_));
 sg13g2_and2_1 _1106_ (.A(net35),
    .B(_0370_),
    .X(_0447_));
 sg13g2_nor2_1 _1107_ (.A(net31),
    .B(_0435_),
    .Y(_0448_));
 sg13g2_a221oi_1 _1108_ (.B2(_0448_),
    .C1(net44),
    .B1(_0447_),
    .A1(_0404_),
    .Y(_0449_),
    .A2(_0446_));
 sg13g2_nor3_1 _1109_ (.A(net35),
    .B(_0162_),
    .C(_0363_),
    .Y(_0450_));
 sg13g2_a221oi_1 _1110_ (.B2(_0448_),
    .C1(_0401_),
    .B1(_0450_),
    .A1(net35),
    .Y(_0451_),
    .A2(_0446_));
 sg13g2_nand3_1 _1111_ (.B(_0396_),
    .C(_0446_),
    .A(_0394_),
    .Y(_0452_));
 sg13g2_o21ai_1 _1112_ (.B1(_0452_),
    .Y(_0453_),
    .A1(_0449_),
    .A2(_0451_));
 sg13g2_nor2b_1 _1113_ (.A(_0418_),
    .B_N(_0448_),
    .Y(_0454_));
 sg13g2_nor2_1 _1114_ (.A(net18),
    .B(_0454_),
    .Y(_0455_));
 sg13g2_a21oi_1 _1115_ (.A1(_0432_),
    .A2(_0453_),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_mux2_1 _1116_ (.A0(_0407_),
    .A1(net18),
    .S(_0456_),
    .X(_0457_));
 sg13g2_mux2_1 _1117_ (.A0(_0444_),
    .A1(_0445_),
    .S(_0457_),
    .X(_0095_));
 sg13g2_and2_1 _1118_ (.A(net26),
    .B(_0008_),
    .X(_0096_));
 sg13g2_xnor2_1 _1119_ (.Y(_0458_),
    .A(\rgb_mixer.pwm0.count[1] ),
    .B(\rgb_mixer.pwm0.count[0] ));
 sg13g2_nor2_1 _1120_ (.A(_0192_),
    .B(_0458_),
    .Y(_0097_));
 sg13g2_inv_1 _1121_ (.Y(_0459_),
    .A(\rgb_mixer.pwm0.count[2] ));
 sg13g2_nand2_1 _1122_ (.Y(_0460_),
    .A(\rgb_mixer.pwm0.count[1] ),
    .B(\rgb_mixer.pwm0.count[0] ));
 sg13g2_xnor2_1 _1123_ (.Y(_0461_),
    .A(_0459_),
    .B(_0460_));
 sg13g2_nor2_1 _1124_ (.A(net22),
    .B(_0461_),
    .Y(_0098_));
 sg13g2_inv_1 _1125_ (.Y(_0462_),
    .A(\rgb_mixer.pwm0.count[3] ));
 sg13g2_nand3_1 _1126_ (.B(\rgb_mixer.pwm0.count[1] ),
    .C(\rgb_mixer.pwm0.count[0] ),
    .A(\rgb_mixer.pwm0.count[2] ),
    .Y(_0463_));
 sg13g2_xnor2_1 _1127_ (.Y(_0464_),
    .A(_0462_),
    .B(_0463_));
 sg13g2_nor2_1 _1128_ (.A(net22),
    .B(_0464_),
    .Y(_0099_));
 sg13g2_buf_1 _1129_ (.A(_0190_),
    .X(_0465_));
 sg13g2_buf_1 _1130_ (.A(\rgb_mixer.pwm0.count[4] ),
    .X(_0466_));
 sg13g2_nor2_2 _1131_ (.A(_0462_),
    .B(_0463_),
    .Y(_0467_));
 sg13g2_xnor2_1 _1132_ (.Y(_0468_),
    .A(_0466_),
    .B(_0467_));
 sg13g2_nor2_1 _1133_ (.A(net20),
    .B(_0468_),
    .Y(_0100_));
 sg13g2_inv_1 _1134_ (.Y(_0469_),
    .A(\rgb_mixer.pwm0.count[5] ));
 sg13g2_nand2_1 _1135_ (.Y(_0470_),
    .A(_0466_),
    .B(_0467_));
 sg13g2_xnor2_1 _1136_ (.Y(_0471_),
    .A(_0469_),
    .B(_0470_));
 sg13g2_nor2_1 _1137_ (.A(net20),
    .B(_0471_),
    .Y(_0101_));
 sg13g2_nand3_1 _1138_ (.B(_0466_),
    .C(_0467_),
    .A(\rgb_mixer.pwm0.count[5] ),
    .Y(_0472_));
 sg13g2_xor2_1 _1139_ (.B(_0472_),
    .A(\rgb_mixer.pwm0.count[6] ),
    .X(_0473_));
 sg13g2_nor2_1 _1140_ (.A(_0465_),
    .B(_0473_),
    .Y(_0102_));
 sg13g2_nand4_1 _1141_ (.B(\rgb_mixer.pwm0.count[5] ),
    .C(_0466_),
    .A(\rgb_mixer.pwm0.count[6] ),
    .Y(_0474_),
    .D(_0467_));
 sg13g2_xor2_1 _1142_ (.B(_0474_),
    .A(\rgb_mixer.pwm0.count[7] ),
    .X(_0475_));
 sg13g2_nor2_1 _1143_ (.A(_0465_),
    .B(_0475_),
    .Y(_0103_));
 sg13g2_nand2b_1 _1144_ (.Y(_0476_),
    .B(net37),
    .A_N(\rgb_mixer.pwm0.count[6] ));
 sg13g2_inv_1 _1145_ (.Y(_0477_),
    .A(\enc0[7] ));
 sg13g2_o21ai_1 _1146_ (.B1(_0477_),
    .Y(_0478_),
    .A1(\rgb_mixer.pwm0.count[7] ),
    .A2(_0476_));
 sg13g2_nand2_1 _1147_ (.Y(_0479_),
    .A(\rgb_mixer.pwm0.count[7] ),
    .B(_0476_));
 sg13g2_a22oi_1 _1148_ (.Y(_0480_),
    .B1(_0478_),
    .B2(_0479_),
    .A2(net38),
    .A1(_0469_));
 sg13g2_inv_1 _1149_ (.Y(_0481_),
    .A(net40));
 sg13g2_nand2_1 _1150_ (.Y(_0482_),
    .A(_0459_),
    .B(net41));
 sg13g2_inv_1 _1151_ (.Y(_0483_),
    .A(\rgb_mixer.pwm0.count[0] ));
 sg13g2_a21oi_1 _1152_ (.A1(_0483_),
    .A2(_0187_),
    .Y(_0484_),
    .B1(net42));
 sg13g2_nand3_1 _1153_ (.B(_0483_),
    .C(_0187_),
    .A(net42),
    .Y(_0485_));
 sg13g2_o21ai_1 _1154_ (.B1(_0485_),
    .Y(_0486_),
    .A1(\rgb_mixer.pwm0.count[1] ),
    .A2(_0484_));
 sg13g2_o21ai_1 _1155_ (.B1(_0486_),
    .Y(_0487_),
    .A1(_0459_),
    .A2(net41));
 sg13g2_a22oi_1 _1156_ (.Y(_0488_),
    .B1(_0482_),
    .B2(_0487_),
    .A2(_0481_),
    .A1(\rgb_mixer.pwm0.count[3] ));
 sg13g2_nand2b_1 _1157_ (.Y(_0489_),
    .B(net39),
    .A_N(_0466_));
 sg13g2_o21ai_1 _1158_ (.B1(_0489_),
    .Y(_0490_),
    .A1(\rgb_mixer.pwm0.count[3] ),
    .A2(_0481_));
 sg13g2_nand2b_1 _1159_ (.Y(_0491_),
    .B(_0466_),
    .A_N(net39));
 sg13g2_o21ai_1 _1160_ (.B1(_0491_),
    .Y(_0492_),
    .A1(_0488_),
    .A2(_0490_));
 sg13g2_nand2b_1 _1161_ (.Y(_0493_),
    .B(\rgb_mixer.pwm0.count[5] ),
    .A_N(net38));
 sg13g2_nor2_1 _1162_ (.A(net37),
    .B(_0493_),
    .Y(_0494_));
 sg13g2_nor2_1 _1163_ (.A(\rgb_mixer.pwm0.count[6] ),
    .B(_0494_),
    .Y(_0495_));
 sg13g2_a21oi_1 _1164_ (.A1(net37),
    .A2(_0493_),
    .Y(_0496_),
    .B1(_0495_));
 sg13g2_a21oi_1 _1165_ (.A1(\rgb_mixer.pwm0.count[7] ),
    .A2(_0496_),
    .Y(_0497_),
    .B1(_0477_));
 sg13g2_nor2_1 _1166_ (.A(\rgb_mixer.pwm0.count[7] ),
    .B(_0496_),
    .Y(_0498_));
 sg13g2_o21ai_1 _1167_ (.B1(net29),
    .Y(_0499_),
    .A1(_0497_),
    .A2(_0498_));
 sg13g2_a21oi_1 _1168_ (.A1(_0480_),
    .A2(_0492_),
    .Y(_0104_),
    .B1(_0499_));
 sg13g2_and2_1 _1169_ (.A(net27),
    .B(_0007_),
    .X(_0105_));
 sg13g2_xnor2_1 _1170_ (.Y(_0500_),
    .A(\rgb_mixer.pwm1.count[1] ),
    .B(\rgb_mixer.pwm1.count[0] ));
 sg13g2_nor2_1 _1171_ (.A(net20),
    .B(_0500_),
    .Y(_0106_));
 sg13g2_nand2_1 _1172_ (.Y(_0501_),
    .A(\rgb_mixer.pwm1.count[1] ),
    .B(\rgb_mixer.pwm1.count[0] ));
 sg13g2_xor2_1 _1173_ (.B(_0501_),
    .A(\rgb_mixer.pwm1.count[2] ),
    .X(_0502_));
 sg13g2_nor2_1 _1174_ (.A(net20),
    .B(_0502_),
    .Y(_0107_));
 sg13g2_inv_1 _1175_ (.Y(_0503_),
    .A(\rgb_mixer.pwm1.count[3] ));
 sg13g2_nand3_1 _1176_ (.B(\rgb_mixer.pwm1.count[1] ),
    .C(\rgb_mixer.pwm1.count[0] ),
    .A(\rgb_mixer.pwm1.count[2] ),
    .Y(_0504_));
 sg13g2_xnor2_1 _1177_ (.Y(_0505_),
    .A(_0503_),
    .B(_0504_));
 sg13g2_nor2_1 _1178_ (.A(net20),
    .B(_0505_),
    .Y(_0108_));
 sg13g2_nor2_1 _1179_ (.A(_0503_),
    .B(_0504_),
    .Y(_0506_));
 sg13g2_xnor2_1 _1180_ (.Y(_0507_),
    .A(\rgb_mixer.pwm1.count[4] ),
    .B(_0506_));
 sg13g2_nor2_1 _1181_ (.A(net20),
    .B(_0507_),
    .Y(_0109_));
 sg13g2_inv_1 _1182_ (.Y(_0508_),
    .A(\rgb_mixer.pwm1.count[5] ));
 sg13g2_nand2_1 _1183_ (.Y(_0509_),
    .A(\rgb_mixer.pwm1.count[4] ),
    .B(_0506_));
 sg13g2_xnor2_1 _1184_ (.Y(_0510_),
    .A(_0508_),
    .B(_0509_));
 sg13g2_nor2_1 _1185_ (.A(net20),
    .B(_0510_),
    .Y(_0110_));
 sg13g2_inv_1 _1186_ (.Y(_0511_),
    .A(\rgb_mixer.pwm1.count[6] ));
 sg13g2_nand3_1 _1187_ (.B(\rgb_mixer.pwm1.count[4] ),
    .C(_0506_),
    .A(\rgb_mixer.pwm1.count[5] ),
    .Y(_0512_));
 sg13g2_xnor2_1 _1188_ (.Y(_0513_),
    .A(_0511_),
    .B(_0512_));
 sg13g2_nor2_1 _1189_ (.A(net20),
    .B(_0513_),
    .Y(_0111_));
 sg13g2_or2_1 _1190_ (.X(_0514_),
    .B(_0512_),
    .A(_0511_));
 sg13g2_xor2_1 _1191_ (.B(_0514_),
    .A(\rgb_mixer.pwm1.count[7] ),
    .X(_0515_));
 sg13g2_nor2_1 _1192_ (.A(net23),
    .B(_0515_),
    .Y(_0112_));
 sg13g2_nand2b_1 _1193_ (.Y(_0516_),
    .B(\rgb_mixer.pwm1.count[7] ),
    .A_N(\enc1[7] ));
 sg13g2_nand2b_1 _1194_ (.Y(_0517_),
    .B(\rgb_mixer.pwm1.count[5] ),
    .A_N(_0325_));
 sg13g2_xnor2_1 _1195_ (.Y(_0518_),
    .A(_0336_),
    .B(\rgb_mixer.pwm1.count[6] ));
 sg13g2_nand2b_1 _1196_ (.Y(_0519_),
    .B(\rgb_mixer.pwm1.count[2] ),
    .A_N(_0298_));
 sg13g2_inv_1 _1197_ (.Y(_0520_),
    .A(\rgb_mixer.pwm1.count[1] ));
 sg13g2_inv_1 _1198_ (.Y(_0521_),
    .A(\rgb_mixer.pwm1.count[0] ));
 sg13g2_a22oi_1 _1199_ (.Y(_0522_),
    .B1(_0521_),
    .B2(_0280_),
    .A2(_0520_),
    .A1(_0290_));
 sg13g2_a21oi_1 _1200_ (.A1(_0291_),
    .A2(\rgb_mixer.pwm1.count[1] ),
    .Y(_0523_),
    .B1(_0522_));
 sg13g2_nor2b_1 _1201_ (.A(\rgb_mixer.pwm1.count[2] ),
    .B_N(_0298_),
    .Y(_0524_));
 sg13g2_a221oi_1 _1202_ (.B2(_0523_),
    .C1(_0524_),
    .B1(_0519_),
    .A1(_0304_),
    .Y(_0525_),
    .A2(_0503_));
 sg13g2_nand2b_1 _1203_ (.Y(_0526_),
    .B(\rgb_mixer.pwm1.count[4] ),
    .A_N(net36));
 sg13g2_o21ai_1 _1204_ (.B1(_0526_),
    .Y(_0527_),
    .A1(_0304_),
    .A2(_0503_));
 sg13g2_nand2b_1 _1205_ (.Y(_0528_),
    .B(net36),
    .A_N(\rgb_mixer.pwm1.count[4] ));
 sg13g2_o21ai_1 _1206_ (.B1(_0528_),
    .Y(_0529_),
    .A1(_0525_),
    .A2(_0527_));
 sg13g2_nand4_1 _1207_ (.B(_0517_),
    .C(_0518_),
    .A(_0516_),
    .Y(_0530_),
    .D(_0529_));
 sg13g2_a22oi_1 _1208_ (.Y(_0531_),
    .B1(_0508_),
    .B2(_0325_),
    .A2(_0511_),
    .A1(_0336_));
 sg13g2_a21oi_1 _1209_ (.A1(_0338_),
    .A2(\rgb_mixer.pwm1.count[6] ),
    .Y(_0532_),
    .B1(_0531_));
 sg13g2_nor2b_1 _1210_ (.A(\rgb_mixer.pwm1.count[7] ),
    .B_N(\enc1[7] ),
    .Y(_0533_));
 sg13g2_a21oi_1 _1211_ (.A1(_0516_),
    .A2(_0532_),
    .Y(_0534_),
    .B1(_0533_));
 sg13g2_a21oi_1 _1212_ (.A1(_0530_),
    .A2(_0534_),
    .Y(_0113_),
    .B1(net21));
 sg13g2_and2_1 _1213_ (.A(net27),
    .B(_0006_),
    .X(_0114_));
 sg13g2_xnor2_1 _1214_ (.Y(_0535_),
    .A(\rgb_mixer.pwm2.count[1] ),
    .B(\rgb_mixer.pwm2.count[0] ));
 sg13g2_nor2_1 _1215_ (.A(net23),
    .B(_0535_),
    .Y(_0115_));
 sg13g2_inv_1 _1216_ (.Y(_0536_),
    .A(\rgb_mixer.pwm2.count[2] ));
 sg13g2_nand2_1 _1217_ (.Y(_0537_),
    .A(\rgb_mixer.pwm2.count[1] ),
    .B(\rgb_mixer.pwm2.count[0] ));
 sg13g2_xnor2_1 _1218_ (.Y(_0538_),
    .A(_0536_),
    .B(_0537_));
 sg13g2_nor2_1 _1219_ (.A(net23),
    .B(_0538_),
    .Y(_0116_));
 sg13g2_inv_1 _1220_ (.Y(_0539_),
    .A(\rgb_mixer.pwm2.count[3] ));
 sg13g2_nand3_1 _1221_ (.B(\rgb_mixer.pwm2.count[1] ),
    .C(\rgb_mixer.pwm2.count[0] ),
    .A(\rgb_mixer.pwm2.count[2] ),
    .Y(_0540_));
 sg13g2_xnor2_1 _1222_ (.Y(_0541_),
    .A(_0539_),
    .B(_0540_));
 sg13g2_nor2_1 _1223_ (.A(net23),
    .B(_0541_),
    .Y(_0117_));
 sg13g2_nor2_1 _1224_ (.A(_0539_),
    .B(_0540_),
    .Y(_0542_));
 sg13g2_xnor2_1 _1225_ (.Y(_0543_),
    .A(\rgb_mixer.pwm2.count[4] ),
    .B(_0542_));
 sg13g2_nor2_1 _1226_ (.A(net23),
    .B(_0543_),
    .Y(_0118_));
 sg13g2_inv_1 _1227_ (.Y(_0544_),
    .A(\rgb_mixer.pwm2.count[5] ));
 sg13g2_nand2_1 _1228_ (.Y(_0545_),
    .A(\rgb_mixer.pwm2.count[4] ),
    .B(_0542_));
 sg13g2_xnor2_1 _1229_ (.Y(_0546_),
    .A(_0544_),
    .B(_0545_));
 sg13g2_nor2_1 _1230_ (.A(net23),
    .B(_0546_),
    .Y(_0119_));
 sg13g2_inv_1 _1231_ (.Y(_0547_),
    .A(\rgb_mixer.pwm2.count[6] ));
 sg13g2_nand3_1 _1232_ (.B(\rgb_mixer.pwm2.count[4] ),
    .C(_0542_),
    .A(\rgb_mixer.pwm2.count[5] ),
    .Y(_0548_));
 sg13g2_xnor2_1 _1233_ (.Y(_0549_),
    .A(_0547_),
    .B(_0548_));
 sg13g2_nor2_1 _1234_ (.A(net23),
    .B(_0549_),
    .Y(_0120_));
 sg13g2_or2_1 _1235_ (.X(_0550_),
    .B(_0548_),
    .A(_0547_));
 sg13g2_xor2_1 _1236_ (.B(_0550_),
    .A(\rgb_mixer.pwm2.count[7] ),
    .X(_0551_));
 sg13g2_nor2_1 _1237_ (.A(net23),
    .B(_0551_),
    .Y(_0121_));
 sg13g2_nand2b_1 _1238_ (.Y(_0552_),
    .B(\rgb_mixer.pwm2.count[7] ),
    .A_N(\enc2[7] ));
 sg13g2_nand2b_1 _1239_ (.Y(_0553_),
    .B(\rgb_mixer.pwm2.count[5] ),
    .A_N(net31));
 sg13g2_xnor2_1 _1240_ (.Y(_0554_),
    .A(_0435_),
    .B(\rgb_mixer.pwm2.count[6] ));
 sg13g2_nand2b_1 _1241_ (.Y(_0555_),
    .B(net34),
    .A_N(\rgb_mixer.pwm2.count[1] ));
 sg13g2_nand2b_1 _1242_ (.Y(_0556_),
    .B(\rgb_mixer.pwm2.count[1] ),
    .A_N(net34));
 sg13g2_nand3b_1 _1243_ (.B(_0556_),
    .C(_0359_),
    .Y(_0557_),
    .A_N(\rgb_mixer.pwm2.count[0] ));
 sg13g2_a22oi_1 _1244_ (.Y(_0558_),
    .B1(_0555_),
    .B2(_0557_),
    .A2(\rgb_mixer.pwm2.count[2] ),
    .A1(_0382_));
 sg13g2_a221oi_1 _1245_ (.B2(_0381_),
    .C1(_0558_),
    .B1(_0536_),
    .A1(net33),
    .Y(_0559_),
    .A2(_0539_));
 sg13g2_nand2b_1 _1246_ (.Y(_0560_),
    .B(\rgb_mixer.pwm2.count[4] ),
    .A_N(net32));
 sg13g2_o21ai_1 _1247_ (.B1(_0560_),
    .Y(_0561_),
    .A1(_0390_),
    .A2(_0539_));
 sg13g2_nand2b_1 _1248_ (.Y(_0562_),
    .B(_0393_),
    .A_N(\rgb_mixer.pwm2.count[4] ));
 sg13g2_o21ai_1 _1249_ (.B1(_0562_),
    .Y(_0563_),
    .A1(_0559_),
    .A2(_0561_));
 sg13g2_nand4_1 _1250_ (.B(_0553_),
    .C(_0554_),
    .A(_0552_),
    .Y(_0564_),
    .D(_0563_));
 sg13g2_a22oi_1 _1251_ (.Y(_0565_),
    .B1(_0544_),
    .B2(_0415_),
    .A2(_0547_),
    .A1(_0435_));
 sg13g2_a21oi_1 _1252_ (.A1(_0436_),
    .A2(\rgb_mixer.pwm2.count[6] ),
    .Y(_0566_),
    .B1(_0565_));
 sg13g2_nor2b_1 _1253_ (.A(\rgb_mixer.pwm2.count[7] ),
    .B_N(\enc2[7] ),
    .Y(_0567_));
 sg13g2_a21oi_1 _1254_ (.A1(_0552_),
    .A2(_0566_),
    .Y(_0568_),
    .B1(_0567_));
 sg13g2_a21oi_1 _1255_ (.A1(_0564_),
    .A2(_0568_),
    .Y(_0122_),
    .B1(net21));
 sg13g2_buf_1 _1256_ (.A(ui_in[6]),
    .X(_0569_));
 sg13g2_buf_2 _1257_ (.A(ui_in[7]),
    .X(_0570_));
 sg13g2_buf_1 _1258_ (.A(_0570_),
    .X(_0571_));
 sg13g2_nor2b_1 _1259_ (.A(net30),
    .B_N(_0187_),
    .Y(_0572_));
 sg13g2_a21oi_1 _1260_ (.A1(_0571_),
    .A2(_0359_),
    .Y(_0573_),
    .B1(_0572_));
 sg13g2_nor2b_1 _1261_ (.A(_0570_),
    .B_N(net47),
    .Y(_0574_));
 sg13g2_buf_2 _1262_ (.A(_0574_),
    .X(_0575_));
 sg13g2_nand2_1 _1263_ (.Y(_0576_),
    .A(_0280_),
    .B(_0575_));
 sg13g2_o21ai_1 _1264_ (.B1(_0576_),
    .Y(net7),
    .A1(net47),
    .A2(_0573_));
 sg13g2_nor2b_1 _1265_ (.A(_0571_),
    .B_N(_0193_),
    .Y(_0577_));
 sg13g2_a21oi_1 _1266_ (.A1(net30),
    .A2(_0367_),
    .Y(_0578_),
    .B1(_0577_));
 sg13g2_nand2_1 _1267_ (.Y(_0579_),
    .A(_0290_),
    .B(_0575_));
 sg13g2_o21ai_1 _1268_ (.B1(_0579_),
    .Y(net8),
    .A1(net47),
    .A2(_0578_));
 sg13g2_nor2b_1 _1269_ (.A(_0570_),
    .B_N(net41),
    .Y(_0580_));
 sg13g2_a21oi_1 _1270_ (.A1(net30),
    .A2(_0381_),
    .Y(_0581_),
    .B1(_0580_));
 sg13g2_nand2_1 _1271_ (.Y(_0582_),
    .A(_0298_),
    .B(_0575_));
 sg13g2_o21ai_1 _1272_ (.B1(_0582_),
    .Y(net9),
    .A1(net47),
    .A2(_0581_));
 sg13g2_nor2_1 _1273_ (.A(_0570_),
    .B(_0481_),
    .Y(_0583_));
 sg13g2_a21oi_1 _1274_ (.A1(net30),
    .A2(_0390_),
    .Y(_0584_),
    .B1(_0583_));
 sg13g2_nand2_1 _1275_ (.Y(_0585_),
    .A(_0304_),
    .B(_0575_));
 sg13g2_o21ai_1 _1276_ (.B1(_0585_),
    .Y(net10),
    .A1(_0569_),
    .A2(_0584_));
 sg13g2_nor2b_1 _1277_ (.A(_0570_),
    .B_N(net39),
    .Y(_0586_));
 sg13g2_a21oi_1 _1278_ (.A1(net30),
    .A2(net32),
    .Y(_0587_),
    .B1(_0586_));
 sg13g2_nand2_1 _1279_ (.Y(_0588_),
    .A(net36),
    .B(_0575_));
 sg13g2_o21ai_1 _1280_ (.B1(_0588_),
    .Y(net11),
    .A1(net47),
    .A2(_0587_));
 sg13g2_nor2b_1 _1281_ (.A(_0570_),
    .B_N(net38),
    .Y(_0589_));
 sg13g2_a21oi_1 _1282_ (.A1(net30),
    .A2(net31),
    .Y(_0590_),
    .B1(_0589_));
 sg13g2_nand2_1 _1283_ (.Y(_0591_),
    .A(_0325_),
    .B(_0575_));
 sg13g2_o21ai_1 _1284_ (.B1(_0591_),
    .Y(net12),
    .A1(net47),
    .A2(_0590_));
 sg13g2_nor2b_1 _1285_ (.A(_0570_),
    .B_N(net37),
    .Y(_0592_));
 sg13g2_a21oi_1 _1286_ (.A1(net30),
    .A2(_0435_),
    .Y(_0593_),
    .B1(_0592_));
 sg13g2_nand2_1 _1287_ (.Y(_0594_),
    .A(_0336_),
    .B(_0575_));
 sg13g2_o21ai_1 _1288_ (.B1(_0594_),
    .Y(net13),
    .A1(net47),
    .A2(_0593_));
 sg13g2_nor2_1 _1289_ (.A(_0570_),
    .B(_0477_),
    .Y(_0595_));
 sg13g2_a21oi_1 _1290_ (.A1(net30),
    .A2(\enc2[7] ),
    .Y(_0596_),
    .B1(_0595_));
 sg13g2_nand2_1 _1291_ (.Y(_0597_),
    .A(\enc1[7] ),
    .B(_0575_));
 sg13g2_o21ai_1 _1292_ (.B1(_0597_),
    .Y(net14),
    .A1(net47),
    .A2(_0596_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _1295__53 (.L_HI(net53));
 sg13g2_buf_1 _1295_ (.A(net53),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1296_ (.A(net54),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1297_ (.A(net55),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1298_ (.A(net56),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1299_ (.A(net57),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1300_ (.A(net58),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1301_ (.A(net59),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1302_ (.A(net60),
    .X(uio_oe[7]));
 sg13g2_buf_1 _1303_ (.A(\rgb_mixer.pwm0.out ),
    .X(net15));
 sg13g2_buf_1 _1304_ (.A(\rgb_mixer.pwm1.out ),
    .X(net16));
 sg13g2_buf_1 _1305_ (.A(\rgb_mixer.pwm2.out ),
    .X(net17));
 sg13g2_buf_1 _1306_ (.A(net48),
    .X(uo_out[3]));
 sg13g2_buf_1 _1307_ (.A(net49),
    .X(uo_out[4]));
 sg13g2_buf_1 _1308_ (.A(net50),
    .X(uo_out[5]));
 sg13g2_buf_1 _1309_ (.A(net51),
    .X(uo_out[6]));
 sg13g2_buf_1 _1310_ (.A(net52),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_a.button_hist[0]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net61),
    .D(_0012_),
    .Q_N(_0696_),
    .Q(\rgb_mixer.debounce0_a.button_hist[0] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_a.button_hist[1]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net62),
    .D(_0013_),
    .Q_N(_0695_),
    .Q(\rgb_mixer.debounce0_a.button_hist[1] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_a.button_hist[2]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net63),
    .D(_0014_),
    .Q_N(_0694_),
    .Q(\rgb_mixer.debounce0_a.button_hist[2] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_a.button_hist[3]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net64),
    .D(_0015_),
    .Q_N(_0693_),
    .Q(\rgb_mixer.debounce0_a.button_hist[3] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_a.button_hist[4]$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net65),
    .D(_0016_),
    .Q_N(_0692_),
    .Q(\rgb_mixer.debounce0_a.button_hist[4] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_a.button_hist[5]$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net66),
    .D(_0017_),
    .Q_N(_0691_),
    .Q(\rgb_mixer.debounce0_a.button_hist[5] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_a.button_hist[6]$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net67),
    .D(_0018_),
    .Q_N(_0690_),
    .Q(\rgb_mixer.debounce0_a.button_hist[6] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_a.button_hist[7]$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net68),
    .D(_0019_),
    .Q_N(_0689_),
    .Q(\rgb_mixer.debounce0_a.button_hist[7] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_a.debounced$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net69),
    .D(_0020_),
    .Q_N(_0688_),
    .Q(\rgb_mixer.debounce0_a.debounced ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_b.button_hist[0]$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net70),
    .D(_0021_),
    .Q_N(_0687_),
    .Q(\rgb_mixer.debounce0_b.button_hist[0] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_b.button_hist[1]$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net71),
    .D(_0022_),
    .Q_N(_0686_),
    .Q(\rgb_mixer.debounce0_b.button_hist[1] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_b.button_hist[2]$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net72),
    .D(_0023_),
    .Q_N(_0685_),
    .Q(\rgb_mixer.debounce0_b.button_hist[2] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_b.button_hist[3]$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net73),
    .D(_0024_),
    .Q_N(_0684_),
    .Q(\rgb_mixer.debounce0_b.button_hist[3] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_b.button_hist[4]$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net74),
    .D(_0025_),
    .Q_N(_0683_),
    .Q(\rgb_mixer.debounce0_b.button_hist[4] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_b.button_hist[5]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net75),
    .D(_0026_),
    .Q_N(_0682_),
    .Q(\rgb_mixer.debounce0_b.button_hist[5] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_b.button_hist[6]$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net76),
    .D(_0027_),
    .Q_N(_0681_),
    .Q(\rgb_mixer.debounce0_b.button_hist[6] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_b.button_hist[7]$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net77),
    .D(_0028_),
    .Q_N(_0680_),
    .Q(\rgb_mixer.debounce0_b.button_hist[7] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce0_b.debounced$_SDFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net78),
    .D(_0029_),
    .Q_N(_0679_),
    .Q(\rgb_mixer.debounce0_b.debounced ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_a.button_hist[0]$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net79),
    .D(_0030_),
    .Q_N(_0678_),
    .Q(\rgb_mixer.debounce1_a.button_hist[0] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_a.button_hist[1]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net80),
    .D(_0031_),
    .Q_N(_0677_),
    .Q(\rgb_mixer.debounce1_a.button_hist[1] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_a.button_hist[2]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net81),
    .D(_0032_),
    .Q_N(_0676_),
    .Q(\rgb_mixer.debounce1_a.button_hist[2] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_a.button_hist[3]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net82),
    .D(_0033_),
    .Q_N(_0675_),
    .Q(\rgb_mixer.debounce1_a.button_hist[3] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_a.button_hist[4]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net83),
    .D(_0034_),
    .Q_N(_0674_),
    .Q(\rgb_mixer.debounce1_a.button_hist[4] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_a.button_hist[5]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net84),
    .D(_0035_),
    .Q_N(_0673_),
    .Q(\rgb_mixer.debounce1_a.button_hist[5] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_a.button_hist[6]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net85),
    .D(_0036_),
    .Q_N(_0672_),
    .Q(\rgb_mixer.debounce1_a.button_hist[6] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_a.button_hist[7]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net86),
    .D(_0037_),
    .Q_N(_0671_),
    .Q(\rgb_mixer.debounce1_a.button_hist[7] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_a.debounced$_SDFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net87),
    .D(_0038_),
    .Q_N(_0670_),
    .Q(\rgb_mixer.debounce1_a.debounced ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_b.button_hist[0]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net88),
    .D(_0039_),
    .Q_N(_0669_),
    .Q(\rgb_mixer.debounce1_b.button_hist[0] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_b.button_hist[1]$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net89),
    .D(_0040_),
    .Q_N(_0668_),
    .Q(\rgb_mixer.debounce1_b.button_hist[1] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_b.button_hist[2]$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net90),
    .D(_0041_),
    .Q_N(_0667_),
    .Q(\rgb_mixer.debounce1_b.button_hist[2] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_b.button_hist[3]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net91),
    .D(_0042_),
    .Q_N(_0666_),
    .Q(\rgb_mixer.debounce1_b.button_hist[3] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_b.button_hist[4]$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net92),
    .D(_0043_),
    .Q_N(_0665_),
    .Q(\rgb_mixer.debounce1_b.button_hist[4] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_b.button_hist[5]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net93),
    .D(_0044_),
    .Q_N(_0664_),
    .Q(\rgb_mixer.debounce1_b.button_hist[5] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_b.button_hist[6]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net94),
    .D(_0045_),
    .Q_N(_0663_),
    .Q(\rgb_mixer.debounce1_b.button_hist[6] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_b.button_hist[7]$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net95),
    .D(_0046_),
    .Q_N(_0662_),
    .Q(\rgb_mixer.debounce1_b.button_hist[7] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce1_b.debounced$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net96),
    .D(_0047_),
    .Q_N(_0661_),
    .Q(\rgb_mixer.debounce1_b.debounced ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_a.button_hist[0]$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net97),
    .D(_0048_),
    .Q_N(_0660_),
    .Q(\rgb_mixer.debounce2_a.button_hist[0] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_a.button_hist[1]$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net98),
    .D(_0049_),
    .Q_N(_0659_),
    .Q(\rgb_mixer.debounce2_a.button_hist[1] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_a.button_hist[2]$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net99),
    .D(_0050_),
    .Q_N(_0658_),
    .Q(\rgb_mixer.debounce2_a.button_hist[2] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_a.button_hist[3]$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net100),
    .D(_0051_),
    .Q_N(_0657_),
    .Q(\rgb_mixer.debounce2_a.button_hist[3] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_a.button_hist[4]$_SDFF_PN0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net101),
    .D(_0052_),
    .Q_N(_0656_),
    .Q(\rgb_mixer.debounce2_a.button_hist[4] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_a.button_hist[5]$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net102),
    .D(_0053_),
    .Q_N(_0655_),
    .Q(\rgb_mixer.debounce2_a.button_hist[5] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_a.button_hist[6]$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net103),
    .D(_0054_),
    .Q_N(_0654_),
    .Q(\rgb_mixer.debounce2_a.button_hist[6] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_a.button_hist[7]$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net104),
    .D(_0055_),
    .Q_N(_0653_),
    .Q(\rgb_mixer.debounce2_a.button_hist[7] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_a.debounced$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net105),
    .D(_0056_),
    .Q_N(_0652_),
    .Q(\rgb_mixer.debounce2_a.debounced ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_b.button_hist[0]$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net106),
    .D(_0057_),
    .Q_N(_0651_),
    .Q(\rgb_mixer.debounce2_b.button_hist[0] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_b.button_hist[1]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net107),
    .D(_0058_),
    .Q_N(_0650_),
    .Q(\rgb_mixer.debounce2_b.button_hist[1] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_b.button_hist[2]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net108),
    .D(_0059_),
    .Q_N(_0649_),
    .Q(\rgb_mixer.debounce2_b.button_hist[2] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_b.button_hist[3]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net109),
    .D(_0060_),
    .Q_N(_0648_),
    .Q(\rgb_mixer.debounce2_b.button_hist[3] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_b.button_hist[4]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net110),
    .D(_0061_),
    .Q_N(_0647_),
    .Q(\rgb_mixer.debounce2_b.button_hist[4] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_b.button_hist[5]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net111),
    .D(_0062_),
    .Q_N(_0646_),
    .Q(\rgb_mixer.debounce2_b.button_hist[5] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_b.button_hist[6]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net112),
    .D(_0063_),
    .Q_N(_0645_),
    .Q(\rgb_mixer.debounce2_b.button_hist[6] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_b.button_hist[7]$_SDFF_PN0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net113),
    .D(_0064_),
    .Q_N(_0644_),
    .Q(\rgb_mixer.debounce2_b.button_hist[7] ));
 sg13g2_dfrbp_1 \rgb_mixer.debounce2_b.debounced$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net114),
    .D(_0065_),
    .Q_N(_0643_),
    .Q(\rgb_mixer.debounce2_b.debounced ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder0.old_a$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net115),
    .D(_0066_),
    .Q_N(_0642_),
    .Q(\rgb_mixer.encoder0.old_a ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder0.old_b$_SDFF_PN0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net116),
    .D(_0067_),
    .Q_N(_0641_),
    .Q(\rgb_mixer.encoder0.old_b ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder0.value[0]$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net117),
    .D(_0068_),
    .Q_N(_0009_),
    .Q(\enc0[0] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder0.value[1]$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net118),
    .D(_0069_),
    .Q_N(_0640_),
    .Q(\enc0[1] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder0.value[2]$_SDFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net119),
    .D(_0070_),
    .Q_N(_0004_),
    .Q(\enc0[2] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder0.value[3]$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net120),
    .D(_0071_),
    .Q_N(_0005_),
    .Q(\enc0[3] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder0.value[4]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net121),
    .D(_0072_),
    .Q_N(_0639_),
    .Q(\enc0[4] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder0.value[5]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net122),
    .D(_0073_),
    .Q_N(_0638_),
    .Q(\enc0[5] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder0.value[6]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net123),
    .D(_0074_),
    .Q_N(_0637_),
    .Q(\enc0[6] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder0.value[7]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net124),
    .D(_0075_),
    .Q_N(_0636_),
    .Q(\enc0[7] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder1.old_a$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net125),
    .D(_0076_),
    .Q_N(_0635_),
    .Q(\rgb_mixer.encoder1.old_a ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder1.old_b$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net126),
    .D(_0077_),
    .Q_N(_0634_),
    .Q(\rgb_mixer.encoder1.old_b ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder1.value[0]$_SDFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net127),
    .D(_0078_),
    .Q_N(_0010_),
    .Q(\enc1[0] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder1.value[1]$_SDFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net128),
    .D(_0079_),
    .Q_N(_0633_),
    .Q(\enc1[1] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder1.value[2]$_SDFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net129),
    .D(_0080_),
    .Q_N(_0002_),
    .Q(\enc1[2] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder1.value[3]$_SDFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net130),
    .D(_0081_),
    .Q_N(_0003_),
    .Q(\enc1[3] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder1.value[4]$_SDFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net131),
    .D(_0082_),
    .Q_N(_0632_),
    .Q(\enc1[4] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder1.value[5]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net132),
    .D(_0083_),
    .Q_N(_0631_),
    .Q(\enc1[5] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder1.value[6]$_SDFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net133),
    .D(_0084_),
    .Q_N(_0630_),
    .Q(\enc1[6] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder1.value[7]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net134),
    .D(_0085_),
    .Q_N(_0629_),
    .Q(\enc1[7] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder2.old_a$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net135),
    .D(_0086_),
    .Q_N(_0628_),
    .Q(\rgb_mixer.encoder2.old_a ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder2.old_b$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net136),
    .D(_0087_),
    .Q_N(_0627_),
    .Q(\rgb_mixer.encoder2.old_b ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder2.value[0]$_SDFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net137),
    .D(_0088_),
    .Q_N(_0011_),
    .Q(\enc2[0] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder2.value[1]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net138),
    .D(_0089_),
    .Q_N(_0626_),
    .Q(\enc2[1] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder2.value[2]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net139),
    .D(_0090_),
    .Q_N(_0000_),
    .Q(\enc2[2] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder2.value[3]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net140),
    .D(_0091_),
    .Q_N(_0001_),
    .Q(\enc2[3] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder2.value[4]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net141),
    .D(_0092_),
    .Q_N(_0625_),
    .Q(\enc2[4] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder2.value[5]$_SDFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net142),
    .D(_0093_),
    .Q_N(_0624_),
    .Q(\enc2[5] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder2.value[6]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net143),
    .D(_0094_),
    .Q_N(_0623_),
    .Q(\enc2[6] ));
 sg13g2_dfrbp_1 \rgb_mixer.encoder2.value[7]$_SDFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net144),
    .D(_0095_),
    .Q_N(_0622_),
    .Q(\enc2[7] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm0.count[0]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net145),
    .D(_0096_),
    .Q_N(_0008_),
    .Q(\rgb_mixer.pwm0.count[0] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm0.count[1]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net146),
    .D(_0097_),
    .Q_N(_0621_),
    .Q(\rgb_mixer.pwm0.count[1] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm0.count[2]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net147),
    .D(_0098_),
    .Q_N(_0620_),
    .Q(\rgb_mixer.pwm0.count[2] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm0.count[3]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net148),
    .D(_0099_),
    .Q_N(_0619_),
    .Q(\rgb_mixer.pwm0.count[3] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm0.count[4]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net149),
    .D(_0100_),
    .Q_N(_0618_),
    .Q(\rgb_mixer.pwm0.count[4] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm0.count[5]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net150),
    .D(_0101_),
    .Q_N(_0617_),
    .Q(\rgb_mixer.pwm0.count[5] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm0.count[6]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net151),
    .D(_0102_),
    .Q_N(_0616_),
    .Q(\rgb_mixer.pwm0.count[6] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm0.count[7]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net152),
    .D(_0103_),
    .Q_N(_0615_),
    .Q(\rgb_mixer.pwm0.count[7] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm0.out$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net153),
    .D(_0104_),
    .Q_N(_0614_),
    .Q(\rgb_mixer.pwm0.out ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm1.count[0]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net154),
    .D(_0105_),
    .Q_N(_0007_),
    .Q(\rgb_mixer.pwm1.count[0] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm1.count[1]$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net155),
    .D(_0106_),
    .Q_N(_0613_),
    .Q(\rgb_mixer.pwm1.count[1] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm1.count[2]$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net156),
    .D(_0107_),
    .Q_N(_0612_),
    .Q(\rgb_mixer.pwm1.count[2] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm1.count[3]$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net157),
    .D(_0108_),
    .Q_N(_0611_),
    .Q(\rgb_mixer.pwm1.count[3] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm1.count[4]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net158),
    .D(_0109_),
    .Q_N(_0610_),
    .Q(\rgb_mixer.pwm1.count[4] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm1.count[5]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net159),
    .D(_0110_),
    .Q_N(_0609_),
    .Q(\rgb_mixer.pwm1.count[5] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm1.count[6]$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net160),
    .D(_0111_),
    .Q_N(_0608_),
    .Q(\rgb_mixer.pwm1.count[6] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm1.count[7]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net161),
    .D(_0112_),
    .Q_N(_0607_),
    .Q(\rgb_mixer.pwm1.count[7] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm1.out$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net162),
    .D(_0113_),
    .Q_N(_0606_),
    .Q(\rgb_mixer.pwm1.out ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm2.count[0]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net163),
    .D(_0114_),
    .Q_N(_0006_),
    .Q(\rgb_mixer.pwm2.count[0] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm2.count[1]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net164),
    .D(_0115_),
    .Q_N(_0605_),
    .Q(\rgb_mixer.pwm2.count[1] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm2.count[2]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net165),
    .D(_0116_),
    .Q_N(_0604_),
    .Q(\rgb_mixer.pwm2.count[2] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm2.count[3]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net166),
    .D(_0117_),
    .Q_N(_0603_),
    .Q(\rgb_mixer.pwm2.count[3] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm2.count[4]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net167),
    .D(_0118_),
    .Q_N(_0602_),
    .Q(\rgb_mixer.pwm2.count[4] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm2.count[5]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net168),
    .D(_0119_),
    .Q_N(_0601_),
    .Q(\rgb_mixer.pwm2.count[5] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm2.count[6]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net169),
    .D(_0120_),
    .Q_N(_0600_),
    .Q(\rgb_mixer.pwm2.count[6] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm2.count[7]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net170),
    .D(_0121_),
    .Q_N(_0599_),
    .Q(\rgb_mixer.pwm2.count[7] ));
 sg13g2_dfrbp_1 \rgb_mixer.pwm2.out$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net171),
    .D(_0122_),
    .Q_N(_0598_),
    .Q(\rgb_mixer.pwm2.out ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[0]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[1]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[2]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[3]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[4]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[5]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[6]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[7]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[0]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[1]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[2]));
 sg13g2_buf_2 fanout18 (.A(_0373_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0294_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0465_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0200_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0192_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0191_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0144_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0135_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0134_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0126_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0159_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0125_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0571_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0415_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0393_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0390_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0367_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0362_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0314_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0256_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0235_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0217_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0215_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0201_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0193_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0176_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0170_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0138_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0124_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0569_),
    .X(net47));
 sg13g2_tielo _1306__48 (.L_LO(net48));
 sg13g2_tielo _1307__49 (.L_LO(net49));
 sg13g2_tielo _1308__50 (.L_LO(net50));
 sg13g2_tielo _1309__51 (.L_LO(net51));
 sg13g2_tielo _1310__52 (.L_LO(net52));
 sg13g2_tiehi _1296__54 (.L_HI(net54));
 sg13g2_tiehi _1297__55 (.L_HI(net55));
 sg13g2_tiehi _1298__56 (.L_HI(net56));
 sg13g2_tiehi _1299__57 (.L_HI(net57));
 sg13g2_tiehi _1300__58 (.L_HI(net58));
 sg13g2_tiehi _1301__59 (.L_HI(net59));
 sg13g2_tiehi _1302__60 (.L_HI(net60));
 sg13g2_tiehi \rgb_mixer.debounce0_a.button_hist[0]$_SDFF_PN0__61  (.L_HI(net61));
 sg13g2_tiehi \rgb_mixer.debounce0_a.button_hist[1]$_SDFF_PN0__62  (.L_HI(net62));
 sg13g2_tiehi \rgb_mixer.debounce0_a.button_hist[2]$_SDFF_PN0__63  (.L_HI(net63));
 sg13g2_tiehi \rgb_mixer.debounce0_a.button_hist[3]$_SDFF_PN0__64  (.L_HI(net64));
 sg13g2_tiehi \rgb_mixer.debounce0_a.button_hist[4]$_SDFF_PN0__65  (.L_HI(net65));
 sg13g2_tiehi \rgb_mixer.debounce0_a.button_hist[5]$_SDFF_PN0__66  (.L_HI(net66));
 sg13g2_tiehi \rgb_mixer.debounce0_a.button_hist[6]$_SDFF_PN0__67  (.L_HI(net67));
 sg13g2_tiehi \rgb_mixer.debounce0_a.button_hist[7]$_SDFF_PN0__68  (.L_HI(net68));
 sg13g2_tiehi \rgb_mixer.debounce0_a.debounced$_SDFFE_PN0P__69  (.L_HI(net69));
 sg13g2_tiehi \rgb_mixer.debounce0_b.button_hist[0]$_SDFF_PN0__70  (.L_HI(net70));
 sg13g2_tiehi \rgb_mixer.debounce0_b.button_hist[1]$_SDFF_PN0__71  (.L_HI(net71));
 sg13g2_tiehi \rgb_mixer.debounce0_b.button_hist[2]$_SDFF_PN0__72  (.L_HI(net72));
 sg13g2_tiehi \rgb_mixer.debounce0_b.button_hist[3]$_SDFF_PN0__73  (.L_HI(net73));
 sg13g2_tiehi \rgb_mixer.debounce0_b.button_hist[4]$_SDFF_PN0__74  (.L_HI(net74));
 sg13g2_tiehi \rgb_mixer.debounce0_b.button_hist[5]$_SDFF_PN0__75  (.L_HI(net75));
 sg13g2_tiehi \rgb_mixer.debounce0_b.button_hist[6]$_SDFF_PN0__76  (.L_HI(net76));
 sg13g2_tiehi \rgb_mixer.debounce0_b.button_hist[7]$_SDFF_PN0__77  (.L_HI(net77));
 sg13g2_tiehi \rgb_mixer.debounce0_b.debounced$_SDFFE_PN0P__78  (.L_HI(net78));
 sg13g2_tiehi \rgb_mixer.debounce1_a.button_hist[0]$_SDFF_PN0__79  (.L_HI(net79));
 sg13g2_tiehi \rgb_mixer.debounce1_a.button_hist[1]$_SDFF_PN0__80  (.L_HI(net80));
 sg13g2_tiehi \rgb_mixer.debounce1_a.button_hist[2]$_SDFF_PN0__81  (.L_HI(net81));
 sg13g2_tiehi \rgb_mixer.debounce1_a.button_hist[3]$_SDFF_PN0__82  (.L_HI(net82));
 sg13g2_tiehi \rgb_mixer.debounce1_a.button_hist[4]$_SDFF_PN0__83  (.L_HI(net83));
 sg13g2_tiehi \rgb_mixer.debounce1_a.button_hist[5]$_SDFF_PN0__84  (.L_HI(net84));
 sg13g2_tiehi \rgb_mixer.debounce1_a.button_hist[6]$_SDFF_PN0__85  (.L_HI(net85));
 sg13g2_tiehi \rgb_mixer.debounce1_a.button_hist[7]$_SDFF_PN0__86  (.L_HI(net86));
 sg13g2_tiehi \rgb_mixer.debounce1_a.debounced$_SDFFE_PN0P__87  (.L_HI(net87));
 sg13g2_tiehi \rgb_mixer.debounce1_b.button_hist[0]$_SDFF_PN0__88  (.L_HI(net88));
 sg13g2_tiehi \rgb_mixer.debounce1_b.button_hist[1]$_SDFF_PN0__89  (.L_HI(net89));
 sg13g2_tiehi \rgb_mixer.debounce1_b.button_hist[2]$_SDFF_PN0__90  (.L_HI(net90));
 sg13g2_tiehi \rgb_mixer.debounce1_b.button_hist[3]$_SDFF_PN0__91  (.L_HI(net91));
 sg13g2_tiehi \rgb_mixer.debounce1_b.button_hist[4]$_SDFF_PN0__92  (.L_HI(net92));
 sg13g2_tiehi \rgb_mixer.debounce1_b.button_hist[5]$_SDFF_PN0__93  (.L_HI(net93));
 sg13g2_tiehi \rgb_mixer.debounce1_b.button_hist[6]$_SDFF_PN0__94  (.L_HI(net94));
 sg13g2_tiehi \rgb_mixer.debounce1_b.button_hist[7]$_SDFF_PN0__95  (.L_HI(net95));
 sg13g2_tiehi \rgb_mixer.debounce1_b.debounced$_SDFFE_PN0P__96  (.L_HI(net96));
 sg13g2_tiehi \rgb_mixer.debounce2_a.button_hist[0]$_SDFF_PN0__97  (.L_HI(net97));
 sg13g2_tiehi \rgb_mixer.debounce2_a.button_hist[1]$_SDFF_PN0__98  (.L_HI(net98));
 sg13g2_tiehi \rgb_mixer.debounce2_a.button_hist[2]$_SDFF_PN0__99  (.L_HI(net99));
 sg13g2_tiehi \rgb_mixer.debounce2_a.button_hist[3]$_SDFF_PN0__100  (.L_HI(net100));
 sg13g2_tiehi \rgb_mixer.debounce2_a.button_hist[4]$_SDFF_PN0__101  (.L_HI(net101));
 sg13g2_tiehi \rgb_mixer.debounce2_a.button_hist[5]$_SDFF_PN0__102  (.L_HI(net102));
 sg13g2_tiehi \rgb_mixer.debounce2_a.button_hist[6]$_SDFF_PN0__103  (.L_HI(net103));
 sg13g2_tiehi \rgb_mixer.debounce2_a.button_hist[7]$_SDFF_PN0__104  (.L_HI(net104));
 sg13g2_tiehi \rgb_mixer.debounce2_a.debounced$_SDFFE_PN0P__105  (.L_HI(net105));
 sg13g2_tiehi \rgb_mixer.debounce2_b.button_hist[0]$_SDFF_PN0__106  (.L_HI(net106));
 sg13g2_tiehi \rgb_mixer.debounce2_b.button_hist[1]$_SDFF_PN0__107  (.L_HI(net107));
 sg13g2_tiehi \rgb_mixer.debounce2_b.button_hist[2]$_SDFF_PN0__108  (.L_HI(net108));
 sg13g2_tiehi \rgb_mixer.debounce2_b.button_hist[3]$_SDFF_PN0__109  (.L_HI(net109));
 sg13g2_tiehi \rgb_mixer.debounce2_b.button_hist[4]$_SDFF_PN0__110  (.L_HI(net110));
 sg13g2_tiehi \rgb_mixer.debounce2_b.button_hist[5]$_SDFF_PN0__111  (.L_HI(net111));
 sg13g2_tiehi \rgb_mixer.debounce2_b.button_hist[6]$_SDFF_PN0__112  (.L_HI(net112));
 sg13g2_tiehi \rgb_mixer.debounce2_b.button_hist[7]$_SDFF_PN0__113  (.L_HI(net113));
 sg13g2_tiehi \rgb_mixer.debounce2_b.debounced$_SDFFE_PN0P__114  (.L_HI(net114));
 sg13g2_tiehi \rgb_mixer.encoder0.old_a$_SDFF_PN0__115  (.L_HI(net115));
 sg13g2_tiehi \rgb_mixer.encoder0.old_b$_SDFF_PN0__116  (.L_HI(net116));
 sg13g2_tiehi \rgb_mixer.encoder0.value[0]$_SDFFE_PN0P__117  (.L_HI(net117));
 sg13g2_tiehi \rgb_mixer.encoder0.value[1]$_SDFFE_PN0P__118  (.L_HI(net118));
 sg13g2_tiehi \rgb_mixer.encoder0.value[2]$_SDFFE_PN0P__119  (.L_HI(net119));
 sg13g2_tiehi \rgb_mixer.encoder0.value[3]$_SDFFE_PN0P__120  (.L_HI(net120));
 sg13g2_tiehi \rgb_mixer.encoder0.value[4]$_SDFFE_PN0P__121  (.L_HI(net121));
 sg13g2_tiehi \rgb_mixer.encoder0.value[5]$_SDFFE_PN0P__122  (.L_HI(net122));
 sg13g2_tiehi \rgb_mixer.encoder0.value[6]$_SDFFE_PN0P__123  (.L_HI(net123));
 sg13g2_tiehi \rgb_mixer.encoder0.value[7]$_SDFFE_PN0P__124  (.L_HI(net124));
 sg13g2_tiehi \rgb_mixer.encoder1.old_a$_SDFF_PN0__125  (.L_HI(net125));
 sg13g2_tiehi \rgb_mixer.encoder1.old_b$_SDFF_PN0__126  (.L_HI(net126));
 sg13g2_tiehi \rgb_mixer.encoder1.value[0]$_SDFFE_PN0P__127  (.L_HI(net127));
 sg13g2_tiehi \rgb_mixer.encoder1.value[1]$_SDFFE_PN0P__128  (.L_HI(net128));
 sg13g2_tiehi \rgb_mixer.encoder1.value[2]$_SDFFE_PN0P__129  (.L_HI(net129));
 sg13g2_tiehi \rgb_mixer.encoder1.value[3]$_SDFFE_PN0P__130  (.L_HI(net130));
 sg13g2_tiehi \rgb_mixer.encoder1.value[4]$_SDFFE_PN0P__131  (.L_HI(net131));
 sg13g2_tiehi \rgb_mixer.encoder1.value[5]$_SDFFE_PN0P__132  (.L_HI(net132));
 sg13g2_tiehi \rgb_mixer.encoder1.value[6]$_SDFFE_PN0P__133  (.L_HI(net133));
 sg13g2_tiehi \rgb_mixer.encoder1.value[7]$_SDFFE_PN0P__134  (.L_HI(net134));
 sg13g2_tiehi \rgb_mixer.encoder2.old_a$_SDFF_PN0__135  (.L_HI(net135));
 sg13g2_tiehi \rgb_mixer.encoder2.old_b$_SDFF_PN0__136  (.L_HI(net136));
 sg13g2_tiehi \rgb_mixer.encoder2.value[0]$_SDFFE_PN0P__137  (.L_HI(net137));
 sg13g2_tiehi \rgb_mixer.encoder2.value[1]$_SDFFE_PN0P__138  (.L_HI(net138));
 sg13g2_tiehi \rgb_mixer.encoder2.value[2]$_SDFFE_PN0P__139  (.L_HI(net139));
 sg13g2_tiehi \rgb_mixer.encoder2.value[3]$_SDFFE_PN0P__140  (.L_HI(net140));
 sg13g2_tiehi \rgb_mixer.encoder2.value[4]$_SDFFE_PN0P__141  (.L_HI(net141));
 sg13g2_tiehi \rgb_mixer.encoder2.value[5]$_SDFFE_PN0P__142  (.L_HI(net142));
 sg13g2_tiehi \rgb_mixer.encoder2.value[6]$_SDFFE_PN0P__143  (.L_HI(net143));
 sg13g2_tiehi \rgb_mixer.encoder2.value[7]$_SDFFE_PN0P__144  (.L_HI(net144));
 sg13g2_tiehi \rgb_mixer.pwm0.count[0]$_SDFF_PN0__145  (.L_HI(net145));
 sg13g2_tiehi \rgb_mixer.pwm0.count[1]$_SDFF_PN0__146  (.L_HI(net146));
 sg13g2_tiehi \rgb_mixer.pwm0.count[2]$_SDFF_PN0__147  (.L_HI(net147));
 sg13g2_tiehi \rgb_mixer.pwm0.count[3]$_SDFF_PN0__148  (.L_HI(net148));
 sg13g2_tiehi \rgb_mixer.pwm0.count[4]$_SDFF_PN0__149  (.L_HI(net149));
 sg13g2_tiehi \rgb_mixer.pwm0.count[5]$_SDFF_PN0__150  (.L_HI(net150));
 sg13g2_tiehi \rgb_mixer.pwm0.count[6]$_SDFF_PN0__151  (.L_HI(net151));
 sg13g2_tiehi \rgb_mixer.pwm0.count[7]$_SDFF_PN0__152  (.L_HI(net152));
 sg13g2_tiehi \rgb_mixer.pwm0.out$_SDFF_PN0__153  (.L_HI(net153));
 sg13g2_tiehi \rgb_mixer.pwm1.count[0]$_SDFF_PN0__154  (.L_HI(net154));
 sg13g2_tiehi \rgb_mixer.pwm1.count[1]$_SDFF_PN0__155  (.L_HI(net155));
 sg13g2_tiehi \rgb_mixer.pwm1.count[2]$_SDFF_PN0__156  (.L_HI(net156));
 sg13g2_tiehi \rgb_mixer.pwm1.count[3]$_SDFF_PN0__157  (.L_HI(net157));
 sg13g2_tiehi \rgb_mixer.pwm1.count[4]$_SDFF_PN0__158  (.L_HI(net158));
 sg13g2_tiehi \rgb_mixer.pwm1.count[5]$_SDFF_PN0__159  (.L_HI(net159));
 sg13g2_tiehi \rgb_mixer.pwm1.count[6]$_SDFF_PN0__160  (.L_HI(net160));
 sg13g2_tiehi \rgb_mixer.pwm1.count[7]$_SDFF_PN0__161  (.L_HI(net161));
 sg13g2_tiehi \rgb_mixer.pwm1.out$_SDFF_PN0__162  (.L_HI(net162));
 sg13g2_tiehi \rgb_mixer.pwm2.count[0]$_SDFF_PN0__163  (.L_HI(net163));
 sg13g2_tiehi \rgb_mixer.pwm2.count[1]$_SDFF_PN0__164  (.L_HI(net164));
 sg13g2_tiehi \rgb_mixer.pwm2.count[2]$_SDFF_PN0__165  (.L_HI(net165));
 sg13g2_tiehi \rgb_mixer.pwm2.count[3]$_SDFF_PN0__166  (.L_HI(net166));
 sg13g2_tiehi \rgb_mixer.pwm2.count[4]$_SDFF_PN0__167  (.L_HI(net167));
 sg13g2_tiehi \rgb_mixer.pwm2.count[5]$_SDFF_PN0__168  (.L_HI(net168));
 sg13g2_tiehi \rgb_mixer.pwm2.count[6]$_SDFF_PN0__169  (.L_HI(net169));
 sg13g2_tiehi \rgb_mixer.pwm2.count[7]$_SDFF_PN0__170  (.L_HI(net170));
 sg13g2_tiehi \rgb_mixer.pwm2.out$_SDFF_PN0__171  (.L_HI(net171));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_4 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_134 ();
 sg13g2_decap_8 FILLER_13_141 ();
 sg13g2_decap_8 FILLER_13_148 ();
 sg13g2_decap_8 FILLER_13_155 ();
 sg13g2_decap_8 FILLER_13_162 ();
 sg13g2_decap_8 FILLER_13_169 ();
 sg13g2_decap_8 FILLER_13_176 ();
 sg13g2_decap_8 FILLER_13_183 ();
 sg13g2_decap_8 FILLER_13_190 ();
 sg13g2_decap_8 FILLER_13_197 ();
 sg13g2_decap_8 FILLER_13_204 ();
 sg13g2_decap_8 FILLER_13_211 ();
 sg13g2_decap_8 FILLER_13_218 ();
 sg13g2_decap_8 FILLER_13_225 ();
 sg13g2_decap_8 FILLER_13_232 ();
 sg13g2_decap_8 FILLER_13_239 ();
 sg13g2_decap_8 FILLER_13_246 ();
 sg13g2_decap_8 FILLER_13_253 ();
 sg13g2_decap_8 FILLER_13_260 ();
 sg13g2_decap_8 FILLER_13_267 ();
 sg13g2_decap_8 FILLER_13_274 ();
 sg13g2_decap_8 FILLER_13_281 ();
 sg13g2_decap_8 FILLER_13_288 ();
 sg13g2_fill_2 FILLER_13_295 ();
 sg13g2_fill_1 FILLER_13_297 ();
 sg13g2_decap_8 FILLER_13_303 ();
 sg13g2_decap_8 FILLER_13_310 ();
 sg13g2_decap_8 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_324 ();
 sg13g2_decap_8 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_338 ();
 sg13g2_decap_8 FILLER_13_345 ();
 sg13g2_decap_8 FILLER_13_352 ();
 sg13g2_decap_8 FILLER_13_359 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_decap_8 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_13_415 ();
 sg13g2_decap_8 FILLER_13_422 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_4 FILLER_14_77 ();
 sg13g2_fill_2 FILLER_14_81 ();
 sg13g2_fill_1 FILLER_14_87 ();
 sg13g2_decap_4 FILLER_14_114 ();
 sg13g2_fill_1 FILLER_14_118 ();
 sg13g2_fill_1 FILLER_14_149 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_decap_4 FILLER_14_165 ();
 sg13g2_fill_2 FILLER_14_169 ();
 sg13g2_fill_2 FILLER_14_180 ();
 sg13g2_decap_8 FILLER_14_192 ();
 sg13g2_decap_8 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_decap_4 FILLER_14_213 ();
 sg13g2_decap_8 FILLER_14_247 ();
 sg13g2_decap_8 FILLER_14_254 ();
 sg13g2_decap_8 FILLER_14_261 ();
 sg13g2_decap_4 FILLER_14_268 ();
 sg13g2_fill_2 FILLER_14_272 ();
 sg13g2_fill_1 FILLER_14_300 ();
 sg13g2_decap_8 FILLER_14_327 ();
 sg13g2_fill_1 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_339 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_decap_8 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_decap_8 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_14_409 ();
 sg13g2_decap_8 FILLER_14_416 ();
 sg13g2_decap_8 FILLER_14_423 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_49 ();
 sg13g2_fill_1 FILLER_15_76 ();
 sg13g2_fill_1 FILLER_15_82 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_120 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_decap_4 FILLER_15_134 ();
 sg13g2_fill_1 FILLER_15_179 ();
 sg13g2_fill_1 FILLER_15_194 ();
 sg13g2_decap_4 FILLER_15_203 ();
 sg13g2_fill_1 FILLER_15_207 ();
 sg13g2_decap_4 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_226 ();
 sg13g2_decap_8 FILLER_15_233 ();
 sg13g2_decap_8 FILLER_15_240 ();
 sg13g2_decap_4 FILLER_15_247 ();
 sg13g2_fill_1 FILLER_15_251 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_300 ();
 sg13g2_fill_1 FILLER_15_307 ();
 sg13g2_decap_8 FILLER_15_312 ();
 sg13g2_decap_4 FILLER_15_319 ();
 sg13g2_fill_2 FILLER_15_354 ();
 sg13g2_fill_1 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_4 FILLER_16_60 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_fill_2 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_97 ();
 sg13g2_fill_2 FILLER_16_120 ();
 sg13g2_fill_1 FILLER_16_147 ();
 sg13g2_decap_4 FILLER_16_153 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_fill_1 FILLER_16_184 ();
 sg13g2_fill_1 FILLER_16_188 ();
 sg13g2_fill_1 FILLER_16_206 ();
 sg13g2_fill_1 FILLER_16_212 ();
 sg13g2_fill_2 FILLER_16_218 ();
 sg13g2_decap_4 FILLER_16_254 ();
 sg13g2_fill_2 FILLER_16_258 ();
 sg13g2_decap_8 FILLER_16_264 ();
 sg13g2_fill_2 FILLER_16_271 ();
 sg13g2_decap_4 FILLER_16_301 ();
 sg13g2_fill_1 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_344 ();
 sg13g2_decap_4 FILLER_16_355 ();
 sg13g2_fill_1 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_fill_2 FILLER_16_376 ();
 sg13g2_fill_1 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_16_412 ();
 sg13g2_decap_8 FILLER_16_419 ();
 sg13g2_decap_4 FILLER_16_426 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_fill_2 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_58 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_fill_1 FILLER_17_70 ();
 sg13g2_decap_4 FILLER_17_83 ();
 sg13g2_fill_2 FILLER_17_87 ();
 sg13g2_decap_8 FILLER_17_109 ();
 sg13g2_decap_8 FILLER_17_116 ();
 sg13g2_decap_8 FILLER_17_123 ();
 sg13g2_decap_4 FILLER_17_146 ();
 sg13g2_fill_1 FILLER_17_179 ();
 sg13g2_fill_2 FILLER_17_185 ();
 sg13g2_decap_8 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_216 ();
 sg13g2_fill_1 FILLER_17_223 ();
 sg13g2_decap_4 FILLER_17_229 ();
 sg13g2_fill_2 FILLER_17_233 ();
 sg13g2_decap_4 FILLER_17_239 ();
 sg13g2_fill_1 FILLER_17_243 ();
 sg13g2_fill_2 FILLER_17_270 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_decap_8 FILLER_17_276 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_fill_1 FILLER_17_290 ();
 sg13g2_decap_4 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_decap_4 FILLER_17_315 ();
 sg13g2_fill_1 FILLER_17_319 ();
 sg13g2_fill_2 FILLER_17_324 ();
 sg13g2_fill_2 FILLER_17_336 ();
 sg13g2_decap_4 FILLER_17_369 ();
 sg13g2_fill_2 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_17_414 ();
 sg13g2_decap_8 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_4 FILLER_18_28 ();
 sg13g2_fill_2 FILLER_18_58 ();
 sg13g2_fill_2 FILLER_18_64 ();
 sg13g2_fill_2 FILLER_18_74 ();
 sg13g2_fill_1 FILLER_18_76 ();
 sg13g2_fill_1 FILLER_18_116 ();
 sg13g2_fill_1 FILLER_18_121 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_4 FILLER_18_133 ();
 sg13g2_fill_2 FILLER_18_153 ();
 sg13g2_fill_2 FILLER_18_159 ();
 sg13g2_fill_1 FILLER_18_161 ();
 sg13g2_fill_1 FILLER_18_167 ();
 sg13g2_decap_8 FILLER_18_173 ();
 sg13g2_decap_8 FILLER_18_180 ();
 sg13g2_decap_8 FILLER_18_187 ();
 sg13g2_decap_8 FILLER_18_194 ();
 sg13g2_decap_8 FILLER_18_205 ();
 sg13g2_decap_8 FILLER_18_212 ();
 sg13g2_decap_8 FILLER_18_219 ();
 sg13g2_decap_8 FILLER_18_226 ();
 sg13g2_fill_2 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_239 ();
 sg13g2_decap_4 FILLER_18_246 ();
 sg13g2_decap_8 FILLER_18_254 ();
 sg13g2_fill_2 FILLER_18_261 ();
 sg13g2_fill_1 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_fill_1 FILLER_18_361 ();
 sg13g2_fill_2 FILLER_18_369 ();
 sg13g2_fill_1 FILLER_18_371 ();
 sg13g2_fill_2 FILLER_18_397 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_4 FILLER_19_21 ();
 sg13g2_fill_1 FILLER_19_25 ();
 sg13g2_decap_8 FILLER_19_31 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_4 FILLER_19_63 ();
 sg13g2_fill_1 FILLER_19_79 ();
 sg13g2_decap_8 FILLER_19_85 ();
 sg13g2_decap_8 FILLER_19_92 ();
 sg13g2_decap_4 FILLER_19_99 ();
 sg13g2_decap_4 FILLER_19_113 ();
 sg13g2_fill_1 FILLER_19_131 ();
 sg13g2_fill_2 FILLER_19_141 ();
 sg13g2_decap_8 FILLER_19_148 ();
 sg13g2_fill_2 FILLER_19_155 ();
 sg13g2_decap_4 FILLER_19_162 ();
 sg13g2_fill_1 FILLER_19_166 ();
 sg13g2_decap_8 FILLER_19_171 ();
 sg13g2_decap_8 FILLER_19_178 ();
 sg13g2_decap_4 FILLER_19_185 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_decap_4 FILLER_19_220 ();
 sg13g2_decap_8 FILLER_19_254 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_decap_8 FILLER_19_268 ();
 sg13g2_fill_2 FILLER_19_275 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_fill_2 FILLER_19_315 ();
 sg13g2_decap_4 FILLER_19_321 ();
 sg13g2_fill_2 FILLER_19_325 ();
 sg13g2_decap_4 FILLER_19_331 ();
 sg13g2_decap_4 FILLER_19_339 ();
 sg13g2_decap_4 FILLER_19_384 ();
 sg13g2_fill_2 FILLER_19_388 ();
 sg13g2_fill_1 FILLER_19_395 ();
 sg13g2_fill_2 FILLER_19_422 ();
 sg13g2_fill_1 FILLER_19_424 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_11 ();
 sg13g2_fill_2 FILLER_20_69 ();
 sg13g2_fill_1 FILLER_20_71 ();
 sg13g2_fill_1 FILLER_20_82 ();
 sg13g2_decap_4 FILLER_20_109 ();
 sg13g2_fill_2 FILLER_20_113 ();
 sg13g2_decap_8 FILLER_20_118 ();
 sg13g2_decap_8 FILLER_20_125 ();
 sg13g2_fill_2 FILLER_20_132 ();
 sg13g2_fill_2 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_155 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_185 ();
 sg13g2_fill_1 FILLER_20_197 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_fill_2 FILLER_20_217 ();
 sg13g2_decap_4 FILLER_20_227 ();
 sg13g2_fill_2 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_245 ();
 sg13g2_decap_4 FILLER_20_250 ();
 sg13g2_fill_2 FILLER_20_254 ();
 sg13g2_decap_8 FILLER_20_292 ();
 sg13g2_decap_4 FILLER_20_299 ();
 sg13g2_fill_1 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_309 ();
 sg13g2_decap_4 FILLER_20_336 ();
 sg13g2_fill_1 FILLER_20_340 ();
 sg13g2_decap_4 FILLER_20_350 ();
 sg13g2_fill_2 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_decap_4 FILLER_20_372 ();
 sg13g2_decap_4 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_4 FILLER_20_396 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_25 ();
 sg13g2_decap_4 FILLER_21_32 ();
 sg13g2_fill_1 FILLER_21_48 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_decap_4 FILLER_21_60 ();
 sg13g2_fill_2 FILLER_21_64 ();
 sg13g2_fill_2 FILLER_21_71 ();
 sg13g2_fill_2 FILLER_21_78 ();
 sg13g2_fill_1 FILLER_21_80 ();
 sg13g2_decap_8 FILLER_21_95 ();
 sg13g2_decap_4 FILLER_21_107 ();
 sg13g2_fill_1 FILLER_21_137 ();
 sg13g2_fill_2 FILLER_21_153 ();
 sg13g2_decap_8 FILLER_21_159 ();
 sg13g2_decap_8 FILLER_21_166 ();
 sg13g2_fill_2 FILLER_21_173 ();
 sg13g2_fill_2 FILLER_21_179 ();
 sg13g2_fill_1 FILLER_21_181 ();
 sg13g2_fill_1 FILLER_21_187 ();
 sg13g2_decap_4 FILLER_21_212 ();
 sg13g2_decap_8 FILLER_21_251 ();
 sg13g2_decap_8 FILLER_21_258 ();
 sg13g2_fill_1 FILLER_21_265 ();
 sg13g2_decap_8 FILLER_21_278 ();
 sg13g2_fill_2 FILLER_21_285 ();
 sg13g2_decap_4 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_313 ();
 sg13g2_fill_2 FILLER_21_319 ();
 sg13g2_fill_1 FILLER_21_347 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_fill_1 FILLER_21_409 ();
 sg13g2_decap_8 FILLER_21_414 ();
 sg13g2_decap_8 FILLER_21_421 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_20 ();
 sg13g2_decap_8 FILLER_22_27 ();
 sg13g2_fill_2 FILLER_22_34 ();
 sg13g2_fill_1 FILLER_22_36 ();
 sg13g2_fill_2 FILLER_22_50 ();
 sg13g2_fill_2 FILLER_22_80 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_decap_4 FILLER_22_101 ();
 sg13g2_fill_1 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_120 ();
 sg13g2_decap_8 FILLER_22_125 ();
 sg13g2_decap_8 FILLER_22_132 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_fill_2 FILLER_22_175 ();
 sg13g2_fill_1 FILLER_22_177 ();
 sg13g2_fill_1 FILLER_22_195 ();
 sg13g2_decap_8 FILLER_22_222 ();
 sg13g2_fill_2 FILLER_22_238 ();
 sg13g2_fill_1 FILLER_22_244 ();
 sg13g2_decap_8 FILLER_22_254 ();
 sg13g2_fill_2 FILLER_22_261 ();
 sg13g2_fill_1 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_268 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_fill_2 FILLER_22_292 ();
 sg13g2_fill_1 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_321 ();
 sg13g2_fill_2 FILLER_22_328 ();
 sg13g2_fill_2 FILLER_22_334 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_4 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_4 FILLER_22_371 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_388 ();
 sg13g2_decap_4 FILLER_22_395 ();
 sg13g2_fill_1 FILLER_22_399 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_fill_1 FILLER_22_409 ();
 sg13g2_decap_8 FILLER_22_414 ();
 sg13g2_decap_8 FILLER_22_421 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_38 ();
 sg13g2_fill_2 FILLER_23_43 ();
 sg13g2_decap_8 FILLER_23_79 ();
 sg13g2_decap_4 FILLER_23_86 ();
 sg13g2_fill_2 FILLER_23_90 ();
 sg13g2_decap_4 FILLER_23_102 ();
 sg13g2_fill_1 FILLER_23_106 ();
 sg13g2_fill_2 FILLER_23_114 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_4 FILLER_23_168 ();
 sg13g2_fill_1 FILLER_23_172 ();
 sg13g2_decap_8 FILLER_23_181 ();
 sg13g2_decap_8 FILLER_23_188 ();
 sg13g2_decap_4 FILLER_23_195 ();
 sg13g2_fill_2 FILLER_23_206 ();
 sg13g2_decap_8 FILLER_23_213 ();
 sg13g2_decap_4 FILLER_23_220 ();
 sg13g2_fill_2 FILLER_23_241 ();
 sg13g2_fill_1 FILLER_23_269 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_4 FILLER_23_287 ();
 sg13g2_fill_1 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_302 ();
 sg13g2_decap_8 FILLER_23_309 ();
 sg13g2_decap_4 FILLER_23_316 ();
 sg13g2_decap_4 FILLER_23_357 ();
 sg13g2_fill_2 FILLER_23_361 ();
 sg13g2_fill_2 FILLER_23_373 ();
 sg13g2_fill_1 FILLER_23_375 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_22 ();
 sg13g2_decap_8 FILLER_24_29 ();
 sg13g2_fill_2 FILLER_24_36 ();
 sg13g2_fill_1 FILLER_24_38 ();
 sg13g2_decap_8 FILLER_24_47 ();
 sg13g2_decap_4 FILLER_24_54 ();
 sg13g2_fill_2 FILLER_24_58 ();
 sg13g2_decap_8 FILLER_24_64 ();
 sg13g2_fill_1 FILLER_24_71 ();
 sg13g2_decap_4 FILLER_24_76 ();
 sg13g2_fill_2 FILLER_24_80 ();
 sg13g2_decap_8 FILLER_24_86 ();
 sg13g2_decap_8 FILLER_24_93 ();
 sg13g2_decap_8 FILLER_24_100 ();
 sg13g2_decap_4 FILLER_24_107 ();
 sg13g2_fill_1 FILLER_24_111 ();
 sg13g2_decap_8 FILLER_24_118 ();
 sg13g2_decap_4 FILLER_24_125 ();
 sg13g2_decap_4 FILLER_24_133 ();
 sg13g2_decap_4 FILLER_24_141 ();
 sg13g2_fill_2 FILLER_24_177 ();
 sg13g2_fill_1 FILLER_24_179 ();
 sg13g2_decap_4 FILLER_24_213 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_fill_2 FILLER_24_228 ();
 sg13g2_decap_4 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_272 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_decap_4 FILLER_24_313 ();
 sg13g2_fill_2 FILLER_24_317 ();
 sg13g2_decap_8 FILLER_24_326 ();
 sg13g2_decap_4 FILLER_24_333 ();
 sg13g2_fill_1 FILLER_24_337 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_349 ();
 sg13g2_decap_4 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_fill_1 FILLER_24_398 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_37 ();
 sg13g2_decap_4 FILLER_25_54 ();
 sg13g2_fill_1 FILLER_25_58 ();
 sg13g2_fill_2 FILLER_25_104 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_fill_2 FILLER_25_133 ();
 sg13g2_fill_1 FILLER_25_139 ();
 sg13g2_fill_1 FILLER_25_145 ();
 sg13g2_fill_2 FILLER_25_150 ();
 sg13g2_fill_2 FILLER_25_156 ();
 sg13g2_fill_2 FILLER_25_166 ();
 sg13g2_fill_1 FILLER_25_168 ();
 sg13g2_decap_4 FILLER_25_173 ();
 sg13g2_fill_2 FILLER_25_177 ();
 sg13g2_fill_2 FILLER_25_183 ();
 sg13g2_fill_1 FILLER_25_185 ();
 sg13g2_decap_4 FILLER_25_190 ();
 sg13g2_fill_2 FILLER_25_194 ();
 sg13g2_fill_1 FILLER_25_206 ();
 sg13g2_decap_8 FILLER_25_213 ();
 sg13g2_decap_8 FILLER_25_220 ();
 sg13g2_fill_1 FILLER_25_227 ();
 sg13g2_fill_1 FILLER_25_236 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_249 ();
 sg13g2_fill_1 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_263 ();
 sg13g2_fill_1 FILLER_25_267 ();
 sg13g2_fill_1 FILLER_25_272 ();
 sg13g2_decap_8 FILLER_25_283 ();
 sg13g2_decap_4 FILLER_25_290 ();
 sg13g2_fill_2 FILLER_25_294 ();
 sg13g2_fill_2 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_331 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_fill_2 FILLER_25_350 ();
 sg13g2_fill_1 FILLER_25_352 ();
 sg13g2_decap_4 FILLER_25_357 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_fill_1 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_405 ();
 sg13g2_fill_1 FILLER_25_412 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_4 FILLER_25_424 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_25 ();
 sg13g2_fill_2 FILLER_26_31 ();
 sg13g2_fill_1 FILLER_26_33 ();
 sg13g2_decap_4 FILLER_26_64 ();
 sg13g2_fill_1 FILLER_26_68 ();
 sg13g2_decap_8 FILLER_26_74 ();
 sg13g2_decap_4 FILLER_26_81 ();
 sg13g2_fill_1 FILLER_26_85 ();
 sg13g2_decap_4 FILLER_26_95 ();
 sg13g2_decap_4 FILLER_26_104 ();
 sg13g2_decap_4 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_fill_1 FILLER_26_170 ();
 sg13g2_decap_8 FILLER_26_186 ();
 sg13g2_decap_4 FILLER_26_193 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_209 ();
 sg13g2_decap_8 FILLER_26_220 ();
 sg13g2_decap_4 FILLER_26_227 ();
 sg13g2_fill_1 FILLER_26_231 ();
 sg13g2_decap_4 FILLER_26_236 ();
 sg13g2_fill_1 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_decap_4 FILLER_26_263 ();
 sg13g2_fill_2 FILLER_26_272 ();
 sg13g2_fill_1 FILLER_26_274 ();
 sg13g2_fill_2 FILLER_26_305 ();
 sg13g2_fill_1 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_330 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_fill_2 FILLER_26_344 ();
 sg13g2_fill_2 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_4 FILLER_26_390 ();
 sg13g2_decap_4 FILLER_26_425 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_11 ();
 sg13g2_decap_4 FILLER_27_39 ();
 sg13g2_fill_2 FILLER_27_43 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_67 ();
 sg13g2_fill_2 FILLER_27_116 ();
 sg13g2_decap_8 FILLER_27_123 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_decap_4 FILLER_27_135 ();
 sg13g2_fill_2 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_149 ();
 sg13g2_fill_2 FILLER_27_158 ();
 sg13g2_fill_1 FILLER_27_160 ();
 sg13g2_decap_8 FILLER_27_169 ();
 sg13g2_fill_2 FILLER_27_176 ();
 sg13g2_fill_2 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_234 ();
 sg13g2_decap_4 FILLER_27_246 ();
 sg13g2_fill_1 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_268 ();
 sg13g2_decap_4 FILLER_27_276 ();
 sg13g2_fill_1 FILLER_27_280 ();
 sg13g2_fill_2 FILLER_27_286 ();
 sg13g2_fill_2 FILLER_27_317 ();
 sg13g2_decap_8 FILLER_27_331 ();
 sg13g2_decap_8 FILLER_27_338 ();
 sg13g2_decap_8 FILLER_27_345 ();
 sg13g2_fill_2 FILLER_27_352 ();
 sg13g2_fill_1 FILLER_27_354 ();
 sg13g2_fill_2 FILLER_27_381 ();
 sg13g2_fill_2 FILLER_27_388 ();
 sg13g2_fill_1 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_27_421 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_4 FILLER_28_25 ();
 sg13g2_decap_8 FILLER_28_33 ();
 sg13g2_decap_8 FILLER_28_40 ();
 sg13g2_decap_8 FILLER_28_81 ();
 sg13g2_decap_8 FILLER_28_88 ();
 sg13g2_decap_8 FILLER_28_95 ();
 sg13g2_decap_8 FILLER_28_102 ();
 sg13g2_fill_2 FILLER_28_109 ();
 sg13g2_decap_8 FILLER_28_116 ();
 sg13g2_fill_1 FILLER_28_149 ();
 sg13g2_decap_4 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_fill_1 FILLER_28_197 ();
 sg13g2_fill_1 FILLER_28_202 ();
 sg13g2_decap_4 FILLER_28_208 ();
 sg13g2_fill_2 FILLER_28_212 ();
 sg13g2_decap_8 FILLER_28_244 ();
 sg13g2_decap_8 FILLER_28_251 ();
 sg13g2_decap_8 FILLER_28_258 ();
 sg13g2_decap_8 FILLER_28_265 ();
 sg13g2_decap_4 FILLER_28_272 ();
 sg13g2_decap_4 FILLER_28_290 ();
 sg13g2_fill_1 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_299 ();
 sg13g2_fill_2 FILLER_28_314 ();
 sg13g2_fill_2 FILLER_28_319 ();
 sg13g2_decap_8 FILLER_28_356 ();
 sg13g2_fill_2 FILLER_28_383 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_4 FILLER_28_396 ();
 sg13g2_fill_1 FILLER_28_405 ();
 sg13g2_fill_1 FILLER_28_410 ();
 sg13g2_decap_8 FILLER_28_415 ();
 sg13g2_decap_8 FILLER_28_422 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_48 ();
 sg13g2_fill_1 FILLER_29_50 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_67 ();
 sg13g2_decap_8 FILLER_29_74 ();
 sg13g2_decap_4 FILLER_29_81 ();
 sg13g2_fill_1 FILLER_29_85 ();
 sg13g2_decap_8 FILLER_29_96 ();
 sg13g2_decap_4 FILLER_29_103 ();
 sg13g2_decap_8 FILLER_29_141 ();
 sg13g2_fill_1 FILLER_29_148 ();
 sg13g2_fill_1 FILLER_29_153 ();
 sg13g2_fill_1 FILLER_29_159 ();
 sg13g2_fill_2 FILLER_29_164 ();
 sg13g2_fill_1 FILLER_29_171 ();
 sg13g2_fill_2 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_fill_1 FILLER_29_214 ();
 sg13g2_decap_4 FILLER_29_219 ();
 sg13g2_decap_8 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_234 ();
 sg13g2_fill_2 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_254 ();
 sg13g2_decap_8 FILLER_29_261 ();
 sg13g2_fill_1 FILLER_29_268 ();
 sg13g2_decap_4 FILLER_29_273 ();
 sg13g2_decap_4 FILLER_29_287 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_decap_8 FILLER_29_319 ();
 sg13g2_fill_2 FILLER_29_326 ();
 sg13g2_fill_1 FILLER_29_331 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_fill_2 FILLER_29_374 ();
 sg13g2_fill_1 FILLER_29_376 ();
 sg13g2_fill_1 FILLER_29_403 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_27 ();
 sg13g2_fill_1 FILLER_30_29 ();
 sg13g2_decap_8 FILLER_30_38 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_4 FILLER_30_120 ();
 sg13g2_fill_2 FILLER_30_128 ();
 sg13g2_decap_8 FILLER_30_134 ();
 sg13g2_decap_8 FILLER_30_141 ();
 sg13g2_decap_4 FILLER_30_148 ();
 sg13g2_fill_2 FILLER_30_152 ();
 sg13g2_decap_8 FILLER_30_159 ();
 sg13g2_decap_4 FILLER_30_171 ();
 sg13g2_fill_1 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_decap_4 FILLER_30_214 ();
 sg13g2_fill_2 FILLER_30_218 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_262 ();
 sg13g2_fill_2 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_271 ();
 sg13g2_decap_8 FILLER_30_277 ();
 sg13g2_decap_8 FILLER_30_284 ();
 sg13g2_decap_8 FILLER_30_291 ();
 sg13g2_fill_2 FILLER_30_298 ();
 sg13g2_fill_1 FILLER_30_300 ();
 sg13g2_decap_8 FILLER_30_305 ();
 sg13g2_decap_4 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_316 ();
 sg13g2_decap_8 FILLER_30_380 ();
 sg13g2_decap_8 FILLER_30_387 ();
 sg13g2_decap_4 FILLER_30_394 ();
 sg13g2_fill_1 FILLER_30_398 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_12 ();
 sg13g2_decap_4 FILLER_31_19 ();
 sg13g2_fill_1 FILLER_31_23 ();
 sg13g2_decap_8 FILLER_31_36 ();
 sg13g2_fill_1 FILLER_31_43 ();
 sg13g2_decap_4 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_57 ();
 sg13g2_decap_8 FILLER_31_64 ();
 sg13g2_decap_4 FILLER_31_71 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_4 FILLER_31_108 ();
 sg13g2_fill_1 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_149 ();
 sg13g2_decap_4 FILLER_31_161 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_decap_8 FILLER_31_172 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_fill_1 FILLER_31_206 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_fill_1 FILLER_31_238 ();
 sg13g2_fill_2 FILLER_31_265 ();
 sg13g2_fill_1 FILLER_31_311 ();
 sg13g2_decap_8 FILLER_31_317 ();
 sg13g2_fill_2 FILLER_31_332 ();
 sg13g2_decap_4 FILLER_31_400 ();
 sg13g2_decap_8 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_31_415 ();
 sg13g2_decap_8 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_4 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_53 ();
 sg13g2_fill_1 FILLER_32_70 ();
 sg13g2_decap_4 FILLER_32_75 ();
 sg13g2_fill_2 FILLER_32_79 ();
 sg13g2_fill_2 FILLER_32_86 ();
 sg13g2_fill_1 FILLER_32_88 ();
 sg13g2_decap_8 FILLER_32_95 ();
 sg13g2_decap_4 FILLER_32_102 ();
 sg13g2_fill_1 FILLER_32_106 ();
 sg13g2_decap_8 FILLER_32_123 ();
 sg13g2_fill_2 FILLER_32_130 ();
 sg13g2_decap_4 FILLER_32_136 ();
 sg13g2_fill_1 FILLER_32_140 ();
 sg13g2_fill_2 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_249 ();
 sg13g2_decap_4 FILLER_32_256 ();
 sg13g2_fill_2 FILLER_32_260 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_fill_1 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_297 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_341 ();
 sg13g2_fill_1 FILLER_32_348 ();
 sg13g2_fill_1 FILLER_32_353 ();
 sg13g2_fill_1 FILLER_32_359 ();
 sg13g2_fill_1 FILLER_32_386 ();
 sg13g2_fill_1 FILLER_32_391 ();
 sg13g2_fill_1 FILLER_32_397 ();
 sg13g2_fill_2 FILLER_32_424 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_13 ();
 sg13g2_decap_4 FILLER_33_19 ();
 sg13g2_fill_2 FILLER_33_23 ();
 sg13g2_decap_8 FILLER_33_41 ();
 sg13g2_decap_8 FILLER_33_48 ();
 sg13g2_fill_2 FILLER_33_55 ();
 sg13g2_fill_1 FILLER_33_57 ();
 sg13g2_fill_1 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_90 ();
 sg13g2_decap_8 FILLER_33_97 ();
 sg13g2_fill_2 FILLER_33_104 ();
 sg13g2_decap_4 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_130 ();
 sg13g2_decap_8 FILLER_33_181 ();
 sg13g2_decap_8 FILLER_33_188 ();
 sg13g2_fill_2 FILLER_33_195 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_235 ();
 sg13g2_decap_4 FILLER_33_242 ();
 sg13g2_decap_4 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_255 ();
 sg13g2_fill_2 FILLER_33_282 ();
 sg13g2_decap_8 FILLER_33_320 ();
 sg13g2_decap_4 FILLER_33_327 ();
 sg13g2_fill_1 FILLER_33_331 ();
 sg13g2_decap_4 FILLER_33_336 ();
 sg13g2_fill_1 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_346 ();
 sg13g2_decap_8 FILLER_33_353 ();
 sg13g2_decap_8 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_33_367 ();
 sg13g2_fill_2 FILLER_33_374 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_33_415 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_28 ();
 sg13g2_fill_2 FILLER_34_33 ();
 sg13g2_fill_1 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_76 ();
 sg13g2_fill_1 FILLER_34_83 ();
 sg13g2_decap_4 FILLER_34_89 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_4 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_114 ();
 sg13g2_fill_2 FILLER_34_121 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_decap_8 FILLER_34_137 ();
 sg13g2_decap_8 FILLER_34_157 ();
 sg13g2_fill_1 FILLER_34_164 ();
 sg13g2_fill_2 FILLER_34_175 ();
 sg13g2_fill_2 FILLER_34_187 ();
 sg13g2_fill_1 FILLER_34_189 ();
 sg13g2_fill_2 FILLER_34_196 ();
 sg13g2_fill_1 FILLER_34_204 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_decap_4 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_263 ();
 sg13g2_decap_8 FILLER_34_274 ();
 sg13g2_decap_8 FILLER_34_281 ();
 sg13g2_decap_4 FILLER_34_288 ();
 sg13g2_decap_4 FILLER_34_301 ();
 sg13g2_fill_1 FILLER_34_305 ();
 sg13g2_fill_2 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_315 ();
 sg13g2_fill_2 FILLER_34_377 ();
 sg13g2_fill_1 FILLER_34_386 ();
 sg13g2_decap_8 FILLER_34_409 ();
 sg13g2_decap_8 FILLER_34_416 ();
 sg13g2_decap_8 FILLER_34_423 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_fill_1 FILLER_35_9 ();
 sg13g2_fill_2 FILLER_35_36 ();
 sg13g2_fill_2 FILLER_35_46 ();
 sg13g2_fill_1 FILLER_35_48 ();
 sg13g2_decap_4 FILLER_35_54 ();
 sg13g2_fill_1 FILLER_35_58 ();
 sg13g2_fill_1 FILLER_35_65 ();
 sg13g2_fill_2 FILLER_35_78 ();
 sg13g2_fill_1 FILLER_35_108 ();
 sg13g2_fill_1 FILLER_35_117 ();
 sg13g2_fill_2 FILLER_35_130 ();
 sg13g2_fill_1 FILLER_35_132 ();
 sg13g2_fill_2 FILLER_35_138 ();
 sg13g2_decap_4 FILLER_35_158 ();
 sg13g2_decap_8 FILLER_35_172 ();
 sg13g2_decap_8 FILLER_35_187 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_fill_1 FILLER_35_210 ();
 sg13g2_fill_2 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_233 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_decap_8 FILLER_35_244 ();
 sg13g2_fill_1 FILLER_35_251 ();
 sg13g2_fill_1 FILLER_35_310 ();
 sg13g2_fill_1 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_349 ();
 sg13g2_fill_1 FILLER_35_356 ();
 sg13g2_fill_2 FILLER_35_361 ();
 sg13g2_fill_1 FILLER_35_363 ();
 sg13g2_decap_8 FILLER_35_368 ();
 sg13g2_decap_4 FILLER_35_375 ();
 sg13g2_decap_4 FILLER_35_384 ();
 sg13g2_fill_1 FILLER_35_403 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_20 ();
 sg13g2_decap_8 FILLER_36_27 ();
 sg13g2_decap_8 FILLER_36_34 ();
 sg13g2_decap_8 FILLER_36_41 ();
 sg13g2_decap_8 FILLER_36_48 ();
 sg13g2_decap_8 FILLER_36_55 ();
 sg13g2_decap_4 FILLER_36_62 ();
 sg13g2_fill_2 FILLER_36_66 ();
 sg13g2_decap_8 FILLER_36_76 ();
 sg13g2_fill_2 FILLER_36_83 ();
 sg13g2_fill_1 FILLER_36_85 ();
 sg13g2_fill_2 FILLER_36_101 ();
 sg13g2_decap_8 FILLER_36_111 ();
 sg13g2_decap_8 FILLER_36_118 ();
 sg13g2_fill_2 FILLER_36_132 ();
 sg13g2_fill_2 FILLER_36_139 ();
 sg13g2_decap_8 FILLER_36_145 ();
 sg13g2_fill_2 FILLER_36_152 ();
 sg13g2_fill_2 FILLER_36_158 ();
 sg13g2_fill_1 FILLER_36_160 ();
 sg13g2_fill_1 FILLER_36_165 ();
 sg13g2_fill_2 FILLER_36_174 ();
 sg13g2_decap_8 FILLER_36_180 ();
 sg13g2_decap_8 FILLER_36_187 ();
 sg13g2_fill_1 FILLER_36_194 ();
 sg13g2_decap_8 FILLER_36_212 ();
 sg13g2_decap_8 FILLER_36_219 ();
 sg13g2_decap_8 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_233 ();
 sg13g2_decap_8 FILLER_36_265 ();
 sg13g2_decap_8 FILLER_36_272 ();
 sg13g2_decap_4 FILLER_36_279 ();
 sg13g2_decap_4 FILLER_36_287 ();
 sg13g2_fill_1 FILLER_36_291 ();
 sg13g2_fill_2 FILLER_36_302 ();
 sg13g2_decap_4 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_decap_4 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_328 ();
 sg13g2_decap_8 FILLER_36_334 ();
 sg13g2_decap_8 FILLER_36_341 ();
 sg13g2_decap_8 FILLER_36_348 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_fill_2 FILLER_36_383 ();
 sg13g2_decap_4 FILLER_36_395 ();
 sg13g2_fill_1 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_fill_2 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_44 ();
 sg13g2_decap_8 FILLER_37_90 ();
 sg13g2_fill_2 FILLER_37_97 ();
 sg13g2_fill_1 FILLER_37_159 ();
 sg13g2_fill_1 FILLER_37_165 ();
 sg13g2_fill_1 FILLER_37_171 ();
 sg13g2_fill_1 FILLER_37_177 ();
 sg13g2_fill_1 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_198 ();
 sg13g2_decap_4 FILLER_37_205 ();
 sg13g2_fill_2 FILLER_37_209 ();
 sg13g2_fill_1 FILLER_37_215 ();
 sg13g2_fill_2 FILLER_37_220 ();
 sg13g2_decap_4 FILLER_37_252 ();
 sg13g2_fill_2 FILLER_37_256 ();
 sg13g2_decap_8 FILLER_37_262 ();
 sg13g2_fill_2 FILLER_37_269 ();
 sg13g2_fill_1 FILLER_37_271 ();
 sg13g2_decap_8 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_283 ();
 sg13g2_fill_1 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_fill_2 FILLER_37_427 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_fill_2 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_55 ();
 sg13g2_decap_4 FILLER_38_62 ();
 sg13g2_fill_2 FILLER_38_66 ();
 sg13g2_fill_2 FILLER_38_89 ();
 sg13g2_fill_1 FILLER_38_103 ();
 sg13g2_fill_1 FILLER_38_112 ();
 sg13g2_fill_1 FILLER_38_133 ();
 sg13g2_fill_1 FILLER_38_142 ();
 sg13g2_fill_2 FILLER_38_147 ();
 sg13g2_fill_2 FILLER_38_153 ();
 sg13g2_fill_2 FILLER_38_159 ();
 sg13g2_fill_1 FILLER_38_161 ();
 sg13g2_fill_2 FILLER_38_184 ();
 sg13g2_decap_4 FILLER_38_190 ();
 sg13g2_fill_1 FILLER_38_194 ();
 sg13g2_fill_2 FILLER_38_216 ();
 sg13g2_fill_1 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_239 ();
 sg13g2_fill_2 FILLER_38_264 ();
 sg13g2_fill_1 FILLER_38_292 ();
 sg13g2_decap_4 FILLER_38_297 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_decap_4 FILLER_38_313 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_decap_8 FILLER_38_327 ();
 sg13g2_decap_4 FILLER_38_334 ();
 sg13g2_fill_2 FILLER_38_338 ();
 sg13g2_fill_1 FILLER_38_345 ();
 sg13g2_fill_2 FILLER_38_350 ();
 sg13g2_fill_1 FILLER_38_383 ();
 sg13g2_fill_2 FILLER_38_388 ();
 sg13g2_fill_2 FILLER_38_394 ();
 sg13g2_fill_2 FILLER_38_400 ();
 sg13g2_fill_1 FILLER_38_402 ();
 sg13g2_decap_8 FILLER_38_412 ();
 sg13g2_decap_8 FILLER_38_419 ();
 sg13g2_decap_4 FILLER_38_426 ();
endmodule
