module tt_um_calonso88_74181 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire clknet_0_clk;
 wire net166;
 wire \alu_74181_i0.a[0] ;
 wire \alu_74181_i0.a[1] ;
 wire \alu_74181_i0.a[2] ;
 wire \alu_74181_i0.a[3] ;
 wire \alu_74181_i0.alu_74181_arith_inst.b[0] ;
 wire \alu_74181_i0.alu_74181_arith_inst.b[1] ;
 wire \alu_74181_i0.alu_74181_arith_inst.b[2] ;
 wire \alu_74181_i0.alu_74181_arith_inst.b[3] ;
 wire \alu_74181_i0.alu_74181_arith_inst.cn ;
 wire \alu_74181_i0.alu_74181_arith_inst.s[0] ;
 wire \alu_74181_i0.alu_74181_arith_inst.s[1] ;
 wire \alu_74181_i0.alu_74181_arith_inst.s[2] ;
 wire \alu_74181_i0.alu_74181_arith_inst.s[3] ;
 wire \alu_74181_i0.m ;
 wire \alu_74181_i1.a[0] ;
 wire \alu_74181_i1.a[1] ;
 wire \alu_74181_i1.a[2] ;
 wire \alu_74181_i1.a[3] ;
 wire \alu_74181_i1.alu_74181_arith_inst.b[0] ;
 wire \alu_74181_i1.alu_74181_arith_inst.b[1] ;
 wire \alu_74181_i1.alu_74181_arith_inst.b[2] ;
 wire \alu_74181_i1.alu_74181_arith_inst.b[3] ;
 wire \config_regs[22] ;
 wire \config_regs[23] ;
 wire \config_regs[24] ;
 wire \config_regs[25] ;
 wire \config_regs[26] ;
 wire \config_regs[27] ;
 wire \config_regs[28] ;
 wire \config_regs[29] ;
 wire \config_regs[30] ;
 wire \config_regs[31] ;
 wire \config_regs[32] ;
 wire \config_regs[33] ;
 wire \config_regs[34] ;
 wire \config_regs[35] ;
 wire \config_regs[36] ;
 wire \config_regs[37] ;
 wire \config_regs[38] ;
 wire \config_regs[39] ;
 wire \config_regs[40] ;
 wire \config_regs[41] ;
 wire \config_regs[42] ;
 wire \config_regs[43] ;
 wire \config_regs[44] ;
 wire \config_regs[45] ;
 wire \config_regs[46] ;
 wire \config_regs[47] ;
 wire \config_regs[48] ;
 wire \config_regs[49] ;
 wire \config_regs[50] ;
 wire \config_regs[51] ;
 wire \config_regs[52] ;
 wire \config_regs[53] ;
 wire \config_regs[54] ;
 wire \config_regs[55] ;
 wire \config_regs[56] ;
 wire \config_regs[57] ;
 wire \config_regs[58] ;
 wire \config_regs[59] ;
 wire \config_regs[60] ;
 wire \config_regs[61] ;
 wire \config_regs[62] ;
 wire \config_regs[63] ;
 wire cpha_sync;
 wire cpol_sync;
 wire spi_clk_sync;
 wire spi_cs_n_sync;
 wire spi_miso;
 wire spi_mosi_sync;
 wire \spi_wrapper_i.reg_addr[0] ;
 wire \spi_wrapper_i.reg_addr[1] ;
 wire \spi_wrapper_i.reg_addr[2] ;
 wire \spi_wrapper_i.reg_addr[3] ;
 wire \spi_wrapper_i.reg_data_o[0] ;
 wire \spi_wrapper_i.reg_data_o[1] ;
 wire \spi_wrapper_i.reg_data_o[2] ;
 wire \spi_wrapper_i.reg_data_o[3] ;
 wire \spi_wrapper_i.reg_data_o[4] ;
 wire \spi_wrapper_i.reg_data_o[5] ;
 wire \spi_wrapper_i.reg_data_o[6] ;
 wire \spi_wrapper_i.reg_data_o[7] ;
 wire \spi_wrapper_i.reg_data_o_vld ;
 wire \spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ;
 wire \spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ;
 wire \spi_wrapper_i.spi_reg_inst.reg_rw ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[0] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[1] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[2] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[3] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[4] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[5] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[6] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer[7] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ;
 wire \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ;
 wire \spi_wrapper_i.spi_reg_inst.state[0] ;
 wire \spi_wrapper_i.spi_reg_inst.state[1] ;
 wire \spi_wrapper_i.spi_reg_inst.state[2] ;
 wire \spi_wrapper_i.spi_reg_inst.state[3] ;
 wire \spi_wrapper_i.spi_reg_inst.state[4] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[0] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[1] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[2] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[3] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[4] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[5] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer[6] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ;
 wire \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ;
 wire \synchronizer_spi_clk_inst.data_sync[1] ;
 wire \synchronizer_spi_cs_n_inst.data_sync[1] ;
 wire \synchronizer_spi_mode_cpha.data_sync[1] ;
 wire \synchronizer_spi_mode_cpol.data_sync[1] ;
 wire \synchronizer_spi_mosi_inst.data_sync[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_1 _1560_ (.A(ena),
    .X(_0749_));
 sg13g2_buf_1 _1561_ (.A(_0749_),
    .X(_0750_));
 sg13g2_nand2_1 _1562_ (.Y(_0751_),
    .A(net132),
    .B(\spi_wrapper_i.spi_reg_inst.state[2] ));
 sg13g2_buf_1 _1563_ (.A(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .X(_0752_));
 sg13g2_buf_2 _1564_ (.A(spi_cs_n_sync),
    .X(_0753_));
 sg13g2_nor2b_1 _1565_ (.A(_0752_),
    .B_N(_0753_),
    .Y(_0754_));
 sg13g2_buf_1 _1566_ (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ),
    .X(_0755_));
 sg13g2_buf_1 _1567_ (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ),
    .X(_0756_));
 sg13g2_buf_1 _1568_ (.A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ),
    .X(_0757_));
 sg13g2_nor3_2 _1569_ (.A(_0756_),
    .B(_0757_),
    .C(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .Y(_0758_));
 sg13g2_mux2_1 _1570_ (.A0(_0754_),
    .A1(_0755_),
    .S(_0758_),
    .X(_0759_));
 sg13g2_nand2_1 _1571_ (.Y(_0760_),
    .A(_0750_),
    .B(_0759_));
 sg13g2_nand2_1 _1572_ (.Y(_0761_),
    .A(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .B(_0760_));
 sg13g2_o21ai_1 _1573_ (.B1(_0761_),
    .Y(_0000_),
    .A1(\spi_wrapper_i.spi_reg_inst.reg_rw ),
    .A2(_0751_));
 sg13g2_inv_1 _1574_ (.Y(_0762_),
    .A(_0749_));
 sg13g2_buf_1 _1575_ (.A(_0762_),
    .X(_0763_));
 sg13g2_buf_2 _1576_ (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ),
    .X(_0764_));
 sg13g2_buf_1 _1577_ (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ),
    .X(_0765_));
 sg13g2_buf_1 _1578_ (.A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ),
    .X(_0766_));
 sg13g2_nor2_1 _1579_ (.A(_0765_),
    .B(_0766_),
    .Y(_0767_));
 sg13g2_nand3b_1 _1580_ (.B(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ),
    .C(_0767_),
    .Y(_0768_),
    .A_N(_0764_));
 sg13g2_nand2_1 _1581_ (.Y(_0769_),
    .A(net132),
    .B(\spi_wrapper_i.spi_reg_inst.state[3] ));
 sg13g2_nor2_1 _1582_ (.A(_0768_),
    .B(_0769_),
    .Y(_0770_));
 sg13g2_buf_1 _1583_ (.A(_0770_),
    .X(_0771_));
 sg13g2_a21o_1 _1584_ (.A2(\spi_wrapper_i.spi_reg_inst.state[2] ),
    .A1(net112),
    .B1(_0771_),
    .X(_0001_));
 sg13g2_inv_1 _1585_ (.Y(_0772_),
    .A(_0752_));
 sg13g2_nor2_1 _1586_ (.A(_0762_),
    .B(_0772_),
    .Y(_0773_));
 sg13g2_a22oi_1 _1587_ (.Y(_0774_),
    .B1(_0773_),
    .B2(\spi_wrapper_i.spi_reg_inst.state[0] ),
    .A2(_0768_),
    .A1(\spi_wrapper_i.spi_reg_inst.state[3] ));
 sg13g2_inv_1 _1588_ (.Y(_0775_),
    .A(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ));
 sg13g2_nor4_2 _1589_ (.A(_0764_),
    .B(_0765_),
    .C(_0775_),
    .Y(_0776_),
    .D(_0766_));
 sg13g2_o21ai_1 _1590_ (.B1(net132),
    .Y(_0777_),
    .A1(_0772_),
    .A2(_0776_));
 sg13g2_nand2_1 _1591_ (.Y(_0778_),
    .A(\spi_wrapper_i.spi_reg_inst.state[3] ),
    .B(_0777_));
 sg13g2_o21ai_1 _1592_ (.B1(_0778_),
    .Y(_0002_),
    .A1(_0753_),
    .A2(_0774_));
 sg13g2_inv_1 _1593_ (.Y(_0779_),
    .A(\spi_wrapper_i.spi_reg_inst.reg_rw ));
 sg13g2_nor2_1 _1594_ (.A(_0754_),
    .B(_0776_),
    .Y(_0780_));
 sg13g2_o21ai_1 _1595_ (.B1(\spi_wrapper_i.spi_reg_inst.state[4] ),
    .Y(_0781_),
    .A1(net112),
    .A2(_0780_));
 sg13g2_o21ai_1 _1596_ (.B1(_0781_),
    .Y(_0003_),
    .A1(_0779_),
    .A2(_0751_));
 sg13g2_buf_1 _1597_ (.A(\alu_74181_i1.a[1] ),
    .X(_0782_));
 sg13g2_buf_1 _1598_ (.A(net131),
    .X(_0783_));
 sg13g2_buf_1 _1599_ (.A(\alu_74181_i0.alu_74181_arith_inst.s[0] ),
    .X(_0784_));
 sg13g2_buf_8 _1600_ (.A(\alu_74181_i0.alu_74181_arith_inst.s[2] ),
    .X(_0785_));
 sg13g2_nor2b_1 _1601_ (.A(net130),
    .B_N(net129),
    .Y(_0786_));
 sg13g2_buf_2 _1602_ (.A(_0786_),
    .X(_0787_));
 sg13g2_buf_2 _1603_ (.A(\alu_74181_i0.alu_74181_arith_inst.s[3] ),
    .X(_0788_));
 sg13g2_buf_8 _1604_ (.A(\alu_74181_i0.alu_74181_arith_inst.s[1] ),
    .X(_0789_));
 sg13g2_buf_8 _1605_ (.A(_0789_),
    .X(_0790_));
 sg13g2_nor2b_1 _1606_ (.A(_0788_),
    .B_N(net110),
    .Y(_0791_));
 sg13g2_buf_2 _1607_ (.A(_0791_),
    .X(_0792_));
 sg13g2_nand2_1 _1608_ (.Y(_0793_),
    .A(_0787_),
    .B(_0792_));
 sg13g2_buf_1 _1609_ (.A(_0793_),
    .X(_0794_));
 sg13g2_buf_2 _1610_ (.A(\alu_74181_i1.alu_74181_arith_inst.b[1] ),
    .X(_0795_));
 sg13g2_buf_1 _1611_ (.A(_0795_),
    .X(_0796_));
 sg13g2_buf_1 _1612_ (.A(net109),
    .X(_0797_));
 sg13g2_buf_1 _1613_ (.A(\alu_74181_i1.alu_74181_arith_inst.b[0] ),
    .X(_0798_));
 sg13g2_buf_2 _1614_ (.A(\alu_74181_i1.a[0] ),
    .X(_0799_));
 sg13g2_nand2b_1 _1615_ (.Y(_0800_),
    .B(_0799_),
    .A_N(_0798_));
 sg13g2_buf_1 _1616_ (.A(_0800_),
    .X(_0801_));
 sg13g2_xor2_1 _1617_ (.B(net83),
    .A(_0797_),
    .X(_0802_));
 sg13g2_buf_1 _1618_ (.A(net129),
    .X(_0803_));
 sg13g2_inv_1 _1619_ (.Y(_0804_),
    .A(net108));
 sg13g2_buf_8 _1620_ (.A(_0788_),
    .X(_0805_));
 sg13g2_inv_2 _1621_ (.Y(_0806_),
    .A(net107));
 sg13g2_nand2_1 _1622_ (.Y(_0807_),
    .A(_0804_),
    .B(net82));
 sg13g2_buf_1 _1623_ (.A(_0807_),
    .X(_0808_));
 sg13g2_o21ai_1 _1624_ (.B1(net41),
    .Y(_0809_),
    .A1(net29),
    .A2(_0802_));
 sg13g2_nor2_1 _1625_ (.A(net111),
    .B(net29),
    .Y(_0810_));
 sg13g2_buf_1 _1626_ (.A(net130),
    .X(_0811_));
 sg13g2_inv_2 _1627_ (.Y(_0812_),
    .A(net110));
 sg13g2_nor2_1 _1628_ (.A(net106),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_buf_2 _1629_ (.A(_0813_),
    .X(_0814_));
 sg13g2_buf_1 _1630_ (.A(net110),
    .X(_0815_));
 sg13g2_nor2_1 _1631_ (.A(net81),
    .B(net84),
    .Y(_0816_));
 sg13g2_buf_1 _1632_ (.A(net106),
    .X(_0817_));
 sg13g2_a221oi_1 _1633_ (.B2(net80),
    .C1(net41),
    .B1(_0816_),
    .A1(net84),
    .Y(_0818_),
    .A2(_0814_));
 sg13g2_a221oi_1 _1634_ (.B2(_0802_),
    .C1(_0818_),
    .B1(_0810_),
    .A1(net111),
    .Y(_0819_),
    .A2(_0809_));
 sg13g2_buf_1 _1635_ (.A(net107),
    .X(_0820_));
 sg13g2_nand2_1 _1636_ (.Y(_0821_),
    .A(net130),
    .B(net129));
 sg13g2_buf_1 _1637_ (.A(_0821_),
    .X(_0822_));
 sg13g2_nor2_1 _1638_ (.A(net79),
    .B(net78),
    .Y(_0823_));
 sg13g2_buf_2 _1639_ (.A(_0823_),
    .X(_0824_));
 sg13g2_buf_8 _1640_ (.A(_0799_),
    .X(_0825_));
 sg13g2_inv_1 _1641_ (.Y(_0826_),
    .A(net105));
 sg13g2_buf_1 _1642_ (.A(_0798_),
    .X(_0827_));
 sg13g2_nor2_2 _1643_ (.A(_0826_),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_inv_1 _1644_ (.Y(_0829_),
    .A(_0782_));
 sg13g2_nand2b_1 _1645_ (.Y(_0830_),
    .B(net110),
    .A_N(net107));
 sg13g2_buf_2 _1646_ (.A(_0830_),
    .X(_0831_));
 sg13g2_nor2_2 _1647_ (.A(net78),
    .B(_0831_),
    .Y(_0832_));
 sg13g2_a21oi_1 _1648_ (.A1(_0829_),
    .A2(_0832_),
    .Y(_0833_),
    .B1(net84));
 sg13g2_xnor2_1 _1649_ (.Y(_0834_),
    .A(_0828_),
    .B(_0833_));
 sg13g2_buf_1 _1650_ (.A(net104),
    .X(_0835_));
 sg13g2_nand2_2 _1651_ (.Y(_0836_),
    .A(net105),
    .B(net77));
 sg13g2_and2_1 _1652_ (.A(_0788_),
    .B(_0789_),
    .X(_0837_));
 sg13g2_buf_2 _1653_ (.A(_0837_),
    .X(_0838_));
 sg13g2_nor2b_1 _1654_ (.A(net108),
    .B_N(net106),
    .Y(_0839_));
 sg13g2_nand2_2 _1655_ (.Y(_0840_),
    .A(_0838_),
    .B(_0839_));
 sg13g2_o21ai_1 _1656_ (.B1(net84),
    .Y(_0841_),
    .A1(net111),
    .A2(_0840_));
 sg13g2_xnor2_1 _1657_ (.Y(_0842_),
    .A(_0836_),
    .B(_0841_));
 sg13g2_nor3_2 _1658_ (.A(net108),
    .B(net82),
    .C(_0812_),
    .Y(_0843_));
 sg13g2_a22oi_1 _1659_ (.Y(_0844_),
    .B1(_0842_),
    .B2(_0843_),
    .A2(_0834_),
    .A1(_0824_));
 sg13g2_nand2_1 _1660_ (.Y(_0845_),
    .A(_0819_),
    .B(_0844_));
 sg13g2_nor2_2 _1661_ (.A(net106),
    .B(_0803_),
    .Y(_0846_));
 sg13g2_nor2b_1 _1662_ (.A(net110),
    .B_N(_0788_),
    .Y(_0847_));
 sg13g2_buf_2 _1663_ (.A(_0847_),
    .X(_0848_));
 sg13g2_a21oi_1 _1664_ (.A1(_0846_),
    .A2(_0848_),
    .Y(_0849_),
    .B1(net109));
 sg13g2_and2_1 _1665_ (.A(\alu_74181_i1.a[1] ),
    .B(_0795_),
    .X(_0850_));
 sg13g2_buf_1 _1666_ (.A(_0850_),
    .X(_0851_));
 sg13g2_and2_1 _1667_ (.A(net104),
    .B(_0851_),
    .X(_0852_));
 sg13g2_buf_1 _1668_ (.A(net105),
    .X(_0853_));
 sg13g2_o21ai_1 _1669_ (.B1(net76),
    .Y(_0854_),
    .A1(_0849_),
    .A2(_0852_));
 sg13g2_inv_1 _1670_ (.Y(_0855_),
    .A(net104));
 sg13g2_nand2b_1 _1671_ (.Y(_0856_),
    .B(_0795_),
    .A_N(net131));
 sg13g2_buf_2 _1672_ (.A(_0856_),
    .X(_0857_));
 sg13g2_nor2_1 _1673_ (.A(_0855_),
    .B(_0857_),
    .Y(_0858_));
 sg13g2_a21oi_1 _1674_ (.A1(_0838_),
    .A2(_0787_),
    .Y(_0859_),
    .B1(net109));
 sg13g2_o21ai_1 _1675_ (.B1(_0826_),
    .Y(_0860_),
    .A1(_0858_),
    .A2(_0859_));
 sg13g2_or2_1 _1676_ (.X(_0861_),
    .B(net129),
    .A(net130));
 sg13g2_buf_2 _1677_ (.A(_0861_),
    .X(_0862_));
 sg13g2_nand2b_1 _1678_ (.Y(_0863_),
    .B(_0788_),
    .A_N(_0789_));
 sg13g2_buf_8 _1679_ (.A(_0863_),
    .X(_0864_));
 sg13g2_o21ai_1 _1680_ (.B1(net111),
    .Y(_0865_),
    .A1(_0862_),
    .A2(net75));
 sg13g2_a21o_1 _1681_ (.A2(_0865_),
    .A1(net84),
    .B1(net77),
    .X(_0866_));
 sg13g2_nand2_1 _1682_ (.Y(_0867_),
    .A(_0846_),
    .B(_0848_));
 sg13g2_nor2_1 _1683_ (.A(net77),
    .B(net111),
    .Y(_0868_));
 sg13g2_nand2_1 _1684_ (.Y(_0869_),
    .A(_0838_),
    .B(_0787_));
 sg13g2_o21ai_1 _1685_ (.B1(_0869_),
    .Y(_0870_),
    .A1(_0867_),
    .A2(_0868_));
 sg13g2_nand4_1 _1686_ (.B(_0860_),
    .C(_0866_),
    .A(_0854_),
    .Y(_0871_),
    .D(_0870_));
 sg13g2_nor2_1 _1687_ (.A(net75),
    .B(_0822_),
    .Y(_0872_));
 sg13g2_buf_1 _1688_ (.A(_0872_),
    .X(_0873_));
 sg13g2_nor2_1 _1689_ (.A(_0799_),
    .B(net104),
    .Y(_0874_));
 sg13g2_nor2_1 _1690_ (.A(net131),
    .B(net109),
    .Y(_0875_));
 sg13g2_xor2_1 _1691_ (.B(_0875_),
    .A(_0874_),
    .X(_0876_));
 sg13g2_inv_1 _1692_ (.Y(_0877_),
    .A(net130));
 sg13g2_xnor2_1 _1693_ (.Y(_0878_),
    .A(net104),
    .B(net109));
 sg13g2_o21ai_1 _1694_ (.B1(_0812_),
    .Y(_0879_),
    .A1(net103),
    .A2(_0878_));
 sg13g2_nand2_1 _1695_ (.Y(_0880_),
    .A(_0848_),
    .B(_0787_));
 sg13g2_xnor2_1 _1696_ (.Y(_0881_),
    .A(net105),
    .B(net131));
 sg13g2_o21ai_1 _1697_ (.B1(net107),
    .Y(_0882_),
    .A1(_0880_),
    .A2(_0881_));
 sg13g2_a221oi_1 _1698_ (.B2(_0804_),
    .C1(_0882_),
    .B1(_0879_),
    .A1(net40),
    .Y(_0883_),
    .A2(_0876_));
 sg13g2_nand2b_1 _1699_ (.Y(_0884_),
    .B(net131),
    .A_N(_0795_));
 sg13g2_buf_1 _1700_ (.A(_0884_),
    .X(_0885_));
 sg13g2_nand2_1 _1701_ (.Y(_0886_),
    .A(_0885_),
    .B(net83));
 sg13g2_nor2_1 _1702_ (.A(_0829_),
    .B(net84),
    .Y(_0887_));
 sg13g2_nand2_1 _1703_ (.Y(_0888_),
    .A(_0887_),
    .B(_0828_));
 sg13g2_nand2b_2 _1704_ (.Y(_0889_),
    .B(_0789_),
    .A_N(net129));
 sg13g2_and2_1 _1705_ (.A(net107),
    .B(_0889_),
    .X(_0890_));
 sg13g2_buf_2 _1706_ (.A(_0890_),
    .X(_0891_));
 sg13g2_a21oi_1 _1707_ (.A1(_0886_),
    .A2(_0888_),
    .Y(_0892_),
    .B1(_0891_));
 sg13g2_a21o_1 _1708_ (.A2(_0883_),
    .A1(_0871_),
    .B1(_0892_),
    .X(_0893_));
 sg13g2_buf_1 _1709_ (.A(_0024_),
    .X(_0894_));
 sg13g2_nand2_2 _1710_ (.Y(_0895_),
    .A(net107),
    .B(_0889_));
 sg13g2_nor3_1 _1711_ (.A(net110),
    .B(net78),
    .C(_0874_),
    .Y(_0896_));
 sg13g2_or2_1 _1712_ (.X(_0897_),
    .B(_0025_),
    .A(net108));
 sg13g2_a21oi_1 _1713_ (.A1(_0812_),
    .A2(_0897_),
    .Y(_0898_),
    .B1(net103));
 sg13g2_nand2b_1 _1714_ (.Y(_0899_),
    .B(net107),
    .A_N(net106));
 sg13g2_xor2_1 _1715_ (.B(_0789_),
    .A(_0785_),
    .X(_0900_));
 sg13g2_a21oi_1 _1716_ (.A1(net108),
    .A2(net110),
    .Y(_0901_),
    .B1(_0827_));
 sg13g2_nor2b_1 _1717_ (.A(_0799_),
    .B_N(_0798_),
    .Y(_0902_));
 sg13g2_buf_2 _1718_ (.A(_0902_),
    .X(_0903_));
 sg13g2_nor4_1 _1719_ (.A(_0899_),
    .B(_0900_),
    .C(_0901_),
    .D(_0903_),
    .Y(_0904_));
 sg13g2_or4_1 _1720_ (.A(_0895_),
    .B(_0896_),
    .C(_0898_),
    .D(_0904_),
    .X(_0905_));
 sg13g2_nand2_1 _1721_ (.Y(_0906_),
    .A(_0895_),
    .B(net83));
 sg13g2_and3_1 _1722_ (.X(_0907_),
    .A(_0894_),
    .B(_0905_),
    .C(_0906_));
 sg13g2_buf_1 _1723_ (.A(_0907_),
    .X(_0908_));
 sg13g2_xnor2_1 _1724_ (.Y(_0909_),
    .A(_0893_),
    .B(_0908_));
 sg13g2_nand2_1 _1725_ (.Y(_0910_),
    .A(net82),
    .B(_0812_));
 sg13g2_buf_2 _1726_ (.A(_0910_),
    .X(_0911_));
 sg13g2_nor2_2 _1727_ (.A(_0862_),
    .B(_0911_),
    .Y(_0912_));
 sg13g2_inv_1 _1728_ (.Y(_0913_),
    .A(_0912_));
 sg13g2_o21ai_1 _1729_ (.B1(_0913_),
    .Y(_0914_),
    .A1(_0845_),
    .A2(_0909_));
 sg13g2_inv_1 _1730_ (.Y(_0915_),
    .A(_0023_));
 sg13g2_or2_1 _1731_ (.X(_0916_),
    .B(_0789_),
    .A(net130));
 sg13g2_buf_1 _1732_ (.A(_0916_),
    .X(_0917_));
 sg13g2_a21o_1 _1733_ (.A2(_0917_),
    .A1(net82),
    .B1(_0804_),
    .X(_0918_));
 sg13g2_and2_1 _1734_ (.A(net75),
    .B(_0918_),
    .X(_0919_));
 sg13g2_buf_1 _1735_ (.A(_0919_),
    .X(_0920_));
 sg13g2_a21oi_1 _1736_ (.A1(_0915_),
    .A2(_0909_),
    .Y(_0921_),
    .B1(net28));
 sg13g2_nor2_1 _1737_ (.A(_0845_),
    .B(_0921_),
    .Y(_0922_));
 sg13g2_a21oi_1 _1738_ (.A1(_0023_),
    .A2(_0914_),
    .Y(_0923_),
    .B1(_0922_));
 sg13g2_buf_2 _1739_ (.A(_0923_),
    .X(_0924_));
 sg13g2_buf_2 _1740_ (.A(\alu_74181_i0.m ),
    .X(_0925_));
 sg13g2_inv_1 _1741_ (.Y(_0926_),
    .A(_0925_));
 sg13g2_buf_1 _1742_ (.A(\config_regs[24] ),
    .X(_0927_));
 sg13g2_buf_4 _1743_ (.X(_0928_),
    .A(\config_regs[25] ));
 sg13g2_inv_1 _1744_ (.Y(_0929_),
    .A(\config_regs[26] ));
 sg13g2_nor2_1 _1745_ (.A(_0928_),
    .B(_0929_),
    .Y(_0930_));
 sg13g2_and2_1 _1746_ (.A(_0927_),
    .B(_0930_),
    .X(_0931_));
 sg13g2_buf_1 _1747_ (.A(_0931_),
    .X(_0932_));
 sg13g2_nand2_1 _1748_ (.Y(_0933_),
    .A(_0926_),
    .B(_0932_));
 sg13g2_nor2_1 _1749_ (.A(net103),
    .B(net110),
    .Y(_0934_));
 sg13g2_nand2_1 _1750_ (.Y(_0935_),
    .A(net82),
    .B(_0801_));
 sg13g2_buf_1 _1751_ (.A(net108),
    .X(_0936_));
 sg13g2_buf_1 _1752_ (.A(net82),
    .X(_0937_));
 sg13g2_a21oi_1 _1753_ (.A1(net81),
    .A2(_0836_),
    .Y(_0938_),
    .B1(net58));
 sg13g2_a221oi_1 _1754_ (.B2(net74),
    .C1(_0938_),
    .B1(_0935_),
    .A1(_0934_),
    .Y(_0939_),
    .A2(_0874_));
 sg13g2_nor2_1 _1755_ (.A(_0804_),
    .B(_0790_),
    .Y(_0940_));
 sg13g2_and2_1 _1756_ (.A(net81),
    .B(_0903_),
    .X(_0941_));
 sg13g2_o21ai_1 _1757_ (.B1(_0877_),
    .Y(_0942_),
    .A1(_0940_),
    .A2(_0941_));
 sg13g2_nor2_1 _1758_ (.A(_0894_),
    .B(_0880_),
    .Y(_0943_));
 sg13g2_o21ai_1 _1759_ (.B1(_0906_),
    .Y(_0944_),
    .A1(_0905_),
    .A2(_0943_));
 sg13g2_xnor2_1 _1760_ (.Y(_0945_),
    .A(net76),
    .B(_0944_));
 sg13g2_nand2_1 _1761_ (.Y(_0946_),
    .A(net75),
    .B(_0918_));
 sg13g2_buf_8 _1762_ (.A(_0946_),
    .X(_0947_));
 sg13g2_a22oi_1 _1763_ (.Y(_0948_),
    .B1(_0945_),
    .B2(_0947_),
    .A2(_0942_),
    .A1(_0939_));
 sg13g2_a21o_1 _1764_ (.A2(_0912_),
    .A1(_0894_),
    .B1(_0948_),
    .X(_0949_));
 sg13g2_buf_1 _1765_ (.A(_0949_),
    .X(_0950_));
 sg13g2_nor2_1 _1766_ (.A(_0933_),
    .B(_0950_),
    .Y(_0951_));
 sg13g2_nand2b_1 _1767_ (.Y(_0952_),
    .B(_0951_),
    .A_N(_0924_));
 sg13g2_buf_1 _1768_ (.A(_0926_),
    .X(_0953_));
 sg13g2_and2_1 _1769_ (.A(net73),
    .B(_0932_),
    .X(_0954_));
 sg13g2_nand2_1 _1770_ (.Y(_0955_),
    .A(_0954_),
    .B(_0924_));
 sg13g2_buf_2 _1771_ (.A(\alu_74181_i0.alu_74181_arith_inst.b[3] ),
    .X(_0956_));
 sg13g2_buf_1 _1772_ (.A(_0956_),
    .X(_0957_));
 sg13g2_buf_1 _1773_ (.A(_0957_),
    .X(_0958_));
 sg13g2_nand2_1 _1774_ (.Y(_0959_),
    .A(_0788_),
    .B(_0789_));
 sg13g2_buf_1 _1775_ (.A(_0959_),
    .X(_0960_));
 sg13g2_buf_1 _1776_ (.A(_0960_),
    .X(_0961_));
 sg13g2_nand2b_1 _1777_ (.Y(_0962_),
    .B(net130),
    .A_N(net129));
 sg13g2_buf_1 _1778_ (.A(_0962_),
    .X(_0963_));
 sg13g2_nor2_2 _1779_ (.A(net57),
    .B(net71),
    .Y(_0964_));
 sg13g2_buf_1 _1780_ (.A(_0964_),
    .X(_0965_));
 sg13g2_buf_1 _1781_ (.A(\alu_74181_i0.alu_74181_arith_inst.b[2] ),
    .X(_0966_));
 sg13g2_buf_1 _1782_ (.A(net128),
    .X(_0967_));
 sg13g2_buf_8 _1783_ (.A(\alu_74181_i0.alu_74181_arith_inst.b[1] ),
    .X(_0968_));
 sg13g2_buf_1 _1784_ (.A(net127),
    .X(_0969_));
 sg13g2_buf_8 _1785_ (.A(\alu_74181_i0.alu_74181_arith_inst.b[0] ),
    .X(_0970_));
 sg13g2_buf_8 _1786_ (.A(\alu_74181_i0.a[0] ),
    .X(_0971_));
 sg13g2_nand2_1 _1787_ (.Y(_0972_),
    .A(_0970_),
    .B(net126));
 sg13g2_buf_2 _1788_ (.A(_0972_),
    .X(_0973_));
 sg13g2_buf_8 _1789_ (.A(\alu_74181_i0.a[1] ),
    .X(_0974_));
 sg13g2_nand2_1 _1790_ (.Y(_0975_),
    .A(_0974_),
    .B(\alu_74181_i0.alu_74181_arith_inst.b[1] ));
 sg13g2_buf_2 _1791_ (.A(_0975_),
    .X(_0976_));
 sg13g2_o21ai_1 _1792_ (.B1(_0976_),
    .Y(_0977_),
    .A1(net100),
    .A2(_0973_));
 sg13g2_buf_1 _1793_ (.A(_0977_),
    .X(_0978_));
 sg13g2_buf_8 _1794_ (.A(\alu_74181_i0.a[2] ),
    .X(_0979_));
 sg13g2_nand2b_1 _1795_ (.Y(_0980_),
    .B(net128),
    .A_N(net124));
 sg13g2_o21ai_1 _1796_ (.B1(_0980_),
    .Y(_0981_),
    .A1(net101),
    .A2(_0978_));
 sg13g2_buf_1 _1797_ (.A(\alu_74181_i0.a[3] ),
    .X(_0982_));
 sg13g2_nand2_2 _1798_ (.Y(_0983_),
    .A(net124),
    .B(net128));
 sg13g2_nand3_1 _1799_ (.B(_0973_),
    .C(_0983_),
    .A(_0976_),
    .Y(_0984_));
 sg13g2_buf_1 _1800_ (.A(_0984_),
    .X(_0985_));
 sg13g2_nand3_1 _1801_ (.B(_0964_),
    .C(_0985_),
    .A(net123),
    .Y(_0986_));
 sg13g2_o21ai_1 _1802_ (.B1(_0986_),
    .Y(_0987_),
    .A1(net27),
    .A2(_0981_));
 sg13g2_inv_2 _1803_ (.Y(_0988_),
    .A(net123));
 sg13g2_inv_1 _1804_ (.Y(_0989_),
    .A(net102));
 sg13g2_a21oi_1 _1805_ (.A1(_0988_),
    .A2(net27),
    .Y(_0990_),
    .B1(_0989_));
 sg13g2_a21oi_1 _1806_ (.A1(net27),
    .A2(_0985_),
    .Y(_0991_),
    .B1(_0990_));
 sg13g2_a22oi_1 _1807_ (.Y(_0992_),
    .B1(_0991_),
    .B2(_0981_),
    .A2(_0987_),
    .A1(net72));
 sg13g2_nand2b_1 _1808_ (.Y(_0993_),
    .B(_0843_),
    .A_N(_0992_));
 sg13g2_nand2b_1 _1809_ (.Y(_0994_),
    .B(_0974_),
    .A_N(_0968_));
 sg13g2_nand2b_1 _1810_ (.Y(_0995_),
    .B(net126),
    .A_N(_0970_));
 sg13g2_buf_2 _1811_ (.A(_0995_),
    .X(_0996_));
 sg13g2_nand2_1 _1812_ (.Y(_0997_),
    .A(_0994_),
    .B(_0996_));
 sg13g2_inv_1 _1813_ (.Y(_0998_),
    .A(_0969_));
 sg13g2_o21ai_1 _1814_ (.B1(_0994_),
    .Y(_0999_),
    .A1(_0998_),
    .A2(_0996_));
 sg13g2_nor2b_1 _1815_ (.A(_0966_),
    .B_N(net124),
    .Y(_1000_));
 sg13g2_a221oi_1 _1816_ (.B2(_0967_),
    .C1(_1000_),
    .B1(_0999_),
    .A1(_0832_),
    .Y(_1001_),
    .A2(_0997_));
 sg13g2_nor2_2 _1817_ (.A(_0970_),
    .B(net126),
    .Y(_1002_));
 sg13g2_nor4_2 _1818_ (.A(_0970_),
    .B(net126),
    .C(net125),
    .Y(_1003_),
    .D(_0968_));
 sg13g2_nor2_2 _1819_ (.A(_0979_),
    .B(net128),
    .Y(_1004_));
 sg13g2_xnor2_1 _1820_ (.Y(_1005_),
    .A(_1003_),
    .B(_1004_));
 sg13g2_and2_1 _1821_ (.A(_0784_),
    .B(net108),
    .X(_1006_));
 sg13g2_buf_2 _1822_ (.A(_1006_),
    .X(_1007_));
 sg13g2_a21oi_1 _1823_ (.A1(_1007_),
    .A2(_0792_),
    .Y(_1008_),
    .B1(net100));
 sg13g2_nand3_1 _1824_ (.B(_1005_),
    .C(_1008_),
    .A(_1002_),
    .Y(_1009_));
 sg13g2_nand2_1 _1825_ (.Y(_1010_),
    .A(_1001_),
    .B(_1009_));
 sg13g2_a21oi_1 _1826_ (.A1(_0988_),
    .A2(_0832_),
    .Y(_1011_),
    .B1(net102));
 sg13g2_nand2_2 _1827_ (.Y(_1012_),
    .A(_1007_),
    .B(_0792_));
 sg13g2_and2_1 _1828_ (.A(_1003_),
    .B(_1004_),
    .X(_1013_));
 sg13g2_buf_1 _1829_ (.A(_1013_),
    .X(_1014_));
 sg13g2_nand2_1 _1830_ (.Y(_1015_),
    .A(_1012_),
    .B(_1014_));
 sg13g2_mux2_1 _1831_ (.A0(_0957_),
    .A1(_1011_),
    .S(_1015_),
    .X(_1016_));
 sg13g2_xnor2_1 _1832_ (.Y(_1017_),
    .A(_1010_),
    .B(_1016_));
 sg13g2_nor2b_1 _1833_ (.A(net124),
    .B_N(net128),
    .Y(_1018_));
 sg13g2_nand2b_1 _1834_ (.Y(_1019_),
    .B(net127),
    .A_N(net125));
 sg13g2_buf_1 _1835_ (.A(_0970_),
    .X(_1020_));
 sg13g2_buf_8 _1836_ (.A(_0971_),
    .X(_1021_));
 sg13g2_nor2b_1 _1837_ (.A(net99),
    .B_N(net98),
    .Y(_1022_));
 sg13g2_buf_1 _1838_ (.A(_1022_),
    .X(_1023_));
 sg13g2_nor2b_1 _1839_ (.A(net127),
    .B_N(net125),
    .Y(_1024_));
 sg13g2_buf_2 _1840_ (.A(_1024_),
    .X(_1025_));
 sg13g2_a21oi_1 _1841_ (.A1(_1019_),
    .A2(net56),
    .Y(_1026_),
    .B1(_1025_));
 sg13g2_nand2b_1 _1842_ (.Y(_1027_),
    .B(net124),
    .A_N(net128));
 sg13g2_o21ai_1 _1843_ (.B1(_1027_),
    .Y(_1028_),
    .A1(_1018_),
    .A2(_1026_));
 sg13g2_xnor2_1 _1844_ (.Y(_1029_),
    .A(net102),
    .B(_1028_));
 sg13g2_o21ai_1 _1845_ (.B1(net41),
    .Y(_1030_),
    .A1(net29),
    .A2(_1029_));
 sg13g2_buf_1 _1846_ (.A(_0982_),
    .X(_1031_));
 sg13g2_nor2_1 _1847_ (.A(net123),
    .B(net29),
    .Y(_1032_));
 sg13g2_nor2_1 _1848_ (.A(_0815_),
    .B(net102),
    .Y(_1033_));
 sg13g2_a221oi_1 _1849_ (.B2(_0811_),
    .C1(_0807_),
    .B1(_1033_),
    .A1(net102),
    .Y(_1034_),
    .A2(_0814_));
 sg13g2_a21o_1 _1850_ (.A2(_1032_),
    .A1(_1029_),
    .B1(_1034_),
    .X(_1035_));
 sg13g2_a221oi_1 _1851_ (.B2(net97),
    .C1(_1035_),
    .B1(_1030_),
    .A1(_0824_),
    .Y(_1036_),
    .A2(_1017_));
 sg13g2_a22oi_1 _1852_ (.Y(_1037_),
    .B1(_0993_),
    .B2(_1036_),
    .A2(_0912_),
    .A1(_0021_));
 sg13g2_nor3_1 _1853_ (.A(_1025_),
    .B(net56),
    .C(_1000_),
    .Y(_1038_));
 sg13g2_a21oi_1 _1854_ (.A1(net107),
    .A2(_0889_),
    .Y(_1039_),
    .B1(_0956_));
 sg13g2_a22oi_1 _1855_ (.Y(_1040_),
    .B1(_1038_),
    .B2(_1039_),
    .A2(_1014_),
    .A1(net40));
 sg13g2_inv_1 _1856_ (.Y(_1041_),
    .A(_1040_));
 sg13g2_nand3_1 _1857_ (.B(_0996_),
    .C(_1027_),
    .A(_0994_),
    .Y(_1042_));
 sg13g2_buf_1 _1858_ (.A(_0017_),
    .X(_1043_));
 sg13g2_nor2_1 _1859_ (.A(net128),
    .B(net127),
    .Y(_1044_));
 sg13g2_and4_1 _1860_ (.A(_1043_),
    .B(_0848_),
    .C(_0839_),
    .D(_1044_),
    .X(_1045_));
 sg13g2_a221oi_1 _1861_ (.B2(_0895_),
    .C1(_1045_),
    .B1(_1042_),
    .A1(_0873_),
    .Y(_1046_),
    .A2(_1014_));
 sg13g2_nor2_1 _1862_ (.A(_0862_),
    .B(net75),
    .Y(_1047_));
 sg13g2_buf_1 _1863_ (.A(_1047_),
    .X(_1048_));
 sg13g2_nand2_1 _1864_ (.Y(_1049_),
    .A(_1043_),
    .B(_1044_));
 sg13g2_nor2_2 _1865_ (.A(net75),
    .B(net71),
    .Y(_1050_));
 sg13g2_a221oi_1 _1866_ (.B2(_1050_),
    .C1(_0956_),
    .B1(_1049_),
    .A1(net39),
    .Y(_1051_),
    .A2(_0985_));
 sg13g2_a21oi_1 _1867_ (.A1(_0956_),
    .A2(_1046_),
    .Y(_1052_),
    .B1(_1051_));
 sg13g2_buf_1 _1868_ (.A(_0016_),
    .X(_1053_));
 sg13g2_nand2b_1 _1869_ (.Y(_1054_),
    .B(net129),
    .A_N(net130));
 sg13g2_nor2_1 _1870_ (.A(_0863_),
    .B(_1054_),
    .Y(_1055_));
 sg13g2_buf_1 _1871_ (.A(_1055_),
    .X(_1056_));
 sg13g2_buf_1 _1872_ (.A(net125),
    .X(_1057_));
 sg13g2_nor2_1 _1873_ (.A(net124),
    .B(net96),
    .Y(_1058_));
 sg13g2_nand4_1 _1874_ (.B(net123),
    .C(net55),
    .A(_1053_),
    .Y(_1059_),
    .D(_1058_));
 sg13g2_and3_1 _1875_ (.X(_1060_),
    .A(_0976_),
    .B(_0973_),
    .C(_0983_));
 sg13g2_nand4_1 _1876_ (.B(_0956_),
    .C(net39),
    .A(net123),
    .Y(_1061_),
    .D(_1060_));
 sg13g2_nor2b_1 _1877_ (.A(net125),
    .B_N(net127),
    .Y(_1062_));
 sg13g2_nor2b_1 _1878_ (.A(net126),
    .B_N(_0970_),
    .Y(_1063_));
 sg13g2_buf_2 _1879_ (.A(_1063_),
    .X(_1064_));
 sg13g2_nand3_1 _1880_ (.B(_1064_),
    .C(_1018_),
    .A(_1062_),
    .Y(_1065_));
 sg13g2_nor2b_2 _1881_ (.A(_0982_),
    .B_N(_0956_),
    .Y(_1066_));
 sg13g2_or3_1 _1882_ (.A(_0869_),
    .B(_1065_),
    .C(_1066_),
    .X(_1067_));
 sg13g2_nor2_1 _1883_ (.A(_0960_),
    .B(_1054_),
    .Y(_1068_));
 sg13g2_buf_1 _1884_ (.A(_1068_),
    .X(_1069_));
 sg13g2_nand3_1 _1885_ (.B(_1065_),
    .C(_1066_),
    .A(net38),
    .Y(_1070_));
 sg13g2_nand4_1 _1886_ (.B(_1061_),
    .C(_1067_),
    .A(_1059_),
    .Y(_1071_),
    .D(_1070_));
 sg13g2_nor3_1 _1887_ (.A(_1041_),
    .B(_1052_),
    .C(_1071_),
    .Y(_1072_));
 sg13g2_buf_1 _1888_ (.A(_0895_),
    .X(_1073_));
 sg13g2_a22oi_1 _1889_ (.Y(_1074_),
    .B1(_1042_),
    .B2(net54),
    .A2(_0985_),
    .A1(net39));
 sg13g2_nand2_1 _1890_ (.Y(_1075_),
    .A(_1053_),
    .B(_1058_));
 sg13g2_nor3_1 _1891_ (.A(_0956_),
    .B(_0864_),
    .C(_0822_),
    .Y(_1076_));
 sg13g2_nand2_1 _1892_ (.Y(_1077_),
    .A(_1003_),
    .B(_1004_));
 sg13g2_a221oi_1 _1893_ (.B2(_1077_),
    .C1(net123),
    .B1(_1076_),
    .A1(net55),
    .Y(_1078_),
    .A2(_1075_));
 sg13g2_nand2_1 _1894_ (.Y(_1079_),
    .A(_1074_),
    .B(_1078_));
 sg13g2_or3_1 _1895_ (.A(_1052_),
    .B(_1071_),
    .C(_1079_),
    .X(_1080_));
 sg13g2_o21ai_1 _1896_ (.B1(_1080_),
    .Y(_1081_),
    .A1(_0988_),
    .A2(_1072_));
 sg13g2_a21oi_1 _1897_ (.A1(net129),
    .A2(_0789_),
    .Y(_1082_),
    .B1(_1020_));
 sg13g2_nor4_2 _1898_ (.A(net106),
    .B(_1064_),
    .C(_0900_),
    .Y(_1083_),
    .D(_1082_));
 sg13g2_o21ai_1 _1899_ (.B1(net108),
    .Y(_1084_),
    .A1(_1020_),
    .A2(net98));
 sg13g2_or2_1 _1900_ (.X(_1085_),
    .B(_0785_),
    .A(_1043_));
 sg13g2_a21oi_1 _1901_ (.A1(_1084_),
    .A2(_1085_),
    .Y(_1086_),
    .B1(net103));
 sg13g2_o21ai_1 _1902_ (.B1(_0805_),
    .Y(_1087_),
    .A1(_0812_),
    .A2(_0787_));
 sg13g2_nor3_2 _1903_ (.A(_1083_),
    .B(_1086_),
    .C(_1087_),
    .Y(_1088_));
 sg13g2_o21ai_1 _1904_ (.B1(_1053_),
    .Y(_1089_),
    .A1(_1023_),
    .A2(_0891_));
 sg13g2_nor2_1 _1905_ (.A(_1088_),
    .B(_1089_),
    .Y(_1090_));
 sg13g2_or2_1 _1906_ (.X(_1091_),
    .B(net127),
    .A(net125));
 sg13g2_buf_1 _1907_ (.A(_1091_),
    .X(_1092_));
 sg13g2_xnor2_1 _1908_ (.Y(_1093_),
    .A(_1092_),
    .B(_1002_));
 sg13g2_xnor2_1 _1909_ (.Y(_1094_),
    .A(_1019_),
    .B(_1064_));
 sg13g2_a22oi_1 _1910_ (.Y(_1095_),
    .B1(_1069_),
    .B2(_1094_),
    .A2(_1093_),
    .A1(_0872_));
 sg13g2_and2_1 _1911_ (.A(_0970_),
    .B(net126),
    .X(_1096_));
 sg13g2_buf_1 _1912_ (.A(_1096_),
    .X(_1097_));
 sg13g2_xnor2_1 _1913_ (.Y(_1098_),
    .A(_0976_),
    .B(_1097_));
 sg13g2_nand2_1 _1914_ (.Y(_1099_),
    .A(_1048_),
    .B(_1098_));
 sg13g2_xor2_1 _1915_ (.B(net96),
    .A(_1021_),
    .X(_1100_));
 sg13g2_xor2_1 _1916_ (.B(net127),
    .A(net99),
    .X(_1101_));
 sg13g2_a221oi_1 _1917_ (.B2(_1101_),
    .C1(_0895_),
    .B1(_1050_),
    .A1(net55),
    .Y(_1102_),
    .A2(_1100_));
 sg13g2_nand3_1 _1918_ (.B(_1099_),
    .C(_1102_),
    .A(_1095_),
    .Y(_1103_));
 sg13g2_buf_1 _1919_ (.A(_1103_),
    .X(_1104_));
 sg13g2_nand2_1 _1920_ (.Y(_1105_),
    .A(_1025_),
    .B(net56));
 sg13g2_a21oi_2 _1921_ (.B1(_0891_),
    .Y(_1106_),
    .A2(_1105_),
    .A1(_0997_));
 sg13g2_nor2_1 _1922_ (.A(net96),
    .B(_1106_),
    .Y(_1107_));
 sg13g2_and2_1 _1923_ (.A(_1104_),
    .B(_1107_),
    .X(_1108_));
 sg13g2_a21o_1 _1924_ (.A2(_0973_),
    .A1(_0976_),
    .B1(_0983_),
    .X(_1109_));
 sg13g2_nand3_1 _1925_ (.B(_0985_),
    .C(_1109_),
    .A(_1048_),
    .Y(_1110_));
 sg13g2_nand2b_1 _1926_ (.Y(_1111_),
    .B(_0872_),
    .A_N(_1005_));
 sg13g2_a21oi_1 _1927_ (.A1(_1062_),
    .A2(_1064_),
    .Y(_1112_),
    .B1(_0980_));
 sg13g2_nand2b_1 _1928_ (.Y(_1113_),
    .B(_0970_),
    .A_N(net126));
 sg13g2_nor3_1 _1929_ (.A(_1019_),
    .B(_1113_),
    .C(_1018_),
    .Y(_1114_));
 sg13g2_o21ai_1 _1930_ (.B1(_1068_),
    .Y(_1115_),
    .A1(_1112_),
    .A2(_1114_));
 sg13g2_and3_1 _1931_ (.X(_1116_),
    .A(_1110_),
    .B(_1111_),
    .C(_1115_));
 sg13g2_buf_2 _1932_ (.A(_0020_),
    .X(_1117_));
 sg13g2_or3_1 _1933_ (.A(net126),
    .B(net124),
    .C(net125),
    .X(_1118_));
 sg13g2_o21ai_1 _1934_ (.B1(net124),
    .Y(_1119_),
    .A1(_0971_),
    .A2(net125));
 sg13g2_and2_1 _1935_ (.A(_1118_),
    .B(_1119_),
    .X(_1120_));
 sg13g2_nor2_1 _1936_ (.A(net99),
    .B(net127),
    .Y(_1121_));
 sg13g2_xnor2_1 _1937_ (.Y(_1122_),
    .A(net128),
    .B(_1121_));
 sg13g2_a221oi_1 _1938_ (.B2(_1050_),
    .C1(_0895_),
    .B1(_1122_),
    .A1(net55),
    .Y(_1123_),
    .A2(_1120_));
 sg13g2_and2_1 _1939_ (.A(_1117_),
    .B(_1123_),
    .X(_1124_));
 sg13g2_o21ai_1 _1940_ (.B1(_1000_),
    .Y(_1125_),
    .A1(_1025_),
    .A2(net56));
 sg13g2_a21oi_1 _1941_ (.A1(_1042_),
    .A2(_1125_),
    .Y(_1126_),
    .B1(_0891_));
 sg13g2_nor2_1 _1942_ (.A(_1117_),
    .B(_1126_),
    .Y(_1127_));
 sg13g2_nand4_1 _1943_ (.B(_1123_),
    .C(_1111_),
    .A(_1110_),
    .Y(_1128_),
    .D(_1115_));
 sg13g2_buf_1 _1944_ (.A(_1128_),
    .X(_1129_));
 sg13g2_and2_1 _1945_ (.A(_1117_),
    .B(_1126_),
    .X(_1130_));
 sg13g2_a221oi_1 _1946_ (.B2(_1129_),
    .C1(_1130_),
    .B1(_1127_),
    .A1(_1116_),
    .Y(_1131_),
    .A2(_1124_));
 sg13g2_nand4_1 _1947_ (.B(_1095_),
    .C(_1099_),
    .A(net96),
    .Y(_1132_),
    .D(_1102_));
 sg13g2_nand2_1 _1948_ (.Y(_1133_),
    .A(net96),
    .B(_1106_));
 sg13g2_a221oi_1 _1949_ (.B2(_1133_),
    .C1(_1130_),
    .B1(_1132_),
    .A1(_1116_),
    .Y(_1134_),
    .A2(_1124_));
 sg13g2_or4_1 _1950_ (.A(_1090_),
    .B(_1108_),
    .C(_1131_),
    .D(_1134_),
    .X(_1135_));
 sg13g2_inv_1 _1951_ (.Y(_1136_),
    .A(_1126_));
 sg13g2_nand4_1 _1952_ (.B(_1129_),
    .C(_1132_),
    .A(_1136_),
    .Y(_1137_),
    .D(_1133_));
 sg13g2_buf_1 _1953_ (.A(_0979_),
    .X(_1138_));
 sg13g2_inv_1 _1954_ (.Y(_1139_),
    .A(_1138_));
 sg13g2_nand3_1 _1955_ (.B(_1136_),
    .C(_1129_),
    .A(_1139_),
    .Y(_1140_));
 sg13g2_nand3_1 _1956_ (.B(_1132_),
    .C(_1133_),
    .A(_1139_),
    .Y(_1141_));
 sg13g2_nand3_1 _1957_ (.B(_1140_),
    .C(_1141_),
    .A(_1137_),
    .Y(_1142_));
 sg13g2_and4_1 _1958_ (.A(_0947_),
    .B(_1081_),
    .C(_1135_),
    .D(_1142_),
    .X(_1143_));
 sg13g2_nor3_1 _1959_ (.A(net28),
    .B(_1081_),
    .C(_1135_),
    .Y(_1144_));
 sg13g2_nor3_1 _1960_ (.A(net28),
    .B(_1081_),
    .C(_1142_),
    .Y(_1145_));
 sg13g2_nor4_1 _1961_ (.A(_1037_),
    .B(_1143_),
    .C(_1144_),
    .D(_1145_),
    .Y(_1146_));
 sg13g2_nand2_1 _1962_ (.Y(_1147_),
    .A(_1012_),
    .B(_1003_));
 sg13g2_o21ai_1 _1963_ (.B1(_1147_),
    .Y(_1148_),
    .A1(net95),
    .A2(_1012_));
 sg13g2_inv_2 _1964_ (.Y(_1149_),
    .A(net101));
 sg13g2_mux2_1 _1965_ (.A0(_1147_),
    .A1(_1148_),
    .S(_1149_),
    .X(_1150_));
 sg13g2_xnor2_1 _1966_ (.Y(_1151_),
    .A(_1021_),
    .B(_1008_));
 sg13g2_o21ai_1 _1967_ (.B1(_0994_),
    .Y(_1152_),
    .A1(net99),
    .A2(_1151_));
 sg13g2_xor2_1 _1968_ (.B(_1152_),
    .A(_1150_),
    .X(_1153_));
 sg13g2_nor2_1 _1969_ (.A(net74),
    .B(_0820_),
    .Y(_1154_));
 sg13g2_nor2_1 _1970_ (.A(net81),
    .B(net101),
    .Y(_1155_));
 sg13g2_a22oi_1 _1971_ (.Y(_1156_),
    .B1(_1155_),
    .B2(_0811_),
    .A2(_0814_),
    .A1(net101));
 sg13g2_nand2_1 _1972_ (.Y(_1157_),
    .A(net95),
    .B(_0973_));
 sg13g2_a21oi_1 _1973_ (.A1(_0964_),
    .A2(_1157_),
    .Y(_1158_),
    .B1(_0978_));
 sg13g2_o21ai_1 _1974_ (.B1(_0973_),
    .Y(_1159_),
    .A1(net95),
    .A2(_0976_));
 sg13g2_and2_1 _1975_ (.A(_0964_),
    .B(_0983_),
    .X(_1160_));
 sg13g2_nor2_1 _1976_ (.A(net74),
    .B(_0806_),
    .Y(_1161_));
 sg13g2_nand2_1 _1977_ (.Y(_1162_),
    .A(net81),
    .B(_1161_));
 sg13g2_a221oi_1 _1978_ (.B2(_1160_),
    .C1(_1162_),
    .B1(_1159_),
    .A1(net101),
    .Y(_1163_),
    .A2(_1158_));
 sg13g2_nand2_1 _1979_ (.Y(_1164_),
    .A(_1149_),
    .B(_0978_));
 sg13g2_a22oi_1 _1980_ (.Y(_1165_),
    .B1(_1163_),
    .B2(_1164_),
    .A2(_1156_),
    .A1(_1154_));
 sg13g2_xnor2_1 _1981_ (.Y(_1166_),
    .A(_1149_),
    .B(_1026_));
 sg13g2_o21ai_1 _1982_ (.B1(_0808_),
    .Y(_1167_),
    .A1(net29),
    .A2(_1166_));
 sg13g2_nand2_1 _1983_ (.Y(_1168_),
    .A(_1138_),
    .B(_1167_));
 sg13g2_nor2_1 _1984_ (.A(_1054_),
    .B(_0831_),
    .Y(_1169_));
 sg13g2_nand3_1 _1985_ (.B(_1169_),
    .C(_1166_),
    .A(_1139_),
    .Y(_1170_));
 sg13g2_nand3_1 _1986_ (.B(_1168_),
    .C(_1170_),
    .A(_1165_),
    .Y(_1171_));
 sg13g2_a21oi_1 _1987_ (.A1(_0824_),
    .A2(_1153_),
    .Y(_1172_),
    .B1(_1171_));
 sg13g2_a21o_1 _1988_ (.A2(_1129_),
    .A1(_1136_),
    .B1(_1139_),
    .X(_1173_));
 sg13g2_nor3_1 _1989_ (.A(_1088_),
    .B(_1106_),
    .C(_1089_),
    .Y(_1174_));
 sg13g2_o21ai_1 _1990_ (.B1(_1104_),
    .Y(_1175_),
    .A1(_1174_),
    .A2(_1107_));
 sg13g2_inv_1 _1991_ (.Y(_1176_),
    .A(_1057_));
 sg13g2_nand2_1 _1992_ (.Y(_1177_),
    .A(_1176_),
    .B(_1090_));
 sg13g2_a22oi_1 _1993_ (.Y(_1178_),
    .B1(_1175_),
    .B2(_1177_),
    .A2(_1173_),
    .A1(_1140_));
 sg13g2_and4_1 _1994_ (.A(_1177_),
    .B(_1140_),
    .C(_1173_),
    .D(_1175_),
    .X(_1179_));
 sg13g2_or3_1 _1995_ (.A(net28),
    .B(_1178_),
    .C(_1179_),
    .X(_1180_));
 sg13g2_nor3_1 _1996_ (.A(net96),
    .B(net78),
    .C(_0831_),
    .Y(_1181_));
 sg13g2_or3_1 _1997_ (.A(net100),
    .B(net56),
    .C(_1181_),
    .X(_1182_));
 sg13g2_o21ai_1 _1998_ (.B1(net56),
    .Y(_1183_),
    .A1(net100),
    .A2(_1181_));
 sg13g2_nand3_1 _1999_ (.B(_1182_),
    .C(_1183_),
    .A(_0824_),
    .Y(_1184_));
 sg13g2_nor3_1 _2000_ (.A(net96),
    .B(_0960_),
    .C(net71),
    .Y(_1185_));
 sg13g2_nor3_1 _2001_ (.A(_0998_),
    .B(_1097_),
    .C(_1185_),
    .Y(_1186_));
 sg13g2_o21ai_1 _2002_ (.B1(_1097_),
    .Y(_1187_),
    .A1(_0998_),
    .A2(_1185_));
 sg13g2_nand3b_1 _2003_ (.B(_1187_),
    .C(_0843_),
    .Y(_1188_),
    .A_N(_1186_));
 sg13g2_buf_1 _2004_ (.A(_1057_),
    .X(_1189_));
 sg13g2_xnor2_1 _2005_ (.Y(_1190_),
    .A(net100),
    .B(net56));
 sg13g2_o21ai_1 _2006_ (.B1(_0807_),
    .Y(_1191_),
    .A1(net29),
    .A2(_1190_));
 sg13g2_nor2_1 _2007_ (.A(net96),
    .B(_0794_),
    .Y(_1192_));
 sg13g2_nor2_1 _2008_ (.A(_0790_),
    .B(net100),
    .Y(_1193_));
 sg13g2_a221oi_1 _2009_ (.B2(net106),
    .C1(_0807_),
    .B1(_1193_),
    .A1(net100),
    .Y(_1194_),
    .A2(_0814_));
 sg13g2_a221oi_1 _2010_ (.B2(_1190_),
    .C1(_1194_),
    .B1(_1192_),
    .A1(net70),
    .Y(_1195_),
    .A2(_1191_));
 sg13g2_and3_1 _2011_ (.X(_1196_),
    .A(_1184_),
    .B(_1188_),
    .C(_1195_));
 sg13g2_nand4_1 _2012_ (.B(_0947_),
    .C(_1104_),
    .A(net70),
    .Y(_1197_),
    .D(_1174_));
 sg13g2_or3_1 _2013_ (.A(_1083_),
    .B(_1086_),
    .C(_1087_),
    .X(_1198_));
 sg13g2_inv_1 _2014_ (.Y(_1199_),
    .A(_1053_));
 sg13g2_a21oi_1 _2015_ (.A1(_0996_),
    .A2(net54),
    .Y(_1200_),
    .B1(_1199_));
 sg13g2_nand2_1 _2016_ (.Y(_1201_),
    .A(_1198_),
    .B(_1200_));
 sg13g2_nor2_1 _2017_ (.A(_0891_),
    .B(_1190_),
    .Y(_1202_));
 sg13g2_nand4_1 _2018_ (.B(_0947_),
    .C(_1201_),
    .A(net70),
    .Y(_1203_),
    .D(_1202_));
 sg13g2_nand3_1 _2019_ (.B(_1197_),
    .C(_1203_),
    .A(_1196_),
    .Y(_1204_));
 sg13g2_and3_1 _2020_ (.X(_1205_),
    .A(_1095_),
    .B(_1099_),
    .C(_1102_));
 sg13g2_buf_1 _2021_ (.A(_1205_),
    .X(_1206_));
 sg13g2_or4_1 _2022_ (.A(_1189_),
    .B(_1106_),
    .C(_1206_),
    .D(_1090_),
    .X(_1207_));
 sg13g2_a21oi_1 _2023_ (.A1(_1198_),
    .A2(_1200_),
    .Y(_1208_),
    .B1(_1176_));
 sg13g2_nor3_1 _2024_ (.A(_1189_),
    .B(_1088_),
    .C(_1089_),
    .Y(_1209_));
 sg13g2_o21ai_1 _2025_ (.B1(_1206_),
    .Y(_1210_),
    .A1(_1208_),
    .A2(_1209_));
 sg13g2_a21oi_1 _2026_ (.A1(_1207_),
    .A2(_1210_),
    .Y(_1211_),
    .B1(net28));
 sg13g2_nand2b_1 _2027_ (.Y(_1212_),
    .B(\alu_74181_i0.alu_74181_arith_inst.cn ),
    .A_N(_0019_));
 sg13g2_nand2_1 _2028_ (.Y(_1213_),
    .A(net82),
    .B(_0996_));
 sg13g2_a21oi_1 _2029_ (.A1(_0815_),
    .A2(_0973_),
    .Y(_1214_),
    .B1(net82));
 sg13g2_a221oi_1 _2030_ (.B2(_0934_),
    .C1(_1214_),
    .B1(_1002_),
    .A1(_0936_),
    .Y(_1215_),
    .A2(_1213_));
 sg13g2_nor2_1 _2031_ (.A(_0812_),
    .B(_1113_),
    .Y(_1216_));
 sg13g2_o21ai_1 _2032_ (.B1(net103),
    .Y(_1217_),
    .A1(_0940_),
    .A2(_1216_));
 sg13g2_nand3b_1 _2033_ (.B(_0803_),
    .C(_0805_),
    .Y(_1218_),
    .A_N(_1053_));
 sg13g2_nor2_1 _2034_ (.A(_0917_),
    .B(_1218_),
    .Y(_1219_));
 sg13g2_nor4_1 _2035_ (.A(_1083_),
    .B(_1086_),
    .C(_1087_),
    .D(_1219_),
    .Y(_1220_));
 sg13g2_a21o_1 _2036_ (.A2(_1073_),
    .A1(_0996_),
    .B1(_1220_),
    .X(_1221_));
 sg13g2_and2_1 _2037_ (.A(net98),
    .B(_0947_),
    .X(_1222_));
 sg13g2_nor3_1 _2038_ (.A(net98),
    .B(_1073_),
    .C(_1220_),
    .Y(_1223_));
 sg13g2_a221oi_1 _2039_ (.B2(_1222_),
    .C1(_1223_),
    .B1(_1221_),
    .A1(_1215_),
    .Y(_1224_),
    .A2(_1217_));
 sg13g2_nor2_1 _2040_ (.A(_1199_),
    .B(_0913_),
    .Y(_1225_));
 sg13g2_and2_1 _2041_ (.A(_0022_),
    .B(_0912_),
    .X(_1226_));
 sg13g2_nor4_1 _2042_ (.A(_1212_),
    .B(_1224_),
    .C(_1225_),
    .D(_1226_),
    .Y(_1227_));
 sg13g2_o21ai_1 _2043_ (.B1(_1227_),
    .Y(_1228_),
    .A1(_1204_),
    .A2(_1211_));
 sg13g2_buf_1 _2044_ (.A(_1228_),
    .X(_1229_));
 sg13g2_a221oi_1 _2045_ (.B2(_1180_),
    .C1(_1229_),
    .B1(_1172_),
    .A1(_1117_),
    .Y(_1230_),
    .A2(_0912_));
 sg13g2_nand2b_1 _2046_ (.Y(_1231_),
    .B(_1230_),
    .A_N(_1146_));
 sg13g2_a21oi_1 _2047_ (.A1(net72),
    .A2(_1009_),
    .Y(_1232_),
    .B1(_0988_));
 sg13g2_nand2b_1 _2048_ (.Y(_1233_),
    .B(_1001_),
    .A_N(_1232_));
 sg13g2_and2_1 _2049_ (.A(net72),
    .B(_1077_),
    .X(_1234_));
 sg13g2_nor2_1 _2050_ (.A(_0988_),
    .B(net72),
    .Y(_1235_));
 sg13g2_a221oi_1 _2051_ (.B2(_1234_),
    .C1(_1235_),
    .B1(_1010_),
    .A1(_1007_),
    .Y(_1236_),
    .A2(_0792_));
 sg13g2_a21oi_1 _2052_ (.A1(_0832_),
    .A2(_1233_),
    .Y(_1237_),
    .B1(_1236_));
 sg13g2_nor2b_1 _2053_ (.A(net72),
    .B_N(_1028_),
    .Y(_1238_));
 sg13g2_nand2b_1 _2054_ (.Y(_1239_),
    .B(_0958_),
    .A_N(_1028_));
 sg13g2_o21ai_1 _2055_ (.B1(_1239_),
    .Y(_1240_),
    .A1(net97),
    .A2(_1238_));
 sg13g2_a21oi_1 _2056_ (.A1(_0787_),
    .A2(_1240_),
    .Y(_1241_),
    .B1(_0839_));
 sg13g2_nor2_1 _2057_ (.A(net101),
    .B(_0978_),
    .Y(_1242_));
 sg13g2_nor4_1 _2058_ (.A(net27),
    .B(_1018_),
    .C(_1242_),
    .D(_1066_),
    .Y(_1243_));
 sg13g2_nand2_1 _2059_ (.Y(_1244_),
    .A(net97),
    .B(net102));
 sg13g2_nand3_1 _2060_ (.B(_1060_),
    .C(_1244_),
    .A(_0965_),
    .Y(_1245_));
 sg13g2_o21ai_1 _2061_ (.B1(_1245_),
    .Y(_1246_),
    .A1(_0965_),
    .A2(_1244_));
 sg13g2_o21ai_1 _2062_ (.B1(_0843_),
    .Y(_1247_),
    .A1(_1243_),
    .A2(_1246_));
 sg13g2_o21ai_1 _2063_ (.B1(_1247_),
    .Y(_1248_),
    .A1(_0831_),
    .A2(_1241_));
 sg13g2_a21oi_1 _2064_ (.A1(_0824_),
    .A2(_1237_),
    .Y(_1249_),
    .B1(_1248_));
 sg13g2_a21oi_1 _2065_ (.A1(_1136_),
    .A2(_1129_),
    .Y(_1250_),
    .B1(_1139_));
 sg13g2_o21ai_1 _2066_ (.B1(_1201_),
    .Y(_1251_),
    .A1(_1106_),
    .A2(_1206_));
 sg13g2_a221oi_1 _2067_ (.B2(_1176_),
    .C1(_1131_),
    .B1(_1251_),
    .A1(_1104_),
    .Y(_1252_),
    .A2(_1174_));
 sg13g2_a22oi_1 _2068_ (.Y(_1253_),
    .B1(_1074_),
    .B2(_1078_),
    .A2(_1040_),
    .A1(net123));
 sg13g2_nor3_1 _2069_ (.A(_1052_),
    .B(_1071_),
    .C(_1253_),
    .Y(_1254_));
 sg13g2_o21ai_1 _2070_ (.B1(_1254_),
    .Y(_1255_),
    .A1(_1250_),
    .A2(_1252_));
 sg13g2_o21ai_1 _2071_ (.B1(net97),
    .Y(_1256_),
    .A1(net55),
    .A2(_1039_));
 sg13g2_or2_1 _2072_ (.X(_1257_),
    .B(net102),
    .A(net123));
 sg13g2_o21ai_1 _2073_ (.B1(_0873_),
    .Y(_1258_),
    .A1(_1077_),
    .A2(_1257_));
 sg13g2_buf_1 _2074_ (.A(_0804_),
    .X(_1259_));
 sg13g2_buf_1 _2075_ (.A(_0812_),
    .X(_1260_));
 sg13g2_nor2_1 _2076_ (.A(net53),
    .B(net52),
    .Y(_1261_));
 sg13g2_nor2_1 _2077_ (.A(net102),
    .B(_1261_),
    .Y(_1262_));
 sg13g2_or4_1 _2078_ (.A(_0899_),
    .B(_0900_),
    .C(_1066_),
    .D(_1262_),
    .X(_1263_));
 sg13g2_nor4_1 _2079_ (.A(net99),
    .B(_0956_),
    .C(_0967_),
    .D(net100),
    .Y(_1264_));
 sg13g2_nor3_1 _2080_ (.A(net75),
    .B(net71),
    .C(_1264_),
    .Y(_1265_));
 sg13g2_a221oi_1 _2081_ (.B2(_1056_),
    .C1(_1265_),
    .B1(_1118_),
    .A1(_1069_),
    .Y(_1266_),
    .A2(_1065_));
 sg13g2_and2_1 _2082_ (.A(_1074_),
    .B(_1266_),
    .X(_1267_));
 sg13g2_nand4_1 _2083_ (.B(_1258_),
    .C(_1263_),
    .A(_1256_),
    .Y(_1268_),
    .D(_1267_));
 sg13g2_buf_1 _2084_ (.A(_1268_),
    .X(_1269_));
 sg13g2_nor3_1 _2085_ (.A(net97),
    .B(net28),
    .C(_1269_),
    .Y(_1270_));
 sg13g2_or2_1 _2086_ (.X(_1271_),
    .B(_1254_),
    .A(_1250_));
 sg13g2_nor4_1 _2087_ (.A(_0920_),
    .B(_1269_),
    .C(_1252_),
    .D(_1271_),
    .Y(_1272_));
 sg13g2_a21oi_1 _2088_ (.A1(_1255_),
    .A2(_1270_),
    .Y(_1273_),
    .B1(_1272_));
 sg13g2_nand3b_1 _2089_ (.B(_1269_),
    .C(_0947_),
    .Y(_1274_),
    .A_N(_1255_));
 sg13g2_or2_1 _2090_ (.X(_1275_),
    .B(_1271_),
    .A(_1252_));
 sg13g2_nand4_1 _2091_ (.B(_0947_),
    .C(_1269_),
    .A(_1031_),
    .Y(_1276_),
    .D(_1275_));
 sg13g2_nand4_1 _2092_ (.B(_1273_),
    .C(_1274_),
    .A(_1249_),
    .Y(_1277_),
    .D(_1276_));
 sg13g2_xor2_1 _2093_ (.B(_1277_),
    .A(_1231_),
    .X(_1278_));
 sg13g2_buf_8 _2094_ (.A(_1278_),
    .X(_1279_));
 sg13g2_mux2_1 _2095_ (.A0(_0952_),
    .A1(_0955_),
    .S(net22),
    .X(_1280_));
 sg13g2_inv_1 _2096_ (.Y(_1281_),
    .A(_0950_));
 sg13g2_nor2_1 _2097_ (.A(_0933_),
    .B(_1281_),
    .Y(_1282_));
 sg13g2_buf_1 _2098_ (.A(_0927_),
    .X(_1283_));
 sg13g2_nand2b_1 _2099_ (.Y(_1284_),
    .B(\config_regs[26] ),
    .A_N(_0928_));
 sg13g2_or2_1 _2100_ (.X(_1285_),
    .B(_1284_),
    .A(_1283_));
 sg13g2_nor2_1 _2101_ (.A(_1224_),
    .B(_1225_),
    .Y(_1286_));
 sg13g2_nand2b_1 _2102_ (.Y(_1287_),
    .B(_1286_),
    .A_N(_1212_));
 sg13g2_and3_1 _2103_ (.X(_1288_),
    .A(_1196_),
    .B(_1197_),
    .C(_1203_));
 sg13g2_a21o_1 _2104_ (.A2(_1210_),
    .A1(_1207_),
    .B1(_0920_),
    .X(_1289_));
 sg13g2_a21oi_1 _2105_ (.A1(_1288_),
    .A2(_1289_),
    .Y(_1290_),
    .B1(_1226_));
 sg13g2_xnor2_1 _2106_ (.Y(_1291_),
    .A(_1287_),
    .B(_1290_));
 sg13g2_buf_1 _2107_ (.A(_0912_),
    .X(_1292_));
 sg13g2_buf_1 _2108_ (.A(net74),
    .X(_1293_));
 sg13g2_buf_1 _2109_ (.A(net51),
    .X(_1294_));
 sg13g2_buf_1 _2110_ (.A(net79),
    .X(_1295_));
 sg13g2_buf_1 _2111_ (.A(net50),
    .X(_1296_));
 sg13g2_a22oi_1 _2112_ (.Y(_1297_),
    .B1(_0934_),
    .B2(net70),
    .A2(_1092_),
    .A1(_0814_));
 sg13g2_nand2_1 _2113_ (.Y(_1298_),
    .A(net36),
    .B(_1297_));
 sg13g2_nor2_1 _2114_ (.A(_1296_),
    .B(_1025_),
    .Y(_1299_));
 sg13g2_o21ai_1 _2115_ (.B1(_1299_),
    .Y(_1300_),
    .A1(net70),
    .A2(_0917_));
 sg13g2_nand3_1 _2116_ (.B(_1298_),
    .C(_1300_),
    .A(net37),
    .Y(_1301_));
 sg13g2_buf_1 _2117_ (.A(net80),
    .X(_1302_));
 sg13g2_buf_1 _2118_ (.A(net81),
    .X(_1303_));
 sg13g2_nand2b_1 _2119_ (.Y(_1304_),
    .B(net53),
    .A_N(_0976_));
 sg13g2_o21ai_1 _2120_ (.B1(_1304_),
    .Y(_1305_),
    .A1(_1303_),
    .A2(_1092_));
 sg13g2_buf_1 _2121_ (.A(net80),
    .X(_1306_));
 sg13g2_nor4_1 _2122_ (.A(net47),
    .B(net51),
    .C(net48),
    .D(_1025_),
    .Y(_1307_));
 sg13g2_a21o_1 _2123_ (.A2(_1305_),
    .A1(net49),
    .B1(_1307_),
    .X(_1308_));
 sg13g2_nand3b_1 _2124_ (.B(_0838_),
    .C(_1294_),
    .Y(_1309_),
    .A_N(_0022_));
 sg13g2_o21ai_1 _2125_ (.B1(_1309_),
    .Y(_1310_),
    .A1(_0911_),
    .A2(_1092_));
 sg13g2_o21ai_1 _2126_ (.B1(_0911_),
    .Y(_1311_),
    .A1(_0027_),
    .A2(_0961_));
 sg13g2_nand2_1 _2127_ (.Y(_1312_),
    .A(_1259_),
    .B(_1311_));
 sg13g2_a22oi_1 _2128_ (.Y(_1313_),
    .B1(_0792_),
    .B2(_1062_),
    .A2(_0848_),
    .A1(net37));
 sg13g2_a21oi_1 _2129_ (.A1(_1312_),
    .A2(_1313_),
    .Y(_1314_),
    .B1(net49));
 sg13g2_a221oi_1 _2130_ (.B2(_1302_),
    .C1(_1314_),
    .B1(_1310_),
    .A1(net36),
    .Y(_1315_),
    .A2(_1308_));
 sg13g2_a221oi_1 _2131_ (.B2(_1315_),
    .C1(net73),
    .B1(_1301_),
    .A1(net70),
    .Y(_1316_),
    .A2(_1292_));
 sg13g2_a21oi_1 _2132_ (.A1(net73),
    .A2(_1291_),
    .Y(_1317_),
    .B1(_1316_));
 sg13g2_mux4_1 _2133_ (.S0(_0928_),
    .A0(net70),
    .A1(_0969_),
    .A2(net111),
    .A3(_0797_),
    .S1(net94),
    .X(_1318_));
 sg13g2_a221oi_1 _2134_ (.B2(net58),
    .C1(net53),
    .B1(_0851_),
    .A1(net49),
    .Y(_1319_),
    .A2(_0838_));
 sg13g2_buf_1 _2135_ (.A(net103),
    .X(_1320_));
 sg13g2_buf_1 _2136_ (.A(net48),
    .X(_1321_));
 sg13g2_a221oi_1 _2137_ (.B2(net36),
    .C1(net37),
    .B1(_0887_),
    .A1(net69),
    .Y(_1322_),
    .A2(net35));
 sg13g2_o21ai_1 _2138_ (.B1(_0857_),
    .Y(_1323_),
    .A1(_0829_),
    .A2(net41));
 sg13g2_a22oi_1 _2139_ (.Y(_1324_),
    .B1(_1323_),
    .B2(net49),
    .A2(_0829_),
    .A1(net35));
 sg13g2_o21ai_1 _2140_ (.B1(_1324_),
    .Y(_1325_),
    .A1(_1319_),
    .A2(_1322_));
 sg13g2_nand2b_1 _2141_ (.Y(_1326_),
    .B(_1161_),
    .A_N(_0026_));
 sg13g2_o21ai_1 _2142_ (.B1(_1326_),
    .Y(_1327_),
    .A1(net50),
    .A2(_0857_));
 sg13g2_nand3_1 _2143_ (.B(net50),
    .C(_0915_),
    .A(net47),
    .Y(_1328_));
 sg13g2_o21ai_1 _2144_ (.B1(_1328_),
    .Y(_1329_),
    .A1(net49),
    .A2(_0857_));
 sg13g2_a22oi_1 _2145_ (.Y(_1330_),
    .B1(_1329_),
    .B2(net37),
    .A2(_1327_),
    .A1(net69));
 sg13g2_nand2b_1 _2146_ (.Y(_1331_),
    .B(net35),
    .A_N(_1330_));
 sg13g2_a221oi_1 _2147_ (.B2(_1331_),
    .C1(net73),
    .B1(_1325_),
    .A1(_0783_),
    .Y(_1332_),
    .A2(net25));
 sg13g2_a22oi_1 _2148_ (.Y(_1333_),
    .B1(_0932_),
    .B2(_1332_),
    .A2(_1318_),
    .A1(_0929_));
 sg13g2_o21ai_1 _2149_ (.B1(_1333_),
    .Y(_1334_),
    .A1(_1285_),
    .A2(_1317_));
 sg13g2_a21oi_1 _2150_ (.A1(_0924_),
    .A2(_1282_),
    .Y(_1335_),
    .B1(_1334_));
 sg13g2_and2_1 _2151_ (.A(_1280_),
    .B(_1335_),
    .X(_1336_));
 sg13g2_buf_1 _2152_ (.A(_1336_),
    .X(_1337_));
 sg13g2_nor2_1 _2153_ (.A(_0915_),
    .B(_0908_),
    .Y(_1338_));
 sg13g2_o21ai_1 _2154_ (.B1(_0893_),
    .Y(_1339_),
    .A1(_0783_),
    .A2(_1338_));
 sg13g2_or3_1 _2155_ (.A(_0023_),
    .B(_0893_),
    .C(_0908_),
    .X(_1340_));
 sg13g2_buf_1 _2156_ (.A(_1340_),
    .X(_1341_));
 sg13g2_buf_1 _2157_ (.A(\alu_74181_i1.alu_74181_arith_inst.b[2] ),
    .X(_1342_));
 sg13g2_buf_1 _2158_ (.A(_1342_),
    .X(_1343_));
 sg13g2_buf_1 _2159_ (.A(net93),
    .X(_1344_));
 sg13g2_nor2b_1 _2160_ (.A(net131),
    .B_N(_0795_),
    .Y(_1345_));
 sg13g2_nand2_1 _2161_ (.Y(_1346_),
    .A(_1345_),
    .B(_0903_));
 sg13g2_nand3_1 _2162_ (.B(net38),
    .C(_1346_),
    .A(net68),
    .Y(_1347_));
 sg13g2_inv_2 _2163_ (.Y(_1348_),
    .A(net93));
 sg13g2_or4_1 _2164_ (.A(net105),
    .B(net104),
    .C(_0782_),
    .D(net109),
    .X(_1349_));
 sg13g2_nand3_1 _2165_ (.B(net40),
    .C(_1349_),
    .A(_1348_),
    .Y(_1350_));
 sg13g2_a22oi_1 _2166_ (.Y(_1351_),
    .B1(net131),
    .B2(_0795_),
    .A2(net104),
    .A1(net105));
 sg13g2_buf_1 _2167_ (.A(_1351_),
    .X(_1352_));
 sg13g2_inv_1 _2168_ (.Y(_1353_),
    .A(_1352_));
 sg13g2_buf_1 _2169_ (.A(\alu_74181_i1.a[2] ),
    .X(_1354_));
 sg13g2_buf_1 _2170_ (.A(_1354_),
    .X(_1355_));
 sg13g2_a221oi_1 _2171_ (.B2(net39),
    .C1(net92),
    .B1(_1353_),
    .A1(net54),
    .Y(_1356_),
    .A2(_0886_));
 sg13g2_nand3_1 _2172_ (.B(_1350_),
    .C(_1356_),
    .A(_1347_),
    .Y(_1357_));
 sg13g2_buf_1 _2173_ (.A(net92),
    .X(_1358_));
 sg13g2_nand3_1 _2174_ (.B(net39),
    .C(_1352_),
    .A(net93),
    .Y(_1359_));
 sg13g2_nand4_1 _2175_ (.B(net54),
    .C(_0885_),
    .A(_1348_),
    .Y(_1360_),
    .D(net83));
 sg13g2_and2_1 _2176_ (.A(_1345_),
    .B(_0903_),
    .X(_1361_));
 sg13g2_nor4_2 _2177_ (.A(net105),
    .B(net104),
    .C(net131),
    .Y(_1362_),
    .D(_0795_));
 sg13g2_a22oi_1 _2178_ (.Y(_1363_),
    .B1(_1362_),
    .B2(net40),
    .A2(_1361_),
    .A1(net38));
 sg13g2_nand4_1 _2179_ (.B(_1359_),
    .C(_1360_),
    .A(net67),
    .Y(_1364_),
    .D(_1363_));
 sg13g2_a221oi_1 _2180_ (.B2(net40),
    .C1(_1348_),
    .B1(_1362_),
    .A1(net54),
    .Y(_1365_),
    .A2(_0886_));
 sg13g2_a221oi_1 _2181_ (.B2(net39),
    .C1(net93),
    .B1(_1353_),
    .A1(net38),
    .Y(_1366_),
    .A2(_1361_));
 sg13g2_nor2_1 _2182_ (.A(_0825_),
    .B(net111),
    .Y(_1367_));
 sg13g2_xnor2_1 _2183_ (.Y(_1368_),
    .A(_1355_),
    .B(_1367_));
 sg13g2_nor2_1 _2184_ (.A(net77),
    .B(net84),
    .Y(_1369_));
 sg13g2_xnor2_1 _2185_ (.Y(_1370_),
    .A(net93),
    .B(_1369_));
 sg13g2_a22oi_1 _2186_ (.Y(_1371_),
    .B1(_1370_),
    .B2(_1050_),
    .A2(_1368_),
    .A1(net55));
 sg13g2_o21ai_1 _2187_ (.B1(_1371_),
    .Y(_1372_),
    .A1(_1365_),
    .A2(_1366_));
 sg13g2_a21oi_1 _2188_ (.A1(_1357_),
    .A2(_1364_),
    .Y(_1373_),
    .B1(_1372_));
 sg13g2_inv_1 _2189_ (.Y(_1374_),
    .A(_1373_));
 sg13g2_a21o_1 _2190_ (.A2(_1341_),
    .A1(_1339_),
    .B1(_1374_),
    .X(_1375_));
 sg13g2_nand3_1 _2191_ (.B(_1341_),
    .C(_1374_),
    .A(_1339_),
    .Y(_1376_));
 sg13g2_mux2_1 _2192_ (.A0(net67),
    .A1(_1346_),
    .S(_0840_),
    .X(_1377_));
 sg13g2_nor3_1 _2193_ (.A(net68),
    .B(net27),
    .C(_1346_),
    .Y(_1378_));
 sg13g2_a21oi_1 _2194_ (.A1(net68),
    .A2(_1377_),
    .Y(_1379_),
    .B1(_1378_));
 sg13g2_o21ai_1 _2195_ (.B1(net109),
    .Y(_1380_),
    .A1(_0960_),
    .A2(net71));
 sg13g2_xnor2_1 _2196_ (.Y(_1381_),
    .A(net76),
    .B(_1380_));
 sg13g2_a21oi_1 _2197_ (.A1(net77),
    .A2(_1381_),
    .Y(_1382_),
    .B1(_0851_));
 sg13g2_xnor2_1 _2198_ (.Y(_1383_),
    .A(_1379_),
    .B(_1382_));
 sg13g2_nand2_1 _2199_ (.Y(_1384_),
    .A(_0843_),
    .B(_1383_));
 sg13g2_nor2_1 _2200_ (.A(net109),
    .B(net83),
    .Y(_1385_));
 sg13g2_a21oi_1 _2201_ (.A1(_0796_),
    .A2(net83),
    .Y(_1386_),
    .B1(_0829_));
 sg13g2_nor3_1 _2202_ (.A(_1348_),
    .B(_1385_),
    .C(_1386_),
    .Y(_1387_));
 sg13g2_o21ai_1 _2203_ (.B1(_1348_),
    .Y(_1388_),
    .A1(_1385_),
    .A2(_1386_));
 sg13g2_nor2b_1 _2204_ (.A(_1387_),
    .B_N(_1388_),
    .Y(_1389_));
 sg13g2_o21ai_1 _2205_ (.B1(net41),
    .Y(_1390_),
    .A1(net29),
    .A2(_1389_));
 sg13g2_a21oi_1 _2206_ (.A1(_1007_),
    .A2(_0792_),
    .Y(_1391_),
    .B1(_0796_));
 sg13g2_xnor2_1 _2207_ (.Y(_1392_),
    .A(_0825_),
    .B(_1391_));
 sg13g2_o21ai_1 _2208_ (.B1(_0885_),
    .Y(_1393_),
    .A1(net77),
    .A2(_1392_));
 sg13g2_a21oi_1 _2209_ (.A1(_1007_),
    .A2(_0792_),
    .Y(_1394_),
    .B1(_1349_));
 sg13g2_nor3_1 _2210_ (.A(net92),
    .B(net78),
    .C(_0831_),
    .Y(_1395_));
 sg13g2_nor3_1 _2211_ (.A(net68),
    .B(_1394_),
    .C(_1395_),
    .Y(_1396_));
 sg13g2_a21oi_1 _2212_ (.A1(net68),
    .A2(_1394_),
    .Y(_1397_),
    .B1(_1396_));
 sg13g2_xor2_1 _2213_ (.B(_1397_),
    .A(_1393_),
    .X(_1398_));
 sg13g2_nor2_1 _2214_ (.A(net67),
    .B(net29),
    .Y(_1399_));
 sg13g2_nor2_1 _2215_ (.A(net81),
    .B(_1344_),
    .Y(_1400_));
 sg13g2_a221oi_1 _2216_ (.B2(net106),
    .C1(_0807_),
    .B1(_1400_),
    .A1(_1344_),
    .Y(_1401_),
    .A2(_0814_));
 sg13g2_a21o_1 _2217_ (.A2(_1399_),
    .A1(_1389_),
    .B1(_1401_),
    .X(_1402_));
 sg13g2_a221oi_1 _2218_ (.B2(_0824_),
    .C1(_1402_),
    .B1(_1398_),
    .A1(net67),
    .Y(_1403_),
    .A2(_1390_));
 sg13g2_nand3_1 _2219_ (.B(_1384_),
    .C(_1403_),
    .A(_0028_),
    .Y(_1404_));
 sg13g2_a21oi_1 _2220_ (.A1(_1375_),
    .A2(_1376_),
    .Y(_1405_),
    .B1(_1404_));
 sg13g2_inv_1 _2221_ (.Y(_1406_),
    .A(_0028_));
 sg13g2_and2_1 _2222_ (.A(_1384_),
    .B(_1403_),
    .X(_1407_));
 sg13g2_and4_1 _2223_ (.A(_1406_),
    .B(_1407_),
    .C(_1375_),
    .D(_1376_),
    .X(_1408_));
 sg13g2_nand3_1 _2224_ (.B(_1384_),
    .C(_1403_),
    .A(net28),
    .Y(_1409_));
 sg13g2_o21ai_1 _2225_ (.B1(_1409_),
    .Y(_1410_),
    .A1(_1406_),
    .A2(_0913_));
 sg13g2_nor3_2 _2226_ (.A(_1405_),
    .B(_1408_),
    .C(_1410_),
    .Y(_1411_));
 sg13g2_nand2_1 _2227_ (.Y(_1412_),
    .A(_0924_),
    .B(_0951_));
 sg13g2_or3_1 _2228_ (.A(net22),
    .B(_1411_),
    .C(_1412_),
    .X(_1413_));
 sg13g2_nand3_1 _2229_ (.B(net22),
    .C(_1411_),
    .A(_0954_),
    .Y(_1414_));
 sg13g2_mux4_1 _2230_ (.S0(_0928_),
    .A0(net95),
    .A1(net101),
    .A2(_1358_),
    .A3(net68),
    .S1(net94),
    .X(_1415_));
 sg13g2_a21oi_1 _2231_ (.A1(_0924_),
    .A2(_1281_),
    .Y(_1416_),
    .B1(_0933_));
 sg13g2_nor2_1 _2232_ (.A(_0927_),
    .B(_0925_),
    .Y(_1417_));
 sg13g2_nand2b_1 _2233_ (.Y(_1418_),
    .B(_1417_),
    .A_N(_1229_));
 sg13g2_nand2_1 _2234_ (.Y(_1419_),
    .A(_1229_),
    .B(_1417_));
 sg13g2_a22oi_1 _2235_ (.Y(_1420_),
    .B1(_1172_),
    .B2(_1180_),
    .A2(_1292_),
    .A1(_1117_));
 sg13g2_mux2_1 _2236_ (.A0(_1418_),
    .A1(_1419_),
    .S(_1420_),
    .X(_1421_));
 sg13g2_nor2_1 _2237_ (.A(net103),
    .B(net79),
    .Y(_1422_));
 sg13g2_nor2_1 _2238_ (.A(net58),
    .B(net68),
    .Y(_1423_));
 sg13g2_o21ai_1 _2239_ (.B1(net67),
    .Y(_1424_),
    .A1(_1422_),
    .A2(_1423_));
 sg13g2_o21ai_1 _2240_ (.B1(_0814_),
    .Y(_1425_),
    .A1(net50),
    .A2(net67));
 sg13g2_a21o_1 _2241_ (.A2(_1425_),
    .A1(_1424_),
    .B1(net51),
    .X(_1426_));
 sg13g2_nor2_1 _2242_ (.A(net92),
    .B(_1343_),
    .Y(_1427_));
 sg13g2_nand2_1 _2243_ (.Y(_1428_),
    .A(net35),
    .B(_1427_));
 sg13g2_nand4_1 _2244_ (.B(net58),
    .C(net67),
    .A(net51),
    .Y(_1429_),
    .D(net68));
 sg13g2_nor2b_1 _2245_ (.A(net92),
    .B_N(net93),
    .Y(_1430_));
 sg13g2_o21ai_1 _2246_ (.B1(net47),
    .Y(_1431_),
    .A1(_1261_),
    .A2(_1430_));
 sg13g2_nand4_1 _2247_ (.B(_1428_),
    .C(_1429_),
    .A(_1426_),
    .Y(_1432_),
    .D(_1431_));
 sg13g2_nand2b_1 _2248_ (.Y(_1433_),
    .B(_1354_),
    .A_N(_1342_));
 sg13g2_buf_1 _2249_ (.A(_1433_),
    .X(_1434_));
 sg13g2_nor2_1 _2250_ (.A(net79),
    .B(_1434_),
    .Y(_1435_));
 sg13g2_a21oi_1 _2251_ (.A1(net50),
    .A2(_1406_),
    .Y(_1436_),
    .B1(_1435_));
 sg13g2_nor2_1 _2252_ (.A(net78),
    .B(_1436_),
    .Y(_1437_));
 sg13g2_nor3_1 _2253_ (.A(net58),
    .B(_0029_),
    .C(_0862_),
    .Y(_1438_));
 sg13g2_o21ai_1 _2254_ (.B1(net35),
    .Y(_1439_),
    .A1(_1437_),
    .A2(_1438_));
 sg13g2_a221oi_1 _2255_ (.B2(_1439_),
    .C1(_0926_),
    .B1(_1432_),
    .A1(_1358_),
    .Y(_1440_),
    .A2(net25));
 sg13g2_nor2_1 _2256_ (.A(net80),
    .B(_0820_),
    .Y(_1441_));
 sg13g2_inv_1 _2257_ (.Y(_1442_),
    .A(_1441_));
 sg13g2_nand3_1 _2258_ (.B(_1295_),
    .C(net95),
    .A(net47),
    .Y(_1443_));
 sg13g2_o21ai_1 _2259_ (.B1(_1443_),
    .Y(_1444_),
    .A1(net95),
    .A2(_1442_));
 sg13g2_nor2_1 _2260_ (.A(_1149_),
    .B(_0889_),
    .Y(_1445_));
 sg13g2_o21ai_1 _2261_ (.B1(_0911_),
    .Y(_1446_),
    .A1(_0030_),
    .A2(_0961_));
 sg13g2_a22oi_1 _2262_ (.Y(_1447_),
    .B1(_1446_),
    .B2(_0846_),
    .A2(_1445_),
    .A1(_1444_));
 sg13g2_nand2_1 _2263_ (.Y(_1448_),
    .A(net80),
    .B(_0940_));
 sg13g2_nand2_1 _2264_ (.Y(_1449_),
    .A(_1448_),
    .B(_0983_));
 sg13g2_nand2_1 _2265_ (.Y(_1450_),
    .A(net74),
    .B(_0848_));
 sg13g2_nand2_1 _2266_ (.Y(_1451_),
    .A(_1450_),
    .B(net41));
 sg13g2_a22oi_1 _2267_ (.Y(_1452_),
    .B1(_1451_),
    .B2(net69),
    .A2(_1449_),
    .A1(_0937_));
 sg13g2_nand2_1 _2268_ (.Y(_1453_),
    .A(net52),
    .B(_1027_));
 sg13g2_a21oi_1 _2269_ (.A1(net57),
    .A2(_0980_),
    .Y(_1454_),
    .B1(net69));
 sg13g2_a221oi_1 _2270_ (.B2(_1259_),
    .C1(_1454_),
    .B1(_1453_),
    .A1(_1321_),
    .Y(_1455_),
    .A2(_1004_));
 sg13g2_nand2_1 _2271_ (.Y(_1456_),
    .A(net103),
    .B(_0848_));
 sg13g2_nor2_1 _2272_ (.A(net101),
    .B(_0911_),
    .Y(_1457_));
 sg13g2_nor2_1 _2273_ (.A(_1117_),
    .B(net57),
    .Y(_1458_));
 sg13g2_o21ai_1 _2274_ (.B1(_1302_),
    .Y(_0153_),
    .A1(_1457_),
    .A2(_1458_));
 sg13g2_nand2_1 _2275_ (.Y(_0154_),
    .A(_1456_),
    .B(_0153_));
 sg13g2_a22oi_1 _2276_ (.Y(_0155_),
    .B1(_0154_),
    .B2(net37),
    .A2(_1455_),
    .A1(_1452_));
 sg13g2_a22oi_1 _2277_ (.Y(_0156_),
    .B1(_1447_),
    .B2(_0155_),
    .A2(net25),
    .A1(net95));
 sg13g2_nor2_1 _2278_ (.A(_0927_),
    .B(net73),
    .Y(_0157_));
 sg13g2_a22oi_1 _2279_ (.Y(_0158_),
    .B1(_0156_),
    .B2(_0157_),
    .A2(_1440_),
    .A1(net94));
 sg13g2_a21oi_1 _2280_ (.A1(_1421_),
    .A2(_0158_),
    .Y(_0159_),
    .B1(_1284_));
 sg13g2_a221oi_1 _2281_ (.B2(_1411_),
    .C1(_0159_),
    .B1(_1416_),
    .A1(_0929_),
    .Y(_0160_),
    .A2(_1415_));
 sg13g2_and3_1 _2282_ (.X(_0161_),
    .A(_1413_),
    .B(_1414_),
    .C(_0160_));
 sg13g2_buf_8 _2283_ (.A(_0161_),
    .X(_0162_));
 sg13g2_mux4_1 _2284_ (.S0(net94),
    .A0(net98),
    .A1(net76),
    .A2(net99),
    .A3(net77),
    .S1(_0928_),
    .X(_0163_));
 sg13g2_xnor2_1 _2285_ (.Y(_0164_),
    .A(\alu_74181_i0.alu_74181_arith_inst.cn ),
    .B(_1286_));
 sg13g2_o21ai_1 _2286_ (.B1(net80),
    .Y(_0165_),
    .A1(net79),
    .A2(net99));
 sg13g2_a22oi_1 _2287_ (.Y(_0166_),
    .B1(_1097_),
    .B2(_0937_),
    .A2(_1002_),
    .A1(net48));
 sg13g2_nand4_1 _2288_ (.B(_0864_),
    .C(_0165_),
    .A(net51),
    .Y(_0167_),
    .D(_0166_));
 sg13g2_nand2_1 _2289_ (.Y(_0168_),
    .A(net74),
    .B(net79));
 sg13g2_a21oi_1 _2290_ (.A1(_0168_),
    .A2(net41),
    .Y(_0169_),
    .B1(net48));
 sg13g2_nor2_1 _2291_ (.A(_1043_),
    .B(_1162_),
    .Y(_0170_));
 sg13g2_o21ai_1 _2292_ (.B1(net69),
    .Y(_0171_),
    .A1(_0169_),
    .A2(_0170_));
 sg13g2_nor2_1 _2293_ (.A(net69),
    .B(_1218_),
    .Y(_0172_));
 sg13g2_nor3_1 _2294_ (.A(net79),
    .B(_0862_),
    .C(_1113_),
    .Y(_0173_));
 sg13g2_o21ai_1 _2295_ (.B1(net48),
    .Y(_0174_),
    .A1(_0172_),
    .A2(_0173_));
 sg13g2_nand3_1 _2296_ (.B(_1002_),
    .C(_1422_),
    .A(net52),
    .Y(_0175_));
 sg13g2_and4_1 _2297_ (.A(_0167_),
    .B(_0171_),
    .C(_0174_),
    .D(_0175_),
    .X(_0176_));
 sg13g2_a21o_1 _2298_ (.A2(net98),
    .A1(_0936_),
    .B1(_1002_),
    .X(_0177_));
 sg13g2_a22oi_1 _2299_ (.Y(_0178_),
    .B1(_0177_),
    .B2(net47),
    .A2(_0996_),
    .A1(_0846_));
 sg13g2_nor2_1 _2300_ (.A(net48),
    .B(_0178_),
    .Y(_0179_));
 sg13g2_nor2_1 _2301_ (.A(_0973_),
    .B(_0963_),
    .Y(_0180_));
 sg13g2_o21ai_1 _2302_ (.B1(_1296_),
    .Y(_0181_),
    .A1(_0179_),
    .A2(_0180_));
 sg13g2_a22oi_1 _2303_ (.Y(_0182_),
    .B1(_0176_),
    .B2(_0181_),
    .A2(net25),
    .A1(net98));
 sg13g2_nand2_1 _2304_ (.Y(_0183_),
    .A(_0925_),
    .B(_0182_));
 sg13g2_o21ai_1 _2305_ (.B1(_0183_),
    .Y(_0184_),
    .A1(_0925_),
    .A2(_0164_));
 sg13g2_a22oi_1 _2306_ (.Y(_0185_),
    .B1(_0903_),
    .B2(_1320_),
    .A2(_0828_),
    .A1(net51));
 sg13g2_nor3_1 _2307_ (.A(_0817_),
    .B(net76),
    .C(net77),
    .Y(_0186_));
 sg13g2_a21oi_1 _2308_ (.A1(net47),
    .A2(_0894_),
    .Y(_0187_),
    .B1(_0186_));
 sg13g2_nand2b_1 _2309_ (.Y(_0188_),
    .B(_0187_),
    .A_N(_0168_));
 sg13g2_o21ai_1 _2310_ (.B1(_0188_),
    .Y(_0189_),
    .A1(net36),
    .A2(_0185_));
 sg13g2_nand2_1 _2311_ (.Y(_0190_),
    .A(net47),
    .B(_0835_));
 sg13g2_a21oi_1 _2312_ (.A1(net50),
    .A2(_0853_),
    .Y(_0191_),
    .B1(_0190_));
 sg13g2_nand2_1 _2313_ (.Y(_0192_),
    .A(net58),
    .B(_0836_));
 sg13g2_a21oi_1 _2314_ (.A1(net69),
    .A2(_0192_),
    .Y(_0193_),
    .B1(_1422_));
 sg13g2_nor3_1 _2315_ (.A(net51),
    .B(_0828_),
    .C(_1441_),
    .Y(_0194_));
 sg13g2_a21oi_1 _2316_ (.A1(net37),
    .A2(_0193_),
    .Y(_0195_),
    .B1(_0194_));
 sg13g2_nor3_1 _2317_ (.A(net35),
    .B(_0191_),
    .C(_0195_),
    .Y(_0196_));
 sg13g2_a21oi_1 _2318_ (.A1(net35),
    .A2(_0189_),
    .Y(_0197_),
    .B1(_0196_));
 sg13g2_o21ai_1 _2319_ (.B1(_0911_),
    .Y(_0198_),
    .A1(_0025_),
    .A2(net57));
 sg13g2_inv_1 _2320_ (.Y(_0199_),
    .A(_0198_));
 sg13g2_o21ai_1 _2321_ (.B1(_1450_),
    .Y(_0200_),
    .A1(net37),
    .A2(_0199_));
 sg13g2_nor2_1 _2322_ (.A(_1162_),
    .B(_0836_),
    .Y(_0201_));
 sg13g2_nor3_1 _2323_ (.A(net53),
    .B(_0835_),
    .C(_0911_),
    .Y(_0202_));
 sg13g2_or3_1 _2324_ (.A(net69),
    .B(_0201_),
    .C(_0202_),
    .X(_0203_));
 sg13g2_o21ai_1 _2325_ (.B1(_0203_),
    .Y(_0204_),
    .A1(net49),
    .A2(_0200_));
 sg13g2_a221oi_1 _2326_ (.B2(_0204_),
    .C1(net73),
    .B1(_0197_),
    .A1(_0853_),
    .Y(_0205_),
    .A2(net25));
 sg13g2_mux2_1 _2327_ (.A0(_0184_),
    .A1(_0205_),
    .S(net94),
    .X(_0206_));
 sg13g2_a22oi_1 _2328_ (.Y(_0207_),
    .B1(_0206_),
    .B2(_0930_),
    .A2(_0163_),
    .A1(_0929_));
 sg13g2_inv_1 _2329_ (.Y(_0208_),
    .A(_1282_));
 sg13g2_inv_1 _2330_ (.Y(_0209_),
    .A(_0951_));
 sg13g2_mux2_1 _2331_ (.A0(_0208_),
    .A1(_0209_),
    .S(_1279_),
    .X(_0210_));
 sg13g2_and2_1 _2332_ (.A(_0207_),
    .B(_0210_),
    .X(_0211_));
 sg13g2_buf_1 _2333_ (.A(_0211_),
    .X(_0212_));
 sg13g2_nor2_1 _2334_ (.A(_0162_),
    .B(net19),
    .Y(_0213_));
 sg13g2_nand2_1 _2335_ (.Y(_0214_),
    .A(_0207_),
    .B(_0210_));
 sg13g2_buf_1 _2336_ (.A(_0214_),
    .X(_0215_));
 sg13g2_xnor2_1 _2337_ (.Y(_0216_),
    .A(_0162_),
    .B(net18));
 sg13g2_nand3_1 _2338_ (.B(_1281_),
    .C(_1411_),
    .A(_0924_),
    .Y(_0217_));
 sg13g2_buf_2 _2339_ (.A(_0004_),
    .X(_0218_));
 sg13g2_buf_1 _2340_ (.A(\alu_74181_i1.alu_74181_arith_inst.b[3] ),
    .X(_0219_));
 sg13g2_buf_1 _2341_ (.A(_0219_),
    .X(_0220_));
 sg13g2_inv_1 _2342_ (.Y(_0221_),
    .A(_0025_));
 sg13g2_or2_1 _2343_ (.X(_0222_),
    .B(_1342_),
    .A(_0795_));
 sg13g2_buf_1 _2344_ (.A(_0222_),
    .X(_0223_));
 sg13g2_nor2_1 _2345_ (.A(_0221_),
    .B(_0223_),
    .Y(_0224_));
 sg13g2_xnor2_1 _2346_ (.Y(_0225_),
    .A(net91),
    .B(_0224_));
 sg13g2_inv_1 _2347_ (.Y(_0226_),
    .A(_1355_));
 sg13g2_nand3_1 _2348_ (.B(_0894_),
    .C(_0226_),
    .A(_0829_),
    .Y(_0227_));
 sg13g2_nor2_1 _2349_ (.A(_0880_),
    .B(_0227_),
    .Y(_0228_));
 sg13g2_buf_1 _2350_ (.A(\alu_74181_i1.a[3] ),
    .X(_0229_));
 sg13g2_buf_1 _2351_ (.A(_0229_),
    .X(_0230_));
 sg13g2_a22oi_1 _2352_ (.Y(_0231_),
    .B1(_0228_),
    .B2(net90),
    .A2(_0225_),
    .A1(_1050_));
 sg13g2_nand2_1 _2353_ (.Y(_0232_),
    .A(net92),
    .B(_1343_));
 sg13g2_and2_1 _2354_ (.A(_1352_),
    .B(_0232_),
    .X(_0233_));
 sg13g2_inv_1 _2355_ (.Y(_0234_),
    .A(_0229_));
 sg13g2_nor3_1 _2356_ (.A(_0234_),
    .B(_0862_),
    .C(net75),
    .Y(_0235_));
 sg13g2_nand3_1 _2357_ (.B(net83),
    .C(_1434_),
    .A(_0885_),
    .Y(_0236_));
 sg13g2_and4_1 _2358_ (.A(_0848_),
    .B(_1007_),
    .C(_1362_),
    .D(_1427_),
    .X(_0237_));
 sg13g2_a221oi_1 _2359_ (.B2(net54),
    .C1(_0237_),
    .B1(_0236_),
    .A1(_0233_),
    .Y(_0238_),
    .A2(_0235_));
 sg13g2_nand2b_1 _2360_ (.Y(_0239_),
    .B(_1342_),
    .A_N(_1354_));
 sg13g2_nor4_2 _2361_ (.A(net105),
    .B(_0855_),
    .C(_0857_),
    .Y(_0240_),
    .D(_0239_));
 sg13g2_nand2_1 _2362_ (.Y(_0241_),
    .A(_1352_),
    .B(_0232_));
 sg13g2_a221oi_1 _2363_ (.B2(net39),
    .C1(net91),
    .B1(_0241_),
    .A1(net38),
    .Y(_0242_),
    .A2(_0240_));
 sg13g2_a21o_1 _2364_ (.A2(_0238_),
    .A1(net91),
    .B1(_0242_),
    .X(_0243_));
 sg13g2_buf_1 _2365_ (.A(_0234_),
    .X(_0244_));
 sg13g2_nor2_1 _2366_ (.A(net66),
    .B(_0219_),
    .Y(_0245_));
 sg13g2_and3_1 _2367_ (.X(_0246_),
    .A(_0885_),
    .B(net83),
    .C(_1434_));
 sg13g2_mux2_1 _2368_ (.A0(net66),
    .A1(_0245_),
    .S(_0246_),
    .X(_0247_));
 sg13g2_nand2_1 _2369_ (.Y(_0248_),
    .A(net54),
    .B(_0247_));
 sg13g2_nand3_1 _2370_ (.B(_0243_),
    .C(_0248_),
    .A(_0231_),
    .Y(_0249_));
 sg13g2_buf_1 _2371_ (.A(_0249_),
    .X(_0250_));
 sg13g2_a21oi_1 _2372_ (.A1(net38),
    .A2(_0240_),
    .Y(_0251_),
    .B1(_0237_));
 sg13g2_inv_2 _2373_ (.Y(_0252_),
    .A(_0219_));
 sg13g2_nand2_1 _2374_ (.Y(_0253_),
    .A(_1362_),
    .B(_1427_));
 sg13g2_nand3_1 _2375_ (.B(net40),
    .C(_0253_),
    .A(_0252_),
    .Y(_0254_));
 sg13g2_nand3_1 _2376_ (.B(_0903_),
    .C(_1430_),
    .A(_1345_),
    .Y(_0255_));
 sg13g2_nand3_1 _2377_ (.B(net38),
    .C(_0255_),
    .A(net91),
    .Y(_0256_));
 sg13g2_a22oi_1 _2378_ (.Y(_0257_),
    .B1(_0241_),
    .B2(net39),
    .A2(_0227_),
    .A1(net55));
 sg13g2_and4_1 _2379_ (.A(net66),
    .B(_0254_),
    .C(_0256_),
    .D(_0257_),
    .X(_0258_));
 sg13g2_a21oi_2 _2380_ (.B1(_0258_),
    .Y(_0259_),
    .A2(_0251_),
    .A1(net90));
 sg13g2_nor3_2 _2381_ (.A(_0226_),
    .B(_1364_),
    .C(_1372_),
    .Y(_0260_));
 sg13g2_nor4_1 _2382_ (.A(_0218_),
    .B(_0250_),
    .C(_0259_),
    .D(_0260_),
    .Y(_0261_));
 sg13g2_nor2_1 _2383_ (.A(_0250_),
    .B(_0259_),
    .Y(_0262_));
 sg13g2_nor2_1 _2384_ (.A(_0218_),
    .B(_0262_),
    .Y(_0263_));
 sg13g2_xnor2_1 _2385_ (.Y(_0264_),
    .A(_1406_),
    .B(_1373_));
 sg13g2_a21oi_1 _2386_ (.A1(_1339_),
    .A2(_1341_),
    .Y(_0265_),
    .B1(_0264_));
 sg13g2_mux2_1 _2387_ (.A0(_0261_),
    .A1(_0263_),
    .S(_0265_),
    .X(_0266_));
 sg13g2_nand2b_1 _2388_ (.Y(_0267_),
    .B(_0260_),
    .A_N(_0262_));
 sg13g2_o21ai_1 _2389_ (.B1(_0947_),
    .Y(_0268_),
    .A1(_0218_),
    .A2(_0267_));
 sg13g2_o21ai_1 _2390_ (.B1(_0239_),
    .Y(_0269_),
    .A1(_1385_),
    .A2(_1386_));
 sg13g2_a21oi_1 _2391_ (.A1(_1434_),
    .A2(_0269_),
    .Y(_0270_),
    .B1(_0220_));
 sg13g2_buf_1 _2392_ (.A(_0220_),
    .X(_0271_));
 sg13g2_and3_1 _2393_ (.X(_0272_),
    .A(net65),
    .B(_1434_),
    .C(_0269_));
 sg13g2_o21ai_1 _2394_ (.B1(_1169_),
    .Y(_0273_),
    .A1(_0270_),
    .A2(_0272_));
 sg13g2_nor2_1 _2395_ (.A(net66),
    .B(_1154_),
    .Y(_0274_));
 sg13g2_nand3_1 _2396_ (.B(_1434_),
    .C(_0269_),
    .A(net65),
    .Y(_0275_));
 sg13g2_nand3b_1 _2397_ (.B(_0275_),
    .C(_1169_),
    .Y(_0276_),
    .A_N(_0270_));
 sg13g2_a22oi_1 _2398_ (.Y(_0277_),
    .B1(_0276_),
    .B2(net66),
    .A2(_0274_),
    .A1(_0273_));
 sg13g2_o21ai_1 _2399_ (.B1(_0223_),
    .Y(_0278_),
    .A1(_0960_),
    .A2(net71));
 sg13g2_nor2_1 _2400_ (.A(net76),
    .B(_0857_),
    .Y(_0279_));
 sg13g2_a22oi_1 _2401_ (.Y(_0280_),
    .B1(_0279_),
    .B2(_0840_),
    .A2(_0278_),
    .A1(net76));
 sg13g2_o21ai_1 _2402_ (.B1(net93),
    .Y(_0281_),
    .A1(net57),
    .A2(net71));
 sg13g2_a21oi_1 _2403_ (.A1(_0851_),
    .A2(_0281_),
    .Y(_0282_),
    .B1(net92));
 sg13g2_o21ai_1 _2404_ (.B1(_0282_),
    .Y(_0283_),
    .A1(_0855_),
    .A2(_0280_));
 sg13g2_nor2b_1 _2405_ (.A(_0836_),
    .B_N(_1380_),
    .Y(_0284_));
 sg13g2_or3_1 _2406_ (.A(net93),
    .B(_0851_),
    .C(_0284_),
    .X(_0285_));
 sg13g2_buf_1 _2407_ (.A(_0285_),
    .X(_0286_));
 sg13g2_nor3_1 _2408_ (.A(_0229_),
    .B(net57),
    .C(net71),
    .Y(_0287_));
 sg13g2_a21oi_1 _2409_ (.A1(_0840_),
    .A2(_0240_),
    .Y(_0288_),
    .B1(_0287_));
 sg13g2_nor3_1 _2410_ (.A(net91),
    .B(_0964_),
    .C(_0255_),
    .Y(_0289_));
 sg13g2_a21o_1 _2411_ (.A2(_0288_),
    .A1(net91),
    .B1(_0289_),
    .X(_0290_));
 sg13g2_nand3_1 _2412_ (.B(_0286_),
    .C(_0290_),
    .A(_0283_),
    .Y(_0291_));
 sg13g2_a21o_1 _2413_ (.A2(_0286_),
    .A1(_0283_),
    .B1(_0290_),
    .X(_0292_));
 sg13g2_a21oi_1 _2414_ (.A1(_0291_),
    .A2(_0292_),
    .Y(_0293_),
    .B1(_1162_));
 sg13g2_nor3_1 _2415_ (.A(_0229_),
    .B(net78),
    .C(_0831_),
    .Y(_0294_));
 sg13g2_nor2_1 _2416_ (.A(net91),
    .B(_0294_),
    .Y(_0295_));
 sg13g2_and2_1 _2417_ (.A(_1362_),
    .B(_1427_),
    .X(_0296_));
 sg13g2_nand2_1 _2418_ (.Y(_0297_),
    .A(_1012_),
    .B(_0296_));
 sg13g2_mux2_1 _2419_ (.A0(net91),
    .A1(_0295_),
    .S(_0297_),
    .X(_0298_));
 sg13g2_and2_1 _2420_ (.A(_0824_),
    .B(_0298_),
    .X(_0299_));
 sg13g2_nor3_1 _2421_ (.A(net79),
    .B(net78),
    .C(_0298_),
    .Y(_0300_));
 sg13g2_o21ai_1 _2422_ (.B1(_1012_),
    .Y(_0301_),
    .A1(_1348_),
    .A2(_1362_));
 sg13g2_or2_1 _2423_ (.X(_0302_),
    .B(_1394_),
    .A(net92));
 sg13g2_a22oi_1 _2424_ (.Y(_0303_),
    .B1(_0302_),
    .B2(_1348_),
    .A2(_0301_),
    .A1(_1393_));
 sg13g2_buf_1 _2425_ (.A(_0303_),
    .X(_0304_));
 sg13g2_mux2_1 _2426_ (.A0(_0299_),
    .A1(_0300_),
    .S(_0304_),
    .X(_0305_));
 sg13g2_nor2_1 _2427_ (.A(net81),
    .B(net65),
    .Y(_0306_));
 sg13g2_a221oi_1 _2428_ (.B2(net80),
    .C1(net41),
    .B1(_0306_),
    .A1(net65),
    .Y(_0307_),
    .A2(_0814_));
 sg13g2_nor4_1 _2429_ (.A(_0277_),
    .B(_0293_),
    .C(_0305_),
    .D(_0307_),
    .Y(_0308_));
 sg13g2_o21ai_1 _2430_ (.B1(_0308_),
    .Y(_0309_),
    .A1(_0266_),
    .A2(_0268_));
 sg13g2_or2_1 _2431_ (.X(_0310_),
    .B(_0260_),
    .A(_0265_));
 sg13g2_inv_1 _2432_ (.Y(_0311_),
    .A(_0218_));
 sg13g2_nor3_1 _2433_ (.A(_0311_),
    .B(_0250_),
    .C(_0259_),
    .Y(_0312_));
 sg13g2_and2_1 _2434_ (.A(_0308_),
    .B(_0312_),
    .X(_0313_));
 sg13g2_or4_1 _2435_ (.A(_0277_),
    .B(_0293_),
    .C(_0305_),
    .D(_0307_),
    .X(_0314_));
 sg13g2_o21ai_1 _2436_ (.B1(_0218_),
    .Y(_0315_),
    .A1(_0250_),
    .A2(_0259_));
 sg13g2_nor4_1 _2437_ (.A(_0314_),
    .B(_0265_),
    .C(_0260_),
    .D(_0315_),
    .Y(_0316_));
 sg13g2_a221oi_1 _2438_ (.B2(_0313_),
    .C1(_0316_),
    .B1(_0310_),
    .A1(_0218_),
    .Y(_0317_),
    .A2(net25));
 sg13g2_and3_1 _2439_ (.X(_0318_),
    .A(_0954_),
    .B(_0309_),
    .C(_0317_));
 sg13g2_o21ai_1 _2440_ (.B1(_0318_),
    .Y(_0319_),
    .A1(net22),
    .A2(_0217_));
 sg13g2_and2_1 _2441_ (.A(_0309_),
    .B(_0317_),
    .X(_0320_));
 sg13g2_buf_1 _2442_ (.A(_0320_),
    .X(_0321_));
 sg13g2_or4_1 _2443_ (.A(_0933_),
    .B(net22),
    .C(_0217_),
    .D(_0321_),
    .X(_0322_));
 sg13g2_mux4_1 _2444_ (.S0(_0928_),
    .A0(net97),
    .A1(net72),
    .A2(net90),
    .A3(_0271_),
    .S1(net94),
    .X(_0323_));
 sg13g2_nand2b_1 _2445_ (.Y(_0324_),
    .B(_1146_),
    .A_N(_1230_));
 sg13g2_and3_1 _2446_ (.X(_0325_),
    .A(net73),
    .B(_1231_),
    .C(_0324_));
 sg13g2_nor2_1 _2447_ (.A(_1283_),
    .B(_1284_),
    .Y(_0326_));
 sg13g2_nand2_1 _2448_ (.Y(_0327_),
    .A(_0817_),
    .B(net72));
 sg13g2_o21ai_1 _2449_ (.B1(_0327_),
    .Y(_0328_),
    .A1(net52),
    .A2(net72));
 sg13g2_nand2_1 _2450_ (.Y(_0329_),
    .A(_0988_),
    .B(_0328_));
 sg13g2_o21ai_1 _2451_ (.B1(net57),
    .Y(_0330_),
    .A1(_0988_),
    .A2(_0808_));
 sg13g2_o21ai_1 _2452_ (.B1(_1456_),
    .Y(_0331_),
    .A1(_1295_),
    .A2(_1244_));
 sg13g2_o21ai_1 _2453_ (.B1(net50),
    .Y(_0332_),
    .A1(net48),
    .A2(_1235_));
 sg13g2_nand2_1 _2454_ (.Y(_0333_),
    .A(net48),
    .B(net97));
 sg13g2_a21oi_1 _2455_ (.A1(_0332_),
    .A2(_0333_),
    .Y(_0334_),
    .B1(_1293_));
 sg13g2_a221oi_1 _2456_ (.B2(_1293_),
    .C1(_0334_),
    .B1(_0331_),
    .A1(_1306_),
    .Y(_0335_),
    .A2(_0330_));
 sg13g2_inv_1 _2457_ (.Y(_0336_),
    .A(_0006_));
 sg13g2_nand2b_1 _2458_ (.Y(_0337_),
    .B(net74),
    .A_N(_0021_));
 sg13g2_o21ai_1 _2459_ (.B1(_0337_),
    .Y(_0338_),
    .A1(net74),
    .A2(_1244_));
 sg13g2_a22oi_1 _2460_ (.Y(_0339_),
    .B1(_0338_),
    .B2(_1306_),
    .A2(_0846_),
    .A1(_0336_));
 sg13g2_nand2_1 _2461_ (.Y(_0340_),
    .A(_1260_),
    .B(_0787_));
 sg13g2_o21ai_1 _2462_ (.B1(_0340_),
    .Y(_0341_),
    .A1(_1260_),
    .A2(_0339_));
 sg13g2_a22oi_1 _2463_ (.Y(_0342_),
    .B1(_0341_),
    .B2(net36),
    .A2(_0335_),
    .A1(_0329_));
 sg13g2_a21oi_1 _2464_ (.A1(net97),
    .A2(net25),
    .Y(_0343_),
    .B1(_0926_));
 sg13g2_nand2b_1 _2465_ (.Y(_0344_),
    .B(_0343_),
    .A_N(_0342_));
 sg13g2_o21ai_1 _2466_ (.B1(_1303_),
    .Y(_0345_),
    .A1(net50),
    .A2(_0252_));
 sg13g2_nand2_1 _2467_ (.Y(_0346_),
    .A(net66),
    .B(_0252_));
 sg13g2_nor2_1 _2468_ (.A(net53),
    .B(net57),
    .Y(_0347_));
 sg13g2_a22oi_1 _2469_ (.Y(_0348_),
    .B1(_0346_),
    .B2(_0347_),
    .A2(_0345_),
    .A1(_0244_));
 sg13g2_nand2_1 _2470_ (.Y(_0349_),
    .A(net90),
    .B(net65));
 sg13g2_inv_1 _2471_ (.Y(_0350_),
    .A(_0005_));
 sg13g2_a221oi_1 _2472_ (.B2(_0311_),
    .C1(net52),
    .B1(_1007_),
    .A1(_0350_),
    .Y(_0351_),
    .A2(_0846_));
 sg13g2_a21oi_1 _2473_ (.A1(net52),
    .A2(_0349_),
    .Y(_0352_),
    .B1(_0351_));
 sg13g2_nand4_1 _2474_ (.B(_0230_),
    .C(_0271_),
    .A(net80),
    .Y(_0353_),
    .D(_0838_));
 sg13g2_o21ai_1 _2475_ (.B1(_0353_),
    .Y(_0354_),
    .A1(net47),
    .A2(_0911_));
 sg13g2_nor2_1 _2476_ (.A(net51),
    .B(_0244_),
    .Y(_0355_));
 sg13g2_a21oi_1 _2477_ (.A1(net58),
    .A2(net90),
    .Y(_0356_),
    .B1(net52));
 sg13g2_nor3_1 _2478_ (.A(net65),
    .B(_0355_),
    .C(_0356_),
    .Y(_0357_));
 sg13g2_a221oi_1 _2479_ (.B2(net53),
    .C1(_0357_),
    .B1(_0354_),
    .A1(net36),
    .Y(_0358_),
    .A2(_0352_));
 sg13g2_o21ai_1 _2480_ (.B1(_0358_),
    .Y(_0359_),
    .A1(net49),
    .A2(_0348_));
 sg13g2_a21oi_1 _2481_ (.A1(_0230_),
    .A2(net25),
    .Y(_0360_),
    .B1(_0926_));
 sg13g2_nand2_1 _2482_ (.Y(_0361_),
    .A(_0359_),
    .B(_0360_));
 sg13g2_mux2_1 _2483_ (.A0(_0344_),
    .A1(_0361_),
    .S(_0927_),
    .X(_0362_));
 sg13g2_nor2_1 _2484_ (.A(_1284_),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_a221oi_1 _2485_ (.B2(_0326_),
    .C1(_0363_),
    .B1(_0325_),
    .A1(_0929_),
    .Y(_0364_),
    .A2(_0323_));
 sg13g2_and3_1 _2486_ (.X(_0365_),
    .A(_0319_),
    .B(_0322_),
    .C(_0364_));
 sg13g2_buf_8 _2487_ (.A(_0365_),
    .X(_0366_));
 sg13g2_buf_8 _2488_ (.A(_0366_),
    .X(_0367_));
 sg13g2_mux2_1 _2489_ (.A0(_0213_),
    .A1(_0216_),
    .S(net16),
    .X(_0368_));
 sg13g2_nor2_1 _2490_ (.A(net21),
    .B(net16),
    .Y(_0369_));
 sg13g2_and2_1 _2491_ (.A(net20),
    .B(net18),
    .X(_0370_));
 sg13g2_buf_1 _2492_ (.A(_0370_),
    .X(_0371_));
 sg13g2_a221oi_1 _2493_ (.B2(_0371_),
    .C1(_0763_),
    .B1(_0369_),
    .A1(net21),
    .Y(_0372_),
    .A2(_0368_));
 sg13g2_a21o_1 _2494_ (.A2(net8),
    .A1(net112),
    .B1(_0372_),
    .X(_0032_));
 sg13g2_nand2b_1 _2495_ (.Y(_0373_),
    .B(net18),
    .A_N(net20));
 sg13g2_nand2b_1 _2496_ (.Y(_0374_),
    .B(net19),
    .A_N(net20));
 sg13g2_nand2_1 _2497_ (.Y(_0375_),
    .A(net21),
    .B(net16));
 sg13g2_mux2_1 _2498_ (.A0(_0373_),
    .A1(_0374_),
    .S(_0375_),
    .X(_0376_));
 sg13g2_nand2_1 _2499_ (.Y(_0377_),
    .A(_0215_),
    .B(_0369_));
 sg13g2_nand2_1 _2500_ (.Y(_0378_),
    .A(_0376_),
    .B(_0377_));
 sg13g2_nand2_1 _2501_ (.Y(_0379_),
    .A(net112),
    .B(net9));
 sg13g2_o21ai_1 _2502_ (.B1(_0379_),
    .Y(_0033_),
    .A1(net112),
    .A2(_0378_));
 sg13g2_nand2_1 _2503_ (.Y(_0380_),
    .A(_1280_),
    .B(_1335_));
 sg13g2_buf_1 _2504_ (.A(_0380_),
    .X(_0381_));
 sg13g2_buf_8 _2505_ (.A(net20),
    .X(_0382_));
 sg13g2_nand3_1 _2506_ (.B(net20),
    .C(net19),
    .A(net16),
    .Y(_0383_));
 sg13g2_o21ai_1 _2507_ (.B1(_0383_),
    .Y(_0384_),
    .A1(net16),
    .A2(net15));
 sg13g2_nor3_1 _2508_ (.A(net16),
    .B(net20),
    .C(net18),
    .Y(_0385_));
 sg13g2_a21o_1 _2509_ (.A2(_0384_),
    .A1(net17),
    .B1(_0385_),
    .X(_0386_));
 sg13g2_nand2_1 _2510_ (.Y(_0387_),
    .A(net112),
    .B(net10));
 sg13g2_o21ai_1 _2511_ (.B1(_0387_),
    .Y(_0034_),
    .A1(_0763_),
    .A2(_0386_));
 sg13g2_nand3_1 _2512_ (.B(_0322_),
    .C(_0364_),
    .A(_0319_),
    .Y(_0388_));
 sg13g2_buf_2 _2513_ (.A(_0388_),
    .X(_0389_));
 sg13g2_nor3_1 _2514_ (.A(net17),
    .B(_0389_),
    .C(net18),
    .Y(_0390_));
 sg13g2_nor2_1 _2515_ (.A(_1337_),
    .B(net19),
    .Y(_0391_));
 sg13g2_nor3_1 _2516_ (.A(net15),
    .B(_0390_),
    .C(_0391_),
    .Y(_0392_));
 sg13g2_nor3_1 _2517_ (.A(_1336_),
    .B(_0366_),
    .C(net18),
    .Y(_0393_));
 sg13g2_o21ai_1 _2518_ (.B1(net15),
    .Y(_0394_),
    .A1(net17),
    .A2(net19));
 sg13g2_nor2_1 _2519_ (.A(_0393_),
    .B(_0394_),
    .Y(_0395_));
 sg13g2_or2_1 _2520_ (.X(_0396_),
    .B(_0395_),
    .A(_0392_));
 sg13g2_buf_1 _2521_ (.A(net132),
    .X(_0397_));
 sg13g2_mux2_1 _2522_ (.A0(net11),
    .A1(_0396_),
    .S(net89),
    .X(_0035_));
 sg13g2_nand2b_1 _2523_ (.Y(_0398_),
    .B(_1337_),
    .A_N(net20));
 sg13g2_a21oi_1 _2524_ (.A1(net19),
    .A2(_0398_),
    .Y(_0399_),
    .B1(_0389_));
 sg13g2_a21oi_1 _2525_ (.A1(net21),
    .A2(_0371_),
    .Y(_0400_),
    .B1(_0399_));
 sg13g2_mux2_1 _2526_ (.A0(net12),
    .A1(_0400_),
    .S(net89),
    .X(_0036_));
 sg13g2_nor2_1 _2527_ (.A(net21),
    .B(_0389_),
    .Y(_0401_));
 sg13g2_a22oi_1 _2528_ (.Y(_0402_),
    .B1(_0401_),
    .B2(_0374_),
    .A2(_0371_),
    .A1(net16));
 sg13g2_nor2_1 _2529_ (.A(net17),
    .B(_0366_),
    .Y(_0403_));
 sg13g2_nand2_1 _2530_ (.Y(_0404_),
    .A(_0213_),
    .B(_0403_));
 sg13g2_and2_1 _2531_ (.A(_0402_),
    .B(_0404_),
    .X(_0405_));
 sg13g2_mux2_1 _2532_ (.A0(net13),
    .A1(_0405_),
    .S(_0397_),
    .X(_0037_));
 sg13g2_nor2_1 _2533_ (.A(_0367_),
    .B(net18),
    .Y(_0406_));
 sg13g2_nor2_1 _2534_ (.A(net17),
    .B(_0382_),
    .Y(_0407_));
 sg13g2_mux2_1 _2535_ (.A0(_0382_),
    .A1(_0213_),
    .S(net17),
    .X(_0408_));
 sg13g2_a221oi_1 _2536_ (.B2(_0367_),
    .C1(_0762_),
    .B1(_0408_),
    .A1(_0406_),
    .Y(_0409_),
    .A2(_0407_));
 sg13g2_a21o_1 _2537_ (.A2(net14),
    .A1(net112),
    .B1(_0409_),
    .X(_0038_));
 sg13g2_buf_1 _2538_ (.A(\spi_wrapper_i.reg_data_o[0] ),
    .X(_0410_));
 sg13g2_buf_2 _2539_ (.A(\spi_wrapper_i.reg_addr[1] ),
    .X(_0411_));
 sg13g2_buf_1 _2540_ (.A(_0411_),
    .X(_0412_));
 sg13g2_buf_1 _2541_ (.A(net88),
    .X(_0413_));
 sg13g2_buf_1 _2542_ (.A(\spi_wrapper_i.reg_addr[0] ),
    .X(_0414_));
 sg13g2_buf_1 _2543_ (.A(net121),
    .X(_0415_));
 sg13g2_buf_1 _2544_ (.A(net87),
    .X(_0416_));
 sg13g2_nand2_1 _2545_ (.Y(_0417_),
    .A(_0749_),
    .B(\spi_wrapper_i.reg_data_o_vld ));
 sg13g2_buf_2 _2546_ (.A(_0417_),
    .X(_0418_));
 sg13g2_or4_1 _2547_ (.A(net64),
    .B(net63),
    .C(\spi_wrapper_i.reg_addr[2] ),
    .D(_0418_),
    .X(_0419_));
 sg13g2_buf_4 _2548_ (.X(_0420_),
    .A(_0419_));
 sg13g2_mux2_1 _2549_ (.A0(_0410_),
    .A1(net98),
    .S(_0420_),
    .X(_0039_));
 sg13g2_buf_1 _2550_ (.A(\spi_wrapper_i.reg_data_o[1] ),
    .X(_0421_));
 sg13g2_mux2_1 _2551_ (.A0(net120),
    .A1(net70),
    .S(_0420_),
    .X(_0040_));
 sg13g2_buf_1 _2552_ (.A(\spi_wrapper_i.reg_data_o[2] ),
    .X(_0422_));
 sg13g2_mux2_1 _2553_ (.A0(net119),
    .A1(net95),
    .S(_0420_),
    .X(_0041_));
 sg13g2_buf_1 _2554_ (.A(\spi_wrapper_i.reg_data_o[3] ),
    .X(_0423_));
 sg13g2_mux2_1 _2555_ (.A0(net118),
    .A1(_1031_),
    .S(_0420_),
    .X(_0042_));
 sg13g2_buf_1 _2556_ (.A(\spi_wrapper_i.reg_data_o[4] ),
    .X(_0424_));
 sg13g2_mux2_1 _2557_ (.A0(net117),
    .A1(net76),
    .S(_0420_),
    .X(_0043_));
 sg13g2_buf_1 _2558_ (.A(\spi_wrapper_i.reg_data_o[5] ),
    .X(_0425_));
 sg13g2_mux2_1 _2559_ (.A0(net116),
    .A1(net111),
    .S(_0420_),
    .X(_0044_));
 sg13g2_buf_1 _2560_ (.A(\spi_wrapper_i.reg_data_o[6] ),
    .X(_0426_));
 sg13g2_mux2_1 _2561_ (.A0(net115),
    .A1(net67),
    .S(_0420_),
    .X(_0045_));
 sg13g2_buf_1 _2562_ (.A(\spi_wrapper_i.reg_data_o[7] ),
    .X(_0427_));
 sg13g2_mux2_1 _2563_ (.A0(net114),
    .A1(net90),
    .S(_0420_),
    .X(_0046_));
 sg13g2_buf_2 _2564_ (.A(_0015_),
    .X(_0428_));
 sg13g2_nand2_2 _2565_ (.Y(_0429_),
    .A(net121),
    .B(_0428_));
 sg13g2_nor3_2 _2566_ (.A(net64),
    .B(_0418_),
    .C(_0429_),
    .Y(_0430_));
 sg13g2_buf_1 _2567_ (.A(_0430_),
    .X(_0431_));
 sg13g2_mux2_1 _2568_ (.A0(net99),
    .A1(net122),
    .S(net34),
    .X(_0047_));
 sg13g2_nand2_1 _2569_ (.Y(_0432_),
    .A(_0421_),
    .B(net34));
 sg13g2_o21ai_1 _2570_ (.B1(_0432_),
    .Y(_0048_),
    .A1(_0998_),
    .A2(net34));
 sg13g2_nand2_1 _2571_ (.Y(_0433_),
    .A(_0422_),
    .B(net34));
 sg13g2_o21ai_1 _2572_ (.B1(_0433_),
    .Y(_0049_),
    .A1(_1149_),
    .A2(_0431_));
 sg13g2_mux2_1 _2573_ (.A0(_0958_),
    .A1(_0423_),
    .S(_0431_),
    .X(_0050_));
 sg13g2_nand2_1 _2574_ (.Y(_0434_),
    .A(net117),
    .B(_0430_));
 sg13g2_o21ai_1 _2575_ (.B1(_0434_),
    .Y(_0051_),
    .A1(_0855_),
    .A2(net34));
 sg13g2_mux2_1 _2576_ (.A0(net84),
    .A1(net116),
    .S(net34),
    .X(_0052_));
 sg13g2_nand2_1 _2577_ (.Y(_0435_),
    .A(net115),
    .B(_0430_));
 sg13g2_o21ai_1 _2578_ (.B1(_0435_),
    .Y(_0053_),
    .A1(_1348_),
    .A2(net34));
 sg13g2_nand2_1 _2579_ (.Y(_0436_),
    .A(net114),
    .B(_0430_));
 sg13g2_o21ai_1 _2580_ (.B1(_0436_),
    .Y(_0054_),
    .A1(_0252_),
    .A2(net34));
 sg13g2_inv_2 _2581_ (.Y(_0437_),
    .A(_0411_));
 sg13g2_buf_1 _2582_ (.A(_0437_),
    .X(_0438_));
 sg13g2_inv_2 _2583_ (.Y(_0439_),
    .A(_0428_));
 sg13g2_buf_1 _2584_ (.A(_0439_),
    .X(_0440_));
 sg13g2_nor4_2 _2585_ (.A(net62),
    .B(net63),
    .C(net61),
    .Y(_0441_),
    .D(_0418_));
 sg13g2_buf_1 _2586_ (.A(_0441_),
    .X(_0442_));
 sg13g2_nand2_1 _2587_ (.Y(_0443_),
    .A(net122),
    .B(net33));
 sg13g2_o21ai_1 _2588_ (.B1(_0443_),
    .Y(_0055_),
    .A1(_1320_),
    .A2(net33));
 sg13g2_nand2_1 _2589_ (.Y(_0444_),
    .A(net120),
    .B(net33));
 sg13g2_o21ai_1 _2590_ (.B1(_0444_),
    .Y(_0056_),
    .A1(net52),
    .A2(net33));
 sg13g2_nand2_1 _2591_ (.Y(_0445_),
    .A(net119),
    .B(_0441_));
 sg13g2_o21ai_1 _2592_ (.B1(_0445_),
    .Y(_0057_),
    .A1(net53),
    .A2(_0442_));
 sg13g2_nand2_1 _2593_ (.Y(_0446_),
    .A(net118),
    .B(_0441_));
 sg13g2_o21ai_1 _2594_ (.B1(_0446_),
    .Y(_0058_),
    .A1(net58),
    .A2(_0442_));
 sg13g2_nand2_1 _2595_ (.Y(_0447_),
    .A(net117),
    .B(_0441_));
 sg13g2_o21ai_1 _2596_ (.B1(_0447_),
    .Y(_0059_),
    .A1(net73),
    .A2(net33));
 sg13g2_mux2_1 _2597_ (.A0(\alu_74181_i0.alu_74181_arith_inst.cn ),
    .A1(net116),
    .S(net33),
    .X(_0060_));
 sg13g2_mux2_1 _2598_ (.A0(\config_regs[22] ),
    .A1(net115),
    .S(net33),
    .X(_0061_));
 sg13g2_mux2_1 _2599_ (.A0(\config_regs[23] ),
    .A1(net114),
    .S(net33),
    .X(_0062_));
 sg13g2_buf_1 _2600_ (.A(_0428_),
    .X(_0448_));
 sg13g2_buf_1 _2601_ (.A(net86),
    .X(_0449_));
 sg13g2_inv_1 _2602_ (.Y(_0450_),
    .A(_0414_));
 sg13g2_nor2_1 _2603_ (.A(_0437_),
    .B(_0450_),
    .Y(_0451_));
 sg13g2_buf_1 _2604_ (.A(_0451_),
    .X(_0452_));
 sg13g2_nand2_1 _2605_ (.Y(_0453_),
    .A(net60),
    .B(net46));
 sg13g2_buf_1 _2606_ (.A(_0453_),
    .X(_0454_));
 sg13g2_nor2_1 _2607_ (.A(_0418_),
    .B(_0454_),
    .Y(_0455_));
 sg13g2_buf_1 _2608_ (.A(_0455_),
    .X(_0456_));
 sg13g2_mux2_1 _2609_ (.A0(net94),
    .A1(net122),
    .S(net23),
    .X(_0063_));
 sg13g2_mux2_1 _2610_ (.A0(_0928_),
    .A1(net120),
    .S(net23),
    .X(_0064_));
 sg13g2_nand2_1 _2611_ (.Y(_0457_),
    .A(net119),
    .B(net23));
 sg13g2_o21ai_1 _2612_ (.B1(_0457_),
    .Y(_0065_),
    .A1(_0929_),
    .A2(_0456_));
 sg13g2_mux2_1 _2613_ (.A0(\config_regs[27] ),
    .A1(net118),
    .S(_0456_),
    .X(_0066_));
 sg13g2_mux2_1 _2614_ (.A0(\config_regs[28] ),
    .A1(net117),
    .S(net23),
    .X(_0067_));
 sg13g2_inv_1 _2615_ (.Y(_0458_),
    .A(\config_regs[29] ));
 sg13g2_nand2_1 _2616_ (.Y(_0459_),
    .A(net116),
    .B(net23));
 sg13g2_o21ai_1 _2617_ (.B1(_0459_),
    .Y(_0068_),
    .A1(_0458_),
    .A2(net23));
 sg13g2_mux2_1 _2618_ (.A0(\config_regs[30] ),
    .A1(net115),
    .S(net23),
    .X(_0069_));
 sg13g2_mux2_1 _2619_ (.A0(\config_regs[31] ),
    .A1(net114),
    .S(net23),
    .X(_0070_));
 sg13g2_inv_1 _2620_ (.Y(_0460_),
    .A(\config_regs[32] ));
 sg13g2_buf_1 _2621_ (.A(net60),
    .X(_0461_));
 sg13g2_nor4_1 _2622_ (.A(net64),
    .B(net63),
    .C(net45),
    .D(_0418_),
    .Y(_0462_));
 sg13g2_buf_1 _2623_ (.A(_0462_),
    .X(_0463_));
 sg13g2_nand2_1 _2624_ (.Y(_0464_),
    .A(net122),
    .B(net26));
 sg13g2_o21ai_1 _2625_ (.B1(_0464_),
    .Y(_0071_),
    .A1(_0460_),
    .A2(net26));
 sg13g2_mux2_1 _2626_ (.A0(\config_regs[33] ),
    .A1(net120),
    .S(net26),
    .X(_0072_));
 sg13g2_mux2_1 _2627_ (.A0(\config_regs[34] ),
    .A1(net119),
    .S(net26),
    .X(_0073_));
 sg13g2_mux2_1 _2628_ (.A0(\config_regs[35] ),
    .A1(net118),
    .S(net26),
    .X(_0074_));
 sg13g2_mux2_1 _2629_ (.A0(\config_regs[36] ),
    .A1(net117),
    .S(_0463_),
    .X(_0075_));
 sg13g2_mux2_1 _2630_ (.A0(\config_regs[37] ),
    .A1(net116),
    .S(net26),
    .X(_0076_));
 sg13g2_mux2_1 _2631_ (.A0(\config_regs[38] ),
    .A1(net115),
    .S(net26),
    .X(_0077_));
 sg13g2_mux2_1 _2632_ (.A0(\config_regs[39] ),
    .A1(net114),
    .S(net26),
    .X(_0078_));
 sg13g2_buf_1 _2633_ (.A(_0450_),
    .X(_0465_));
 sg13g2_nor4_1 _2634_ (.A(net64),
    .B(net59),
    .C(net45),
    .D(_0418_),
    .Y(_0466_));
 sg13g2_buf_4 _2635_ (.X(_0467_),
    .A(_0466_));
 sg13g2_mux2_1 _2636_ (.A0(\config_regs[40] ),
    .A1(net122),
    .S(_0467_),
    .X(_0079_));
 sg13g2_mux2_1 _2637_ (.A0(\config_regs[41] ),
    .A1(net120),
    .S(_0467_),
    .X(_0080_));
 sg13g2_mux2_1 _2638_ (.A0(\config_regs[42] ),
    .A1(net119),
    .S(_0467_),
    .X(_0081_));
 sg13g2_mux2_1 _2639_ (.A0(\config_regs[43] ),
    .A1(net118),
    .S(_0467_),
    .X(_0082_));
 sg13g2_mux2_1 _2640_ (.A0(\config_regs[44] ),
    .A1(net117),
    .S(_0467_),
    .X(_0083_));
 sg13g2_mux2_1 _2641_ (.A0(\config_regs[45] ),
    .A1(net116),
    .S(_0467_),
    .X(_0084_));
 sg13g2_mux2_1 _2642_ (.A0(\config_regs[46] ),
    .A1(net115),
    .S(_0467_),
    .X(_0085_));
 sg13g2_mux2_1 _2643_ (.A0(\config_regs[47] ),
    .A1(net114),
    .S(_0467_),
    .X(_0086_));
 sg13g2_nor4_1 _2644_ (.A(net62),
    .B(net63),
    .C(net45),
    .D(_0418_),
    .Y(_0468_));
 sg13g2_buf_4 _2645_ (.X(_0469_),
    .A(_0468_));
 sg13g2_mux2_1 _2646_ (.A0(\config_regs[48] ),
    .A1(net122),
    .S(_0469_),
    .X(_0087_));
 sg13g2_mux2_1 _2647_ (.A0(\config_regs[49] ),
    .A1(net120),
    .S(_0469_),
    .X(_0088_));
 sg13g2_mux2_1 _2648_ (.A0(\config_regs[50] ),
    .A1(net119),
    .S(_0469_),
    .X(_0089_));
 sg13g2_mux2_1 _2649_ (.A0(\config_regs[51] ),
    .A1(net118),
    .S(_0469_),
    .X(_0090_));
 sg13g2_mux2_1 _2650_ (.A0(\config_regs[52] ),
    .A1(net117),
    .S(_0469_),
    .X(_0091_));
 sg13g2_mux2_1 _2651_ (.A0(\config_regs[53] ),
    .A1(net116),
    .S(_0469_),
    .X(_0092_));
 sg13g2_mux2_1 _2652_ (.A0(\config_regs[54] ),
    .A1(net115),
    .S(_0469_),
    .X(_0093_));
 sg13g2_mux2_1 _2653_ (.A0(\config_regs[55] ),
    .A1(net114),
    .S(_0469_),
    .X(_0094_));
 sg13g2_nand2_1 _2654_ (.Y(_0470_),
    .A(net64),
    .B(net87));
 sg13g2_nor3_1 _2655_ (.A(net45),
    .B(_0418_),
    .C(_0470_),
    .Y(_0471_));
 sg13g2_buf_4 _2656_ (.X(_0472_),
    .A(_0471_));
 sg13g2_mux2_1 _2657_ (.A0(\config_regs[56] ),
    .A1(net122),
    .S(_0472_),
    .X(_0095_));
 sg13g2_mux2_1 _2658_ (.A0(\config_regs[57] ),
    .A1(net120),
    .S(_0472_),
    .X(_0096_));
 sg13g2_mux2_1 _2659_ (.A0(\config_regs[58] ),
    .A1(net119),
    .S(_0472_),
    .X(_0097_));
 sg13g2_mux2_1 _2660_ (.A0(\config_regs[59] ),
    .A1(net118),
    .S(_0472_),
    .X(_0098_));
 sg13g2_mux2_1 _2661_ (.A0(\config_regs[60] ),
    .A1(net117),
    .S(_0472_),
    .X(_0099_));
 sg13g2_mux2_1 _2662_ (.A0(\config_regs[61] ),
    .A1(net116),
    .S(_0472_),
    .X(_0100_));
 sg13g2_mux2_1 _2663_ (.A0(\config_regs[62] ),
    .A1(net115),
    .S(_0472_),
    .X(_0101_));
 sg13g2_mux2_1 _2664_ (.A0(\config_regs[63] ),
    .A1(net114),
    .S(_0472_),
    .X(_0102_));
 sg13g2_nand2_1 _2665_ (.Y(_0473_),
    .A(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .B(net42));
 sg13g2_o21ai_1 _2666_ (.B1(_0473_),
    .Y(_0103_),
    .A1(net59),
    .A2(net42));
 sg13g2_nand2_1 _2667_ (.Y(_0474_),
    .A(\spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .B(net42));
 sg13g2_o21ai_1 _2668_ (.B1(_0474_),
    .Y(_0104_),
    .A1(net62),
    .A2(net42));
 sg13g2_mux2_1 _2669_ (.A0(\spi_wrapper_i.reg_addr[2] ),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .S(net42),
    .X(_0105_));
 sg13g2_buf_1 _2670_ (.A(\spi_wrapper_i.reg_addr[3] ),
    .X(_0475_));
 sg13g2_inv_1 _2671_ (.Y(_0476_),
    .A(_0475_));
 sg13g2_nand2_1 _2672_ (.Y(_0477_),
    .A(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .B(net42));
 sg13g2_o21ai_1 _2673_ (.B1(_0477_),
    .Y(_0106_),
    .A1(_0476_),
    .A2(_0771_));
 sg13g2_nand2_1 _2674_ (.Y(_0478_),
    .A(net132),
    .B(\spi_wrapper_i.spi_reg_inst.state[4] ));
 sg13g2_nor2_1 _2675_ (.A(_0768_),
    .B(_0478_),
    .Y(_0479_));
 sg13g2_buf_1 _2676_ (.A(_0479_),
    .X(_0480_));
 sg13g2_mux2_1 _2677_ (.A0(net122),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .S(net32),
    .X(_0107_));
 sg13g2_mux2_1 _2678_ (.A0(net120),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .S(net32),
    .X(_0108_));
 sg13g2_mux2_1 _2679_ (.A0(net119),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .S(net32),
    .X(_0109_));
 sg13g2_mux2_1 _2680_ (.A0(net118),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .S(net32),
    .X(_0110_));
 sg13g2_mux2_1 _2681_ (.A0(_0424_),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[4] ),
    .S(net32),
    .X(_0111_));
 sg13g2_mux2_1 _2682_ (.A0(_0425_),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[5] ),
    .S(net32),
    .X(_0112_));
 sg13g2_mux2_1 _2683_ (.A0(_0426_),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[6] ),
    .S(net32),
    .X(_0113_));
 sg13g2_mux2_1 _2684_ (.A0(_0427_),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[7] ),
    .S(net32),
    .X(_0114_));
 sg13g2_a22oi_1 _2685_ (.Y(_0481_),
    .B1(_0480_),
    .B2(\spi_wrapper_i.spi_reg_inst.reg_rw ),
    .A2(\spi_wrapper_i.reg_data_o_vld ),
    .A1(net112));
 sg13g2_inv_1 _2686_ (.Y(_0115_),
    .A(_0481_));
 sg13g2_nand2_1 _2687_ (.Y(_0482_),
    .A(\spi_wrapper_i.spi_reg_inst.rx_buffer[7] ),
    .B(net42));
 sg13g2_o21ai_1 _2688_ (.B1(_0482_),
    .Y(_0116_),
    .A1(_0779_),
    .A2(net42));
 sg13g2_buf_1 _2689_ (.A(_0750_),
    .X(_0483_));
 sg13g2_nand2_1 _2690_ (.Y(_0484_),
    .A(net85),
    .B(_0753_));
 sg13g2_o21ai_1 _2691_ (.B1(_0484_),
    .Y(_0117_),
    .A1(net89),
    .A2(_0772_));
 sg13g2_mux2_1 _2692_ (.A0(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .A1(spi_clk_sync),
    .S(net89),
    .X(_0118_));
 sg13g2_nor2b_1 _2693_ (.A(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .B_N(spi_clk_sync),
    .Y(_0485_));
 sg13g2_nor2b_1 _2694_ (.A(spi_clk_sync),
    .B_N(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .Y(_0486_));
 sg13g2_xor2_1 _2695_ (.B(cpol_sync),
    .A(cpha_sync),
    .X(_0487_));
 sg13g2_mux2_1 _2696_ (.A0(_0485_),
    .A1(_0486_),
    .S(_0487_),
    .X(_0488_));
 sg13g2_and2_1 _2697_ (.A(_0014_),
    .B(_0488_),
    .X(_0489_));
 sg13g2_and2_1 _2698_ (.A(_0749_),
    .B(_0489_),
    .X(_0490_));
 sg13g2_buf_1 _2699_ (.A(_0490_),
    .X(_0491_));
 sg13g2_mux2_1 _2700_ (.A0(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .A1(spi_mosi_sync),
    .S(_0491_),
    .X(_0119_));
 sg13g2_nand2_1 _2701_ (.Y(_0492_),
    .A(net132),
    .B(_0489_));
 sg13g2_buf_1 _2702_ (.A(_0492_),
    .X(_0493_));
 sg13g2_mux2_1 _2703_ (.A0(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .S(net31),
    .X(_0120_));
 sg13g2_mux2_1 _2704_ (.A0(\spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .S(net31),
    .X(_0121_));
 sg13g2_mux2_1 _2705_ (.A0(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .S(net31),
    .X(_0122_));
 sg13g2_mux2_1 _2706_ (.A0(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[4] ),
    .S(net31),
    .X(_0123_));
 sg13g2_mux2_1 _2707_ (.A0(\spi_wrapper_i.spi_reg_inst.rx_buffer[4] ),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[5] ),
    .S(net31),
    .X(_0124_));
 sg13g2_mux2_1 _2708_ (.A0(\spi_wrapper_i.spi_reg_inst.rx_buffer[5] ),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[6] ),
    .S(net31),
    .X(_0125_));
 sg13g2_mux2_1 _2709_ (.A0(\spi_wrapper_i.spi_reg_inst.rx_buffer[6] ),
    .A1(\spi_wrapper_i.spi_reg_inst.rx_buffer[7] ),
    .S(net31),
    .X(_0126_));
 sg13g2_nor3_1 _2710_ (.A(_0765_),
    .B(_0776_),
    .C(net31),
    .Y(_0494_));
 sg13g2_a21o_1 _2711_ (.A2(_0493_),
    .A1(_0765_),
    .B1(_0494_),
    .X(_0127_));
 sg13g2_and2_1 _2712_ (.A(_0765_),
    .B(_0491_),
    .X(_0495_));
 sg13g2_buf_1 _2713_ (.A(_0495_),
    .X(_0496_));
 sg13g2_xor2_1 _2714_ (.B(_0496_),
    .A(_0764_),
    .X(_0128_));
 sg13g2_nand2_1 _2715_ (.Y(_0497_),
    .A(_0764_),
    .B(_0496_));
 sg13g2_xnor2_1 _2716_ (.Y(_0129_),
    .A(_0766_),
    .B(_0497_));
 sg13g2_a21oi_1 _2717_ (.A1(_0766_),
    .A2(_0496_),
    .Y(_0498_),
    .B1(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ));
 sg13g2_a21oi_1 _2718_ (.A1(net132),
    .A2(_0767_),
    .Y(_0499_),
    .B1(_0775_));
 sg13g2_nand4_1 _2719_ (.B(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ),
    .C(_0766_),
    .A(_0764_),
    .Y(_0500_),
    .D(_0496_));
 sg13g2_o21ai_1 _2720_ (.B1(_0500_),
    .Y(_0501_),
    .A1(_0764_),
    .A2(_0499_));
 sg13g2_nor2_1 _2721_ (.A(_0498_),
    .B(_0501_),
    .Y(_0130_));
 sg13g2_nand3b_1 _2722_ (.B(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .C(_0758_),
    .Y(_0502_),
    .A_N(_0755_));
 sg13g2_buf_1 _2723_ (.A(_0502_),
    .X(_0503_));
 sg13g2_inv_1 _2724_ (.Y(_0504_),
    .A(net44));
 sg13g2_nand2b_1 _2725_ (.Y(_0505_),
    .B(_0752_),
    .A_N(_0753_));
 sg13g2_nor2_2 _2726_ (.A(_0411_),
    .B(net121),
    .Y(_0506_));
 sg13g2_nand2_2 _2727_ (.Y(_0507_),
    .A(net60),
    .B(_0506_));
 sg13g2_mux4_1 _2728_ (.S0(net86),
    .A0(\config_regs[48] ),
    .A1(net49),
    .A2(\config_regs[56] ),
    .A3(net94),
    .S1(net87),
    .X(_0508_));
 sg13g2_nand2_1 _2729_ (.Y(_0509_),
    .A(_0428_),
    .B(_1043_));
 sg13g2_o21ai_1 _2730_ (.B1(_0509_),
    .Y(_0510_),
    .A1(net86),
    .A2(\config_regs[40] ));
 sg13g2_nor2_1 _2731_ (.A(net121),
    .B(_0428_),
    .Y(_0511_));
 sg13g2_a221oi_1 _2732_ (.B2(_0460_),
    .C1(net88),
    .B1(_0511_),
    .A1(net87),
    .Y(_0512_),
    .A2(_0510_));
 sg13g2_a21o_1 _2733_ (.A2(_0508_),
    .A1(net88),
    .B1(_0512_),
    .X(_0513_));
 sg13g2_o21ai_1 _2734_ (.B1(_0513_),
    .Y(_0514_),
    .A1(_1199_),
    .A2(_0507_));
 sg13g2_o21ai_1 _2735_ (.B1(net113),
    .Y(_0515_),
    .A1(_0184_),
    .A2(_0507_));
 sg13g2_o21ai_1 _2736_ (.B1(_0515_),
    .Y(_0516_),
    .A1(net113),
    .A2(_0514_));
 sg13g2_nand4_1 _2737_ (.B(_0504_),
    .C(_0505_),
    .A(net85),
    .Y(_0517_),
    .D(_0516_));
 sg13g2_xnor2_1 _2738_ (.Y(_0518_),
    .A(net17),
    .B(_0366_));
 sg13g2_nand4_1 _2739_ (.B(_0371_),
    .C(net46),
    .A(net45),
    .Y(_0519_),
    .D(_0518_));
 sg13g2_nor2_1 _2740_ (.A(net18),
    .B(_0454_),
    .Y(_0520_));
 sg13g2_o21ai_1 _2741_ (.B1(_0520_),
    .Y(_0521_),
    .A1(_0389_),
    .A2(_0398_));
 sg13g2_or3_1 _2742_ (.A(_0373_),
    .B(_0403_),
    .C(_0454_),
    .X(_0522_));
 sg13g2_a21o_1 _2743_ (.A2(net8),
    .A1(net61),
    .B1(_0465_),
    .X(_0523_));
 sg13g2_nor2_1 _2744_ (.A(_0437_),
    .B(_0439_),
    .Y(_0524_));
 sg13g2_nor2_1 _2745_ (.A(_0411_),
    .B(net86),
    .Y(_0525_));
 sg13g2_a21oi_1 _2746_ (.A1(net19),
    .A2(_0524_),
    .Y(_0526_),
    .B1(_0525_));
 sg13g2_a21oi_1 _2747_ (.A1(_0523_),
    .A2(_0526_),
    .Y(_0527_),
    .B1(_0476_));
 sg13g2_and4_1 _2748_ (.A(_0519_),
    .B(_0521_),
    .C(_0522_),
    .D(_0527_),
    .X(_0528_));
 sg13g2_mux2_1 _2749_ (.A0(_0486_),
    .A1(_0485_),
    .S(_0487_),
    .X(_0529_));
 sg13g2_nand2_1 _2750_ (.Y(_0530_),
    .A(_0014_),
    .B(_0529_));
 sg13g2_nand3_1 _2751_ (.B(net44),
    .C(_0505_),
    .A(_0530_),
    .Y(_0531_));
 sg13g2_nand2_1 _2752_ (.Y(_0532_),
    .A(_0749_),
    .B(_0531_));
 sg13g2_buf_1 _2753_ (.A(_0532_),
    .X(_0533_));
 sg13g2_nand2_1 _2754_ (.Y(_0534_),
    .A(\spi_wrapper_i.spi_reg_inst.tx_buffer[0] ),
    .B(net24));
 sg13g2_o21ai_1 _2755_ (.B1(_0534_),
    .Y(_0131_),
    .A1(_0517_),
    .A2(_0528_));
 sg13g2_buf_1 _2756_ (.A(net44),
    .X(_0535_));
 sg13g2_nor2_1 _2757_ (.A(_0753_),
    .B(_0772_),
    .Y(_0536_));
 sg13g2_nor2_2 _2758_ (.A(_0536_),
    .B(_0533_),
    .Y(_0537_));
 sg13g2_nand2_1 _2759_ (.Y(_0538_),
    .A(net113),
    .B(_0537_));
 sg13g2_a21oi_1 _2760_ (.A1(_0007_),
    .A2(net30),
    .Y(_0539_),
    .B1(_0538_));
 sg13g2_nand2b_1 _2761_ (.Y(_0540_),
    .B(_0539_),
    .A_N(_0454_));
 sg13g2_nor2_2 _2762_ (.A(_0450_),
    .B(net86),
    .Y(_0541_));
 sg13g2_nor2_1 _2763_ (.A(net121),
    .B(_0439_),
    .Y(_0542_));
 sg13g2_a22oi_1 _2764_ (.Y(_0543_),
    .B1(_0542_),
    .B2(net17),
    .A2(_0541_),
    .A1(net9));
 sg13g2_and2_1 _2765_ (.A(_0448_),
    .B(_0506_),
    .X(_0544_));
 sg13g2_buf_1 _2766_ (.A(_0544_),
    .X(_0545_));
 sg13g2_nand2b_1 _2767_ (.Y(_0546_),
    .B(net43),
    .A_N(_1317_));
 sg13g2_o21ai_1 _2768_ (.B1(_0546_),
    .Y(_0547_),
    .A1(net62),
    .A2(_0543_));
 sg13g2_inv_1 _2769_ (.Y(_0548_),
    .A(_0537_));
 sg13g2_inv_1 _2770_ (.Y(_0549_),
    .A(_0007_));
 sg13g2_nand2_1 _2771_ (.Y(_0550_),
    .A(_0411_),
    .B(\config_regs[49] ));
 sg13g2_nand2_1 _2772_ (.Y(_0551_),
    .A(_0437_),
    .B(\config_regs[33] ));
 sg13g2_a21oi_1 _2773_ (.A1(_0550_),
    .A2(_0551_),
    .Y(_0552_),
    .B1(net60));
 sg13g2_a21oi_1 _2774_ (.A1(_0449_),
    .A2(_1321_),
    .Y(_0553_),
    .B1(_0552_));
 sg13g2_nor2_1 _2775_ (.A(_0411_),
    .B(_0450_),
    .Y(_0554_));
 sg13g2_nand2_1 _2776_ (.Y(_0555_),
    .A(net121),
    .B(_0928_));
 sg13g2_a22oi_1 _2777_ (.Y(_0556_),
    .B1(_0555_),
    .B2(_0412_),
    .A2(_0554_),
    .A1(_0027_));
 sg13g2_mux2_1 _2778_ (.A0(\config_regs[41] ),
    .A1(\config_regs[57] ),
    .S(net88),
    .X(_0557_));
 sg13g2_a22oi_1 _2779_ (.Y(_0558_),
    .B1(_0541_),
    .B2(_0557_),
    .A2(_0556_),
    .A1(net45));
 sg13g2_o21ai_1 _2780_ (.B1(_0558_),
    .Y(_0559_),
    .A1(net63),
    .A2(_0553_));
 sg13g2_nand2_1 _2781_ (.Y(_0560_),
    .A(_0476_),
    .B(_0504_));
 sg13g2_a21oi_1 _2782_ (.A1(_0022_),
    .A2(net43),
    .Y(_0561_),
    .B1(_0560_));
 sg13g2_a22oi_1 _2783_ (.Y(_0562_),
    .B1(_0559_),
    .B2(_0561_),
    .A2(_0535_),
    .A1(_0549_));
 sg13g2_nor2_1 _2784_ (.A(_0548_),
    .B(_0562_),
    .Y(_0563_));
 sg13g2_a221oi_1 _2785_ (.B2(_0547_),
    .C1(_0563_),
    .B1(_0539_),
    .A1(\spi_wrapper_i.spi_reg_inst.tx_buffer[1] ),
    .Y(_0564_),
    .A2(net24));
 sg13g2_o21ai_1 _2786_ (.B1(_0564_),
    .Y(_0132_),
    .A1(_0378_),
    .A2(_0540_));
 sg13g2_xnor2_1 _2787_ (.Y(_0565_),
    .A(_1229_),
    .B(_1420_));
 sg13g2_and2_1 _2788_ (.A(_0925_),
    .B(_0156_),
    .X(_0566_));
 sg13g2_a21oi_1 _2789_ (.A1(_0953_),
    .A2(_0565_),
    .Y(_0567_),
    .B1(_0566_));
 sg13g2_a221oi_1 _2790_ (.B2(_0567_),
    .C1(_0538_),
    .B1(net43),
    .A1(_0008_),
    .Y(_0568_),
    .A2(net44));
 sg13g2_nand2b_1 _2791_ (.Y(_0569_),
    .B(_0568_),
    .A_N(_0454_));
 sg13g2_a21oi_1 _2792_ (.A1(net64),
    .A2(net15),
    .Y(_0570_),
    .B1(_0416_));
 sg13g2_nand4_1 _2793_ (.B(_0857_),
    .C(_0239_),
    .A(_0885_),
    .Y(_0571_),
    .D(_1434_));
 sg13g2_a21oi_1 _2794_ (.A1(_0346_),
    .A2(_0349_),
    .Y(_0572_),
    .B1(_0571_));
 sg13g2_nor4_1 _2795_ (.A(net88),
    .B(_0828_),
    .C(_0903_),
    .D(_0429_),
    .Y(_0573_));
 sg13g2_nor2_1 _2796_ (.A(_0437_),
    .B(_0428_),
    .Y(_0574_));
 sg13g2_a221oi_1 _2797_ (.B2(net10),
    .C1(_0511_),
    .B1(_0574_),
    .A1(_0572_),
    .Y(_0575_),
    .A2(_0573_));
 sg13g2_nand2b_1 _2798_ (.Y(_0576_),
    .B(_0575_),
    .A_N(_0570_));
 sg13g2_inv_1 _2799_ (.Y(_0577_),
    .A(_0008_));
 sg13g2_mux2_1 _2800_ (.A0(\config_regs[50] ),
    .A1(_1294_),
    .S(net60),
    .X(_0578_));
 sg13g2_a22oi_1 _2801_ (.Y(_0579_),
    .B1(_0578_),
    .B2(net59),
    .A2(_0541_),
    .A1(\config_regs[58] ));
 sg13g2_a22oi_1 _2802_ (.Y(_0580_),
    .B1(_0525_),
    .B2(\config_regs[42] ),
    .A2(_0524_),
    .A1(\config_regs[26] ));
 sg13g2_inv_1 _2803_ (.Y(_0581_),
    .A(_0580_));
 sg13g2_o21ai_1 _2804_ (.B1(net59),
    .Y(_0582_),
    .A1(_0448_),
    .A2(\config_regs[34] ));
 sg13g2_o21ai_1 _2805_ (.B1(_0582_),
    .Y(_0583_),
    .A1(_0439_),
    .A2(_0030_));
 sg13g2_a22oi_1 _2806_ (.Y(_0584_),
    .B1(_0583_),
    .B2(_0438_),
    .A2(_0581_),
    .A1(net87));
 sg13g2_o21ai_1 _2807_ (.B1(_0584_),
    .Y(_0585_),
    .A1(net62),
    .A2(_0579_));
 sg13g2_a21oi_1 _2808_ (.A1(_1117_),
    .A2(net43),
    .Y(_0586_),
    .B1(_0560_));
 sg13g2_a22oi_1 _2809_ (.Y(_0587_),
    .B1(_0585_),
    .B2(_0586_),
    .A2(net30),
    .A1(_0577_));
 sg13g2_nor2_1 _2810_ (.A(_0548_),
    .B(_0587_),
    .Y(_0588_));
 sg13g2_a221oi_1 _2811_ (.B2(_0576_),
    .C1(_0588_),
    .B1(_0568_),
    .A1(\spi_wrapper_i.spi_reg_inst.tx_buffer[2] ),
    .Y(_0589_),
    .A2(net24));
 sg13g2_o21ai_1 _2812_ (.B1(_0589_),
    .Y(_0133_),
    .A1(_0386_),
    .A2(_0569_));
 sg13g2_nand2_1 _2813_ (.Y(_0590_),
    .A(_0344_),
    .B(_0545_));
 sg13g2_and2_1 _2814_ (.A(_0009_),
    .B(net44),
    .X(_0591_));
 sg13g2_a21oi_1 _2815_ (.A1(net11),
    .A2(net46),
    .Y(_0592_),
    .B1(_0461_));
 sg13g2_nor3_1 _2816_ (.A(_0538_),
    .B(_0591_),
    .C(_0592_),
    .Y(_0593_));
 sg13g2_o21ai_1 _2817_ (.B1(_0593_),
    .Y(_0594_),
    .A1(_0325_),
    .A2(_0590_));
 sg13g2_nor4_1 _2818_ (.A(net15),
    .B(_0390_),
    .C(_0391_),
    .D(_0470_),
    .Y(_0595_));
 sg13g2_nor2_1 _2819_ (.A(_0381_),
    .B(net19),
    .Y(_0596_));
 sg13g2_nand2_1 _2820_ (.Y(_0597_),
    .A(net15),
    .B(_0452_));
 sg13g2_nor3_1 _2821_ (.A(_0596_),
    .B(_0393_),
    .C(_0597_),
    .Y(_0598_));
 sg13g2_nor2_1 _2822_ (.A(net40),
    .B(net38),
    .Y(_0599_));
 sg13g2_nand2_1 _2823_ (.Y(_0600_),
    .A(_0252_),
    .B(net54));
 sg13g2_o21ai_1 _2824_ (.B1(net40),
    .Y(_0601_),
    .A1(net65),
    .A2(_0253_));
 sg13g2_a22oi_1 _2825_ (.Y(_0602_),
    .B1(_0601_),
    .B2(net66),
    .A2(_0600_),
    .A1(_0599_));
 sg13g2_nand3b_1 _2826_ (.B(_0252_),
    .C(_0855_),
    .Y(_0603_),
    .A_N(_0223_));
 sg13g2_nand3_1 _2827_ (.B(net66),
    .C(_1367_),
    .A(_0226_),
    .Y(_0604_));
 sg13g2_a22oi_1 _2828_ (.Y(_0605_),
    .B1(_0604_),
    .B2(net55),
    .A2(_0603_),
    .A1(_1050_));
 sg13g2_o21ai_1 _2829_ (.B1(_0605_),
    .Y(_0606_),
    .A1(_0891_),
    .A2(_0246_));
 sg13g2_a21oi_1 _2830_ (.A1(net65),
    .A2(_0240_),
    .Y(_0607_),
    .B1(_0869_));
 sg13g2_a21oi_1 _2831_ (.A1(_0233_),
    .A2(_0349_),
    .Y(_0608_),
    .B1(_0867_));
 sg13g2_nor4_1 _2832_ (.A(_0602_),
    .B(_0606_),
    .C(_0607_),
    .D(_0608_),
    .Y(_0609_));
 sg13g2_o21ai_1 _2833_ (.B1(_0310_),
    .Y(_0610_),
    .A1(_0263_),
    .A2(_0312_));
 sg13g2_nand2_1 _2834_ (.Y(_0611_),
    .A(net90),
    .B(_0262_));
 sg13g2_nand2_1 _2835_ (.Y(_0612_),
    .A(_0610_),
    .B(_0611_));
 sg13g2_xnor2_1 _2836_ (.Y(_0613_),
    .A(_0609_),
    .B(_0612_));
 sg13g2_nor3_1 _2837_ (.A(_0832_),
    .B(_0304_),
    .C(_0296_),
    .Y(_0614_));
 sg13g2_a21oi_1 _2838_ (.A1(_0832_),
    .A2(_0304_),
    .Y(_0615_),
    .B1(_0614_));
 sg13g2_a22oi_1 _2839_ (.Y(_0616_),
    .B1(_0245_),
    .B2(_1012_),
    .A2(_0294_),
    .A1(_0304_));
 sg13g2_o21ai_1 _2840_ (.B1(_0616_),
    .Y(_0617_),
    .A1(_0252_),
    .A2(_0615_));
 sg13g2_nand2_1 _2841_ (.Y(_0618_),
    .A(_0283_),
    .B(_0286_));
 sg13g2_nor3_1 _2842_ (.A(net27),
    .B(_0618_),
    .C(_0240_),
    .Y(_0619_));
 sg13g2_a21o_1 _2843_ (.A2(_0618_),
    .A1(net27),
    .B1(_0619_),
    .X(_0620_));
 sg13g2_o21ai_1 _2844_ (.B1(net36),
    .Y(_0621_),
    .A1(net27),
    .A2(_0349_));
 sg13g2_a221oi_1 _2845_ (.B2(_0252_),
    .C1(_0621_),
    .B1(_0620_),
    .A1(_0618_),
    .Y(_0622_),
    .A2(_0287_));
 sg13g2_nand2_1 _2846_ (.Y(_0623_),
    .A(net53),
    .B(_1442_));
 sg13g2_o21ai_1 _2847_ (.B1(_0275_),
    .Y(_0624_),
    .A1(net90),
    .A2(_0270_));
 sg13g2_nand3_1 _2848_ (.B(_1441_),
    .C(_0624_),
    .A(net37),
    .Y(_0625_));
 sg13g2_o21ai_1 _2849_ (.B1(_0625_),
    .Y(_0626_),
    .A1(_0622_),
    .A2(_0623_));
 sg13g2_a22oi_1 _2850_ (.Y(_0627_),
    .B1(_0626_),
    .B2(net35),
    .A2(_0617_),
    .A1(_0824_));
 sg13g2_o21ai_1 _2851_ (.B1(_0627_),
    .Y(_0628_),
    .A1(net28),
    .A2(_0613_));
 sg13g2_nor2_1 _2852_ (.A(_1279_),
    .B(_0217_),
    .Y(_0629_));
 sg13g2_nand2_1 _2853_ (.Y(_0630_),
    .A(_0629_),
    .B(_0321_));
 sg13g2_xor2_1 _2854_ (.B(_0630_),
    .A(_0628_),
    .X(_0631_));
 sg13g2_nand2_1 _2855_ (.Y(_0632_),
    .A(_0465_),
    .B(_0389_));
 sg13g2_a22oi_1 _2856_ (.Y(_0633_),
    .B1(_0632_),
    .B2(_0413_),
    .A2(_0631_),
    .A1(net63));
 sg13g2_nor4_1 _2857_ (.A(net61),
    .B(_0595_),
    .C(_0598_),
    .D(_0633_),
    .Y(_0634_));
 sg13g2_a221oi_1 _2858_ (.B2(\config_regs[59] ),
    .C1(_0449_),
    .B1(net46),
    .A1(\config_regs[35] ),
    .Y(_0635_),
    .A2(_0506_));
 sg13g2_a221oi_1 _2859_ (.B2(net46),
    .C1(net61),
    .B1(\config_regs[27] ),
    .A1(net59),
    .Y(_0636_),
    .A2(net36));
 sg13g2_a22oi_1 _2860_ (.Y(_0637_),
    .B1(\config_regs[43] ),
    .B2(_0541_),
    .A2(_0336_),
    .A1(net60));
 sg13g2_nor2_1 _2861_ (.A(net88),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_nand2_1 _2862_ (.Y(_0639_),
    .A(_0437_),
    .B(net86));
 sg13g2_nand2_1 _2863_ (.Y(_0640_),
    .A(\config_regs[51] ),
    .B(_0574_));
 sg13g2_a21oi_1 _2864_ (.A1(_0639_),
    .A2(_0640_),
    .Y(_0641_),
    .B1(_0415_));
 sg13g2_nor2_1 _2865_ (.A(_0638_),
    .B(_0641_),
    .Y(_0642_));
 sg13g2_o21ai_1 _2866_ (.B1(_0642_),
    .Y(_0643_),
    .A1(_0635_),
    .A2(_0636_));
 sg13g2_a21oi_1 _2867_ (.A1(_0021_),
    .A2(_0545_),
    .Y(_0644_),
    .B1(net113));
 sg13g2_a21oi_1 _2868_ (.A1(_0643_),
    .A2(_0644_),
    .Y(_0645_),
    .B1(net30));
 sg13g2_nor2_1 _2869_ (.A(_0591_),
    .B(_0645_),
    .Y(_0646_));
 sg13g2_a22oi_1 _2870_ (.Y(_0647_),
    .B1(_0537_),
    .B2(_0646_),
    .A2(net24),
    .A1(\spi_wrapper_i.spi_reg_inst.tx_buffer[3] ));
 sg13g2_o21ai_1 _2871_ (.B1(_0647_),
    .Y(_0134_),
    .A1(_0594_),
    .A2(_0634_));
 sg13g2_nor2_1 _2872_ (.A(_0389_),
    .B(net15),
    .Y(_0648_));
 sg13g2_o21ai_1 _2873_ (.B1(net21),
    .Y(_0649_),
    .A1(_0371_),
    .A2(_0648_));
 sg13g2_nor2_1 _2874_ (.A(_0389_),
    .B(_0212_),
    .Y(_0650_));
 sg13g2_nor2_1 _2875_ (.A(_0650_),
    .B(_0454_),
    .Y(_0651_));
 sg13g2_nand2b_1 _2876_ (.Y(_0652_),
    .B(net63),
    .A_N(net12));
 sg13g2_nand3_1 _2877_ (.B(net61),
    .C(_0652_),
    .A(net64),
    .Y(_0653_));
 sg13g2_o21ai_1 _2878_ (.B1(_0653_),
    .Y(_0654_),
    .A1(net64),
    .A2(_0511_));
 sg13g2_a22oi_1 _2879_ (.Y(_0655_),
    .B1(_0654_),
    .B2(_0429_),
    .A2(_0651_),
    .A1(_0649_));
 sg13g2_xnor2_1 _2880_ (.Y(_0656_),
    .A(_0950_),
    .B(net22));
 sg13g2_nor2_1 _2881_ (.A(_0205_),
    .B(_0507_),
    .Y(_0657_));
 sg13g2_o21ai_1 _2882_ (.B1(_0657_),
    .Y(_0658_),
    .A1(_0925_),
    .A2(_0656_));
 sg13g2_a21oi_1 _2883_ (.A1(_0010_),
    .A2(net30),
    .Y(_0659_),
    .B1(_0538_));
 sg13g2_nand2_1 _2884_ (.Y(_0660_),
    .A(_0658_),
    .B(_0659_));
 sg13g2_a221oi_1 _2885_ (.B2(\config_regs[60] ),
    .C1(net60),
    .B1(net46),
    .A1(\config_regs[36] ),
    .Y(_0661_),
    .A2(_0506_));
 sg13g2_inv_1 _2886_ (.Y(_0662_),
    .A(_0018_));
 sg13g2_a221oi_1 _2887_ (.B2(\config_regs[28] ),
    .C1(net61),
    .B1(net46),
    .A1(net59),
    .Y(_0663_),
    .A2(_0662_));
 sg13g2_a22oi_1 _2888_ (.Y(_0664_),
    .B1(\config_regs[44] ),
    .B2(_0541_),
    .A2(_0221_),
    .A1(net60));
 sg13g2_nor2_1 _2889_ (.A(_0412_),
    .B(_0664_),
    .Y(_0665_));
 sg13g2_nand2_1 _2890_ (.Y(_0666_),
    .A(\config_regs[52] ),
    .B(_0574_));
 sg13g2_a21oi_1 _2891_ (.A1(_0639_),
    .A2(_0666_),
    .Y(_0667_),
    .B1(_0415_));
 sg13g2_nor2_1 _2892_ (.A(_0665_),
    .B(_0667_),
    .Y(_0668_));
 sg13g2_o21ai_1 _2893_ (.B1(_0668_),
    .Y(_0669_),
    .A1(_0661_),
    .A2(_0663_));
 sg13g2_a21oi_1 _2894_ (.A1(_0894_),
    .A2(net43),
    .Y(_0670_),
    .B1(net113));
 sg13g2_a21oi_1 _2895_ (.A1(_0669_),
    .A2(_0670_),
    .Y(_0671_),
    .B1(net30));
 sg13g2_a21oi_1 _2896_ (.A1(_0010_),
    .A2(net30),
    .Y(_0672_),
    .B1(_0671_));
 sg13g2_a22oi_1 _2897_ (.Y(_0673_),
    .B1(_0537_),
    .B2(_0672_),
    .A2(net24),
    .A1(\spi_wrapper_i.spi_reg_inst.tx_buffer[4] ));
 sg13g2_o21ai_1 _2898_ (.B1(_0673_),
    .Y(_0135_),
    .A1(_0655_),
    .A2(_0660_));
 sg13g2_a21oi_1 _2899_ (.A1(_0402_),
    .A2(_0404_),
    .Y(_0674_),
    .B1(net61));
 sg13g2_nor2_1 _2900_ (.A(_0950_),
    .B(net22),
    .Y(_0675_));
 sg13g2_xor2_1 _2901_ (.B(_0675_),
    .A(_0924_),
    .X(_0676_));
 sg13g2_nand2_1 _2902_ (.Y(_0677_),
    .A(_0953_),
    .B(_0676_));
 sg13g2_nor2_1 _2903_ (.A(_1332_),
    .B(_0507_),
    .Y(_0678_));
 sg13g2_a221oi_1 _2904_ (.B2(_0678_),
    .C1(_0538_),
    .B1(_0677_),
    .A1(_0011_),
    .Y(_0679_),
    .A2(net44));
 sg13g2_or2_1 _2905_ (.X(_0680_),
    .B(net13),
    .A(_0461_));
 sg13g2_nand3_1 _2906_ (.B(_0679_),
    .C(_0680_),
    .A(_0452_),
    .Y(_0681_));
 sg13g2_mux4_1 _2907_ (.S0(_0437_),
    .A0(_0019_),
    .A1(_0023_),
    .A2(_0458_),
    .A3(_0026_),
    .S1(net121),
    .X(_0682_));
 sg13g2_mux4_1 _2908_ (.S0(net121),
    .A0(\config_regs[37] ),
    .A1(\config_regs[45] ),
    .A2(\config_regs[53] ),
    .A3(\config_regs[61] ),
    .S1(_0411_),
    .X(_0683_));
 sg13g2_nand2_1 _2909_ (.Y(_0684_),
    .A(_0439_),
    .B(_0683_));
 sg13g2_o21ai_1 _2910_ (.B1(_0684_),
    .Y(_0685_),
    .A1(_0439_),
    .A2(_0682_));
 sg13g2_a21oi_1 _2911_ (.A1(_0476_),
    .A2(_0685_),
    .Y(_0686_),
    .B1(net44));
 sg13g2_a21oi_1 _2912_ (.A1(_0011_),
    .A2(_0503_),
    .Y(_0687_),
    .B1(_0686_));
 sg13g2_and2_1 _2913_ (.A(_0537_),
    .B(_0687_),
    .X(_0688_));
 sg13g2_a221oi_1 _2914_ (.B2(_0679_),
    .C1(_0688_),
    .B1(net43),
    .A1(\spi_wrapper_i.spi_reg_inst.tx_buffer[5] ),
    .Y(_0689_),
    .A2(_0533_));
 sg13g2_o21ai_1 _2915_ (.B1(_0689_),
    .Y(_0136_),
    .A1(_0674_),
    .A2(_0681_));
 sg13g2_nand2_1 _2916_ (.Y(_0690_),
    .A(\spi_wrapper_i.spi_reg_inst.tx_buffer[6] ),
    .B(net24));
 sg13g2_a21oi_1 _2917_ (.A1(_0012_),
    .A2(_0535_),
    .Y(_0691_),
    .B1(_0536_));
 sg13g2_nand2b_1 _2918_ (.Y(_0692_),
    .B(_0691_),
    .A_N(net24));
 sg13g2_nor2_1 _2919_ (.A(net62),
    .B(net87),
    .Y(_0693_));
 sg13g2_a22oi_1 _2920_ (.Y(_0694_),
    .B1(_0554_),
    .B2(\config_regs[46] ),
    .A2(_0693_),
    .A1(\config_regs[54] ));
 sg13g2_mux2_1 _2921_ (.A0(\config_regs[62] ),
    .A1(\config_regs[30] ),
    .S(net86),
    .X(_0695_));
 sg13g2_nand2b_1 _2922_ (.Y(_0696_),
    .B(_0411_),
    .A_N(\config_regs[22] ));
 sg13g2_nor2_1 _2923_ (.A(_0029_),
    .B(_0429_),
    .Y(_0697_));
 sg13g2_a21oi_1 _2924_ (.A1(\config_regs[38] ),
    .A2(_0511_),
    .Y(_0698_),
    .B1(_0697_));
 sg13g2_nor2_1 _2925_ (.A(net88),
    .B(_0698_),
    .Y(_0699_));
 sg13g2_a221oi_1 _2926_ (.B2(_0542_),
    .C1(_0699_),
    .B1(_0696_),
    .A1(net46),
    .Y(_0700_),
    .A2(_0695_));
 sg13g2_o21ai_1 _2927_ (.B1(_0700_),
    .Y(_0701_),
    .A1(net45),
    .A2(_0694_));
 sg13g2_a21oi_1 _2928_ (.A1(_0028_),
    .A2(net43),
    .Y(_0702_),
    .B1(net113));
 sg13g2_a221oi_1 _2929_ (.B2(_0702_),
    .C1(net44),
    .B1(_0701_),
    .A1(_0762_),
    .Y(_0703_),
    .A2(\spi_wrapper_i.spi_reg_inst.tx_buffer[6] ));
 sg13g2_nor4_1 _2930_ (.A(_1025_),
    .B(_1062_),
    .C(net56),
    .D(_1064_),
    .Y(_0704_));
 sg13g2_nand3_1 _2931_ (.B(_1027_),
    .C(_0704_),
    .A(_0980_),
    .Y(_0705_));
 sg13g2_or4_1 _2932_ (.A(_0440_),
    .B(_1066_),
    .C(_1235_),
    .D(_0705_),
    .X(_0706_));
 sg13g2_nand3_1 _2933_ (.B(net63),
    .C(_0706_),
    .A(net62),
    .Y(_0707_));
 sg13g2_o21ai_1 _2934_ (.B1(_0440_),
    .Y(_0708_),
    .A1(net59),
    .A2(net14));
 sg13g2_nand2_1 _2935_ (.Y(_0709_),
    .A(_0413_),
    .B(_0708_));
 sg13g2_nor2_1 _2936_ (.A(net21),
    .B(net15),
    .Y(_0710_));
 sg13g2_a21oi_1 _2937_ (.A1(_0650_),
    .A2(_0710_),
    .Y(_0711_),
    .B1(_0454_));
 sg13g2_and2_1 _2938_ (.A(net16),
    .B(net20),
    .X(_0712_));
 sg13g2_o21ai_1 _2939_ (.B1(net21),
    .Y(_0713_),
    .A1(_0712_),
    .A2(_0385_));
 sg13g2_a22oi_1 _2940_ (.Y(_0714_),
    .B1(_0711_),
    .B2(_0713_),
    .A2(_0709_),
    .A1(_0707_));
 sg13g2_and2_1 _2941_ (.A(_0924_),
    .B(_0675_),
    .X(_0715_));
 sg13g2_xnor2_1 _2942_ (.Y(_0716_),
    .A(_1411_),
    .B(_0715_));
 sg13g2_nor2_1 _2943_ (.A(_1440_),
    .B(_0507_),
    .Y(_0717_));
 sg13g2_o21ai_1 _2944_ (.B1(_0717_),
    .Y(_0718_),
    .A1(_0925_),
    .A2(_0716_));
 sg13g2_inv_1 _2945_ (.Y(_0719_),
    .A(_0703_));
 sg13g2_a21oi_1 _2946_ (.A1(_0475_),
    .A2(_0718_),
    .Y(_0720_),
    .B1(_0719_));
 sg13g2_a221oi_1 _2947_ (.B2(_0714_),
    .C1(_0720_),
    .B1(_0703_),
    .A1(_0690_),
    .Y(_0137_),
    .A2(_0692_));
 sg13g2_o21ai_1 _2948_ (.B1(_0416_),
    .Y(_0721_),
    .A1(net61),
    .A2(net22));
 sg13g2_xnor2_1 _2949_ (.Y(_0722_),
    .A(_0629_),
    .B(_0321_));
 sg13g2_a21oi_1 _2950_ (.A1(_0359_),
    .A2(_0360_),
    .Y(_0723_),
    .B1(_0507_));
 sg13g2_o21ai_1 _2951_ (.B1(_0723_),
    .Y(_0724_),
    .A1(_0925_),
    .A2(_0722_));
 sg13g2_nand4_1 _2952_ (.B(net113),
    .C(_0721_),
    .A(_0438_),
    .Y(_0725_),
    .D(_0724_));
 sg13g2_mux2_1 _2953_ (.A0(\config_regs[55] ),
    .A1(\config_regs[63] ),
    .S(net87),
    .X(_0726_));
 sg13g2_a22oi_1 _2954_ (.Y(_0727_),
    .B1(_0726_),
    .B2(net88),
    .A2(_0554_),
    .A1(\config_regs[47] ));
 sg13g2_o21ai_1 _2955_ (.B1(net59),
    .Y(_0728_),
    .A1(net86),
    .A2(\config_regs[39] ));
 sg13g2_o21ai_1 _2956_ (.B1(_0728_),
    .Y(_0729_),
    .A1(_0439_),
    .A2(_0005_));
 sg13g2_mux2_1 _2957_ (.A0(\config_regs[23] ),
    .A1(\config_regs[31] ),
    .S(net87),
    .X(_0730_));
 sg13g2_a22oi_1 _2958_ (.Y(_0731_),
    .B1(_0730_),
    .B2(_0524_),
    .A2(_0729_),
    .A1(net62));
 sg13g2_o21ai_1 _2959_ (.B1(_0731_),
    .Y(_0732_),
    .A1(net45),
    .A2(_0727_));
 sg13g2_a21oi_1 _2960_ (.A1(_0218_),
    .A2(net43),
    .Y(_0733_),
    .B1(net113));
 sg13g2_a21oi_1 _2961_ (.A1(_0732_),
    .A2(_0733_),
    .Y(_0734_),
    .B1(net30));
 sg13g2_a221oi_1 _2962_ (.B2(_0734_),
    .C1(_0548_),
    .B1(_0725_),
    .A1(_0013_),
    .Y(_0735_),
    .A2(net30));
 sg13g2_a21o_1 _2963_ (.A2(net24),
    .A1(spi_miso),
    .B1(_0735_),
    .X(_0138_));
 sg13g2_nor2_1 _2964_ (.A(_0756_),
    .B(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .Y(_0736_));
 sg13g2_a21oi_1 _2965_ (.A1(_0755_),
    .A2(_0736_),
    .Y(_0737_),
    .B1(_0757_));
 sg13g2_mux2_1 _2966_ (.A0(_0757_),
    .A1(_0737_),
    .S(_0491_),
    .X(_0139_));
 sg13g2_nand2_1 _2967_ (.Y(_0738_),
    .A(_0757_),
    .B(_0491_));
 sg13g2_xnor2_1 _2968_ (.Y(_0140_),
    .A(_0756_),
    .B(_0738_));
 sg13g2_nand3_1 _2969_ (.B(_0757_),
    .C(_0491_),
    .A(_0756_),
    .Y(_0739_));
 sg13g2_xnor2_1 _2970_ (.Y(_0141_),
    .A(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .B(_0739_));
 sg13g2_and4_1 _2971_ (.A(_0756_),
    .B(_0757_),
    .C(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .D(_0489_),
    .X(_0740_));
 sg13g2_a21o_1 _2972_ (.A2(_0740_),
    .A1(_0755_),
    .B1(_0758_),
    .X(_0741_));
 sg13g2_a21oi_1 _2973_ (.A1(net85),
    .A2(_0740_),
    .Y(_0742_),
    .B1(_0755_));
 sg13g2_a21oi_1 _2974_ (.A1(_0397_),
    .A2(_0741_),
    .Y(_0142_),
    .B1(_0742_));
 sg13g2_mux2_1 _2975_ (.A0(\synchronizer_spi_clk_inst.data_sync[1] ),
    .A1(net5),
    .S(net89),
    .X(_0143_));
 sg13g2_mux2_1 _2976_ (.A0(spi_clk_sync),
    .A1(\synchronizer_spi_clk_inst.data_sync[1] ),
    .S(net89),
    .X(_0144_));
 sg13g2_mux2_1 _2977_ (.A0(\synchronizer_spi_cs_n_inst.data_sync[1] ),
    .A1(net4),
    .S(net89),
    .X(_0145_));
 sg13g2_mux2_1 _2978_ (.A0(_0753_),
    .A1(\synchronizer_spi_cs_n_inst.data_sync[1] ),
    .S(net89),
    .X(_0146_));
 sg13g2_mux2_1 _2979_ (.A0(\synchronizer_spi_mode_cpha.data_sync[1] ),
    .A1(net3),
    .S(net85),
    .X(_0147_));
 sg13g2_mux2_1 _2980_ (.A0(cpha_sync),
    .A1(\synchronizer_spi_mode_cpha.data_sync[1] ),
    .S(net85),
    .X(_0148_));
 sg13g2_mux2_1 _2981_ (.A0(\synchronizer_spi_mode_cpol.data_sync[1] ),
    .A1(net2),
    .S(_0483_),
    .X(_0149_));
 sg13g2_mux2_1 _2982_ (.A0(cpol_sync),
    .A1(\synchronizer_spi_mode_cpol.data_sync[1] ),
    .S(_0483_),
    .X(_0150_));
 sg13g2_mux2_1 _2983_ (.A0(\synchronizer_spi_mosi_inst.data_sync[1] ),
    .A1(net6),
    .S(net85),
    .X(_0151_));
 sg13g2_mux2_1 _2984_ (.A0(spi_mosi_sync),
    .A1(\synchronizer_spi_mosi_inst.data_sync[1] ),
    .S(net85),
    .X(_0152_));
 sg13g2_nor3_1 _2985_ (.A(_0752_),
    .B(_0776_),
    .C(_0769_),
    .Y(_0743_));
 sg13g2_o21ai_1 _2986_ (.B1(_0753_),
    .Y(_0744_),
    .A1(\spi_wrapper_i.spi_reg_inst.state[0] ),
    .A2(_0743_));
 sg13g2_nand2_1 _2987_ (.Y(_0745_),
    .A(net132),
    .B(_0752_));
 sg13g2_nor2_1 _2988_ (.A(_0780_),
    .B(_0478_),
    .Y(_0746_));
 sg13g2_a21oi_1 _2989_ (.A1(\spi_wrapper_i.spi_reg_inst.state[0] ),
    .A2(_0745_),
    .Y(_0747_),
    .B1(_0746_));
 sg13g2_nand3_1 _2990_ (.B(\spi_wrapper_i.spi_reg_inst.state[1] ),
    .C(_0759_),
    .A(net85),
    .Y(_0748_));
 sg13g2_and3_1 _2991_ (.X(_0031_),
    .A(_0744_),
    .B(_0747_),
    .C(_0748_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _2994__166 (.L_HI(net166));
 sg13g2_buf_1 _2994_ (.A(net166),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2995_ (.A(net167),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2996_ (.A(net168),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2997_ (.A(net169),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2998_ (.A(net155),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2999_ (.A(net156),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3000_ (.A(net157),
    .X(uio_oe[6]));
 sg13g2_buf_1 _3001_ (.A(net170),
    .X(uio_oe[7]));
 sg13g2_buf_1 _3002_ (.A(net158),
    .X(uio_out[0]));
 sg13g2_buf_1 _3003_ (.A(net159),
    .X(uio_out[1]));
 sg13g2_buf_1 _3004_ (.A(net160),
    .X(uio_out[2]));
 sg13g2_buf_1 _3005_ (.A(spi_miso),
    .X(net7));
 sg13g2_buf_1 _3006_ (.A(net161),
    .X(uio_out[4]));
 sg13g2_buf_1 _3007_ (.A(net162),
    .X(uio_out[5]));
 sg13g2_buf_1 _3008_ (.A(net163),
    .X(uio_out[6]));
 sg13g2_buf_1 _3009_ (.A(net164),
    .X(uio_out[7]));
 sg13g2_buf_1 _3010_ (.A(net165),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \reclocking_7seg.data_sync[0]$_DFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net150),
    .D(_0032_),
    .Q_N(_1553_),
    .Q(net8));
 sg13g2_dfrbp_1 \reclocking_7seg.data_sync[1]$_DFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net148),
    .D(_0033_),
    .Q_N(_1552_),
    .Q(net9));
 sg13g2_dfrbp_1 \reclocking_7seg.data_sync[2]$_DFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net150),
    .D(_0034_),
    .Q_N(_1551_),
    .Q(net10));
 sg13g2_dfrbp_1 \reclocking_7seg.data_sync[3]$_DFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net147),
    .D(_0035_),
    .Q_N(_1550_),
    .Q(net11));
 sg13g2_dfrbp_1 \reclocking_7seg.data_sync[4]$_DFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net150),
    .D(_0036_),
    .Q_N(_1549_),
    .Q(net12));
 sg13g2_dfrbp_1 \reclocking_7seg.data_sync[5]$_DFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net150),
    .D(_0037_),
    .Q_N(_1548_),
    .Q(net13));
 sg13g2_dfrbp_1 \reclocking_7seg.data_sync[6]$_DFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net150),
    .D(_0038_),
    .Q_N(_1547_),
    .Q(net14));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[0][0]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net147),
    .D(_0039_),
    .Q_N(_0016_),
    .Q(\alu_74181_i0.a[0] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[0][1]$_DFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net147),
    .D(_0040_),
    .Q_N(_0022_),
    .Q(\alu_74181_i0.a[1] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[0][2]$_DFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net147),
    .D(_0041_),
    .Q_N(_0020_),
    .Q(\alu_74181_i0.a[2] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[0][3]$_DFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net147),
    .D(_0042_),
    .Q_N(_0021_),
    .Q(\alu_74181_i0.a[3] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[0][4]$_DFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net133),
    .D(_0043_),
    .Q_N(_0024_),
    .Q(\alu_74181_i1.a[0] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[0][5]$_DFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net133),
    .D(_0044_),
    .Q_N(_0023_),
    .Q(\alu_74181_i1.a[1] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[0][6]$_DFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net133),
    .D(_0045_),
    .Q_N(_0028_),
    .Q(\alu_74181_i1.a[2] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[0][7]$_DFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net134),
    .D(_0046_),
    .Q_N(_0004_),
    .Q(\alu_74181_i1.a[3] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[1][0]$_DFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net134),
    .D(_0047_),
    .Q_N(_0017_),
    .Q(\alu_74181_i0.alu_74181_arith_inst.b[0] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[1][1]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net154),
    .D(_0048_),
    .Q_N(_0027_),
    .Q(\alu_74181_i0.alu_74181_arith_inst.b[1] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[1][2]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net154),
    .D(_0049_),
    .Q_N(_0030_),
    .Q(\alu_74181_i0.alu_74181_arith_inst.b[2] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[1][3]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net154),
    .D(_0050_),
    .Q_N(_0006_),
    .Q(\alu_74181_i0.alu_74181_arith_inst.b[3] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[1][4]$_DFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net133),
    .D(_0051_),
    .Q_N(_0025_),
    .Q(\alu_74181_i1.alu_74181_arith_inst.b[0] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[1][5]$_DFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net133),
    .D(_0052_),
    .Q_N(_0026_),
    .Q(\alu_74181_i1.alu_74181_arith_inst.b[1] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[1][6]$_DFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net133),
    .D(_0053_),
    .Q_N(_0029_),
    .Q(\alu_74181_i1.alu_74181_arith_inst.b[2] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[1][7]$_DFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net134),
    .D(_0054_),
    .Q_N(_0005_),
    .Q(\alu_74181_i1.alu_74181_arith_inst.b[3] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[2][0]$_DFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net133),
    .D(_0055_),
    .Q_N(_1546_),
    .Q(\alu_74181_i0.alu_74181_arith_inst.s[0] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[2][1]$_DFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net134),
    .D(_0056_),
    .Q_N(_1545_),
    .Q(\alu_74181_i0.alu_74181_arith_inst.s[1] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[2][2]$_DFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net133),
    .D(_0057_),
    .Q_N(_1544_),
    .Q(\alu_74181_i0.alu_74181_arith_inst.s[2] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[2][3]$_DFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net138),
    .D(_0058_),
    .Q_N(_1543_),
    .Q(\alu_74181_i0.alu_74181_arith_inst.s[3] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[2][4]$_DFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net138),
    .D(_0059_),
    .Q_N(_0018_),
    .Q(\alu_74181_i0.m ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[2][5]$_DFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net135),
    .D(_0060_),
    .Q_N(_0019_),
    .Q(\alu_74181_i0.alu_74181_arith_inst.cn ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[2][6]$_DFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net136),
    .D(_0061_),
    .Q_N(_1542_),
    .Q(\config_regs[22] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[2][7]$_DFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net135),
    .D(_0062_),
    .Q_N(_1541_),
    .Q(\config_regs[23] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[3][0]$_DFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net138),
    .D(_0063_),
    .Q_N(_1540_),
    .Q(\config_regs[24] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[3][1]$_DFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net135),
    .D(_0064_),
    .Q_N(_1539_),
    .Q(\config_regs[25] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[3][2]$_DFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net138),
    .D(_0065_),
    .Q_N(_1538_),
    .Q(\config_regs[26] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[3][3]$_DFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net138),
    .D(_0066_),
    .Q_N(_1537_),
    .Q(\config_regs[27] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[3][4]$_DFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net138),
    .D(_0067_),
    .Q_N(_1536_),
    .Q(\config_regs[28] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[3][5]$_DFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net135),
    .D(_0068_),
    .Q_N(_1535_),
    .Q(\config_regs[29] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[3][6]$_DFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net136),
    .D(_0069_),
    .Q_N(_1534_),
    .Q(\config_regs[30] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[3][7]$_DFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net135),
    .D(_0070_),
    .Q_N(_1533_),
    .Q(\config_regs[31] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[4][0]$_DFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net139),
    .D(_0071_),
    .Q_N(_1532_),
    .Q(\config_regs[32] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[4][1]$_DFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net141),
    .D(_0072_),
    .Q_N(_1531_),
    .Q(\config_regs[33] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[4][2]$_DFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net143),
    .D(_0073_),
    .Q_N(_1530_),
    .Q(\config_regs[34] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[4][3]$_DFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net145),
    .D(_0074_),
    .Q_N(_1529_),
    .Q(\config_regs[35] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[4][4]$_DFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net145),
    .D(_0075_),
    .Q_N(_1528_),
    .Q(\config_regs[36] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[4][5]$_DFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net140),
    .D(_0076_),
    .Q_N(_1527_),
    .Q(\config_regs[37] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[4][6]$_DFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net139),
    .D(_0077_),
    .Q_N(_1526_),
    .Q(\config_regs[38] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[4][7]$_DFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net142),
    .D(_0078_),
    .Q_N(_1525_),
    .Q(\config_regs[39] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[5][0]$_DFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net136),
    .D(_0079_),
    .Q_N(_1524_),
    .Q(\config_regs[40] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[5][1]$_DFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net135),
    .D(_0080_),
    .Q_N(_1523_),
    .Q(\config_regs[41] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[5][2]$_DFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net148),
    .D(_0081_),
    .Q_N(_1522_),
    .Q(\config_regs[42] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[5][3]$_DFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net148),
    .D(_0082_),
    .Q_N(_1521_),
    .Q(\config_regs[43] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[5][4]$_DFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net136),
    .D(_0083_),
    .Q_N(_1520_),
    .Q(\config_regs[44] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[5][5]$_DFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net139),
    .D(_0084_),
    .Q_N(_1519_),
    .Q(\config_regs[45] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[5][6]$_DFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net142),
    .D(_0085_),
    .Q_N(_1518_),
    .Q(\config_regs[46] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[5][7]$_DFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net139),
    .D(_0086_),
    .Q_N(_1517_),
    .Q(\config_regs[47] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[6][0]$_DFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net145),
    .D(_0087_),
    .Q_N(_1516_),
    .Q(\config_regs[48] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[6][1]$_DFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net139),
    .D(_0088_),
    .Q_N(_1515_),
    .Q(\config_regs[49] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[6][2]$_DFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net145),
    .D(_0089_),
    .Q_N(_1514_),
    .Q(\config_regs[50] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[6][3]$_DFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net145),
    .D(_0090_),
    .Q_N(_1513_),
    .Q(\config_regs[51] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[6][4]$_DFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net145),
    .D(_0091_),
    .Q_N(_1512_),
    .Q(\config_regs[52] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[6][5]$_DFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net139),
    .D(_0092_),
    .Q_N(_1511_),
    .Q(\config_regs[53] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[6][6]$_DFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net142),
    .D(_0093_),
    .Q_N(_1510_),
    .Q(\config_regs[54] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[6][7]$_DFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net139),
    .D(_0094_),
    .Q_N(_1509_),
    .Q(\config_regs[55] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[7][0]$_DFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net138),
    .D(_0095_),
    .Q_N(_1508_),
    .Q(\config_regs[56] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[7][1]$_DFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net135),
    .D(_0096_),
    .Q_N(_1507_),
    .Q(\config_regs[57] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[7][2]$_DFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net148),
    .D(_0097_),
    .Q_N(_1506_),
    .Q(\config_regs[58] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[7][3]$_DFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net145),
    .D(_0098_),
    .Q_N(_1505_),
    .Q(\config_regs[59] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[7][4]$_DFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net145),
    .D(_0099_),
    .Q_N(_1504_),
    .Q(\config_regs[60] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[7][5]$_DFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net140),
    .D(_0100_),
    .Q_N(_1503_),
    .Q(\config_regs[61] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[7][6]$_DFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net135),
    .D(_0101_),
    .Q_N(_1502_),
    .Q(\config_regs[62] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.config_mem[7][7]$_DFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net139),
    .D(_0102_),
    .Q_N(_1501_),
    .Q(\config_regs[63] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.addr[0]$_DFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net143),
    .D(_0103_),
    .Q_N(_1500_),
    .Q(\spi_wrapper_i.reg_addr[0] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.addr[1]$_DFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net143),
    .D(_0104_),
    .Q_N(_1499_),
    .Q(\spi_wrapper_i.reg_addr[1] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.addr[2]$_DFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net143),
    .D(_0105_),
    .Q_N(_0015_),
    .Q(\spi_wrapper_i.reg_addr[2] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.addr[3]$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net143),
    .D(_0106_),
    .Q_N(_1498_),
    .Q(\spi_wrapper_i.reg_addr[3] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.data[0]$_DFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net141),
    .D(_0107_),
    .Q_N(_1497_),
    .Q(\spi_wrapper_i.reg_data_o[0] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.data[1]$_DFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net141),
    .D(_0108_),
    .Q_N(_1496_),
    .Q(\spi_wrapper_i.reg_data_o[1] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.data[2]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net143),
    .D(_0109_),
    .Q_N(_1495_),
    .Q(\spi_wrapper_i.reg_data_o[2] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.data[3]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net144),
    .D(_0110_),
    .Q_N(_1494_),
    .Q(\spi_wrapper_i.reg_data_o[3] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.data[4]$_DFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net140),
    .D(_0111_),
    .Q_N(_1493_),
    .Q(\spi_wrapper_i.reg_data_o[4] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.data[5]$_DFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net140),
    .D(_0112_),
    .Q_N(_1492_),
    .Q(\spi_wrapper_i.reg_data_o[5] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.data[6]$_DFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net140),
    .D(_0113_),
    .Q_N(_1491_),
    .Q(\spi_wrapper_i.reg_data_o[6] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.data[7]$_DFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net140),
    .D(_0114_),
    .Q_N(_1490_),
    .Q(\spi_wrapper_i.reg_data_o[7] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.dv$_DFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net149),
    .D(_0115_),
    .Q_N(_1489_),
    .Q(\spi_wrapper_i.reg_data_o_vld ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.reg_rw$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net144),
    .D(_0116_),
    .Q_N(_1488_),
    .Q(\spi_wrapper_i.spi_reg_inst.reg_rw ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rising_edge_detector_eof.data_dly$_DFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net148),
    .D(_0117_),
    .Q_N(_1487_),
    .Q(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rising_edge_detector_spi_clk.data_dly$_DFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net151),
    .D(_0118_),
    .Q_N(_1486_),
    .Q(\spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rx_buffer[0]$_DFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net151),
    .D(_0119_),
    .Q_N(_1485_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[0] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rx_buffer[1]$_DFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net141),
    .D(_0120_),
    .Q_N(_1484_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[1] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rx_buffer[2]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net143),
    .D(_0121_),
    .Q_N(_1483_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[2] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rx_buffer[3]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net143),
    .D(_0122_),
    .Q_N(_1482_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[3] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rx_buffer[4]$_DFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net141),
    .D(_0123_),
    .Q_N(_1481_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[4] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rx_buffer[5]$_DFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net140),
    .D(_0124_),
    .Q_N(_1480_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[5] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rx_buffer[6]$_DFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net140),
    .D(_0125_),
    .Q_N(_1479_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[6] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rx_buffer[7]$_DFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net141),
    .D(_0126_),
    .Q_N(_1478_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer[7] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0]$_DFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net149),
    .D(_0127_),
    .Q_N(_1477_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1]$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net144),
    .D(_0128_),
    .Q_N(_1476_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2]$_DFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net149),
    .D(_0129_),
    .Q_N(_1475_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3]$_DFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net144),
    .D(_0130_),
    .Q_N(_1474_),
    .Q(\spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.state[0]$_DFF_PN1_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net149),
    .D(_0031_),
    .Q_N(\spi_wrapper_i.spi_reg_inst.state[0] ),
    .Q(_1557_));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.state[1]$_DFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net149),
    .D(_0000_),
    .Q_N(_1554_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[1] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.state[2]$_DFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net144),
    .D(_0001_),
    .Q_N(_1555_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[2] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.state[3]$_DFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net151),
    .D(_0002_),
    .Q_N(_1556_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[3] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.state[4]$_DFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net149),
    .D(_0003_),
    .Q_N(_1473_),
    .Q(\spi_wrapper_i.spi_reg_inst.state[4] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.tx_buffer[0]$_DFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net148),
    .D(_0131_),
    .Q_N(_0007_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[0] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.tx_buffer[1]$_DFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net148),
    .D(_0132_),
    .Q_N(_0008_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[1] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.tx_buffer[2]$_DFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net150),
    .D(_0133_),
    .Q_N(_0009_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[2] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.tx_buffer[3]$_DFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net147),
    .D(_0134_),
    .Q_N(_0010_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[3] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.tx_buffer[4]$_DFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net147),
    .D(_0135_),
    .Q_N(_0011_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[4] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.tx_buffer[5]$_DFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net150),
    .D(_0136_),
    .Q_N(_0012_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[5] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.tx_buffer[6]$_DFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net147),
    .D(_0137_),
    .Q_N(_0013_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer[6] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.tx_buffer[7]$_DFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net148),
    .D(_0138_),
    .Q_N(_1472_),
    .Q(spi_miso));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0]$_DFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net151),
    .D(_0139_),
    .Q_N(_1471_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1]$_DFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net151),
    .D(_0140_),
    .Q_N(_1470_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2]$_DFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net152),
    .D(_0141_),
    .Q_N(_1469_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ));
 sg13g2_dfrbp_1 \spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3]$_DFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net152),
    .D(_0142_),
    .Q_N(_1468_),
    .Q(\spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ));
 sg13g2_dfrbp_1 \synchronizer_spi_clk_inst.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net150),
    .D(_0143_),
    .Q_N(_1467_),
    .Q(\synchronizer_spi_clk_inst.data_sync[1] ));
 sg13g2_dfrbp_1 \synchronizer_spi_clk_inst.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net153),
    .D(_0144_),
    .Q_N(_1466_),
    .Q(spi_clk_sync));
 sg13g2_dfrbp_1 \synchronizer_spi_cs_n_inst.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net151),
    .D(_0145_),
    .Q_N(_1465_),
    .Q(\synchronizer_spi_cs_n_inst.data_sync[1] ));
 sg13g2_dfrbp_1 \synchronizer_spi_cs_n_inst.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net151),
    .D(_0146_),
    .Q_N(_0014_),
    .Q(spi_cs_n_sync));
 sg13g2_dfrbp_1 \synchronizer_spi_mode_cpha.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net152),
    .D(_0147_),
    .Q_N(_1464_),
    .Q(\synchronizer_spi_mode_cpha.data_sync[1] ));
 sg13g2_dfrbp_1 \synchronizer_spi_mode_cpha.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net152),
    .D(_0148_),
    .Q_N(_1463_),
    .Q(cpha_sync));
 sg13g2_dfrbp_1 \synchronizer_spi_mode_cpol.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net152),
    .D(_0149_),
    .Q_N(_1462_),
    .Q(\synchronizer_spi_mode_cpol.data_sync[1] ));
 sg13g2_dfrbp_1 \synchronizer_spi_mode_cpol.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net152),
    .D(_0150_),
    .Q_N(_1461_),
    .Q(cpol_sync));
 sg13g2_dfrbp_1 \synchronizer_spi_mosi_inst.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net149),
    .D(_0151_),
    .Q_N(_1460_),
    .Q(\synchronizer_spi_mosi_inst.data_sync[1] ));
 sg13g2_dfrbp_1 \synchronizer_spi_mosi_inst.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net151),
    .D(_0152_),
    .Q_N(_1459_),
    .Q(spi_mosi_sync));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[4]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[5]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[6]),
    .X(net6));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[3]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[0]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[1]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[2]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[3]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[4]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[5]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[6]));
 sg13g2_buf_2 fanout15 (.A(_0382_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0367_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0381_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0215_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0212_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0162_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_1337_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_1279_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0456_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0533_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1292_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0463_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0965_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0920_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0794_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0535_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0493_),
    .X(net31));
 sg13g2_buf_4 fanout32 (.X(net32),
    .A(_0480_));
 sg13g2_buf_2 fanout33 (.A(_0442_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0431_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1321_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1296_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1294_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1069_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1048_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0873_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0808_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0771_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0545_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0503_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0461_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0452_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1306_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1303_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1302_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1295_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_1293_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_1260_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1259_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1073_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1056_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1023_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0961_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0937_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0465_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0449_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0440_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0438_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0416_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0413_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0271_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0244_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1358_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1344_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1320_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1189_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0963_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0958_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0953_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0936_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0864_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0853_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0835_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0822_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0820_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0817_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0815_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0806_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0801_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0797_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0483_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0448_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0415_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0412_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0397_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0230_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0220_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_1355_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_1343_),
    .X(net93));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(_1283_));
 sg13g2_buf_2 fanout95 (.A(_1138_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_1057_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_1031_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_1021_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_1020_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_0969_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_0967_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_0957_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_0877_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_0827_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_0825_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_0811_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_0805_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_0803_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_0796_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_0790_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_0783_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_0763_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_0475_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0427_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_0426_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_0425_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_0424_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_0423_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_0422_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_0421_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_0414_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_0410_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_0982_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_0979_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_0974_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_0971_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_0968_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_0966_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_0785_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_0784_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_0782_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_0750_),
    .X(net132));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(net137));
 sg13g2_buf_2 fanout134 (.A(net137),
    .X(net134));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(net137));
 sg13g2_buf_2 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_1 fanout137 (.A(net138),
    .X(net137));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(net1));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(net142));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(net141));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(net142));
 sg13g2_buf_2 fanout142 (.A(net146),
    .X(net142));
 sg13g2_buf_4 fanout143 (.X(net143),
    .A(net146));
 sg13g2_buf_2 fanout144 (.A(net146),
    .X(net144));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(net146));
 sg13g2_buf_1 fanout146 (.A(net1),
    .X(net146));
 sg13g2_buf_4 fanout147 (.X(net147),
    .A(net154));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(net154));
 sg13g2_buf_4 fanout149 (.X(net149),
    .A(net154));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(net153));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(net153));
 sg13g2_buf_2 fanout152 (.A(net153),
    .X(net152));
 sg13g2_buf_1 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(net1),
    .X(net154));
 sg13g2_tielo _2998__155 (.L_LO(net155));
 sg13g2_tielo _2999__156 (.L_LO(net156));
 sg13g2_tielo _3000__157 (.L_LO(net157));
 sg13g2_tielo _3002__158 (.L_LO(net158));
 sg13g2_tielo _3003__159 (.L_LO(net159));
 sg13g2_tielo _3004__160 (.L_LO(net160));
 sg13g2_tielo _3006__161 (.L_LO(net161));
 sg13g2_tielo _3007__162 (.L_LO(net162));
 sg13g2_tielo _3008__163 (.L_LO(net163));
 sg13g2_tielo _3009__164 (.L_LO(net164));
 sg13g2_tielo _3010__165 (.L_LO(net165));
 sg13g2_tiehi _2995__167 (.L_HI(net167));
 sg13g2_tiehi _2996__168 (.L_HI(net168));
 sg13g2_tiehi _2997__169 (.L_HI(net169));
 sg13g2_tiehi _3001__170 (.L_HI(net170));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_31__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_fill_2 FILLER_0_63 ();
 sg13g2_fill_1 FILLER_0_65 ();
 sg13g2_fill_2 FILLER_0_76 ();
 sg13g2_fill_1 FILLER_0_78 ();
 sg13g2_fill_2 FILLER_0_92 ();
 sg13g2_fill_1 FILLER_0_94 ();
 sg13g2_decap_8 FILLER_0_104 ();
 sg13g2_decap_8 FILLER_0_111 ();
 sg13g2_decap_8 FILLER_0_118 ();
 sg13g2_decap_8 FILLER_0_125 ();
 sg13g2_decap_8 FILLER_0_132 ();
 sg13g2_decap_8 FILLER_0_139 ();
 sg13g2_decap_8 FILLER_0_146 ();
 sg13g2_decap_4 FILLER_0_153 ();
 sg13g2_fill_2 FILLER_0_157 ();
 sg13g2_decap_4 FILLER_0_172 ();
 sg13g2_fill_1 FILLER_0_176 ();
 sg13g2_decap_4 FILLER_0_182 ();
 sg13g2_fill_1 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_200 ();
 sg13g2_fill_2 FILLER_0_207 ();
 sg13g2_decap_8 FILLER_0_214 ();
 sg13g2_fill_2 FILLER_0_221 ();
 sg13g2_fill_2 FILLER_0_248 ();
 sg13g2_decap_8 FILLER_0_255 ();
 sg13g2_decap_8 FILLER_0_262 ();
 sg13g2_decap_8 FILLER_0_269 ();
 sg13g2_decap_8 FILLER_0_276 ();
 sg13g2_decap_8 FILLER_0_283 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_fill_2 FILLER_0_297 ();
 sg13g2_fill_1 FILLER_0_304 ();
 sg13g2_decap_8 FILLER_0_317 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_decap_4 FILLER_0_331 ();
 sg13g2_fill_2 FILLER_0_335 ();
 sg13g2_decap_4 FILLER_0_341 ();
 sg13g2_fill_2 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_fill_2 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_0_412 ();
 sg13g2_decap_8 FILLER_0_419 ();
 sg13g2_decap_4 FILLER_0_426 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_4 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_46 ();
 sg13g2_fill_2 FILLER_1_64 ();
 sg13g2_fill_1 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_76 ();
 sg13g2_decap_4 FILLER_1_89 ();
 sg13g2_fill_2 FILLER_1_97 ();
 sg13g2_fill_1 FILLER_1_99 ();
 sg13g2_fill_2 FILLER_1_105 ();
 sg13g2_fill_1 FILLER_1_107 ();
 sg13g2_decap_4 FILLER_1_125 ();
 sg13g2_fill_1 FILLER_1_129 ();
 sg13g2_fill_2 FILLER_1_144 ();
 sg13g2_fill_2 FILLER_1_151 ();
 sg13g2_fill_1 FILLER_1_153 ();
 sg13g2_fill_2 FILLER_1_159 ();
 sg13g2_fill_1 FILLER_1_161 ();
 sg13g2_fill_2 FILLER_1_167 ();
 sg13g2_fill_1 FILLER_1_169 ();
 sg13g2_fill_2 FILLER_1_175 ();
 sg13g2_fill_2 FILLER_1_198 ();
 sg13g2_decap_4 FILLER_1_205 ();
 sg13g2_fill_1 FILLER_1_216 ();
 sg13g2_fill_2 FILLER_1_253 ();
 sg13g2_decap_4 FILLER_1_267 ();
 sg13g2_fill_1 FILLER_1_283 ();
 sg13g2_fill_2 FILLER_1_297 ();
 sg13g2_fill_2 FILLER_1_309 ();
 sg13g2_decap_4 FILLER_1_321 ();
 sg13g2_fill_1 FILLER_1_325 ();
 sg13g2_fill_1 FILLER_1_340 ();
 sg13g2_decap_8 FILLER_1_368 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_fill_1 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_decap_8 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_fill_2 FILLER_2_35 ();
 sg13g2_fill_1 FILLER_2_37 ();
 sg13g2_decap_4 FILLER_2_46 ();
 sg13g2_fill_1 FILLER_2_62 ();
 sg13g2_fill_1 FILLER_2_78 ();
 sg13g2_fill_2 FILLER_2_87 ();
 sg13g2_fill_1 FILLER_2_106 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_4 FILLER_2_124 ();
 sg13g2_fill_2 FILLER_2_128 ();
 sg13g2_fill_1 FILLER_2_144 ();
 sg13g2_fill_1 FILLER_2_150 ();
 sg13g2_fill_1 FILLER_2_156 ();
 sg13g2_fill_1 FILLER_2_167 ();
 sg13g2_decap_8 FILLER_2_173 ();
 sg13g2_decap_4 FILLER_2_180 ();
 sg13g2_fill_2 FILLER_2_184 ();
 sg13g2_fill_2 FILLER_2_201 ();
 sg13g2_fill_1 FILLER_2_203 ();
 sg13g2_fill_1 FILLER_2_207 ();
 sg13g2_fill_2 FILLER_2_238 ();
 sg13g2_fill_2 FILLER_2_245 ();
 sg13g2_fill_2 FILLER_2_275 ();
 sg13g2_fill_2 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_295 ();
 sg13g2_decap_4 FILLER_2_302 ();
 sg13g2_fill_1 FILLER_2_326 ();
 sg13g2_fill_2 FILLER_2_332 ();
 sg13g2_decap_8 FILLER_2_339 ();
 sg13g2_fill_2 FILLER_2_346 ();
 sg13g2_fill_1 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_fill_2 FILLER_2_378 ();
 sg13g2_fill_1 FILLER_2_380 ();
 sg13g2_fill_1 FILLER_2_389 ();
 sg13g2_fill_1 FILLER_2_398 ();
 sg13g2_decap_8 FILLER_2_404 ();
 sg13g2_decap_8 FILLER_2_411 ();
 sg13g2_decap_8 FILLER_2_418 ();
 sg13g2_decap_4 FILLER_2_425 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_7 ();
 sg13g2_fill_1 FILLER_3_9 ();
 sg13g2_fill_2 FILLER_3_26 ();
 sg13g2_fill_1 FILLER_3_32 ();
 sg13g2_fill_1 FILLER_3_44 ();
 sg13g2_fill_1 FILLER_3_49 ();
 sg13g2_fill_1 FILLER_3_91 ();
 sg13g2_fill_2 FILLER_3_122 ();
 sg13g2_fill_1 FILLER_3_124 ();
 sg13g2_fill_1 FILLER_3_133 ();
 sg13g2_fill_1 FILLER_3_142 ();
 sg13g2_fill_2 FILLER_3_148 ();
 sg13g2_decap_4 FILLER_3_158 ();
 sg13g2_fill_1 FILLER_3_171 ();
 sg13g2_fill_1 FILLER_3_181 ();
 sg13g2_fill_2 FILLER_3_190 ();
 sg13g2_fill_1 FILLER_3_201 ();
 sg13g2_fill_2 FILLER_3_211 ();
 sg13g2_fill_2 FILLER_3_226 ();
 sg13g2_fill_2 FILLER_3_233 ();
 sg13g2_fill_1 FILLER_3_235 ();
 sg13g2_fill_1 FILLER_3_245 ();
 sg13g2_fill_2 FILLER_3_262 ();
 sg13g2_decap_4 FILLER_3_280 ();
 sg13g2_fill_2 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_fill_2 FILLER_3_298 ();
 sg13g2_fill_1 FILLER_3_300 ();
 sg13g2_decap_8 FILLER_3_313 ();
 sg13g2_fill_2 FILLER_3_320 ();
 sg13g2_fill_1 FILLER_3_322 ();
 sg13g2_fill_1 FILLER_3_328 ();
 sg13g2_decap_4 FILLER_3_337 ();
 sg13g2_fill_1 FILLER_3_346 ();
 sg13g2_fill_1 FILLER_3_366 ();
 sg13g2_fill_1 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_402 ();
 sg13g2_decap_8 FILLER_3_409 ();
 sg13g2_decap_8 FILLER_3_416 ();
 sg13g2_decap_8 FILLER_3_423 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_2 ();
 sg13g2_fill_2 FILLER_4_35 ();
 sg13g2_fill_1 FILLER_4_51 ();
 sg13g2_fill_2 FILLER_4_74 ();
 sg13g2_decap_8 FILLER_4_81 ();
 sg13g2_fill_1 FILLER_4_88 ();
 sg13g2_fill_1 FILLER_4_101 ();
 sg13g2_fill_2 FILLER_4_113 ();
 sg13g2_fill_1 FILLER_4_123 ();
 sg13g2_decap_4 FILLER_4_134 ();
 sg13g2_fill_1 FILLER_4_138 ();
 sg13g2_fill_2 FILLER_4_152 ();
 sg13g2_fill_1 FILLER_4_154 ();
 sg13g2_fill_1 FILLER_4_162 ();
 sg13g2_decap_8 FILLER_4_167 ();
 sg13g2_fill_2 FILLER_4_174 ();
 sg13g2_decap_4 FILLER_4_180 ();
 sg13g2_fill_2 FILLER_4_184 ();
 sg13g2_fill_1 FILLER_4_195 ();
 sg13g2_fill_1 FILLER_4_223 ();
 sg13g2_fill_1 FILLER_4_232 ();
 sg13g2_fill_2 FILLER_4_242 ();
 sg13g2_decap_8 FILLER_4_262 ();
 sg13g2_fill_1 FILLER_4_269 ();
 sg13g2_decap_8 FILLER_4_279 ();
 sg13g2_fill_2 FILLER_4_286 ();
 sg13g2_fill_2 FILLER_4_297 ();
 sg13g2_fill_1 FILLER_4_299 ();
 sg13g2_decap_4 FILLER_4_318 ();
 sg13g2_decap_4 FILLER_4_327 ();
 sg13g2_fill_2 FILLER_4_363 ();
 sg13g2_fill_1 FILLER_4_370 ();
 sg13g2_fill_2 FILLER_4_376 ();
 sg13g2_fill_1 FILLER_4_378 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_fill_1 FILLER_4_409 ();
 sg13g2_fill_1 FILLER_4_415 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_7 ();
 sg13g2_fill_2 FILLER_5_23 ();
 sg13g2_fill_1 FILLER_5_44 ();
 sg13g2_fill_2 FILLER_5_50 ();
 sg13g2_fill_2 FILLER_5_56 ();
 sg13g2_fill_1 FILLER_5_58 ();
 sg13g2_fill_2 FILLER_5_64 ();
 sg13g2_fill_1 FILLER_5_66 ();
 sg13g2_fill_2 FILLER_5_73 ();
 sg13g2_fill_1 FILLER_5_115 ();
 sg13g2_decap_4 FILLER_5_121 ();
 sg13g2_fill_2 FILLER_5_125 ();
 sg13g2_fill_1 FILLER_5_132 ();
 sg13g2_decap_4 FILLER_5_152 ();
 sg13g2_fill_1 FILLER_5_156 ();
 sg13g2_fill_2 FILLER_5_170 ();
 sg13g2_fill_1 FILLER_5_172 ();
 sg13g2_fill_2 FILLER_5_194 ();
 sg13g2_fill_1 FILLER_5_201 ();
 sg13g2_fill_1 FILLER_5_207 ();
 sg13g2_fill_2 FILLER_5_216 ();
 sg13g2_fill_2 FILLER_5_223 ();
 sg13g2_decap_4 FILLER_5_229 ();
 sg13g2_fill_1 FILLER_5_233 ();
 sg13g2_fill_2 FILLER_5_239 ();
 sg13g2_fill_1 FILLER_5_247 ();
 sg13g2_fill_2 FILLER_5_255 ();
 sg13g2_fill_2 FILLER_5_263 ();
 sg13g2_fill_2 FILLER_5_281 ();
 sg13g2_fill_1 FILLER_5_283 ();
 sg13g2_decap_4 FILLER_5_312 ();
 sg13g2_fill_2 FILLER_5_316 ();
 sg13g2_fill_1 FILLER_5_335 ();
 sg13g2_fill_2 FILLER_5_347 ();
 sg13g2_fill_1 FILLER_5_377 ();
 sg13g2_fill_1 FILLER_5_383 ();
 sg13g2_decap_4 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_20 ();
 sg13g2_fill_1 FILLER_6_26 ();
 sg13g2_fill_2 FILLER_6_33 ();
 sg13g2_fill_2 FILLER_6_43 ();
 sg13g2_fill_1 FILLER_6_45 ();
 sg13g2_fill_1 FILLER_6_51 ();
 sg13g2_fill_2 FILLER_6_57 ();
 sg13g2_fill_1 FILLER_6_59 ();
 sg13g2_fill_1 FILLER_6_64 ();
 sg13g2_fill_1 FILLER_6_69 ();
 sg13g2_fill_2 FILLER_6_80 ();
 sg13g2_fill_1 FILLER_6_87 ();
 sg13g2_fill_2 FILLER_6_96 ();
 sg13g2_fill_1 FILLER_6_98 ();
 sg13g2_fill_1 FILLER_6_103 ();
 sg13g2_decap_8 FILLER_6_109 ();
 sg13g2_fill_1 FILLER_6_140 ();
 sg13g2_fill_2 FILLER_6_146 ();
 sg13g2_fill_2 FILLER_6_154 ();
 sg13g2_fill_2 FILLER_6_166 ();
 sg13g2_fill_1 FILLER_6_168 ();
 sg13g2_fill_2 FILLER_6_207 ();
 sg13g2_fill_1 FILLER_6_229 ();
 sg13g2_decap_4 FILLER_6_234 ();
 sg13g2_fill_2 FILLER_6_246 ();
 sg13g2_fill_1 FILLER_6_248 ();
 sg13g2_fill_2 FILLER_6_258 ();
 sg13g2_fill_1 FILLER_6_260 ();
 sg13g2_fill_2 FILLER_6_265 ();
 sg13g2_fill_1 FILLER_6_278 ();
 sg13g2_decap_8 FILLER_6_283 ();
 sg13g2_fill_2 FILLER_6_290 ();
 sg13g2_fill_1 FILLER_6_292 ();
 sg13g2_fill_1 FILLER_6_318 ();
 sg13g2_fill_1 FILLER_6_324 ();
 sg13g2_fill_2 FILLER_6_331 ();
 sg13g2_fill_2 FILLER_6_341 ();
 sg13g2_fill_1 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_348 ();
 sg13g2_fill_2 FILLER_6_371 ();
 sg13g2_fill_1 FILLER_6_373 ();
 sg13g2_fill_1 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_423 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_4 ();
 sg13g2_fill_2 FILLER_7_13 ();
 sg13g2_fill_1 FILLER_7_35 ();
 sg13g2_fill_1 FILLER_7_41 ();
 sg13g2_fill_1 FILLER_7_47 ();
 sg13g2_fill_2 FILLER_7_53 ();
 sg13g2_fill_2 FILLER_7_71 ();
 sg13g2_fill_1 FILLER_7_73 ();
 sg13g2_fill_1 FILLER_7_78 ();
 sg13g2_fill_2 FILLER_7_95 ();
 sg13g2_fill_1 FILLER_7_97 ();
 sg13g2_decap_8 FILLER_7_107 ();
 sg13g2_fill_1 FILLER_7_123 ();
 sg13g2_fill_1 FILLER_7_129 ();
 sg13g2_fill_2 FILLER_7_135 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_fill_2 FILLER_7_147 ();
 sg13g2_fill_1 FILLER_7_149 ();
 sg13g2_fill_1 FILLER_7_162 ();
 sg13g2_decap_4 FILLER_7_177 ();
 sg13g2_fill_1 FILLER_7_181 ();
 sg13g2_decap_4 FILLER_7_186 ();
 sg13g2_fill_2 FILLER_7_201 ();
 sg13g2_fill_2 FILLER_7_235 ();
 sg13g2_fill_1 FILLER_7_237 ();
 sg13g2_decap_4 FILLER_7_246 ();
 sg13g2_fill_2 FILLER_7_250 ();
 sg13g2_fill_2 FILLER_7_256 ();
 sg13g2_decap_4 FILLER_7_262 ();
 sg13g2_fill_2 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_279 ();
 sg13g2_fill_1 FILLER_7_296 ();
 sg13g2_fill_1 FILLER_7_301 ();
 sg13g2_fill_1 FILLER_7_306 ();
 sg13g2_fill_2 FILLER_7_312 ();
 sg13g2_fill_1 FILLER_7_329 ();
 sg13g2_fill_1 FILLER_7_339 ();
 sg13g2_fill_1 FILLER_7_362 ();
 sg13g2_fill_2 FILLER_7_391 ();
 sg13g2_fill_1 FILLER_7_399 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_2 FILLER_7_414 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_decap_4 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_4 ();
 sg13g2_fill_1 FILLER_8_10 ();
 sg13g2_fill_1 FILLER_8_20 ();
 sg13g2_fill_1 FILLER_8_25 ();
 sg13g2_fill_1 FILLER_8_32 ();
 sg13g2_fill_1 FILLER_8_59 ();
 sg13g2_fill_2 FILLER_8_72 ();
 sg13g2_fill_1 FILLER_8_82 ();
 sg13g2_fill_2 FILLER_8_88 ();
 sg13g2_fill_2 FILLER_8_103 ();
 sg13g2_fill_1 FILLER_8_105 ();
 sg13g2_fill_1 FILLER_8_114 ();
 sg13g2_fill_1 FILLER_8_132 ();
 sg13g2_decap_8 FILLER_8_137 ();
 sg13g2_decap_8 FILLER_8_144 ();
 sg13g2_fill_1 FILLER_8_165 ();
 sg13g2_fill_2 FILLER_8_197 ();
 sg13g2_fill_2 FILLER_8_203 ();
 sg13g2_fill_2 FILLER_8_215 ();
 sg13g2_fill_2 FILLER_8_221 ();
 sg13g2_fill_2 FILLER_8_227 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_fill_2 FILLER_8_260 ();
 sg13g2_fill_2 FILLER_8_266 ();
 sg13g2_fill_1 FILLER_8_268 ();
 sg13g2_fill_2 FILLER_8_282 ();
 sg13g2_fill_2 FILLER_8_289 ();
 sg13g2_fill_2 FILLER_8_316 ();
 sg13g2_fill_1 FILLER_8_318 ();
 sg13g2_decap_4 FILLER_8_329 ();
 sg13g2_fill_2 FILLER_8_333 ();
 sg13g2_fill_1 FILLER_8_346 ();
 sg13g2_fill_1 FILLER_8_357 ();
 sg13g2_fill_1 FILLER_8_373 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_4 FILLER_8_412 ();
 sg13g2_fill_2 FILLER_8_416 ();
 sg13g2_decap_8 FILLER_8_423 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_7 ();
 sg13g2_decap_4 FILLER_9_40 ();
 sg13g2_fill_2 FILLER_9_48 ();
 sg13g2_fill_1 FILLER_9_55 ();
 sg13g2_fill_2 FILLER_9_61 ();
 sg13g2_fill_1 FILLER_9_68 ();
 sg13g2_fill_1 FILLER_9_79 ();
 sg13g2_fill_2 FILLER_9_85 ();
 sg13g2_fill_1 FILLER_9_100 ();
 sg13g2_decap_8 FILLER_9_124 ();
 sg13g2_decap_8 FILLER_9_131 ();
 sg13g2_fill_2 FILLER_9_138 ();
 sg13g2_fill_1 FILLER_9_140 ();
 sg13g2_fill_2 FILLER_9_165 ();
 sg13g2_fill_1 FILLER_9_173 ();
 sg13g2_fill_2 FILLER_9_182 ();
 sg13g2_fill_1 FILLER_9_184 ();
 sg13g2_decap_8 FILLER_9_211 ();
 sg13g2_fill_1 FILLER_9_218 ();
 sg13g2_fill_2 FILLER_9_242 ();
 sg13g2_fill_1 FILLER_9_244 ();
 sg13g2_fill_2 FILLER_9_275 ();
 sg13g2_decap_4 FILLER_9_282 ();
 sg13g2_fill_2 FILLER_9_328 ();
 sg13g2_fill_1 FILLER_9_330 ();
 sg13g2_decap_8 FILLER_9_341 ();
 sg13g2_decap_4 FILLER_9_369 ();
 sg13g2_fill_1 FILLER_9_383 ();
 sg13g2_decap_4 FILLER_9_394 ();
 sg13g2_fill_2 FILLER_9_398 ();
 sg13g2_decap_8 FILLER_9_418 ();
 sg13g2_decap_4 FILLER_9_425 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_11 ();
 sg13g2_fill_1 FILLER_10_33 ();
 sg13g2_fill_2 FILLER_10_44 ();
 sg13g2_fill_1 FILLER_10_96 ();
 sg13g2_fill_1 FILLER_10_100 ();
 sg13g2_fill_1 FILLER_10_105 ();
 sg13g2_decap_4 FILLER_10_120 ();
 sg13g2_decap_4 FILLER_10_134 ();
 sg13g2_fill_2 FILLER_10_167 ();
 sg13g2_fill_2 FILLER_10_187 ();
 sg13g2_decap_8 FILLER_10_213 ();
 sg13g2_fill_1 FILLER_10_238 ();
 sg13g2_fill_1 FILLER_10_244 ();
 sg13g2_decap_4 FILLER_10_255 ();
 sg13g2_fill_1 FILLER_10_264 ();
 sg13g2_decap_4 FILLER_10_275 ();
 sg13g2_fill_1 FILLER_10_300 ();
 sg13g2_fill_1 FILLER_10_319 ();
 sg13g2_fill_1 FILLER_10_333 ();
 sg13g2_fill_1 FILLER_10_375 ();
 sg13g2_decap_4 FILLER_10_389 ();
 sg13g2_fill_1 FILLER_10_400 ();
 sg13g2_decap_8 FILLER_10_422 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_4 FILLER_11_31 ();
 sg13g2_fill_2 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_46 ();
 sg13g2_fill_1 FILLER_11_62 ();
 sg13g2_fill_1 FILLER_11_72 ();
 sg13g2_fill_1 FILLER_11_81 ();
 sg13g2_fill_2 FILLER_11_97 ();
 sg13g2_fill_1 FILLER_11_99 ();
 sg13g2_fill_2 FILLER_11_106 ();
 sg13g2_fill_1 FILLER_11_114 ();
 sg13g2_fill_2 FILLER_11_124 ();
 sg13g2_fill_2 FILLER_11_150 ();
 sg13g2_fill_1 FILLER_11_158 ();
 sg13g2_fill_1 FILLER_11_163 ();
 sg13g2_fill_1 FILLER_11_169 ();
 sg13g2_fill_1 FILLER_11_175 ();
 sg13g2_decap_4 FILLER_11_180 ();
 sg13g2_fill_2 FILLER_11_184 ();
 sg13g2_fill_1 FILLER_11_190 ();
 sg13g2_decap_8 FILLER_11_225 ();
 sg13g2_fill_1 FILLER_11_240 ();
 sg13g2_fill_1 FILLER_11_266 ();
 sg13g2_fill_2 FILLER_11_276 ();
 sg13g2_fill_1 FILLER_11_278 ();
 sg13g2_fill_1 FILLER_11_290 ();
 sg13g2_fill_1 FILLER_11_295 ();
 sg13g2_fill_1 FILLER_11_301 ();
 sg13g2_decap_4 FILLER_11_311 ();
 sg13g2_fill_2 FILLER_11_315 ();
 sg13g2_fill_1 FILLER_11_325 ();
 sg13g2_fill_1 FILLER_11_331 ();
 sg13g2_fill_1 FILLER_11_337 ();
 sg13g2_fill_2 FILLER_11_348 ();
 sg13g2_decap_4 FILLER_11_357 ();
 sg13g2_fill_1 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_369 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_decap_4 FILLER_11_383 ();
 sg13g2_fill_1 FILLER_11_387 ();
 sg13g2_decap_4 FILLER_11_424 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_59 ();
 sg13g2_decap_4 FILLER_12_67 ();
 sg13g2_fill_2 FILLER_12_71 ();
 sg13g2_fill_1 FILLER_12_77 ();
 sg13g2_fill_2 FILLER_12_81 ();
 sg13g2_fill_1 FILLER_12_88 ();
 sg13g2_fill_2 FILLER_12_93 ();
 sg13g2_decap_8 FILLER_12_103 ();
 sg13g2_fill_1 FILLER_12_110 ();
 sg13g2_fill_2 FILLER_12_121 ();
 sg13g2_fill_1 FILLER_12_123 ();
 sg13g2_fill_1 FILLER_12_128 ();
 sg13g2_fill_2 FILLER_12_134 ();
 sg13g2_fill_2 FILLER_12_140 ();
 sg13g2_fill_1 FILLER_12_146 ();
 sg13g2_fill_2 FILLER_12_151 ();
 sg13g2_fill_1 FILLER_12_158 ();
 sg13g2_decap_4 FILLER_12_169 ();
 sg13g2_fill_1 FILLER_12_177 ();
 sg13g2_fill_2 FILLER_12_186 ();
 sg13g2_fill_1 FILLER_12_188 ();
 sg13g2_decap_8 FILLER_12_200 ();
 sg13g2_fill_2 FILLER_12_207 ();
 sg13g2_fill_1 FILLER_12_209 ();
 sg13g2_fill_2 FILLER_12_233 ();
 sg13g2_fill_2 FILLER_12_249 ();
 sg13g2_decap_4 FILLER_12_268 ();
 sg13g2_fill_2 FILLER_12_277 ();
 sg13g2_decap_4 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_292 ();
 sg13g2_decap_4 FILLER_12_299 ();
 sg13g2_fill_1 FILLER_12_303 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_4 FILLER_12_322 ();
 sg13g2_fill_1 FILLER_12_344 ();
 sg13g2_decap_4 FILLER_12_350 ();
 sg13g2_fill_2 FILLER_12_354 ();
 sg13g2_fill_2 FILLER_12_360 ();
 sg13g2_fill_2 FILLER_12_404 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_2 ();
 sg13g2_decap_4 FILLER_13_39 ();
 sg13g2_fill_1 FILLER_13_43 ();
 sg13g2_decap_8 FILLER_13_48 ();
 sg13g2_decap_4 FILLER_13_55 ();
 sg13g2_fill_1 FILLER_13_64 ();
 sg13g2_fill_1 FILLER_13_110 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_fill_2 FILLER_13_131 ();
 sg13g2_fill_2 FILLER_13_138 ();
 sg13g2_fill_1 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_13_164 ();
 sg13g2_fill_1 FILLER_13_170 ();
 sg13g2_decap_4 FILLER_13_176 ();
 sg13g2_fill_1 FILLER_13_192 ();
 sg13g2_decap_4 FILLER_13_198 ();
 sg13g2_fill_2 FILLER_13_211 ();
 sg13g2_fill_1 FILLER_13_213 ();
 sg13g2_fill_2 FILLER_13_224 ();
 sg13g2_decap_4 FILLER_13_231 ();
 sg13g2_fill_1 FILLER_13_245 ();
 sg13g2_fill_2 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_260 ();
 sg13g2_fill_2 FILLER_13_276 ();
 sg13g2_decap_8 FILLER_13_288 ();
 sg13g2_fill_2 FILLER_13_295 ();
 sg13g2_fill_2 FILLER_13_303 ();
 sg13g2_decap_8 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_324 ();
 sg13g2_fill_2 FILLER_13_331 ();
 sg13g2_fill_1 FILLER_13_336 ();
 sg13g2_fill_1 FILLER_13_342 ();
 sg13g2_fill_1 FILLER_13_347 ();
 sg13g2_fill_2 FILLER_13_361 ();
 sg13g2_decap_4 FILLER_13_386 ();
 sg13g2_fill_2 FILLER_13_408 ();
 sg13g2_fill_1 FILLER_13_410 ();
 sg13g2_decap_8 FILLER_13_421 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_fill_2 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_30 ();
 sg13g2_decap_8 FILLER_14_57 ();
 sg13g2_fill_1 FILLER_14_90 ();
 sg13g2_decap_4 FILLER_14_107 ();
 sg13g2_decap_8 FILLER_14_131 ();
 sg13g2_fill_2 FILLER_14_148 ();
 sg13g2_fill_1 FILLER_14_150 ();
 sg13g2_fill_1 FILLER_14_165 ();
 sg13g2_fill_1 FILLER_14_191 ();
 sg13g2_fill_1 FILLER_14_211 ();
 sg13g2_decap_4 FILLER_14_217 ();
 sg13g2_fill_1 FILLER_14_221 ();
 sg13g2_fill_2 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_236 ();
 sg13g2_fill_2 FILLER_14_243 ();
 sg13g2_fill_1 FILLER_14_250 ();
 sg13g2_fill_2 FILLER_14_302 ();
 sg13g2_fill_1 FILLER_14_304 ();
 sg13g2_fill_1 FILLER_14_310 ();
 sg13g2_fill_2 FILLER_14_346 ();
 sg13g2_fill_2 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_decap_8 FILLER_14_374 ();
 sg13g2_decap_4 FILLER_14_381 ();
 sg13g2_fill_2 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_416 ();
 sg13g2_decap_8 FILLER_14_423 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_9 ();
 sg13g2_decap_8 FILLER_15_20 ();
 sg13g2_fill_2 FILLER_15_27 ();
 sg13g2_fill_1 FILLER_15_29 ();
 sg13g2_decap_8 FILLER_15_34 ();
 sg13g2_decap_8 FILLER_15_41 ();
 sg13g2_fill_1 FILLER_15_48 ();
 sg13g2_decap_8 FILLER_15_54 ();
 sg13g2_decap_4 FILLER_15_61 ();
 sg13g2_fill_2 FILLER_15_65 ();
 sg13g2_fill_1 FILLER_15_106 ();
 sg13g2_fill_1 FILLER_15_110 ();
 sg13g2_fill_1 FILLER_15_121 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_4 FILLER_15_133 ();
 sg13g2_fill_2 FILLER_15_137 ();
 sg13g2_fill_1 FILLER_15_150 ();
 sg13g2_fill_1 FILLER_15_161 ();
 sg13g2_fill_2 FILLER_15_167 ();
 sg13g2_fill_1 FILLER_15_169 ();
 sg13g2_fill_2 FILLER_15_178 ();
 sg13g2_decap_4 FILLER_15_185 ();
 sg13g2_decap_8 FILLER_15_197 ();
 sg13g2_decap_4 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_281 ();
 sg13g2_fill_2 FILLER_15_290 ();
 sg13g2_fill_1 FILLER_15_292 ();
 sg13g2_fill_1 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_321 ();
 sg13g2_fill_1 FILLER_15_328 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_4 FILLER_15_367 ();
 sg13g2_fill_2 FILLER_15_371 ();
 sg13g2_fill_1 FILLER_15_400 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_decap_4 FILLER_15_426 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_15 ();
 sg13g2_fill_1 FILLER_16_22 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_82 ();
 sg13g2_decap_8 FILLER_16_89 ();
 sg13g2_decap_8 FILLER_16_96 ();
 sg13g2_decap_4 FILLER_16_108 ();
 sg13g2_fill_2 FILLER_16_132 ();
 sg13g2_fill_1 FILLER_16_139 ();
 sg13g2_fill_1 FILLER_16_145 ();
 sg13g2_fill_2 FILLER_16_151 ();
 sg13g2_fill_1 FILLER_16_169 ();
 sg13g2_fill_2 FILLER_16_184 ();
 sg13g2_fill_2 FILLER_16_194 ();
 sg13g2_decap_4 FILLER_16_201 ();
 sg13g2_decap_4 FILLER_16_213 ();
 sg13g2_decap_4 FILLER_16_224 ();
 sg13g2_fill_2 FILLER_16_240 ();
 sg13g2_fill_1 FILLER_16_267 ();
 sg13g2_fill_1 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_fill_1 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_315 ();
 sg13g2_fill_1 FILLER_16_317 ();
 sg13g2_decap_4 FILLER_16_349 ();
 sg13g2_decap_4 FILLER_16_367 ();
 sg13g2_fill_1 FILLER_16_371 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_1 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_16_421 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_28 ();
 sg13g2_fill_2 FILLER_17_66 ();
 sg13g2_fill_1 FILLER_17_68 ();
 sg13g2_decap_4 FILLER_17_73 ();
 sg13g2_fill_2 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_94 ();
 sg13g2_fill_2 FILLER_17_101 ();
 sg13g2_fill_1 FILLER_17_108 ();
 sg13g2_decap_4 FILLER_17_113 ();
 sg13g2_fill_2 FILLER_17_122 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_142 ();
 sg13g2_fill_2 FILLER_17_151 ();
 sg13g2_fill_1 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_204 ();
 sg13g2_decap_8 FILLER_17_211 ();
 sg13g2_decap_4 FILLER_17_218 ();
 sg13g2_fill_2 FILLER_17_222 ();
 sg13g2_decap_4 FILLER_17_261 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_4 FILLER_17_287 ();
 sg13g2_fill_1 FILLER_17_291 ();
 sg13g2_fill_2 FILLER_17_301 ();
 sg13g2_fill_1 FILLER_17_303 ();
 sg13g2_fill_1 FILLER_17_311 ();
 sg13g2_fill_1 FILLER_17_322 ();
 sg13g2_fill_2 FILLER_17_359 ();
 sg13g2_fill_2 FILLER_17_365 ();
 sg13g2_fill_1 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_fill_2 FILLER_18_12 ();
 sg13g2_fill_1 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_29 ();
 sg13g2_fill_1 FILLER_18_31 ();
 sg13g2_fill_2 FILLER_18_36 ();
 sg13g2_fill_2 FILLER_18_151 ();
 sg13g2_fill_2 FILLER_18_156 ();
 sg13g2_decap_8 FILLER_18_176 ();
 sg13g2_decap_8 FILLER_18_183 ();
 sg13g2_decap_8 FILLER_18_190 ();
 sg13g2_decap_8 FILLER_18_197 ();
 sg13g2_fill_2 FILLER_18_204 ();
 sg13g2_fill_1 FILLER_18_206 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_222 ();
 sg13g2_fill_2 FILLER_18_229 ();
 sg13g2_decap_4 FILLER_18_245 ();
 sg13g2_fill_2 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_255 ();
 sg13g2_fill_1 FILLER_18_262 ();
 sg13g2_fill_2 FILLER_18_267 ();
 sg13g2_fill_1 FILLER_18_273 ();
 sg13g2_fill_2 FILLER_18_288 ();
 sg13g2_fill_1 FILLER_18_290 ();
 sg13g2_fill_2 FILLER_18_306 ();
 sg13g2_fill_1 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_321 ();
 sg13g2_fill_1 FILLER_18_328 ();
 sg13g2_fill_2 FILLER_18_337 ();
 sg13g2_fill_1 FILLER_18_353 ();
 sg13g2_fill_1 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_417 ();
 sg13g2_decap_4 FILLER_18_424 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_decap_4 FILLER_19_55 ();
 sg13g2_decap_8 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_74 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_83 ();
 sg13g2_decap_4 FILLER_19_88 ();
 sg13g2_fill_2 FILLER_19_92 ();
 sg13g2_decap_8 FILLER_19_115 ();
 sg13g2_decap_4 FILLER_19_122 ();
 sg13g2_fill_1 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_144 ();
 sg13g2_fill_1 FILLER_19_151 ();
 sg13g2_decap_8 FILLER_19_156 ();
 sg13g2_decap_4 FILLER_19_163 ();
 sg13g2_fill_2 FILLER_19_186 ();
 sg13g2_fill_2 FILLER_19_198 ();
 sg13g2_fill_1 FILLER_19_200 ();
 sg13g2_fill_2 FILLER_19_227 ();
 sg13g2_fill_1 FILLER_19_229 ();
 sg13g2_fill_2 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_236 ();
 sg13g2_fill_2 FILLER_19_241 ();
 sg13g2_fill_2 FILLER_19_256 ();
 sg13g2_fill_1 FILLER_19_264 ();
 sg13g2_fill_2 FILLER_19_275 ();
 sg13g2_fill_2 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_304 ();
 sg13g2_fill_1 FILLER_19_310 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_322 ();
 sg13g2_fill_2 FILLER_19_337 ();
 sg13g2_decap_4 FILLER_19_342 ();
 sg13g2_fill_1 FILLER_19_362 ();
 sg13g2_fill_2 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_8 FILLER_19_403 ();
 sg13g2_decap_8 FILLER_19_410 ();
 sg13g2_decap_8 FILLER_19_417 ();
 sg13g2_decap_4 FILLER_19_424 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_4 FILLER_20_28 ();
 sg13g2_decap_4 FILLER_20_58 ();
 sg13g2_decap_4 FILLER_20_98 ();
 sg13g2_fill_2 FILLER_20_102 ();
 sg13g2_decap_4 FILLER_20_108 ();
 sg13g2_fill_2 FILLER_20_112 ();
 sg13g2_fill_1 FILLER_20_124 ();
 sg13g2_fill_2 FILLER_20_134 ();
 sg13g2_fill_1 FILLER_20_136 ();
 sg13g2_fill_2 FILLER_20_163 ();
 sg13g2_fill_1 FILLER_20_165 ();
 sg13g2_fill_1 FILLER_20_192 ();
 sg13g2_fill_1 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_203 ();
 sg13g2_fill_1 FILLER_20_217 ();
 sg13g2_fill_1 FILLER_20_221 ();
 sg13g2_fill_2 FILLER_20_248 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_fill_1 FILLER_20_276 ();
 sg13g2_fill_1 FILLER_20_281 ();
 sg13g2_fill_2 FILLER_20_290 ();
 sg13g2_fill_2 FILLER_20_297 ();
 sg13g2_decap_4 FILLER_20_303 ();
 sg13g2_fill_2 FILLER_20_315 ();
 sg13g2_fill_1 FILLER_20_317 ();
 sg13g2_fill_1 FILLER_20_322 ();
 sg13g2_fill_1 FILLER_20_331 ();
 sg13g2_fill_1 FILLER_20_337 ();
 sg13g2_fill_1 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_decap_4 FILLER_20_393 ();
 sg13g2_fill_1 FILLER_20_397 ();
 sg13g2_decap_8 FILLER_20_416 ();
 sg13g2_decap_8 FILLER_20_423 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_decap_4 FILLER_21_44 ();
 sg13g2_fill_2 FILLER_21_48 ();
 sg13g2_fill_2 FILLER_21_60 ();
 sg13g2_decap_4 FILLER_21_102 ();
 sg13g2_fill_1 FILLER_21_106 ();
 sg13g2_fill_1 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_138 ();
 sg13g2_fill_1 FILLER_21_156 ();
 sg13g2_decap_8 FILLER_21_160 ();
 sg13g2_decap_8 FILLER_21_167 ();
 sg13g2_decap_4 FILLER_21_174 ();
 sg13g2_fill_1 FILLER_21_178 ();
 sg13g2_decap_4 FILLER_21_192 ();
 sg13g2_fill_1 FILLER_21_196 ();
 sg13g2_decap_4 FILLER_21_228 ();
 sg13g2_fill_2 FILLER_21_232 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_decap_4 FILLER_21_257 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_decap_8 FILLER_21_275 ();
 sg13g2_decap_8 FILLER_21_282 ();
 sg13g2_fill_2 FILLER_21_289 ();
 sg13g2_decap_8 FILLER_21_299 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_fill_2 FILLER_21_313 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_fill_2 FILLER_21_330 ();
 sg13g2_fill_2 FILLER_21_337 ();
 sg13g2_fill_1 FILLER_21_339 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_4 FILLER_21_382 ();
 sg13g2_fill_1 FILLER_21_386 ();
 sg13g2_fill_2 FILLER_21_392 ();
 sg13g2_fill_1 FILLER_21_394 ();
 sg13g2_fill_1 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_404 ();
 sg13g2_decap_8 FILLER_21_411 ();
 sg13g2_decap_8 FILLER_21_418 ();
 sg13g2_decap_4 FILLER_21_425 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_33 ();
 sg13g2_decap_8 FILLER_22_40 ();
 sg13g2_fill_2 FILLER_22_47 ();
 sg13g2_fill_1 FILLER_22_49 ();
 sg13g2_fill_2 FILLER_22_68 ();
 sg13g2_fill_1 FILLER_22_70 ();
 sg13g2_fill_2 FILLER_22_81 ();
 sg13g2_decap_8 FILLER_22_92 ();
 sg13g2_decap_8 FILLER_22_99 ();
 sg13g2_fill_2 FILLER_22_115 ();
 sg13g2_fill_1 FILLER_22_122 ();
 sg13g2_fill_1 FILLER_22_127 ();
 sg13g2_fill_2 FILLER_22_132 ();
 sg13g2_fill_2 FILLER_22_158 ();
 sg13g2_fill_1 FILLER_22_160 ();
 sg13g2_fill_2 FILLER_22_195 ();
 sg13g2_fill_1 FILLER_22_197 ();
 sg13g2_decap_4 FILLER_22_206 ();
 sg13g2_decap_4 FILLER_22_214 ();
 sg13g2_fill_1 FILLER_22_218 ();
 sg13g2_decap_4 FILLER_22_224 ();
 sg13g2_fill_2 FILLER_22_228 ();
 sg13g2_fill_2 FILLER_22_234 ();
 sg13g2_fill_1 FILLER_22_252 ();
 sg13g2_decap_4 FILLER_22_257 ();
 sg13g2_fill_2 FILLER_22_266 ();
 sg13g2_fill_1 FILLER_22_273 ();
 sg13g2_fill_2 FILLER_22_280 ();
 sg13g2_fill_1 FILLER_22_296 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_fill_2 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_4 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_360 ();
 sg13g2_decap_4 FILLER_22_367 ();
 sg13g2_fill_1 FILLER_22_389 ();
 sg13g2_fill_2 FILLER_22_394 ();
 sg13g2_fill_2 FILLER_22_401 ();
 sg13g2_decap_4 FILLER_22_408 ();
 sg13g2_fill_1 FILLER_22_412 ();
 sg13g2_decap_4 FILLER_22_426 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_4 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_18 ();
 sg13g2_fill_1 FILLER_23_131 ();
 sg13g2_fill_1 FILLER_23_136 ();
 sg13g2_decap_8 FILLER_23_149 ();
 sg13g2_fill_1 FILLER_23_156 ();
 sg13g2_fill_1 FILLER_23_208 ();
 sg13g2_fill_2 FILLER_23_214 ();
 sg13g2_fill_2 FILLER_23_226 ();
 sg13g2_fill_1 FILLER_23_228 ();
 sg13g2_decap_4 FILLER_23_239 ();
 sg13g2_fill_1 FILLER_23_243 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_fill_2 FILLER_23_265 ();
 sg13g2_fill_2 FILLER_23_293 ();
 sg13g2_fill_1 FILLER_23_330 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_fill_2 FILLER_23_365 ();
 sg13g2_fill_1 FILLER_23_372 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_fill_1 FILLER_23_388 ();
 sg13g2_decap_4 FILLER_23_399 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_45 ();
 sg13g2_fill_2 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_92 ();
 sg13g2_fill_1 FILLER_24_97 ();
 sg13g2_fill_2 FILLER_24_104 ();
 sg13g2_fill_2 FILLER_24_114 ();
 sg13g2_fill_2 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_122 ();
 sg13g2_decap_8 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_144 ();
 sg13g2_fill_1 FILLER_24_158 ();
 sg13g2_decap_4 FILLER_24_183 ();
 sg13g2_decap_8 FILLER_24_206 ();
 sg13g2_decap_4 FILLER_24_213 ();
 sg13g2_fill_2 FILLER_24_260 ();
 sg13g2_fill_1 FILLER_24_262 ();
 sg13g2_decap_8 FILLER_24_312 ();
 sg13g2_fill_1 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_326 ();
 sg13g2_decap_4 FILLER_24_333 ();
 sg13g2_decap_8 FILLER_24_351 ();
 sg13g2_fill_2 FILLER_24_368 ();
 sg13g2_fill_2 FILLER_24_375 ();
 sg13g2_fill_1 FILLER_24_377 ();
 sg13g2_fill_1 FILLER_24_383 ();
 sg13g2_fill_2 FILLER_24_388 ();
 sg13g2_fill_1 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_422 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_9 ();
 sg13g2_fill_2 FILLER_25_20 ();
 sg13g2_decap_8 FILLER_25_36 ();
 sg13g2_decap_8 FILLER_25_43 ();
 sg13g2_decap_8 FILLER_25_50 ();
 sg13g2_decap_4 FILLER_25_57 ();
 sg13g2_fill_1 FILLER_25_72 ();
 sg13g2_fill_1 FILLER_25_78 ();
 sg13g2_fill_1 FILLER_25_89 ();
 sg13g2_fill_1 FILLER_25_106 ();
 sg13g2_fill_2 FILLER_25_120 ();
 sg13g2_fill_1 FILLER_25_122 ();
 sg13g2_decap_4 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_159 ();
 sg13g2_fill_1 FILLER_25_174 ();
 sg13g2_fill_1 FILLER_25_185 ();
 sg13g2_fill_2 FILLER_25_190 ();
 sg13g2_decap_4 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_200 ();
 sg13g2_decap_4 FILLER_25_220 ();
 sg13g2_fill_2 FILLER_25_224 ();
 sg13g2_fill_2 FILLER_25_236 ();
 sg13g2_fill_1 FILLER_25_238 ();
 sg13g2_fill_2 FILLER_25_255 ();
 sg13g2_fill_1 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_282 ();
 sg13g2_fill_1 FILLER_25_286 ();
 sg13g2_fill_1 FILLER_25_291 ();
 sg13g2_fill_2 FILLER_25_305 ();
 sg13g2_fill_1 FILLER_25_338 ();
 sg13g2_decap_4 FILLER_25_382 ();
 sg13g2_fill_2 FILLER_25_386 ();
 sg13g2_fill_2 FILLER_25_392 ();
 sg13g2_fill_1 FILLER_25_394 ();
 sg13g2_fill_1 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_4 FILLER_25_424 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_39 ();
 sg13g2_fill_1 FILLER_26_50 ();
 sg13g2_fill_1 FILLER_26_87 ();
 sg13g2_fill_1 FILLER_26_92 ();
 sg13g2_fill_2 FILLER_26_119 ();
 sg13g2_decap_4 FILLER_26_136 ();
 sg13g2_fill_2 FILLER_26_140 ();
 sg13g2_decap_4 FILLER_26_147 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_fill_2 FILLER_26_213 ();
 sg13g2_fill_1 FILLER_26_215 ();
 sg13g2_decap_8 FILLER_26_225 ();
 sg13g2_decap_4 FILLER_26_232 ();
 sg13g2_fill_1 FILLER_26_236 ();
 sg13g2_decap_4 FILLER_26_242 ();
 sg13g2_fill_1 FILLER_26_246 ();
 sg13g2_fill_1 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_290 ();
 sg13g2_fill_2 FILLER_26_310 ();
 sg13g2_fill_1 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_341 ();
 sg13g2_fill_1 FILLER_26_352 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_fill_1 FILLER_26_363 ();
 sg13g2_fill_1 FILLER_26_369 ();
 sg13g2_fill_1 FILLER_26_375 ();
 sg13g2_fill_1 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_26_412 ();
 sg13g2_decap_8 FILLER_26_419 ();
 sg13g2_decap_4 FILLER_26_426 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_37 ();
 sg13g2_fill_2 FILLER_27_44 ();
 sg13g2_decap_4 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_86 ();
 sg13g2_decap_4 FILLER_27_156 ();
 sg13g2_decap_8 FILLER_27_174 ();
 sg13g2_decap_4 FILLER_27_181 ();
 sg13g2_fill_1 FILLER_27_185 ();
 sg13g2_fill_2 FILLER_27_190 ();
 sg13g2_decap_4 FILLER_27_202 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_4 FILLER_27_224 ();
 sg13g2_fill_2 FILLER_27_228 ();
 sg13g2_fill_2 FILLER_27_240 ();
 sg13g2_fill_1 FILLER_27_247 ();
 sg13g2_fill_2 FILLER_27_253 ();
 sg13g2_fill_1 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_271 ();
 sg13g2_fill_2 FILLER_27_277 ();
 sg13g2_decap_4 FILLER_27_294 ();
 sg13g2_fill_2 FILLER_27_306 ();
 sg13g2_fill_1 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_318 ();
 sg13g2_fill_2 FILLER_27_325 ();
 sg13g2_fill_2 FILLER_27_335 ();
 sg13g2_fill_2 FILLER_27_354 ();
 sg13g2_fill_1 FILLER_27_356 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_fill_1 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_11 ();
 sg13g2_decap_4 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_53 ();
 sg13g2_decap_4 FILLER_28_59 ();
 sg13g2_fill_2 FILLER_28_63 ();
 sg13g2_fill_1 FILLER_28_109 ();
 sg13g2_fill_2 FILLER_28_136 ();
 sg13g2_fill_1 FILLER_28_138 ();
 sg13g2_fill_2 FILLER_28_143 ();
 sg13g2_fill_2 FILLER_28_151 ();
 sg13g2_fill_2 FILLER_28_157 ();
 sg13g2_fill_1 FILLER_28_159 ();
 sg13g2_fill_1 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_233 ();
 sg13g2_decap_8 FILLER_28_240 ();
 sg13g2_fill_1 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_decap_8 FILLER_28_330 ();
 sg13g2_decap_8 FILLER_28_337 ();
 sg13g2_decap_4 FILLER_28_344 ();
 sg13g2_fill_2 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_32 ();
 sg13g2_fill_2 FILLER_29_79 ();
 sg13g2_decap_4 FILLER_29_85 ();
 sg13g2_decap_4 FILLER_29_94 ();
 sg13g2_fill_2 FILLER_29_98 ();
 sg13g2_decap_4 FILLER_29_109 ();
 sg13g2_fill_1 FILLER_29_113 ();
 sg13g2_decap_4 FILLER_29_117 ();
 sg13g2_fill_2 FILLER_29_121 ();
 sg13g2_decap_4 FILLER_29_128 ();
 sg13g2_fill_2 FILLER_29_132 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_decap_8 FILLER_29_163 ();
 sg13g2_decap_8 FILLER_29_170 ();
 sg13g2_decap_4 FILLER_29_177 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_fill_2 FILLER_29_196 ();
 sg13g2_fill_1 FILLER_29_198 ();
 sg13g2_fill_2 FILLER_29_235 ();
 sg13g2_fill_1 FILLER_29_237 ();
 sg13g2_fill_1 FILLER_29_273 ();
 sg13g2_decap_4 FILLER_29_287 ();
 sg13g2_fill_1 FILLER_29_291 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_fill_2 FILLER_29_304 ();
 sg13g2_fill_1 FILLER_29_306 ();
 sg13g2_fill_2 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_313 ();
 sg13g2_fill_2 FILLER_29_318 ();
 sg13g2_decap_4 FILLER_29_351 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_8 FILLER_29_403 ();
 sg13g2_decap_8 FILLER_29_410 ();
 sg13g2_decap_8 FILLER_29_417 ();
 sg13g2_decap_4 FILLER_29_424 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_2 FILLER_30_39 ();
 sg13g2_fill_1 FILLER_30_41 ();
 sg13g2_fill_1 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_116 ();
 sg13g2_fill_1 FILLER_30_118 ();
 sg13g2_decap_8 FILLER_30_145 ();
 sg13g2_fill_2 FILLER_30_152 ();
 sg13g2_fill_1 FILLER_30_154 ();
 sg13g2_decap_4 FILLER_30_194 ();
 sg13g2_fill_2 FILLER_30_198 ();
 sg13g2_decap_8 FILLER_30_236 ();
 sg13g2_fill_1 FILLER_30_243 ();
 sg13g2_decap_8 FILLER_30_251 ();
 sg13g2_decap_8 FILLER_30_258 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_fill_2 FILLER_30_297 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_4 FILLER_30_364 ();
 sg13g2_fill_2 FILLER_30_368 ();
 sg13g2_fill_2 FILLER_30_374 ();
 sg13g2_fill_1 FILLER_30_376 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_30_417 ();
 sg13g2_decap_4 FILLER_30_424 ();
 sg13g2_fill_2 FILLER_30_428 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_decap_4 FILLER_31_51 ();
 sg13g2_fill_2 FILLER_31_89 ();
 sg13g2_decap_8 FILLER_31_103 ();
 sg13g2_decap_8 FILLER_31_160 ();
 sg13g2_decap_4 FILLER_31_167 ();
 sg13g2_decap_8 FILLER_31_207 ();
 sg13g2_fill_2 FILLER_31_214 ();
 sg13g2_fill_2 FILLER_31_221 ();
 sg13g2_fill_1 FILLER_31_223 ();
 sg13g2_fill_2 FILLER_31_228 ();
 sg13g2_fill_1 FILLER_31_230 ();
 sg13g2_decap_4 FILLER_31_235 ();
 sg13g2_fill_2 FILLER_31_239 ();
 sg13g2_decap_4 FILLER_31_267 ();
 sg13g2_fill_2 FILLER_31_271 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_fill_2 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_341 ();
 sg13g2_fill_1 FILLER_31_384 ();
 sg13g2_fill_2 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_423 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_16 ();
 sg13g2_fill_1 FILLER_32_22 ();
 sg13g2_decap_4 FILLER_32_59 ();
 sg13g2_fill_2 FILLER_32_78 ();
 sg13g2_fill_1 FILLER_32_80 ();
 sg13g2_decap_4 FILLER_32_107 ();
 sg13g2_fill_2 FILLER_32_137 ();
 sg13g2_decap_4 FILLER_32_143 ();
 sg13g2_decap_4 FILLER_32_152 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_decap_4 FILLER_32_207 ();
 sg13g2_decap_4 FILLER_32_240 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_decap_8 FILLER_32_271 ();
 sg13g2_decap_8 FILLER_32_282 ();
 sg13g2_fill_2 FILLER_32_289 ();
 sg13g2_fill_1 FILLER_32_291 ();
 sg13g2_decap_4 FILLER_32_299 ();
 sg13g2_decap_4 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_368 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_72 ();
 sg13g2_decap_8 FILLER_33_79 ();
 sg13g2_decap_4 FILLER_33_86 ();
 sg13g2_decap_4 FILLER_33_95 ();
 sg13g2_fill_1 FILLER_33_99 ();
 sg13g2_fill_2 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_107 ();
 sg13g2_decap_8 FILLER_33_153 ();
 sg13g2_decap_4 FILLER_33_160 ();
 sg13g2_fill_2 FILLER_33_164 ();
 sg13g2_decap_8 FILLER_33_170 ();
 sg13g2_decap_8 FILLER_33_212 ();
 sg13g2_fill_2 FILLER_33_219 ();
 sg13g2_fill_2 FILLER_33_224 ();
 sg13g2_fill_1 FILLER_33_226 ();
 sg13g2_fill_1 FILLER_33_233 ();
 sg13g2_decap_8 FILLER_33_249 ();
 sg13g2_decap_8 FILLER_33_256 ();
 sg13g2_fill_2 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_fill_2 FILLER_33_283 ();
 sg13g2_fill_1 FILLER_33_285 ();
 sg13g2_fill_2 FILLER_33_296 ();
 sg13g2_fill_1 FILLER_33_298 ();
 sg13g2_fill_2 FILLER_33_304 ();
 sg13g2_fill_2 FILLER_33_336 ();
 sg13g2_fill_1 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_391 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_33_415 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_fill_1 FILLER_34_10 ();
 sg13g2_decap_8 FILLER_34_45 ();
 sg13g2_fill_2 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_58 ();
 sg13g2_decap_4 FILLER_34_95 ();
 sg13g2_fill_1 FILLER_34_99 ();
 sg13g2_fill_2 FILLER_34_104 ();
 sg13g2_fill_1 FILLER_34_106 ();
 sg13g2_fill_1 FILLER_34_115 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_decap_8 FILLER_34_151 ();
 sg13g2_decap_8 FILLER_34_158 ();
 sg13g2_fill_2 FILLER_34_222 ();
 sg13g2_fill_1 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_228 ();
 sg13g2_fill_1 FILLER_34_230 ();
 sg13g2_fill_1 FILLER_34_257 ();
 sg13g2_fill_2 FILLER_34_263 ();
 sg13g2_fill_1 FILLER_34_269 ();
 sg13g2_fill_2 FILLER_34_274 ();
 sg13g2_fill_1 FILLER_34_276 ();
 sg13g2_decap_8 FILLER_34_311 ();
 sg13g2_decap_8 FILLER_34_318 ();
 sg13g2_decap_8 FILLER_34_325 ();
 sg13g2_decap_8 FILLER_34_332 ();
 sg13g2_fill_2 FILLER_34_339 ();
 sg13g2_fill_1 FILLER_34_341 ();
 sg13g2_fill_2 FILLER_34_368 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_11 ();
 sg13g2_decap_8 FILLER_35_52 ();
 sg13g2_decap_8 FILLER_35_59 ();
 sg13g2_decap_8 FILLER_35_66 ();
 sg13g2_decap_8 FILLER_35_73 ();
 sg13g2_decap_4 FILLER_35_80 ();
 sg13g2_decap_4 FILLER_35_110 ();
 sg13g2_decap_4 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_179 ();
 sg13g2_decap_4 FILLER_35_186 ();
 sg13g2_fill_2 FILLER_35_190 ();
 sg13g2_decap_8 FILLER_35_205 ();
 sg13g2_decap_4 FILLER_35_212 ();
 sg13g2_fill_1 FILLER_35_216 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_fill_2 FILLER_35_234 ();
 sg13g2_fill_1 FILLER_35_236 ();
 sg13g2_fill_2 FILLER_35_241 ();
 sg13g2_fill_1 FILLER_35_243 ();
 sg13g2_fill_2 FILLER_35_252 ();
 sg13g2_fill_1 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_268 ();
 sg13g2_fill_2 FILLER_35_278 ();
 sg13g2_fill_2 FILLER_35_290 ();
 sg13g2_fill_2 FILLER_35_331 ();
 sg13g2_fill_1 FILLER_35_333 ();
 sg13g2_fill_2 FILLER_35_343 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_358 ();
 sg13g2_decap_4 FILLER_35_386 ();
 sg13g2_fill_2 FILLER_35_390 ();
 sg13g2_decap_4 FILLER_35_400 ();
 sg13g2_decap_4 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_35_420 ();
 sg13g2_fill_2 FILLER_35_427 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_2 ();
 sg13g2_decap_4 FILLER_36_23 ();
 sg13g2_fill_2 FILLER_36_27 ();
 sg13g2_decap_4 FILLER_36_69 ();
 sg13g2_fill_1 FILLER_36_73 ();
 sg13g2_fill_1 FILLER_36_113 ();
 sg13g2_decap_8 FILLER_36_124 ();
 sg13g2_fill_2 FILLER_36_131 ();
 sg13g2_fill_2 FILLER_36_187 ();
 sg13g2_fill_2 FILLER_36_194 ();
 sg13g2_fill_1 FILLER_36_196 ();
 sg13g2_fill_1 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_229 ();
 sg13g2_fill_1 FILLER_36_237 ();
 sg13g2_fill_1 FILLER_36_259 ();
 sg13g2_fill_2 FILLER_36_282 ();
 sg13g2_fill_1 FILLER_36_284 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_fill_1 FILLER_36_350 ();
 sg13g2_fill_2 FILLER_36_381 ();
 sg13g2_fill_1 FILLER_36_383 ();
 sg13g2_fill_2 FILLER_36_392 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_38 ();
 sg13g2_fill_1 FILLER_37_45 ();
 sg13g2_decap_4 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_fill_1 FILLER_37_108 ();
 sg13g2_fill_2 FILLER_37_139 ();
 sg13g2_decap_4 FILLER_37_167 ();
 sg13g2_fill_2 FILLER_37_171 ();
 sg13g2_decap_4 FILLER_37_177 ();
 sg13g2_decap_4 FILLER_37_185 ();
 sg13g2_fill_2 FILLER_37_197 ();
 sg13g2_fill_1 FILLER_37_203 ();
 sg13g2_fill_1 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_fill_1 FILLER_37_240 ();
 sg13g2_fill_2 FILLER_37_264 ();
 sg13g2_fill_1 FILLER_37_286 ();
 sg13g2_fill_2 FILLER_37_297 ();
 sg13g2_fill_2 FILLER_37_353 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_fill_1 FILLER_37_379 ();
 sg13g2_fill_1 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_416 ();
 sg13g2_fill_2 FILLER_37_422 ();
 sg13g2_fill_2 FILLER_37_428 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_4 FILLER_38_61 ();
 sg13g2_fill_1 FILLER_38_109 ();
 sg13g2_fill_1 FILLER_38_114 ();
 sg13g2_fill_2 FILLER_38_209 ();
 sg13g2_fill_1 FILLER_38_293 ();
 sg13g2_decap_8 FILLER_38_320 ();
 sg13g2_fill_2 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_334 ();
 sg13g2_decap_8 FILLER_38_341 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_fill_1 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_fill_1 FILLER_38_429 ();
endmodule
